module basic_3000_30000_3500_6_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_2294,In_672);
nor U1 (N_1,In_866,In_336);
nor U2 (N_2,In_1820,In_2465);
or U3 (N_3,In_1020,In_2277);
nor U4 (N_4,In_353,In_951);
nand U5 (N_5,In_948,In_2934);
or U6 (N_6,In_2303,In_1817);
or U7 (N_7,In_1093,In_2125);
or U8 (N_8,In_1750,In_2314);
or U9 (N_9,In_2564,In_2760);
nor U10 (N_10,In_1454,In_1071);
or U11 (N_11,In_2598,In_2814);
and U12 (N_12,In_2223,In_488);
or U13 (N_13,In_2468,In_2791);
or U14 (N_14,In_1525,In_1213);
nor U15 (N_15,In_586,In_1881);
nand U16 (N_16,In_182,In_2280);
xnor U17 (N_17,In_388,In_2501);
nor U18 (N_18,In_2964,In_1884);
nand U19 (N_19,In_403,In_275);
xor U20 (N_20,In_2696,In_2843);
or U21 (N_21,In_1047,In_2706);
and U22 (N_22,In_2785,In_1401);
or U23 (N_23,In_1963,In_1479);
or U24 (N_24,In_215,In_663);
and U25 (N_25,In_533,In_1159);
and U26 (N_26,In_2879,In_2080);
xnor U27 (N_27,In_1938,In_2110);
or U28 (N_28,In_2678,In_2493);
or U29 (N_29,In_1393,In_1860);
and U30 (N_30,In_2630,In_1675);
and U31 (N_31,In_2351,In_2903);
or U32 (N_32,In_794,In_2744);
nor U33 (N_33,In_2768,In_2010);
nor U34 (N_34,In_2723,In_1925);
nand U35 (N_35,In_1802,In_1024);
and U36 (N_36,In_2543,In_1420);
and U37 (N_37,In_2460,In_933);
nand U38 (N_38,In_919,In_1599);
or U39 (N_39,In_486,In_621);
nor U40 (N_40,In_334,In_1759);
xnor U41 (N_41,In_1697,In_2137);
and U42 (N_42,In_1859,In_382);
or U43 (N_43,In_818,In_1873);
nor U44 (N_44,In_138,In_1235);
nor U45 (N_45,In_993,In_1439);
or U46 (N_46,In_2755,In_851);
and U47 (N_47,In_543,In_1927);
xnor U48 (N_48,In_1397,In_2360);
or U49 (N_49,In_2166,In_1257);
xnor U50 (N_50,In_2756,In_240);
or U51 (N_51,In_2956,In_1296);
nor U52 (N_52,In_654,In_1359);
xnor U53 (N_53,In_149,In_131);
nor U54 (N_54,In_986,In_1382);
and U55 (N_55,In_1299,In_2611);
nor U56 (N_56,In_1219,In_1617);
nor U57 (N_57,In_250,In_2919);
nand U58 (N_58,In_27,In_791);
or U59 (N_59,In_2936,In_1051);
and U60 (N_60,In_222,In_1017);
and U61 (N_61,In_517,In_1991);
and U62 (N_62,In_1433,In_1696);
or U63 (N_63,In_2368,In_2121);
nor U64 (N_64,In_2429,In_1847);
xor U65 (N_65,In_1259,In_764);
nand U66 (N_66,In_2372,In_1554);
and U67 (N_67,In_1288,In_2712);
and U68 (N_68,In_2235,In_479);
and U69 (N_69,In_831,In_116);
xnor U70 (N_70,In_2373,In_1946);
or U71 (N_71,In_9,In_386);
nor U72 (N_72,In_2567,In_1958);
or U73 (N_73,In_1669,In_2011);
xnor U74 (N_74,In_2306,In_566);
and U75 (N_75,In_104,In_2152);
nor U76 (N_76,In_1425,In_1521);
nor U77 (N_77,In_1123,In_883);
nand U78 (N_78,In_2423,In_180);
and U79 (N_79,In_2848,In_1004);
and U80 (N_80,In_2838,In_963);
and U81 (N_81,In_2927,In_2688);
nor U82 (N_82,In_2247,In_1854);
nor U83 (N_83,In_692,In_1723);
nand U84 (N_84,In_970,In_610);
or U85 (N_85,In_2150,In_1740);
or U86 (N_86,In_1006,In_1297);
and U87 (N_87,In_1830,In_2859);
nor U88 (N_88,In_436,In_2466);
nand U89 (N_89,In_2911,In_541);
xnor U90 (N_90,In_296,In_519);
and U91 (N_91,In_2194,In_786);
nand U92 (N_92,In_1849,In_2731);
and U93 (N_93,In_1780,In_1527);
or U94 (N_94,In_2279,In_530);
nor U95 (N_95,In_1418,In_1000);
or U96 (N_96,In_584,In_669);
nand U97 (N_97,In_1950,In_318);
or U98 (N_98,In_591,In_2681);
nor U99 (N_99,In_2232,In_1320);
xnor U100 (N_100,In_161,In_2617);
and U101 (N_101,In_1325,In_345);
or U102 (N_102,In_920,In_2989);
nand U103 (N_103,In_1409,In_1920);
or U104 (N_104,In_376,In_930);
and U105 (N_105,In_463,In_617);
nand U106 (N_106,In_996,In_2535);
or U107 (N_107,In_1404,In_1346);
xor U108 (N_108,In_2063,In_1277);
and U109 (N_109,In_2789,In_1825);
nand U110 (N_110,In_2658,In_2478);
nor U111 (N_111,In_2335,In_2728);
nor U112 (N_112,In_2652,In_226);
and U113 (N_113,In_2537,In_2325);
nand U114 (N_114,In_15,In_915);
xnor U115 (N_115,In_999,In_1548);
or U116 (N_116,In_1162,In_1821);
or U117 (N_117,In_2812,In_1836);
or U118 (N_118,In_2578,In_1310);
or U119 (N_119,In_2454,In_1887);
nand U120 (N_120,In_1134,In_384);
nor U121 (N_121,In_2308,In_2776);
xnor U122 (N_122,In_1270,In_1236);
and U123 (N_123,In_761,In_1304);
nand U124 (N_124,In_1465,In_629);
nor U125 (N_125,In_482,In_2356);
nor U126 (N_126,In_1505,In_1423);
nand U127 (N_127,In_1200,In_1339);
xnor U128 (N_128,In_534,In_2973);
xnor U129 (N_129,In_1130,In_832);
nor U130 (N_130,In_767,In_735);
nor U131 (N_131,In_1922,In_619);
and U132 (N_132,In_1399,In_2562);
nor U133 (N_133,In_1755,In_2419);
or U134 (N_134,In_2014,In_1);
nor U135 (N_135,In_1536,In_2620);
and U136 (N_136,In_2614,In_2746);
xor U137 (N_137,In_10,In_2691);
nor U138 (N_138,In_220,In_2437);
nor U139 (N_139,In_2604,In_2340);
or U140 (N_140,In_755,In_1440);
nand U141 (N_141,In_2718,In_1009);
nor U142 (N_142,In_532,In_2969);
and U143 (N_143,In_448,In_2778);
nand U144 (N_144,In_1874,In_2425);
and U145 (N_145,In_1819,In_2023);
nand U146 (N_146,In_2570,In_772);
nand U147 (N_147,In_233,In_415);
or U148 (N_148,In_724,In_58);
xor U149 (N_149,In_2684,In_2054);
and U150 (N_150,In_242,In_19);
nand U151 (N_151,In_773,In_1862);
and U152 (N_152,In_1165,In_1208);
xnor U153 (N_153,In_1010,In_2378);
nand U154 (N_154,In_606,In_1263);
nor U155 (N_155,In_1625,In_274);
and U156 (N_156,In_356,In_2975);
or U157 (N_157,In_1774,In_184);
or U158 (N_158,In_814,In_905);
nor U159 (N_159,In_2645,In_2055);
or U160 (N_160,In_2820,In_1302);
and U161 (N_161,In_1402,In_151);
and U162 (N_162,In_1983,In_2855);
nor U163 (N_163,In_754,In_314);
nor U164 (N_164,In_327,In_1701);
nor U165 (N_165,In_738,In_727);
and U166 (N_166,In_351,In_864);
nor U167 (N_167,In_2742,In_2762);
nand U168 (N_168,In_1704,In_521);
or U169 (N_169,In_2153,In_1065);
or U170 (N_170,In_2628,In_1980);
nand U171 (N_171,In_2822,In_763);
nor U172 (N_172,In_1113,In_784);
nand U173 (N_173,In_759,In_1545);
xnor U174 (N_174,In_542,In_1201);
nand U175 (N_175,In_1804,In_1223);
xor U176 (N_176,In_2680,In_2738);
and U177 (N_177,In_2026,In_2496);
or U178 (N_178,In_2866,In_1923);
and U179 (N_179,In_1658,In_2845);
or U180 (N_180,In_932,In_304);
xnor U181 (N_181,In_676,In_1467);
and U182 (N_182,In_1550,In_561);
or U183 (N_183,In_2574,In_1108);
and U184 (N_184,In_941,In_1636);
nor U185 (N_185,In_290,In_1491);
nor U186 (N_186,In_1823,In_715);
and U187 (N_187,In_1031,In_526);
nor U188 (N_188,In_1516,In_2986);
nand U189 (N_189,In_2271,In_1916);
and U190 (N_190,In_2606,In_2787);
or U191 (N_191,In_1543,In_217);
or U192 (N_192,In_827,In_983);
and U193 (N_193,In_1224,In_1097);
and U194 (N_194,In_2109,In_651);
and U195 (N_195,In_697,In_1842);
nor U196 (N_196,In_2082,In_469);
nor U197 (N_197,In_1040,In_2829);
and U198 (N_198,In_769,In_1736);
or U199 (N_199,In_1171,In_656);
xor U200 (N_200,In_1987,In_1993);
or U201 (N_201,In_1023,In_2093);
or U202 (N_202,In_241,In_859);
or U203 (N_203,In_1688,In_782);
and U204 (N_204,In_2181,In_554);
xor U205 (N_205,In_1081,In_1630);
or U206 (N_206,In_1225,In_2490);
and U207 (N_207,In_2477,In_123);
nand U208 (N_208,In_2920,In_1044);
nor U209 (N_209,In_2346,In_1622);
nor U210 (N_210,In_234,In_344);
nand U211 (N_211,In_473,In_2726);
xnor U212 (N_212,In_2128,In_1385);
or U213 (N_213,In_2753,In_2329);
nor U214 (N_214,In_1511,In_2725);
nand U215 (N_215,In_648,In_107);
or U216 (N_216,In_2263,In_802);
nand U217 (N_217,In_2521,In_1947);
or U218 (N_218,In_1074,In_1955);
nor U219 (N_219,In_229,In_2893);
or U220 (N_220,In_1260,In_1187);
xor U221 (N_221,In_631,In_1099);
and U222 (N_222,In_1561,In_2650);
and U223 (N_223,In_1114,In_1341);
xor U224 (N_224,In_1915,In_496);
and U225 (N_225,In_823,In_103);
or U226 (N_226,In_2268,In_2724);
nor U227 (N_227,In_1727,In_2944);
and U228 (N_228,In_1809,In_173);
nor U229 (N_229,In_2951,In_740);
nand U230 (N_230,In_1744,In_1939);
or U231 (N_231,In_1076,In_1067);
and U232 (N_232,In_1475,In_730);
nor U233 (N_233,In_1487,In_349);
and U234 (N_234,In_585,In_2663);
xor U235 (N_235,In_882,In_689);
nand U236 (N_236,In_1365,In_1091);
nor U237 (N_237,In_1142,In_1757);
nand U238 (N_238,In_926,In_1309);
and U239 (N_239,In_1743,In_2230);
and U240 (N_240,In_1756,In_276);
nor U241 (N_241,In_2516,In_1117);
nor U242 (N_242,In_537,In_2143);
nor U243 (N_243,In_2160,In_2615);
or U244 (N_244,In_2510,In_87);
and U245 (N_245,In_2997,In_1753);
nand U246 (N_246,In_1292,In_1853);
or U247 (N_247,In_929,In_2795);
or U248 (N_248,In_1871,In_1066);
nand U249 (N_249,In_671,In_2215);
nor U250 (N_250,In_855,In_475);
and U251 (N_251,In_1883,In_342);
nand U252 (N_252,In_1893,In_1607);
and U253 (N_253,In_2906,In_465);
and U254 (N_254,In_310,In_602);
xnor U255 (N_255,In_1770,In_2900);
xor U256 (N_256,In_981,In_1678);
and U257 (N_257,In_1992,In_1553);
nor U258 (N_258,In_175,In_643);
or U259 (N_259,In_1778,In_2884);
nor U260 (N_260,In_780,In_1459);
nand U261 (N_261,In_305,In_801);
nand U262 (N_262,In_1900,In_474);
and U263 (N_263,In_1090,In_574);
nand U264 (N_264,In_2441,In_657);
nand U265 (N_265,In_748,In_547);
nor U266 (N_266,In_2074,In_223);
nand U267 (N_267,In_1226,In_1775);
and U268 (N_268,In_1438,In_80);
nor U269 (N_269,In_2933,In_1929);
nor U270 (N_270,In_1713,In_1319);
nand U271 (N_271,In_102,In_257);
or U272 (N_272,In_467,In_940);
xnor U273 (N_273,In_393,In_2081);
nor U274 (N_274,In_2909,In_355);
nand U275 (N_275,In_942,In_1073);
xnor U276 (N_276,In_1652,In_2371);
nor U277 (N_277,In_1338,In_2896);
nand U278 (N_278,In_2719,In_1986);
nor U279 (N_279,In_1068,In_1250);
nand U280 (N_280,In_1711,In_361);
nor U281 (N_281,In_2307,In_427);
nand U282 (N_282,In_1904,In_2509);
or U283 (N_283,In_1928,In_725);
and U284 (N_284,In_1656,In_2261);
and U285 (N_285,In_1141,In_52);
nor U286 (N_286,In_1665,In_1406);
xor U287 (N_287,In_2069,In_2366);
or U288 (N_288,In_2267,In_641);
or U289 (N_289,In_2375,In_2355);
and U290 (N_290,In_2018,In_758);
nor U291 (N_291,In_272,In_1764);
nand U292 (N_292,In_2282,In_61);
and U293 (N_293,In_2624,In_2332);
and U294 (N_294,In_1272,In_1643);
or U295 (N_295,In_1212,In_2524);
nand U296 (N_296,In_2456,In_1025);
nor U297 (N_297,In_2002,In_760);
nor U298 (N_298,In_1832,In_1841);
xnor U299 (N_299,In_634,In_573);
or U300 (N_300,In_251,In_2698);
nand U301 (N_301,In_916,In_1481);
nand U302 (N_302,In_2849,In_1934);
xor U303 (N_303,In_1390,In_1243);
xor U304 (N_304,In_298,In_380);
nor U305 (N_305,In_2387,In_68);
nor U306 (N_306,In_1412,In_1840);
and U307 (N_307,In_273,In_1542);
and U308 (N_308,In_279,In_1258);
nor U309 (N_309,In_209,In_1677);
xor U310 (N_310,In_1644,In_2212);
nand U311 (N_311,In_2583,In_563);
nand U312 (N_312,In_1450,In_2326);
nand U313 (N_313,In_1602,In_164);
or U314 (N_314,In_246,In_2891);
or U315 (N_315,In_901,In_331);
and U316 (N_316,In_2291,In_675);
nor U317 (N_317,In_2702,In_2968);
or U318 (N_318,In_330,In_409);
or U319 (N_319,In_419,In_795);
nand U320 (N_320,In_421,In_2670);
nand U321 (N_321,In_79,In_200);
nor U322 (N_322,In_2508,In_2185);
nand U323 (N_323,In_159,In_53);
or U324 (N_324,In_2112,In_1662);
and U325 (N_325,In_876,In_659);
and U326 (N_326,In_143,In_745);
nand U327 (N_327,In_2971,In_1549);
nor U328 (N_328,In_987,In_1174);
or U329 (N_329,In_1957,In_2358);
nand U330 (N_330,In_1869,In_2021);
and U331 (N_331,In_191,In_1591);
or U332 (N_332,In_1612,In_807);
nor U333 (N_333,In_1518,In_1910);
nor U334 (N_334,In_976,In_1571);
nor U335 (N_335,In_127,In_2489);
nand U336 (N_336,In_2184,In_881);
or U337 (N_337,In_798,In_1924);
nor U338 (N_338,In_841,In_1728);
nand U339 (N_339,In_278,In_1970);
nor U340 (N_340,In_2586,In_2293);
and U341 (N_341,In_452,In_31);
and U342 (N_342,In_1034,In_1973);
or U343 (N_343,In_1749,In_214);
and U344 (N_344,In_364,In_2974);
nand U345 (N_345,In_958,In_1715);
nand U346 (N_346,In_2107,In_2283);
or U347 (N_347,In_1218,In_2357);
or U348 (N_348,In_1654,In_2272);
or U349 (N_349,In_1541,In_1158);
or U350 (N_350,In_1801,In_2210);
nand U351 (N_351,In_156,In_1038);
nand U352 (N_352,In_1524,In_694);
or U353 (N_353,In_1912,In_950);
and U354 (N_354,In_548,In_826);
nor U355 (N_355,In_379,In_890);
or U356 (N_356,In_1800,In_1761);
or U357 (N_357,In_2816,In_871);
nor U358 (N_358,In_2948,In_2205);
or U359 (N_359,In_1335,In_460);
nor U360 (N_360,In_1328,In_2794);
or U361 (N_361,In_1805,In_2047);
or U362 (N_362,In_2459,In_1803);
or U363 (N_363,In_2139,In_2027);
nor U364 (N_364,In_1741,In_1507);
and U365 (N_365,In_1814,In_295);
nand U366 (N_366,In_1054,In_618);
nand U367 (N_367,In_28,In_1633);
nand U368 (N_368,In_2888,In_2344);
and U369 (N_369,In_450,In_1110);
nand U370 (N_370,In_471,In_2146);
or U371 (N_371,In_1348,In_89);
or U372 (N_372,In_2648,In_712);
nor U373 (N_373,In_653,In_1428);
nand U374 (N_374,In_2452,In_1349);
or U375 (N_375,In_1316,In_1529);
and U376 (N_376,In_2539,In_374);
nand U377 (N_377,In_2122,In_1313);
nand U378 (N_378,In_1911,In_1026);
and U379 (N_379,In_2260,In_1173);
nor U380 (N_380,In_2905,In_1735);
nor U381 (N_381,In_2061,In_900);
and U382 (N_382,In_1135,In_1264);
nor U383 (N_383,In_1868,In_2597);
and U384 (N_384,In_1818,In_360);
and U385 (N_385,In_1289,In_1028);
or U386 (N_386,In_2046,In_2037);
nand U387 (N_387,In_2671,In_2033);
nand U388 (N_388,In_2379,In_2013);
xor U389 (N_389,In_135,In_194);
xor U390 (N_390,In_137,In_1886);
nand U391 (N_391,In_2310,In_2156);
or U392 (N_392,In_2130,In_462);
nor U393 (N_393,In_1584,In_1522);
xor U394 (N_394,In_1532,In_2799);
nor U395 (N_395,In_1345,In_778);
or U396 (N_396,In_2542,In_25);
nor U397 (N_397,In_2715,In_1945);
nand U398 (N_398,In_1011,In_1210);
nor U399 (N_399,In_181,In_1935);
xor U400 (N_400,In_2882,In_1391);
xor U401 (N_401,In_1844,In_2781);
nor U402 (N_402,In_190,In_1298);
and U403 (N_403,In_2077,In_1777);
nand U404 (N_404,In_2792,In_2409);
nand U405 (N_405,In_637,In_1072);
and U406 (N_406,In_2970,In_549);
nand U407 (N_407,In_601,In_1358);
and U408 (N_408,In_1870,In_64);
nor U409 (N_409,In_1228,In_2320);
and U410 (N_410,In_690,In_1087);
and U411 (N_411,In_2221,In_2175);
xnor U412 (N_412,In_1661,In_1285);
nor U413 (N_413,In_2402,In_1480);
nand U414 (N_414,In_2674,In_368);
or U415 (N_415,In_2603,In_2017);
or U416 (N_416,In_2050,In_1793);
or U417 (N_417,In_381,In_2644);
nand U418 (N_418,In_1514,In_2505);
nand U419 (N_419,In_2083,In_1866);
nor U420 (N_420,In_2149,In_2031);
nor U421 (N_421,In_308,In_2533);
nand U422 (N_422,In_2334,In_1300);
or U423 (N_423,In_811,In_2939);
and U424 (N_424,In_2921,In_1729);
nand U425 (N_425,In_1621,In_2589);
and U426 (N_426,In_1948,In_2231);
nand U427 (N_427,In_765,In_2228);
xor U428 (N_428,In_2370,In_146);
and U429 (N_429,In_2549,In_2312);
nand U430 (N_430,In_1673,In_2337);
nor U431 (N_431,In_1052,In_1687);
nand U432 (N_432,In_2904,In_984);
xor U433 (N_433,In_2883,In_2552);
and U434 (N_434,In_2827,In_749);
nand U435 (N_435,In_283,In_545);
nor U436 (N_436,In_2197,In_1271);
nor U437 (N_437,In_105,In_598);
or U438 (N_438,In_418,In_702);
or U439 (N_439,In_2581,In_650);
xor U440 (N_440,In_626,In_2016);
nand U441 (N_441,In_168,In_2127);
and U442 (N_442,In_433,In_2869);
and U443 (N_443,In_1537,In_396);
or U444 (N_444,In_1387,In_887);
nor U445 (N_445,In_846,In_2457);
or U446 (N_446,In_370,In_134);
nand U447 (N_447,In_48,In_2824);
or U448 (N_448,In_1918,In_605);
nor U449 (N_449,In_998,In_1730);
nor U450 (N_450,In_1693,In_2867);
xnor U451 (N_451,In_1850,In_2446);
nand U452 (N_452,In_2625,In_1610);
or U453 (N_453,In_2138,In_2514);
or U454 (N_454,In_503,In_2873);
xor U455 (N_455,In_2548,In_1301);
and U456 (N_456,In_1482,In_2251);
and U457 (N_457,In_1494,In_1655);
nand U458 (N_458,In_2204,In_316);
or U459 (N_459,In_2323,In_1593);
and U460 (N_460,In_301,In_18);
nand U461 (N_461,In_29,In_443);
nor U462 (N_462,In_2853,In_2965);
nand U463 (N_463,In_964,In_484);
nand U464 (N_464,In_969,In_2155);
or U465 (N_465,In_1937,In_1831);
and U466 (N_466,In_2856,In_91);
xnor U467 (N_467,In_248,In_2546);
and U468 (N_468,In_338,In_2664);
or U469 (N_469,In_806,In_1510);
or U470 (N_470,In_2714,In_198);
and U471 (N_471,In_115,In_1177);
nand U472 (N_472,In_1523,In_1352);
nor U473 (N_473,In_167,In_445);
nand U474 (N_474,In_2498,In_646);
or U475 (N_475,In_302,In_2404);
nand U476 (N_476,In_511,In_2158);
nand U477 (N_477,In_2512,In_444);
xnor U478 (N_478,In_1460,In_1811);
nor U479 (N_479,In_2745,In_645);
or U480 (N_480,In_346,In_1186);
or U481 (N_481,In_717,In_2651);
nor U482 (N_482,In_1045,In_157);
or U483 (N_483,In_2550,In_2704);
xnor U484 (N_484,In_1990,In_1417);
nand U485 (N_485,In_323,In_2841);
or U486 (N_486,In_2995,In_106);
nand U487 (N_487,In_0,In_824);
nor U488 (N_488,In_119,In_428);
nor U489 (N_489,In_2020,In_2438);
or U490 (N_490,In_670,In_2519);
and U491 (N_491,In_26,In_1430);
or U492 (N_492,In_2295,In_39);
nor U493 (N_493,In_2248,In_2421);
nand U494 (N_494,In_1620,In_945);
xnor U495 (N_495,In_1379,In_2608);
xor U496 (N_496,In_1679,In_1104);
nand U497 (N_497,In_819,In_432);
nand U498 (N_498,In_2411,In_124);
and U499 (N_499,In_2953,In_1217);
xnor U500 (N_500,In_2266,In_2507);
or U501 (N_501,In_1503,In_263);
nor U502 (N_502,In_1734,In_2709);
nor U503 (N_503,In_111,In_2610);
nor U504 (N_504,In_513,In_678);
and U505 (N_505,In_2835,In_238);
nor U506 (N_506,In_2183,In_1092);
nand U507 (N_507,In_320,In_700);
nor U508 (N_508,In_2802,In_2207);
nand U509 (N_509,In_369,In_485);
nand U510 (N_510,In_2476,In_2443);
nor U511 (N_511,In_122,In_2214);
and U512 (N_512,In_2865,In_781);
nor U513 (N_513,In_2328,In_1603);
nand U514 (N_514,In_1196,In_2765);
nor U515 (N_515,In_1776,In_2763);
nand U516 (N_516,In_1834,In_2863);
and U517 (N_517,In_2428,In_478);
nand U518 (N_518,In_322,In_1905);
nor U519 (N_519,In_2612,In_294);
nand U520 (N_520,In_1360,In_2798);
nand U521 (N_521,In_2559,In_1999);
and U522 (N_522,In_2417,In_2068);
xnor U523 (N_523,In_2043,In_2176);
or U524 (N_524,In_1977,In_1616);
nand U525 (N_525,In_363,In_321);
or U526 (N_526,In_1180,In_1105);
or U527 (N_527,In_2902,In_550);
and U528 (N_528,In_2631,In_1576);
nor U529 (N_529,In_1237,In_2474);
nor U530 (N_530,In_1155,In_2233);
or U531 (N_531,In_1016,In_1663);
or U532 (N_532,In_1798,In_162);
and U533 (N_533,In_2032,In_982);
nand U534 (N_534,In_422,In_101);
and U535 (N_535,In_2898,In_258);
nand U536 (N_536,In_2079,In_129);
nand U537 (N_537,In_1455,In_1242);
nand U538 (N_538,In_1362,In_2318);
and U539 (N_539,In_844,In_437);
xnor U540 (N_540,In_2376,In_2761);
nand U541 (N_541,In_2195,In_1628);
nor U542 (N_542,In_1880,In_611);
nand U543 (N_543,In_737,In_512);
and U544 (N_544,In_2433,In_303);
and U545 (N_545,In_2024,In_2871);
and U546 (N_546,In_1221,In_2052);
nand U547 (N_547,In_37,In_2561);
or U548 (N_548,In_1253,In_1227);
nor U549 (N_549,In_721,In_680);
nand U550 (N_550,In_2942,In_414);
or U551 (N_551,In_2912,In_1552);
and U552 (N_552,In_2692,In_1458);
and U553 (N_553,In_2632,In_1317);
and U554 (N_554,In_1485,In_329);
or U555 (N_555,In_252,In_2639);
or U556 (N_556,In_2613,In_1446);
nand U557 (N_557,In_397,In_2804);
nand U558 (N_558,In_291,In_718);
and U559 (N_559,In_1116,In_2525);
and U560 (N_560,In_2062,In_1120);
nand U561 (N_561,In_85,In_97);
nor U562 (N_562,In_935,In_2929);
and U563 (N_563,In_1468,In_518);
xor U564 (N_564,In_2599,In_2359);
nor U565 (N_565,In_693,In_1931);
nand U566 (N_566,In_2317,In_140);
xnor U567 (N_567,In_2420,In_2000);
or U568 (N_568,In_328,In_228);
nor U569 (N_569,In_1055,In_2398);
and U570 (N_570,In_2713,In_171);
and U571 (N_571,In_268,In_2952);
xor U572 (N_572,In_98,In_2432);
or U573 (N_573,In_1233,In_716);
nor U574 (N_574,In_2264,In_1828);
nand U575 (N_575,In_1036,In_2497);
nand U576 (N_576,In_2287,In_1861);
or U577 (N_577,In_1206,In_2622);
nand U578 (N_578,In_2649,In_1626);
and U579 (N_579,In_896,In_2740);
nand U580 (N_580,In_1432,In_1540);
xnor U581 (N_581,In_466,In_42);
xnor U582 (N_582,In_2281,In_1416);
and U583 (N_583,In_1472,In_2817);
or U584 (N_584,In_365,In_1824);
and U585 (N_585,In_2805,In_72);
nand U586 (N_586,In_2163,In_2515);
nand U587 (N_587,In_1855,In_1167);
xnor U588 (N_588,In_756,In_2837);
nand U589 (N_589,In_1079,In_2730);
or U590 (N_590,In_885,In_1053);
nand U591 (N_591,In_166,In_1153);
nand U592 (N_592,In_2687,In_685);
or U593 (N_593,In_1118,In_509);
and U594 (N_594,In_1737,In_785);
nor U595 (N_595,In_1965,In_2994);
xnor U596 (N_596,In_753,In_803);
or U597 (N_597,In_158,In_74);
nor U598 (N_598,In_2101,In_2788);
xnor U599 (N_599,In_2142,In_2627);
nor U600 (N_600,In_2012,In_489);
nand U601 (N_601,In_2145,In_1822);
nand U602 (N_602,In_614,In_2132);
nor U603 (N_603,In_1790,In_1515);
nor U604 (N_604,In_1722,In_2634);
and U605 (N_605,In_1563,In_994);
nand U606 (N_606,In_1720,In_2555);
nand U607 (N_607,In_1672,In_193);
nor U608 (N_608,In_1386,In_2573);
nand U609 (N_609,In_451,In_2757);
nand U610 (N_610,In_2447,In_2380);
and U611 (N_611,In_1995,In_2250);
or U612 (N_612,In_630,In_2665);
or U613 (N_613,In_1030,In_2923);
and U614 (N_614,In_1070,In_1839);
nor U615 (N_615,In_1484,In_747);
nor U616 (N_616,In_255,In_2470);
or U617 (N_617,In_1998,In_1107);
nor U618 (N_618,In_1502,In_1216);
or U619 (N_619,In_2526,In_95);
nor U620 (N_620,In_1660,In_1974);
nor U621 (N_621,In_1789,In_1451);
and U622 (N_622,In_615,In_572);
xnor U623 (N_623,In_1477,In_2252);
nand U624 (N_624,In_734,In_2162);
and U625 (N_625,In_1978,In_1666);
and U626 (N_626,In_2743,In_2662);
nor U627 (N_627,In_205,In_1029);
and U628 (N_628,In_434,In_1982);
or U629 (N_629,In_2100,In_1077);
or U630 (N_630,In_1415,In_2657);
nor U631 (N_631,In_1240,In_1083);
or U632 (N_632,In_358,In_949);
xor U633 (N_633,In_2168,In_2240);
nor U634 (N_634,In_873,In_2647);
or U635 (N_635,In_1291,In_1588);
or U636 (N_636,In_2414,In_16);
xor U637 (N_637,In_552,In_1520);
or U638 (N_638,In_22,In_2937);
and U639 (N_639,In_2741,In_581);
and U640 (N_640,In_2754,In_2315);
or U641 (N_641,In_284,In_1241);
nor U642 (N_642,In_793,In_49);
nor U643 (N_643,In_1222,In_1969);
and U644 (N_644,In_1373,In_212);
nor U645 (N_645,In_2553,In_347);
or U646 (N_646,In_593,In_865);
or U647 (N_647,In_628,In_1342);
nand U648 (N_648,In_306,In_2571);
or U649 (N_649,In_809,In_2721);
and U650 (N_650,In_1649,In_739);
and U651 (N_651,In_505,In_1064);
nand U652 (N_652,In_1632,In_902);
and U653 (N_653,In_2572,In_821);
or U654 (N_654,In_588,In_1572);
nor U655 (N_655,In_2300,In_77);
xnor U656 (N_656,In_2844,In_1500);
or U657 (N_657,In_2418,In_2557);
nor U658 (N_658,In_2273,In_51);
and U659 (N_659,In_2983,In_2872);
or U660 (N_660,In_1082,In_1333);
nand U661 (N_661,In_441,In_76);
nor U662 (N_662,In_1526,In_2198);
nor U663 (N_663,In_1203,In_1670);
nor U664 (N_664,In_2846,In_1337);
xor U665 (N_665,In_2659,In_1330);
nand U666 (N_666,In_1719,In_2473);
or U667 (N_667,In_232,In_2399);
and U668 (N_668,In_2367,In_2187);
or U669 (N_669,In_1702,In_966);
and U670 (N_670,In_943,In_55);
nor U671 (N_671,In_1245,In_2087);
or U672 (N_672,In_2288,In_1012);
xnor U673 (N_673,In_2106,In_2436);
and U674 (N_674,In_2769,In_1609);
nand U675 (N_675,In_2685,In_2880);
or U676 (N_676,In_577,In_906);
and U677 (N_677,In_2426,In_2290);
or U678 (N_678,In_2455,In_2259);
or U679 (N_679,In_1363,In_392);
nor U680 (N_680,In_2522,In_2779);
or U681 (N_681,In_493,In_2941);
nand U682 (N_682,In_2494,In_1131);
and U683 (N_683,In_627,In_2991);
nand U684 (N_684,In_1334,In_211);
xor U685 (N_685,In_2193,In_1027);
nand U686 (N_686,In_2299,In_2784);
and U687 (N_687,In_603,In_1078);
nor U688 (N_688,In_2528,In_1361);
nand U689 (N_689,In_93,In_1197);
nor U690 (N_690,In_1019,In_1686);
or U691 (N_691,In_2154,In_1340);
nand U692 (N_692,In_1567,In_1568);
nand U693 (N_693,In_708,In_589);
xnor U694 (N_694,In_2940,In_1914);
and U695 (N_695,In_1182,In_2895);
nand U696 (N_696,In_1642,In_2269);
or U697 (N_697,In_2479,In_20);
xor U698 (N_698,In_938,In_1569);
or U699 (N_699,In_1703,In_729);
or U700 (N_700,In_952,In_1369);
xnor U701 (N_701,In_2065,In_231);
and U702 (N_702,In_1555,In_1650);
nor U703 (N_703,In_2727,In_580);
nand U704 (N_704,In_2683,In_425);
nand U705 (N_705,In_1112,In_2737);
xor U706 (N_706,In_1647,In_647);
and U707 (N_707,In_2722,In_2416);
and U708 (N_708,In_1049,In_1700);
or U709 (N_709,In_2600,In_812);
or U710 (N_710,In_1255,In_751);
nor U711 (N_711,In_2808,In_2369);
or U712 (N_712,In_863,In_723);
nor U713 (N_713,In_1137,In_2556);
nor U714 (N_714,In_2405,In_487);
or U715 (N_715,In_1426,In_2499);
or U716 (N_716,In_2336,In_558);
and U717 (N_717,In_1464,In_1967);
nor U718 (N_718,In_1347,In_2103);
nand U719 (N_719,In_2926,In_2157);
and U720 (N_720,In_1042,In_1848);
nand U721 (N_721,In_1239,In_1493);
nor U722 (N_722,In_247,In_2029);
or U723 (N_723,In_1207,In_2487);
nor U724 (N_724,In_2462,In_2339);
nor U725 (N_725,In_208,In_2413);
or U726 (N_726,In_1558,In_2803);
or U727 (N_727,In_2852,In_560);
xor U728 (N_728,In_1976,In_185);
nand U729 (N_729,In_169,In_2042);
xor U730 (N_730,In_2915,In_2025);
nor U731 (N_731,In_564,In_221);
or U732 (N_732,In_774,In_2302);
nand U733 (N_733,In_2381,In_2464);
xnor U734 (N_734,In_858,In_886);
and U735 (N_735,In_1403,In_661);
and U736 (N_736,In_775,In_836);
nor U737 (N_737,In_894,In_1230);
xor U738 (N_738,In_2333,In_609);
and U739 (N_739,In_1303,In_2120);
nand U740 (N_740,In_2959,In_2220);
or U741 (N_741,In_2225,In_399);
or U742 (N_742,In_1752,In_1495);
and U743 (N_743,In_594,In_2495);
nand U744 (N_744,In_1985,In_1127);
nor U745 (N_745,In_1808,In_2609);
nand U746 (N_746,In_974,In_2733);
or U747 (N_747,In_707,In_2091);
nand U748 (N_748,In_2988,In_965);
nand U749 (N_749,In_2222,In_2059);
and U750 (N_750,In_1282,In_1530);
nor U751 (N_751,In_216,In_2253);
nor U752 (N_752,In_928,In_1128);
xnor U753 (N_753,In_108,In_1232);
and U754 (N_754,In_2635,In_677);
or U755 (N_755,In_575,In_559);
and U756 (N_756,In_1872,In_1681);
xor U757 (N_757,In_2582,In_691);
and U758 (N_758,In_424,In_2602);
nand U759 (N_759,In_828,In_1721);
and U760 (N_760,In_1022,In_2345);
nor U761 (N_761,In_5,In_2985);
nand U762 (N_762,In_458,In_2219);
nor U763 (N_763,In_925,In_69);
and U764 (N_764,In_2580,In_1926);
nor U765 (N_765,In_1007,In_536);
nor U766 (N_766,In_2397,In_1634);
and U767 (N_767,In_1144,In_1598);
nor U768 (N_768,In_2887,In_2238);
nand U769 (N_769,In_1574,In_1132);
and U770 (N_770,In_662,In_2945);
and U771 (N_771,In_917,In_1807);
nand U772 (N_772,In_1897,In_2412);
or U773 (N_773,In_1714,In_1096);
and U774 (N_774,In_2851,In_2710);
or U775 (N_775,In_2056,In_1471);
and U776 (N_776,In_402,In_1246);
or U777 (N_777,In_1806,In_1953);
or U778 (N_778,In_2506,In_389);
nor U779 (N_779,In_666,In_1682);
nand U780 (N_780,In_14,In_848);
xor U781 (N_781,In_907,In_1149);
or U782 (N_782,In_546,In_847);
nor U783 (N_783,In_1577,In_2390);
nor U784 (N_784,In_1857,In_2917);
xor U785 (N_785,In_1898,In_332);
or U786 (N_786,In_1538,In_2908);
nor U787 (N_787,In_132,In_2642);
or U788 (N_788,In_612,In_1816);
nor U789 (N_789,In_1294,In_2842);
nand U790 (N_790,In_1899,In_842);
and U791 (N_791,In_528,In_2924);
or U792 (N_792,In_679,In_1546);
or U793 (N_793,In_544,In_1792);
nand U794 (N_794,In_2258,In_1276);
nand U795 (N_795,In_120,In_766);
nand U796 (N_796,In_2672,In_1244);
nand U797 (N_797,In_1395,In_75);
or U798 (N_798,In_2513,In_2200);
or U799 (N_799,In_352,In_1344);
nand U800 (N_800,In_623,In_1095);
nor U801 (N_801,In_2191,In_2861);
nor U802 (N_802,In_2773,In_1278);
xor U803 (N_803,In_771,In_1452);
and U804 (N_804,In_1229,In_2485);
xnor U805 (N_805,In_2111,In_2044);
nand U806 (N_806,In_219,In_1930);
or U807 (N_807,In_54,In_1706);
or U808 (N_808,In_682,In_2171);
and U809 (N_809,In_1050,In_1708);
and U810 (N_810,In_2839,In_38);
or U811 (N_811,In_2752,In_1851);
xnor U812 (N_812,In_2246,In_1150);
nand U813 (N_813,In_1751,In_2289);
nor U814 (N_814,In_1357,In_837);
and U815 (N_815,In_1512,In_1181);
nand U816 (N_816,In_2832,In_2699);
nand U817 (N_817,In_269,In_571);
or U818 (N_818,In_910,In_2739);
and U819 (N_819,In_884,In_1786);
or U820 (N_820,In_1381,In_790);
nand U821 (N_821,In_1234,In_6);
and U822 (N_822,In_1901,In_2140);
or U823 (N_823,In_1683,In_2534);
xnor U824 (N_824,In_1466,In_150);
and U825 (N_825,In_625,In_1763);
nand U826 (N_826,In_2932,In_1198);
or U827 (N_827,In_245,In_459);
or U828 (N_828,In_2857,In_673);
nand U829 (N_829,In_254,In_655);
nand U830 (N_830,In_373,In_642);
nor U831 (N_831,In_939,In_562);
nand U832 (N_832,In_455,In_435);
or U833 (N_833,In_280,In_870);
and U834 (N_834,In_2868,In_498);
nor U835 (N_835,In_206,In_2504);
nor U836 (N_836,In_47,In_2422);
nor U837 (N_837,In_1575,In_1583);
or U838 (N_838,In_2265,In_1254);
and U839 (N_839,In_2777,In_1069);
and U840 (N_840,In_2925,In_2979);
and U841 (N_841,In_2030,In_2596);
or U842 (N_842,In_703,In_377);
nor U843 (N_843,In_529,In_1293);
nor U844 (N_844,In_411,In_2469);
or U845 (N_845,In_1919,In_307);
nor U846 (N_846,In_2881,In_1739);
and U847 (N_847,In_1367,In_186);
nor U848 (N_848,In_2825,In_2396);
and U849 (N_849,In_1718,In_266);
or U850 (N_850,In_979,In_2996);
or U851 (N_851,In_520,In_2575);
nor U852 (N_852,In_1231,In_1648);
nor U853 (N_853,In_1747,In_337);
or U854 (N_854,In_2159,In_1470);
nor U855 (N_855,In_704,In_109);
nor U856 (N_856,In_1676,In_2938);
nor U857 (N_857,In_1637,In_1731);
nor U858 (N_858,In_350,In_282);
and U859 (N_859,In_2407,In_862);
or U860 (N_860,In_438,In_1273);
nor U861 (N_861,In_2676,In_2208);
and U862 (N_862,In_431,In_1709);
or U863 (N_863,In_235,In_741);
or U864 (N_864,In_401,In_1590);
or U865 (N_865,In_2783,In_967);
nor U866 (N_866,In_1398,In_340);
nor U867 (N_867,In_1408,In_1447);
and U868 (N_868,In_335,In_946);
or U869 (N_869,In_579,In_2623);
or U870 (N_870,In_2957,In_341);
and U871 (N_871,In_2588,In_2257);
and U872 (N_872,In_956,In_2931);
xor U873 (N_873,In_2151,In_491);
nand U874 (N_874,In_1889,In_2982);
nand U875 (N_875,In_2073,In_507);
or U876 (N_876,In_2463,In_366);
or U877 (N_877,In_1890,In_911);
nand U878 (N_878,In_849,In_2347);
and U879 (N_879,In_1148,In_1896);
and U880 (N_880,In_1707,In_776);
nor U881 (N_881,In_196,In_899);
nor U882 (N_882,In_2431,In_1265);
nor U883 (N_883,In_1377,In_2764);
nand U884 (N_884,In_1499,In_2899);
nor U885 (N_885,In_1879,In_2815);
and U886 (N_886,In_2352,In_1566);
nand U887 (N_887,In_210,In_1624);
or U888 (N_888,In_218,In_2117);
nor U889 (N_889,In_359,In_833);
nand U890 (N_890,In_1979,In_2601);
or U891 (N_891,In_1799,In_60);
nand U892 (N_892,In_1215,In_281);
or U893 (N_893,In_2907,In_1444);
nor U894 (N_894,In_1600,In_1326);
or U895 (N_895,In_324,In_720);
or U896 (N_896,In_2135,In_343);
and U897 (N_897,In_1972,In_1940);
or U898 (N_898,In_872,In_1084);
and U899 (N_899,In_456,In_1063);
nand U900 (N_900,In_2401,In_2242);
or U901 (N_901,In_1578,In_971);
or U902 (N_902,In_1837,In_2707);
and U903 (N_903,In_1101,In_391);
nand U904 (N_904,In_1169,In_923);
nand U905 (N_905,In_977,In_1308);
nand U906 (N_906,In_2182,In_2560);
nand U907 (N_907,In_12,In_1907);
xor U908 (N_908,In_1544,In_957);
nor U909 (N_909,In_1556,In_2566);
or U910 (N_910,In_1353,In_1587);
or U911 (N_911,In_2966,In_620);
and U912 (N_912,In_2192,In_155);
or U913 (N_913,In_2840,In_90);
or U914 (N_914,In_2686,In_889);
or U915 (N_915,In_315,In_239);
or U916 (N_916,In_1478,In_1157);
nor U917 (N_917,In_387,In_1954);
nor U918 (N_918,In_1838,In_2113);
nand U919 (N_919,In_813,In_2978);
or U920 (N_920,In_962,In_2305);
and U921 (N_921,In_583,In_2040);
nand U922 (N_922,In_699,In_36);
nor U923 (N_923,In_400,In_997);
nand U924 (N_924,In_1768,In_1269);
or U925 (N_925,In_1037,In_2675);
nor U926 (N_926,In_599,In_1631);
and U927 (N_927,In_2236,In_1003);
and U928 (N_928,In_2690,In_860);
nand U929 (N_929,In_991,In_937);
nor U930 (N_930,In_398,In_726);
nand U931 (N_931,In_1315,In_893);
nor U932 (N_932,In_719,In_1094);
and U933 (N_933,In_1891,In_1580);
or U934 (N_934,In_2237,In_1933);
or U935 (N_935,In_2518,In_82);
xnor U936 (N_936,In_1392,In_63);
xnor U937 (N_937,In_446,In_1509);
xor U938 (N_938,In_2009,In_2796);
and U939 (N_939,In_696,In_1698);
or U940 (N_940,In_265,In_2243);
or U941 (N_941,In_539,In_510);
and U942 (N_942,In_385,In_705);
and U943 (N_943,In_810,In_616);
or U944 (N_944,In_2090,In_2133);
nand U945 (N_945,In_2540,In_1441);
nor U946 (N_946,In_2531,In_2104);
and U947 (N_947,In_1498,In_126);
or U948 (N_948,In_877,In_1080);
nand U949 (N_949,In_2584,In_1115);
nor U950 (N_950,In_121,In_2656);
nor U951 (N_951,In_1667,In_2262);
and U952 (N_952,In_891,In_722);
nand U953 (N_953,In_1765,In_1314);
or U954 (N_954,In_2876,In_1111);
nand U955 (N_955,In_1434,In_1350);
nand U956 (N_956,In_1185,In_494);
and U957 (N_957,In_2324,In_1421);
nand U958 (N_958,In_237,In_2800);
and U959 (N_959,In_1653,In_148);
nor U960 (N_960,In_1021,In_2394);
nor U961 (N_961,In_2216,In_1160);
xor U962 (N_962,In_2095,In_2492);
nand U963 (N_963,In_1895,In_84);
and U964 (N_964,In_1247,In_2165);
xor U965 (N_965,In_259,In_177);
nand U966 (N_966,In_2797,In_1960);
or U967 (N_967,In_1018,In_2595);
nand U968 (N_968,In_2053,In_556);
and U969 (N_969,In_2408,In_2036);
xnor U970 (N_970,In_2958,In_70);
and U971 (N_971,In_1483,In_914);
and U972 (N_972,In_2666,In_2392);
or U973 (N_973,In_1909,In_2206);
nand U974 (N_974,In_1172,In_1547);
nand U975 (N_975,In_1179,In_947);
nand U976 (N_976,In_2695,In_2705);
nand U977 (N_977,In_2209,In_1492);
or U978 (N_978,In_1290,In_2035);
and U979 (N_979,In_652,In_1122);
nor U980 (N_980,In_73,In_2129);
and U981 (N_981,In_1378,In_2854);
and U982 (N_982,In_449,In_2255);
xor U983 (N_983,In_130,In_954);
or U984 (N_984,In_2177,In_1903);
and U985 (N_985,In_1248,In_1061);
or U986 (N_986,In_2072,In_1738);
and U987 (N_987,In_2918,In_2234);
nor U988 (N_988,In_531,In_30);
nand U989 (N_989,In_632,In_1209);
and U990 (N_990,In_1205,In_1354);
nor U991 (N_991,In_1136,In_1457);
xor U992 (N_992,In_2089,In_800);
nand U993 (N_993,In_2554,In_1646);
nand U994 (N_994,In_141,In_1932);
nand U995 (N_995,In_1321,In_32);
xnor U996 (N_996,In_2607,In_476);
or U997 (N_997,In_2790,In_2806);
xor U998 (N_998,In_2565,In_1410);
nand U999 (N_999,In_1126,In_2211);
nand U1000 (N_1000,In_1435,In_875);
or U1001 (N_1001,In_65,In_1497);
or U1002 (N_1002,In_815,In_856);
nor U1003 (N_1003,In_207,In_2993);
xor U1004 (N_1004,In_13,In_1892);
and U1005 (N_1005,In_2224,In_2343);
nor U1006 (N_1006,In_1619,In_1211);
or U1007 (N_1007,In_921,In_1048);
and U1008 (N_1008,In_2998,In_1785);
nand U1009 (N_1009,In_592,In_112);
or U1010 (N_1010,In_2278,In_33);
or U1011 (N_1011,In_565,In_2071);
nand U1012 (N_1012,In_2592,In_1582);
nor U1013 (N_1013,In_2461,In_1431);
and U1014 (N_1014,In_2249,In_354);
or U1015 (N_1015,In_2099,In_845);
nor U1016 (N_1016,In_783,In_375);
or U1017 (N_1017,In_44,In_136);
and U1018 (N_1018,In_1311,In_861);
and U1019 (N_1019,In_978,In_2481);
or U1020 (N_1020,In_1748,In_243);
nand U1021 (N_1021,In_2102,In_913);
and U1022 (N_1022,In_1086,In_608);
or U1023 (N_1023,In_1147,In_857);
nor U1024 (N_1024,In_960,In_1613);
and U1025 (N_1025,In_287,In_927);
and U1026 (N_1026,In_1100,In_1194);
nor U1027 (N_1027,In_635,In_869);
nand U1028 (N_1028,In_2448,In_596);
nor U1029 (N_1029,In_2075,In_527);
nand U1030 (N_1030,In_1364,In_410);
or U1031 (N_1031,In_2202,In_1585);
nand U1032 (N_1032,In_1088,In_59);
and U1033 (N_1033,In_203,In_1570);
nor U1034 (N_1034,In_62,In_687);
and U1035 (N_1035,In_540,In_2703);
and U1036 (N_1036,In_2502,In_2541);
nor U1037 (N_1037,In_1462,In_407);
xor U1038 (N_1038,In_2388,In_23);
nand U1039 (N_1039,In_762,In_1988);
and U1040 (N_1040,In_2330,In_499);
and U1041 (N_1041,In_1355,In_1102);
nand U1042 (N_1042,In_1422,In_2331);
nor U1043 (N_1043,In_2039,In_1388);
or U1044 (N_1044,In_853,In_2818);
nor U1045 (N_1045,In_165,In_2001);
xnor U1046 (N_1046,In_188,In_11);
nand U1047 (N_1047,In_2775,In_2786);
nor U1048 (N_1048,In_2834,In_2860);
nand U1049 (N_1049,In_1961,In_2393);
and U1050 (N_1050,In_1959,In_1639);
nand U1051 (N_1051,In_874,In_440);
or U1052 (N_1052,In_2807,In_163);
and U1053 (N_1053,In_1202,In_1956);
and U1054 (N_1054,In_990,In_2530);
or U1055 (N_1055,In_1640,In_1684);
and U1056 (N_1056,In_289,In_2527);
nand U1057 (N_1057,In_1138,In_1305);
and U1058 (N_1058,In_1539,In_2935);
nand U1059 (N_1059,In_2486,In_2605);
nor U1060 (N_1060,In_2285,In_502);
or U1061 (N_1061,In_1089,In_2517);
and U1062 (N_1062,In_1473,In_17);
nand U1063 (N_1063,In_768,In_153);
nand U1064 (N_1064,In_1921,In_1175);
or U1065 (N_1065,In_333,In_249);
and U1066 (N_1066,In_1039,In_972);
and U1067 (N_1067,In_805,In_936);
or U1068 (N_1068,In_867,In_1195);
and U1069 (N_1069,In_1085,In_2638);
nor U1070 (N_1070,In_1579,In_1716);
and U1071 (N_1071,In_1062,In_1779);
and U1072 (N_1072,In_1615,In_2823);
nand U1073 (N_1073,In_2660,In_2451);
nand U1074 (N_1074,In_1517,In_1327);
nor U1075 (N_1075,In_2115,In_1256);
nor U1076 (N_1076,In_1262,In_2767);
or U1077 (N_1077,In_2955,In_1394);
nand U1078 (N_1078,In_2363,In_2735);
and U1079 (N_1079,In_2875,In_1689);
and U1080 (N_1080,In_1878,In_46);
nor U1081 (N_1081,In_649,In_4);
and U1082 (N_1082,In_1060,In_145);
nor U1083 (N_1083,In_597,In_2467);
or U1084 (N_1084,In_1506,In_2729);
nand U1085 (N_1085,In_2188,In_297);
nand U1086 (N_1086,In_367,In_2365);
nor U1087 (N_1087,In_128,In_834);
xnor U1088 (N_1088,In_2870,In_227);
nor U1089 (N_1089,In_1564,In_582);
xnor U1090 (N_1090,In_439,In_2977);
xor U1091 (N_1091,In_78,In_820);
and U1092 (N_1092,In_2654,In_86);
nor U1093 (N_1093,In_2590,In_2097);
or U1094 (N_1094,In_1129,In_1875);
and U1095 (N_1095,In_453,In_2694);
and U1096 (N_1096,In_2377,In_985);
and U1097 (N_1097,In_2594,In_256);
and U1098 (N_1098,In_1562,In_1274);
nand U1099 (N_1099,In_1486,In_2003);
or U1100 (N_1100,In_733,In_1843);
or U1101 (N_1101,In_2124,In_1156);
or U1102 (N_1102,In_2587,In_743);
nand U1103 (N_1103,In_1374,In_639);
nand U1104 (N_1104,In_412,In_2708);
or U1105 (N_1105,In_931,In_2256);
nand U1106 (N_1106,In_2734,In_1592);
and U1107 (N_1107,In_1154,In_2491);
nand U1108 (N_1108,In_139,In_912);
nor U1109 (N_1109,In_1489,In_1008);
xnor U1110 (N_1110,In_1773,In_2161);
and U1111 (N_1111,In_357,In_1797);
nand U1112 (N_1112,In_270,In_1815);
and U1113 (N_1113,In_2475,In_2736);
and U1114 (N_1114,In_2545,In_2910);
or U1115 (N_1115,In_622,In_1331);
nand U1116 (N_1116,In_770,In_1133);
and U1117 (N_1117,In_2987,In_1951);
or U1118 (N_1118,In_924,In_1124);
nand U1119 (N_1119,In_1033,In_1742);
and U1120 (N_1120,In_2772,In_2190);
nand U1121 (N_1121,In_1178,In_213);
xnor U1122 (N_1122,In_1442,In_578);
nand U1123 (N_1123,In_2990,In_2167);
or U1124 (N_1124,In_988,In_1214);
and U1125 (N_1125,In_2136,In_311);
nand U1126 (N_1126,In_71,In_2045);
nor U1127 (N_1127,In_2828,In_1894);
or U1128 (N_1128,In_447,In_1827);
and U1129 (N_1129,In_1557,In_1146);
and U1130 (N_1130,In_2164,In_1936);
or U1131 (N_1131,In_681,In_551);
or U1132 (N_1132,In_2362,In_624);
nand U1133 (N_1133,In_1002,In_2213);
nand U1134 (N_1134,In_684,In_56);
xor U1135 (N_1135,In_1508,In_24);
nor U1136 (N_1136,In_96,In_2229);
or U1137 (N_1137,In_2015,In_1559);
nor U1138 (N_1138,In_1461,In_1504);
nor U1139 (N_1139,In_202,In_483);
xnor U1140 (N_1140,In_2007,In_2450);
nor U1141 (N_1141,In_2766,In_898);
nand U1142 (N_1142,In_2147,In_413);
nand U1143 (N_1143,In_2637,In_835);
and U1144 (N_1144,In_2640,In_2619);
or U1145 (N_1145,In_1001,In_394);
nand U1146 (N_1146,In_57,In_199);
and U1147 (N_1147,In_633,In_2276);
or U1148 (N_1148,In_2984,In_817);
nand U1149 (N_1149,In_514,In_2275);
nor U1150 (N_1150,In_371,In_2717);
nand U1151 (N_1151,In_2226,In_515);
nand U1152 (N_1152,In_2105,In_1190);
nor U1153 (N_1153,In_816,In_2831);
nor U1154 (N_1154,In_2811,In_736);
and U1155 (N_1155,In_1906,In_1437);
nand U1156 (N_1156,In_2389,In_1075);
and U1157 (N_1157,In_1651,In_426);
nor U1158 (N_1158,In_1534,In_1758);
nor U1159 (N_1159,In_595,In_2616);
nand U1160 (N_1160,In_201,In_2439);
or U1161 (N_1161,In_1623,In_2406);
and U1162 (N_1162,In_1519,In_2189);
nor U1163 (N_1163,In_1732,In_497);
nor U1164 (N_1164,In_557,In_638);
nor U1165 (N_1165,In_230,In_895);
and U1166 (N_1166,In_423,In_879);
and U1167 (N_1167,In_495,In_587);
xor U1168 (N_1168,In_1199,In_420);
and U1169 (N_1169,In_2780,In_1766);
and U1170 (N_1170,In_2892,In_416);
xnor U1171 (N_1171,In_2008,In_2889);
nor U1172 (N_1172,In_757,In_1351);
or U1173 (N_1173,In_2296,In_2196);
and U1174 (N_1174,In_1152,In_838);
or U1175 (N_1175,In_1760,In_1176);
or U1176 (N_1176,In_553,In_660);
or U1177 (N_1177,In_1204,In_2341);
nor U1178 (N_1178,In_1400,In_2148);
nand U1179 (N_1179,In_2864,In_2350);
nand U1180 (N_1180,In_2395,In_1005);
xor U1181 (N_1181,In_1405,In_45);
and U1182 (N_1182,In_2569,In_2361);
nand U1183 (N_1183,In_2144,In_2480);
or U1184 (N_1184,In_2801,In_477);
and U1185 (N_1185,In_378,In_348);
nor U1186 (N_1186,In_1674,In_535);
nor U1187 (N_1187,In_1645,In_2066);
nand U1188 (N_1188,In_2826,In_1139);
nor U1189 (N_1189,In_178,In_118);
nand U1190 (N_1190,In_1456,In_2629);
and U1191 (N_1191,In_1106,In_429);
xnor U1192 (N_1192,In_2700,In_1989);
or U1193 (N_1193,In_288,In_688);
nand U1194 (N_1194,In_1997,In_1771);
and U1195 (N_1195,In_34,In_2999);
and U1196 (N_1196,In_2070,In_1835);
and U1197 (N_1197,In_2673,In_516);
nand U1198 (N_1198,In_267,In_147);
nand U1199 (N_1199,In_1691,In_1635);
or U1200 (N_1200,In_312,In_1170);
or U1201 (N_1201,In_839,In_868);
or U1202 (N_1202,In_2770,In_1618);
and U1203 (N_1203,In_417,In_2410);
and U1204 (N_1204,In_1671,In_195);
nor U1205 (N_1205,In_313,In_1772);
and U1206 (N_1206,In_2415,In_1601);
nand U1207 (N_1207,In_2963,In_1266);
nor U1208 (N_1208,In_405,In_525);
xor U1209 (N_1209,In_1280,In_67);
nand U1210 (N_1210,In_1692,In_1784);
nor U1211 (N_1211,In_1885,In_1605);
or U1212 (N_1212,In_1287,In_1641);
nor U1213 (N_1213,In_1306,In_472);
nor U1214 (N_1214,In_555,In_2850);
and U1215 (N_1215,In_2400,In_686);
or U1216 (N_1216,In_2349,In_2298);
and U1217 (N_1217,In_2041,In_395);
and U1218 (N_1218,In_176,In_644);
nand U1219 (N_1219,In_1705,In_607);
or U1220 (N_1220,In_2928,In_2005);
xor U1221 (N_1221,In_2304,In_2862);
nor U1222 (N_1222,In_2636,In_2424);
nand U1223 (N_1223,In_897,In_710);
nor U1224 (N_1224,In_1307,In_383);
and U1225 (N_1225,In_2544,In_1984);
xnor U1226 (N_1226,In_286,In_1833);
nand U1227 (N_1227,In_461,In_1041);
nand U1228 (N_1228,In_1551,In_2810);
nand U1229 (N_1229,In_1867,In_504);
and U1230 (N_1230,In_21,In_2286);
and U1231 (N_1231,In_1589,In_1463);
xnor U1232 (N_1232,In_2774,In_1414);
xor U1233 (N_1233,In_570,In_1275);
or U1234 (N_1234,In_2536,In_204);
nand U1235 (N_1235,In_2449,In_2309);
xnor U1236 (N_1236,In_1573,In_2950);
or U1237 (N_1237,In_492,In_2894);
nand U1238 (N_1238,In_2946,In_1812);
and U1239 (N_1239,In_2771,In_1448);
nor U1240 (N_1240,In_934,In_1608);
nor U1241 (N_1241,In_1324,In_2051);
nor U1242 (N_1242,In_822,In_2170);
nand U1243 (N_1243,In_1191,In_1376);
xor U1244 (N_1244,In_1188,In_2981);
and U1245 (N_1245,In_1962,In_142);
nor U1246 (N_1246,In_2444,In_1411);
nand U1247 (N_1247,In_1166,In_567);
and U1248 (N_1248,In_2836,In_1638);
nand U1249 (N_1249,In_2858,In_293);
or U1250 (N_1250,In_2383,In_1913);
or U1251 (N_1251,In_2327,In_698);
xor U1252 (N_1252,In_961,In_1994);
or U1253 (N_1253,In_2048,In_285);
and U1254 (N_1254,In_1295,In_1533);
nor U1255 (N_1255,In_1413,In_490);
nand U1256 (N_1256,In_892,In_2203);
nor U1257 (N_1257,In_2626,In_1852);
xor U1258 (N_1258,In_523,In_1888);
nor U1259 (N_1259,In_752,In_2961);
nor U1260 (N_1260,In_2813,In_1864);
or U1261 (N_1261,In_2482,In_1058);
nand U1262 (N_1262,In_1193,In_746);
nor U1263 (N_1263,In_2885,In_2483);
and U1264 (N_1264,In_1745,In_2301);
nand U1265 (N_1265,In_2049,In_1796);
or U1266 (N_1266,In_2384,In_2338);
xnor U1267 (N_1267,In_1787,In_2689);
or U1268 (N_1268,In_1846,In_2529);
nand U1269 (N_1269,In_2747,In_2471);
xor U1270 (N_1270,In_2947,In_1882);
and U1271 (N_1271,In_980,In_989);
and U1272 (N_1272,In_292,In_309);
nand U1273 (N_1273,In_2440,In_2434);
nand U1274 (N_1274,In_1389,In_2577);
nand U1275 (N_1275,In_2954,In_2641);
or U1276 (N_1276,In_2201,In_683);
xor U1277 (N_1277,In_1035,In_271);
or U1278 (N_1278,In_2568,In_81);
or U1279 (N_1279,In_2354,In_796);
and U1280 (N_1280,In_1332,In_2914);
or U1281 (N_1281,In_2391,In_339);
or U1282 (N_1282,In_1121,In_299);
and U1283 (N_1283,In_277,In_1865);
and U1284 (N_1284,In_2096,In_2386);
or U1285 (N_1285,In_992,In_1140);
xnor U1286 (N_1286,In_464,In_2313);
nand U1287 (N_1287,In_390,In_1685);
and U1288 (N_1288,In_2750,In_1375);
and U1289 (N_1289,In_2661,In_1427);
or U1290 (N_1290,In_2385,In_2821);
and U1291 (N_1291,In_2653,In_2716);
or U1292 (N_1292,In_658,In_1845);
xnor U1293 (N_1293,In_779,In_1059);
and U1294 (N_1294,In_1318,In_706);
or U1295 (N_1295,In_2520,In_1449);
and U1296 (N_1296,In_2878,In_501);
and U1297 (N_1297,In_1443,In_2114);
and U1298 (N_1298,In_2633,In_187);
nand U1299 (N_1299,In_183,In_2621);
and U1300 (N_1300,In_468,In_2319);
nand U1301 (N_1301,In_1560,In_2178);
and U1302 (N_1302,In_2679,In_1791);
nor U1303 (N_1303,In_3,In_2547);
nor U1304 (N_1304,In_2643,In_117);
and U1305 (N_1305,In_1767,In_1595);
nor U1306 (N_1306,In_442,In_787);
and U1307 (N_1307,In_1788,In_2430);
or U1308 (N_1308,In_903,In_1996);
xor U1309 (N_1309,In_125,In_1810);
or U1310 (N_1310,In_2019,In_1733);
or U1311 (N_1311,In_2141,In_1496);
nor U1312 (N_1312,In_2078,In_1429);
or U1313 (N_1313,In_1710,In_2532);
nor U1314 (N_1314,In_1098,In_953);
xnor U1315 (N_1315,In_160,In_1343);
or U1316 (N_1316,In_1964,In_1917);
nor U1317 (N_1317,In_2118,In_2284);
and U1318 (N_1318,In_728,In_2972);
or U1319 (N_1319,In_8,In_1046);
xor U1320 (N_1320,In_1261,In_1436);
or U1321 (N_1321,In_172,In_1981);
nand U1322 (N_1322,In_174,In_2034);
or U1323 (N_1323,In_1384,In_568);
nor U1324 (N_1324,In_2274,In_244);
nor U1325 (N_1325,In_1902,In_2311);
and U1326 (N_1326,In_2241,In_2591);
nor U1327 (N_1327,In_1876,In_2538);
nand U1328 (N_1328,In_2126,In_2353);
nor U1329 (N_1329,In_1145,In_667);
xor U1330 (N_1330,In_1783,In_430);
nor U1331 (N_1331,In_2134,In_1109);
xnor U1332 (N_1332,In_1143,In_1762);
nand U1333 (N_1333,In_1531,In_2076);
and U1334 (N_1334,In_1057,In_2751);
or U1335 (N_1335,In_576,In_1281);
nand U1336 (N_1336,In_1161,In_406);
nor U1337 (N_1337,In_1863,In_92);
and U1338 (N_1338,In_522,In_973);
nor U1339 (N_1339,In_664,In_852);
and U1340 (N_1340,In_1252,In_2227);
or U1341 (N_1341,In_959,In_2503);
and U1342 (N_1342,In_636,In_731);
and U1343 (N_1343,In_1944,In_750);
or U1344 (N_1344,In_1664,In_524);
nand U1345 (N_1345,In_2922,In_1356);
or U1346 (N_1346,In_480,In_854);
and U1347 (N_1347,In_995,In_500);
or U1348 (N_1348,In_1368,In_1813);
nor U1349 (N_1349,In_1015,In_1424);
nor U1350 (N_1350,In_2916,In_2173);
nand U1351 (N_1351,In_2901,In_1597);
nor U1352 (N_1352,In_2218,In_1366);
nor U1353 (N_1353,In_904,In_1192);
nor U1354 (N_1354,In_197,In_1746);
and U1355 (N_1355,In_2576,In_2913);
nand U1356 (N_1356,In_1581,In_133);
or U1357 (N_1357,In_1407,In_110);
nand U1358 (N_1358,In_1724,In_362);
nand U1359 (N_1359,In_1151,In_2693);
or U1360 (N_1360,In_2748,In_909);
or U1361 (N_1361,In_2976,In_1943);
nor U1362 (N_1362,In_955,In_2551);
nor U1363 (N_1363,In_1611,In_1586);
or U1364 (N_1364,In_1371,In_1322);
xor U1365 (N_1365,In_2348,In_2488);
nor U1366 (N_1366,In_674,In_152);
nand U1367 (N_1367,In_192,In_2217);
nand U1368 (N_1368,In_179,In_2830);
nor U1369 (N_1369,In_2809,In_319);
xor U1370 (N_1370,In_850,In_2793);
and U1371 (N_1371,In_262,In_2316);
and U1372 (N_1372,In_224,In_799);
and U1373 (N_1373,In_1184,In_1629);
or U1374 (N_1374,In_1627,In_1251);
and U1375 (N_1375,In_1032,In_43);
or U1376 (N_1376,In_66,In_326);
or U1377 (N_1377,In_2088,In_1668);
nor U1378 (N_1378,In_2382,In_1014);
nor U1379 (N_1379,In_600,In_1323);
nor U1380 (N_1380,In_2179,In_2297);
nand U1381 (N_1381,In_2364,In_1513);
and U1382 (N_1382,In_888,In_2245);
nor U1383 (N_1383,In_2847,In_1474);
or U1384 (N_1384,In_2585,In_1726);
nor U1385 (N_1385,In_2292,In_300);
or U1386 (N_1386,In_261,In_1056);
and U1387 (N_1387,In_2322,In_2668);
nand U1388 (N_1388,In_2874,In_538);
or U1389 (N_1389,In_2098,In_2169);
nand U1390 (N_1390,In_372,In_2094);
xor U1391 (N_1391,In_1336,In_880);
nor U1392 (N_1392,In_1795,In_1535);
nor U1393 (N_1393,In_2084,In_2057);
nand U1394 (N_1394,In_2711,In_2655);
and U1395 (N_1395,In_2886,In_918);
nor U1396 (N_1396,In_590,In_2980);
nand U1397 (N_1397,In_1657,In_7);
nor U1398 (N_1398,In_1794,In_2819);
and U1399 (N_1399,In_1501,In_1488);
and U1400 (N_1400,In_1712,In_2472);
nand U1401 (N_1401,In_2342,In_2697);
nor U1402 (N_1402,In_2720,In_264);
nand U1403 (N_1403,In_2403,In_404);
or U1404 (N_1404,In_922,In_2004);
or U1405 (N_1405,In_114,In_1249);
nand U1406 (N_1406,In_99,In_1286);
or U1407 (N_1407,In_2180,In_2967);
or U1408 (N_1408,In_2239,In_2992);
nand U1409 (N_1409,In_744,In_695);
or U1410 (N_1410,In_1949,In_2500);
nor U1411 (N_1411,In_714,In_2759);
or U1412 (N_1412,In_1125,In_1968);
nor U1413 (N_1413,In_2108,In_1754);
or U1414 (N_1414,In_613,In_908);
or U1415 (N_1415,In_2667,In_2833);
and U1416 (N_1416,In_1942,In_2435);
or U1417 (N_1417,In_508,In_2);
nand U1418 (N_1418,In_2092,In_604);
nand U1419 (N_1419,In_1877,In_2782);
nand U1420 (N_1420,In_742,In_1013);
nor U1421 (N_1421,In_2669,In_2374);
xnor U1422 (N_1422,In_1279,In_668);
nand U1423 (N_1423,In_35,In_2618);
and U1424 (N_1424,In_788,In_1168);
or U1425 (N_1425,In_1043,In_1383);
nor U1426 (N_1426,In_2119,In_2458);
nor U1427 (N_1427,In_1445,In_2199);
nand U1428 (N_1428,In_2186,In_2058);
nor U1429 (N_1429,In_1268,In_1163);
nor U1430 (N_1430,In_1690,In_2445);
or U1431 (N_1431,In_792,In_2677);
or U1432 (N_1432,In_2174,In_797);
nand U1433 (N_1433,In_2116,In_1283);
xor U1434 (N_1434,In_189,In_1164);
and U1435 (N_1435,In_506,In_1238);
and U1436 (N_1436,In_1220,In_1419);
or U1437 (N_1437,In_713,In_1103);
or U1438 (N_1438,In_2321,In_804);
nor U1439 (N_1439,In_1594,In_2682);
and U1440 (N_1440,In_1453,In_2270);
nand U1441 (N_1441,In_709,In_2890);
nor U1442 (N_1442,In_94,In_1725);
and U1443 (N_1443,In_878,In_2172);
and U1444 (N_1444,In_113,In_88);
or U1445 (N_1445,In_2579,In_1490);
nor U1446 (N_1446,In_325,In_1941);
nor U1447 (N_1447,In_843,In_1858);
or U1448 (N_1448,In_808,In_1476);
nor U1449 (N_1449,In_2131,In_1614);
nor U1450 (N_1450,In_100,In_2028);
and U1451 (N_1451,In_1284,In_50);
xnor U1452 (N_1452,In_1528,In_2086);
or U1453 (N_1453,In_2960,In_1975);
and U1454 (N_1454,In_1782,In_1966);
and U1455 (N_1455,In_840,In_1380);
nor U1456 (N_1456,In_1694,In_2511);
nor U1457 (N_1457,In_1189,In_1596);
nor U1458 (N_1458,In_40,In_1370);
and U1459 (N_1459,In_2427,In_260);
xor U1460 (N_1460,In_1695,In_1659);
and U1461 (N_1461,In_2749,In_1469);
or U1462 (N_1462,In_144,In_1604);
and U1463 (N_1463,In_569,In_1717);
or U1464 (N_1464,In_2484,In_1971);
or U1465 (N_1465,In_789,In_830);
or U1466 (N_1466,In_1119,In_2563);
or U1467 (N_1467,In_968,In_2038);
xnor U1468 (N_1468,In_2067,In_2523);
or U1469 (N_1469,In_457,In_1826);
and U1470 (N_1470,In_701,In_944);
nand U1471 (N_1471,In_225,In_829);
nand U1472 (N_1472,In_825,In_1829);
or U1473 (N_1473,In_1680,In_236);
nor U1474 (N_1474,In_1856,In_640);
or U1475 (N_1475,In_2442,In_2897);
or U1476 (N_1476,In_170,In_1183);
nor U1477 (N_1477,In_2244,In_317);
or U1478 (N_1478,In_2646,In_732);
xnor U1479 (N_1479,In_2732,In_1781);
nor U1480 (N_1480,In_777,In_1372);
nor U1481 (N_1481,In_665,In_2453);
and U1482 (N_1482,In_2558,In_154);
xnor U1483 (N_1483,In_2593,In_2758);
nand U1484 (N_1484,In_41,In_1267);
xnor U1485 (N_1485,In_2060,In_2022);
nand U1486 (N_1486,In_1952,In_1908);
and U1487 (N_1487,In_1565,In_470);
or U1488 (N_1488,In_2877,In_454);
nand U1489 (N_1489,In_2254,In_1699);
and U1490 (N_1490,In_1769,In_1396);
or U1491 (N_1491,In_2949,In_408);
nand U1492 (N_1492,In_83,In_2962);
nor U1493 (N_1493,In_711,In_2701);
and U1494 (N_1494,In_2064,In_481);
nor U1495 (N_1495,In_975,In_2123);
or U1496 (N_1496,In_2930,In_2085);
nand U1497 (N_1497,In_1606,In_2943);
and U1498 (N_1498,In_2006,In_253);
or U1499 (N_1499,In_1312,In_1329);
nor U1500 (N_1500,In_2649,In_361);
or U1501 (N_1501,In_2777,In_2435);
and U1502 (N_1502,In_652,In_2426);
and U1503 (N_1503,In_2382,In_796);
xnor U1504 (N_1504,In_2406,In_2812);
and U1505 (N_1505,In_2117,In_138);
nand U1506 (N_1506,In_978,In_1396);
nor U1507 (N_1507,In_1834,In_2053);
nor U1508 (N_1508,In_2916,In_2551);
nand U1509 (N_1509,In_2607,In_395);
nand U1510 (N_1510,In_2025,In_760);
and U1511 (N_1511,In_2316,In_1506);
nand U1512 (N_1512,In_1280,In_1816);
or U1513 (N_1513,In_768,In_1611);
nand U1514 (N_1514,In_2757,In_2276);
nand U1515 (N_1515,In_837,In_2163);
nand U1516 (N_1516,In_1722,In_894);
nor U1517 (N_1517,In_1401,In_2650);
nand U1518 (N_1518,In_2250,In_445);
nand U1519 (N_1519,In_2695,In_614);
xor U1520 (N_1520,In_257,In_1708);
nand U1521 (N_1521,In_431,In_404);
or U1522 (N_1522,In_2583,In_220);
nor U1523 (N_1523,In_1847,In_949);
and U1524 (N_1524,In_1142,In_1409);
and U1525 (N_1525,In_84,In_842);
nand U1526 (N_1526,In_2048,In_2896);
or U1527 (N_1527,In_332,In_2247);
and U1528 (N_1528,In_1897,In_1839);
and U1529 (N_1529,In_2913,In_1254);
nor U1530 (N_1530,In_1175,In_2548);
xor U1531 (N_1531,In_325,In_2935);
xnor U1532 (N_1532,In_2608,In_1729);
and U1533 (N_1533,In_1738,In_1108);
or U1534 (N_1534,In_1841,In_2887);
nor U1535 (N_1535,In_1001,In_304);
nor U1536 (N_1536,In_288,In_1204);
or U1537 (N_1537,In_102,In_2468);
nor U1538 (N_1538,In_1477,In_1566);
and U1539 (N_1539,In_2506,In_214);
nand U1540 (N_1540,In_2698,In_2856);
nor U1541 (N_1541,In_1213,In_2687);
and U1542 (N_1542,In_2679,In_2021);
nor U1543 (N_1543,In_791,In_841);
xor U1544 (N_1544,In_1613,In_2008);
nor U1545 (N_1545,In_531,In_629);
nand U1546 (N_1546,In_2164,In_1318);
and U1547 (N_1547,In_826,In_769);
and U1548 (N_1548,In_295,In_805);
and U1549 (N_1549,In_2798,In_2577);
nor U1550 (N_1550,In_934,In_1003);
nor U1551 (N_1551,In_2008,In_1936);
or U1552 (N_1552,In_276,In_2135);
and U1553 (N_1553,In_1410,In_2368);
or U1554 (N_1554,In_2173,In_2579);
nor U1555 (N_1555,In_2942,In_1964);
and U1556 (N_1556,In_284,In_1225);
and U1557 (N_1557,In_209,In_1456);
nand U1558 (N_1558,In_234,In_1080);
nor U1559 (N_1559,In_1678,In_405);
and U1560 (N_1560,In_104,In_424);
or U1561 (N_1561,In_1003,In_559);
or U1562 (N_1562,In_665,In_288);
or U1563 (N_1563,In_58,In_2895);
or U1564 (N_1564,In_694,In_304);
nand U1565 (N_1565,In_737,In_1096);
and U1566 (N_1566,In_2004,In_655);
nand U1567 (N_1567,In_2461,In_2891);
nor U1568 (N_1568,In_271,In_165);
nor U1569 (N_1569,In_1111,In_1490);
and U1570 (N_1570,In_1911,In_1901);
nand U1571 (N_1571,In_2544,In_2115);
and U1572 (N_1572,In_2090,In_2320);
nor U1573 (N_1573,In_2689,In_1282);
nor U1574 (N_1574,In_1356,In_454);
xnor U1575 (N_1575,In_773,In_2468);
or U1576 (N_1576,In_265,In_2627);
and U1577 (N_1577,In_1949,In_1963);
or U1578 (N_1578,In_439,In_970);
nor U1579 (N_1579,In_2506,In_1566);
nor U1580 (N_1580,In_2772,In_36);
or U1581 (N_1581,In_1145,In_897);
nand U1582 (N_1582,In_29,In_762);
or U1583 (N_1583,In_2677,In_1293);
nand U1584 (N_1584,In_156,In_694);
nand U1585 (N_1585,In_2839,In_2912);
nand U1586 (N_1586,In_1585,In_1043);
xnor U1587 (N_1587,In_2249,In_284);
and U1588 (N_1588,In_1495,In_1034);
and U1589 (N_1589,In_2830,In_573);
or U1590 (N_1590,In_910,In_448);
and U1591 (N_1591,In_2048,In_605);
or U1592 (N_1592,In_2793,In_1212);
nor U1593 (N_1593,In_2556,In_833);
and U1594 (N_1594,In_1682,In_2682);
or U1595 (N_1595,In_1646,In_911);
or U1596 (N_1596,In_950,In_2540);
xnor U1597 (N_1597,In_1902,In_1924);
and U1598 (N_1598,In_1646,In_321);
or U1599 (N_1599,In_790,In_1256);
xor U1600 (N_1600,In_2066,In_2415);
or U1601 (N_1601,In_820,In_1030);
or U1602 (N_1602,In_2037,In_2839);
nand U1603 (N_1603,In_1907,In_311);
or U1604 (N_1604,In_583,In_635);
nand U1605 (N_1605,In_553,In_1323);
nand U1606 (N_1606,In_152,In_1171);
nor U1607 (N_1607,In_764,In_1315);
or U1608 (N_1608,In_50,In_2150);
nand U1609 (N_1609,In_1877,In_492);
or U1610 (N_1610,In_1025,In_342);
or U1611 (N_1611,In_70,In_2116);
or U1612 (N_1612,In_936,In_679);
nor U1613 (N_1613,In_900,In_1312);
and U1614 (N_1614,In_1523,In_2228);
nor U1615 (N_1615,In_2896,In_1959);
and U1616 (N_1616,In_2432,In_989);
and U1617 (N_1617,In_1908,In_1850);
nor U1618 (N_1618,In_2015,In_2314);
xnor U1619 (N_1619,In_1284,In_2326);
nor U1620 (N_1620,In_1745,In_2575);
nand U1621 (N_1621,In_1828,In_2847);
nand U1622 (N_1622,In_686,In_1145);
nand U1623 (N_1623,In_2367,In_1001);
nand U1624 (N_1624,In_1242,In_1493);
nor U1625 (N_1625,In_2800,In_646);
nor U1626 (N_1626,In_1166,In_149);
nand U1627 (N_1627,In_1624,In_145);
nor U1628 (N_1628,In_919,In_230);
nor U1629 (N_1629,In_2972,In_465);
and U1630 (N_1630,In_749,In_1423);
or U1631 (N_1631,In_1919,In_639);
xnor U1632 (N_1632,In_998,In_1515);
xnor U1633 (N_1633,In_964,In_2994);
nor U1634 (N_1634,In_1707,In_1074);
or U1635 (N_1635,In_2482,In_199);
xor U1636 (N_1636,In_1839,In_223);
and U1637 (N_1637,In_1571,In_612);
nand U1638 (N_1638,In_2410,In_2196);
xnor U1639 (N_1639,In_2704,In_2792);
nand U1640 (N_1640,In_2796,In_1374);
nor U1641 (N_1641,In_2093,In_2920);
or U1642 (N_1642,In_2880,In_647);
nor U1643 (N_1643,In_1677,In_2930);
or U1644 (N_1644,In_2611,In_1951);
or U1645 (N_1645,In_2272,In_88);
xor U1646 (N_1646,In_2741,In_1849);
and U1647 (N_1647,In_2323,In_2675);
or U1648 (N_1648,In_1468,In_1673);
or U1649 (N_1649,In_2791,In_1252);
nor U1650 (N_1650,In_1573,In_661);
or U1651 (N_1651,In_1224,In_1131);
nor U1652 (N_1652,In_1680,In_1799);
nand U1653 (N_1653,In_2241,In_2235);
nand U1654 (N_1654,In_830,In_52);
nand U1655 (N_1655,In_2235,In_709);
or U1656 (N_1656,In_676,In_122);
and U1657 (N_1657,In_1528,In_2132);
and U1658 (N_1658,In_2121,In_42);
nor U1659 (N_1659,In_2100,In_2875);
or U1660 (N_1660,In_2652,In_889);
or U1661 (N_1661,In_1185,In_1761);
nor U1662 (N_1662,In_2762,In_1570);
nand U1663 (N_1663,In_2003,In_903);
nand U1664 (N_1664,In_919,In_339);
or U1665 (N_1665,In_1686,In_2498);
nor U1666 (N_1666,In_28,In_2591);
nor U1667 (N_1667,In_1988,In_1037);
nand U1668 (N_1668,In_1915,In_879);
nor U1669 (N_1669,In_849,In_2991);
or U1670 (N_1670,In_2867,In_793);
xnor U1671 (N_1671,In_1543,In_2653);
or U1672 (N_1672,In_1726,In_2153);
nand U1673 (N_1673,In_2137,In_1754);
or U1674 (N_1674,In_1756,In_1831);
or U1675 (N_1675,In_943,In_2493);
or U1676 (N_1676,In_450,In_109);
nand U1677 (N_1677,In_2433,In_1131);
or U1678 (N_1678,In_1423,In_505);
or U1679 (N_1679,In_250,In_543);
nand U1680 (N_1680,In_666,In_2174);
nand U1681 (N_1681,In_1300,In_1417);
nor U1682 (N_1682,In_1449,In_1273);
nor U1683 (N_1683,In_2242,In_1246);
and U1684 (N_1684,In_287,In_271);
or U1685 (N_1685,In_1911,In_322);
xnor U1686 (N_1686,In_1307,In_1890);
or U1687 (N_1687,In_2837,In_599);
and U1688 (N_1688,In_891,In_1550);
nor U1689 (N_1689,In_508,In_457);
and U1690 (N_1690,In_1262,In_1134);
xnor U1691 (N_1691,In_1173,In_1688);
or U1692 (N_1692,In_1181,In_113);
xor U1693 (N_1693,In_1766,In_1296);
and U1694 (N_1694,In_1758,In_2635);
and U1695 (N_1695,In_306,In_575);
and U1696 (N_1696,In_2669,In_2202);
nand U1697 (N_1697,In_1291,In_1299);
nor U1698 (N_1698,In_1518,In_2376);
and U1699 (N_1699,In_2549,In_2216);
nand U1700 (N_1700,In_1099,In_1079);
xnor U1701 (N_1701,In_2777,In_2276);
nand U1702 (N_1702,In_2279,In_1271);
nor U1703 (N_1703,In_1716,In_1095);
nand U1704 (N_1704,In_2758,In_554);
or U1705 (N_1705,In_371,In_1957);
nor U1706 (N_1706,In_2965,In_1427);
nand U1707 (N_1707,In_1783,In_652);
or U1708 (N_1708,In_2109,In_2071);
nor U1709 (N_1709,In_97,In_514);
nor U1710 (N_1710,In_2439,In_365);
nand U1711 (N_1711,In_1982,In_1302);
nand U1712 (N_1712,In_1053,In_160);
nor U1713 (N_1713,In_596,In_2437);
nor U1714 (N_1714,In_2251,In_1579);
nor U1715 (N_1715,In_2882,In_703);
nor U1716 (N_1716,In_233,In_2561);
nand U1717 (N_1717,In_80,In_1559);
and U1718 (N_1718,In_2473,In_1268);
nand U1719 (N_1719,In_1458,In_2620);
nand U1720 (N_1720,In_2734,In_1031);
xor U1721 (N_1721,In_2326,In_202);
nand U1722 (N_1722,In_2224,In_2778);
nand U1723 (N_1723,In_1715,In_256);
or U1724 (N_1724,In_1054,In_1082);
nand U1725 (N_1725,In_82,In_1395);
and U1726 (N_1726,In_897,In_823);
and U1727 (N_1727,In_1202,In_54);
nor U1728 (N_1728,In_45,In_1759);
nor U1729 (N_1729,In_1429,In_651);
nor U1730 (N_1730,In_588,In_179);
and U1731 (N_1731,In_140,In_189);
nand U1732 (N_1732,In_1589,In_680);
or U1733 (N_1733,In_2496,In_1533);
nor U1734 (N_1734,In_495,In_2200);
nor U1735 (N_1735,In_2475,In_1739);
xnor U1736 (N_1736,In_221,In_1753);
nand U1737 (N_1737,In_179,In_2720);
nor U1738 (N_1738,In_214,In_914);
or U1739 (N_1739,In_778,In_2040);
or U1740 (N_1740,In_263,In_2869);
nand U1741 (N_1741,In_1331,In_50);
nand U1742 (N_1742,In_2462,In_2477);
and U1743 (N_1743,In_1987,In_259);
or U1744 (N_1744,In_1095,In_1531);
nand U1745 (N_1745,In_2577,In_2366);
xnor U1746 (N_1746,In_2006,In_1533);
nor U1747 (N_1747,In_1881,In_1220);
nand U1748 (N_1748,In_1768,In_1644);
or U1749 (N_1749,In_2491,In_213);
nor U1750 (N_1750,In_1291,In_2558);
nand U1751 (N_1751,In_984,In_362);
nor U1752 (N_1752,In_706,In_925);
nor U1753 (N_1753,In_54,In_454);
nor U1754 (N_1754,In_2278,In_835);
nor U1755 (N_1755,In_52,In_229);
nand U1756 (N_1756,In_428,In_1430);
or U1757 (N_1757,In_835,In_1065);
nor U1758 (N_1758,In_2961,In_1362);
and U1759 (N_1759,In_2230,In_1309);
and U1760 (N_1760,In_2719,In_560);
or U1761 (N_1761,In_1694,In_337);
nand U1762 (N_1762,In_158,In_2400);
nand U1763 (N_1763,In_750,In_1339);
or U1764 (N_1764,In_1460,In_329);
nor U1765 (N_1765,In_2201,In_2647);
or U1766 (N_1766,In_2703,In_653);
xor U1767 (N_1767,In_154,In_665);
nand U1768 (N_1768,In_1222,In_1894);
or U1769 (N_1769,In_1056,In_2192);
or U1770 (N_1770,In_2384,In_1062);
and U1771 (N_1771,In_860,In_2465);
nor U1772 (N_1772,In_1829,In_2466);
or U1773 (N_1773,In_820,In_2240);
nor U1774 (N_1774,In_1125,In_2395);
nor U1775 (N_1775,In_1517,In_641);
and U1776 (N_1776,In_1769,In_1302);
nor U1777 (N_1777,In_1596,In_1732);
and U1778 (N_1778,In_2604,In_1349);
nand U1779 (N_1779,In_1811,In_2653);
and U1780 (N_1780,In_440,In_1224);
or U1781 (N_1781,In_2778,In_3);
nand U1782 (N_1782,In_2094,In_2552);
nand U1783 (N_1783,In_1911,In_1482);
or U1784 (N_1784,In_2490,In_2878);
nand U1785 (N_1785,In_1539,In_2088);
and U1786 (N_1786,In_1343,In_2517);
or U1787 (N_1787,In_675,In_1702);
nor U1788 (N_1788,In_1054,In_272);
nand U1789 (N_1789,In_474,In_2613);
nand U1790 (N_1790,In_1684,In_2777);
and U1791 (N_1791,In_449,In_1968);
or U1792 (N_1792,In_1274,In_2417);
nor U1793 (N_1793,In_167,In_1939);
and U1794 (N_1794,In_1570,In_952);
nand U1795 (N_1795,In_1757,In_2971);
nor U1796 (N_1796,In_97,In_2440);
and U1797 (N_1797,In_2134,In_2087);
nand U1798 (N_1798,In_2660,In_2129);
nor U1799 (N_1799,In_2039,In_980);
nor U1800 (N_1800,In_2628,In_2630);
nor U1801 (N_1801,In_1192,In_781);
xnor U1802 (N_1802,In_2921,In_2544);
nor U1803 (N_1803,In_28,In_2241);
and U1804 (N_1804,In_2927,In_2991);
nand U1805 (N_1805,In_1540,In_2695);
nor U1806 (N_1806,In_2061,In_1387);
and U1807 (N_1807,In_880,In_1536);
and U1808 (N_1808,In_2307,In_2080);
or U1809 (N_1809,In_373,In_1443);
nand U1810 (N_1810,In_1165,In_740);
nor U1811 (N_1811,In_2367,In_401);
and U1812 (N_1812,In_2308,In_1025);
or U1813 (N_1813,In_1529,In_490);
nor U1814 (N_1814,In_2269,In_580);
or U1815 (N_1815,In_1243,In_274);
or U1816 (N_1816,In_2199,In_254);
nand U1817 (N_1817,In_2774,In_1531);
nand U1818 (N_1818,In_2478,In_1336);
and U1819 (N_1819,In_1020,In_1970);
nand U1820 (N_1820,In_2136,In_1686);
or U1821 (N_1821,In_1124,In_659);
or U1822 (N_1822,In_515,In_658);
and U1823 (N_1823,In_57,In_939);
or U1824 (N_1824,In_726,In_2158);
nor U1825 (N_1825,In_204,In_1091);
nand U1826 (N_1826,In_1024,In_1483);
nor U1827 (N_1827,In_477,In_364);
nor U1828 (N_1828,In_505,In_2087);
nor U1829 (N_1829,In_50,In_1639);
and U1830 (N_1830,In_2200,In_1304);
nand U1831 (N_1831,In_735,In_777);
and U1832 (N_1832,In_2278,In_2426);
or U1833 (N_1833,In_415,In_93);
nand U1834 (N_1834,In_2094,In_646);
nor U1835 (N_1835,In_356,In_162);
and U1836 (N_1836,In_2110,In_2660);
nand U1837 (N_1837,In_1210,In_6);
nor U1838 (N_1838,In_488,In_2398);
nor U1839 (N_1839,In_51,In_1906);
nand U1840 (N_1840,In_1660,In_1902);
and U1841 (N_1841,In_1676,In_2438);
or U1842 (N_1842,In_1745,In_2560);
nor U1843 (N_1843,In_1697,In_32);
nand U1844 (N_1844,In_905,In_2439);
nand U1845 (N_1845,In_625,In_2079);
nor U1846 (N_1846,In_2785,In_343);
nand U1847 (N_1847,In_2028,In_2295);
nand U1848 (N_1848,In_335,In_1947);
nand U1849 (N_1849,In_157,In_2162);
nand U1850 (N_1850,In_1761,In_1838);
and U1851 (N_1851,In_2323,In_1776);
nand U1852 (N_1852,In_2797,In_2298);
nor U1853 (N_1853,In_1805,In_2113);
or U1854 (N_1854,In_1972,In_146);
and U1855 (N_1855,In_305,In_2022);
nor U1856 (N_1856,In_981,In_1570);
and U1857 (N_1857,In_2053,In_2586);
and U1858 (N_1858,In_210,In_586);
nor U1859 (N_1859,In_2230,In_103);
nand U1860 (N_1860,In_2115,In_2675);
or U1861 (N_1861,In_2149,In_89);
and U1862 (N_1862,In_604,In_1674);
nand U1863 (N_1863,In_191,In_718);
and U1864 (N_1864,In_2080,In_3);
nand U1865 (N_1865,In_489,In_358);
nand U1866 (N_1866,In_1317,In_1205);
or U1867 (N_1867,In_2578,In_949);
xor U1868 (N_1868,In_1754,In_1231);
nand U1869 (N_1869,In_2586,In_829);
nor U1870 (N_1870,In_1323,In_377);
nor U1871 (N_1871,In_135,In_1256);
nor U1872 (N_1872,In_453,In_1967);
nor U1873 (N_1873,In_1483,In_1249);
or U1874 (N_1874,In_1786,In_525);
nor U1875 (N_1875,In_1187,In_2155);
or U1876 (N_1876,In_11,In_710);
and U1877 (N_1877,In_2714,In_2240);
or U1878 (N_1878,In_594,In_885);
and U1879 (N_1879,In_1921,In_2089);
and U1880 (N_1880,In_891,In_2153);
nor U1881 (N_1881,In_753,In_721);
or U1882 (N_1882,In_1223,In_0);
or U1883 (N_1883,In_1408,In_1691);
and U1884 (N_1884,In_2058,In_2202);
nand U1885 (N_1885,In_711,In_1020);
or U1886 (N_1886,In_1214,In_2745);
nor U1887 (N_1887,In_2436,In_1772);
nand U1888 (N_1888,In_870,In_1382);
nor U1889 (N_1889,In_75,In_641);
and U1890 (N_1890,In_1037,In_167);
nand U1891 (N_1891,In_257,In_2123);
nand U1892 (N_1892,In_748,In_2550);
and U1893 (N_1893,In_743,In_2176);
nor U1894 (N_1894,In_2680,In_2701);
xor U1895 (N_1895,In_2909,In_292);
nor U1896 (N_1896,In_2258,In_1192);
or U1897 (N_1897,In_847,In_1733);
nor U1898 (N_1898,In_1613,In_1411);
or U1899 (N_1899,In_230,In_1490);
or U1900 (N_1900,In_1343,In_2534);
nor U1901 (N_1901,In_2102,In_676);
nand U1902 (N_1902,In_2645,In_563);
nor U1903 (N_1903,In_1488,In_655);
and U1904 (N_1904,In_301,In_1259);
or U1905 (N_1905,In_30,In_110);
and U1906 (N_1906,In_1004,In_1958);
xor U1907 (N_1907,In_2340,In_1346);
nor U1908 (N_1908,In_733,In_2841);
and U1909 (N_1909,In_2824,In_1007);
or U1910 (N_1910,In_2481,In_966);
nand U1911 (N_1911,In_2808,In_991);
nor U1912 (N_1912,In_372,In_2236);
nor U1913 (N_1913,In_835,In_124);
xnor U1914 (N_1914,In_444,In_1560);
nor U1915 (N_1915,In_2731,In_2814);
nor U1916 (N_1916,In_1850,In_1323);
and U1917 (N_1917,In_2686,In_234);
nand U1918 (N_1918,In_2670,In_1897);
and U1919 (N_1919,In_167,In_663);
nor U1920 (N_1920,In_1084,In_2531);
nor U1921 (N_1921,In_1038,In_2870);
or U1922 (N_1922,In_1574,In_1689);
nor U1923 (N_1923,In_2804,In_584);
xor U1924 (N_1924,In_1528,In_271);
or U1925 (N_1925,In_658,In_138);
and U1926 (N_1926,In_359,In_336);
nand U1927 (N_1927,In_1564,In_592);
nor U1928 (N_1928,In_1607,In_1144);
or U1929 (N_1929,In_2935,In_173);
nand U1930 (N_1930,In_2661,In_2434);
or U1931 (N_1931,In_972,In_2209);
or U1932 (N_1932,In_1407,In_1962);
nand U1933 (N_1933,In_1320,In_1142);
or U1934 (N_1934,In_1081,In_2968);
nor U1935 (N_1935,In_2642,In_1912);
nand U1936 (N_1936,In_905,In_776);
or U1937 (N_1937,In_2177,In_307);
nand U1938 (N_1938,In_1670,In_1568);
nand U1939 (N_1939,In_2041,In_1575);
nand U1940 (N_1940,In_2278,In_1386);
or U1941 (N_1941,In_1710,In_1146);
and U1942 (N_1942,In_2724,In_332);
nor U1943 (N_1943,In_776,In_1755);
and U1944 (N_1944,In_2295,In_645);
nor U1945 (N_1945,In_1410,In_1839);
nor U1946 (N_1946,In_1124,In_2620);
nand U1947 (N_1947,In_641,In_2367);
or U1948 (N_1948,In_2542,In_2608);
and U1949 (N_1949,In_2845,In_1706);
or U1950 (N_1950,In_1875,In_2953);
or U1951 (N_1951,In_1192,In_1912);
and U1952 (N_1952,In_2800,In_1782);
and U1953 (N_1953,In_1814,In_1590);
or U1954 (N_1954,In_1711,In_2991);
and U1955 (N_1955,In_1146,In_1066);
and U1956 (N_1956,In_2013,In_2958);
nand U1957 (N_1957,In_1300,In_2732);
and U1958 (N_1958,In_1043,In_1898);
or U1959 (N_1959,In_1877,In_2140);
nand U1960 (N_1960,In_1971,In_2984);
and U1961 (N_1961,In_1577,In_2548);
and U1962 (N_1962,In_1242,In_1640);
and U1963 (N_1963,In_289,In_1088);
nand U1964 (N_1964,In_307,In_1428);
and U1965 (N_1965,In_1350,In_2638);
and U1966 (N_1966,In_580,In_1455);
nand U1967 (N_1967,In_1035,In_1698);
xor U1968 (N_1968,In_531,In_1653);
xor U1969 (N_1969,In_1616,In_545);
nand U1970 (N_1970,In_1103,In_1329);
and U1971 (N_1971,In_1995,In_1346);
nand U1972 (N_1972,In_123,In_132);
or U1973 (N_1973,In_2817,In_1777);
and U1974 (N_1974,In_1419,In_494);
and U1975 (N_1975,In_1609,In_570);
nor U1976 (N_1976,In_2418,In_1483);
nand U1977 (N_1977,In_925,In_2139);
nand U1978 (N_1978,In_1122,In_2460);
nand U1979 (N_1979,In_1990,In_114);
and U1980 (N_1980,In_1670,In_1680);
and U1981 (N_1981,In_1264,In_1563);
and U1982 (N_1982,In_1687,In_2002);
xor U1983 (N_1983,In_1956,In_1177);
nor U1984 (N_1984,In_2793,In_284);
nor U1985 (N_1985,In_1576,In_50);
nand U1986 (N_1986,In_1032,In_1030);
nor U1987 (N_1987,In_1033,In_287);
nor U1988 (N_1988,In_2642,In_1490);
nand U1989 (N_1989,In_297,In_2830);
and U1990 (N_1990,In_1089,In_2639);
nor U1991 (N_1991,In_1266,In_2672);
nand U1992 (N_1992,In_507,In_286);
nor U1993 (N_1993,In_2918,In_729);
and U1994 (N_1994,In_2187,In_910);
or U1995 (N_1995,In_2973,In_2562);
nor U1996 (N_1996,In_98,In_2996);
nor U1997 (N_1997,In_447,In_2924);
and U1998 (N_1998,In_48,In_140);
or U1999 (N_1999,In_2943,In_1669);
or U2000 (N_2000,In_2124,In_1606);
or U2001 (N_2001,In_2229,In_2784);
nand U2002 (N_2002,In_1278,In_2325);
nor U2003 (N_2003,In_754,In_409);
and U2004 (N_2004,In_2560,In_306);
or U2005 (N_2005,In_2326,In_2823);
nand U2006 (N_2006,In_2773,In_2639);
and U2007 (N_2007,In_2020,In_1901);
and U2008 (N_2008,In_709,In_232);
nand U2009 (N_2009,In_479,In_809);
or U2010 (N_2010,In_292,In_2408);
nand U2011 (N_2011,In_598,In_2053);
and U2012 (N_2012,In_2665,In_1900);
nor U2013 (N_2013,In_2637,In_1198);
or U2014 (N_2014,In_1760,In_2461);
or U2015 (N_2015,In_702,In_1568);
nand U2016 (N_2016,In_2851,In_400);
or U2017 (N_2017,In_2958,In_2959);
nor U2018 (N_2018,In_804,In_1296);
and U2019 (N_2019,In_1018,In_1132);
nor U2020 (N_2020,In_2853,In_804);
and U2021 (N_2021,In_1824,In_2394);
or U2022 (N_2022,In_2897,In_1062);
and U2023 (N_2023,In_1015,In_1373);
or U2024 (N_2024,In_2509,In_1951);
or U2025 (N_2025,In_2276,In_2168);
or U2026 (N_2026,In_2403,In_882);
nand U2027 (N_2027,In_1796,In_526);
nor U2028 (N_2028,In_2519,In_1016);
nand U2029 (N_2029,In_1483,In_2796);
nand U2030 (N_2030,In_906,In_1472);
xnor U2031 (N_2031,In_97,In_423);
nor U2032 (N_2032,In_849,In_869);
nor U2033 (N_2033,In_2791,In_2722);
nand U2034 (N_2034,In_1836,In_581);
or U2035 (N_2035,In_1991,In_2596);
nor U2036 (N_2036,In_1582,In_1549);
and U2037 (N_2037,In_1729,In_98);
nor U2038 (N_2038,In_1823,In_1932);
nand U2039 (N_2039,In_1726,In_1137);
nor U2040 (N_2040,In_2193,In_969);
nand U2041 (N_2041,In_1601,In_624);
and U2042 (N_2042,In_2685,In_1265);
nor U2043 (N_2043,In_21,In_1311);
and U2044 (N_2044,In_1112,In_2030);
and U2045 (N_2045,In_2081,In_837);
or U2046 (N_2046,In_2632,In_1996);
or U2047 (N_2047,In_2197,In_789);
or U2048 (N_2048,In_439,In_580);
and U2049 (N_2049,In_778,In_448);
or U2050 (N_2050,In_2591,In_1545);
nor U2051 (N_2051,In_2417,In_114);
and U2052 (N_2052,In_166,In_289);
xnor U2053 (N_2053,In_1243,In_1104);
nand U2054 (N_2054,In_1178,In_121);
nor U2055 (N_2055,In_1947,In_2316);
nor U2056 (N_2056,In_467,In_1182);
or U2057 (N_2057,In_985,In_2676);
xor U2058 (N_2058,In_94,In_1619);
or U2059 (N_2059,In_2033,In_2469);
nor U2060 (N_2060,In_1067,In_2405);
nand U2061 (N_2061,In_1309,In_1694);
and U2062 (N_2062,In_688,In_848);
and U2063 (N_2063,In_1620,In_2490);
and U2064 (N_2064,In_978,In_272);
nor U2065 (N_2065,In_2066,In_2124);
nand U2066 (N_2066,In_424,In_2798);
nand U2067 (N_2067,In_75,In_549);
xnor U2068 (N_2068,In_849,In_1353);
nand U2069 (N_2069,In_1085,In_2426);
xor U2070 (N_2070,In_31,In_1585);
nor U2071 (N_2071,In_1647,In_1302);
or U2072 (N_2072,In_394,In_1455);
nand U2073 (N_2073,In_2542,In_1110);
and U2074 (N_2074,In_885,In_151);
nor U2075 (N_2075,In_858,In_527);
or U2076 (N_2076,In_2768,In_2711);
nand U2077 (N_2077,In_577,In_2822);
and U2078 (N_2078,In_155,In_395);
xnor U2079 (N_2079,In_1813,In_926);
and U2080 (N_2080,In_2343,In_1181);
nor U2081 (N_2081,In_1021,In_827);
or U2082 (N_2082,In_1698,In_2760);
and U2083 (N_2083,In_517,In_2094);
or U2084 (N_2084,In_2388,In_1917);
nor U2085 (N_2085,In_2793,In_2058);
xor U2086 (N_2086,In_1253,In_969);
and U2087 (N_2087,In_1225,In_936);
or U2088 (N_2088,In_1876,In_2149);
and U2089 (N_2089,In_721,In_1872);
and U2090 (N_2090,In_198,In_2481);
nand U2091 (N_2091,In_1301,In_962);
nor U2092 (N_2092,In_2909,In_2032);
nor U2093 (N_2093,In_1986,In_2447);
and U2094 (N_2094,In_1412,In_910);
and U2095 (N_2095,In_1819,In_820);
nand U2096 (N_2096,In_2730,In_693);
or U2097 (N_2097,In_29,In_1165);
or U2098 (N_2098,In_2912,In_224);
and U2099 (N_2099,In_1454,In_2719);
and U2100 (N_2100,In_2685,In_467);
and U2101 (N_2101,In_863,In_930);
and U2102 (N_2102,In_2926,In_2854);
and U2103 (N_2103,In_2046,In_1753);
and U2104 (N_2104,In_2088,In_770);
or U2105 (N_2105,In_1706,In_1664);
nor U2106 (N_2106,In_2892,In_2400);
and U2107 (N_2107,In_1874,In_1597);
or U2108 (N_2108,In_2514,In_2724);
xor U2109 (N_2109,In_2306,In_622);
nor U2110 (N_2110,In_2168,In_1589);
nand U2111 (N_2111,In_2934,In_2947);
or U2112 (N_2112,In_784,In_2981);
nor U2113 (N_2113,In_1014,In_2443);
or U2114 (N_2114,In_795,In_1869);
nor U2115 (N_2115,In_432,In_652);
or U2116 (N_2116,In_574,In_2);
or U2117 (N_2117,In_1076,In_1650);
nor U2118 (N_2118,In_932,In_143);
nand U2119 (N_2119,In_1874,In_1647);
nand U2120 (N_2120,In_1197,In_1994);
and U2121 (N_2121,In_2492,In_2851);
or U2122 (N_2122,In_2231,In_2669);
nand U2123 (N_2123,In_2346,In_1641);
nor U2124 (N_2124,In_2091,In_60);
nand U2125 (N_2125,In_2176,In_1741);
nor U2126 (N_2126,In_711,In_2978);
nor U2127 (N_2127,In_2207,In_2407);
xor U2128 (N_2128,In_1606,In_1341);
and U2129 (N_2129,In_1696,In_888);
or U2130 (N_2130,In_629,In_2150);
nand U2131 (N_2131,In_887,In_565);
and U2132 (N_2132,In_2773,In_621);
and U2133 (N_2133,In_2055,In_1117);
and U2134 (N_2134,In_1574,In_96);
nor U2135 (N_2135,In_1858,In_2439);
or U2136 (N_2136,In_1455,In_1644);
xor U2137 (N_2137,In_1352,In_27);
xor U2138 (N_2138,In_2004,In_2296);
nand U2139 (N_2139,In_57,In_1093);
nor U2140 (N_2140,In_60,In_795);
nand U2141 (N_2141,In_1145,In_971);
xnor U2142 (N_2142,In_431,In_1042);
nand U2143 (N_2143,In_592,In_385);
and U2144 (N_2144,In_1085,In_2288);
nand U2145 (N_2145,In_2161,In_670);
or U2146 (N_2146,In_570,In_1652);
and U2147 (N_2147,In_1532,In_2519);
nand U2148 (N_2148,In_499,In_2566);
xor U2149 (N_2149,In_1710,In_2622);
or U2150 (N_2150,In_264,In_855);
xor U2151 (N_2151,In_823,In_2602);
xnor U2152 (N_2152,In_1707,In_1645);
nor U2153 (N_2153,In_2763,In_2216);
nand U2154 (N_2154,In_1434,In_1178);
or U2155 (N_2155,In_2730,In_2852);
nand U2156 (N_2156,In_575,In_914);
or U2157 (N_2157,In_196,In_2388);
or U2158 (N_2158,In_2646,In_2276);
nand U2159 (N_2159,In_600,In_92);
nor U2160 (N_2160,In_364,In_2237);
or U2161 (N_2161,In_2140,In_2141);
and U2162 (N_2162,In_2661,In_2688);
and U2163 (N_2163,In_1039,In_2963);
or U2164 (N_2164,In_2683,In_351);
or U2165 (N_2165,In_1737,In_1050);
and U2166 (N_2166,In_2283,In_2849);
and U2167 (N_2167,In_2181,In_1221);
nand U2168 (N_2168,In_109,In_1203);
nand U2169 (N_2169,In_2677,In_1615);
or U2170 (N_2170,In_721,In_630);
or U2171 (N_2171,In_2867,In_101);
nand U2172 (N_2172,In_1913,In_504);
nand U2173 (N_2173,In_479,In_956);
or U2174 (N_2174,In_2841,In_690);
or U2175 (N_2175,In_2162,In_311);
nor U2176 (N_2176,In_2577,In_1015);
nor U2177 (N_2177,In_1625,In_471);
nand U2178 (N_2178,In_1524,In_341);
and U2179 (N_2179,In_2811,In_123);
nor U2180 (N_2180,In_1268,In_2184);
and U2181 (N_2181,In_2642,In_2677);
or U2182 (N_2182,In_242,In_1300);
nand U2183 (N_2183,In_1008,In_10);
nor U2184 (N_2184,In_770,In_1983);
or U2185 (N_2185,In_1071,In_223);
nand U2186 (N_2186,In_2119,In_2665);
and U2187 (N_2187,In_2619,In_344);
nor U2188 (N_2188,In_2739,In_1698);
and U2189 (N_2189,In_2223,In_1212);
nand U2190 (N_2190,In_1809,In_843);
nor U2191 (N_2191,In_1000,In_2366);
nand U2192 (N_2192,In_1313,In_1763);
nor U2193 (N_2193,In_340,In_2125);
nor U2194 (N_2194,In_477,In_435);
or U2195 (N_2195,In_2367,In_1959);
and U2196 (N_2196,In_2772,In_794);
nand U2197 (N_2197,In_1276,In_2054);
and U2198 (N_2198,In_475,In_1136);
nor U2199 (N_2199,In_557,In_2156);
xnor U2200 (N_2200,In_183,In_1816);
and U2201 (N_2201,In_2017,In_129);
and U2202 (N_2202,In_1244,In_2967);
xor U2203 (N_2203,In_1495,In_2874);
nor U2204 (N_2204,In_2562,In_374);
xnor U2205 (N_2205,In_1396,In_1316);
nor U2206 (N_2206,In_1495,In_2050);
and U2207 (N_2207,In_1274,In_2543);
and U2208 (N_2208,In_457,In_1464);
nor U2209 (N_2209,In_2360,In_1202);
and U2210 (N_2210,In_2641,In_2464);
or U2211 (N_2211,In_1169,In_1849);
nand U2212 (N_2212,In_480,In_2568);
nor U2213 (N_2213,In_2905,In_2513);
nand U2214 (N_2214,In_831,In_640);
nor U2215 (N_2215,In_1229,In_2749);
and U2216 (N_2216,In_2995,In_1702);
and U2217 (N_2217,In_1875,In_2866);
nand U2218 (N_2218,In_2926,In_1436);
and U2219 (N_2219,In_1009,In_1544);
or U2220 (N_2220,In_1000,In_2674);
xor U2221 (N_2221,In_2860,In_2194);
nor U2222 (N_2222,In_1594,In_2373);
nor U2223 (N_2223,In_865,In_1620);
xor U2224 (N_2224,In_2223,In_32);
nor U2225 (N_2225,In_738,In_48);
or U2226 (N_2226,In_417,In_71);
or U2227 (N_2227,In_1139,In_2691);
and U2228 (N_2228,In_1163,In_473);
nand U2229 (N_2229,In_2734,In_1247);
nor U2230 (N_2230,In_2860,In_1794);
nand U2231 (N_2231,In_1015,In_2648);
nor U2232 (N_2232,In_742,In_377);
nor U2233 (N_2233,In_56,In_1425);
and U2234 (N_2234,In_2224,In_2102);
or U2235 (N_2235,In_2475,In_2337);
nand U2236 (N_2236,In_2067,In_1386);
nand U2237 (N_2237,In_2109,In_436);
nor U2238 (N_2238,In_1600,In_851);
nand U2239 (N_2239,In_1572,In_2739);
nor U2240 (N_2240,In_2526,In_1838);
or U2241 (N_2241,In_1535,In_962);
nor U2242 (N_2242,In_2881,In_823);
xor U2243 (N_2243,In_2794,In_788);
and U2244 (N_2244,In_2465,In_728);
or U2245 (N_2245,In_1484,In_1245);
xnor U2246 (N_2246,In_33,In_752);
xnor U2247 (N_2247,In_1952,In_486);
nand U2248 (N_2248,In_2932,In_2770);
nand U2249 (N_2249,In_2666,In_1470);
or U2250 (N_2250,In_2118,In_2277);
nor U2251 (N_2251,In_1611,In_2288);
or U2252 (N_2252,In_1358,In_1518);
xor U2253 (N_2253,In_1440,In_2248);
nand U2254 (N_2254,In_1433,In_574);
or U2255 (N_2255,In_2575,In_1856);
nor U2256 (N_2256,In_997,In_11);
nand U2257 (N_2257,In_2239,In_2402);
or U2258 (N_2258,In_844,In_2913);
or U2259 (N_2259,In_1145,In_2540);
nor U2260 (N_2260,In_1863,In_1348);
nor U2261 (N_2261,In_267,In_1341);
and U2262 (N_2262,In_790,In_2863);
nor U2263 (N_2263,In_1415,In_1327);
xor U2264 (N_2264,In_1627,In_2699);
and U2265 (N_2265,In_2823,In_1180);
nand U2266 (N_2266,In_2385,In_1714);
nand U2267 (N_2267,In_2493,In_1657);
or U2268 (N_2268,In_1681,In_2393);
nor U2269 (N_2269,In_1923,In_2097);
xor U2270 (N_2270,In_1013,In_1757);
or U2271 (N_2271,In_1567,In_1467);
or U2272 (N_2272,In_1048,In_2680);
nor U2273 (N_2273,In_2353,In_383);
nor U2274 (N_2274,In_1994,In_777);
nand U2275 (N_2275,In_477,In_1912);
nor U2276 (N_2276,In_1575,In_14);
and U2277 (N_2277,In_122,In_2621);
xnor U2278 (N_2278,In_2490,In_1465);
nor U2279 (N_2279,In_1387,In_341);
xor U2280 (N_2280,In_2196,In_610);
nand U2281 (N_2281,In_833,In_142);
or U2282 (N_2282,In_2507,In_1600);
and U2283 (N_2283,In_1462,In_776);
xor U2284 (N_2284,In_1633,In_1375);
and U2285 (N_2285,In_243,In_235);
nor U2286 (N_2286,In_971,In_2838);
and U2287 (N_2287,In_2066,In_1951);
and U2288 (N_2288,In_2381,In_2138);
nor U2289 (N_2289,In_585,In_141);
nor U2290 (N_2290,In_857,In_421);
and U2291 (N_2291,In_2640,In_683);
nand U2292 (N_2292,In_473,In_1152);
or U2293 (N_2293,In_1341,In_2271);
xnor U2294 (N_2294,In_2926,In_2781);
xor U2295 (N_2295,In_2027,In_2999);
nor U2296 (N_2296,In_54,In_1968);
nor U2297 (N_2297,In_1032,In_762);
nor U2298 (N_2298,In_2621,In_1852);
and U2299 (N_2299,In_12,In_1484);
and U2300 (N_2300,In_835,In_489);
or U2301 (N_2301,In_1984,In_1466);
nand U2302 (N_2302,In_1607,In_991);
or U2303 (N_2303,In_169,In_2683);
and U2304 (N_2304,In_1704,In_466);
nor U2305 (N_2305,In_1114,In_902);
or U2306 (N_2306,In_68,In_2252);
nand U2307 (N_2307,In_2053,In_644);
and U2308 (N_2308,In_1036,In_1465);
xor U2309 (N_2309,In_284,In_2517);
or U2310 (N_2310,In_1011,In_1007);
and U2311 (N_2311,In_1809,In_326);
nor U2312 (N_2312,In_1440,In_2601);
or U2313 (N_2313,In_874,In_2093);
nor U2314 (N_2314,In_1384,In_448);
xnor U2315 (N_2315,In_1961,In_1858);
nand U2316 (N_2316,In_2239,In_1221);
or U2317 (N_2317,In_1629,In_2028);
and U2318 (N_2318,In_953,In_2150);
xor U2319 (N_2319,In_302,In_1540);
and U2320 (N_2320,In_2083,In_609);
and U2321 (N_2321,In_1078,In_1881);
nand U2322 (N_2322,In_992,In_528);
nor U2323 (N_2323,In_751,In_1117);
and U2324 (N_2324,In_1651,In_233);
or U2325 (N_2325,In_882,In_11);
xor U2326 (N_2326,In_953,In_655);
xnor U2327 (N_2327,In_2463,In_2047);
or U2328 (N_2328,In_2367,In_2142);
nand U2329 (N_2329,In_502,In_482);
or U2330 (N_2330,In_2984,In_1515);
or U2331 (N_2331,In_2579,In_2720);
and U2332 (N_2332,In_1203,In_2298);
nor U2333 (N_2333,In_1428,In_2884);
nand U2334 (N_2334,In_852,In_576);
or U2335 (N_2335,In_1893,In_53);
nor U2336 (N_2336,In_2468,In_2800);
or U2337 (N_2337,In_792,In_895);
xor U2338 (N_2338,In_1681,In_2565);
or U2339 (N_2339,In_127,In_1424);
nand U2340 (N_2340,In_1514,In_1037);
and U2341 (N_2341,In_2788,In_42);
and U2342 (N_2342,In_2332,In_165);
nor U2343 (N_2343,In_1142,In_809);
or U2344 (N_2344,In_2348,In_2621);
and U2345 (N_2345,In_1891,In_1535);
or U2346 (N_2346,In_1762,In_204);
nor U2347 (N_2347,In_1710,In_2884);
nand U2348 (N_2348,In_1008,In_2403);
and U2349 (N_2349,In_1979,In_1803);
nor U2350 (N_2350,In_1788,In_768);
and U2351 (N_2351,In_1320,In_2654);
nand U2352 (N_2352,In_643,In_1108);
xor U2353 (N_2353,In_1069,In_2947);
and U2354 (N_2354,In_160,In_2469);
and U2355 (N_2355,In_1757,In_2378);
or U2356 (N_2356,In_618,In_329);
xor U2357 (N_2357,In_1382,In_1842);
and U2358 (N_2358,In_278,In_2388);
nand U2359 (N_2359,In_2979,In_2577);
and U2360 (N_2360,In_2509,In_1081);
and U2361 (N_2361,In_2639,In_2719);
nor U2362 (N_2362,In_1754,In_1066);
or U2363 (N_2363,In_1296,In_717);
nand U2364 (N_2364,In_1527,In_2806);
nor U2365 (N_2365,In_2963,In_2962);
and U2366 (N_2366,In_1944,In_806);
xnor U2367 (N_2367,In_2636,In_2622);
or U2368 (N_2368,In_2520,In_1856);
nor U2369 (N_2369,In_511,In_1068);
nand U2370 (N_2370,In_2209,In_1598);
nand U2371 (N_2371,In_1823,In_75);
nand U2372 (N_2372,In_751,In_57);
xnor U2373 (N_2373,In_2239,In_2425);
nor U2374 (N_2374,In_2423,In_2141);
and U2375 (N_2375,In_654,In_700);
nor U2376 (N_2376,In_1516,In_706);
and U2377 (N_2377,In_579,In_2378);
and U2378 (N_2378,In_866,In_144);
and U2379 (N_2379,In_926,In_1326);
nor U2380 (N_2380,In_2751,In_531);
and U2381 (N_2381,In_1500,In_859);
nand U2382 (N_2382,In_1676,In_1612);
and U2383 (N_2383,In_209,In_2562);
and U2384 (N_2384,In_2590,In_2849);
nor U2385 (N_2385,In_2008,In_986);
and U2386 (N_2386,In_279,In_2123);
nor U2387 (N_2387,In_2655,In_1127);
nor U2388 (N_2388,In_893,In_1323);
and U2389 (N_2389,In_217,In_1538);
nor U2390 (N_2390,In_1526,In_1357);
and U2391 (N_2391,In_228,In_1160);
and U2392 (N_2392,In_896,In_2322);
and U2393 (N_2393,In_2867,In_42);
and U2394 (N_2394,In_1539,In_247);
nor U2395 (N_2395,In_2456,In_976);
or U2396 (N_2396,In_2603,In_2757);
or U2397 (N_2397,In_846,In_15);
and U2398 (N_2398,In_2674,In_2024);
xnor U2399 (N_2399,In_248,In_2136);
and U2400 (N_2400,In_643,In_2692);
and U2401 (N_2401,In_2266,In_826);
xnor U2402 (N_2402,In_2219,In_1878);
or U2403 (N_2403,In_1866,In_1494);
nor U2404 (N_2404,In_595,In_855);
nand U2405 (N_2405,In_2966,In_968);
xor U2406 (N_2406,In_110,In_2854);
nand U2407 (N_2407,In_333,In_2892);
and U2408 (N_2408,In_1695,In_2360);
and U2409 (N_2409,In_1860,In_1086);
nor U2410 (N_2410,In_2281,In_2312);
nand U2411 (N_2411,In_2258,In_314);
nor U2412 (N_2412,In_855,In_777);
nor U2413 (N_2413,In_615,In_1252);
xnor U2414 (N_2414,In_593,In_259);
nor U2415 (N_2415,In_1760,In_2912);
nor U2416 (N_2416,In_2131,In_1964);
or U2417 (N_2417,In_2749,In_799);
nor U2418 (N_2418,In_1083,In_1779);
xnor U2419 (N_2419,In_457,In_1997);
nor U2420 (N_2420,In_1867,In_2860);
xor U2421 (N_2421,In_1859,In_2782);
nand U2422 (N_2422,In_1555,In_911);
nor U2423 (N_2423,In_2156,In_1514);
and U2424 (N_2424,In_686,In_899);
or U2425 (N_2425,In_926,In_1109);
or U2426 (N_2426,In_1814,In_1833);
nor U2427 (N_2427,In_1229,In_2690);
nor U2428 (N_2428,In_1028,In_1088);
and U2429 (N_2429,In_1431,In_1555);
or U2430 (N_2430,In_2371,In_2672);
nor U2431 (N_2431,In_2494,In_629);
and U2432 (N_2432,In_55,In_1261);
or U2433 (N_2433,In_1724,In_834);
nand U2434 (N_2434,In_552,In_2165);
or U2435 (N_2435,In_2128,In_1142);
nor U2436 (N_2436,In_1859,In_1631);
or U2437 (N_2437,In_2785,In_2303);
nor U2438 (N_2438,In_2804,In_2511);
and U2439 (N_2439,In_1458,In_1367);
and U2440 (N_2440,In_2705,In_1972);
or U2441 (N_2441,In_2090,In_2674);
and U2442 (N_2442,In_366,In_385);
and U2443 (N_2443,In_1028,In_730);
nor U2444 (N_2444,In_2059,In_1299);
nand U2445 (N_2445,In_2955,In_2872);
and U2446 (N_2446,In_1025,In_749);
and U2447 (N_2447,In_1677,In_176);
nor U2448 (N_2448,In_1741,In_1251);
xnor U2449 (N_2449,In_739,In_2453);
nor U2450 (N_2450,In_2901,In_17);
nand U2451 (N_2451,In_2093,In_2585);
xor U2452 (N_2452,In_2287,In_2621);
and U2453 (N_2453,In_2101,In_943);
and U2454 (N_2454,In_2470,In_2688);
or U2455 (N_2455,In_1623,In_1943);
and U2456 (N_2456,In_1393,In_428);
and U2457 (N_2457,In_990,In_210);
nor U2458 (N_2458,In_1352,In_1357);
or U2459 (N_2459,In_2757,In_47);
and U2460 (N_2460,In_2411,In_2068);
xor U2461 (N_2461,In_225,In_615);
and U2462 (N_2462,In_1270,In_595);
xnor U2463 (N_2463,In_1777,In_227);
xnor U2464 (N_2464,In_1366,In_2176);
and U2465 (N_2465,In_2501,In_2075);
and U2466 (N_2466,In_464,In_2130);
nand U2467 (N_2467,In_425,In_1935);
nor U2468 (N_2468,In_363,In_2324);
nand U2469 (N_2469,In_1864,In_724);
nor U2470 (N_2470,In_201,In_1349);
xor U2471 (N_2471,In_2462,In_1765);
nand U2472 (N_2472,In_2648,In_2530);
nand U2473 (N_2473,In_904,In_2942);
or U2474 (N_2474,In_2651,In_475);
or U2475 (N_2475,In_2169,In_928);
and U2476 (N_2476,In_2999,In_1486);
and U2477 (N_2477,In_99,In_2186);
or U2478 (N_2478,In_2065,In_1285);
nand U2479 (N_2479,In_1219,In_2604);
and U2480 (N_2480,In_1561,In_2880);
nand U2481 (N_2481,In_2200,In_420);
and U2482 (N_2482,In_2396,In_1506);
nor U2483 (N_2483,In_493,In_913);
nor U2484 (N_2484,In_2632,In_771);
nor U2485 (N_2485,In_2150,In_905);
or U2486 (N_2486,In_278,In_1815);
or U2487 (N_2487,In_1880,In_910);
nand U2488 (N_2488,In_395,In_2474);
nor U2489 (N_2489,In_334,In_866);
nor U2490 (N_2490,In_1784,In_150);
or U2491 (N_2491,In_915,In_1763);
nand U2492 (N_2492,In_1899,In_2466);
nor U2493 (N_2493,In_2907,In_388);
xor U2494 (N_2494,In_1852,In_2101);
or U2495 (N_2495,In_930,In_236);
nor U2496 (N_2496,In_2760,In_500);
nor U2497 (N_2497,In_552,In_2980);
nand U2498 (N_2498,In_244,In_1047);
or U2499 (N_2499,In_236,In_224);
or U2500 (N_2500,In_480,In_97);
or U2501 (N_2501,In_716,In_966);
or U2502 (N_2502,In_2194,In_2110);
and U2503 (N_2503,In_1149,In_220);
and U2504 (N_2504,In_93,In_2877);
nor U2505 (N_2505,In_600,In_2020);
nor U2506 (N_2506,In_588,In_1272);
nand U2507 (N_2507,In_1771,In_1904);
nand U2508 (N_2508,In_237,In_2287);
nand U2509 (N_2509,In_1391,In_1952);
and U2510 (N_2510,In_422,In_824);
xor U2511 (N_2511,In_1594,In_1399);
nor U2512 (N_2512,In_514,In_306);
nor U2513 (N_2513,In_1122,In_2105);
and U2514 (N_2514,In_671,In_1193);
and U2515 (N_2515,In_504,In_435);
and U2516 (N_2516,In_2779,In_2772);
xnor U2517 (N_2517,In_1706,In_2425);
nand U2518 (N_2518,In_1962,In_2220);
or U2519 (N_2519,In_720,In_2171);
or U2520 (N_2520,In_2875,In_2365);
or U2521 (N_2521,In_262,In_2199);
or U2522 (N_2522,In_912,In_814);
nor U2523 (N_2523,In_1806,In_1746);
xor U2524 (N_2524,In_2364,In_2210);
and U2525 (N_2525,In_553,In_557);
nand U2526 (N_2526,In_2268,In_2066);
and U2527 (N_2527,In_1492,In_1709);
or U2528 (N_2528,In_1077,In_591);
nand U2529 (N_2529,In_413,In_981);
nand U2530 (N_2530,In_952,In_1950);
or U2531 (N_2531,In_1388,In_2579);
or U2532 (N_2532,In_261,In_1500);
xor U2533 (N_2533,In_1811,In_358);
nor U2534 (N_2534,In_7,In_1390);
and U2535 (N_2535,In_665,In_301);
nand U2536 (N_2536,In_1270,In_1000);
nor U2537 (N_2537,In_1310,In_741);
nand U2538 (N_2538,In_726,In_268);
nor U2539 (N_2539,In_2595,In_1733);
nor U2540 (N_2540,In_1148,In_1297);
or U2541 (N_2541,In_2385,In_1377);
xnor U2542 (N_2542,In_1117,In_2358);
or U2543 (N_2543,In_1387,In_1207);
nand U2544 (N_2544,In_206,In_2252);
nand U2545 (N_2545,In_491,In_2429);
and U2546 (N_2546,In_1583,In_639);
nor U2547 (N_2547,In_2211,In_1083);
nor U2548 (N_2548,In_2844,In_1975);
nor U2549 (N_2549,In_1029,In_3);
xor U2550 (N_2550,In_1704,In_959);
xnor U2551 (N_2551,In_342,In_1932);
nor U2552 (N_2552,In_2392,In_2584);
nor U2553 (N_2553,In_2587,In_1001);
and U2554 (N_2554,In_1306,In_1952);
and U2555 (N_2555,In_1804,In_2488);
nand U2556 (N_2556,In_2300,In_2638);
xor U2557 (N_2557,In_2398,In_2372);
nor U2558 (N_2558,In_2814,In_1255);
nor U2559 (N_2559,In_162,In_307);
nor U2560 (N_2560,In_832,In_268);
nand U2561 (N_2561,In_1459,In_735);
or U2562 (N_2562,In_1781,In_2319);
nand U2563 (N_2563,In_2252,In_1201);
or U2564 (N_2564,In_2777,In_1990);
and U2565 (N_2565,In_2362,In_418);
nor U2566 (N_2566,In_1186,In_2408);
nand U2567 (N_2567,In_2108,In_931);
xor U2568 (N_2568,In_184,In_1378);
and U2569 (N_2569,In_1307,In_2853);
nor U2570 (N_2570,In_1682,In_846);
xnor U2571 (N_2571,In_2896,In_2216);
or U2572 (N_2572,In_2083,In_1056);
or U2573 (N_2573,In_103,In_1218);
nand U2574 (N_2574,In_1412,In_2708);
or U2575 (N_2575,In_2732,In_2669);
or U2576 (N_2576,In_1254,In_2812);
and U2577 (N_2577,In_1714,In_968);
and U2578 (N_2578,In_1044,In_2241);
or U2579 (N_2579,In_2517,In_2974);
or U2580 (N_2580,In_2716,In_2478);
or U2581 (N_2581,In_2508,In_979);
and U2582 (N_2582,In_1920,In_2672);
and U2583 (N_2583,In_2611,In_525);
and U2584 (N_2584,In_2138,In_1995);
or U2585 (N_2585,In_1003,In_862);
and U2586 (N_2586,In_97,In_1694);
and U2587 (N_2587,In_122,In_974);
nor U2588 (N_2588,In_1076,In_2634);
and U2589 (N_2589,In_945,In_1616);
nand U2590 (N_2590,In_1045,In_1256);
nor U2591 (N_2591,In_43,In_228);
nand U2592 (N_2592,In_911,In_1571);
nor U2593 (N_2593,In_2259,In_1);
xor U2594 (N_2594,In_2022,In_956);
and U2595 (N_2595,In_2621,In_736);
and U2596 (N_2596,In_2877,In_47);
and U2597 (N_2597,In_1596,In_1512);
and U2598 (N_2598,In_2607,In_1705);
and U2599 (N_2599,In_615,In_2220);
nand U2600 (N_2600,In_1181,In_953);
and U2601 (N_2601,In_1710,In_2182);
and U2602 (N_2602,In_1940,In_1493);
nand U2603 (N_2603,In_2441,In_1391);
and U2604 (N_2604,In_1511,In_1288);
nor U2605 (N_2605,In_760,In_2089);
or U2606 (N_2606,In_757,In_956);
or U2607 (N_2607,In_898,In_1859);
nand U2608 (N_2608,In_737,In_2147);
or U2609 (N_2609,In_2530,In_1330);
and U2610 (N_2610,In_2189,In_1598);
nor U2611 (N_2611,In_527,In_2549);
and U2612 (N_2612,In_24,In_114);
nor U2613 (N_2613,In_2901,In_1983);
and U2614 (N_2614,In_205,In_1494);
or U2615 (N_2615,In_906,In_56);
nor U2616 (N_2616,In_1107,In_2075);
nand U2617 (N_2617,In_273,In_2289);
nor U2618 (N_2618,In_1168,In_1656);
nor U2619 (N_2619,In_704,In_2321);
xor U2620 (N_2620,In_1850,In_1707);
nand U2621 (N_2621,In_2907,In_1304);
nand U2622 (N_2622,In_2591,In_2564);
and U2623 (N_2623,In_2613,In_1799);
or U2624 (N_2624,In_874,In_2152);
nand U2625 (N_2625,In_1970,In_2201);
xnor U2626 (N_2626,In_551,In_182);
nor U2627 (N_2627,In_2773,In_2181);
or U2628 (N_2628,In_90,In_1089);
and U2629 (N_2629,In_1716,In_1315);
nand U2630 (N_2630,In_945,In_1481);
nand U2631 (N_2631,In_1469,In_2163);
nand U2632 (N_2632,In_2981,In_1864);
nand U2633 (N_2633,In_330,In_1975);
nand U2634 (N_2634,In_2682,In_1727);
nand U2635 (N_2635,In_211,In_1043);
nand U2636 (N_2636,In_1623,In_147);
nand U2637 (N_2637,In_2340,In_228);
or U2638 (N_2638,In_1430,In_2091);
nand U2639 (N_2639,In_123,In_1253);
nand U2640 (N_2640,In_163,In_524);
or U2641 (N_2641,In_2528,In_2558);
nor U2642 (N_2642,In_640,In_2160);
nor U2643 (N_2643,In_146,In_1318);
and U2644 (N_2644,In_728,In_1147);
xnor U2645 (N_2645,In_877,In_2362);
nand U2646 (N_2646,In_1751,In_2121);
nand U2647 (N_2647,In_909,In_2151);
and U2648 (N_2648,In_108,In_1026);
or U2649 (N_2649,In_1281,In_2586);
nand U2650 (N_2650,In_1456,In_1559);
nand U2651 (N_2651,In_2326,In_2367);
and U2652 (N_2652,In_2693,In_2111);
nand U2653 (N_2653,In_903,In_1444);
nor U2654 (N_2654,In_1626,In_2664);
and U2655 (N_2655,In_842,In_57);
and U2656 (N_2656,In_2173,In_2406);
and U2657 (N_2657,In_1338,In_1770);
nand U2658 (N_2658,In_2617,In_2696);
and U2659 (N_2659,In_1721,In_1487);
or U2660 (N_2660,In_47,In_2467);
or U2661 (N_2661,In_1476,In_2249);
nor U2662 (N_2662,In_1211,In_2788);
and U2663 (N_2663,In_1190,In_1068);
nor U2664 (N_2664,In_954,In_1519);
nor U2665 (N_2665,In_1218,In_1940);
xnor U2666 (N_2666,In_64,In_1395);
and U2667 (N_2667,In_738,In_2026);
and U2668 (N_2668,In_2422,In_1683);
nand U2669 (N_2669,In_288,In_1383);
nand U2670 (N_2670,In_2621,In_1257);
or U2671 (N_2671,In_1908,In_1342);
nor U2672 (N_2672,In_1985,In_249);
or U2673 (N_2673,In_1779,In_1086);
or U2674 (N_2674,In_854,In_2654);
nor U2675 (N_2675,In_2734,In_189);
nor U2676 (N_2676,In_2062,In_2575);
and U2677 (N_2677,In_2272,In_487);
nor U2678 (N_2678,In_1105,In_2357);
nand U2679 (N_2679,In_1373,In_1844);
and U2680 (N_2680,In_2255,In_2201);
nor U2681 (N_2681,In_541,In_2328);
and U2682 (N_2682,In_570,In_1551);
nand U2683 (N_2683,In_951,In_1949);
xor U2684 (N_2684,In_865,In_1539);
xnor U2685 (N_2685,In_143,In_717);
nor U2686 (N_2686,In_886,In_612);
nor U2687 (N_2687,In_1834,In_1871);
and U2688 (N_2688,In_1878,In_2767);
nor U2689 (N_2689,In_849,In_273);
or U2690 (N_2690,In_1418,In_256);
nor U2691 (N_2691,In_706,In_968);
and U2692 (N_2692,In_1534,In_2978);
xor U2693 (N_2693,In_954,In_1733);
and U2694 (N_2694,In_1060,In_487);
nor U2695 (N_2695,In_1624,In_1678);
or U2696 (N_2696,In_523,In_274);
or U2697 (N_2697,In_1363,In_32);
and U2698 (N_2698,In_321,In_576);
or U2699 (N_2699,In_2527,In_352);
xor U2700 (N_2700,In_1464,In_1347);
nand U2701 (N_2701,In_2556,In_1812);
or U2702 (N_2702,In_1792,In_2182);
and U2703 (N_2703,In_2722,In_516);
nor U2704 (N_2704,In_2855,In_306);
nand U2705 (N_2705,In_1448,In_789);
nand U2706 (N_2706,In_2532,In_902);
and U2707 (N_2707,In_1706,In_1054);
nor U2708 (N_2708,In_35,In_1961);
and U2709 (N_2709,In_2053,In_908);
nor U2710 (N_2710,In_233,In_1215);
nand U2711 (N_2711,In_2697,In_1567);
nand U2712 (N_2712,In_1787,In_1867);
or U2713 (N_2713,In_1239,In_858);
and U2714 (N_2714,In_12,In_907);
nor U2715 (N_2715,In_1382,In_401);
and U2716 (N_2716,In_206,In_1930);
nor U2717 (N_2717,In_2588,In_177);
or U2718 (N_2718,In_2054,In_2904);
nand U2719 (N_2719,In_1069,In_2198);
or U2720 (N_2720,In_946,In_796);
and U2721 (N_2721,In_2765,In_2282);
nor U2722 (N_2722,In_53,In_2894);
or U2723 (N_2723,In_681,In_310);
and U2724 (N_2724,In_1590,In_2266);
nor U2725 (N_2725,In_1998,In_163);
or U2726 (N_2726,In_2403,In_505);
or U2727 (N_2727,In_1577,In_1912);
and U2728 (N_2728,In_2480,In_447);
and U2729 (N_2729,In_2312,In_2555);
xnor U2730 (N_2730,In_1031,In_2860);
nand U2731 (N_2731,In_2787,In_1859);
nor U2732 (N_2732,In_2961,In_1765);
and U2733 (N_2733,In_385,In_1552);
nor U2734 (N_2734,In_231,In_2921);
nand U2735 (N_2735,In_2232,In_765);
nand U2736 (N_2736,In_362,In_835);
nand U2737 (N_2737,In_2178,In_2171);
and U2738 (N_2738,In_2068,In_1688);
or U2739 (N_2739,In_300,In_178);
and U2740 (N_2740,In_754,In_2375);
and U2741 (N_2741,In_2642,In_1507);
or U2742 (N_2742,In_2789,In_699);
or U2743 (N_2743,In_2846,In_59);
and U2744 (N_2744,In_1109,In_1339);
or U2745 (N_2745,In_219,In_85);
or U2746 (N_2746,In_2360,In_2643);
and U2747 (N_2747,In_2412,In_2234);
xor U2748 (N_2748,In_881,In_1751);
or U2749 (N_2749,In_387,In_863);
or U2750 (N_2750,In_2919,In_801);
nor U2751 (N_2751,In_1284,In_276);
and U2752 (N_2752,In_1578,In_2337);
xor U2753 (N_2753,In_217,In_893);
or U2754 (N_2754,In_2822,In_913);
or U2755 (N_2755,In_1778,In_2143);
nor U2756 (N_2756,In_119,In_650);
nor U2757 (N_2757,In_2248,In_832);
or U2758 (N_2758,In_614,In_203);
xor U2759 (N_2759,In_87,In_2975);
nand U2760 (N_2760,In_1253,In_1538);
and U2761 (N_2761,In_1313,In_197);
or U2762 (N_2762,In_2875,In_2644);
and U2763 (N_2763,In_598,In_1319);
nor U2764 (N_2764,In_1738,In_631);
nor U2765 (N_2765,In_1641,In_2150);
xnor U2766 (N_2766,In_1983,In_1373);
nand U2767 (N_2767,In_594,In_2519);
and U2768 (N_2768,In_2838,In_87);
nand U2769 (N_2769,In_911,In_891);
nand U2770 (N_2770,In_2918,In_2319);
nand U2771 (N_2771,In_378,In_1170);
nor U2772 (N_2772,In_2307,In_1808);
nand U2773 (N_2773,In_601,In_560);
nor U2774 (N_2774,In_2267,In_1349);
xor U2775 (N_2775,In_537,In_1081);
nand U2776 (N_2776,In_841,In_111);
nor U2777 (N_2777,In_349,In_2071);
and U2778 (N_2778,In_2976,In_1025);
nor U2779 (N_2779,In_2678,In_1327);
and U2780 (N_2780,In_2734,In_1378);
nor U2781 (N_2781,In_1483,In_1582);
xor U2782 (N_2782,In_2761,In_1397);
nor U2783 (N_2783,In_2100,In_433);
or U2784 (N_2784,In_880,In_1814);
nand U2785 (N_2785,In_295,In_2448);
nand U2786 (N_2786,In_24,In_1360);
xnor U2787 (N_2787,In_1870,In_1708);
xnor U2788 (N_2788,In_944,In_2728);
and U2789 (N_2789,In_952,In_1559);
or U2790 (N_2790,In_1126,In_2514);
nand U2791 (N_2791,In_2974,In_304);
nor U2792 (N_2792,In_1486,In_2884);
nand U2793 (N_2793,In_1019,In_2289);
and U2794 (N_2794,In_392,In_2658);
nand U2795 (N_2795,In_2592,In_2641);
nand U2796 (N_2796,In_2131,In_2178);
nand U2797 (N_2797,In_2319,In_410);
nand U2798 (N_2798,In_1284,In_133);
and U2799 (N_2799,In_2390,In_1317);
nor U2800 (N_2800,In_2817,In_2478);
and U2801 (N_2801,In_1227,In_2983);
or U2802 (N_2802,In_618,In_2143);
nand U2803 (N_2803,In_426,In_1038);
nor U2804 (N_2804,In_1169,In_148);
nor U2805 (N_2805,In_2969,In_2459);
nand U2806 (N_2806,In_2926,In_738);
or U2807 (N_2807,In_2618,In_681);
xnor U2808 (N_2808,In_1990,In_1746);
xnor U2809 (N_2809,In_1337,In_68);
nor U2810 (N_2810,In_2271,In_2459);
nand U2811 (N_2811,In_2719,In_2961);
nor U2812 (N_2812,In_1906,In_2764);
xor U2813 (N_2813,In_815,In_2279);
or U2814 (N_2814,In_975,In_2899);
and U2815 (N_2815,In_1141,In_1827);
or U2816 (N_2816,In_2145,In_2368);
nor U2817 (N_2817,In_456,In_1424);
nor U2818 (N_2818,In_1832,In_2248);
xnor U2819 (N_2819,In_1438,In_2993);
or U2820 (N_2820,In_935,In_2742);
and U2821 (N_2821,In_2292,In_591);
or U2822 (N_2822,In_1707,In_2936);
nand U2823 (N_2823,In_488,In_1970);
nand U2824 (N_2824,In_216,In_520);
nand U2825 (N_2825,In_2522,In_1799);
or U2826 (N_2826,In_880,In_1433);
or U2827 (N_2827,In_2849,In_2383);
or U2828 (N_2828,In_179,In_2110);
nor U2829 (N_2829,In_1025,In_111);
xnor U2830 (N_2830,In_2820,In_1030);
nor U2831 (N_2831,In_1774,In_2944);
nor U2832 (N_2832,In_1367,In_303);
nand U2833 (N_2833,In_2168,In_1099);
nand U2834 (N_2834,In_1287,In_96);
or U2835 (N_2835,In_943,In_261);
and U2836 (N_2836,In_1321,In_528);
xor U2837 (N_2837,In_1897,In_770);
nand U2838 (N_2838,In_2627,In_846);
nand U2839 (N_2839,In_563,In_2577);
xor U2840 (N_2840,In_2507,In_1045);
nor U2841 (N_2841,In_2498,In_2724);
or U2842 (N_2842,In_2159,In_1646);
nor U2843 (N_2843,In_2048,In_396);
or U2844 (N_2844,In_377,In_2041);
and U2845 (N_2845,In_226,In_1097);
or U2846 (N_2846,In_1406,In_95);
nor U2847 (N_2847,In_1258,In_2767);
nand U2848 (N_2848,In_1816,In_1490);
or U2849 (N_2849,In_458,In_113);
or U2850 (N_2850,In_1846,In_2873);
nor U2851 (N_2851,In_195,In_1966);
or U2852 (N_2852,In_2322,In_1642);
or U2853 (N_2853,In_2113,In_917);
or U2854 (N_2854,In_1407,In_154);
nand U2855 (N_2855,In_1275,In_2548);
or U2856 (N_2856,In_2953,In_1572);
xnor U2857 (N_2857,In_2627,In_831);
and U2858 (N_2858,In_2012,In_2369);
or U2859 (N_2859,In_113,In_1339);
nor U2860 (N_2860,In_2989,In_2069);
or U2861 (N_2861,In_1486,In_2313);
nand U2862 (N_2862,In_2616,In_342);
nor U2863 (N_2863,In_2137,In_1847);
and U2864 (N_2864,In_145,In_72);
and U2865 (N_2865,In_2469,In_2835);
and U2866 (N_2866,In_2939,In_376);
nor U2867 (N_2867,In_965,In_18);
xnor U2868 (N_2868,In_354,In_2573);
nor U2869 (N_2869,In_417,In_2449);
nand U2870 (N_2870,In_346,In_2820);
nand U2871 (N_2871,In_625,In_2217);
or U2872 (N_2872,In_69,In_1926);
or U2873 (N_2873,In_765,In_2762);
xnor U2874 (N_2874,In_2205,In_2591);
nand U2875 (N_2875,In_1662,In_1771);
xor U2876 (N_2876,In_941,In_1957);
nand U2877 (N_2877,In_580,In_1571);
nand U2878 (N_2878,In_2853,In_4);
nand U2879 (N_2879,In_1704,In_1209);
or U2880 (N_2880,In_665,In_1764);
or U2881 (N_2881,In_2247,In_630);
or U2882 (N_2882,In_2141,In_2298);
nor U2883 (N_2883,In_1056,In_936);
and U2884 (N_2884,In_745,In_917);
or U2885 (N_2885,In_1066,In_1157);
nand U2886 (N_2886,In_426,In_1602);
xnor U2887 (N_2887,In_1180,In_374);
nand U2888 (N_2888,In_1032,In_2365);
and U2889 (N_2889,In_2154,In_1919);
nand U2890 (N_2890,In_2670,In_1682);
or U2891 (N_2891,In_858,In_2423);
or U2892 (N_2892,In_1280,In_2310);
nor U2893 (N_2893,In_1487,In_99);
and U2894 (N_2894,In_910,In_2183);
or U2895 (N_2895,In_2277,In_2599);
nor U2896 (N_2896,In_1199,In_770);
or U2897 (N_2897,In_857,In_1769);
nand U2898 (N_2898,In_2968,In_2321);
nand U2899 (N_2899,In_1153,In_439);
and U2900 (N_2900,In_359,In_2509);
or U2901 (N_2901,In_2030,In_1038);
or U2902 (N_2902,In_1075,In_905);
nand U2903 (N_2903,In_437,In_2439);
nor U2904 (N_2904,In_261,In_355);
xnor U2905 (N_2905,In_1028,In_1267);
or U2906 (N_2906,In_261,In_2632);
or U2907 (N_2907,In_2228,In_1687);
and U2908 (N_2908,In_421,In_2068);
nor U2909 (N_2909,In_1607,In_444);
nand U2910 (N_2910,In_2206,In_2629);
nand U2911 (N_2911,In_250,In_2354);
or U2912 (N_2912,In_401,In_2844);
and U2913 (N_2913,In_681,In_1580);
nand U2914 (N_2914,In_2513,In_112);
nor U2915 (N_2915,In_2746,In_2883);
or U2916 (N_2916,In_533,In_900);
nand U2917 (N_2917,In_2705,In_1231);
or U2918 (N_2918,In_1816,In_2915);
nand U2919 (N_2919,In_1976,In_315);
and U2920 (N_2920,In_1006,In_121);
nand U2921 (N_2921,In_737,In_2521);
nand U2922 (N_2922,In_2946,In_1677);
and U2923 (N_2923,In_618,In_2785);
or U2924 (N_2924,In_65,In_950);
nand U2925 (N_2925,In_2028,In_963);
and U2926 (N_2926,In_2286,In_1163);
nor U2927 (N_2927,In_197,In_2131);
nand U2928 (N_2928,In_1038,In_946);
nor U2929 (N_2929,In_1337,In_20);
nand U2930 (N_2930,In_2551,In_853);
or U2931 (N_2931,In_1975,In_2694);
and U2932 (N_2932,In_876,In_624);
nand U2933 (N_2933,In_724,In_1416);
or U2934 (N_2934,In_2458,In_837);
or U2935 (N_2935,In_437,In_2194);
or U2936 (N_2936,In_1805,In_128);
nor U2937 (N_2937,In_1773,In_777);
nand U2938 (N_2938,In_1868,In_1470);
and U2939 (N_2939,In_2167,In_676);
nand U2940 (N_2940,In_1149,In_1027);
or U2941 (N_2941,In_1232,In_845);
xor U2942 (N_2942,In_1212,In_124);
nor U2943 (N_2943,In_2108,In_1770);
nor U2944 (N_2944,In_925,In_2776);
or U2945 (N_2945,In_617,In_468);
nand U2946 (N_2946,In_1976,In_1401);
and U2947 (N_2947,In_2429,In_2801);
or U2948 (N_2948,In_2867,In_2776);
or U2949 (N_2949,In_993,In_2987);
or U2950 (N_2950,In_136,In_1559);
or U2951 (N_2951,In_2384,In_1008);
nand U2952 (N_2952,In_1248,In_2822);
nor U2953 (N_2953,In_596,In_1804);
nand U2954 (N_2954,In_2658,In_1571);
nand U2955 (N_2955,In_1514,In_205);
xor U2956 (N_2956,In_1274,In_1552);
nor U2957 (N_2957,In_160,In_2151);
or U2958 (N_2958,In_2753,In_750);
nand U2959 (N_2959,In_538,In_2692);
nor U2960 (N_2960,In_2316,In_2811);
nor U2961 (N_2961,In_623,In_751);
xnor U2962 (N_2962,In_2376,In_247);
nand U2963 (N_2963,In_2238,In_2249);
or U2964 (N_2964,In_2158,In_2847);
nand U2965 (N_2965,In_427,In_69);
nand U2966 (N_2966,In_1002,In_2833);
or U2967 (N_2967,In_2855,In_1415);
nor U2968 (N_2968,In_989,In_2662);
or U2969 (N_2969,In_1261,In_808);
nor U2970 (N_2970,In_601,In_43);
nor U2971 (N_2971,In_8,In_206);
and U2972 (N_2972,In_2776,In_777);
or U2973 (N_2973,In_1542,In_1838);
and U2974 (N_2974,In_1454,In_1075);
nand U2975 (N_2975,In_2641,In_2451);
nor U2976 (N_2976,In_2323,In_1072);
xnor U2977 (N_2977,In_1398,In_1840);
nor U2978 (N_2978,In_1143,In_2326);
and U2979 (N_2979,In_1973,In_888);
nor U2980 (N_2980,In_896,In_2341);
nand U2981 (N_2981,In_1389,In_2892);
nand U2982 (N_2982,In_685,In_2104);
nor U2983 (N_2983,In_832,In_585);
nand U2984 (N_2984,In_1971,In_774);
or U2985 (N_2985,In_2671,In_2369);
nor U2986 (N_2986,In_1223,In_1892);
nand U2987 (N_2987,In_1677,In_86);
and U2988 (N_2988,In_1715,In_63);
nor U2989 (N_2989,In_1183,In_2478);
or U2990 (N_2990,In_2120,In_2449);
nor U2991 (N_2991,In_2146,In_1280);
nand U2992 (N_2992,In_1787,In_796);
or U2993 (N_2993,In_2629,In_2753);
nand U2994 (N_2994,In_2396,In_1094);
and U2995 (N_2995,In_1780,In_797);
nor U2996 (N_2996,In_2417,In_1199);
nor U2997 (N_2997,In_592,In_2240);
xnor U2998 (N_2998,In_2342,In_2251);
and U2999 (N_2999,In_1753,In_1095);
or U3000 (N_3000,In_2984,In_1998);
nor U3001 (N_3001,In_2076,In_31);
nor U3002 (N_3002,In_419,In_901);
nand U3003 (N_3003,In_2255,In_2086);
nand U3004 (N_3004,In_2977,In_1534);
or U3005 (N_3005,In_1349,In_759);
and U3006 (N_3006,In_115,In_2119);
xor U3007 (N_3007,In_1313,In_666);
or U3008 (N_3008,In_523,In_2909);
and U3009 (N_3009,In_936,In_1701);
or U3010 (N_3010,In_2572,In_2365);
nor U3011 (N_3011,In_590,In_768);
xnor U3012 (N_3012,In_555,In_1314);
and U3013 (N_3013,In_670,In_2334);
nor U3014 (N_3014,In_1645,In_1128);
or U3015 (N_3015,In_1795,In_2864);
nand U3016 (N_3016,In_769,In_1998);
or U3017 (N_3017,In_2970,In_2414);
or U3018 (N_3018,In_1724,In_2105);
nor U3019 (N_3019,In_2167,In_1483);
or U3020 (N_3020,In_718,In_1880);
nand U3021 (N_3021,In_2468,In_1639);
nand U3022 (N_3022,In_910,In_1864);
nor U3023 (N_3023,In_2587,In_962);
and U3024 (N_3024,In_621,In_2227);
nor U3025 (N_3025,In_1136,In_2493);
nor U3026 (N_3026,In_320,In_1599);
nor U3027 (N_3027,In_2648,In_879);
or U3028 (N_3028,In_49,In_2540);
xor U3029 (N_3029,In_1101,In_544);
xnor U3030 (N_3030,In_2083,In_867);
nand U3031 (N_3031,In_2303,In_859);
nor U3032 (N_3032,In_1717,In_2480);
nand U3033 (N_3033,In_2826,In_2973);
or U3034 (N_3034,In_2436,In_1761);
or U3035 (N_3035,In_1006,In_1906);
and U3036 (N_3036,In_2963,In_2262);
and U3037 (N_3037,In_2000,In_25);
nor U3038 (N_3038,In_1325,In_2094);
nor U3039 (N_3039,In_1726,In_1099);
or U3040 (N_3040,In_1997,In_9);
or U3041 (N_3041,In_1206,In_1236);
nor U3042 (N_3042,In_1178,In_1439);
nor U3043 (N_3043,In_804,In_2703);
xnor U3044 (N_3044,In_859,In_2414);
nand U3045 (N_3045,In_2814,In_1963);
or U3046 (N_3046,In_428,In_627);
nor U3047 (N_3047,In_2722,In_119);
or U3048 (N_3048,In_1785,In_53);
nor U3049 (N_3049,In_1257,In_2974);
nor U3050 (N_3050,In_1129,In_2447);
or U3051 (N_3051,In_118,In_2500);
and U3052 (N_3052,In_970,In_1262);
nand U3053 (N_3053,In_2037,In_2619);
nor U3054 (N_3054,In_1821,In_2252);
xnor U3055 (N_3055,In_2578,In_1132);
and U3056 (N_3056,In_962,In_273);
xor U3057 (N_3057,In_430,In_2656);
or U3058 (N_3058,In_1722,In_2794);
or U3059 (N_3059,In_2229,In_1353);
xor U3060 (N_3060,In_1533,In_2914);
nand U3061 (N_3061,In_1766,In_597);
and U3062 (N_3062,In_2129,In_960);
or U3063 (N_3063,In_2681,In_30);
nand U3064 (N_3064,In_1478,In_1488);
or U3065 (N_3065,In_1563,In_272);
nand U3066 (N_3066,In_2472,In_2497);
or U3067 (N_3067,In_96,In_2820);
xor U3068 (N_3068,In_1525,In_2758);
and U3069 (N_3069,In_334,In_2859);
and U3070 (N_3070,In_2854,In_844);
or U3071 (N_3071,In_2339,In_1725);
nor U3072 (N_3072,In_2729,In_2283);
nand U3073 (N_3073,In_2126,In_1576);
nand U3074 (N_3074,In_1655,In_2085);
nand U3075 (N_3075,In_1366,In_1264);
or U3076 (N_3076,In_1035,In_991);
or U3077 (N_3077,In_1385,In_1064);
nand U3078 (N_3078,In_454,In_1212);
and U3079 (N_3079,In_75,In_2789);
and U3080 (N_3080,In_0,In_945);
nor U3081 (N_3081,In_585,In_1130);
nand U3082 (N_3082,In_2132,In_2007);
nand U3083 (N_3083,In_1346,In_1413);
or U3084 (N_3084,In_2025,In_2313);
nor U3085 (N_3085,In_2884,In_2821);
and U3086 (N_3086,In_2072,In_256);
nor U3087 (N_3087,In_1060,In_1787);
nor U3088 (N_3088,In_730,In_2073);
and U3089 (N_3089,In_2378,In_2256);
and U3090 (N_3090,In_644,In_2076);
and U3091 (N_3091,In_1481,In_2052);
nor U3092 (N_3092,In_2356,In_1378);
and U3093 (N_3093,In_579,In_2320);
or U3094 (N_3094,In_199,In_558);
and U3095 (N_3095,In_506,In_103);
nand U3096 (N_3096,In_46,In_933);
or U3097 (N_3097,In_8,In_480);
nand U3098 (N_3098,In_976,In_520);
and U3099 (N_3099,In_792,In_2323);
or U3100 (N_3100,In_2684,In_126);
and U3101 (N_3101,In_2466,In_1373);
or U3102 (N_3102,In_2145,In_1678);
nor U3103 (N_3103,In_2542,In_833);
nand U3104 (N_3104,In_234,In_712);
nand U3105 (N_3105,In_2711,In_964);
or U3106 (N_3106,In_255,In_2882);
xnor U3107 (N_3107,In_2699,In_2687);
xnor U3108 (N_3108,In_1634,In_1364);
nor U3109 (N_3109,In_474,In_2927);
nor U3110 (N_3110,In_508,In_1347);
or U3111 (N_3111,In_954,In_2914);
nor U3112 (N_3112,In_2054,In_2636);
and U3113 (N_3113,In_1892,In_249);
or U3114 (N_3114,In_2412,In_1562);
or U3115 (N_3115,In_284,In_2322);
and U3116 (N_3116,In_847,In_1854);
nand U3117 (N_3117,In_173,In_2584);
and U3118 (N_3118,In_1570,In_1532);
nor U3119 (N_3119,In_1791,In_476);
or U3120 (N_3120,In_1889,In_2045);
nor U3121 (N_3121,In_1979,In_1708);
or U3122 (N_3122,In_1745,In_1024);
nand U3123 (N_3123,In_1845,In_2171);
or U3124 (N_3124,In_1745,In_2036);
nor U3125 (N_3125,In_1938,In_2726);
and U3126 (N_3126,In_1095,In_788);
xor U3127 (N_3127,In_721,In_1407);
and U3128 (N_3128,In_344,In_411);
xor U3129 (N_3129,In_2959,In_1258);
and U3130 (N_3130,In_11,In_1030);
and U3131 (N_3131,In_444,In_1237);
and U3132 (N_3132,In_2220,In_555);
and U3133 (N_3133,In_168,In_2451);
and U3134 (N_3134,In_21,In_103);
or U3135 (N_3135,In_599,In_30);
nor U3136 (N_3136,In_2685,In_2128);
nand U3137 (N_3137,In_1550,In_2645);
xnor U3138 (N_3138,In_114,In_2443);
and U3139 (N_3139,In_842,In_548);
or U3140 (N_3140,In_1116,In_509);
or U3141 (N_3141,In_1702,In_2032);
nor U3142 (N_3142,In_855,In_143);
and U3143 (N_3143,In_821,In_1941);
or U3144 (N_3144,In_442,In_209);
nand U3145 (N_3145,In_1194,In_2465);
and U3146 (N_3146,In_939,In_2273);
and U3147 (N_3147,In_2060,In_415);
nand U3148 (N_3148,In_1789,In_1638);
and U3149 (N_3149,In_693,In_1693);
and U3150 (N_3150,In_2080,In_1960);
nand U3151 (N_3151,In_31,In_229);
nor U3152 (N_3152,In_530,In_1271);
xnor U3153 (N_3153,In_1987,In_1421);
nor U3154 (N_3154,In_356,In_600);
xnor U3155 (N_3155,In_44,In_10);
nor U3156 (N_3156,In_1398,In_779);
nor U3157 (N_3157,In_1982,In_2352);
and U3158 (N_3158,In_961,In_2611);
nand U3159 (N_3159,In_2046,In_2334);
or U3160 (N_3160,In_1829,In_1800);
xnor U3161 (N_3161,In_1124,In_2719);
and U3162 (N_3162,In_2374,In_1988);
or U3163 (N_3163,In_954,In_842);
nor U3164 (N_3164,In_1386,In_1931);
xor U3165 (N_3165,In_2551,In_843);
or U3166 (N_3166,In_1300,In_1200);
nor U3167 (N_3167,In_1793,In_118);
or U3168 (N_3168,In_2875,In_1135);
nor U3169 (N_3169,In_2075,In_1540);
or U3170 (N_3170,In_237,In_2461);
nor U3171 (N_3171,In_1067,In_1773);
xnor U3172 (N_3172,In_1436,In_184);
nor U3173 (N_3173,In_564,In_1235);
nand U3174 (N_3174,In_2622,In_1375);
nand U3175 (N_3175,In_2206,In_25);
and U3176 (N_3176,In_1050,In_1867);
and U3177 (N_3177,In_2628,In_2737);
nor U3178 (N_3178,In_2052,In_819);
or U3179 (N_3179,In_2061,In_923);
or U3180 (N_3180,In_611,In_2428);
nand U3181 (N_3181,In_2457,In_2318);
nand U3182 (N_3182,In_2672,In_152);
or U3183 (N_3183,In_404,In_2079);
or U3184 (N_3184,In_1183,In_587);
or U3185 (N_3185,In_1317,In_1298);
nor U3186 (N_3186,In_2797,In_2085);
and U3187 (N_3187,In_1232,In_2306);
or U3188 (N_3188,In_1816,In_2220);
nand U3189 (N_3189,In_2586,In_2489);
or U3190 (N_3190,In_550,In_315);
nor U3191 (N_3191,In_1345,In_447);
xor U3192 (N_3192,In_391,In_1272);
or U3193 (N_3193,In_2160,In_892);
xnor U3194 (N_3194,In_203,In_1209);
nor U3195 (N_3195,In_2838,In_262);
and U3196 (N_3196,In_707,In_1657);
nand U3197 (N_3197,In_872,In_332);
or U3198 (N_3198,In_1387,In_2127);
nor U3199 (N_3199,In_2755,In_1906);
and U3200 (N_3200,In_208,In_1442);
or U3201 (N_3201,In_892,In_583);
and U3202 (N_3202,In_2102,In_2796);
xor U3203 (N_3203,In_1686,In_477);
nand U3204 (N_3204,In_2336,In_1842);
xor U3205 (N_3205,In_2579,In_1164);
nor U3206 (N_3206,In_2808,In_433);
or U3207 (N_3207,In_854,In_1021);
nor U3208 (N_3208,In_2271,In_2419);
nor U3209 (N_3209,In_352,In_2752);
and U3210 (N_3210,In_2165,In_553);
or U3211 (N_3211,In_431,In_1094);
nand U3212 (N_3212,In_617,In_2645);
nor U3213 (N_3213,In_1250,In_375);
nor U3214 (N_3214,In_235,In_1939);
xnor U3215 (N_3215,In_769,In_2164);
nand U3216 (N_3216,In_76,In_2456);
nand U3217 (N_3217,In_1430,In_1066);
xnor U3218 (N_3218,In_1532,In_450);
nand U3219 (N_3219,In_906,In_1220);
nand U3220 (N_3220,In_1675,In_396);
or U3221 (N_3221,In_150,In_2111);
nor U3222 (N_3222,In_1713,In_1697);
and U3223 (N_3223,In_2113,In_41);
nand U3224 (N_3224,In_1991,In_56);
and U3225 (N_3225,In_748,In_712);
or U3226 (N_3226,In_1100,In_1635);
xnor U3227 (N_3227,In_2564,In_775);
or U3228 (N_3228,In_2498,In_417);
nor U3229 (N_3229,In_596,In_394);
and U3230 (N_3230,In_992,In_1267);
or U3231 (N_3231,In_254,In_422);
xor U3232 (N_3232,In_2109,In_2316);
and U3233 (N_3233,In_2684,In_2831);
nand U3234 (N_3234,In_2360,In_1210);
nand U3235 (N_3235,In_461,In_336);
nor U3236 (N_3236,In_2277,In_2712);
nor U3237 (N_3237,In_2737,In_2799);
or U3238 (N_3238,In_1622,In_566);
nor U3239 (N_3239,In_2105,In_428);
or U3240 (N_3240,In_2883,In_611);
or U3241 (N_3241,In_341,In_2771);
nand U3242 (N_3242,In_2584,In_1476);
nand U3243 (N_3243,In_508,In_958);
and U3244 (N_3244,In_1176,In_1051);
nand U3245 (N_3245,In_2497,In_2309);
and U3246 (N_3246,In_1138,In_635);
xor U3247 (N_3247,In_1966,In_690);
and U3248 (N_3248,In_72,In_1973);
or U3249 (N_3249,In_2906,In_862);
nand U3250 (N_3250,In_2514,In_2094);
xor U3251 (N_3251,In_2012,In_2089);
xor U3252 (N_3252,In_224,In_592);
nand U3253 (N_3253,In_2693,In_199);
xnor U3254 (N_3254,In_2523,In_1003);
xor U3255 (N_3255,In_2788,In_1389);
and U3256 (N_3256,In_902,In_2670);
or U3257 (N_3257,In_18,In_2871);
and U3258 (N_3258,In_2303,In_1148);
or U3259 (N_3259,In_911,In_198);
nand U3260 (N_3260,In_2476,In_1981);
nand U3261 (N_3261,In_2938,In_2422);
xor U3262 (N_3262,In_1977,In_2208);
xor U3263 (N_3263,In_1436,In_1366);
nor U3264 (N_3264,In_1245,In_1498);
nor U3265 (N_3265,In_382,In_1936);
and U3266 (N_3266,In_1934,In_1408);
and U3267 (N_3267,In_168,In_810);
nor U3268 (N_3268,In_453,In_358);
nand U3269 (N_3269,In_743,In_455);
nand U3270 (N_3270,In_1542,In_1697);
nor U3271 (N_3271,In_2060,In_2096);
and U3272 (N_3272,In_218,In_2102);
nor U3273 (N_3273,In_1786,In_1412);
and U3274 (N_3274,In_1180,In_1690);
or U3275 (N_3275,In_1679,In_536);
nor U3276 (N_3276,In_971,In_1828);
and U3277 (N_3277,In_2452,In_2850);
nor U3278 (N_3278,In_1862,In_1985);
and U3279 (N_3279,In_683,In_1689);
nand U3280 (N_3280,In_544,In_1883);
nor U3281 (N_3281,In_1011,In_123);
nor U3282 (N_3282,In_2149,In_1528);
nor U3283 (N_3283,In_1257,In_2039);
and U3284 (N_3284,In_1753,In_164);
nand U3285 (N_3285,In_1446,In_1889);
xor U3286 (N_3286,In_867,In_478);
or U3287 (N_3287,In_436,In_1778);
xor U3288 (N_3288,In_1987,In_1288);
nand U3289 (N_3289,In_2750,In_714);
xnor U3290 (N_3290,In_2901,In_2672);
and U3291 (N_3291,In_1499,In_1415);
nor U3292 (N_3292,In_2901,In_1251);
and U3293 (N_3293,In_615,In_1254);
nand U3294 (N_3294,In_1471,In_1565);
xor U3295 (N_3295,In_1979,In_2496);
nor U3296 (N_3296,In_2699,In_338);
nand U3297 (N_3297,In_1478,In_2533);
nand U3298 (N_3298,In_654,In_2815);
or U3299 (N_3299,In_1201,In_2844);
xor U3300 (N_3300,In_1078,In_2450);
nand U3301 (N_3301,In_1968,In_1186);
or U3302 (N_3302,In_2887,In_859);
and U3303 (N_3303,In_2863,In_83);
nand U3304 (N_3304,In_1980,In_1728);
and U3305 (N_3305,In_2919,In_725);
and U3306 (N_3306,In_2736,In_324);
nand U3307 (N_3307,In_62,In_2947);
xnor U3308 (N_3308,In_291,In_2157);
xnor U3309 (N_3309,In_2309,In_1523);
and U3310 (N_3310,In_1336,In_2660);
and U3311 (N_3311,In_1953,In_1394);
nor U3312 (N_3312,In_1087,In_1813);
and U3313 (N_3313,In_1607,In_1785);
nor U3314 (N_3314,In_1035,In_199);
xor U3315 (N_3315,In_37,In_552);
or U3316 (N_3316,In_1824,In_371);
xor U3317 (N_3317,In_1560,In_1276);
nor U3318 (N_3318,In_1224,In_2826);
nor U3319 (N_3319,In_2617,In_676);
nor U3320 (N_3320,In_1707,In_629);
and U3321 (N_3321,In_2046,In_1769);
xnor U3322 (N_3322,In_2385,In_361);
nor U3323 (N_3323,In_871,In_1044);
nor U3324 (N_3324,In_555,In_2215);
nand U3325 (N_3325,In_601,In_616);
and U3326 (N_3326,In_1102,In_1183);
xor U3327 (N_3327,In_277,In_2107);
or U3328 (N_3328,In_2201,In_1012);
and U3329 (N_3329,In_747,In_742);
nor U3330 (N_3330,In_1404,In_1145);
nor U3331 (N_3331,In_1868,In_2590);
or U3332 (N_3332,In_2317,In_1048);
and U3333 (N_3333,In_1853,In_1137);
and U3334 (N_3334,In_2301,In_2586);
xor U3335 (N_3335,In_715,In_1463);
or U3336 (N_3336,In_1131,In_2402);
nand U3337 (N_3337,In_2533,In_607);
nand U3338 (N_3338,In_1232,In_769);
or U3339 (N_3339,In_2912,In_221);
or U3340 (N_3340,In_504,In_2188);
nor U3341 (N_3341,In_531,In_419);
nand U3342 (N_3342,In_1844,In_1341);
nor U3343 (N_3343,In_779,In_2319);
xor U3344 (N_3344,In_207,In_963);
or U3345 (N_3345,In_1199,In_973);
or U3346 (N_3346,In_1418,In_2164);
xnor U3347 (N_3347,In_1721,In_836);
or U3348 (N_3348,In_572,In_2470);
and U3349 (N_3349,In_1172,In_1288);
nand U3350 (N_3350,In_2795,In_44);
and U3351 (N_3351,In_1677,In_62);
nand U3352 (N_3352,In_2056,In_1720);
or U3353 (N_3353,In_2311,In_283);
nor U3354 (N_3354,In_2503,In_989);
and U3355 (N_3355,In_1652,In_2592);
nor U3356 (N_3356,In_283,In_665);
or U3357 (N_3357,In_140,In_2206);
xnor U3358 (N_3358,In_703,In_2185);
and U3359 (N_3359,In_2582,In_299);
and U3360 (N_3360,In_2643,In_2331);
and U3361 (N_3361,In_2419,In_575);
nand U3362 (N_3362,In_1586,In_771);
or U3363 (N_3363,In_2278,In_2249);
xnor U3364 (N_3364,In_1915,In_2011);
or U3365 (N_3365,In_187,In_1446);
or U3366 (N_3366,In_2575,In_1679);
nand U3367 (N_3367,In_2534,In_2599);
or U3368 (N_3368,In_213,In_2203);
nor U3369 (N_3369,In_2234,In_2757);
or U3370 (N_3370,In_1112,In_514);
or U3371 (N_3371,In_257,In_2823);
nor U3372 (N_3372,In_2962,In_1704);
or U3373 (N_3373,In_1448,In_2293);
nand U3374 (N_3374,In_1688,In_1276);
nor U3375 (N_3375,In_222,In_599);
xnor U3376 (N_3376,In_894,In_1371);
and U3377 (N_3377,In_2929,In_1646);
or U3378 (N_3378,In_741,In_2486);
nand U3379 (N_3379,In_620,In_139);
and U3380 (N_3380,In_1213,In_123);
or U3381 (N_3381,In_169,In_761);
nor U3382 (N_3382,In_2161,In_1288);
or U3383 (N_3383,In_1912,In_2491);
and U3384 (N_3384,In_2350,In_1196);
and U3385 (N_3385,In_1565,In_1247);
nand U3386 (N_3386,In_1481,In_1838);
or U3387 (N_3387,In_692,In_489);
and U3388 (N_3388,In_1774,In_2256);
nor U3389 (N_3389,In_1429,In_720);
nor U3390 (N_3390,In_374,In_2827);
and U3391 (N_3391,In_1069,In_1669);
xor U3392 (N_3392,In_585,In_1129);
or U3393 (N_3393,In_2853,In_1877);
and U3394 (N_3394,In_2827,In_513);
or U3395 (N_3395,In_1921,In_1896);
and U3396 (N_3396,In_1926,In_746);
or U3397 (N_3397,In_1422,In_1040);
nor U3398 (N_3398,In_22,In_1894);
and U3399 (N_3399,In_347,In_368);
xor U3400 (N_3400,In_1858,In_2793);
and U3401 (N_3401,In_2679,In_2754);
and U3402 (N_3402,In_430,In_1392);
xor U3403 (N_3403,In_1255,In_946);
nor U3404 (N_3404,In_2302,In_2885);
or U3405 (N_3405,In_2653,In_2408);
nor U3406 (N_3406,In_2533,In_1496);
and U3407 (N_3407,In_1571,In_2310);
nand U3408 (N_3408,In_2853,In_1591);
nor U3409 (N_3409,In_1261,In_74);
or U3410 (N_3410,In_2169,In_2007);
or U3411 (N_3411,In_1949,In_1928);
xnor U3412 (N_3412,In_855,In_691);
nand U3413 (N_3413,In_1836,In_1453);
or U3414 (N_3414,In_507,In_2060);
or U3415 (N_3415,In_2570,In_1646);
or U3416 (N_3416,In_2550,In_195);
xnor U3417 (N_3417,In_1336,In_972);
xor U3418 (N_3418,In_145,In_2675);
xnor U3419 (N_3419,In_1656,In_1489);
xor U3420 (N_3420,In_2007,In_1708);
and U3421 (N_3421,In_115,In_920);
or U3422 (N_3422,In_2505,In_2401);
nand U3423 (N_3423,In_1311,In_1174);
nand U3424 (N_3424,In_1793,In_777);
or U3425 (N_3425,In_2060,In_1851);
or U3426 (N_3426,In_2699,In_2208);
and U3427 (N_3427,In_945,In_2206);
nand U3428 (N_3428,In_48,In_807);
or U3429 (N_3429,In_1050,In_256);
or U3430 (N_3430,In_1131,In_2207);
or U3431 (N_3431,In_801,In_37);
or U3432 (N_3432,In_685,In_1118);
and U3433 (N_3433,In_20,In_392);
nor U3434 (N_3434,In_2682,In_1415);
and U3435 (N_3435,In_832,In_484);
or U3436 (N_3436,In_573,In_29);
nand U3437 (N_3437,In_2373,In_2973);
xor U3438 (N_3438,In_460,In_2118);
or U3439 (N_3439,In_1198,In_1579);
or U3440 (N_3440,In_2024,In_1454);
nor U3441 (N_3441,In_1411,In_2513);
nor U3442 (N_3442,In_883,In_281);
nor U3443 (N_3443,In_2389,In_1782);
and U3444 (N_3444,In_2302,In_1642);
and U3445 (N_3445,In_1266,In_1652);
nand U3446 (N_3446,In_2054,In_483);
nor U3447 (N_3447,In_2567,In_1424);
or U3448 (N_3448,In_2633,In_1040);
nand U3449 (N_3449,In_1457,In_2762);
and U3450 (N_3450,In_2026,In_990);
or U3451 (N_3451,In_2446,In_2470);
and U3452 (N_3452,In_992,In_1872);
nor U3453 (N_3453,In_1820,In_2254);
nand U3454 (N_3454,In_2532,In_1505);
or U3455 (N_3455,In_53,In_1745);
nand U3456 (N_3456,In_88,In_1588);
or U3457 (N_3457,In_2741,In_2703);
xnor U3458 (N_3458,In_2,In_1824);
and U3459 (N_3459,In_2383,In_2657);
and U3460 (N_3460,In_1582,In_1936);
and U3461 (N_3461,In_1159,In_2562);
nor U3462 (N_3462,In_435,In_324);
nor U3463 (N_3463,In_400,In_742);
and U3464 (N_3464,In_718,In_1204);
nand U3465 (N_3465,In_2083,In_2728);
nor U3466 (N_3466,In_1153,In_2399);
nand U3467 (N_3467,In_2403,In_2937);
nand U3468 (N_3468,In_2335,In_1273);
nand U3469 (N_3469,In_2448,In_519);
xor U3470 (N_3470,In_2922,In_969);
nand U3471 (N_3471,In_1079,In_2050);
nand U3472 (N_3472,In_22,In_1248);
nand U3473 (N_3473,In_2875,In_475);
nand U3474 (N_3474,In_190,In_2053);
xor U3475 (N_3475,In_2813,In_677);
and U3476 (N_3476,In_1990,In_574);
nand U3477 (N_3477,In_691,In_1072);
or U3478 (N_3478,In_2343,In_2524);
or U3479 (N_3479,In_1870,In_1783);
nor U3480 (N_3480,In_1477,In_197);
and U3481 (N_3481,In_1864,In_2213);
or U3482 (N_3482,In_1776,In_99);
nor U3483 (N_3483,In_2781,In_2846);
and U3484 (N_3484,In_1366,In_1567);
nand U3485 (N_3485,In_1635,In_241);
nor U3486 (N_3486,In_1959,In_432);
nand U3487 (N_3487,In_72,In_1176);
and U3488 (N_3488,In_2008,In_2807);
and U3489 (N_3489,In_2410,In_813);
and U3490 (N_3490,In_2161,In_1104);
or U3491 (N_3491,In_333,In_2428);
nand U3492 (N_3492,In_7,In_409);
nand U3493 (N_3493,In_1081,In_919);
nand U3494 (N_3494,In_1071,In_83);
xnor U3495 (N_3495,In_587,In_180);
nand U3496 (N_3496,In_1021,In_357);
xnor U3497 (N_3497,In_721,In_1886);
nand U3498 (N_3498,In_1907,In_2997);
or U3499 (N_3499,In_282,In_2092);
and U3500 (N_3500,In_1615,In_2219);
and U3501 (N_3501,In_626,In_1963);
nand U3502 (N_3502,In_1442,In_814);
and U3503 (N_3503,In_2481,In_297);
or U3504 (N_3504,In_1698,In_1590);
nor U3505 (N_3505,In_566,In_2448);
nand U3506 (N_3506,In_2064,In_658);
and U3507 (N_3507,In_704,In_1498);
nor U3508 (N_3508,In_2566,In_387);
nand U3509 (N_3509,In_1631,In_2888);
nor U3510 (N_3510,In_870,In_2171);
nand U3511 (N_3511,In_600,In_2262);
nor U3512 (N_3512,In_2236,In_559);
nor U3513 (N_3513,In_2200,In_1567);
and U3514 (N_3514,In_1669,In_787);
or U3515 (N_3515,In_2264,In_1682);
and U3516 (N_3516,In_2434,In_356);
nor U3517 (N_3517,In_2635,In_1003);
or U3518 (N_3518,In_2878,In_866);
xnor U3519 (N_3519,In_1568,In_1457);
or U3520 (N_3520,In_2220,In_1982);
or U3521 (N_3521,In_1148,In_1564);
nand U3522 (N_3522,In_2394,In_376);
or U3523 (N_3523,In_1072,In_1326);
nor U3524 (N_3524,In_278,In_1763);
nor U3525 (N_3525,In_2802,In_460);
or U3526 (N_3526,In_280,In_2141);
and U3527 (N_3527,In_2442,In_1700);
nor U3528 (N_3528,In_1684,In_2252);
and U3529 (N_3529,In_121,In_2874);
nand U3530 (N_3530,In_2824,In_1446);
xor U3531 (N_3531,In_108,In_1040);
or U3532 (N_3532,In_2095,In_1457);
nand U3533 (N_3533,In_393,In_2282);
nand U3534 (N_3534,In_2150,In_2100);
nand U3535 (N_3535,In_978,In_1018);
xor U3536 (N_3536,In_43,In_422);
and U3537 (N_3537,In_494,In_687);
nand U3538 (N_3538,In_213,In_328);
and U3539 (N_3539,In_777,In_139);
xnor U3540 (N_3540,In_363,In_894);
xnor U3541 (N_3541,In_1107,In_2223);
xnor U3542 (N_3542,In_1695,In_510);
or U3543 (N_3543,In_226,In_573);
nor U3544 (N_3544,In_1829,In_1620);
and U3545 (N_3545,In_2703,In_2309);
nor U3546 (N_3546,In_2944,In_2778);
and U3547 (N_3547,In_1595,In_958);
or U3548 (N_3548,In_351,In_2445);
or U3549 (N_3549,In_2706,In_325);
nand U3550 (N_3550,In_729,In_446);
or U3551 (N_3551,In_1929,In_974);
and U3552 (N_3552,In_1508,In_1348);
xnor U3553 (N_3553,In_152,In_646);
nor U3554 (N_3554,In_1826,In_2890);
nand U3555 (N_3555,In_1258,In_2266);
nand U3556 (N_3556,In_2252,In_533);
xnor U3557 (N_3557,In_2319,In_602);
nand U3558 (N_3558,In_171,In_498);
and U3559 (N_3559,In_2941,In_490);
or U3560 (N_3560,In_690,In_2712);
and U3561 (N_3561,In_249,In_2897);
and U3562 (N_3562,In_2125,In_796);
and U3563 (N_3563,In_2231,In_573);
nand U3564 (N_3564,In_907,In_2059);
nand U3565 (N_3565,In_1170,In_2201);
nand U3566 (N_3566,In_234,In_438);
and U3567 (N_3567,In_2733,In_537);
or U3568 (N_3568,In_425,In_1110);
nor U3569 (N_3569,In_2398,In_1108);
nand U3570 (N_3570,In_2473,In_2775);
and U3571 (N_3571,In_2603,In_2289);
and U3572 (N_3572,In_1605,In_227);
nor U3573 (N_3573,In_1028,In_1050);
and U3574 (N_3574,In_2742,In_875);
nor U3575 (N_3575,In_376,In_122);
nand U3576 (N_3576,In_2528,In_470);
and U3577 (N_3577,In_1909,In_2861);
or U3578 (N_3578,In_1434,In_973);
and U3579 (N_3579,In_2383,In_267);
or U3580 (N_3580,In_2612,In_1684);
or U3581 (N_3581,In_2979,In_2670);
and U3582 (N_3582,In_2206,In_1942);
and U3583 (N_3583,In_12,In_2275);
nor U3584 (N_3584,In_946,In_1357);
xor U3585 (N_3585,In_1034,In_374);
xor U3586 (N_3586,In_1005,In_2384);
or U3587 (N_3587,In_2950,In_893);
xor U3588 (N_3588,In_1403,In_1979);
and U3589 (N_3589,In_708,In_915);
nor U3590 (N_3590,In_1001,In_2907);
nor U3591 (N_3591,In_1252,In_1531);
and U3592 (N_3592,In_2270,In_2747);
or U3593 (N_3593,In_1414,In_472);
or U3594 (N_3594,In_811,In_119);
nand U3595 (N_3595,In_2714,In_2866);
nor U3596 (N_3596,In_1876,In_536);
nor U3597 (N_3597,In_1081,In_953);
nor U3598 (N_3598,In_1366,In_1429);
or U3599 (N_3599,In_204,In_982);
xor U3600 (N_3600,In_250,In_2741);
nor U3601 (N_3601,In_1623,In_1361);
nor U3602 (N_3602,In_1727,In_323);
nand U3603 (N_3603,In_2180,In_2469);
nand U3604 (N_3604,In_1371,In_1201);
or U3605 (N_3605,In_2805,In_626);
nand U3606 (N_3606,In_566,In_628);
or U3607 (N_3607,In_2192,In_2800);
or U3608 (N_3608,In_1277,In_1886);
or U3609 (N_3609,In_1847,In_1639);
or U3610 (N_3610,In_1043,In_239);
or U3611 (N_3611,In_1585,In_1710);
nand U3612 (N_3612,In_1575,In_1075);
nand U3613 (N_3613,In_1995,In_665);
nand U3614 (N_3614,In_2090,In_1617);
nor U3615 (N_3615,In_897,In_667);
nand U3616 (N_3616,In_17,In_779);
nand U3617 (N_3617,In_1841,In_913);
or U3618 (N_3618,In_700,In_2964);
nor U3619 (N_3619,In_1173,In_1025);
or U3620 (N_3620,In_1552,In_1221);
and U3621 (N_3621,In_1507,In_1592);
or U3622 (N_3622,In_2390,In_1309);
nand U3623 (N_3623,In_2022,In_2795);
or U3624 (N_3624,In_1696,In_1158);
nand U3625 (N_3625,In_2288,In_2933);
and U3626 (N_3626,In_675,In_2733);
nor U3627 (N_3627,In_2227,In_629);
and U3628 (N_3628,In_70,In_2621);
nand U3629 (N_3629,In_2139,In_2595);
or U3630 (N_3630,In_1569,In_1007);
or U3631 (N_3631,In_2949,In_1240);
nor U3632 (N_3632,In_2249,In_2189);
or U3633 (N_3633,In_900,In_2381);
nand U3634 (N_3634,In_1708,In_1166);
nand U3635 (N_3635,In_320,In_1917);
nand U3636 (N_3636,In_2578,In_1532);
xor U3637 (N_3637,In_670,In_775);
nor U3638 (N_3638,In_2132,In_52);
or U3639 (N_3639,In_1184,In_996);
nand U3640 (N_3640,In_2729,In_2964);
or U3641 (N_3641,In_2448,In_1240);
nor U3642 (N_3642,In_17,In_831);
and U3643 (N_3643,In_1051,In_441);
and U3644 (N_3644,In_1697,In_1770);
nor U3645 (N_3645,In_2698,In_293);
nand U3646 (N_3646,In_118,In_1634);
nor U3647 (N_3647,In_2575,In_2571);
xor U3648 (N_3648,In_2638,In_1280);
and U3649 (N_3649,In_2238,In_2484);
or U3650 (N_3650,In_1431,In_1320);
nor U3651 (N_3651,In_1965,In_2808);
nand U3652 (N_3652,In_795,In_1015);
or U3653 (N_3653,In_394,In_1342);
and U3654 (N_3654,In_453,In_1757);
and U3655 (N_3655,In_360,In_1836);
or U3656 (N_3656,In_2321,In_1965);
xor U3657 (N_3657,In_959,In_2619);
xnor U3658 (N_3658,In_1948,In_1180);
or U3659 (N_3659,In_1360,In_439);
nand U3660 (N_3660,In_1159,In_2937);
nand U3661 (N_3661,In_2414,In_2392);
or U3662 (N_3662,In_2452,In_1034);
or U3663 (N_3663,In_1221,In_888);
nor U3664 (N_3664,In_1021,In_1412);
or U3665 (N_3665,In_2158,In_1850);
xnor U3666 (N_3666,In_823,In_1001);
nand U3667 (N_3667,In_682,In_1737);
and U3668 (N_3668,In_2229,In_436);
and U3669 (N_3669,In_1462,In_2691);
nor U3670 (N_3670,In_379,In_103);
nor U3671 (N_3671,In_2447,In_2085);
nor U3672 (N_3672,In_2480,In_689);
xnor U3673 (N_3673,In_908,In_2693);
nor U3674 (N_3674,In_770,In_2765);
xor U3675 (N_3675,In_1400,In_80);
nor U3676 (N_3676,In_888,In_1243);
or U3677 (N_3677,In_322,In_2603);
nand U3678 (N_3678,In_2440,In_2384);
nand U3679 (N_3679,In_1134,In_2493);
and U3680 (N_3680,In_1942,In_649);
nor U3681 (N_3681,In_2631,In_1028);
or U3682 (N_3682,In_1070,In_2049);
or U3683 (N_3683,In_1763,In_2565);
and U3684 (N_3684,In_2435,In_2727);
xor U3685 (N_3685,In_2203,In_2486);
xor U3686 (N_3686,In_2839,In_2778);
nor U3687 (N_3687,In_490,In_2801);
nand U3688 (N_3688,In_1989,In_559);
and U3689 (N_3689,In_2570,In_1764);
or U3690 (N_3690,In_2796,In_2546);
nor U3691 (N_3691,In_2483,In_1388);
nor U3692 (N_3692,In_2556,In_1465);
nand U3693 (N_3693,In_1805,In_1646);
or U3694 (N_3694,In_36,In_246);
xnor U3695 (N_3695,In_70,In_2821);
or U3696 (N_3696,In_607,In_1979);
nand U3697 (N_3697,In_1657,In_2659);
and U3698 (N_3698,In_545,In_1230);
or U3699 (N_3699,In_464,In_514);
or U3700 (N_3700,In_2403,In_1913);
nand U3701 (N_3701,In_959,In_876);
xnor U3702 (N_3702,In_313,In_2236);
xnor U3703 (N_3703,In_54,In_1965);
nand U3704 (N_3704,In_247,In_1982);
nor U3705 (N_3705,In_1113,In_436);
and U3706 (N_3706,In_675,In_2123);
nand U3707 (N_3707,In_512,In_841);
nor U3708 (N_3708,In_599,In_2029);
nor U3709 (N_3709,In_1593,In_797);
nand U3710 (N_3710,In_29,In_2175);
and U3711 (N_3711,In_2758,In_661);
nor U3712 (N_3712,In_909,In_2596);
xnor U3713 (N_3713,In_112,In_2570);
nor U3714 (N_3714,In_599,In_2420);
or U3715 (N_3715,In_1296,In_1021);
xnor U3716 (N_3716,In_2816,In_1721);
nand U3717 (N_3717,In_211,In_1356);
xnor U3718 (N_3718,In_2544,In_1638);
nand U3719 (N_3719,In_84,In_2406);
nor U3720 (N_3720,In_1997,In_1781);
or U3721 (N_3721,In_2331,In_980);
xor U3722 (N_3722,In_127,In_1479);
nor U3723 (N_3723,In_1507,In_2784);
nand U3724 (N_3724,In_456,In_1990);
nor U3725 (N_3725,In_510,In_2400);
xnor U3726 (N_3726,In_2086,In_2880);
nor U3727 (N_3727,In_2196,In_231);
and U3728 (N_3728,In_1053,In_2315);
nor U3729 (N_3729,In_1082,In_93);
and U3730 (N_3730,In_1151,In_2611);
xor U3731 (N_3731,In_2181,In_2502);
nor U3732 (N_3732,In_1107,In_1989);
nand U3733 (N_3733,In_2169,In_1863);
and U3734 (N_3734,In_1970,In_679);
nand U3735 (N_3735,In_2565,In_2006);
and U3736 (N_3736,In_1820,In_2579);
and U3737 (N_3737,In_210,In_162);
and U3738 (N_3738,In_1058,In_2810);
or U3739 (N_3739,In_2975,In_198);
nand U3740 (N_3740,In_1906,In_1507);
and U3741 (N_3741,In_739,In_1638);
xnor U3742 (N_3742,In_2378,In_679);
and U3743 (N_3743,In_1080,In_2149);
or U3744 (N_3744,In_2768,In_2455);
nand U3745 (N_3745,In_1090,In_876);
and U3746 (N_3746,In_108,In_1456);
and U3747 (N_3747,In_787,In_849);
and U3748 (N_3748,In_1328,In_1187);
and U3749 (N_3749,In_1323,In_2813);
nor U3750 (N_3750,In_2585,In_844);
and U3751 (N_3751,In_661,In_2970);
nor U3752 (N_3752,In_1878,In_188);
or U3753 (N_3753,In_2059,In_687);
or U3754 (N_3754,In_1592,In_2740);
and U3755 (N_3755,In_1442,In_265);
or U3756 (N_3756,In_1005,In_751);
nor U3757 (N_3757,In_174,In_107);
nor U3758 (N_3758,In_2188,In_2293);
and U3759 (N_3759,In_1592,In_960);
and U3760 (N_3760,In_1813,In_1382);
or U3761 (N_3761,In_1454,In_1832);
or U3762 (N_3762,In_444,In_1884);
nor U3763 (N_3763,In_1875,In_1606);
nand U3764 (N_3764,In_548,In_1010);
or U3765 (N_3765,In_7,In_708);
nand U3766 (N_3766,In_1162,In_829);
or U3767 (N_3767,In_1093,In_2155);
nand U3768 (N_3768,In_2466,In_476);
or U3769 (N_3769,In_1038,In_2896);
nor U3770 (N_3770,In_2986,In_1543);
or U3771 (N_3771,In_577,In_2970);
and U3772 (N_3772,In_1953,In_1021);
nand U3773 (N_3773,In_300,In_1557);
nand U3774 (N_3774,In_845,In_1751);
and U3775 (N_3775,In_2220,In_2990);
or U3776 (N_3776,In_447,In_2745);
nor U3777 (N_3777,In_1334,In_1722);
or U3778 (N_3778,In_2877,In_1653);
nor U3779 (N_3779,In_103,In_140);
nand U3780 (N_3780,In_644,In_2035);
xnor U3781 (N_3781,In_1935,In_2841);
xor U3782 (N_3782,In_1452,In_1578);
and U3783 (N_3783,In_45,In_2096);
and U3784 (N_3784,In_2296,In_2181);
nor U3785 (N_3785,In_450,In_285);
or U3786 (N_3786,In_2314,In_1500);
nor U3787 (N_3787,In_1639,In_1904);
nor U3788 (N_3788,In_2473,In_1601);
or U3789 (N_3789,In_2931,In_1308);
nor U3790 (N_3790,In_2030,In_1266);
nand U3791 (N_3791,In_1955,In_2032);
nor U3792 (N_3792,In_2749,In_523);
xor U3793 (N_3793,In_2913,In_1874);
and U3794 (N_3794,In_567,In_1267);
nor U3795 (N_3795,In_1024,In_1270);
nor U3796 (N_3796,In_57,In_508);
nor U3797 (N_3797,In_2875,In_1283);
nor U3798 (N_3798,In_479,In_837);
or U3799 (N_3799,In_293,In_851);
or U3800 (N_3800,In_98,In_361);
nor U3801 (N_3801,In_118,In_2207);
or U3802 (N_3802,In_918,In_1111);
or U3803 (N_3803,In_1282,In_814);
and U3804 (N_3804,In_1571,In_2106);
nand U3805 (N_3805,In_1863,In_2766);
nor U3806 (N_3806,In_2093,In_1592);
xor U3807 (N_3807,In_2114,In_2309);
or U3808 (N_3808,In_1400,In_2674);
and U3809 (N_3809,In_1771,In_1016);
xnor U3810 (N_3810,In_57,In_886);
nand U3811 (N_3811,In_1398,In_2268);
nand U3812 (N_3812,In_1635,In_813);
xnor U3813 (N_3813,In_596,In_2554);
nand U3814 (N_3814,In_484,In_77);
nor U3815 (N_3815,In_518,In_827);
xnor U3816 (N_3816,In_1070,In_747);
and U3817 (N_3817,In_1076,In_336);
nor U3818 (N_3818,In_2514,In_186);
nand U3819 (N_3819,In_2723,In_1456);
nor U3820 (N_3820,In_1306,In_2756);
or U3821 (N_3821,In_2545,In_1835);
and U3822 (N_3822,In_1811,In_189);
nand U3823 (N_3823,In_1733,In_133);
xnor U3824 (N_3824,In_19,In_1761);
and U3825 (N_3825,In_1109,In_121);
and U3826 (N_3826,In_1125,In_702);
or U3827 (N_3827,In_716,In_487);
xor U3828 (N_3828,In_792,In_2032);
nand U3829 (N_3829,In_860,In_696);
nor U3830 (N_3830,In_216,In_1787);
xor U3831 (N_3831,In_1509,In_2053);
or U3832 (N_3832,In_2156,In_1857);
nor U3833 (N_3833,In_1885,In_2023);
or U3834 (N_3834,In_666,In_2377);
nor U3835 (N_3835,In_785,In_2423);
or U3836 (N_3836,In_586,In_161);
nor U3837 (N_3837,In_563,In_715);
nor U3838 (N_3838,In_37,In_2527);
nand U3839 (N_3839,In_870,In_2270);
xor U3840 (N_3840,In_733,In_932);
and U3841 (N_3841,In_809,In_513);
and U3842 (N_3842,In_1208,In_1372);
and U3843 (N_3843,In_2559,In_2766);
nor U3844 (N_3844,In_2719,In_629);
nand U3845 (N_3845,In_1410,In_1952);
xnor U3846 (N_3846,In_818,In_1268);
nand U3847 (N_3847,In_1419,In_2179);
nor U3848 (N_3848,In_828,In_1427);
nand U3849 (N_3849,In_2039,In_778);
xnor U3850 (N_3850,In_1066,In_2745);
nand U3851 (N_3851,In_44,In_421);
or U3852 (N_3852,In_1443,In_69);
or U3853 (N_3853,In_1358,In_2735);
nor U3854 (N_3854,In_908,In_1695);
and U3855 (N_3855,In_57,In_2285);
nor U3856 (N_3856,In_2896,In_951);
nand U3857 (N_3857,In_1457,In_1629);
and U3858 (N_3858,In_2292,In_568);
nor U3859 (N_3859,In_206,In_2540);
and U3860 (N_3860,In_860,In_1555);
nand U3861 (N_3861,In_179,In_1265);
nand U3862 (N_3862,In_1832,In_2841);
and U3863 (N_3863,In_664,In_1511);
nor U3864 (N_3864,In_2735,In_1730);
or U3865 (N_3865,In_523,In_1538);
nand U3866 (N_3866,In_2338,In_2154);
xnor U3867 (N_3867,In_1414,In_2849);
nand U3868 (N_3868,In_2637,In_652);
or U3869 (N_3869,In_1270,In_2493);
xor U3870 (N_3870,In_2305,In_522);
nor U3871 (N_3871,In_749,In_1290);
or U3872 (N_3872,In_2188,In_1706);
or U3873 (N_3873,In_1266,In_2054);
nand U3874 (N_3874,In_2430,In_1149);
nand U3875 (N_3875,In_1201,In_1343);
nor U3876 (N_3876,In_934,In_2854);
nor U3877 (N_3877,In_1284,In_2071);
xnor U3878 (N_3878,In_2463,In_1236);
nand U3879 (N_3879,In_2065,In_2483);
nor U3880 (N_3880,In_1661,In_2181);
nand U3881 (N_3881,In_1664,In_2734);
and U3882 (N_3882,In_1402,In_1810);
or U3883 (N_3883,In_1043,In_2737);
and U3884 (N_3884,In_548,In_1538);
nor U3885 (N_3885,In_2679,In_474);
or U3886 (N_3886,In_1914,In_227);
xor U3887 (N_3887,In_123,In_665);
and U3888 (N_3888,In_330,In_2522);
nand U3889 (N_3889,In_1607,In_2305);
or U3890 (N_3890,In_1384,In_394);
nand U3891 (N_3891,In_2609,In_19);
nand U3892 (N_3892,In_2046,In_1057);
nor U3893 (N_3893,In_2802,In_1489);
and U3894 (N_3894,In_1905,In_355);
nand U3895 (N_3895,In_2087,In_2070);
nor U3896 (N_3896,In_1611,In_882);
and U3897 (N_3897,In_1024,In_1161);
or U3898 (N_3898,In_1598,In_1117);
nor U3899 (N_3899,In_1498,In_994);
and U3900 (N_3900,In_1091,In_70);
and U3901 (N_3901,In_2257,In_539);
and U3902 (N_3902,In_765,In_1445);
nor U3903 (N_3903,In_2159,In_269);
nand U3904 (N_3904,In_2498,In_1185);
xor U3905 (N_3905,In_2246,In_1668);
nand U3906 (N_3906,In_1825,In_1667);
and U3907 (N_3907,In_1982,In_731);
xnor U3908 (N_3908,In_2586,In_1908);
xor U3909 (N_3909,In_723,In_2568);
nand U3910 (N_3910,In_2069,In_2218);
or U3911 (N_3911,In_2681,In_1118);
nand U3912 (N_3912,In_220,In_2304);
nand U3913 (N_3913,In_2064,In_600);
nor U3914 (N_3914,In_2673,In_918);
nor U3915 (N_3915,In_375,In_1866);
or U3916 (N_3916,In_1258,In_1491);
nand U3917 (N_3917,In_2794,In_223);
or U3918 (N_3918,In_506,In_1186);
nor U3919 (N_3919,In_735,In_1639);
xor U3920 (N_3920,In_2449,In_147);
nand U3921 (N_3921,In_2453,In_1007);
nor U3922 (N_3922,In_1707,In_2475);
nor U3923 (N_3923,In_36,In_2406);
nor U3924 (N_3924,In_256,In_1771);
or U3925 (N_3925,In_2566,In_442);
or U3926 (N_3926,In_534,In_2930);
nand U3927 (N_3927,In_2727,In_1615);
nor U3928 (N_3928,In_2082,In_2459);
and U3929 (N_3929,In_1645,In_1947);
and U3930 (N_3930,In_2930,In_644);
or U3931 (N_3931,In_2852,In_1334);
nor U3932 (N_3932,In_1220,In_2477);
nor U3933 (N_3933,In_1719,In_1099);
and U3934 (N_3934,In_1475,In_389);
and U3935 (N_3935,In_2163,In_1223);
or U3936 (N_3936,In_2198,In_1268);
or U3937 (N_3937,In_2630,In_2008);
nand U3938 (N_3938,In_346,In_2140);
nor U3939 (N_3939,In_1288,In_343);
nand U3940 (N_3940,In_1052,In_1957);
nand U3941 (N_3941,In_1467,In_1743);
nand U3942 (N_3942,In_2170,In_555);
or U3943 (N_3943,In_2516,In_2671);
nor U3944 (N_3944,In_846,In_140);
or U3945 (N_3945,In_1630,In_1235);
xor U3946 (N_3946,In_880,In_2602);
and U3947 (N_3947,In_1627,In_41);
nor U3948 (N_3948,In_1270,In_2179);
or U3949 (N_3949,In_137,In_2514);
nor U3950 (N_3950,In_1981,In_754);
and U3951 (N_3951,In_1471,In_325);
and U3952 (N_3952,In_2206,In_1498);
nand U3953 (N_3953,In_596,In_100);
nor U3954 (N_3954,In_1271,In_2545);
nand U3955 (N_3955,In_2724,In_91);
or U3956 (N_3956,In_1172,In_117);
and U3957 (N_3957,In_1072,In_517);
xnor U3958 (N_3958,In_562,In_2738);
nor U3959 (N_3959,In_1318,In_2307);
or U3960 (N_3960,In_14,In_2267);
or U3961 (N_3961,In_530,In_1239);
and U3962 (N_3962,In_748,In_305);
xnor U3963 (N_3963,In_1303,In_1205);
and U3964 (N_3964,In_473,In_463);
nor U3965 (N_3965,In_1501,In_1145);
or U3966 (N_3966,In_1844,In_1195);
nand U3967 (N_3967,In_2590,In_2791);
or U3968 (N_3968,In_1078,In_2323);
nand U3969 (N_3969,In_1281,In_2257);
or U3970 (N_3970,In_461,In_2918);
or U3971 (N_3971,In_2108,In_624);
or U3972 (N_3972,In_2194,In_2144);
or U3973 (N_3973,In_104,In_825);
nand U3974 (N_3974,In_103,In_2540);
nor U3975 (N_3975,In_1280,In_2602);
and U3976 (N_3976,In_2228,In_1230);
and U3977 (N_3977,In_1539,In_649);
xor U3978 (N_3978,In_1500,In_1032);
nand U3979 (N_3979,In_1261,In_868);
or U3980 (N_3980,In_1903,In_682);
and U3981 (N_3981,In_630,In_382);
and U3982 (N_3982,In_2157,In_1893);
and U3983 (N_3983,In_11,In_833);
or U3984 (N_3984,In_1865,In_544);
or U3985 (N_3985,In_56,In_1376);
and U3986 (N_3986,In_2795,In_2227);
nor U3987 (N_3987,In_2745,In_335);
and U3988 (N_3988,In_1573,In_1737);
and U3989 (N_3989,In_1531,In_1114);
and U3990 (N_3990,In_536,In_974);
nand U3991 (N_3991,In_93,In_408);
xnor U3992 (N_3992,In_2042,In_2740);
or U3993 (N_3993,In_805,In_596);
xnor U3994 (N_3994,In_550,In_310);
nor U3995 (N_3995,In_2173,In_483);
or U3996 (N_3996,In_879,In_2773);
nand U3997 (N_3997,In_2245,In_1246);
nand U3998 (N_3998,In_2690,In_374);
nand U3999 (N_3999,In_1566,In_2563);
nor U4000 (N_4000,In_378,In_1667);
or U4001 (N_4001,In_716,In_656);
or U4002 (N_4002,In_320,In_1630);
or U4003 (N_4003,In_958,In_1783);
nor U4004 (N_4004,In_595,In_1661);
nor U4005 (N_4005,In_2406,In_2940);
and U4006 (N_4006,In_23,In_1608);
nand U4007 (N_4007,In_227,In_1325);
or U4008 (N_4008,In_1003,In_1216);
or U4009 (N_4009,In_1142,In_175);
and U4010 (N_4010,In_759,In_158);
nor U4011 (N_4011,In_2378,In_2308);
and U4012 (N_4012,In_1971,In_2258);
or U4013 (N_4013,In_471,In_1509);
nor U4014 (N_4014,In_1648,In_1505);
and U4015 (N_4015,In_1740,In_1791);
and U4016 (N_4016,In_738,In_1022);
xnor U4017 (N_4017,In_2249,In_1381);
nand U4018 (N_4018,In_950,In_623);
xnor U4019 (N_4019,In_440,In_2208);
nor U4020 (N_4020,In_204,In_2491);
and U4021 (N_4021,In_655,In_98);
nor U4022 (N_4022,In_2565,In_1349);
xor U4023 (N_4023,In_1310,In_2109);
nor U4024 (N_4024,In_1392,In_2542);
nand U4025 (N_4025,In_1911,In_1485);
nand U4026 (N_4026,In_596,In_1000);
and U4027 (N_4027,In_527,In_387);
and U4028 (N_4028,In_95,In_2419);
nand U4029 (N_4029,In_270,In_2794);
and U4030 (N_4030,In_2219,In_2311);
and U4031 (N_4031,In_648,In_839);
and U4032 (N_4032,In_2157,In_610);
and U4033 (N_4033,In_2509,In_325);
nand U4034 (N_4034,In_2104,In_192);
or U4035 (N_4035,In_2151,In_1368);
or U4036 (N_4036,In_923,In_1624);
xor U4037 (N_4037,In_1088,In_1708);
nor U4038 (N_4038,In_147,In_2922);
or U4039 (N_4039,In_2198,In_2361);
and U4040 (N_4040,In_9,In_1045);
or U4041 (N_4041,In_2166,In_553);
and U4042 (N_4042,In_1928,In_964);
nand U4043 (N_4043,In_2661,In_265);
xor U4044 (N_4044,In_342,In_325);
nand U4045 (N_4045,In_545,In_1154);
nor U4046 (N_4046,In_1552,In_1555);
nand U4047 (N_4047,In_2997,In_1592);
nor U4048 (N_4048,In_1891,In_2610);
xor U4049 (N_4049,In_1450,In_425);
or U4050 (N_4050,In_1230,In_2812);
xor U4051 (N_4051,In_2796,In_1010);
or U4052 (N_4052,In_1629,In_2130);
nand U4053 (N_4053,In_2797,In_1820);
xnor U4054 (N_4054,In_1288,In_1825);
xor U4055 (N_4055,In_2674,In_1497);
or U4056 (N_4056,In_2858,In_222);
or U4057 (N_4057,In_1291,In_2850);
xnor U4058 (N_4058,In_2359,In_2071);
nor U4059 (N_4059,In_2975,In_2315);
and U4060 (N_4060,In_2823,In_1445);
and U4061 (N_4061,In_1797,In_68);
nor U4062 (N_4062,In_1284,In_2497);
nand U4063 (N_4063,In_2481,In_2240);
and U4064 (N_4064,In_2117,In_1747);
and U4065 (N_4065,In_2672,In_841);
nor U4066 (N_4066,In_2005,In_1981);
nand U4067 (N_4067,In_829,In_2347);
and U4068 (N_4068,In_221,In_2530);
nor U4069 (N_4069,In_115,In_2497);
nand U4070 (N_4070,In_823,In_2467);
nor U4071 (N_4071,In_1896,In_1588);
nand U4072 (N_4072,In_492,In_948);
or U4073 (N_4073,In_947,In_1824);
and U4074 (N_4074,In_2732,In_2191);
nor U4075 (N_4075,In_1916,In_544);
nand U4076 (N_4076,In_1334,In_1871);
and U4077 (N_4077,In_1120,In_808);
nand U4078 (N_4078,In_1212,In_452);
xnor U4079 (N_4079,In_1297,In_1190);
or U4080 (N_4080,In_1104,In_980);
or U4081 (N_4081,In_2151,In_985);
xor U4082 (N_4082,In_101,In_1974);
or U4083 (N_4083,In_2970,In_440);
and U4084 (N_4084,In_1125,In_2205);
nand U4085 (N_4085,In_706,In_70);
nor U4086 (N_4086,In_1001,In_1876);
nand U4087 (N_4087,In_2073,In_50);
nand U4088 (N_4088,In_474,In_1463);
xor U4089 (N_4089,In_1947,In_1637);
or U4090 (N_4090,In_1790,In_1825);
and U4091 (N_4091,In_1691,In_2770);
nand U4092 (N_4092,In_2501,In_302);
nand U4093 (N_4093,In_437,In_1225);
or U4094 (N_4094,In_46,In_2677);
nor U4095 (N_4095,In_2946,In_2919);
nor U4096 (N_4096,In_1682,In_2734);
or U4097 (N_4097,In_2483,In_1229);
nor U4098 (N_4098,In_223,In_495);
or U4099 (N_4099,In_2999,In_647);
and U4100 (N_4100,In_837,In_1513);
or U4101 (N_4101,In_609,In_557);
and U4102 (N_4102,In_1273,In_884);
nor U4103 (N_4103,In_2647,In_913);
or U4104 (N_4104,In_272,In_2223);
and U4105 (N_4105,In_291,In_1214);
and U4106 (N_4106,In_915,In_535);
xor U4107 (N_4107,In_677,In_1009);
and U4108 (N_4108,In_2974,In_1760);
nor U4109 (N_4109,In_653,In_2338);
and U4110 (N_4110,In_1589,In_178);
or U4111 (N_4111,In_2335,In_783);
nand U4112 (N_4112,In_1014,In_147);
and U4113 (N_4113,In_7,In_1465);
nor U4114 (N_4114,In_2358,In_1862);
nor U4115 (N_4115,In_1538,In_86);
or U4116 (N_4116,In_1953,In_2961);
and U4117 (N_4117,In_906,In_2991);
or U4118 (N_4118,In_2246,In_1948);
or U4119 (N_4119,In_877,In_2102);
nor U4120 (N_4120,In_1796,In_54);
nand U4121 (N_4121,In_1343,In_365);
or U4122 (N_4122,In_1293,In_2687);
nor U4123 (N_4123,In_788,In_783);
nand U4124 (N_4124,In_829,In_476);
and U4125 (N_4125,In_593,In_1584);
and U4126 (N_4126,In_2496,In_2167);
and U4127 (N_4127,In_623,In_1433);
and U4128 (N_4128,In_373,In_2031);
and U4129 (N_4129,In_1333,In_1901);
xnor U4130 (N_4130,In_985,In_1491);
or U4131 (N_4131,In_2642,In_2461);
or U4132 (N_4132,In_1750,In_55);
or U4133 (N_4133,In_1154,In_661);
and U4134 (N_4134,In_382,In_1244);
and U4135 (N_4135,In_1009,In_2115);
xnor U4136 (N_4136,In_2917,In_15);
nor U4137 (N_4137,In_1392,In_2329);
or U4138 (N_4138,In_302,In_139);
nand U4139 (N_4139,In_822,In_160);
nand U4140 (N_4140,In_148,In_2726);
xor U4141 (N_4141,In_593,In_1553);
xor U4142 (N_4142,In_1809,In_1705);
nor U4143 (N_4143,In_1468,In_2158);
and U4144 (N_4144,In_160,In_2160);
and U4145 (N_4145,In_340,In_327);
nand U4146 (N_4146,In_2921,In_850);
nor U4147 (N_4147,In_1365,In_1667);
nand U4148 (N_4148,In_2081,In_1154);
nand U4149 (N_4149,In_874,In_502);
nor U4150 (N_4150,In_1196,In_1874);
nand U4151 (N_4151,In_669,In_2675);
xnor U4152 (N_4152,In_2476,In_390);
and U4153 (N_4153,In_1622,In_1838);
nand U4154 (N_4154,In_2950,In_2108);
and U4155 (N_4155,In_2151,In_2769);
or U4156 (N_4156,In_1809,In_120);
nor U4157 (N_4157,In_1383,In_1256);
nand U4158 (N_4158,In_1818,In_571);
nand U4159 (N_4159,In_793,In_2737);
nand U4160 (N_4160,In_1552,In_1895);
and U4161 (N_4161,In_127,In_1056);
and U4162 (N_4162,In_1206,In_1229);
nand U4163 (N_4163,In_169,In_643);
nand U4164 (N_4164,In_2693,In_2880);
or U4165 (N_4165,In_2377,In_1786);
nand U4166 (N_4166,In_849,In_1234);
nor U4167 (N_4167,In_51,In_2559);
nand U4168 (N_4168,In_2859,In_467);
nand U4169 (N_4169,In_2646,In_179);
nor U4170 (N_4170,In_1359,In_2020);
and U4171 (N_4171,In_78,In_750);
xor U4172 (N_4172,In_2669,In_2097);
and U4173 (N_4173,In_2443,In_701);
nand U4174 (N_4174,In_2962,In_1038);
xor U4175 (N_4175,In_2565,In_2236);
nand U4176 (N_4176,In_426,In_1367);
nand U4177 (N_4177,In_1288,In_2490);
nand U4178 (N_4178,In_2933,In_1611);
and U4179 (N_4179,In_938,In_2881);
and U4180 (N_4180,In_1922,In_1373);
or U4181 (N_4181,In_130,In_296);
nand U4182 (N_4182,In_2159,In_1635);
nand U4183 (N_4183,In_127,In_1700);
nor U4184 (N_4184,In_791,In_2301);
nand U4185 (N_4185,In_2156,In_2307);
nor U4186 (N_4186,In_2640,In_2862);
or U4187 (N_4187,In_1233,In_2438);
and U4188 (N_4188,In_423,In_2623);
nand U4189 (N_4189,In_2194,In_813);
or U4190 (N_4190,In_518,In_2969);
or U4191 (N_4191,In_1692,In_2098);
nand U4192 (N_4192,In_2010,In_2281);
nor U4193 (N_4193,In_2557,In_2991);
or U4194 (N_4194,In_815,In_899);
nand U4195 (N_4195,In_1724,In_2113);
xor U4196 (N_4196,In_1049,In_1831);
or U4197 (N_4197,In_307,In_1502);
or U4198 (N_4198,In_631,In_1477);
nor U4199 (N_4199,In_1274,In_2033);
or U4200 (N_4200,In_653,In_549);
or U4201 (N_4201,In_239,In_1423);
and U4202 (N_4202,In_2231,In_456);
or U4203 (N_4203,In_1259,In_676);
and U4204 (N_4204,In_171,In_1403);
or U4205 (N_4205,In_2784,In_994);
nand U4206 (N_4206,In_406,In_1603);
nand U4207 (N_4207,In_2518,In_2980);
nor U4208 (N_4208,In_2347,In_1216);
nand U4209 (N_4209,In_2038,In_2914);
nand U4210 (N_4210,In_1616,In_25);
nand U4211 (N_4211,In_1526,In_2573);
nand U4212 (N_4212,In_456,In_1333);
and U4213 (N_4213,In_1985,In_174);
and U4214 (N_4214,In_1292,In_93);
nand U4215 (N_4215,In_2280,In_1638);
and U4216 (N_4216,In_2507,In_947);
and U4217 (N_4217,In_2287,In_2817);
nand U4218 (N_4218,In_1671,In_339);
or U4219 (N_4219,In_2257,In_380);
or U4220 (N_4220,In_2509,In_355);
and U4221 (N_4221,In_203,In_2680);
or U4222 (N_4222,In_677,In_2695);
and U4223 (N_4223,In_731,In_1868);
and U4224 (N_4224,In_1263,In_1840);
nor U4225 (N_4225,In_36,In_1566);
nand U4226 (N_4226,In_2945,In_679);
nor U4227 (N_4227,In_1046,In_2144);
or U4228 (N_4228,In_1977,In_2217);
nor U4229 (N_4229,In_2903,In_101);
xor U4230 (N_4230,In_2098,In_212);
nand U4231 (N_4231,In_2713,In_2578);
or U4232 (N_4232,In_2774,In_1394);
nand U4233 (N_4233,In_2357,In_2144);
nand U4234 (N_4234,In_1796,In_913);
and U4235 (N_4235,In_687,In_1505);
nor U4236 (N_4236,In_2027,In_107);
nand U4237 (N_4237,In_15,In_621);
and U4238 (N_4238,In_804,In_2196);
and U4239 (N_4239,In_2196,In_2393);
and U4240 (N_4240,In_2722,In_388);
nand U4241 (N_4241,In_2926,In_1617);
or U4242 (N_4242,In_2802,In_344);
and U4243 (N_4243,In_1721,In_2349);
nand U4244 (N_4244,In_1806,In_164);
nor U4245 (N_4245,In_868,In_799);
nand U4246 (N_4246,In_43,In_114);
nand U4247 (N_4247,In_378,In_2007);
and U4248 (N_4248,In_1333,In_1621);
or U4249 (N_4249,In_1889,In_819);
nand U4250 (N_4250,In_1814,In_2056);
or U4251 (N_4251,In_1176,In_1962);
or U4252 (N_4252,In_64,In_2225);
nand U4253 (N_4253,In_2527,In_2246);
nand U4254 (N_4254,In_34,In_256);
or U4255 (N_4255,In_1492,In_1961);
and U4256 (N_4256,In_2511,In_2911);
and U4257 (N_4257,In_2061,In_358);
nor U4258 (N_4258,In_1234,In_2811);
or U4259 (N_4259,In_1085,In_2641);
nand U4260 (N_4260,In_2315,In_2746);
nand U4261 (N_4261,In_1339,In_2598);
or U4262 (N_4262,In_1882,In_2802);
nand U4263 (N_4263,In_2892,In_2980);
nand U4264 (N_4264,In_2766,In_2765);
xnor U4265 (N_4265,In_135,In_2399);
nand U4266 (N_4266,In_407,In_1952);
nand U4267 (N_4267,In_2299,In_2074);
xnor U4268 (N_4268,In_14,In_1572);
and U4269 (N_4269,In_1261,In_2750);
nand U4270 (N_4270,In_2928,In_739);
or U4271 (N_4271,In_1628,In_2439);
nand U4272 (N_4272,In_608,In_2774);
nand U4273 (N_4273,In_188,In_945);
and U4274 (N_4274,In_682,In_2379);
or U4275 (N_4275,In_1249,In_2435);
or U4276 (N_4276,In_495,In_2772);
nor U4277 (N_4277,In_943,In_662);
nor U4278 (N_4278,In_1044,In_2847);
and U4279 (N_4279,In_920,In_2838);
and U4280 (N_4280,In_1948,In_919);
nand U4281 (N_4281,In_1158,In_2449);
xnor U4282 (N_4282,In_2983,In_1009);
and U4283 (N_4283,In_1065,In_827);
nand U4284 (N_4284,In_2848,In_2232);
and U4285 (N_4285,In_2541,In_1260);
and U4286 (N_4286,In_411,In_2800);
nor U4287 (N_4287,In_553,In_1591);
or U4288 (N_4288,In_2837,In_1833);
and U4289 (N_4289,In_2046,In_1195);
or U4290 (N_4290,In_2505,In_502);
nand U4291 (N_4291,In_1963,In_1470);
nand U4292 (N_4292,In_306,In_2525);
nand U4293 (N_4293,In_2596,In_364);
nand U4294 (N_4294,In_2154,In_2144);
and U4295 (N_4295,In_1906,In_884);
and U4296 (N_4296,In_2863,In_1070);
and U4297 (N_4297,In_1257,In_1383);
nor U4298 (N_4298,In_362,In_1429);
and U4299 (N_4299,In_1802,In_2941);
nand U4300 (N_4300,In_1652,In_946);
nand U4301 (N_4301,In_764,In_2230);
xor U4302 (N_4302,In_1281,In_1046);
nand U4303 (N_4303,In_622,In_529);
nand U4304 (N_4304,In_1952,In_2078);
xor U4305 (N_4305,In_22,In_1265);
and U4306 (N_4306,In_949,In_1082);
nor U4307 (N_4307,In_764,In_999);
or U4308 (N_4308,In_519,In_946);
and U4309 (N_4309,In_2224,In_2894);
and U4310 (N_4310,In_730,In_53);
xor U4311 (N_4311,In_2848,In_955);
or U4312 (N_4312,In_1403,In_491);
or U4313 (N_4313,In_757,In_222);
nand U4314 (N_4314,In_931,In_1937);
nand U4315 (N_4315,In_1055,In_1989);
and U4316 (N_4316,In_1970,In_2736);
or U4317 (N_4317,In_1971,In_1402);
or U4318 (N_4318,In_1769,In_2189);
nand U4319 (N_4319,In_1587,In_1751);
xnor U4320 (N_4320,In_101,In_2381);
nand U4321 (N_4321,In_1335,In_2151);
nor U4322 (N_4322,In_1744,In_2770);
xor U4323 (N_4323,In_894,In_2991);
nor U4324 (N_4324,In_1382,In_1080);
nand U4325 (N_4325,In_2257,In_10);
nor U4326 (N_4326,In_1097,In_1967);
or U4327 (N_4327,In_2503,In_2653);
nor U4328 (N_4328,In_2636,In_2363);
nand U4329 (N_4329,In_787,In_866);
nor U4330 (N_4330,In_2214,In_308);
or U4331 (N_4331,In_1073,In_1126);
nor U4332 (N_4332,In_2777,In_389);
and U4333 (N_4333,In_8,In_2261);
nor U4334 (N_4334,In_1061,In_1798);
nand U4335 (N_4335,In_2162,In_2149);
nor U4336 (N_4336,In_1251,In_424);
nor U4337 (N_4337,In_2889,In_600);
and U4338 (N_4338,In_1943,In_42);
and U4339 (N_4339,In_621,In_1698);
or U4340 (N_4340,In_2205,In_2192);
or U4341 (N_4341,In_274,In_2157);
nand U4342 (N_4342,In_2466,In_888);
xnor U4343 (N_4343,In_2068,In_2675);
nor U4344 (N_4344,In_2293,In_2746);
and U4345 (N_4345,In_2091,In_527);
or U4346 (N_4346,In_2997,In_361);
nor U4347 (N_4347,In_1433,In_1784);
nor U4348 (N_4348,In_501,In_2859);
nand U4349 (N_4349,In_2871,In_1557);
or U4350 (N_4350,In_2865,In_2752);
nor U4351 (N_4351,In_151,In_1098);
nor U4352 (N_4352,In_1019,In_2869);
nor U4353 (N_4353,In_2181,In_133);
nand U4354 (N_4354,In_1583,In_176);
and U4355 (N_4355,In_1301,In_369);
xor U4356 (N_4356,In_2395,In_2409);
and U4357 (N_4357,In_475,In_2133);
nand U4358 (N_4358,In_1106,In_1451);
nor U4359 (N_4359,In_1206,In_1699);
nor U4360 (N_4360,In_803,In_2681);
or U4361 (N_4361,In_2096,In_239);
xnor U4362 (N_4362,In_1206,In_313);
nor U4363 (N_4363,In_1708,In_1575);
or U4364 (N_4364,In_1473,In_2062);
or U4365 (N_4365,In_1034,In_31);
nor U4366 (N_4366,In_1425,In_1483);
or U4367 (N_4367,In_490,In_1970);
nand U4368 (N_4368,In_36,In_2658);
nor U4369 (N_4369,In_1031,In_1085);
nand U4370 (N_4370,In_803,In_1768);
or U4371 (N_4371,In_2871,In_84);
nand U4372 (N_4372,In_2355,In_1771);
and U4373 (N_4373,In_194,In_196);
nand U4374 (N_4374,In_1076,In_575);
xnor U4375 (N_4375,In_2054,In_1059);
xnor U4376 (N_4376,In_1133,In_2902);
and U4377 (N_4377,In_428,In_1571);
and U4378 (N_4378,In_1870,In_1428);
nor U4379 (N_4379,In_1302,In_1112);
nor U4380 (N_4380,In_897,In_2621);
and U4381 (N_4381,In_1664,In_1341);
nand U4382 (N_4382,In_1505,In_475);
or U4383 (N_4383,In_1857,In_1093);
or U4384 (N_4384,In_1644,In_2632);
or U4385 (N_4385,In_2158,In_1758);
and U4386 (N_4386,In_1436,In_646);
nor U4387 (N_4387,In_1573,In_1483);
nand U4388 (N_4388,In_2035,In_1445);
or U4389 (N_4389,In_2870,In_2471);
xor U4390 (N_4390,In_1030,In_2648);
nor U4391 (N_4391,In_2379,In_2093);
and U4392 (N_4392,In_1644,In_543);
and U4393 (N_4393,In_1388,In_2330);
nand U4394 (N_4394,In_19,In_1217);
or U4395 (N_4395,In_1806,In_2617);
nand U4396 (N_4396,In_2071,In_1867);
or U4397 (N_4397,In_2565,In_1889);
and U4398 (N_4398,In_1719,In_824);
xor U4399 (N_4399,In_2310,In_769);
or U4400 (N_4400,In_1723,In_2879);
nand U4401 (N_4401,In_1606,In_1650);
xor U4402 (N_4402,In_978,In_2753);
or U4403 (N_4403,In_1998,In_623);
or U4404 (N_4404,In_1947,In_841);
or U4405 (N_4405,In_2856,In_1048);
nor U4406 (N_4406,In_1017,In_863);
nand U4407 (N_4407,In_319,In_1402);
nand U4408 (N_4408,In_2753,In_551);
or U4409 (N_4409,In_1335,In_2152);
or U4410 (N_4410,In_2354,In_932);
nor U4411 (N_4411,In_1008,In_237);
and U4412 (N_4412,In_154,In_810);
or U4413 (N_4413,In_1536,In_2523);
nor U4414 (N_4414,In_2254,In_1608);
or U4415 (N_4415,In_860,In_1475);
nand U4416 (N_4416,In_1548,In_2800);
nor U4417 (N_4417,In_2667,In_2405);
and U4418 (N_4418,In_1129,In_2655);
nand U4419 (N_4419,In_1664,In_2325);
nor U4420 (N_4420,In_2235,In_1384);
or U4421 (N_4421,In_513,In_674);
nor U4422 (N_4422,In_104,In_722);
and U4423 (N_4423,In_2692,In_2613);
or U4424 (N_4424,In_1123,In_2812);
and U4425 (N_4425,In_601,In_2962);
nand U4426 (N_4426,In_402,In_1625);
nand U4427 (N_4427,In_123,In_2424);
and U4428 (N_4428,In_1465,In_2614);
or U4429 (N_4429,In_532,In_1764);
nor U4430 (N_4430,In_2695,In_2468);
xnor U4431 (N_4431,In_484,In_2886);
nand U4432 (N_4432,In_491,In_2393);
and U4433 (N_4433,In_1566,In_2841);
xnor U4434 (N_4434,In_2391,In_2798);
or U4435 (N_4435,In_2131,In_449);
and U4436 (N_4436,In_1993,In_47);
or U4437 (N_4437,In_1382,In_2973);
and U4438 (N_4438,In_2320,In_1525);
xnor U4439 (N_4439,In_482,In_2759);
nand U4440 (N_4440,In_927,In_1840);
nand U4441 (N_4441,In_1514,In_2521);
or U4442 (N_4442,In_322,In_2974);
nand U4443 (N_4443,In_2110,In_1407);
and U4444 (N_4444,In_2969,In_2627);
and U4445 (N_4445,In_1881,In_1776);
nor U4446 (N_4446,In_347,In_1762);
nand U4447 (N_4447,In_734,In_2541);
and U4448 (N_4448,In_2838,In_884);
nand U4449 (N_4449,In_1604,In_1473);
nor U4450 (N_4450,In_2526,In_221);
and U4451 (N_4451,In_2175,In_1529);
nand U4452 (N_4452,In_2071,In_1971);
xnor U4453 (N_4453,In_503,In_1945);
nor U4454 (N_4454,In_1140,In_406);
or U4455 (N_4455,In_1546,In_1949);
nand U4456 (N_4456,In_205,In_1721);
nand U4457 (N_4457,In_2065,In_829);
nor U4458 (N_4458,In_2471,In_817);
and U4459 (N_4459,In_216,In_2214);
xnor U4460 (N_4460,In_1701,In_2193);
nand U4461 (N_4461,In_2708,In_2189);
nor U4462 (N_4462,In_1132,In_371);
or U4463 (N_4463,In_1778,In_797);
nor U4464 (N_4464,In_2336,In_1480);
or U4465 (N_4465,In_1850,In_4);
and U4466 (N_4466,In_2797,In_293);
and U4467 (N_4467,In_2847,In_2504);
and U4468 (N_4468,In_2094,In_2921);
nand U4469 (N_4469,In_456,In_2046);
and U4470 (N_4470,In_1833,In_90);
and U4471 (N_4471,In_128,In_520);
xnor U4472 (N_4472,In_189,In_1780);
and U4473 (N_4473,In_1741,In_2395);
and U4474 (N_4474,In_1459,In_167);
or U4475 (N_4475,In_1947,In_1737);
nor U4476 (N_4476,In_401,In_1564);
nand U4477 (N_4477,In_2267,In_451);
or U4478 (N_4478,In_1446,In_522);
nor U4479 (N_4479,In_2362,In_1134);
or U4480 (N_4480,In_1720,In_1146);
xnor U4481 (N_4481,In_1324,In_658);
nand U4482 (N_4482,In_712,In_2601);
nor U4483 (N_4483,In_1760,In_667);
nand U4484 (N_4484,In_400,In_287);
and U4485 (N_4485,In_376,In_2123);
or U4486 (N_4486,In_2544,In_863);
nor U4487 (N_4487,In_342,In_2171);
and U4488 (N_4488,In_1430,In_961);
nor U4489 (N_4489,In_1143,In_190);
xnor U4490 (N_4490,In_1028,In_1675);
or U4491 (N_4491,In_2845,In_2014);
nand U4492 (N_4492,In_337,In_1548);
nor U4493 (N_4493,In_2620,In_1653);
nand U4494 (N_4494,In_2422,In_1106);
nor U4495 (N_4495,In_676,In_2276);
or U4496 (N_4496,In_1598,In_1066);
or U4497 (N_4497,In_2873,In_794);
xor U4498 (N_4498,In_1684,In_1677);
or U4499 (N_4499,In_2802,In_2671);
or U4500 (N_4500,In_1263,In_2925);
or U4501 (N_4501,In_2971,In_2757);
or U4502 (N_4502,In_1012,In_886);
and U4503 (N_4503,In_1227,In_482);
nor U4504 (N_4504,In_70,In_954);
nand U4505 (N_4505,In_2656,In_2446);
or U4506 (N_4506,In_1157,In_1638);
xnor U4507 (N_4507,In_1333,In_2905);
nor U4508 (N_4508,In_1285,In_252);
xnor U4509 (N_4509,In_2740,In_154);
nor U4510 (N_4510,In_734,In_1603);
nor U4511 (N_4511,In_1133,In_1065);
and U4512 (N_4512,In_2583,In_2550);
nor U4513 (N_4513,In_984,In_2788);
nand U4514 (N_4514,In_2369,In_1424);
xor U4515 (N_4515,In_2037,In_887);
and U4516 (N_4516,In_470,In_2958);
and U4517 (N_4517,In_2582,In_1096);
and U4518 (N_4518,In_943,In_957);
nand U4519 (N_4519,In_1047,In_1096);
or U4520 (N_4520,In_652,In_168);
nor U4521 (N_4521,In_1597,In_2677);
nand U4522 (N_4522,In_2814,In_2241);
nand U4523 (N_4523,In_191,In_401);
nor U4524 (N_4524,In_2330,In_1457);
nor U4525 (N_4525,In_2682,In_473);
nand U4526 (N_4526,In_1385,In_140);
xor U4527 (N_4527,In_2969,In_1371);
and U4528 (N_4528,In_254,In_1432);
nand U4529 (N_4529,In_2592,In_2804);
or U4530 (N_4530,In_1618,In_2873);
and U4531 (N_4531,In_2593,In_2542);
or U4532 (N_4532,In_1498,In_2505);
xor U4533 (N_4533,In_223,In_1191);
nand U4534 (N_4534,In_1533,In_456);
nand U4535 (N_4535,In_1038,In_2302);
nand U4536 (N_4536,In_918,In_1600);
nor U4537 (N_4537,In_1739,In_546);
xor U4538 (N_4538,In_1674,In_260);
nand U4539 (N_4539,In_67,In_1853);
or U4540 (N_4540,In_1426,In_1659);
nand U4541 (N_4541,In_1312,In_1114);
or U4542 (N_4542,In_2829,In_2854);
or U4543 (N_4543,In_157,In_2631);
and U4544 (N_4544,In_716,In_971);
nor U4545 (N_4545,In_118,In_472);
nand U4546 (N_4546,In_250,In_456);
or U4547 (N_4547,In_1276,In_2208);
and U4548 (N_4548,In_2647,In_1586);
nor U4549 (N_4549,In_240,In_2288);
and U4550 (N_4550,In_1723,In_2166);
nor U4551 (N_4551,In_2660,In_2772);
and U4552 (N_4552,In_2384,In_2706);
and U4553 (N_4553,In_439,In_1321);
nand U4554 (N_4554,In_1853,In_1873);
nand U4555 (N_4555,In_459,In_238);
nor U4556 (N_4556,In_1762,In_2174);
nand U4557 (N_4557,In_637,In_271);
xor U4558 (N_4558,In_2216,In_2972);
or U4559 (N_4559,In_2837,In_622);
nor U4560 (N_4560,In_2241,In_924);
nor U4561 (N_4561,In_1978,In_531);
nor U4562 (N_4562,In_2153,In_1305);
or U4563 (N_4563,In_2872,In_1353);
or U4564 (N_4564,In_1833,In_1854);
and U4565 (N_4565,In_703,In_2281);
or U4566 (N_4566,In_157,In_1354);
or U4567 (N_4567,In_2538,In_765);
nor U4568 (N_4568,In_1092,In_1162);
nand U4569 (N_4569,In_541,In_2481);
or U4570 (N_4570,In_2875,In_2277);
or U4571 (N_4571,In_754,In_2593);
nand U4572 (N_4572,In_311,In_2528);
nor U4573 (N_4573,In_2467,In_1339);
nand U4574 (N_4574,In_2966,In_2402);
nor U4575 (N_4575,In_2724,In_303);
nand U4576 (N_4576,In_1698,In_518);
or U4577 (N_4577,In_2593,In_2299);
and U4578 (N_4578,In_1517,In_2753);
and U4579 (N_4579,In_1387,In_1067);
xor U4580 (N_4580,In_70,In_2177);
xor U4581 (N_4581,In_845,In_2897);
nor U4582 (N_4582,In_1483,In_2601);
nand U4583 (N_4583,In_979,In_452);
or U4584 (N_4584,In_1350,In_1601);
nor U4585 (N_4585,In_1870,In_2050);
or U4586 (N_4586,In_2037,In_2515);
nand U4587 (N_4587,In_2177,In_1970);
nand U4588 (N_4588,In_1394,In_1932);
nor U4589 (N_4589,In_2421,In_2555);
nor U4590 (N_4590,In_570,In_2383);
nand U4591 (N_4591,In_387,In_1235);
or U4592 (N_4592,In_2698,In_2951);
nor U4593 (N_4593,In_2765,In_2676);
nor U4594 (N_4594,In_1954,In_1991);
and U4595 (N_4595,In_1045,In_656);
and U4596 (N_4596,In_2544,In_1412);
nand U4597 (N_4597,In_489,In_703);
xnor U4598 (N_4598,In_454,In_2470);
and U4599 (N_4599,In_2264,In_1596);
nand U4600 (N_4600,In_817,In_1603);
nor U4601 (N_4601,In_1952,In_914);
or U4602 (N_4602,In_2764,In_2832);
or U4603 (N_4603,In_903,In_233);
xnor U4604 (N_4604,In_190,In_713);
nor U4605 (N_4605,In_247,In_239);
xor U4606 (N_4606,In_2211,In_1044);
or U4607 (N_4607,In_1184,In_1103);
nor U4608 (N_4608,In_1465,In_2700);
and U4609 (N_4609,In_854,In_1081);
and U4610 (N_4610,In_182,In_1301);
and U4611 (N_4611,In_1192,In_96);
nor U4612 (N_4612,In_1430,In_1058);
nand U4613 (N_4613,In_2761,In_1024);
and U4614 (N_4614,In_1507,In_1289);
and U4615 (N_4615,In_1562,In_884);
and U4616 (N_4616,In_1929,In_173);
nor U4617 (N_4617,In_93,In_1179);
xnor U4618 (N_4618,In_1121,In_2645);
or U4619 (N_4619,In_1403,In_2719);
xnor U4620 (N_4620,In_2628,In_2344);
nor U4621 (N_4621,In_355,In_1591);
nor U4622 (N_4622,In_506,In_617);
or U4623 (N_4623,In_1974,In_2787);
or U4624 (N_4624,In_126,In_864);
nand U4625 (N_4625,In_2270,In_231);
nor U4626 (N_4626,In_1221,In_620);
and U4627 (N_4627,In_1209,In_1259);
or U4628 (N_4628,In_205,In_2005);
nor U4629 (N_4629,In_548,In_288);
or U4630 (N_4630,In_1904,In_633);
and U4631 (N_4631,In_834,In_2631);
nand U4632 (N_4632,In_2632,In_2466);
or U4633 (N_4633,In_1671,In_943);
xor U4634 (N_4634,In_1830,In_1611);
nor U4635 (N_4635,In_1930,In_942);
or U4636 (N_4636,In_25,In_1391);
or U4637 (N_4637,In_272,In_2288);
nor U4638 (N_4638,In_2110,In_405);
and U4639 (N_4639,In_2272,In_215);
xor U4640 (N_4640,In_2455,In_288);
and U4641 (N_4641,In_459,In_2862);
or U4642 (N_4642,In_924,In_1135);
nand U4643 (N_4643,In_750,In_1235);
nor U4644 (N_4644,In_56,In_1914);
xor U4645 (N_4645,In_1899,In_786);
nor U4646 (N_4646,In_1229,In_1809);
nor U4647 (N_4647,In_761,In_1151);
or U4648 (N_4648,In_1750,In_1476);
xnor U4649 (N_4649,In_2290,In_2026);
and U4650 (N_4650,In_273,In_2810);
or U4651 (N_4651,In_2186,In_1729);
xor U4652 (N_4652,In_2650,In_2062);
nand U4653 (N_4653,In_714,In_2247);
or U4654 (N_4654,In_1184,In_2702);
nand U4655 (N_4655,In_2038,In_932);
nand U4656 (N_4656,In_2697,In_2547);
nand U4657 (N_4657,In_777,In_201);
xor U4658 (N_4658,In_1125,In_2187);
nor U4659 (N_4659,In_2720,In_1115);
nand U4660 (N_4660,In_2629,In_2508);
nand U4661 (N_4661,In_258,In_496);
nor U4662 (N_4662,In_2378,In_1069);
xor U4663 (N_4663,In_20,In_1783);
nor U4664 (N_4664,In_2311,In_1509);
nand U4665 (N_4665,In_1285,In_332);
nand U4666 (N_4666,In_1654,In_815);
nor U4667 (N_4667,In_2380,In_1210);
or U4668 (N_4668,In_2385,In_1079);
or U4669 (N_4669,In_1890,In_2522);
nand U4670 (N_4670,In_121,In_2765);
nand U4671 (N_4671,In_2721,In_503);
xnor U4672 (N_4672,In_332,In_2232);
nor U4673 (N_4673,In_133,In_1327);
nor U4674 (N_4674,In_1081,In_100);
and U4675 (N_4675,In_2266,In_2855);
nand U4676 (N_4676,In_829,In_2216);
or U4677 (N_4677,In_1770,In_2395);
nand U4678 (N_4678,In_103,In_2359);
nor U4679 (N_4679,In_1438,In_2285);
or U4680 (N_4680,In_1386,In_561);
or U4681 (N_4681,In_1252,In_630);
nand U4682 (N_4682,In_1739,In_598);
nand U4683 (N_4683,In_2549,In_2873);
nor U4684 (N_4684,In_2918,In_1205);
nor U4685 (N_4685,In_1216,In_1520);
and U4686 (N_4686,In_2498,In_2010);
nand U4687 (N_4687,In_2505,In_2221);
or U4688 (N_4688,In_2403,In_2864);
nand U4689 (N_4689,In_2453,In_238);
nor U4690 (N_4690,In_398,In_1363);
nor U4691 (N_4691,In_1163,In_350);
nand U4692 (N_4692,In_2926,In_1907);
or U4693 (N_4693,In_709,In_1523);
and U4694 (N_4694,In_529,In_245);
nand U4695 (N_4695,In_2344,In_950);
and U4696 (N_4696,In_871,In_368);
nor U4697 (N_4697,In_1941,In_497);
or U4698 (N_4698,In_128,In_1951);
and U4699 (N_4699,In_2885,In_830);
nor U4700 (N_4700,In_2674,In_1137);
or U4701 (N_4701,In_2065,In_141);
nor U4702 (N_4702,In_1254,In_1415);
nand U4703 (N_4703,In_2782,In_1141);
nand U4704 (N_4704,In_2091,In_872);
nand U4705 (N_4705,In_1515,In_2536);
or U4706 (N_4706,In_352,In_1756);
or U4707 (N_4707,In_2920,In_2064);
nand U4708 (N_4708,In_598,In_1311);
xor U4709 (N_4709,In_1816,In_2560);
xnor U4710 (N_4710,In_2133,In_76);
or U4711 (N_4711,In_112,In_2650);
or U4712 (N_4712,In_897,In_1428);
nand U4713 (N_4713,In_2283,In_1947);
nand U4714 (N_4714,In_227,In_49);
or U4715 (N_4715,In_2130,In_942);
or U4716 (N_4716,In_2168,In_1664);
or U4717 (N_4717,In_2877,In_902);
nand U4718 (N_4718,In_1462,In_2778);
nand U4719 (N_4719,In_2866,In_472);
and U4720 (N_4720,In_932,In_1418);
and U4721 (N_4721,In_2709,In_2719);
or U4722 (N_4722,In_2278,In_1441);
and U4723 (N_4723,In_30,In_897);
and U4724 (N_4724,In_1444,In_2489);
nor U4725 (N_4725,In_2525,In_1687);
or U4726 (N_4726,In_2497,In_536);
or U4727 (N_4727,In_2816,In_1494);
xnor U4728 (N_4728,In_222,In_1932);
or U4729 (N_4729,In_403,In_2452);
xor U4730 (N_4730,In_269,In_2921);
nor U4731 (N_4731,In_2160,In_749);
nand U4732 (N_4732,In_1900,In_525);
nor U4733 (N_4733,In_1406,In_210);
nand U4734 (N_4734,In_1314,In_346);
xnor U4735 (N_4735,In_2905,In_1164);
nand U4736 (N_4736,In_1865,In_445);
and U4737 (N_4737,In_728,In_1239);
or U4738 (N_4738,In_1382,In_2359);
nor U4739 (N_4739,In_2537,In_2020);
or U4740 (N_4740,In_1598,In_1133);
and U4741 (N_4741,In_1581,In_1515);
nand U4742 (N_4742,In_2238,In_1112);
nor U4743 (N_4743,In_904,In_2923);
or U4744 (N_4744,In_2479,In_2521);
nor U4745 (N_4745,In_1977,In_1184);
nand U4746 (N_4746,In_1822,In_249);
nor U4747 (N_4747,In_2481,In_2471);
or U4748 (N_4748,In_1817,In_82);
nand U4749 (N_4749,In_945,In_2278);
or U4750 (N_4750,In_1936,In_1303);
nor U4751 (N_4751,In_1607,In_1106);
or U4752 (N_4752,In_1847,In_1348);
nor U4753 (N_4753,In_2739,In_2348);
nor U4754 (N_4754,In_690,In_2977);
and U4755 (N_4755,In_1176,In_53);
or U4756 (N_4756,In_132,In_1113);
nand U4757 (N_4757,In_775,In_434);
nand U4758 (N_4758,In_167,In_2458);
nor U4759 (N_4759,In_643,In_835);
or U4760 (N_4760,In_2896,In_357);
or U4761 (N_4761,In_1255,In_46);
and U4762 (N_4762,In_187,In_205);
or U4763 (N_4763,In_135,In_300);
nand U4764 (N_4764,In_734,In_1928);
and U4765 (N_4765,In_519,In_814);
and U4766 (N_4766,In_98,In_2822);
nor U4767 (N_4767,In_1199,In_1852);
and U4768 (N_4768,In_600,In_1021);
and U4769 (N_4769,In_1719,In_984);
nor U4770 (N_4770,In_101,In_977);
nor U4771 (N_4771,In_1243,In_944);
nor U4772 (N_4772,In_830,In_2854);
nand U4773 (N_4773,In_636,In_919);
or U4774 (N_4774,In_1695,In_940);
nand U4775 (N_4775,In_2422,In_1926);
or U4776 (N_4776,In_522,In_1622);
xor U4777 (N_4777,In_2193,In_660);
xnor U4778 (N_4778,In_2206,In_1977);
nor U4779 (N_4779,In_1599,In_541);
or U4780 (N_4780,In_1580,In_1980);
xor U4781 (N_4781,In_2452,In_58);
or U4782 (N_4782,In_2302,In_520);
or U4783 (N_4783,In_2784,In_844);
or U4784 (N_4784,In_2197,In_2408);
nor U4785 (N_4785,In_1065,In_1615);
xor U4786 (N_4786,In_486,In_2047);
nand U4787 (N_4787,In_378,In_31);
or U4788 (N_4788,In_641,In_2540);
nand U4789 (N_4789,In_697,In_1039);
nor U4790 (N_4790,In_204,In_1436);
nor U4791 (N_4791,In_2016,In_2946);
nor U4792 (N_4792,In_2688,In_2214);
nand U4793 (N_4793,In_2609,In_1762);
xor U4794 (N_4794,In_2511,In_1513);
nand U4795 (N_4795,In_619,In_1741);
xor U4796 (N_4796,In_912,In_1868);
nor U4797 (N_4797,In_285,In_154);
nor U4798 (N_4798,In_268,In_2712);
nor U4799 (N_4799,In_1724,In_865);
xnor U4800 (N_4800,In_737,In_2839);
and U4801 (N_4801,In_2561,In_1035);
nand U4802 (N_4802,In_2548,In_1444);
or U4803 (N_4803,In_2687,In_286);
or U4804 (N_4804,In_2215,In_766);
nand U4805 (N_4805,In_2860,In_2349);
nor U4806 (N_4806,In_1511,In_1898);
nor U4807 (N_4807,In_2208,In_2130);
and U4808 (N_4808,In_2344,In_2415);
and U4809 (N_4809,In_2221,In_670);
nor U4810 (N_4810,In_2344,In_36);
or U4811 (N_4811,In_631,In_1788);
nor U4812 (N_4812,In_1252,In_1775);
or U4813 (N_4813,In_1338,In_2030);
nor U4814 (N_4814,In_1778,In_1586);
and U4815 (N_4815,In_2597,In_336);
nor U4816 (N_4816,In_328,In_2139);
or U4817 (N_4817,In_2581,In_336);
or U4818 (N_4818,In_1867,In_1580);
or U4819 (N_4819,In_2968,In_1908);
or U4820 (N_4820,In_2845,In_2851);
or U4821 (N_4821,In_57,In_2341);
nor U4822 (N_4822,In_1218,In_922);
or U4823 (N_4823,In_303,In_418);
nand U4824 (N_4824,In_2228,In_1821);
nor U4825 (N_4825,In_2702,In_2174);
nand U4826 (N_4826,In_668,In_2842);
or U4827 (N_4827,In_726,In_2947);
and U4828 (N_4828,In_2362,In_207);
nor U4829 (N_4829,In_2368,In_2706);
xnor U4830 (N_4830,In_2969,In_1372);
and U4831 (N_4831,In_1949,In_676);
nor U4832 (N_4832,In_2266,In_1706);
or U4833 (N_4833,In_2801,In_882);
and U4834 (N_4834,In_600,In_2200);
xnor U4835 (N_4835,In_344,In_2408);
and U4836 (N_4836,In_1524,In_2817);
and U4837 (N_4837,In_2823,In_2793);
nand U4838 (N_4838,In_1027,In_1877);
xnor U4839 (N_4839,In_2815,In_1538);
nor U4840 (N_4840,In_1880,In_2788);
nand U4841 (N_4841,In_1797,In_783);
xor U4842 (N_4842,In_158,In_2879);
or U4843 (N_4843,In_1900,In_2251);
and U4844 (N_4844,In_2440,In_219);
or U4845 (N_4845,In_2043,In_1247);
or U4846 (N_4846,In_516,In_1168);
or U4847 (N_4847,In_814,In_2916);
and U4848 (N_4848,In_1120,In_748);
nor U4849 (N_4849,In_1054,In_444);
xor U4850 (N_4850,In_1685,In_414);
or U4851 (N_4851,In_1900,In_1646);
nor U4852 (N_4852,In_2774,In_958);
nor U4853 (N_4853,In_1187,In_1660);
nand U4854 (N_4854,In_179,In_1368);
nor U4855 (N_4855,In_915,In_2126);
nor U4856 (N_4856,In_2800,In_2500);
or U4857 (N_4857,In_1247,In_1912);
or U4858 (N_4858,In_2660,In_1814);
nand U4859 (N_4859,In_370,In_2364);
xnor U4860 (N_4860,In_2200,In_2510);
or U4861 (N_4861,In_933,In_1351);
and U4862 (N_4862,In_295,In_1537);
nand U4863 (N_4863,In_2813,In_1419);
or U4864 (N_4864,In_771,In_449);
nand U4865 (N_4865,In_870,In_1088);
nor U4866 (N_4866,In_1022,In_1597);
nor U4867 (N_4867,In_1294,In_2720);
nand U4868 (N_4868,In_1039,In_2716);
and U4869 (N_4869,In_40,In_2165);
nand U4870 (N_4870,In_1170,In_570);
nor U4871 (N_4871,In_461,In_1097);
nor U4872 (N_4872,In_1812,In_2770);
or U4873 (N_4873,In_1082,In_2493);
nor U4874 (N_4874,In_2706,In_686);
and U4875 (N_4875,In_2369,In_2375);
or U4876 (N_4876,In_1333,In_976);
or U4877 (N_4877,In_1605,In_1095);
and U4878 (N_4878,In_2746,In_2598);
nand U4879 (N_4879,In_1861,In_465);
nand U4880 (N_4880,In_29,In_2058);
nand U4881 (N_4881,In_1864,In_1869);
nand U4882 (N_4882,In_1306,In_1133);
or U4883 (N_4883,In_589,In_632);
xor U4884 (N_4884,In_2480,In_2581);
nand U4885 (N_4885,In_2511,In_1607);
and U4886 (N_4886,In_2639,In_2838);
and U4887 (N_4887,In_1450,In_337);
nand U4888 (N_4888,In_2911,In_2758);
nand U4889 (N_4889,In_2734,In_792);
nand U4890 (N_4890,In_127,In_882);
and U4891 (N_4891,In_1088,In_189);
or U4892 (N_4892,In_2233,In_621);
nand U4893 (N_4893,In_2195,In_1536);
nor U4894 (N_4894,In_568,In_404);
xor U4895 (N_4895,In_77,In_427);
nor U4896 (N_4896,In_2779,In_2127);
nand U4897 (N_4897,In_418,In_2892);
or U4898 (N_4898,In_139,In_2036);
nor U4899 (N_4899,In_1744,In_800);
xnor U4900 (N_4900,In_2331,In_2600);
nand U4901 (N_4901,In_1464,In_1574);
or U4902 (N_4902,In_993,In_692);
or U4903 (N_4903,In_1536,In_350);
nand U4904 (N_4904,In_1224,In_678);
and U4905 (N_4905,In_32,In_1657);
nand U4906 (N_4906,In_1060,In_2106);
or U4907 (N_4907,In_1731,In_1866);
nor U4908 (N_4908,In_810,In_1948);
nor U4909 (N_4909,In_1045,In_2225);
or U4910 (N_4910,In_134,In_5);
nor U4911 (N_4911,In_2902,In_2623);
or U4912 (N_4912,In_2134,In_2782);
xnor U4913 (N_4913,In_264,In_2341);
nand U4914 (N_4914,In_2793,In_1994);
and U4915 (N_4915,In_1211,In_887);
and U4916 (N_4916,In_790,In_101);
nand U4917 (N_4917,In_2480,In_1716);
nor U4918 (N_4918,In_2610,In_888);
and U4919 (N_4919,In_2281,In_1562);
nor U4920 (N_4920,In_2025,In_230);
xnor U4921 (N_4921,In_2821,In_854);
and U4922 (N_4922,In_2715,In_89);
nor U4923 (N_4923,In_1394,In_2928);
or U4924 (N_4924,In_2496,In_1057);
nor U4925 (N_4925,In_2559,In_801);
nand U4926 (N_4926,In_2618,In_2867);
or U4927 (N_4927,In_2493,In_447);
or U4928 (N_4928,In_1892,In_1365);
or U4929 (N_4929,In_1612,In_1611);
and U4930 (N_4930,In_1779,In_1253);
nor U4931 (N_4931,In_1783,In_637);
xnor U4932 (N_4932,In_613,In_2158);
and U4933 (N_4933,In_2424,In_1429);
or U4934 (N_4934,In_49,In_2880);
nor U4935 (N_4935,In_2636,In_195);
nor U4936 (N_4936,In_2336,In_1528);
nand U4937 (N_4937,In_960,In_1212);
or U4938 (N_4938,In_2684,In_1097);
nor U4939 (N_4939,In_1280,In_2038);
nor U4940 (N_4940,In_1633,In_742);
nand U4941 (N_4941,In_721,In_2178);
or U4942 (N_4942,In_952,In_613);
xnor U4943 (N_4943,In_316,In_2101);
xnor U4944 (N_4944,In_340,In_319);
nor U4945 (N_4945,In_2280,In_727);
or U4946 (N_4946,In_2572,In_2593);
or U4947 (N_4947,In_2112,In_2933);
nand U4948 (N_4948,In_1526,In_2472);
nand U4949 (N_4949,In_80,In_2403);
nand U4950 (N_4950,In_2793,In_1569);
nand U4951 (N_4951,In_1102,In_646);
or U4952 (N_4952,In_306,In_1222);
nor U4953 (N_4953,In_478,In_391);
or U4954 (N_4954,In_2874,In_481);
nor U4955 (N_4955,In_1058,In_346);
and U4956 (N_4956,In_1964,In_1882);
nor U4957 (N_4957,In_287,In_1248);
nand U4958 (N_4958,In_474,In_1855);
nand U4959 (N_4959,In_1358,In_2575);
and U4960 (N_4960,In_80,In_75);
or U4961 (N_4961,In_1281,In_463);
nand U4962 (N_4962,In_1649,In_2014);
or U4963 (N_4963,In_550,In_489);
nor U4964 (N_4964,In_290,In_1627);
nand U4965 (N_4965,In_561,In_1762);
nor U4966 (N_4966,In_1085,In_60);
and U4967 (N_4967,In_1827,In_90);
nor U4968 (N_4968,In_224,In_1999);
or U4969 (N_4969,In_72,In_2804);
nor U4970 (N_4970,In_140,In_2937);
or U4971 (N_4971,In_1683,In_1574);
and U4972 (N_4972,In_2288,In_5);
nand U4973 (N_4973,In_254,In_1210);
nor U4974 (N_4974,In_376,In_2589);
nor U4975 (N_4975,In_1813,In_2822);
nor U4976 (N_4976,In_1338,In_130);
nor U4977 (N_4977,In_2919,In_719);
nand U4978 (N_4978,In_2644,In_1861);
nand U4979 (N_4979,In_817,In_1788);
nand U4980 (N_4980,In_1682,In_2367);
nand U4981 (N_4981,In_140,In_1458);
nand U4982 (N_4982,In_1608,In_710);
nand U4983 (N_4983,In_869,In_1382);
nand U4984 (N_4984,In_779,In_1852);
nor U4985 (N_4985,In_1353,In_928);
xnor U4986 (N_4986,In_2194,In_597);
or U4987 (N_4987,In_1778,In_757);
or U4988 (N_4988,In_637,In_1409);
and U4989 (N_4989,In_1539,In_2643);
and U4990 (N_4990,In_2337,In_2046);
nor U4991 (N_4991,In_600,In_1871);
xnor U4992 (N_4992,In_72,In_2182);
and U4993 (N_4993,In_196,In_2763);
nand U4994 (N_4994,In_1878,In_2658);
and U4995 (N_4995,In_2064,In_2580);
nand U4996 (N_4996,In_1933,In_77);
nand U4997 (N_4997,In_2053,In_2614);
nand U4998 (N_4998,In_2649,In_2942);
nand U4999 (N_4999,In_352,In_1488);
nor U5000 (N_5000,N_313,N_1804);
nor U5001 (N_5001,N_1734,N_3616);
or U5002 (N_5002,N_4810,N_4434);
nand U5003 (N_5003,N_1886,N_253);
nand U5004 (N_5004,N_1395,N_11);
nand U5005 (N_5005,N_4887,N_1276);
and U5006 (N_5006,N_849,N_3934);
nor U5007 (N_5007,N_2027,N_1347);
or U5008 (N_5008,N_4501,N_490);
or U5009 (N_5009,N_4042,N_4975);
and U5010 (N_5010,N_2899,N_3343);
and U5011 (N_5011,N_3831,N_3344);
or U5012 (N_5012,N_63,N_121);
nor U5013 (N_5013,N_3681,N_2057);
and U5014 (N_5014,N_4385,N_2787);
nor U5015 (N_5015,N_4354,N_70);
nand U5016 (N_5016,N_1805,N_1718);
and U5017 (N_5017,N_3846,N_378);
or U5018 (N_5018,N_1437,N_3209);
nor U5019 (N_5019,N_693,N_3745);
nor U5020 (N_5020,N_977,N_827);
or U5021 (N_5021,N_577,N_4784);
and U5022 (N_5022,N_4232,N_724);
nand U5023 (N_5023,N_2611,N_3392);
and U5024 (N_5024,N_2644,N_2880);
or U5025 (N_5025,N_896,N_613);
nand U5026 (N_5026,N_1569,N_3419);
nand U5027 (N_5027,N_4352,N_3446);
xnor U5028 (N_5028,N_3526,N_3986);
and U5029 (N_5029,N_4814,N_4266);
or U5030 (N_5030,N_4590,N_1965);
xnor U5031 (N_5031,N_1962,N_830);
or U5032 (N_5032,N_2193,N_4224);
nand U5033 (N_5033,N_4956,N_1611);
xnor U5034 (N_5034,N_4473,N_4688);
or U5035 (N_5035,N_2491,N_3900);
xor U5036 (N_5036,N_3769,N_910);
nand U5037 (N_5037,N_4998,N_1217);
nor U5038 (N_5038,N_2390,N_4250);
nand U5039 (N_5039,N_3161,N_2044);
xor U5040 (N_5040,N_307,N_1911);
or U5041 (N_5041,N_4018,N_846);
nor U5042 (N_5042,N_2817,N_1952);
and U5043 (N_5043,N_4973,N_3386);
nand U5044 (N_5044,N_3198,N_1359);
nor U5045 (N_5045,N_2726,N_4374);
or U5046 (N_5046,N_2933,N_3000);
xor U5047 (N_5047,N_4336,N_3875);
and U5048 (N_5048,N_609,N_1213);
xor U5049 (N_5049,N_4401,N_1361);
nand U5050 (N_5050,N_3612,N_4782);
or U5051 (N_5051,N_3087,N_236);
and U5052 (N_5052,N_248,N_447);
or U5053 (N_5053,N_4111,N_2495);
nand U5054 (N_5054,N_170,N_9);
or U5055 (N_5055,N_4309,N_4669);
nand U5056 (N_5056,N_1788,N_46);
and U5057 (N_5057,N_344,N_3157);
or U5058 (N_5058,N_3369,N_4117);
nor U5059 (N_5059,N_2586,N_1625);
nand U5060 (N_5060,N_4282,N_1023);
or U5061 (N_5061,N_2357,N_4320);
and U5062 (N_5062,N_274,N_1507);
nand U5063 (N_5063,N_1021,N_3840);
nand U5064 (N_5064,N_2159,N_4755);
nor U5065 (N_5065,N_1224,N_3762);
xnor U5066 (N_5066,N_4217,N_989);
or U5067 (N_5067,N_2781,N_841);
nand U5068 (N_5068,N_4758,N_1552);
nand U5069 (N_5069,N_2831,N_2975);
or U5070 (N_5070,N_1615,N_2146);
or U5071 (N_5071,N_800,N_303);
or U5072 (N_5072,N_2411,N_1461);
nand U5073 (N_5073,N_2095,N_2062);
nor U5074 (N_5074,N_1424,N_1046);
and U5075 (N_5075,N_4721,N_3431);
and U5076 (N_5076,N_2373,N_297);
or U5077 (N_5077,N_231,N_635);
nand U5078 (N_5078,N_1303,N_2459);
nand U5079 (N_5079,N_1606,N_4799);
nor U5080 (N_5080,N_2779,N_587);
xor U5081 (N_5081,N_3667,N_938);
or U5082 (N_5082,N_3210,N_2805);
or U5083 (N_5083,N_942,N_3034);
nor U5084 (N_5084,N_3852,N_527);
nor U5085 (N_5085,N_4351,N_4378);
or U5086 (N_5086,N_402,N_990);
and U5087 (N_5087,N_3258,N_4933);
nor U5088 (N_5088,N_2409,N_3314);
nor U5089 (N_5089,N_2101,N_2456);
nor U5090 (N_5090,N_1139,N_1057);
nor U5091 (N_5091,N_744,N_2296);
nand U5092 (N_5092,N_1402,N_3976);
and U5093 (N_5093,N_405,N_2500);
nor U5094 (N_5094,N_4740,N_741);
or U5095 (N_5095,N_4813,N_222);
and U5096 (N_5096,N_756,N_3341);
nor U5097 (N_5097,N_1555,N_105);
or U5098 (N_5098,N_3636,N_4929);
nor U5099 (N_5099,N_3893,N_3094);
or U5100 (N_5100,N_1842,N_3791);
nor U5101 (N_5101,N_1319,N_4729);
and U5102 (N_5102,N_295,N_3531);
or U5103 (N_5103,N_4444,N_1505);
and U5104 (N_5104,N_1000,N_2043);
or U5105 (N_5105,N_2842,N_3178);
nor U5106 (N_5106,N_948,N_4459);
and U5107 (N_5107,N_1933,N_2825);
xor U5108 (N_5108,N_3383,N_4928);
nand U5109 (N_5109,N_4122,N_4618);
nand U5110 (N_5110,N_450,N_3036);
nor U5111 (N_5111,N_2808,N_1257);
or U5112 (N_5112,N_862,N_970);
nand U5113 (N_5113,N_4854,N_3701);
and U5114 (N_5114,N_608,N_4511);
xor U5115 (N_5115,N_221,N_389);
xnor U5116 (N_5116,N_665,N_3371);
nor U5117 (N_5117,N_2271,N_3236);
or U5118 (N_5118,N_2153,N_3364);
and U5119 (N_5119,N_3155,N_469);
or U5120 (N_5120,N_1195,N_391);
or U5121 (N_5121,N_895,N_1206);
nor U5122 (N_5122,N_4718,N_2964);
nor U5123 (N_5123,N_1918,N_4253);
or U5124 (N_5124,N_4941,N_4964);
nor U5125 (N_5125,N_3175,N_4684);
nor U5126 (N_5126,N_212,N_4872);
and U5127 (N_5127,N_3981,N_1603);
or U5128 (N_5128,N_2157,N_3948);
nand U5129 (N_5129,N_4291,N_3412);
and U5130 (N_5130,N_3650,N_2510);
and U5131 (N_5131,N_1680,N_1586);
nor U5132 (N_5132,N_1940,N_2670);
nand U5133 (N_5133,N_3190,N_1752);
or U5134 (N_5134,N_1450,N_2548);
or U5135 (N_5135,N_336,N_1454);
and U5136 (N_5136,N_2946,N_1494);
or U5137 (N_5137,N_4347,N_3759);
nor U5138 (N_5138,N_597,N_1921);
nor U5139 (N_5139,N_1644,N_3674);
and U5140 (N_5140,N_4389,N_1444);
and U5141 (N_5141,N_1588,N_416);
or U5142 (N_5142,N_3628,N_1455);
nand U5143 (N_5143,N_4880,N_1714);
xor U5144 (N_5144,N_1553,N_2662);
or U5145 (N_5145,N_3538,N_921);
and U5146 (N_5146,N_1131,N_2818);
or U5147 (N_5147,N_4619,N_2713);
or U5148 (N_5148,N_4948,N_3851);
nand U5149 (N_5149,N_2361,N_123);
or U5150 (N_5150,N_1299,N_3376);
or U5151 (N_5151,N_2689,N_2783);
nand U5152 (N_5152,N_2681,N_4314);
or U5153 (N_5153,N_2244,N_1687);
or U5154 (N_5154,N_3377,N_652);
nand U5155 (N_5155,N_4835,N_2738);
nor U5156 (N_5156,N_4907,N_4139);
nor U5157 (N_5157,N_3891,N_1813);
or U5158 (N_5158,N_3618,N_1763);
or U5159 (N_5159,N_473,N_2520);
or U5160 (N_5160,N_1433,N_2737);
nand U5161 (N_5161,N_2201,N_3604);
nand U5162 (N_5162,N_4962,N_2503);
xnor U5163 (N_5163,N_3323,N_1639);
or U5164 (N_5164,N_2824,N_3133);
or U5165 (N_5165,N_213,N_3266);
and U5166 (N_5166,N_406,N_3630);
or U5167 (N_5167,N_1683,N_2859);
and U5168 (N_5168,N_1595,N_4938);
nand U5169 (N_5169,N_631,N_737);
and U5170 (N_5170,N_1945,N_658);
nand U5171 (N_5171,N_4337,N_622);
nor U5172 (N_5172,N_3201,N_2351);
nand U5173 (N_5173,N_2403,N_1891);
nor U5174 (N_5174,N_2154,N_1104);
nand U5175 (N_5175,N_1272,N_1121);
or U5176 (N_5176,N_195,N_760);
nor U5177 (N_5177,N_4040,N_3448);
or U5178 (N_5178,N_2544,N_135);
and U5179 (N_5179,N_2528,N_3219);
or U5180 (N_5180,N_4142,N_3045);
or U5181 (N_5181,N_3651,N_2121);
or U5182 (N_5182,N_3480,N_1358);
and U5183 (N_5183,N_1915,N_1253);
nand U5184 (N_5184,N_991,N_3284);
nand U5185 (N_5185,N_264,N_2498);
nand U5186 (N_5186,N_512,N_489);
or U5187 (N_5187,N_2698,N_1829);
xnor U5188 (N_5188,N_3283,N_4935);
and U5189 (N_5189,N_1240,N_2733);
nor U5190 (N_5190,N_2900,N_3);
nor U5191 (N_5191,N_865,N_1246);
and U5192 (N_5192,N_4919,N_754);
or U5193 (N_5193,N_3066,N_1503);
or U5194 (N_5194,N_3415,N_4882);
nor U5195 (N_5195,N_3914,N_4070);
nand U5196 (N_5196,N_1992,N_1113);
nand U5197 (N_5197,N_4708,N_2185);
or U5198 (N_5198,N_1202,N_245);
or U5199 (N_5199,N_2269,N_2002);
or U5200 (N_5200,N_3204,N_3334);
or U5201 (N_5201,N_2522,N_3351);
nor U5202 (N_5202,N_1176,N_4791);
or U5203 (N_5203,N_31,N_3430);
and U5204 (N_5204,N_695,N_4110);
xor U5205 (N_5205,N_1235,N_306);
nor U5206 (N_5206,N_2915,N_3876);
nand U5207 (N_5207,N_1579,N_2898);
and U5208 (N_5208,N_2813,N_751);
nand U5209 (N_5209,N_550,N_2284);
nor U5210 (N_5210,N_3718,N_2213);
and U5211 (N_5211,N_4976,N_4769);
or U5212 (N_5212,N_1037,N_2716);
and U5213 (N_5213,N_4229,N_4779);
nor U5214 (N_5214,N_1968,N_3613);
and U5215 (N_5215,N_833,N_4234);
nand U5216 (N_5216,N_4360,N_1501);
or U5217 (N_5217,N_1912,N_4596);
nand U5218 (N_5218,N_1153,N_3324);
or U5219 (N_5219,N_1493,N_1719);
and U5220 (N_5220,N_1695,N_3911);
nor U5221 (N_5221,N_552,N_848);
and U5222 (N_5222,N_2655,N_3179);
and U5223 (N_5223,N_965,N_2616);
nor U5224 (N_5224,N_3693,N_4044);
nor U5225 (N_5225,N_4055,N_2582);
nor U5226 (N_5226,N_1955,N_2345);
xor U5227 (N_5227,N_64,N_2);
nand U5228 (N_5228,N_4920,N_777);
or U5229 (N_5229,N_2490,N_706);
or U5230 (N_5230,N_1720,N_4299);
or U5231 (N_5231,N_3043,N_1273);
nand U5232 (N_5232,N_3584,N_917);
nand U5233 (N_5233,N_423,N_171);
nor U5234 (N_5234,N_4700,N_3873);
nand U5235 (N_5235,N_1990,N_4436);
and U5236 (N_5236,N_3465,N_3352);
nand U5237 (N_5237,N_3231,N_215);
nand U5238 (N_5238,N_3261,N_2626);
nor U5239 (N_5239,N_2906,N_2417);
nor U5240 (N_5240,N_191,N_4133);
nand U5241 (N_5241,N_2207,N_2181);
or U5242 (N_5242,N_1214,N_409);
or U5243 (N_5243,N_529,N_4005);
and U5244 (N_5244,N_4141,N_1283);
nor U5245 (N_5245,N_2455,N_4179);
nand U5246 (N_5246,N_3990,N_3682);
or U5247 (N_5247,N_1049,N_1201);
or U5248 (N_5248,N_3505,N_3092);
nand U5249 (N_5249,N_79,N_4908);
and U5250 (N_5250,N_4999,N_3763);
and U5251 (N_5251,N_3128,N_4553);
nand U5252 (N_5252,N_82,N_1372);
or U5253 (N_5253,N_941,N_4711);
xnor U5254 (N_5254,N_1295,N_1407);
nand U5255 (N_5255,N_3235,N_971);
and U5256 (N_5256,N_2126,N_179);
nand U5257 (N_5257,N_311,N_4983);
xor U5258 (N_5258,N_369,N_4623);
or U5259 (N_5259,N_4969,N_1400);
nor U5260 (N_5260,N_201,N_2923);
or U5261 (N_5261,N_4621,N_3320);
nand U5262 (N_5262,N_4519,N_2647);
nand U5263 (N_5263,N_2748,N_3458);
or U5264 (N_5264,N_2612,N_2467);
nand U5265 (N_5265,N_1060,N_1197);
nand U5266 (N_5266,N_2341,N_3440);
nor U5267 (N_5267,N_484,N_2111);
and U5268 (N_5268,N_3040,N_2051);
or U5269 (N_5269,N_4630,N_2005);
nor U5270 (N_5270,N_4824,N_451);
nor U5271 (N_5271,N_1741,N_4426);
or U5272 (N_5272,N_766,N_4372);
and U5273 (N_5273,N_4727,N_206);
and U5274 (N_5274,N_3308,N_559);
nand U5275 (N_5275,N_668,N_2451);
or U5276 (N_5276,N_1277,N_4380);
nor U5277 (N_5277,N_700,N_870);
xnor U5278 (N_5278,N_858,N_3321);
or U5279 (N_5279,N_3031,N_1738);
xor U5280 (N_5280,N_2212,N_1421);
and U5281 (N_5281,N_58,N_1840);
nor U5282 (N_5282,N_778,N_1182);
nand U5283 (N_5283,N_3638,N_4893);
or U5284 (N_5284,N_655,N_332);
nor U5285 (N_5285,N_2888,N_1094);
nor U5286 (N_5286,N_1546,N_4079);
nand U5287 (N_5287,N_1960,N_459);
nor U5288 (N_5288,N_37,N_4716);
nand U5289 (N_5289,N_3626,N_1298);
and U5290 (N_5290,N_18,N_3938);
nand U5291 (N_5291,N_3683,N_4656);
nor U5292 (N_5292,N_2067,N_2601);
and U5293 (N_5293,N_716,N_3821);
nand U5294 (N_5294,N_3785,N_1848);
or U5295 (N_5295,N_4696,N_216);
nor U5296 (N_5296,N_1472,N_3265);
nand U5297 (N_5297,N_1868,N_2200);
nor U5298 (N_5298,N_4858,N_1244);
nand U5299 (N_5299,N_547,N_208);
xnor U5300 (N_5300,N_1492,N_1950);
nor U5301 (N_5301,N_3275,N_2585);
nand U5302 (N_5302,N_3025,N_1963);
nor U5303 (N_5303,N_1793,N_4734);
nand U5304 (N_5304,N_1999,N_4068);
and U5305 (N_5305,N_1574,N_379);
nand U5306 (N_5306,N_946,N_4206);
nand U5307 (N_5307,N_2856,N_1670);
nand U5308 (N_5308,N_4588,N_2176);
or U5309 (N_5309,N_3479,N_435);
and U5310 (N_5310,N_612,N_1498);
nand U5311 (N_5311,N_1536,N_4506);
xor U5312 (N_5312,N_663,N_1301);
nor U5313 (N_5313,N_540,N_4617);
nor U5314 (N_5314,N_1123,N_1535);
xor U5315 (N_5315,N_4633,N_2381);
nor U5316 (N_5316,N_4805,N_793);
or U5317 (N_5317,N_2120,N_3437);
and U5318 (N_5318,N_1203,N_4248);
nor U5319 (N_5319,N_536,N_1701);
xnor U5320 (N_5320,N_4572,N_1550);
nor U5321 (N_5321,N_4402,N_4322);
and U5322 (N_5322,N_3606,N_3012);
and U5323 (N_5323,N_1497,N_1027);
and U5324 (N_5324,N_2668,N_3809);
and U5325 (N_5325,N_229,N_1653);
nor U5326 (N_5326,N_3060,N_3228);
nor U5327 (N_5327,N_4147,N_2930);
nand U5328 (N_5328,N_4335,N_4802);
nand U5329 (N_5329,N_4756,N_2047);
or U5330 (N_5330,N_316,N_3143);
and U5331 (N_5331,N_497,N_258);
and U5332 (N_5332,N_319,N_2097);
or U5333 (N_5333,N_3238,N_4143);
nand U5334 (N_5334,N_1510,N_1102);
nand U5335 (N_5335,N_732,N_439);
nor U5336 (N_5336,N_3950,N_2919);
or U5337 (N_5337,N_3889,N_2545);
nand U5338 (N_5338,N_4667,N_2460);
xnor U5339 (N_5339,N_1907,N_538);
or U5340 (N_5340,N_36,N_4176);
or U5341 (N_5341,N_3273,N_2191);
or U5342 (N_5342,N_1927,N_4660);
nand U5343 (N_5343,N_3356,N_3885);
or U5344 (N_5344,N_4049,N_2519);
or U5345 (N_5345,N_3473,N_2718);
nand U5346 (N_5346,N_2725,N_725);
and U5347 (N_5347,N_4647,N_2897);
nand U5348 (N_5348,N_1864,N_2010);
and U5349 (N_5349,N_2109,N_2569);
nor U5350 (N_5350,N_2116,N_2504);
or U5351 (N_5351,N_3573,N_2727);
nand U5352 (N_5352,N_2627,N_752);
nand U5353 (N_5353,N_3892,N_3050);
nor U5354 (N_5354,N_3887,N_2326);
or U5355 (N_5355,N_3342,N_2033);
or U5356 (N_5356,N_1570,N_610);
or U5357 (N_5357,N_4287,N_1392);
and U5358 (N_5358,N_4991,N_2717);
and U5359 (N_5359,N_34,N_3138);
nor U5360 (N_5360,N_1879,N_1414);
and U5361 (N_5361,N_3183,N_1533);
and U5362 (N_5362,N_4869,N_2087);
and U5363 (N_5363,N_2571,N_47);
or U5364 (N_5364,N_768,N_2458);
and U5365 (N_5365,N_496,N_3168);
and U5366 (N_5366,N_243,N_3089);
nor U5367 (N_5367,N_3117,N_4532);
xnor U5368 (N_5368,N_4350,N_4736);
or U5369 (N_5369,N_2184,N_3869);
nor U5370 (N_5370,N_1596,N_797);
nand U5371 (N_5371,N_4267,N_4943);
or U5372 (N_5372,N_2079,N_1418);
nor U5373 (N_5373,N_1045,N_1167);
or U5374 (N_5374,N_653,N_1818);
nor U5375 (N_5375,N_1883,N_1621);
nand U5376 (N_5376,N_3227,N_2436);
or U5377 (N_5377,N_1396,N_3129);
xor U5378 (N_5378,N_685,N_1173);
nor U5379 (N_5379,N_1685,N_2376);
xor U5380 (N_5380,N_4086,N_1649);
nand U5381 (N_5381,N_23,N_183);
or U5382 (N_5382,N_3224,N_2881);
nand U5383 (N_5383,N_3753,N_2579);
xnor U5384 (N_5384,N_66,N_28);
nor U5385 (N_5385,N_4911,N_2792);
nor U5386 (N_5386,N_2526,N_3353);
and U5387 (N_5387,N_2093,N_1026);
nor U5388 (N_5388,N_1591,N_4742);
xnor U5389 (N_5389,N_2938,N_2695);
nand U5390 (N_5390,N_955,N_2209);
and U5391 (N_5391,N_3735,N_4323);
nor U5392 (N_5392,N_1162,N_4095);
nor U5393 (N_5393,N_1810,N_4388);
and U5394 (N_5394,N_1177,N_2761);
nor U5395 (N_5395,N_4724,N_3080);
nand U5396 (N_5396,N_629,N_4741);
nor U5397 (N_5397,N_1245,N_4892);
xor U5398 (N_5398,N_1654,N_2066);
or U5399 (N_5399,N_4978,N_73);
nand U5400 (N_5400,N_3196,N_3101);
nand U5401 (N_5401,N_4862,N_2833);
xor U5402 (N_5402,N_4628,N_2648);
and U5403 (N_5403,N_692,N_2337);
and U5404 (N_5404,N_2192,N_4842);
and U5405 (N_5405,N_603,N_4289);
or U5406 (N_5406,N_3244,N_543);
and U5407 (N_5407,N_323,N_493);
and U5408 (N_5408,N_1149,N_1093);
nand U5409 (N_5409,N_3528,N_2583);
nand U5410 (N_5410,N_2420,N_4706);
nor U5411 (N_5411,N_234,N_3591);
and U5412 (N_5412,N_2550,N_3064);
or U5413 (N_5413,N_202,N_4302);
and U5414 (N_5414,N_3492,N_1811);
nor U5415 (N_5415,N_1529,N_2145);
and U5416 (N_5416,N_4989,N_2036);
or U5417 (N_5417,N_3629,N_3478);
or U5418 (N_5418,N_1011,N_3367);
nand U5419 (N_5419,N_4828,N_3609);
nor U5420 (N_5420,N_2966,N_4985);
and U5421 (N_5421,N_4029,N_4857);
nand U5422 (N_5422,N_736,N_2298);
or U5423 (N_5423,N_4405,N_4598);
nand U5424 (N_5424,N_4204,N_4896);
and U5425 (N_5425,N_4123,N_511);
nor U5426 (N_5426,N_4771,N_2018);
or U5427 (N_5427,N_3061,N_824);
xor U5428 (N_5428,N_2000,N_1511);
and U5429 (N_5429,N_1315,N_108);
or U5430 (N_5430,N_1003,N_2396);
nor U5431 (N_5431,N_625,N_968);
nand U5432 (N_5432,N_886,N_4889);
and U5433 (N_5433,N_2714,N_3096);
nand U5434 (N_5434,N_4987,N_3277);
and U5435 (N_5435,N_1619,N_238);
nor U5436 (N_5436,N_3535,N_1264);
and U5437 (N_5437,N_2492,N_3520);
nor U5438 (N_5438,N_2853,N_1029);
nor U5439 (N_5439,N_2139,N_1089);
and U5440 (N_5440,N_1211,N_1078);
nand U5441 (N_5441,N_277,N_136);
or U5442 (N_5442,N_906,N_1025);
nor U5443 (N_5443,N_4730,N_1067);
and U5444 (N_5444,N_3725,N_249);
and U5445 (N_5445,N_4750,N_3729);
or U5446 (N_5446,N_709,N_4376);
and U5447 (N_5447,N_1913,N_1863);
nand U5448 (N_5448,N_4502,N_891);
xnor U5449 (N_5449,N_1766,N_2630);
xnor U5450 (N_5450,N_3347,N_1185);
or U5451 (N_5451,N_3588,N_3029);
nor U5452 (N_5452,N_3713,N_2052);
nand U5453 (N_5453,N_2908,N_677);
or U5454 (N_5454,N_8,N_2677);
nand U5455 (N_5455,N_1977,N_2001);
nor U5456 (N_5456,N_1629,N_301);
nor U5457 (N_5457,N_3062,N_1608);
nand U5458 (N_5458,N_275,N_32);
or U5459 (N_5459,N_4279,N_4344);
and U5460 (N_5460,N_1753,N_3105);
nand U5461 (N_5461,N_755,N_349);
nor U5462 (N_5462,N_448,N_241);
and U5463 (N_5463,N_4797,N_3744);
nor U5464 (N_5464,N_4059,N_342);
or U5465 (N_5465,N_3985,N_338);
and U5466 (N_5466,N_2775,N_4109);
nand U5467 (N_5467,N_257,N_1378);
and U5468 (N_5468,N_4608,N_1145);
xnor U5469 (N_5469,N_632,N_1739);
nand U5470 (N_5470,N_2650,N_844);
nor U5471 (N_5471,N_3030,N_2961);
nand U5472 (N_5472,N_1432,N_4512);
or U5473 (N_5473,N_805,N_2928);
or U5474 (N_5474,N_50,N_591);
or U5475 (N_5475,N_1226,N_3907);
and U5476 (N_5476,N_1765,N_4474);
or U5477 (N_5477,N_1083,N_1607);
nand U5478 (N_5478,N_4582,N_4903);
or U5479 (N_5479,N_3634,N_3818);
and U5480 (N_5480,N_3391,N_590);
and U5481 (N_5481,N_3263,N_2252);
nor U5482 (N_5482,N_592,N_314);
nor U5483 (N_5483,N_4475,N_2890);
nand U5484 (N_5484,N_3903,N_4697);
nor U5485 (N_5485,N_1946,N_4230);
or U5486 (N_5486,N_879,N_2424);
or U5487 (N_5487,N_623,N_4007);
and U5488 (N_5488,N_4577,N_2871);
nor U5489 (N_5489,N_2136,N_3269);
nand U5490 (N_5490,N_4952,N_4045);
or U5491 (N_5491,N_2049,N_4632);
nand U5492 (N_5492,N_1541,N_2663);
nor U5493 (N_5493,N_2724,N_2442);
and U5494 (N_5494,N_641,N_2473);
nand U5495 (N_5495,N_1613,N_2158);
and U5496 (N_5496,N_1682,N_589);
nand U5497 (N_5497,N_3009,N_1008);
xnor U5498 (N_5498,N_4800,N_1098);
nor U5499 (N_5499,N_244,N_2584);
nand U5500 (N_5500,N_1478,N_1849);
or U5501 (N_5501,N_1759,N_4167);
and U5502 (N_5502,N_1034,N_638);
or U5503 (N_5503,N_318,N_292);
and U5504 (N_5504,N_44,N_4054);
and U5505 (N_5505,N_1696,N_3992);
or U5506 (N_5506,N_3624,N_4789);
and U5507 (N_5507,N_4020,N_382);
nor U5508 (N_5508,N_4427,N_3393);
nand U5509 (N_5509,N_2661,N_4550);
nor U5510 (N_5510,N_4208,N_2563);
and U5511 (N_5511,N_2774,N_3287);
nand U5512 (N_5512,N_3281,N_194);
nor U5513 (N_5513,N_516,N_3648);
nor U5514 (N_5514,N_4316,N_4362);
or U5515 (N_5515,N_77,N_2387);
nand U5516 (N_5516,N_1733,N_783);
xor U5517 (N_5517,N_4855,N_675);
and U5518 (N_5518,N_818,N_1697);
or U5519 (N_5519,N_674,N_3004);
xor U5520 (N_5520,N_3229,N_823);
xor U5521 (N_5521,N_2554,N_3988);
and U5522 (N_5522,N_109,N_345);
or U5523 (N_5523,N_2314,N_530);
nor U5524 (N_5524,N_2007,N_2107);
nor U5525 (N_5525,N_293,N_2084);
or U5526 (N_5526,N_1627,N_4877);
or U5527 (N_5527,N_4571,N_15);
and U5528 (N_5528,N_2452,N_4682);
or U5529 (N_5529,N_4787,N_723);
or U5530 (N_5530,N_2266,N_1188);
and U5531 (N_5531,N_4184,N_4996);
xnor U5532 (N_5532,N_934,N_3047);
nand U5533 (N_5533,N_2719,N_1548);
and U5534 (N_5534,N_3983,N_1275);
nand U5535 (N_5535,N_139,N_3163);
nor U5536 (N_5536,N_4333,N_3326);
nor U5537 (N_5537,N_4548,N_1561);
nor U5538 (N_5538,N_645,N_3814);
nand U5539 (N_5539,N_2312,N_1242);
nand U5540 (N_5540,N_2304,N_634);
nand U5541 (N_5541,N_1125,N_2895);
or U5542 (N_5542,N_267,N_93);
or U5543 (N_5543,N_1311,N_3305);
and U5544 (N_5544,N_2308,N_650);
nor U5545 (N_5545,N_2872,N_3390);
nor U5546 (N_5546,N_2349,N_3216);
or U5547 (N_5547,N_1906,N_3511);
nor U5548 (N_5548,N_585,N_1512);
or U5549 (N_5549,N_1473,N_2777);
nor U5550 (N_5550,N_1019,N_2592);
and U5551 (N_5551,N_1479,N_4757);
nor U5552 (N_5552,N_2023,N_2083);
nor U5553 (N_5553,N_4085,N_4524);
nor U5554 (N_5554,N_4406,N_2362);
xnor U5555 (N_5555,N_365,N_3790);
nand U5556 (N_5556,N_3810,N_4479);
xnor U5557 (N_5557,N_4754,N_498);
xnor U5558 (N_5558,N_256,N_425);
nor U5559 (N_5559,N_3699,N_3056);
and U5560 (N_5560,N_2489,N_3394);
and U5561 (N_5561,N_408,N_4125);
or U5562 (N_5562,N_2753,N_2851);
xnor U5563 (N_5563,N_3741,N_803);
and U5564 (N_5564,N_2279,N_837);
nor U5565 (N_5565,N_918,N_501);
nand U5566 (N_5566,N_856,N_4022);
nand U5567 (N_5567,N_1799,N_145);
nor U5568 (N_5568,N_3730,N_3687);
or U5569 (N_5569,N_3502,N_4240);
or U5570 (N_5570,N_4024,N_3280);
and U5571 (N_5571,N_2178,N_1334);
nand U5572 (N_5572,N_2280,N_2924);
nor U5573 (N_5573,N_4820,N_651);
nor U5574 (N_5574,N_494,N_1484);
and U5575 (N_5575,N_3566,N_4542);
nor U5576 (N_5576,N_3951,N_4574);
or U5577 (N_5577,N_1142,N_3118);
nand U5578 (N_5578,N_4284,N_664);
and U5579 (N_5579,N_1964,N_952);
or U5580 (N_5580,N_2956,N_2998);
and U5581 (N_5581,N_4442,N_2081);
nor U5582 (N_5582,N_2977,N_3671);
and U5583 (N_5583,N_4078,N_1379);
or U5584 (N_5584,N_2202,N_761);
or U5585 (N_5585,N_3468,N_3781);
or U5586 (N_5586,N_471,N_3749);
xor U5587 (N_5587,N_3643,N_3349);
nor U5588 (N_5588,N_4915,N_368);
nand U5589 (N_5589,N_966,N_1779);
and U5590 (N_5590,N_3476,N_3614);
nor U5591 (N_5591,N_4804,N_3700);
nand U5592 (N_5592,N_1134,N_2470);
xor U5593 (N_5593,N_2437,N_1168);
or U5594 (N_5594,N_506,N_4249);
nand U5595 (N_5595,N_4261,N_4177);
nand U5596 (N_5596,N_3136,N_681);
nor U5597 (N_5597,N_1795,N_4056);
nand U5598 (N_5598,N_5,N_1594);
and U5599 (N_5599,N_774,N_1363);
nand U5600 (N_5600,N_4946,N_2514);
or U5601 (N_5601,N_2782,N_449);
nand U5602 (N_5602,N_4692,N_3569);
or U5603 (N_5603,N_4001,N_2760);
nor U5604 (N_5604,N_4870,N_2183);
nor U5605 (N_5605,N_3568,N_1580);
and U5606 (N_5606,N_888,N_1356);
nor U5607 (N_5607,N_2840,N_4178);
and U5608 (N_5608,N_940,N_1282);
or U5609 (N_5609,N_4589,N_3708);
nor U5610 (N_5610,N_2377,N_4439);
and U5611 (N_5611,N_2543,N_3193);
or U5612 (N_5612,N_2652,N_4516);
nand U5613 (N_5613,N_639,N_1525);
and U5614 (N_5614,N_4080,N_1647);
nand U5615 (N_5615,N_3474,N_4643);
nand U5616 (N_5616,N_3270,N_164);
and U5617 (N_5617,N_3169,N_1411);
or U5618 (N_5618,N_3125,N_4627);
or U5619 (N_5619,N_4859,N_3093);
nand U5620 (N_5620,N_98,N_572);
or U5621 (N_5621,N_3329,N_2040);
or U5622 (N_5622,N_2289,N_721);
xor U5623 (N_5623,N_2285,N_1828);
xnor U5624 (N_5624,N_2640,N_654);
and U5625 (N_5625,N_4830,N_455);
and U5626 (N_5626,N_1169,N_3217);
and U5627 (N_5627,N_2844,N_399);
and U5628 (N_5628,N_2415,N_3655);
nand U5629 (N_5629,N_3654,N_3822);
and U5630 (N_5630,N_546,N_738);
xnor U5631 (N_5631,N_2599,N_3888);
and U5632 (N_5632,N_2884,N_2048);
or U5633 (N_5633,N_1269,N_4012);
or U5634 (N_5634,N_2931,N_4605);
nor U5635 (N_5635,N_671,N_210);
nand U5636 (N_5636,N_1831,N_920);
nor U5637 (N_5637,N_1204,N_4980);
nor U5638 (N_5638,N_1809,N_1079);
nand U5639 (N_5639,N_1120,N_4203);
or U5640 (N_5640,N_3770,N_682);
nor U5641 (N_5641,N_331,N_4225);
nand U5642 (N_5642,N_2903,N_4415);
or U5643 (N_5643,N_2602,N_2963);
nor U5644 (N_5644,N_2960,N_1662);
nor U5645 (N_5645,N_436,N_4592);
nand U5646 (N_5646,N_4864,N_4437);
and U5647 (N_5647,N_4847,N_2429);
or U5648 (N_5648,N_3286,N_3119);
nor U5649 (N_5649,N_2874,N_3787);
xnor U5650 (N_5650,N_4714,N_3104);
nand U5651 (N_5651,N_2828,N_2309);
xor U5652 (N_5652,N_3510,N_2135);
nand U5653 (N_5653,N_4747,N_2021);
and U5654 (N_5654,N_2597,N_980);
and U5655 (N_5655,N_1768,N_4092);
xor U5656 (N_5656,N_3370,N_4215);
or U5657 (N_5657,N_1645,N_122);
nor U5658 (N_5658,N_1114,N_1453);
or U5659 (N_5659,N_317,N_3184);
and U5660 (N_5660,N_1538,N_4435);
nand U5661 (N_5661,N_3558,N_579);
or U5662 (N_5662,N_157,N_3855);
nor U5663 (N_5663,N_4701,N_982);
nor U5664 (N_5664,N_770,N_957);
and U5665 (N_5665,N_1254,N_1587);
nor U5666 (N_5666,N_4159,N_2982);
nand U5667 (N_5667,N_3906,N_2524);
nor U5668 (N_5668,N_3844,N_3223);
nor U5669 (N_5669,N_4382,N_254);
nand U5670 (N_5670,N_1563,N_1944);
nand U5671 (N_5671,N_743,N_604);
xnor U5672 (N_5672,N_158,N_2485);
and U5673 (N_5673,N_2720,N_3659);
nor U5674 (N_5674,N_4515,N_1745);
nor U5675 (N_5675,N_227,N_1292);
nand U5676 (N_5676,N_4957,N_3955);
nand U5677 (N_5677,N_3932,N_4293);
nor U5678 (N_5678,N_1866,N_315);
nor U5679 (N_5679,N_383,N_4982);
or U5680 (N_5680,N_16,N_2182);
nor U5681 (N_5681,N_2393,N_3524);
nor U5682 (N_5682,N_1066,N_3315);
nor U5683 (N_5683,N_2061,N_4418);
xnor U5684 (N_5684,N_4599,N_3276);
nor U5685 (N_5685,N_2955,N_962);
and U5686 (N_5686,N_4759,N_1252);
nor U5687 (N_5687,N_3515,N_266);
nor U5688 (N_5688,N_1291,N_2697);
nor U5689 (N_5689,N_4431,N_4008);
nand U5690 (N_5690,N_3707,N_1578);
or U5691 (N_5691,N_3167,N_2746);
nand U5692 (N_5692,N_4646,N_570);
xnor U5693 (N_5693,N_2168,N_821);
nand U5694 (N_5694,N_466,N_3989);
xor U5695 (N_5695,N_308,N_350);
and U5696 (N_5696,N_3147,N_53);
nand U5697 (N_5697,N_120,N_515);
and U5698 (N_5698,N_1815,N_825);
and U5699 (N_5699,N_2696,N_1539);
and U5700 (N_5700,N_84,N_1187);
nor U5701 (N_5701,N_3698,N_2481);
or U5702 (N_5702,N_1051,N_2433);
xor U5703 (N_5703,N_2106,N_1887);
and U5704 (N_5704,N_2287,N_4452);
and U5705 (N_5705,N_39,N_4698);
nor U5706 (N_5706,N_1063,N_3943);
and U5707 (N_5707,N_3107,N_4798);
or U5708 (N_5708,N_3137,N_4668);
nor U5709 (N_5709,N_2921,N_556);
nor U5710 (N_5710,N_3037,N_1726);
nand U5711 (N_5711,N_914,N_1735);
nor U5712 (N_5712,N_614,N_1038);
and U5713 (N_5713,N_595,N_1560);
nand U5714 (N_5714,N_3074,N_4745);
nor U5715 (N_5715,N_4984,N_2523);
or U5716 (N_5716,N_1502,N_2854);
and U5717 (N_5717,N_3575,N_381);
nor U5718 (N_5718,N_199,N_4171);
nor U5719 (N_5719,N_953,N_101);
nor U5720 (N_5720,N_3969,N_2624);
and U5721 (N_5721,N_2076,N_2418);
and U5722 (N_5722,N_541,N_75);
nand U5723 (N_5723,N_1221,N_2758);
nor U5724 (N_5724,N_995,N_2297);
and U5725 (N_5725,N_1600,N_3920);
or U5726 (N_5726,N_3172,N_2127);
nor U5727 (N_5727,N_3673,N_3354);
or U5728 (N_5728,N_3188,N_2598);
nand U5729 (N_5729,N_930,N_4918);
nor U5730 (N_5730,N_2555,N_3327);
nor U5731 (N_5731,N_2531,N_1822);
xor U5732 (N_5732,N_1551,N_3084);
nor U5733 (N_5733,N_1704,N_2795);
xnor U5734 (N_5734,N_1671,N_1837);
nor U5735 (N_5735,N_3754,N_3052);
xor U5736 (N_5736,N_2637,N_1661);
nor U5737 (N_5737,N_2756,N_3237);
nand U5738 (N_5738,N_4258,N_757);
or U5739 (N_5739,N_1441,N_730);
nand U5740 (N_5740,N_1881,N_396);
or U5741 (N_5741,N_1256,N_4611);
nand U5742 (N_5742,N_1890,N_4329);
nand U5743 (N_5743,N_525,N_3159);
and U5744 (N_5744,N_2468,N_2858);
nand U5745 (N_5745,N_374,N_3572);
nand U5746 (N_5746,N_1429,N_390);
and U5747 (N_5747,N_4272,N_1584);
or U5748 (N_5748,N_2987,N_2711);
xor U5749 (N_5749,N_1043,N_745);
nor U5750 (N_5750,N_3580,N_1081);
and U5751 (N_5751,N_3429,N_1711);
xnor U5752 (N_5752,N_1313,N_174);
nor U5753 (N_5753,N_3467,N_3670);
nand U5754 (N_5754,N_1486,N_4464);
or U5755 (N_5755,N_2538,N_1679);
or U5756 (N_5756,N_2386,N_3848);
and U5757 (N_5757,N_3049,N_4988);
or U5758 (N_5758,N_2743,N_2723);
nand U5759 (N_5759,N_1756,N_1033);
nand U5760 (N_5760,N_232,N_4124);
xor U5761 (N_5761,N_814,N_3368);
nand U5762 (N_5762,N_851,N_49);
nor U5763 (N_5763,N_1851,N_4432);
or U5764 (N_5764,N_2226,N_3902);
or U5765 (N_5765,N_4732,N_4233);
xor U5766 (N_5766,N_3203,N_184);
xor U5767 (N_5767,N_3635,N_4255);
or U5768 (N_5768,N_3957,N_3578);
nand U5769 (N_5769,N_4637,N_4932);
nand U5770 (N_5770,N_4888,N_2450);
nor U5771 (N_5771,N_4665,N_403);
and U5772 (N_5772,N_4321,N_4326);
or U5773 (N_5773,N_2749,N_290);
nand U5774 (N_5774,N_4462,N_2194);
and U5775 (N_5775,N_518,N_57);
nor U5776 (N_5776,N_4116,N_3847);
nand U5777 (N_5777,N_4861,N_1354);
nand U5778 (N_5778,N_4538,N_4879);
or U5779 (N_5779,N_2688,N_351);
or U5780 (N_5780,N_1702,N_2623);
or U5781 (N_5781,N_288,N_1979);
nor U5782 (N_5782,N_3069,N_628);
xor U5783 (N_5783,N_1523,N_1564);
and U5784 (N_5784,N_1018,N_1056);
nand U5785 (N_5785,N_507,N_226);
xnor U5786 (N_5786,N_4545,N_2827);
or U5787 (N_5787,N_163,N_2138);
or U5788 (N_5788,N_1419,N_2156);
nor U5789 (N_5789,N_2016,N_3271);
nor U5790 (N_5790,N_1889,N_26);
and U5791 (N_5791,N_4075,N_4901);
xor U5792 (N_5792,N_133,N_4694);
nand U5793 (N_5793,N_3783,N_1664);
nor U5794 (N_5794,N_1814,N_961);
nor U5795 (N_5795,N_1589,N_4944);
nor U5796 (N_5796,N_261,N_134);
and U5797 (N_5797,N_176,N_4648);
nand U5798 (N_5798,N_3679,N_1634);
nor U5799 (N_5799,N_840,N_242);
or U5800 (N_5800,N_1412,N_1101);
or U5801 (N_5801,N_1919,N_1308);
and U5802 (N_5802,N_4495,N_2735);
or U5803 (N_5803,N_2412,N_3523);
or U5804 (N_5804,N_3127,N_3010);
or U5805 (N_5805,N_4476,N_2745);
nor U5806 (N_5806,N_2148,N_407);
nor U5807 (N_5807,N_4968,N_2552);
xor U5808 (N_5808,N_4891,N_2108);
or U5809 (N_5809,N_2570,N_2365);
or U5810 (N_5810,N_3832,N_2734);
nand U5811 (N_5811,N_2392,N_3557);
nand U5812 (N_5812,N_269,N_1465);
xnor U5813 (N_5813,N_2003,N_3181);
nand U5814 (N_5814,N_4130,N_531);
or U5815 (N_5815,N_3070,N_4615);
nand U5816 (N_5816,N_2292,N_3607);
nor U5817 (N_5817,N_3898,N_899);
or U5818 (N_5818,N_4650,N_3842);
nor U5819 (N_5819,N_414,N_1956);
or U5820 (N_5820,N_355,N_925);
nor U5821 (N_5821,N_4642,N_1103);
xor U5822 (N_5822,N_3375,N_3487);
and U5823 (N_5823,N_3082,N_4186);
nor U5824 (N_5824,N_1110,N_1342);
xor U5825 (N_5825,N_522,N_4172);
nor U5826 (N_5826,N_3500,N_1143);
or U5827 (N_5827,N_161,N_3747);
or U5828 (N_5828,N_3453,N_3139);
or U5829 (N_5829,N_3126,N_4905);
nor U5830 (N_5830,N_363,N_4205);
and U5831 (N_5831,N_1761,N_404);
nor U5832 (N_5832,N_4639,N_4554);
or U5833 (N_5833,N_237,N_4099);
or U5834 (N_5834,N_1495,N_263);
and U5835 (N_5835,N_3382,N_2354);
nor U5836 (N_5836,N_4513,N_4503);
or U5837 (N_5837,N_4387,N_495);
and U5838 (N_5838,N_394,N_3692);
and U5839 (N_5839,N_710,N_17);
nand U5840 (N_5840,N_1327,N_4546);
and U5841 (N_5841,N_3798,N_1732);
or U5842 (N_5842,N_1156,N_4053);
or U5843 (N_5843,N_4737,N_775);
and U5844 (N_5844,N_2283,N_1898);
and U5845 (N_5845,N_3776,N_4166);
or U5846 (N_5846,N_3312,N_1194);
nand U5847 (N_5847,N_1754,N_2353);
xor U5848 (N_5848,N_1897,N_1349);
nor U5849 (N_5849,N_807,N_2820);
and U5850 (N_5850,N_2762,N_422);
and U5851 (N_5851,N_1767,N_2077);
nor U5852 (N_5852,N_728,N_1853);
or U5853 (N_5853,N_48,N_2069);
or U5854 (N_5854,N_3489,N_3645);
xnor U5855 (N_5855,N_1474,N_421);
nand U5856 (N_5856,N_1852,N_588);
nor U5857 (N_5857,N_4702,N_2220);
and U5858 (N_5858,N_220,N_2873);
and U5859 (N_5859,N_3335,N_4878);
nor U5860 (N_5860,N_4311,N_4105);
and U5861 (N_5861,N_3697,N_1030);
and U5862 (N_5862,N_4195,N_1446);
nand U5863 (N_5863,N_1322,N_3705);
xor U5864 (N_5864,N_3857,N_4894);
xnor U5865 (N_5865,N_4,N_83);
nor U5866 (N_5866,N_4331,N_3617);
and U5867 (N_5867,N_661,N_670);
nand U5868 (N_5868,N_867,N_959);
xor U5869 (N_5869,N_3853,N_2912);
nand U5870 (N_5870,N_4868,N_3423);
or U5871 (N_5871,N_131,N_4295);
xnor U5872 (N_5872,N_111,N_2505);
or U5873 (N_5873,N_2480,N_4686);
nor U5874 (N_5874,N_4528,N_3469);
nand U5875 (N_5875,N_1157,N_2210);
nor U5876 (N_5876,N_1986,N_3864);
or U5877 (N_5877,N_4849,N_2891);
nand U5878 (N_5878,N_284,N_3806);
and U5879 (N_5879,N_3091,N_720);
nor U5880 (N_5880,N_2474,N_2050);
xnor U5881 (N_5881,N_1666,N_185);
and U5882 (N_5882,N_3746,N_2232);
xor U5883 (N_5883,N_3131,N_3947);
and U5884 (N_5884,N_2276,N_55);
or U5885 (N_5885,N_1136,N_1300);
or U5886 (N_5886,N_3942,N_3764);
nand U5887 (N_5887,N_1118,N_4015);
or U5888 (N_5888,N_2197,N_528);
and U5889 (N_5889,N_3765,N_2860);
nor U5890 (N_5890,N_1797,N_3623);
nor U5891 (N_5891,N_1184,N_1575);
nand U5892 (N_5892,N_4101,N_3816);
nand U5893 (N_5893,N_4461,N_3425);
and U5894 (N_5894,N_594,N_4677);
nand U5895 (N_5895,N_2317,N_3441);
xor U5896 (N_5896,N_334,N_3051);
nand U5897 (N_5897,N_3860,N_4504);
and U5898 (N_5898,N_1020,N_2363);
or U5899 (N_5899,N_4445,N_3962);
or U5900 (N_5900,N_3213,N_4867);
or U5901 (N_5901,N_4190,N_1205);
or U5902 (N_5902,N_2810,N_2323);
and U5903 (N_5903,N_4201,N_912);
and U5904 (N_5904,N_1996,N_2434);
nand U5905 (N_5905,N_561,N_3829);
nand U5906 (N_5906,N_1905,N_1445);
nand U5907 (N_5907,N_1540,N_4772);
nor U5908 (N_5908,N_2302,N_2099);
nand U5909 (N_5909,N_4917,N_1928);
and U5910 (N_5910,N_4396,N_2482);
or U5911 (N_5911,N_997,N_96);
and U5912 (N_5912,N_1351,N_4774);
and U5913 (N_5913,N_2604,N_1183);
and U5914 (N_5914,N_2245,N_2477);
and U5915 (N_5915,N_4884,N_3022);
or U5916 (N_5916,N_3288,N_3738);
xor U5917 (N_5917,N_517,N_3576);
or U5918 (N_5918,N_836,N_3954);
xor U5919 (N_5919,N_2506,N_2837);
and U5920 (N_5920,N_2088,N_2228);
or U5921 (N_5921,N_3800,N_2114);
or U5922 (N_5922,N_992,N_2263);
and U5923 (N_5923,N_1346,N_4477);
or U5924 (N_5924,N_1337,N_4866);
and U5925 (N_5925,N_3768,N_3331);
nor U5926 (N_5926,N_2622,N_2293);
xnor U5927 (N_5927,N_4152,N_2015);
nand U5928 (N_5928,N_3359,N_1724);
or U5929 (N_5929,N_1280,N_3971);
nand U5930 (N_5930,N_4102,N_4341);
nand U5931 (N_5931,N_1086,N_3778);
nand U5932 (N_5932,N_1916,N_3307);
nand U5933 (N_5933,N_3325,N_2117);
nand U5934 (N_5934,N_1459,N_2180);
nand U5935 (N_5935,N_2794,N_4180);
nor U5936 (N_5936,N_2125,N_3711);
xnor U5937 (N_5937,N_4422,N_582);
and U5938 (N_5938,N_1844,N_923);
nor U5939 (N_5939,N_1181,N_4927);
nand U5940 (N_5940,N_182,N_3867);
nor U5941 (N_5941,N_3363,N_4277);
nor U5942 (N_5942,N_593,N_1161);
and U5943 (N_5943,N_1908,N_4087);
nor U5944 (N_5944,N_4164,N_791);
nor U5945 (N_5945,N_4094,N_3678);
xnor U5946 (N_5946,N_1544,N_1393);
xor U5947 (N_5947,N_1410,N_4624);
nor U5948 (N_5948,N_2564,N_1305);
nor U5949 (N_5949,N_2591,N_1803);
and U5950 (N_5950,N_3053,N_2305);
nor U5951 (N_5951,N_764,N_3239);
or U5952 (N_5952,N_1624,N_852);
or U5953 (N_5953,N_3194,N_1072);
nor U5954 (N_5954,N_4222,N_4096);
nand U5955 (N_5955,N_999,N_219);
and U5956 (N_5956,N_2123,N_4645);
nand U5957 (N_5957,N_2802,N_1821);
nand U5958 (N_5958,N_204,N_2692);
nor U5959 (N_5959,N_3123,N_2744);
and U5960 (N_5960,N_3262,N_1084);
or U5961 (N_5961,N_230,N_4175);
nor U5962 (N_5962,N_779,N_3389);
or U5963 (N_5963,N_2613,N_1515);
xor U5964 (N_5964,N_4749,N_2034);
or U5965 (N_5965,N_3786,N_3455);
xor U5966 (N_5966,N_4865,N_4368);
nand U5967 (N_5967,N_2850,N_62);
and U5968 (N_5968,N_4863,N_4127);
or U5969 (N_5969,N_2189,N_3384);
or U5970 (N_5970,N_3755,N_2449);
nand U5971 (N_5971,N_4493,N_1792);
nor U5972 (N_5972,N_2257,N_4922);
nand U5973 (N_5973,N_1297,N_4874);
and U5974 (N_5974,N_3760,N_2942);
or U5975 (N_5975,N_712,N_3886);
nor U5976 (N_5976,N_1709,N_621);
nand U5977 (N_5977,N_467,N_4790);
nor U5978 (N_5978,N_1751,N_1385);
nor U5979 (N_5979,N_4795,N_3076);
xnor U5980 (N_5980,N_4071,N_3593);
nor U5981 (N_5981,N_2683,N_1583);
nor U5982 (N_5982,N_3365,N_919);
nor U5983 (N_5983,N_68,N_2219);
nand U5984 (N_5984,N_926,N_1914);
nand U5985 (N_5985,N_571,N_2203);
and U5986 (N_5986,N_2215,N_4898);
or U5987 (N_5987,N_4600,N_1069);
and U5988 (N_5988,N_4100,N_4246);
nand U5989 (N_5989,N_3180,N_1341);
nand U5990 (N_5990,N_568,N_2502);
and U5991 (N_5991,N_1436,N_4460);
nand U5992 (N_5992,N_2878,N_4283);
or U5993 (N_5993,N_1774,N_1749);
and U5994 (N_5994,N_88,N_3940);
or U5995 (N_5995,N_767,N_1007);
nand U5996 (N_5996,N_4254,N_871);
xnor U5997 (N_5997,N_4120,N_2425);
nor U5998 (N_5998,N_2445,N_2170);
and U5999 (N_5999,N_1383,N_1179);
nor U6000 (N_6000,N_4383,N_3355);
or U6001 (N_6001,N_4430,N_4549);
or U6002 (N_6002,N_4625,N_3215);
and U6003 (N_6003,N_947,N_1876);
and U6004 (N_6004,N_2634,N_2190);
and U6005 (N_6005,N_1775,N_2223);
nand U6006 (N_6006,N_2372,N_835);
nand U6007 (N_6007,N_1128,N_1646);
and U6008 (N_6008,N_2444,N_2100);
or U6009 (N_6009,N_2527,N_509);
or U6010 (N_6010,N_4183,N_4954);
nor U6011 (N_6011,N_715,N_410);
nand U6012 (N_6012,N_2968,N_765);
or U6013 (N_6013,N_4456,N_4520);
nand U6014 (N_6014,N_1485,N_4271);
or U6015 (N_6015,N_1861,N_2845);
nand U6016 (N_6016,N_2399,N_2789);
or U6017 (N_6017,N_3805,N_3627);
and U6018 (N_6018,N_4594,N_3140);
nand U6019 (N_6019,N_2581,N_1232);
and U6020 (N_6020,N_3961,N_1112);
nor U6021 (N_6021,N_1309,N_4450);
and U6022 (N_6022,N_1170,N_666);
nand U6023 (N_6023,N_1573,N_1978);
and U6024 (N_6024,N_3532,N_1549);
and U6025 (N_6025,N_4580,N_372);
nor U6026 (N_6026,N_3863,N_2741);
and U6027 (N_6027,N_279,N_3788);
nor U6028 (N_6028,N_309,N_2916);
nand U6029 (N_6029,N_2566,N_1373);
xor U6030 (N_6030,N_2739,N_1262);
or U6031 (N_6031,N_893,N_1227);
or U6032 (N_6032,N_2608,N_4457);
nor U6033 (N_6033,N_4397,N_915);
xor U6034 (N_6034,N_411,N_1784);
nor U6035 (N_6035,N_2932,N_4014);
nor U6036 (N_6036,N_10,N_676);
nand U6037 (N_6037,N_1635,N_3709);
xor U6038 (N_6038,N_1878,N_3923);
and U6039 (N_6039,N_1812,N_211);
nor U6040 (N_6040,N_4371,N_1260);
or U6041 (N_6041,N_3132,N_945);
and U6042 (N_6042,N_4364,N_4379);
nand U6043 (N_6043,N_127,N_1159);
nand U6044 (N_6044,N_4338,N_3661);
nand U6045 (N_6045,N_1616,N_151);
or U6046 (N_6046,N_2621,N_4043);
and U6047 (N_6047,N_1622,N_2636);
nor U6048 (N_6048,N_4060,N_4118);
and U6049 (N_6049,N_4569,N_2893);
and U6050 (N_6050,N_3780,N_1875);
or U6051 (N_6051,N_173,N_2075);
xor U6052 (N_6052,N_1892,N_3944);
or U6053 (N_6053,N_2660,N_4342);
or U6054 (N_6054,N_1489,N_3380);
xnor U6055 (N_6055,N_4616,N_2558);
nor U6056 (N_6056,N_2382,N_4265);
and U6057 (N_6057,N_4556,N_320);
and U6058 (N_6058,N_4950,N_3426);
nand U6059 (N_6059,N_1522,N_954);
and U6060 (N_6060,N_2068,N_4561);
nor U6061 (N_6061,N_1509,N_1931);
nand U6062 (N_6062,N_283,N_2731);
or U6063 (N_6063,N_2553,N_1065);
nor U6064 (N_6064,N_4411,N_1819);
and U6065 (N_6065,N_1200,N_3583);
or U6066 (N_6066,N_3563,N_1266);
nor U6067 (N_6067,N_2397,N_981);
or U6068 (N_6068,N_4663,N_2336);
nor U6069 (N_6069,N_2620,N_2769);
nor U6070 (N_6070,N_2246,N_1850);
xor U6071 (N_6071,N_3734,N_2922);
xor U6072 (N_6072,N_4093,N_3859);
xor U6073 (N_6073,N_2499,N_2969);
nand U6074 (N_6074,N_2463,N_3490);
nor U6075 (N_6075,N_4312,N_2486);
and U6076 (N_6076,N_2798,N_41);
nor U6077 (N_6077,N_4025,N_3255);
or U6078 (N_6078,N_2012,N_2307);
nand U6079 (N_6079,N_3631,N_1547);
and U6080 (N_6080,N_328,N_4570);
and U6081 (N_6081,N_3434,N_817);
and U6082 (N_6082,N_3208,N_2826);
or U6083 (N_6083,N_247,N_2199);
or U6084 (N_6084,N_4812,N_1972);
and U6085 (N_6085,N_3254,N_1690);
and U6086 (N_6086,N_4274,N_3019);
nor U6087 (N_6087,N_2401,N_30);
and U6088 (N_6088,N_4010,N_627);
xor U6089 (N_6089,N_481,N_4811);
or U6090 (N_6090,N_1335,N_4735);
or U6091 (N_6091,N_4304,N_4381);
nor U6092 (N_6092,N_3250,N_535);
and U6093 (N_6093,N_1909,N_780);
nor U6094 (N_6094,N_142,N_2978);
nand U6095 (N_6095,N_2699,N_2443);
xnor U6096 (N_6096,N_2572,N_1467);
xor U6097 (N_6097,N_4189,N_4357);
and U6098 (N_6098,N_2150,N_2848);
nor U6099 (N_6099,N_875,N_4154);
and U6100 (N_6100,N_322,N_3395);
nand U6101 (N_6101,N_3603,N_3622);
and U6102 (N_6102,N_564,N_488);
nand U6103 (N_6103,N_4514,N_4602);
nor U6104 (N_6104,N_1943,N_1590);
or U6105 (N_6105,N_4153,N_569);
or U6106 (N_6106,N_4306,N_3400);
nor U6107 (N_6107,N_4004,N_2882);
and U6108 (N_6108,N_4319,N_2568);
or U6109 (N_6109,N_773,N_4563);
and U6110 (N_6110,N_3015,N_3905);
nor U6111 (N_6111,N_2488,N_2089);
nor U6112 (N_6112,N_558,N_300);
and U6113 (N_6113,N_3153,N_1769);
nor U6114 (N_6114,N_4163,N_4358);
nor U6115 (N_6115,N_2290,N_14);
nor U6116 (N_6116,N_2174,N_3702);
nand U6117 (N_6117,N_3014,N_380);
and U6118 (N_6118,N_1427,N_3547);
nand U6119 (N_6119,N_1294,N_1234);
or U6120 (N_6120,N_3894,N_3297);
and U6121 (N_6121,N_1545,N_106);
nor U6122 (N_6122,N_4032,N_4494);
nand U6123 (N_6123,N_4595,N_3205);
nand U6124 (N_6124,N_110,N_901);
nor U6125 (N_6125,N_3956,N_4238);
xnor U6126 (N_6126,N_2578,N_2628);
nor U6127 (N_6127,N_3917,N_19);
nand U6128 (N_6128,N_877,N_1332);
xnor U6129 (N_6129,N_4343,N_1449);
nor U6130 (N_6130,N_1316,N_2112);
xnor U6131 (N_6131,N_3918,N_1223);
and U6132 (N_6132,N_2022,N_4585);
nor U6133 (N_6133,N_4303,N_3706);
xnor U6134 (N_6134,N_4386,N_932);
xor U6135 (N_6135,N_3792,N_1387);
and U6136 (N_6136,N_1602,N_1806);
nor U6137 (N_6137,N_1457,N_2224);
xor U6138 (N_6138,N_393,N_4058);
or U6139 (N_6139,N_2788,N_3021);
nor U6140 (N_6140,N_1333,N_4767);
or U6141 (N_6141,N_2770,N_1648);
nand U6142 (N_6142,N_578,N_750);
and U6143 (N_6143,N_102,N_3865);
or U6144 (N_6144,N_601,N_480);
nand U6145 (N_6145,N_3733,N_1116);
or U6146 (N_6146,N_4144,N_13);
nor U6147 (N_6147,N_1903,N_539);
nand U6148 (N_6148,N_2318,N_235);
and U6149 (N_6149,N_3534,N_4786);
xnor U6150 (N_6150,N_4334,N_3994);
and U6151 (N_6151,N_3095,N_1731);
and U6152 (N_6152,N_2835,N_2954);
and U6153 (N_6153,N_2119,N_2606);
and U6154 (N_6154,N_2970,N_2533);
nand U6155 (N_6155,N_3114,N_878);
xor U6156 (N_6156,N_1323,N_2917);
and U6157 (N_6157,N_2865,N_3067);
or U6158 (N_6158,N_4860,N_2147);
or U6159 (N_6159,N_1154,N_2780);
or U6160 (N_6160,N_329,N_2404);
and U6161 (N_6161,N_186,N_1140);
nand U6162 (N_6162,N_2042,N_4448);
nand U6163 (N_6163,N_520,N_883);
or U6164 (N_6164,N_687,N_924);
or U6165 (N_6165,N_1598,N_2985);
and U6166 (N_6166,N_1991,N_4239);
nand U6167 (N_6167,N_1674,N_1997);
and U6168 (N_6168,N_3998,N_3839);
and U6169 (N_6169,N_3345,N_2380);
xor U6170 (N_6170,N_1293,N_1458);
nand U6171 (N_6171,N_4555,N_963);
or U6172 (N_6172,N_2422,N_280);
xnor U6173 (N_6173,N_4530,N_128);
nand U6174 (N_6174,N_1047,N_2225);
and U6175 (N_6175,N_4081,N_986);
or U6176 (N_6176,N_1151,N_816);
xnor U6177 (N_6177,N_3694,N_2708);
nand U6178 (N_6178,N_1100,N_508);
nor U6179 (N_6179,N_2965,N_1099);
and U6180 (N_6180,N_2665,N_3403);
and U6181 (N_6181,N_326,N_1776);
nor U6182 (N_6182,N_4077,N_2129);
nand U6183 (N_6183,N_4559,N_3241);
nor U6184 (N_6184,N_1017,N_3728);
or U6185 (N_6185,N_4076,N_1279);
and U6186 (N_6186,N_1742,N_4537);
nand U6187 (N_6187,N_443,N_3685);
xnor U6188 (N_6188,N_1703,N_4227);
or U6189 (N_6189,N_3130,N_960);
or U6190 (N_6190,N_691,N_1577);
or U6191 (N_6191,N_281,N_4252);
and U6192 (N_6192,N_3933,N_4613);
xnor U6193 (N_6193,N_2577,N_4510);
nor U6194 (N_6194,N_465,N_224);
nand U6195 (N_6195,N_811,N_3085);
nand U6196 (N_6196,N_4410,N_1016);
nand U6197 (N_6197,N_1236,N_4340);
nor U6198 (N_6198,N_2053,N_2144);
nor U6199 (N_6199,N_3508,N_4640);
nand U6200 (N_6200,N_2806,N_197);
and U6201 (N_6201,N_2994,N_987);
nor U6202 (N_6202,N_2217,N_1499);
and U6203 (N_6203,N_3267,N_1722);
nand U6204 (N_6204,N_662,N_1865);
or U6205 (N_6205,N_40,N_4707);
and U6206 (N_6206,N_4808,N_787);
nand U6207 (N_6207,N_3211,N_2419);
or U6208 (N_6208,N_1566,N_2952);
and U6209 (N_6209,N_1302,N_1764);
nor U6210 (N_6210,N_486,N_1080);
or U6211 (N_6211,N_2306,N_1873);
nand U6212 (N_6212,N_2883,N_1712);
xor U6213 (N_6213,N_2149,N_3825);
nand U6214 (N_6214,N_4788,N_698);
and U6215 (N_6215,N_4064,N_4875);
nor U6216 (N_6216,N_2920,N_1318);
nand U6217 (N_6217,N_514,N_3731);
nand U6218 (N_6218,N_1800,N_3912);
nor U6219 (N_6219,N_545,N_3120);
nor U6220 (N_6220,N_1877,N_1669);
or U6221 (N_6221,N_3980,N_2134);
and U6222 (N_6222,N_2771,N_1630);
nand U6223 (N_6223,N_4885,N_2674);
nor U6224 (N_6224,N_4453,N_699);
and U6225 (N_6225,N_4966,N_3555);
nand U6226 (N_6226,N_1838,N_1477);
nor U6227 (N_6227,N_885,N_3234);
or U6228 (N_6228,N_3221,N_1328);
and U6229 (N_6229,N_43,N_327);
nor U6230 (N_6230,N_2398,N_384);
nor U6231 (N_6231,N_3977,N_2332);
nor U6232 (N_6232,N_117,N_4119);
and U6233 (N_6233,N_1382,N_3018);
or U6234 (N_6234,N_4031,N_441);
or U6235 (N_6235,N_3192,N_4226);
nor U6236 (N_6236,N_2248,N_3527);
and U6237 (N_6237,N_432,N_2605);
and U6238 (N_6238,N_2846,N_1178);
nor U6239 (N_6239,N_2934,N_734);
and U6240 (N_6240,N_137,N_4262);
nand U6241 (N_6241,N_3079,N_1324);
nor U6242 (N_6242,N_3068,N_4792);
and U6243 (N_6243,N_1796,N_2541);
nand U6244 (N_6244,N_2834,N_1375);
and U6245 (N_6245,N_3807,N_2643);
nand U6246 (N_6246,N_2615,N_3158);
nor U6247 (N_6247,N_4662,N_272);
nand U6248 (N_6248,N_4017,N_2694);
nand U6249 (N_6249,N_4566,N_1355);
or U6250 (N_6250,N_4850,N_979);
nand U6251 (N_6251,N_3509,N_4216);
xor U6252 (N_6252,N_3658,N_4416);
nand U6253 (N_6253,N_2728,N_1597);
and U6254 (N_6254,N_680,N_1364);
and U6255 (N_6255,N_487,N_4809);
and U6256 (N_6256,N_3186,N_4009);
and U6257 (N_6257,N_4490,N_2249);
nand U6258 (N_6258,N_1314,N_3633);
or U6259 (N_6259,N_4471,N_2693);
and U6260 (N_6260,N_1263,N_4169);
nor U6261 (N_6261,N_943,N_1158);
nand U6262 (N_6262,N_3450,N_1902);
and U6263 (N_6263,N_4072,N_3828);
and U6264 (N_6264,N_2124,N_2843);
or U6265 (N_6265,N_1250,N_2340);
xor U6266 (N_6266,N_2479,N_1321);
nand U6267 (N_6267,N_4664,N_4041);
nor U6268 (N_6268,N_310,N_3752);
nand U6269 (N_6269,N_4257,N_1862);
xor U6270 (N_6270,N_4818,N_321);
and U6271 (N_6271,N_4002,N_1623);
and U6272 (N_6272,N_3559,N_3703);
xor U6273 (N_6273,N_3590,N_1691);
nand U6274 (N_6274,N_557,N_1650);
or U6275 (N_6275,N_3122,N_1174);
nand U6276 (N_6276,N_3197,N_3882);
or U6277 (N_6277,N_884,N_4576);
or U6278 (N_6278,N_1348,N_461);
nor U6279 (N_6279,N_1012,N_2241);
nand U6280 (N_6280,N_2331,N_3979);
and U6281 (N_6281,N_813,N_4909);
and U6282 (N_6282,N_1468,N_2335);
or U6283 (N_6283,N_1516,N_387);
or U6284 (N_6284,N_3185,N_1462);
nand U6285 (N_6285,N_1925,N_1035);
nand U6286 (N_6286,N_4584,N_3574);
nor U6287 (N_6287,N_1138,N_2173);
xnor U6288 (N_6288,N_2750,N_1658);
or U6289 (N_6289,N_2328,N_3507);
nand U6290 (N_6290,N_881,N_4019);
nor U6291 (N_6291,N_4746,N_1998);
and U6292 (N_6292,N_554,N_4155);
nor U6293 (N_6293,N_3849,N_637);
xor U6294 (N_6294,N_1340,N_553);
nor U6295 (N_6295,N_4052,N_2679);
and U6296 (N_6296,N_335,N_3506);
and U6297 (N_6297,N_2179,N_285);
or U6298 (N_6298,N_4560,N_239);
nor U6299 (N_6299,N_1727,N_2763);
or U6300 (N_6300,N_4465,N_424);
and U6301 (N_6301,N_4900,N_4214);
or U6302 (N_6302,N_985,N_1922);
nor U6303 (N_6303,N_3513,N_1744);
or U6304 (N_6304,N_4726,N_2281);
nand U6305 (N_6305,N_1420,N_4699);
and U6306 (N_6306,N_12,N_574);
nor U6307 (N_6307,N_3253,N_2265);
or U6308 (N_6308,N_1678,N_3826);
or U6309 (N_6309,N_1377,N_950);
and U6310 (N_6310,N_3784,N_339);
and U6311 (N_6311,N_1166,N_1526);
or U6312 (N_6312,N_4443,N_908);
nand U6313 (N_6313,N_4604,N_4112);
nor U6314 (N_6314,N_3858,N_3447);
nand U6315 (N_6315,N_2575,N_616);
and U6316 (N_6316,N_178,N_259);
and U6317 (N_6317,N_4533,N_3537);
and U6318 (N_6318,N_3899,N_1655);
or U6319 (N_6319,N_2453,N_3268);
and U6320 (N_6320,N_1171,N_4886);
and U6321 (N_6321,N_4173,N_1699);
and U6322 (N_6322,N_1469,N_4036);
nand U6323 (N_6323,N_703,N_2513);
nor U6324 (N_6324,N_2905,N_1147);
nor U6325 (N_6325,N_3960,N_4223);
xnor U6326 (N_6326,N_4829,N_2400);
nand U6327 (N_6327,N_3340,N_897);
nand U6328 (N_6328,N_2535,N_1705);
nand U6329 (N_6329,N_2346,N_1820);
nor U6330 (N_6330,N_2614,N_2979);
or U6331 (N_6331,N_2709,N_2807);
nand U6332 (N_6332,N_4629,N_4297);
nand U6333 (N_6333,N_434,N_2330);
nand U6334 (N_6334,N_1471,N_4499);
and U6335 (N_6335,N_3561,N_4403);
nand U6336 (N_6336,N_3072,N_4738);
nor U6337 (N_6337,N_3436,N_532);
xor U6338 (N_6338,N_3605,N_3102);
and U6339 (N_6339,N_3793,N_4815);
nand U6340 (N_6340,N_1514,N_200);
and U6341 (N_6341,N_1391,N_104);
or U6342 (N_6342,N_1278,N_472);
or U6343 (N_6343,N_4373,N_1399);
nand U6344 (N_6344,N_4531,N_1938);
or U6345 (N_6345,N_1186,N_994);
nor U6346 (N_6346,N_278,N_3156);
and U6347 (N_6347,N_898,N_826);
and U6348 (N_6348,N_2115,N_4722);
nor U6349 (N_6349,N_3936,N_428);
nand U6350 (N_6350,N_2925,N_1374);
or U6351 (N_6351,N_4906,N_2260);
xor U6352 (N_6352,N_2675,N_1772);
nand U6353 (N_6353,N_916,N_4209);
nand U6354 (N_6354,N_2625,N_3160);
xor U6355 (N_6355,N_3318,N_4719);
nand U6356 (N_6356,N_3020,N_4168);
nand U6357 (N_6357,N_2024,N_3723);
and U6358 (N_6358,N_1439,N_620);
and U6359 (N_6359,N_4575,N_1326);
or U6360 (N_6360,N_4890,N_1032);
nand U6361 (N_6361,N_549,N_3966);
or U6362 (N_6362,N_2992,N_640);
xnor U6363 (N_6363,N_1934,N_2937);
or U6364 (N_6364,N_2141,N_2465);
nand U6365 (N_6365,N_159,N_3200);
nor U6366 (N_6366,N_812,N_1443);
or U6367 (N_6367,N_4793,N_4228);
xnor U6368 (N_6368,N_1146,N_3924);
nand U6369 (N_6369,N_1675,N_600);
nand U6370 (N_6370,N_2704,N_3443);
nor U6371 (N_6371,N_2832,N_576);
or U6372 (N_6372,N_3794,N_4469);
and U6373 (N_6373,N_3757,N_1660);
xnor U6374 (N_6374,N_1859,N_4027);
nor U6375 (N_6375,N_129,N_4720);
nand U6376 (N_6376,N_1287,N_1531);
nor U6377 (N_6377,N_25,N_4951);
and U6378 (N_6378,N_2211,N_144);
or U6379 (N_6379,N_1339,N_2140);
or U6380 (N_6380,N_2587,N_1228);
and U6381 (N_6381,N_4011,N_1628);
nor U6382 (N_6382,N_573,N_678);
nor U6383 (N_6383,N_4607,N_4260);
and U6384 (N_6384,N_2913,N_4370);
nor U6385 (N_6385,N_3551,N_4992);
nor U6386 (N_6386,N_1518,N_2300);
and U6387 (N_6387,N_903,N_1948);
xnor U6388 (N_6388,N_4243,N_2371);
and U6389 (N_6389,N_1344,N_2765);
and U6390 (N_6390,N_1074,N_3775);
and U6391 (N_6391,N_4690,N_2358);
or U6392 (N_6392,N_354,N_4638);
and U6393 (N_6393,N_4407,N_719);
nand U6394 (N_6394,N_3298,N_3499);
or U6395 (N_6395,N_2234,N_1605);
and U6396 (N_6396,N_4841,N_492);
nor U6397 (N_6397,N_3439,N_38);
and U6398 (N_6398,N_4963,N_4307);
nor U6399 (N_6399,N_2230,N_228);
or U6400 (N_6400,N_2011,N_4778);
nand U6401 (N_6401,N_2494,N_4761);
or U6402 (N_6402,N_4425,N_299);
nor U6403 (N_6403,N_1847,N_1370);
nand U6404 (N_6404,N_474,N_2264);
or U6405 (N_6405,N_2347,N_3379);
or U6406 (N_6406,N_4925,N_2402);
and U6407 (N_6407,N_4247,N_4497);
nor U6408 (N_6408,N_3491,N_3843);
and U6409 (N_6409,N_2639,N_1401);
xnor U6410 (N_6410,N_4244,N_4591);
nand U6411 (N_6411,N_4717,N_4428);
nand U6412 (N_6412,N_4451,N_2006);
nand U6413 (N_6413,N_2187,N_4097);
nand U6414 (N_6414,N_2532,N_537);
nand U6415 (N_6415,N_463,N_3599);
or U6416 (N_6416,N_3901,N_141);
nor U6417 (N_6417,N_3877,N_974);
or U6418 (N_6418,N_902,N_2379);
nand U6419 (N_6419,N_1406,N_2233);
xnor U6420 (N_6420,N_1434,N_1939);
xnor U6421 (N_6421,N_2029,N_3660);
and U6422 (N_6422,N_1855,N_1656);
or U6423 (N_6423,N_2823,N_3913);
nand U6424 (N_6424,N_1267,N_4286);
and U6425 (N_6425,N_500,N_4914);
nand U6426 (N_6426,N_2164,N_1836);
nor U6427 (N_6427,N_2350,N_847);
or U6428 (N_6428,N_2701,N_894);
nor U6429 (N_6429,N_475,N_4328);
and U6430 (N_6430,N_152,N_4467);
and U6431 (N_6431,N_3779,N_3567);
or U6432 (N_6432,N_1974,N_4489);
nand U6433 (N_6433,N_126,N_2344);
and U6434 (N_6434,N_3240,N_3421);
or U6435 (N_6435,N_4131,N_4308);
and U6436 (N_6436,N_147,N_3742);
and U6437 (N_6437,N_758,N_3596);
xnor U6438 (N_6438,N_4658,N_3387);
nand U6439 (N_6439,N_2009,N_4349);
and U6440 (N_6440,N_2529,N_302);
nor U6441 (N_6441,N_1854,N_3098);
or U6442 (N_6442,N_1274,N_2163);
and U6443 (N_6443,N_2478,N_1371);
nor U6444 (N_6444,N_646,N_4050);
and U6445 (N_6445,N_3121,N_2370);
nor U6446 (N_6446,N_1251,N_1976);
or U6447 (N_6447,N_2959,N_2712);
and U6448 (N_6448,N_2037,N_4654);
nand U6449 (N_6449,N_1716,N_4899);
or U6450 (N_6450,N_2557,N_2118);
xor U6451 (N_6451,N_2811,N_324);
xor U6452 (N_6452,N_1085,N_1115);
xnor U6453 (N_6453,N_1270,N_3684);
and U6454 (N_6454,N_944,N_3715);
nor U6455 (N_6455,N_2815,N_2722);
nand U6456 (N_6456,N_1369,N_3795);
or U6457 (N_6457,N_1312,N_3544);
nor U6458 (N_6458,N_1480,N_4256);
and U6459 (N_6459,N_3837,N_1380);
nor U6460 (N_6460,N_3582,N_1247);
and U6461 (N_6461,N_2617,N_427);
and U6462 (N_6462,N_690,N_479);
nor U6463 (N_6463,N_1857,N_1899);
nand U6464 (N_6464,N_3404,N_2098);
or U6465 (N_6465,N_2128,N_4398);
nand U6466 (N_6466,N_3259,N_3774);
nor U6467 (N_6467,N_4480,N_4807);
nand U6468 (N_6468,N_1336,N_271);
nand U6469 (N_6469,N_3833,N_1285);
nand U6470 (N_6470,N_1860,N_2198);
nor U6471 (N_6471,N_2819,N_3106);
xnor U6472 (N_6472,N_3339,N_2803);
and U6473 (N_6473,N_1024,N_2539);
and U6474 (N_6474,N_2791,N_2031);
nor U6475 (N_6475,N_771,N_599);
and U6476 (N_6476,N_4290,N_67);
nand U6477 (N_6477,N_4039,N_2742);
nor U6478 (N_6478,N_3148,N_3758);
xnor U6479 (N_6479,N_4676,N_3789);
xnor U6480 (N_6480,N_1782,N_3571);
xor U6481 (N_6481,N_2706,N_71);
and U6482 (N_6482,N_1508,N_2270);
or U6483 (N_6483,N_1165,N_784);
nor U6484 (N_6484,N_1593,N_3570);
or U6485 (N_6485,N_636,N_3579);
and U6486 (N_6486,N_2957,N_2322);
nor U6487 (N_6487,N_483,N_1175);
xor U6488 (N_6488,N_2256,N_2730);
xor U6489 (N_6489,N_2131,N_656);
or U6490 (N_6490,N_697,N_2026);
nand U6491 (N_6491,N_1002,N_3486);
nor U6492 (N_6492,N_3879,N_3162);
nor U6493 (N_6493,N_3602,N_2238);
nand U6494 (N_6494,N_772,N_3460);
nand U6495 (N_6495,N_688,N_3212);
nand U6496 (N_6496,N_3615,N_524);
or U6497 (N_6497,N_3218,N_4752);
and U6498 (N_6498,N_3817,N_832);
and U6499 (N_6499,N_3115,N_1689);
nand U6500 (N_6500,N_4219,N_4679);
nand U6501 (N_6501,N_4199,N_2231);
nor U6502 (N_6502,N_3407,N_2039);
and U6503 (N_6503,N_1163,N_4399);
xor U6504 (N_6504,N_3845,N_4631);
and U6505 (N_6505,N_2072,N_4547);
and U6506 (N_6506,N_4703,N_3665);
or U6507 (N_6507,N_4876,N_2369);
nor U6508 (N_6508,N_2454,N_4151);
or U6509 (N_6509,N_880,N_3134);
and U6510 (N_6510,N_2275,N_1941);
xor U6511 (N_6511,N_4947,N_3002);
xor U6512 (N_6512,N_4725,N_4568);
nor U6513 (N_6513,N_1288,N_4562);
and U6514 (N_6514,N_175,N_4404);
nor U6515 (N_6515,N_1618,N_2221);
or U6516 (N_6516,N_2512,N_3978);
nand U6517 (N_6517,N_1193,N_4241);
nor U6518 (N_6518,N_2800,N_2060);
nor U6519 (N_6519,N_4478,N_3637);
nand U6520 (N_6520,N_4840,N_1781);
nand U6521 (N_6521,N_4518,N_4409);
or U6522 (N_6522,N_3771,N_3462);
nand U6523 (N_6523,N_717,N_2277);
or U6524 (N_6524,N_4796,N_2751);
nand U6525 (N_6525,N_1207,N_4806);
nor U6526 (N_6526,N_2359,N_795);
xnor U6527 (N_6527,N_672,N_3552);
nand U6528 (N_6528,N_2776,N_3716);
or U6529 (N_6529,N_4961,N_544);
or U6530 (N_6530,N_4345,N_1040);
xor U6531 (N_6531,N_2329,N_3454);
and U6532 (N_6532,N_3546,N_1216);
or U6533 (N_6533,N_20,N_857);
nor U6534 (N_6534,N_2867,N_205);
or U6535 (N_6535,N_3553,N_3152);
nor U6536 (N_6536,N_2195,N_2618);
nand U6537 (N_6537,N_2852,N_1191);
or U6538 (N_6538,N_4269,N_54);
nor U6539 (N_6539,N_2801,N_3299);
and U6540 (N_6540,N_4593,N_859);
xor U6541 (N_6541,N_2239,N_3396);
nand U6542 (N_6542,N_1306,N_4827);
and U6543 (N_6543,N_1180,N_1750);
or U6544 (N_6544,N_4424,N_3921);
nor U6545 (N_6545,N_362,N_99);
or U6546 (N_6546,N_1130,N_2902);
and U6547 (N_6547,N_4852,N_2355);
and U6548 (N_6548,N_1966,N_4583);
nand U6549 (N_6549,N_2673,N_460);
xor U6550 (N_6550,N_3488,N_273);
and U6551 (N_6551,N_1794,N_4066);
and U6552 (N_6552,N_831,N_2766);
or U6553 (N_6553,N_1808,N_125);
nand U6554 (N_6554,N_2291,N_2167);
xnor U6555 (N_6555,N_3608,N_3620);
nand U6556 (N_6556,N_4748,N_504);
or U6557 (N_6557,N_1557,N_4392);
nand U6558 (N_6558,N_1054,N_2595);
or U6559 (N_6559,N_4972,N_4104);
and U6560 (N_6560,N_2327,N_4921);
nor U6561 (N_6561,N_1435,N_3108);
and U6562 (N_6562,N_2991,N_3688);
nor U6563 (N_6563,N_287,N_1215);
nor U6564 (N_6564,N_4082,N_165);
nor U6565 (N_6565,N_1009,N_2004);
nor U6566 (N_6566,N_2646,N_1787);
or U6567 (N_6567,N_4578,N_1894);
nand U6568 (N_6568,N_3063,N_1365);
nand U6569 (N_6569,N_1721,N_3663);
or U6570 (N_6570,N_3970,N_2483);
nor U6571 (N_6571,N_3543,N_4292);
nand U6572 (N_6572,N_114,N_834);
nand U6573 (N_6573,N_4525,N_502);
or U6574 (N_6574,N_657,N_4523);
nor U6575 (N_6575,N_4579,N_2869);
and U6576 (N_6576,N_440,N_1281);
nand U6577 (N_6577,N_426,N_1893);
and U6578 (N_6578,N_45,N_225);
nor U6579 (N_6579,N_1620,N_1694);
nand U6580 (N_6580,N_2594,N_1957);
nand U6581 (N_6581,N_103,N_2645);
or U6582 (N_6582,N_3495,N_3982);
nor U6583 (N_6583,N_446,N_904);
or U6584 (N_6584,N_60,N_353);
nand U6585 (N_6585,N_2707,N_3797);
nand U6586 (N_6586,N_1329,N_3972);
or U6587 (N_6587,N_3959,N_3516);
xnor U6588 (N_6588,N_4977,N_4723);
xnor U6589 (N_6589,N_81,N_4710);
and U6590 (N_6590,N_4150,N_2656);
or U6591 (N_6591,N_3187,N_430);
or U6592 (N_6592,N_1537,N_2997);
nor U6593 (N_6593,N_2659,N_1398);
and U6594 (N_6594,N_359,N_4848);
nor U6595 (N_6595,N_4916,N_1707);
nor U6596 (N_6596,N_2671,N_207);
or U6597 (N_6597,N_4136,N_4801);
xor U6598 (N_6598,N_3796,N_4367);
and U6599 (N_6599,N_337,N_347);
nor U6600 (N_6600,N_2672,N_3804);
or U6601 (N_6601,N_1463,N_2988);
nand U6602 (N_6602,N_2385,N_972);
xnor U6603 (N_6603,N_3987,N_2186);
and U6604 (N_6604,N_2829,N_3310);
and U6605 (N_6605,N_1039,N_1783);
nand U6606 (N_6606,N_521,N_1317);
nand U6607 (N_6607,N_2325,N_392);
or U6608 (N_6608,N_113,N_4543);
and U6609 (N_6609,N_1641,N_3494);
nand U6610 (N_6610,N_3290,N_939);
or U6611 (N_6611,N_1425,N_4923);
nand U6612 (N_6612,N_4487,N_3145);
or U6613 (N_6613,N_1633,N_4301);
nor U6614 (N_6614,N_2421,N_1481);
and U6615 (N_6615,N_874,N_705);
nor U6616 (N_6616,N_3740,N_2530);
or U6617 (N_6617,N_575,N_398);
or U6618 (N_6618,N_619,N_6);
or U6619 (N_6619,N_931,N_1798);
and U6620 (N_6620,N_1614,N_2567);
or U6621 (N_6621,N_1521,N_2999);
and U6622 (N_6622,N_2517,N_3803);
and U6623 (N_6623,N_4067,N_138);
nor U6624 (N_6624,N_3597,N_3503);
or U6625 (N_6625,N_1091,N_115);
and U6626 (N_6626,N_2237,N_2172);
or U6627 (N_6627,N_626,N_935);
or U6628 (N_6628,N_4128,N_160);
or U6629 (N_6629,N_4113,N_0);
nand U6630 (N_6630,N_395,N_1070);
and U6631 (N_6631,N_3333,N_3023);
and U6632 (N_6632,N_4211,N_1572);
or U6633 (N_6633,N_2364,N_189);
nor U6634 (N_6634,N_1192,N_798);
nand U6635 (N_6635,N_413,N_2521);
nor U6636 (N_6636,N_29,N_4212);
nand U6637 (N_6637,N_4107,N_2262);
and U6638 (N_6638,N_1816,N_2055);
or U6639 (N_6639,N_3081,N_4655);
and U6640 (N_6640,N_3449,N_2352);
or U6641 (N_6641,N_1708,N_262);
and U6642 (N_6642,N_1289,N_4353);
nand U6643 (N_6643,N_4614,N_3274);
nand U6644 (N_6644,N_4156,N_1087);
nor U6645 (N_6645,N_2793,N_2732);
xor U6646 (N_6646,N_707,N_815);
nor U6647 (N_6647,N_838,N_1830);
nor U6648 (N_6648,N_789,N_2151);
xnor U6649 (N_6649,N_2038,N_3378);
nand U6650 (N_6650,N_3748,N_696);
and U6651 (N_6651,N_3005,N_155);
and U6652 (N_6652,N_747,N_1350);
nor U6653 (N_6653,N_2929,N_4324);
xnor U6654 (N_6654,N_90,N_4325);
nor U6655 (N_6655,N_4486,N_4419);
or U6656 (N_6656,N_1233,N_3026);
and U6657 (N_6657,N_2809,N_4505);
nand U6658 (N_6658,N_2918,N_3642);
or U6659 (N_6659,N_3110,N_819);
and U6660 (N_6660,N_3295,N_2475);
nor U6661 (N_6661,N_3006,N_4536);
nand U6662 (N_6662,N_4016,N_2551);
xor U6663 (N_6663,N_679,N_2008);
nor U6664 (N_6664,N_1135,N_1988);
and U6665 (N_6665,N_973,N_1920);
and U6666 (N_6666,N_2759,N_2836);
nor U6667 (N_6667,N_3007,N_1005);
nor U6668 (N_6668,N_1802,N_4115);
nand U6669 (N_6669,N_740,N_3854);
nor U6670 (N_6670,N_1376,N_1137);
or U6671 (N_6671,N_4833,N_415);
nand U6672 (N_6672,N_4508,N_340);
or U6673 (N_6673,N_1651,N_4763);
or U6674 (N_6674,N_2430,N_855);
and U6675 (N_6675,N_1534,N_911);
or U6676 (N_6676,N_2090,N_505);
nand U6677 (N_6677,N_3493,N_1198);
and U6678 (N_6678,N_3872,N_4883);
or U6679 (N_6679,N_2431,N_4873);
or U6680 (N_6680,N_2476,N_3484);
or U6681 (N_6681,N_4995,N_3301);
nor U6682 (N_6682,N_4913,N_1004);
nor U6683 (N_6683,N_3919,N_2240);
nor U6684 (N_6684,N_1672,N_2074);
nand U6685 (N_6685,N_1360,N_1148);
nand U6686 (N_6686,N_2395,N_2995);
xnor U6687 (N_6687,N_3100,N_1413);
or U6688 (N_6688,N_1248,N_3027);
nor U6689 (N_6689,N_2446,N_3581);
or U6690 (N_6690,N_2740,N_1935);
and U6691 (N_6691,N_2927,N_618);
and U6692 (N_6692,N_4202,N_2949);
nand U6693 (N_6693,N_3452,N_2666);
and U6694 (N_6694,N_2822,N_1366);
nor U6695 (N_6695,N_3904,N_3398);
nor U6696 (N_6696,N_2839,N_3639);
nor U6697 (N_6697,N_842,N_1464);
nand U6698 (N_6698,N_4395,N_2879);
nor U6699 (N_6699,N_4145,N_146);
and U6700 (N_6700,N_4160,N_4529);
nor U6701 (N_6701,N_4047,N_3533);
or U6702 (N_6702,N_3984,N_2019);
or U6703 (N_6703,N_2962,N_956);
nor U6704 (N_6704,N_1048,N_156);
nor U6705 (N_6705,N_1075,N_526);
and U6706 (N_6706,N_3589,N_2588);
and U6707 (N_6707,N_2338,N_4783);
and U6708 (N_6708,N_1442,N_3164);
nor U6709 (N_6709,N_1827,N_726);
or U6710 (N_6710,N_4753,N_2641);
or U6711 (N_6711,N_1090,N_4770);
nand U6712 (N_6712,N_4090,N_3109);
nor U6713 (N_6713,N_1417,N_464);
nand U6714 (N_6714,N_3974,N_615);
nand U6715 (N_6715,N_3686,N_3868);
nand U6716 (N_6716,N_3895,N_3540);
and U6717 (N_6717,N_2205,N_4953);
xnor U6718 (N_6718,N_792,N_364);
or U6719 (N_6719,N_3346,N_4026);
or U6720 (N_6720,N_4751,N_4837);
nor U6721 (N_6721,N_4114,N_86);
or U6722 (N_6722,N_3953,N_4744);
nor U6723 (N_6723,N_1824,N_4361);
nor U6724 (N_6724,N_2511,N_3195);
or U6725 (N_6725,N_829,N_4558);
xor U6726 (N_6726,N_2972,N_2736);
nand U6727 (N_6727,N_2721,N_4620);
and U6728 (N_6728,N_4366,N_4162);
nor U6729 (N_6729,N_2667,N_503);
or U6730 (N_6730,N_1706,N_2559);
and U6731 (N_6731,N_3861,N_3497);
and U6732 (N_6732,N_2814,N_4013);
nand U6733 (N_6733,N_1064,N_4601);
and U6734 (N_6734,N_4715,N_2014);
nand U6735 (N_6735,N_2632,N_2432);
nor U6736 (N_6736,N_2764,N_4539);
nor U6737 (N_6737,N_3717,N_4776);
nor U6738 (N_6738,N_1440,N_3928);
nand U6739 (N_6739,N_2565,N_2631);
nand U6740 (N_6740,N_3963,N_1807);
or U6741 (N_6741,N_3587,N_4089);
and U6742 (N_6742,N_4994,N_4509);
and U6743 (N_6743,N_2360,N_3225);
nand U6744 (N_6744,N_3144,N_2218);
nand U6745 (N_6745,N_188,N_1995);
nor U6746 (N_6746,N_2574,N_1888);
and U6747 (N_6747,N_3272,N_3946);
nor U6748 (N_6748,N_607,N_1686);
nand U6749 (N_6749,N_1225,N_3504);
or U6750 (N_6750,N_4816,N_4773);
and U6751 (N_6751,N_1296,N_250);
or U6752 (N_6752,N_4844,N_3874);
or U6753 (N_6753,N_3750,N_1872);
nand U6754 (N_6754,N_3827,N_4766);
and U6755 (N_6755,N_3600,N_2096);
nand U6756 (N_6756,N_4731,N_2155);
nor U6757 (N_6757,N_2165,N_3038);
nand U6758 (N_6758,N_4997,N_1835);
or U6759 (N_6759,N_2911,N_2130);
and U6760 (N_6760,N_1389,N_2700);
or U6761 (N_6761,N_2904,N_667);
nand U6762 (N_6762,N_2497,N_3808);
nor U6763 (N_6763,N_2315,N_853);
xnor U6764 (N_6764,N_3011,N_3695);
nand U6765 (N_6765,N_1320,N_304);
and U6766 (N_6766,N_4063,N_1390);
nand U6767 (N_6767,N_2160,N_2268);
and U6768 (N_6768,N_3226,N_753);
or U6769 (N_6769,N_1904,N_3586);
nor U6770 (N_6770,N_1241,N_2243);
nand U6771 (N_6771,N_1770,N_2313);
nor U6772 (N_6772,N_3433,N_3256);
and U6773 (N_6773,N_4644,N_1626);
or U6774 (N_6774,N_4912,N_3017);
and U6775 (N_6775,N_4165,N_3366);
or U6776 (N_6776,N_4826,N_2045);
or U6777 (N_6777,N_1164,N_2367);
nand U6778 (N_6778,N_2562,N_3939);
nor U6779 (N_6779,N_361,N_4048);
nand U6780 (N_6780,N_2609,N_4485);
or U6781 (N_6781,N_2166,N_3417);
or U6782 (N_6782,N_367,N_312);
nor U6783 (N_6783,N_1801,N_3935);
nand U6784 (N_6784,N_4764,N_3418);
nand U6785 (N_6785,N_3916,N_4728);
and U6786 (N_6786,N_2394,N_2658);
xor U6787 (N_6787,N_3884,N_642);
and U6788 (N_6788,N_3111,N_1924);
xnor U6789 (N_6789,N_611,N_1880);
nor U6790 (N_6790,N_3564,N_4821);
or U6791 (N_6791,N_581,N_4429);
or U6792 (N_6792,N_1748,N_4270);
nand U6793 (N_6793,N_2348,N_4565);
and U6794 (N_6794,N_3949,N_198);
or U6795 (N_6795,N_3003,N_87);
or U6796 (N_6796,N_4780,N_2301);
xnor U6797 (N_6797,N_2715,N_388);
xor U6798 (N_6798,N_4174,N_3296);
and U6799 (N_6799,N_3058,N_1874);
nor U6800 (N_6800,N_4622,N_2896);
and U6801 (N_6801,N_4993,N_1010);
nor U6802 (N_6802,N_1222,N_437);
nor U6803 (N_6803,N_2561,N_192);
nand U6804 (N_6804,N_4446,N_969);
nor U6805 (N_6805,N_169,N_1405);
xnor U6806 (N_6806,N_684,N_1491);
xnor U6807 (N_6807,N_1212,N_2950);
nor U6808 (N_6808,N_2892,N_2973);
and U6809 (N_6809,N_2222,N_3336);
xor U6810 (N_6810,N_3680,N_2573);
nor U6811 (N_6811,N_2058,N_4526);
nor U6812 (N_6812,N_3915,N_850);
nor U6813 (N_6813,N_3720,N_3910);
and U6814 (N_6814,N_3028,N_742);
nand U6815 (N_6815,N_2772,N_305);
and U6816 (N_6816,N_356,N_2161);
and U6817 (N_6817,N_357,N_251);
nand U6818 (N_6818,N_4051,N_2947);
or U6819 (N_6819,N_808,N_3171);
and U6820 (N_6820,N_3088,N_453);
nand U6821 (N_6821,N_3202,N_3862);
and U6822 (N_6822,N_2945,N_3177);
nor U6823 (N_6823,N_3059,N_551);
and U6824 (N_6824,N_2680,N_4447);
or U6825 (N_6825,N_4298,N_1528);
or U6826 (N_6826,N_4207,N_1152);
or U6827 (N_6827,N_4108,N_69);
nand U6828 (N_6828,N_132,N_4522);
and U6829 (N_6829,N_1755,N_937);
nand U6830 (N_6830,N_3766,N_1559);
nor U6831 (N_6831,N_2847,N_861);
or U6832 (N_6832,N_3414,N_4851);
and U6833 (N_6833,N_519,N_3585);
and U6834 (N_6834,N_763,N_2868);
nor U6835 (N_6835,N_1985,N_4958);
or U6836 (N_6836,N_1408,N_1036);
or U6837 (N_6837,N_2703,N_606);
nor U6838 (N_6838,N_3337,N_4412);
and U6839 (N_6839,N_341,N_255);
or U6840 (N_6840,N_2408,N_1496);
nand U6841 (N_6841,N_1133,N_2757);
nand U6842 (N_6842,N_1737,N_1430);
nor U6843 (N_6843,N_1504,N_190);
nor U6844 (N_6844,N_3496,N_2547);
nand U6845 (N_6845,N_2462,N_863);
and U6846 (N_6846,N_4691,N_786);
nor U6847 (N_6847,N_1403,N_4458);
nand U6848 (N_6848,N_1982,N_4121);
and U6849 (N_6849,N_4421,N_3357);
nand U6850 (N_6850,N_2812,N_218);
xnor U6851 (N_6851,N_1076,N_3401);
nand U6852 (N_6852,N_2629,N_2103);
or U6853 (N_6853,N_3385,N_4313);
or U6854 (N_6854,N_462,N_702);
xnor U6855 (N_6855,N_3065,N_3897);
and U6856 (N_6856,N_2261,N_1044);
or U6857 (N_6857,N_2059,N_1490);
xor U6858 (N_6858,N_2094,N_3927);
nand U6859 (N_6859,N_2247,N_1663);
and U6860 (N_6860,N_4970,N_291);
or U6861 (N_6861,N_1210,N_4170);
nand U6862 (N_6862,N_4061,N_193);
or U6863 (N_6863,N_1258,N_3348);
nor U6864 (N_6864,N_1506,N_85);
or U6865 (N_6865,N_1343,N_1230);
and U6866 (N_6866,N_776,N_3456);
or U6867 (N_6867,N_1249,N_233);
and U6868 (N_6868,N_2910,N_1345);
nand U6869 (N_6869,N_118,N_2797);
or U6870 (N_6870,N_2576,N_4597);
and U6871 (N_6871,N_1845,N_3871);
or U6872 (N_6872,N_1470,N_2849);
nor U6873 (N_6873,N_4777,N_3252);
and U6874 (N_6874,N_3432,N_3232);
nor U6875 (N_6875,N_3459,N_2303);
and U6876 (N_6876,N_162,N_694);
or U6877 (N_6877,N_2152,N_4106);
nand U6878 (N_6878,N_2790,N_97);
or U6879 (N_6879,N_882,N_3381);
xor U6880 (N_6880,N_433,N_4294);
and U6881 (N_6881,N_2070,N_689);
nor U6882 (N_6882,N_1958,N_4003);
nand U6883 (N_6883,N_3319,N_3993);
and U6884 (N_6884,N_444,N_683);
nand U6885 (N_6885,N_975,N_887);
nor U6886 (N_6886,N_1096,N_4924);
nor U6887 (N_6887,N_746,N_2405);
and U6888 (N_6888,N_3967,N_2940);
or U6889 (N_6889,N_3802,N_3214);
and U6890 (N_6890,N_2907,N_4146);
and U6891 (N_6891,N_1209,N_2406);
nor U6892 (N_6892,N_2684,N_1562);
nor U6893 (N_6893,N_1268,N_148);
and U6894 (N_6894,N_3890,N_3420);
nor U6895 (N_6895,N_4672,N_419);
xor U6896 (N_6896,N_2175,N_1882);
xnor U6897 (N_6897,N_2754,N_602);
nor U6898 (N_6898,N_4635,N_456);
nor U6899 (N_6899,N_2687,N_1846);
and U6900 (N_6900,N_4138,N_4384);
and U6901 (N_6901,N_4705,N_1144);
and U6902 (N_6902,N_1681,N_907);
nand U6903 (N_6903,N_2876,N_3260);
nand U6904 (N_6904,N_1052,N_3300);
and U6905 (N_6905,N_3475,N_2082);
or U6906 (N_6906,N_4192,N_4666);
or U6907 (N_6907,N_1513,N_1581);
nand U6908 (N_6908,N_1980,N_3413);
and U6909 (N_6909,N_3830,N_294);
and U6910 (N_6910,N_4420,N_1989);
nor U6911 (N_6911,N_4567,N_4949);
and U6912 (N_6912,N_4678,N_3471);
or U6913 (N_6913,N_1643,N_1394);
and U6914 (N_6914,N_868,N_4500);
or U6915 (N_6915,N_3409,N_1068);
and U6916 (N_6916,N_3182,N_1357);
xnor U6917 (N_6917,N_711,N_1640);
xor U6918 (N_6918,N_2747,N_4231);
and U6919 (N_6919,N_1981,N_4030);
nand U6920 (N_6920,N_107,N_2676);
nor U6921 (N_6921,N_7,N_2654);
xnor U6922 (N_6922,N_1219,N_2110);
nor U6923 (N_6923,N_196,N_4765);
nor U6924 (N_6924,N_2286,N_4359);
nand U6925 (N_6925,N_348,N_3291);
or U6926 (N_6926,N_1386,N_4390);
xnor U6927 (N_6927,N_4843,N_2951);
nor U6928 (N_6928,N_286,N_4157);
and U6929 (N_6929,N_2590,N_130);
and U6930 (N_6930,N_2875,N_1729);
and U6931 (N_6931,N_2664,N_499);
xor U6932 (N_6932,N_2334,N_270);
or U6933 (N_6933,N_3656,N_3220);
and U6934 (N_6934,N_3411,N_187);
or U6935 (N_6935,N_4355,N_2830);
nor U6936 (N_6936,N_3416,N_928);
nor U6937 (N_6937,N_922,N_3279);
nor U6938 (N_6938,N_2958,N_4083);
nor U6939 (N_6939,N_1843,N_2926);
nand U6940 (N_6940,N_3646,N_2423);
and U6941 (N_6941,N_4185,N_1556);
and U6942 (N_6942,N_4091,N_3016);
xor U6943 (N_6943,N_4218,N_2864);
and U6944 (N_6944,N_3958,N_325);
and U6945 (N_6945,N_4897,N_3170);
nor U6946 (N_6946,N_1758,N_2086);
nor U6947 (N_6947,N_4959,N_1786);
and U6948 (N_6948,N_2941,N_802);
and U6949 (N_6949,N_3743,N_3464);
or U6950 (N_6950,N_3399,N_2091);
nand U6951 (N_6951,N_3756,N_485);
nand U6952 (N_6952,N_3264,N_860);
nor U6953 (N_6953,N_2206,N_993);
or U6954 (N_6954,N_2702,N_4931);
nand U6955 (N_6955,N_2976,N_4137);
or U6956 (N_6956,N_333,N_3820);
nor U6957 (N_6957,N_822,N_978);
or U6958 (N_6958,N_1071,N_1791);
and U6959 (N_6959,N_580,N_1961);
nor U6960 (N_6960,N_2516,N_4871);
nor U6961 (N_6961,N_3850,N_4675);
nand U6962 (N_6962,N_644,N_2509);
nor U6963 (N_6963,N_4652,N_3472);
nor U6964 (N_6964,N_3525,N_3293);
and U6965 (N_6965,N_586,N_1746);
xor U6966 (N_6966,N_3929,N_3408);
and U6967 (N_6967,N_2255,N_4034);
nand U6968 (N_6968,N_2669,N_3991);
or U6969 (N_6969,N_2339,N_1106);
and U6970 (N_6970,N_1109,N_1841);
nand U6971 (N_6971,N_2413,N_4670);
nor U6972 (N_6972,N_2282,N_3649);
nor U6973 (N_6973,N_1871,N_78);
or U6974 (N_6974,N_2773,N_3438);
or U6975 (N_6975,N_373,N_2525);
or U6976 (N_6976,N_2796,N_1255);
nor U6977 (N_6977,N_1736,N_1959);
nor U6978 (N_6978,N_1895,N_1338);
and U6979 (N_6979,N_1015,N_35);
nand U6980 (N_6980,N_2914,N_3595);
xnor U6981 (N_6981,N_1058,N_100);
nor U6982 (N_6982,N_1673,N_1638);
nand U6983 (N_6983,N_3870,N_2196);
nor U6984 (N_6984,N_4552,N_1428);
nand U6985 (N_6985,N_2041,N_1220);
nand U6986 (N_6986,N_2484,N_2651);
and U6987 (N_6987,N_4482,N_3675);
nand U6988 (N_6988,N_2342,N_3463);
or U6989 (N_6989,N_2768,N_794);
and U6990 (N_6990,N_3246,N_3294);
xor U6991 (N_6991,N_1723,N_718);
and U6992 (N_6992,N_1910,N_2227);
nand U6993 (N_6993,N_377,N_2866);
nand U6994 (N_6994,N_1460,N_3176);
or U6995 (N_6995,N_438,N_282);
nand U6996 (N_6996,N_2235,N_673);
and U6997 (N_6997,N_4369,N_4573);
nor U6998 (N_6998,N_3592,N_2508);
or U6999 (N_6999,N_1466,N_4472);
nor U7000 (N_7000,N_4273,N_4768);
or U7001 (N_7001,N_2448,N_1730);
nand U7002 (N_7002,N_2729,N_2272);
or U7003 (N_7003,N_1160,N_4339);
or U7004 (N_7004,N_3141,N_1088);
nand U7005 (N_7005,N_1994,N_4440);
and U7006 (N_7006,N_598,N_2785);
nor U7007 (N_7007,N_864,N_1368);
or U7008 (N_7008,N_1231,N_1834);
and U7009 (N_7009,N_2133,N_3397);
xor U7010 (N_7010,N_2944,N_3704);
and U7011 (N_7011,N_3647,N_1452);
nand U7012 (N_7012,N_1762,N_1119);
nand U7013 (N_7013,N_648,N_1409);
or U7014 (N_7014,N_3044,N_2983);
nor U7015 (N_7015,N_4213,N_203);
nor U7016 (N_7016,N_1127,N_3836);
and U7017 (N_7017,N_988,N_366);
nand U7018 (N_7018,N_2102,N_2441);
and U7019 (N_7019,N_454,N_714);
nand U7020 (N_7020,N_56,N_1558);
and U7021 (N_7021,N_2560,N_4693);
xor U7022 (N_7022,N_2653,N_1122);
and U7023 (N_7023,N_3666,N_3046);
nor U7024 (N_7024,N_119,N_4074);
nor U7025 (N_7025,N_3529,N_4695);
and U7026 (N_7026,N_909,N_1239);
or U7027 (N_7027,N_1832,N_4557);
nor U7028 (N_7028,N_3427,N_3360);
nand U7029 (N_7029,N_1126,N_4158);
nand U7030 (N_7030,N_3199,N_2993);
and U7031 (N_7031,N_80,N_1757);
xor U7032 (N_7032,N_2319,N_1229);
or U7033 (N_7033,N_1476,N_2537);
nor U7034 (N_7034,N_3812,N_3142);
or U7035 (N_7035,N_4685,N_1971);
xor U7036 (N_7036,N_2705,N_4413);
xnor U7037 (N_7037,N_2288,N_523);
nand U7038 (N_7038,N_1108,N_4263);
nor U7039 (N_7039,N_876,N_3124);
xor U7040 (N_7040,N_2767,N_4743);
and U7041 (N_7041,N_2428,N_809);
or U7042 (N_7042,N_2267,N_3174);
nor U7043 (N_7043,N_1610,N_4785);
or U7044 (N_7044,N_1825,N_458);
nand U7045 (N_7045,N_2013,N_701);
nor U7046 (N_7046,N_3278,N_343);
nand U7047 (N_7047,N_1092,N_4937);
nand U7048 (N_7048,N_1568,N_782);
nor U7049 (N_7049,N_3676,N_3696);
nand U7050 (N_7050,N_3773,N_1870);
nor U7051 (N_7051,N_2855,N_2366);
or U7052 (N_7052,N_3512,N_4534);
nor U7053 (N_7053,N_3035,N_4327);
nor U7054 (N_7054,N_4455,N_4408);
or U7055 (N_7055,N_153,N_2540);
or U7056 (N_7056,N_4822,N_1896);
nand U7057 (N_7057,N_2857,N_3640);
nand U7058 (N_7058,N_3530,N_2469);
and U7059 (N_7059,N_2974,N_1208);
or U7060 (N_7060,N_2142,N_2841);
nand U7061 (N_7061,N_2046,N_3601);
or U7062 (N_7062,N_3032,N_596);
nand U7063 (N_7063,N_3350,N_1189);
or U7064 (N_7064,N_4986,N_927);
or U7065 (N_7065,N_3541,N_1657);
or U7066 (N_7066,N_3251,N_2549);
or U7067 (N_7067,N_2967,N_3282);
nor U7068 (N_7068,N_4965,N_3466);
nand U7069 (N_7069,N_2887,N_2786);
nor U7070 (N_7070,N_998,N_3724);
and U7071 (N_7071,N_1993,N_4491);
xnor U7072 (N_7072,N_4317,N_583);
nand U7073 (N_7073,N_4315,N_1936);
xnor U7074 (N_7074,N_3519,N_3083);
nand U7075 (N_7075,N_4377,N_1667);
and U7076 (N_7076,N_167,N_4496);
xnor U7077 (N_7077,N_51,N_1517);
nand U7078 (N_7078,N_3521,N_4674);
nor U7079 (N_7079,N_4945,N_1381);
nand U7080 (N_7080,N_143,N_729);
and U7081 (N_7081,N_739,N_630);
and U7082 (N_7082,N_4671,N_4285);
nor U7083 (N_7083,N_2894,N_94);
nor U7084 (N_7084,N_4540,N_177);
or U7085 (N_7085,N_1676,N_3001);
and U7086 (N_7086,N_2080,N_4981);
xnor U7087 (N_7087,N_4974,N_4488);
nand U7088 (N_7088,N_1642,N_400);
and U7089 (N_7089,N_1771,N_4712);
or U7090 (N_7090,N_4028,N_892);
xor U7091 (N_7091,N_3736,N_4365);
and U7092 (N_7092,N_3303,N_3328);
or U7093 (N_7093,N_3799,N_1500);
nor U7094 (N_7094,N_563,N_4653);
nand U7095 (N_7095,N_181,N_3243);
nand U7096 (N_7096,N_4148,N_3033);
and U7097 (N_7097,N_1953,N_4033);
or U7098 (N_7098,N_649,N_214);
nand U7099 (N_7099,N_42,N_3166);
or U7100 (N_7100,N_4103,N_3625);
and U7101 (N_7101,N_704,N_1111);
xnor U7102 (N_7102,N_2321,N_33);
and U7103 (N_7103,N_2122,N_2515);
nor U7104 (N_7104,N_265,N_4251);
and U7105 (N_7105,N_4330,N_2384);
nor U7106 (N_7106,N_2216,N_1693);
and U7107 (N_7107,N_4733,N_268);
or U7108 (N_7108,N_2889,N_1050);
and U7109 (N_7109,N_3945,N_3482);
xor U7110 (N_7110,N_4838,N_468);
or U7111 (N_7111,N_854,N_3995);
and U7112 (N_7112,N_2063,N_154);
nand U7113 (N_7113,N_3801,N_4794);
and U7114 (N_7114,N_1777,N_1937);
or U7115 (N_7115,N_2440,N_2320);
nor U7116 (N_7116,N_116,N_3451);
xor U7117 (N_7117,N_2534,N_4006);
or U7118 (N_7118,N_4188,N_4856);
nor U7119 (N_7119,N_3997,N_1482);
xor U7120 (N_7120,N_4062,N_2635);
xor U7121 (N_7121,N_4417,N_1659);
nand U7122 (N_7122,N_2032,N_2054);
or U7123 (N_7123,N_1717,N_1601);
nand U7124 (N_7124,N_2546,N_3230);
nor U7125 (N_7125,N_1259,N_2861);
nand U7126 (N_7126,N_806,N_3483);
nand U7127 (N_7127,N_76,N_1951);
or U7128 (N_7128,N_2487,N_510);
nor U7129 (N_7129,N_769,N_2607);
or U7130 (N_7130,N_2278,N_731);
nand U7131 (N_7131,N_3099,N_4098);
xnor U7132 (N_7132,N_59,N_4895);
and U7133 (N_7133,N_2536,N_1668);
or U7134 (N_7134,N_4564,N_1969);
xor U7135 (N_7135,N_1599,N_4481);
nand U7136 (N_7136,N_1237,N_2981);
and U7137 (N_7137,N_4910,N_3922);
or U7138 (N_7138,N_4126,N_4904);
and U7139 (N_7139,N_4634,N_401);
or U7140 (N_7140,N_3761,N_4073);
nor U7141 (N_7141,N_4220,N_4649);
and U7142 (N_7142,N_3690,N_3245);
nor U7143 (N_7143,N_1582,N_2295);
nor U7144 (N_7144,N_3973,N_1530);
nor U7145 (N_7145,N_4606,N_2250);
and U7146 (N_7146,N_346,N_1438);
xor U7147 (N_7147,N_3677,N_3834);
nor U7148 (N_7148,N_89,N_1105);
nor U7149 (N_7149,N_74,N_1196);
nand U7150 (N_7150,N_2388,N_418);
xnor U7151 (N_7151,N_872,N_3247);
nand U7152 (N_7152,N_1218,N_4276);
nor U7153 (N_7153,N_4823,N_2064);
xnor U7154 (N_7154,N_2073,N_2472);
nand U7155 (N_7155,N_2556,N_3611);
and U7156 (N_7156,N_4268,N_869);
nand U7157 (N_7157,N_890,N_3815);
or U7158 (N_7158,N_4610,N_1062);
nor U7159 (N_7159,N_804,N_3952);
xnor U7160 (N_7160,N_1984,N_2177);
or U7161 (N_7161,N_3461,N_1923);
and U7162 (N_7162,N_2259,N_1082);
nand U7163 (N_7163,N_1917,N_3008);
and U7164 (N_7164,N_900,N_1284);
nand U7165 (N_7165,N_2375,N_360);
nor U7166 (N_7166,N_3444,N_4484);
and U7167 (N_7167,N_3964,N_1416);
nand U7168 (N_7168,N_2986,N_4681);
nand U7169 (N_7169,N_3996,N_2989);
nor U7170 (N_7170,N_660,N_429);
xor U7171 (N_7171,N_2496,N_4587);
nand U7172 (N_7172,N_1141,N_3457);
nor U7173 (N_7173,N_1858,N_2678);
and U7174 (N_7174,N_2137,N_4433);
xnor U7175 (N_7175,N_3565,N_1073);
nor U7176 (N_7176,N_3405,N_4310);
and U7177 (N_7177,N_3410,N_3078);
and U7178 (N_7178,N_796,N_1129);
and U7179 (N_7179,N_2471,N_2251);
nor U7180 (N_7180,N_2580,N_1567);
and U7181 (N_7181,N_1637,N_3968);
or U7182 (N_7182,N_976,N_3292);
nor U7183 (N_7183,N_4000,N_417);
or U7184 (N_7184,N_1773,N_1604);
nor U7185 (N_7185,N_4760,N_4391);
nor U7186 (N_7186,N_4934,N_3556);
nand U7187 (N_7187,N_1199,N_3664);
and U7188 (N_7188,N_624,N_566);
and U7189 (N_7189,N_1053,N_1124);
nor U7190 (N_7190,N_289,N_3048);
nand U7191 (N_7191,N_3477,N_2939);
and U7192 (N_7192,N_246,N_4603);
nor U7193 (N_7193,N_3165,N_3013);
nand U7194 (N_7194,N_748,N_1947);
or U7195 (N_7195,N_1520,N_759);
or U7196 (N_7196,N_1856,N_4046);
nor U7197 (N_7197,N_4960,N_933);
and U7198 (N_7198,N_4661,N_3657);
or U7199 (N_7199,N_2311,N_2464);
nand U7200 (N_7200,N_2078,N_457);
and U7201 (N_7201,N_560,N_3937);
and U7202 (N_7202,N_140,N_3653);
nor U7203 (N_7203,N_749,N_3883);
or U7204 (N_7204,N_2685,N_2507);
and U7205 (N_7205,N_810,N_4902);
nand U7206 (N_7206,N_2242,N_4197);
xor U7207 (N_7207,N_4940,N_3481);
or U7208 (N_7208,N_3554,N_2710);
and U7209 (N_7209,N_4065,N_1636);
and U7210 (N_7210,N_1527,N_3777);
and U7211 (N_7211,N_4521,N_2600);
and U7212 (N_7212,N_358,N_3925);
nand U7213 (N_7213,N_4507,N_4990);
and U7214 (N_7214,N_4775,N_2610);
nand U7215 (N_7215,N_2493,N_3233);
nor U7216 (N_7216,N_4264,N_1542);
xor U7217 (N_7217,N_3248,N_4296);
and U7218 (N_7218,N_2996,N_4221);
and U7219 (N_7219,N_352,N_2092);
or U7220 (N_7220,N_785,N_2236);
or U7221 (N_7221,N_845,N_124);
and U7222 (N_7222,N_2253,N_2113);
or U7223 (N_7223,N_4281,N_1028);
or U7224 (N_7224,N_3424,N_4853);
and U7225 (N_7225,N_1970,N_2778);
and U7226 (N_7226,N_3767,N_3721);
nand U7227 (N_7227,N_3641,N_330);
nor U7228 (N_7228,N_1740,N_4161);
xor U7229 (N_7229,N_2690,N_3442);
xnor U7230 (N_7230,N_1290,N_1307);
nor U7231 (N_7231,N_1543,N_431);
and U7232 (N_7232,N_3835,N_3662);
nand U7233 (N_7233,N_2343,N_3173);
nor U7234 (N_7234,N_1426,N_2056);
and U7235 (N_7235,N_1692,N_555);
or U7236 (N_7236,N_4181,N_1885);
or U7237 (N_7237,N_1617,N_1243);
nor U7238 (N_7238,N_3710,N_24);
and U7239 (N_7239,N_4834,N_3402);
or U7240 (N_7240,N_2162,N_983);
nand U7241 (N_7241,N_452,N_3926);
and U7242 (N_7242,N_913,N_2542);
or U7243 (N_7243,N_478,N_2642);
xor U7244 (N_7244,N_3689,N_3550);
xnor U7245 (N_7245,N_3151,N_3103);
and U7246 (N_7246,N_2886,N_1388);
and U7247 (N_7247,N_3257,N_605);
or U7248 (N_7248,N_397,N_1826);
or U7249 (N_7249,N_386,N_2799);
or U7250 (N_7250,N_3539,N_217);
nor U7251 (N_7251,N_2909,N_562);
or U7252 (N_7252,N_1352,N_534);
xnor U7253 (N_7253,N_2274,N_1713);
nand U7254 (N_7254,N_1448,N_2294);
and U7255 (N_7255,N_2368,N_2389);
nand U7256 (N_7256,N_172,N_2501);
nand U7257 (N_7257,N_4194,N_476);
or U7258 (N_7258,N_21,N_1949);
nand U7259 (N_7259,N_2407,N_1823);
xor U7260 (N_7260,N_3361,N_4135);
and U7261 (N_7261,N_4236,N_565);
xnor U7262 (N_7262,N_3598,N_4673);
or U7263 (N_7263,N_4936,N_1059);
or U7264 (N_7264,N_1665,N_1817);
nand U7265 (N_7265,N_3039,N_2936);
nor U7266 (N_7266,N_1612,N_4832);
or U7267 (N_7267,N_1677,N_643);
nor U7268 (N_7268,N_3054,N_1867);
or U7269 (N_7269,N_984,N_542);
and U7270 (N_7270,N_4930,N_3317);
or U7271 (N_7271,N_3896,N_958);
nor U7272 (N_7272,N_3518,N_3931);
nand U7273 (N_7273,N_4187,N_839);
and U7274 (N_7274,N_3075,N_112);
nand U7275 (N_7275,N_708,N_2324);
and U7276 (N_7276,N_4781,N_2378);
nand U7277 (N_7277,N_298,N_4527);
and U7278 (N_7278,N_4245,N_1987);
or U7279 (N_7279,N_4242,N_2439);
xnor U7280 (N_7280,N_3330,N_4140);
or U7281 (N_7281,N_1014,N_4517);
nand U7282 (N_7282,N_633,N_4084);
or U7283 (N_7283,N_168,N_584);
nor U7284 (N_7284,N_276,N_1404);
or U7285 (N_7285,N_4689,N_3309);
or U7286 (N_7286,N_2943,N_1006);
or U7287 (N_7287,N_1042,N_3975);
xor U7288 (N_7288,N_3071,N_820);
and U7289 (N_7289,N_799,N_1475);
and U7290 (N_7290,N_65,N_4346);
nor U7291 (N_7291,N_1869,N_1456);
nor U7292 (N_7292,N_3819,N_949);
or U7293 (N_7293,N_3549,N_4498);
and U7294 (N_7294,N_4441,N_4657);
nor U7295 (N_7295,N_3536,N_2901);
nand U7296 (N_7296,N_4454,N_477);
and U7297 (N_7297,N_1747,N_647);
xnor U7298 (N_7298,N_1565,N_4196);
and U7299 (N_7299,N_1929,N_3751);
nor U7300 (N_7300,N_3522,N_4463);
nor U7301 (N_7301,N_2863,N_2638);
or U7302 (N_7302,N_2143,N_1725);
and U7303 (N_7303,N_1155,N_4394);
nor U7304 (N_7304,N_762,N_1700);
nor U7305 (N_7305,N_1884,N_2214);
nand U7306 (N_7306,N_3560,N_1688);
or U7307 (N_7307,N_3116,N_3669);
or U7308 (N_7308,N_733,N_4492);
nand U7309 (N_7309,N_2870,N_4132);
or U7310 (N_7310,N_3097,N_4210);
nor U7311 (N_7311,N_445,N_209);
nand U7312 (N_7312,N_149,N_3545);
xnor U7313 (N_7313,N_3514,N_3908);
or U7314 (N_7314,N_4237,N_2990);
or U7315 (N_7315,N_4129,N_22);
nand U7316 (N_7316,N_3332,N_4134);
or U7317 (N_7317,N_1576,N_2229);
xor U7318 (N_7318,N_3652,N_4803);
or U7319 (N_7319,N_1900,N_4280);
xor U7320 (N_7320,N_1095,N_3501);
xor U7321 (N_7321,N_2104,N_3714);
or U7322 (N_7322,N_1286,N_1571);
and U7323 (N_7323,N_3930,N_2065);
xor U7324 (N_7324,N_2169,N_4149);
nand U7325 (N_7325,N_1743,N_2105);
nand U7326 (N_7326,N_2877,N_4200);
nor U7327 (N_7327,N_2682,N_3548);
and U7328 (N_7328,N_2035,N_1839);
and U7329 (N_7329,N_4836,N_3517);
and U7330 (N_7330,N_4375,N_2030);
and U7331 (N_7331,N_4348,N_1967);
nor U7332 (N_7332,N_1760,N_2752);
nand U7333 (N_7333,N_4819,N_3999);
nor U7334 (N_7334,N_686,N_735);
or U7335 (N_7335,N_4551,N_2374);
xor U7336 (N_7336,N_3073,N_4470);
nand U7337 (N_7337,N_4259,N_533);
nand U7338 (N_7338,N_3322,N_1447);
nor U7339 (N_7339,N_3242,N_3672);
and U7340 (N_7340,N_2935,N_2316);
nand U7341 (N_7341,N_3838,N_1975);
xor U7342 (N_7342,N_1778,N_967);
and U7343 (N_7343,N_3374,N_4400);
nor U7344 (N_7344,N_905,N_4762);
and U7345 (N_7345,N_1353,N_3435);
nand U7346 (N_7346,N_1631,N_4423);
and U7347 (N_7347,N_1,N_929);
nor U7348 (N_7348,N_3304,N_669);
and U7349 (N_7349,N_1715,N_3498);
nor U7350 (N_7350,N_4038,N_4739);
nor U7351 (N_7351,N_3362,N_166);
and U7352 (N_7352,N_3057,N_4544);
and U7353 (N_7353,N_3737,N_4198);
nor U7354 (N_7354,N_4191,N_3024);
nand U7355 (N_7355,N_1785,N_1592);
xnor U7356 (N_7356,N_3813,N_1833);
nand U7357 (N_7357,N_2356,N_2017);
and U7358 (N_7358,N_1942,N_1367);
or U7359 (N_7359,N_3338,N_4193);
or U7360 (N_7360,N_2804,N_2971);
nor U7361 (N_7361,N_4825,N_2414);
nor U7362 (N_7362,N_4641,N_4687);
or U7363 (N_7363,N_375,N_4182);
or U7364 (N_7364,N_4845,N_3306);
and U7365 (N_7365,N_2984,N_4332);
nand U7366 (N_7366,N_3041,N_4305);
nand U7367 (N_7367,N_61,N_3422);
nand U7368 (N_7368,N_4088,N_3811);
and U7369 (N_7369,N_3289,N_2208);
nand U7370 (N_7370,N_4979,N_3090);
or U7371 (N_7371,N_2633,N_1041);
nor U7372 (N_7372,N_1983,N_385);
or U7373 (N_7373,N_3726,N_3207);
nor U7374 (N_7374,N_1780,N_3285);
or U7375 (N_7375,N_3086,N_3965);
or U7376 (N_7376,N_1150,N_491);
and U7377 (N_7377,N_1422,N_801);
nor U7378 (N_7378,N_2619,N_4483);
nor U7379 (N_7379,N_2948,N_2593);
or U7380 (N_7380,N_4680,N_1684);
xor U7381 (N_7381,N_3577,N_936);
or U7382 (N_7382,N_781,N_2784);
nand U7383 (N_7383,N_3824,N_4967);
or U7384 (N_7384,N_1190,N_4817);
and U7385 (N_7385,N_3189,N_2410);
and U7386 (N_7386,N_1451,N_873);
or U7387 (N_7387,N_2953,N_3782);
or U7388 (N_7388,N_1238,N_1728);
nand U7389 (N_7389,N_2204,N_4939);
or U7390 (N_7390,N_2596,N_3856);
or U7391 (N_7391,N_2333,N_1013);
nand U7392 (N_7392,N_3719,N_843);
and U7393 (N_7393,N_951,N_2885);
and U7394 (N_7394,N_252,N_2980);
nand U7395 (N_7395,N_4021,N_4881);
nor U7396 (N_7396,N_4636,N_3146);
nand U7397 (N_7397,N_2691,N_1532);
nor U7398 (N_7398,N_2649,N_4275);
nand U7399 (N_7399,N_2816,N_3154);
nand U7400 (N_7400,N_240,N_3055);
or U7401 (N_7401,N_52,N_1554);
or U7402 (N_7402,N_3562,N_2427);
xor U7403 (N_7403,N_3772,N_713);
and U7404 (N_7404,N_72,N_3739);
or U7405 (N_7405,N_3358,N_4955);
nor U7406 (N_7406,N_4626,N_150);
and U7407 (N_7407,N_4971,N_2603);
and U7408 (N_7408,N_470,N_1710);
and U7409 (N_7409,N_3373,N_1585);
nand U7410 (N_7410,N_4609,N_1930);
nand U7411 (N_7411,N_2028,N_3668);
nand U7412 (N_7412,N_442,N_4468);
nor U7413 (N_7413,N_2686,N_223);
xnor U7414 (N_7414,N_3722,N_3727);
or U7415 (N_7415,N_2416,N_828);
or U7416 (N_7416,N_3150,N_3222);
xnor U7417 (N_7417,N_2461,N_420);
nand U7418 (N_7418,N_567,N_1698);
nand U7419 (N_7419,N_2589,N_2457);
nor U7420 (N_7420,N_376,N_2657);
nand U7421 (N_7421,N_4704,N_1061);
nor U7422 (N_7422,N_548,N_3610);
nand U7423 (N_7423,N_2171,N_1790);
nand U7424 (N_7424,N_4466,N_4288);
xor U7425 (N_7425,N_2838,N_4300);
nand U7426 (N_7426,N_4586,N_2435);
or U7427 (N_7427,N_513,N_3619);
and U7428 (N_7428,N_1415,N_3470);
and U7429 (N_7429,N_1097,N_3316);
and U7430 (N_7430,N_3249,N_2188);
and U7431 (N_7431,N_3878,N_1789);
nor U7432 (N_7432,N_4035,N_2383);
or U7433 (N_7433,N_1055,N_1331);
and U7434 (N_7434,N_2862,N_2466);
nor U7435 (N_7435,N_3406,N_4356);
nor U7436 (N_7436,N_180,N_4713);
and U7437 (N_7437,N_260,N_790);
or U7438 (N_7438,N_1107,N_482);
and U7439 (N_7439,N_1362,N_95);
or U7440 (N_7440,N_1261,N_3632);
nor U7441 (N_7441,N_1652,N_4235);
and U7442 (N_7442,N_296,N_2426);
or U7443 (N_7443,N_1519,N_3941);
nand U7444 (N_7444,N_92,N_1022);
nand U7445 (N_7445,N_3485,N_889);
or U7446 (N_7446,N_2391,N_3881);
nor U7447 (N_7447,N_788,N_3712);
nand U7448 (N_7448,N_1609,N_2258);
or U7449 (N_7449,N_412,N_4393);
nand U7450 (N_7450,N_2518,N_2310);
or U7451 (N_7451,N_27,N_3691);
nand U7452 (N_7452,N_3135,N_1271);
nor U7453 (N_7453,N_3206,N_3313);
nor U7454 (N_7454,N_1117,N_4069);
and U7455 (N_7455,N_4612,N_371);
nor U7456 (N_7456,N_3042,N_3732);
and U7457 (N_7457,N_964,N_659);
nand U7458 (N_7458,N_91,N_1901);
nor U7459 (N_7459,N_3302,N_2821);
nor U7460 (N_7460,N_1954,N_1926);
nand U7461 (N_7461,N_3113,N_1423);
nor U7462 (N_7462,N_4449,N_2299);
nand U7463 (N_7463,N_1524,N_1397);
and U7464 (N_7464,N_1132,N_1487);
or U7465 (N_7465,N_2273,N_3372);
nor U7466 (N_7466,N_3445,N_3823);
nor U7467 (N_7467,N_722,N_1172);
nor U7468 (N_7468,N_1483,N_4363);
and U7469 (N_7469,N_4541,N_996);
and U7470 (N_7470,N_2755,N_1488);
and U7471 (N_7471,N_3880,N_3542);
nand U7472 (N_7472,N_2025,N_1325);
and U7473 (N_7473,N_727,N_3428);
xnor U7474 (N_7474,N_2447,N_1310);
and U7475 (N_7475,N_2071,N_4683);
and U7476 (N_7476,N_3621,N_4535);
nor U7477 (N_7477,N_1304,N_3077);
and U7478 (N_7478,N_1077,N_4318);
nand U7479 (N_7479,N_3311,N_866);
nand U7480 (N_7480,N_4057,N_617);
nor U7481 (N_7481,N_3841,N_4581);
and U7482 (N_7482,N_4831,N_3644);
nor U7483 (N_7483,N_2085,N_1932);
or U7484 (N_7484,N_1001,N_1330);
or U7485 (N_7485,N_4846,N_2438);
nor U7486 (N_7486,N_4438,N_3191);
or U7487 (N_7487,N_4709,N_2132);
and U7488 (N_7488,N_370,N_1384);
xor U7489 (N_7489,N_4414,N_3388);
nand U7490 (N_7490,N_1265,N_1031);
or U7491 (N_7491,N_1431,N_2254);
or U7492 (N_7492,N_3594,N_4839);
and U7493 (N_7493,N_2020,N_1973);
nand U7494 (N_7494,N_1632,N_3149);
nand U7495 (N_7495,N_4651,N_3866);
xor U7496 (N_7496,N_4037,N_4023);
and U7497 (N_7497,N_3909,N_4278);
nand U7498 (N_7498,N_3112,N_4659);
xor U7499 (N_7499,N_4942,N_4926);
nand U7500 (N_7500,N_1969,N_4004);
and U7501 (N_7501,N_203,N_4574);
and U7502 (N_7502,N_8,N_4575);
and U7503 (N_7503,N_2748,N_4921);
nand U7504 (N_7504,N_2465,N_3914);
nor U7505 (N_7505,N_1026,N_2435);
and U7506 (N_7506,N_4956,N_1665);
nand U7507 (N_7507,N_2345,N_2038);
nand U7508 (N_7508,N_1249,N_4621);
or U7509 (N_7509,N_2449,N_4660);
xnor U7510 (N_7510,N_1190,N_1712);
and U7511 (N_7511,N_4106,N_1088);
xnor U7512 (N_7512,N_3950,N_3149);
nor U7513 (N_7513,N_4367,N_4272);
or U7514 (N_7514,N_3663,N_2075);
or U7515 (N_7515,N_1098,N_366);
nor U7516 (N_7516,N_3602,N_4860);
or U7517 (N_7517,N_2018,N_1098);
nand U7518 (N_7518,N_325,N_4082);
nand U7519 (N_7519,N_1028,N_4378);
nand U7520 (N_7520,N_2395,N_1220);
and U7521 (N_7521,N_2253,N_4736);
or U7522 (N_7522,N_4734,N_1704);
or U7523 (N_7523,N_3931,N_4894);
xor U7524 (N_7524,N_201,N_3827);
or U7525 (N_7525,N_2257,N_933);
nand U7526 (N_7526,N_1064,N_4666);
or U7527 (N_7527,N_664,N_73);
xor U7528 (N_7528,N_1362,N_1880);
nor U7529 (N_7529,N_3366,N_3688);
and U7530 (N_7530,N_4556,N_1220);
and U7531 (N_7531,N_2383,N_3284);
nand U7532 (N_7532,N_1199,N_84);
and U7533 (N_7533,N_3967,N_2835);
nor U7534 (N_7534,N_4592,N_1993);
nor U7535 (N_7535,N_2950,N_2176);
and U7536 (N_7536,N_4284,N_2693);
nor U7537 (N_7537,N_963,N_2041);
and U7538 (N_7538,N_4646,N_590);
or U7539 (N_7539,N_437,N_4572);
and U7540 (N_7540,N_1532,N_949);
and U7541 (N_7541,N_120,N_1926);
nor U7542 (N_7542,N_2722,N_2702);
nor U7543 (N_7543,N_2301,N_2368);
xnor U7544 (N_7544,N_2923,N_3689);
nor U7545 (N_7545,N_3812,N_3325);
and U7546 (N_7546,N_1128,N_147);
nand U7547 (N_7547,N_3442,N_4528);
nor U7548 (N_7548,N_189,N_1551);
or U7549 (N_7549,N_2757,N_1912);
nor U7550 (N_7550,N_1,N_1629);
nor U7551 (N_7551,N_1481,N_1193);
nor U7552 (N_7552,N_3074,N_610);
xnor U7553 (N_7553,N_2614,N_625);
nand U7554 (N_7554,N_277,N_3983);
nor U7555 (N_7555,N_4621,N_2900);
and U7556 (N_7556,N_623,N_249);
nor U7557 (N_7557,N_2342,N_1160);
nand U7558 (N_7558,N_3929,N_3411);
nand U7559 (N_7559,N_4818,N_1833);
nor U7560 (N_7560,N_627,N_3358);
or U7561 (N_7561,N_2573,N_534);
or U7562 (N_7562,N_2774,N_1512);
or U7563 (N_7563,N_518,N_957);
or U7564 (N_7564,N_998,N_4509);
nand U7565 (N_7565,N_4662,N_3487);
nand U7566 (N_7566,N_1090,N_130);
nand U7567 (N_7567,N_4896,N_3610);
and U7568 (N_7568,N_447,N_538);
and U7569 (N_7569,N_659,N_1590);
or U7570 (N_7570,N_1627,N_4828);
nand U7571 (N_7571,N_526,N_2444);
nor U7572 (N_7572,N_2319,N_628);
or U7573 (N_7573,N_556,N_2030);
or U7574 (N_7574,N_4180,N_2892);
nand U7575 (N_7575,N_4376,N_81);
and U7576 (N_7576,N_279,N_1922);
nor U7577 (N_7577,N_2801,N_1759);
nor U7578 (N_7578,N_4411,N_1947);
nand U7579 (N_7579,N_1234,N_4540);
nand U7580 (N_7580,N_3313,N_962);
or U7581 (N_7581,N_2516,N_1713);
nand U7582 (N_7582,N_2639,N_3938);
nand U7583 (N_7583,N_166,N_4332);
nand U7584 (N_7584,N_4437,N_1663);
or U7585 (N_7585,N_1965,N_3849);
nand U7586 (N_7586,N_4215,N_2225);
and U7587 (N_7587,N_4036,N_398);
nor U7588 (N_7588,N_4213,N_1633);
or U7589 (N_7589,N_2774,N_2755);
nand U7590 (N_7590,N_747,N_52);
nand U7591 (N_7591,N_682,N_4784);
or U7592 (N_7592,N_3839,N_4235);
nor U7593 (N_7593,N_174,N_3294);
nand U7594 (N_7594,N_1488,N_3485);
and U7595 (N_7595,N_4195,N_3643);
nand U7596 (N_7596,N_2565,N_817);
xor U7597 (N_7597,N_3460,N_80);
or U7598 (N_7598,N_3980,N_4195);
or U7599 (N_7599,N_4144,N_1040);
and U7600 (N_7600,N_785,N_1420);
nand U7601 (N_7601,N_2499,N_4337);
or U7602 (N_7602,N_2774,N_2775);
nand U7603 (N_7603,N_4493,N_3841);
xnor U7604 (N_7604,N_2488,N_3426);
xor U7605 (N_7605,N_4580,N_2515);
or U7606 (N_7606,N_548,N_2239);
or U7607 (N_7607,N_4145,N_4848);
xnor U7608 (N_7608,N_4535,N_4136);
xor U7609 (N_7609,N_2922,N_2963);
or U7610 (N_7610,N_96,N_1607);
or U7611 (N_7611,N_3156,N_3880);
nor U7612 (N_7612,N_4622,N_2449);
and U7613 (N_7613,N_4981,N_1022);
and U7614 (N_7614,N_1226,N_2764);
nor U7615 (N_7615,N_276,N_2740);
or U7616 (N_7616,N_2437,N_1459);
or U7617 (N_7617,N_2201,N_707);
nand U7618 (N_7618,N_3727,N_441);
or U7619 (N_7619,N_2978,N_1764);
or U7620 (N_7620,N_2384,N_1595);
or U7621 (N_7621,N_3805,N_4725);
and U7622 (N_7622,N_3396,N_4941);
or U7623 (N_7623,N_883,N_2531);
nand U7624 (N_7624,N_3090,N_1450);
nor U7625 (N_7625,N_1895,N_1734);
and U7626 (N_7626,N_4395,N_3080);
or U7627 (N_7627,N_3609,N_4208);
xnor U7628 (N_7628,N_1775,N_759);
nor U7629 (N_7629,N_3374,N_228);
nand U7630 (N_7630,N_2831,N_438);
nor U7631 (N_7631,N_1224,N_4831);
nand U7632 (N_7632,N_1827,N_2559);
and U7633 (N_7633,N_883,N_2046);
nor U7634 (N_7634,N_49,N_3765);
nand U7635 (N_7635,N_1593,N_3313);
nand U7636 (N_7636,N_253,N_4704);
or U7637 (N_7637,N_4652,N_1668);
nand U7638 (N_7638,N_2823,N_4408);
or U7639 (N_7639,N_4933,N_1573);
nand U7640 (N_7640,N_1191,N_868);
nand U7641 (N_7641,N_4932,N_252);
and U7642 (N_7642,N_963,N_3243);
and U7643 (N_7643,N_3489,N_4564);
and U7644 (N_7644,N_2910,N_1247);
and U7645 (N_7645,N_1867,N_3107);
and U7646 (N_7646,N_264,N_578);
nand U7647 (N_7647,N_1545,N_2883);
or U7648 (N_7648,N_3516,N_3613);
nand U7649 (N_7649,N_1592,N_149);
and U7650 (N_7650,N_4158,N_2304);
xnor U7651 (N_7651,N_1319,N_2031);
xnor U7652 (N_7652,N_602,N_2647);
nand U7653 (N_7653,N_3186,N_1031);
and U7654 (N_7654,N_4756,N_3395);
or U7655 (N_7655,N_4329,N_3783);
nand U7656 (N_7656,N_3806,N_2193);
or U7657 (N_7657,N_11,N_4387);
and U7658 (N_7658,N_116,N_1934);
and U7659 (N_7659,N_780,N_4652);
nand U7660 (N_7660,N_3909,N_1420);
nand U7661 (N_7661,N_4414,N_1840);
nor U7662 (N_7662,N_1363,N_4774);
and U7663 (N_7663,N_511,N_3999);
nand U7664 (N_7664,N_2809,N_2277);
nand U7665 (N_7665,N_840,N_1905);
xor U7666 (N_7666,N_1694,N_1682);
and U7667 (N_7667,N_3554,N_1975);
or U7668 (N_7668,N_1179,N_4226);
nand U7669 (N_7669,N_4628,N_3817);
and U7670 (N_7670,N_1489,N_781);
and U7671 (N_7671,N_369,N_871);
nor U7672 (N_7672,N_3484,N_4901);
nor U7673 (N_7673,N_1122,N_2876);
nand U7674 (N_7674,N_2103,N_2848);
nand U7675 (N_7675,N_1680,N_839);
nand U7676 (N_7676,N_891,N_47);
or U7677 (N_7677,N_4486,N_1688);
and U7678 (N_7678,N_323,N_1716);
or U7679 (N_7679,N_3468,N_904);
nand U7680 (N_7680,N_3128,N_3053);
or U7681 (N_7681,N_1815,N_2698);
or U7682 (N_7682,N_3560,N_2617);
nor U7683 (N_7683,N_1095,N_2592);
and U7684 (N_7684,N_2105,N_4121);
and U7685 (N_7685,N_4956,N_1552);
and U7686 (N_7686,N_65,N_4973);
xnor U7687 (N_7687,N_1002,N_1759);
nor U7688 (N_7688,N_4751,N_4766);
and U7689 (N_7689,N_3570,N_65);
or U7690 (N_7690,N_2678,N_840);
and U7691 (N_7691,N_1847,N_2556);
nand U7692 (N_7692,N_4645,N_4976);
nand U7693 (N_7693,N_1860,N_382);
and U7694 (N_7694,N_1320,N_1960);
nor U7695 (N_7695,N_4158,N_1716);
nand U7696 (N_7696,N_98,N_283);
or U7697 (N_7697,N_1221,N_2737);
or U7698 (N_7698,N_4439,N_3652);
or U7699 (N_7699,N_798,N_859);
xor U7700 (N_7700,N_522,N_186);
xnor U7701 (N_7701,N_4548,N_1526);
or U7702 (N_7702,N_2652,N_1474);
nor U7703 (N_7703,N_1364,N_401);
and U7704 (N_7704,N_3072,N_2117);
nand U7705 (N_7705,N_4599,N_1133);
nor U7706 (N_7706,N_810,N_3037);
nor U7707 (N_7707,N_3337,N_2859);
nor U7708 (N_7708,N_3454,N_1040);
or U7709 (N_7709,N_3042,N_451);
and U7710 (N_7710,N_2240,N_3864);
and U7711 (N_7711,N_2924,N_2394);
nand U7712 (N_7712,N_3739,N_2619);
nand U7713 (N_7713,N_690,N_1677);
nand U7714 (N_7714,N_2675,N_2781);
nor U7715 (N_7715,N_3256,N_2590);
xor U7716 (N_7716,N_3582,N_2001);
nand U7717 (N_7717,N_2719,N_3116);
nand U7718 (N_7718,N_1915,N_1117);
and U7719 (N_7719,N_2791,N_889);
or U7720 (N_7720,N_4963,N_4045);
and U7721 (N_7721,N_2830,N_2184);
and U7722 (N_7722,N_1064,N_297);
xor U7723 (N_7723,N_4391,N_1697);
xor U7724 (N_7724,N_436,N_4153);
nor U7725 (N_7725,N_1931,N_878);
and U7726 (N_7726,N_904,N_3156);
or U7727 (N_7727,N_2617,N_3940);
nor U7728 (N_7728,N_1334,N_3390);
and U7729 (N_7729,N_376,N_3304);
nor U7730 (N_7730,N_4822,N_2886);
nor U7731 (N_7731,N_223,N_3194);
nand U7732 (N_7732,N_2019,N_3191);
or U7733 (N_7733,N_1225,N_3528);
nand U7734 (N_7734,N_1627,N_1233);
nand U7735 (N_7735,N_3240,N_2540);
nor U7736 (N_7736,N_480,N_1075);
or U7737 (N_7737,N_2215,N_3141);
and U7738 (N_7738,N_1769,N_1485);
or U7739 (N_7739,N_3466,N_484);
nand U7740 (N_7740,N_2143,N_4594);
nor U7741 (N_7741,N_2202,N_3380);
and U7742 (N_7742,N_2253,N_3705);
and U7743 (N_7743,N_2479,N_4663);
xor U7744 (N_7744,N_806,N_1894);
and U7745 (N_7745,N_4967,N_4171);
and U7746 (N_7746,N_4447,N_4243);
nand U7747 (N_7747,N_4861,N_3037);
nor U7748 (N_7748,N_2717,N_4987);
nor U7749 (N_7749,N_1332,N_313);
or U7750 (N_7750,N_1591,N_2578);
nand U7751 (N_7751,N_3757,N_3389);
nor U7752 (N_7752,N_1344,N_1495);
or U7753 (N_7753,N_3523,N_209);
xor U7754 (N_7754,N_2266,N_1780);
xnor U7755 (N_7755,N_1322,N_1391);
or U7756 (N_7756,N_1881,N_3455);
or U7757 (N_7757,N_1008,N_4865);
nor U7758 (N_7758,N_1728,N_2436);
nand U7759 (N_7759,N_2276,N_3748);
nand U7760 (N_7760,N_1971,N_2857);
xnor U7761 (N_7761,N_2080,N_668);
and U7762 (N_7762,N_1836,N_2873);
nand U7763 (N_7763,N_314,N_3643);
xor U7764 (N_7764,N_95,N_4454);
or U7765 (N_7765,N_1000,N_4097);
nand U7766 (N_7766,N_1826,N_3469);
nand U7767 (N_7767,N_1262,N_4142);
xnor U7768 (N_7768,N_1637,N_4013);
nand U7769 (N_7769,N_450,N_831);
and U7770 (N_7770,N_642,N_4385);
or U7771 (N_7771,N_4876,N_4329);
nand U7772 (N_7772,N_3649,N_2997);
or U7773 (N_7773,N_1999,N_1281);
or U7774 (N_7774,N_3507,N_2632);
xnor U7775 (N_7775,N_4195,N_855);
xnor U7776 (N_7776,N_2144,N_2383);
nand U7777 (N_7777,N_3918,N_1911);
nor U7778 (N_7778,N_4996,N_4483);
xor U7779 (N_7779,N_3126,N_2674);
nand U7780 (N_7780,N_370,N_3440);
and U7781 (N_7781,N_3730,N_986);
or U7782 (N_7782,N_356,N_2150);
nand U7783 (N_7783,N_2199,N_3977);
xor U7784 (N_7784,N_1990,N_4478);
nand U7785 (N_7785,N_3502,N_2587);
nor U7786 (N_7786,N_318,N_2540);
and U7787 (N_7787,N_2632,N_3775);
nand U7788 (N_7788,N_1720,N_3676);
nand U7789 (N_7789,N_3129,N_266);
and U7790 (N_7790,N_2867,N_2558);
or U7791 (N_7791,N_635,N_3832);
nor U7792 (N_7792,N_254,N_4681);
nor U7793 (N_7793,N_1928,N_1405);
nand U7794 (N_7794,N_4148,N_3831);
xor U7795 (N_7795,N_3262,N_1820);
and U7796 (N_7796,N_2837,N_1842);
nor U7797 (N_7797,N_2591,N_3528);
nor U7798 (N_7798,N_1299,N_3110);
or U7799 (N_7799,N_645,N_3524);
and U7800 (N_7800,N_2965,N_1249);
nand U7801 (N_7801,N_1379,N_3454);
nand U7802 (N_7802,N_3537,N_254);
nor U7803 (N_7803,N_1592,N_1046);
and U7804 (N_7804,N_1338,N_1255);
and U7805 (N_7805,N_2331,N_4656);
and U7806 (N_7806,N_4334,N_2622);
nand U7807 (N_7807,N_2065,N_1029);
and U7808 (N_7808,N_4983,N_2214);
and U7809 (N_7809,N_383,N_1726);
and U7810 (N_7810,N_3346,N_86);
and U7811 (N_7811,N_602,N_653);
nor U7812 (N_7812,N_2891,N_2153);
and U7813 (N_7813,N_638,N_4689);
and U7814 (N_7814,N_4675,N_3298);
nor U7815 (N_7815,N_4359,N_4622);
or U7816 (N_7816,N_2260,N_194);
nor U7817 (N_7817,N_171,N_1045);
nor U7818 (N_7818,N_4363,N_3111);
nor U7819 (N_7819,N_2169,N_2099);
xnor U7820 (N_7820,N_919,N_2385);
nand U7821 (N_7821,N_1320,N_2230);
and U7822 (N_7822,N_4579,N_4048);
nor U7823 (N_7823,N_1404,N_111);
or U7824 (N_7824,N_1781,N_1800);
xor U7825 (N_7825,N_1456,N_3748);
nand U7826 (N_7826,N_4103,N_1715);
and U7827 (N_7827,N_2705,N_4386);
nor U7828 (N_7828,N_1190,N_4626);
xor U7829 (N_7829,N_1404,N_1256);
nand U7830 (N_7830,N_3178,N_631);
and U7831 (N_7831,N_2863,N_2363);
nand U7832 (N_7832,N_4413,N_1499);
nand U7833 (N_7833,N_2539,N_3876);
nor U7834 (N_7834,N_1128,N_1746);
nand U7835 (N_7835,N_3248,N_4604);
and U7836 (N_7836,N_2800,N_3205);
and U7837 (N_7837,N_2173,N_101);
and U7838 (N_7838,N_2201,N_3446);
nand U7839 (N_7839,N_3873,N_686);
xnor U7840 (N_7840,N_487,N_2691);
xnor U7841 (N_7841,N_4322,N_2482);
or U7842 (N_7842,N_2374,N_2107);
and U7843 (N_7843,N_572,N_3040);
or U7844 (N_7844,N_3116,N_3825);
nor U7845 (N_7845,N_4644,N_1868);
or U7846 (N_7846,N_610,N_413);
nand U7847 (N_7847,N_3793,N_2425);
and U7848 (N_7848,N_1148,N_4777);
nand U7849 (N_7849,N_4955,N_1106);
or U7850 (N_7850,N_2325,N_2119);
or U7851 (N_7851,N_1299,N_4584);
nor U7852 (N_7852,N_1813,N_997);
or U7853 (N_7853,N_184,N_3439);
or U7854 (N_7854,N_2477,N_3938);
nand U7855 (N_7855,N_152,N_3938);
nand U7856 (N_7856,N_4518,N_2084);
or U7857 (N_7857,N_3317,N_4352);
nor U7858 (N_7858,N_560,N_4575);
nor U7859 (N_7859,N_1530,N_1926);
or U7860 (N_7860,N_3276,N_1651);
nand U7861 (N_7861,N_4242,N_510);
nand U7862 (N_7862,N_808,N_794);
nand U7863 (N_7863,N_2410,N_3823);
or U7864 (N_7864,N_1697,N_4983);
xor U7865 (N_7865,N_716,N_136);
nand U7866 (N_7866,N_4775,N_2637);
nand U7867 (N_7867,N_910,N_3731);
nand U7868 (N_7868,N_668,N_1107);
and U7869 (N_7869,N_772,N_2414);
nand U7870 (N_7870,N_397,N_2103);
or U7871 (N_7871,N_395,N_1858);
and U7872 (N_7872,N_4673,N_3464);
nand U7873 (N_7873,N_3253,N_4808);
and U7874 (N_7874,N_4975,N_4982);
and U7875 (N_7875,N_2406,N_427);
nand U7876 (N_7876,N_3958,N_35);
nand U7877 (N_7877,N_2866,N_3791);
nor U7878 (N_7878,N_2054,N_4991);
nor U7879 (N_7879,N_4211,N_796);
nand U7880 (N_7880,N_1792,N_3834);
and U7881 (N_7881,N_3570,N_3842);
or U7882 (N_7882,N_3625,N_1465);
nand U7883 (N_7883,N_3538,N_585);
nor U7884 (N_7884,N_4324,N_4846);
nor U7885 (N_7885,N_4642,N_645);
xnor U7886 (N_7886,N_3138,N_399);
and U7887 (N_7887,N_2464,N_2264);
nand U7888 (N_7888,N_1986,N_4270);
and U7889 (N_7889,N_2552,N_4131);
nand U7890 (N_7890,N_3151,N_1545);
or U7891 (N_7891,N_1524,N_3534);
nor U7892 (N_7892,N_978,N_1107);
nand U7893 (N_7893,N_2716,N_388);
nor U7894 (N_7894,N_3368,N_3192);
or U7895 (N_7895,N_2538,N_4763);
nor U7896 (N_7896,N_3966,N_1357);
or U7897 (N_7897,N_1832,N_2219);
or U7898 (N_7898,N_2897,N_2935);
nor U7899 (N_7899,N_4244,N_1883);
nor U7900 (N_7900,N_2550,N_2588);
nand U7901 (N_7901,N_4633,N_2895);
or U7902 (N_7902,N_1439,N_4560);
nand U7903 (N_7903,N_1161,N_1538);
or U7904 (N_7904,N_4081,N_3823);
and U7905 (N_7905,N_4422,N_1345);
nor U7906 (N_7906,N_3725,N_2319);
nor U7907 (N_7907,N_873,N_1584);
nor U7908 (N_7908,N_3941,N_3091);
or U7909 (N_7909,N_1166,N_967);
nand U7910 (N_7910,N_1988,N_1857);
nand U7911 (N_7911,N_4370,N_2899);
nand U7912 (N_7912,N_3694,N_1464);
or U7913 (N_7913,N_3922,N_2839);
nor U7914 (N_7914,N_3037,N_1975);
nand U7915 (N_7915,N_2273,N_4877);
nor U7916 (N_7916,N_1550,N_4489);
xnor U7917 (N_7917,N_2519,N_3821);
xnor U7918 (N_7918,N_533,N_77);
and U7919 (N_7919,N_2899,N_3452);
nand U7920 (N_7920,N_2462,N_4817);
nor U7921 (N_7921,N_3958,N_3333);
nand U7922 (N_7922,N_3380,N_1617);
and U7923 (N_7923,N_1718,N_2041);
nand U7924 (N_7924,N_2294,N_145);
nor U7925 (N_7925,N_4681,N_1552);
and U7926 (N_7926,N_2679,N_101);
xnor U7927 (N_7927,N_763,N_3104);
nor U7928 (N_7928,N_1658,N_118);
and U7929 (N_7929,N_3958,N_2369);
or U7930 (N_7930,N_1304,N_997);
and U7931 (N_7931,N_1067,N_1486);
nor U7932 (N_7932,N_3317,N_3140);
nand U7933 (N_7933,N_190,N_1533);
nand U7934 (N_7934,N_4002,N_4150);
or U7935 (N_7935,N_1634,N_3523);
xnor U7936 (N_7936,N_3623,N_1947);
nand U7937 (N_7937,N_2778,N_3362);
or U7938 (N_7938,N_2674,N_423);
nor U7939 (N_7939,N_1133,N_1475);
xor U7940 (N_7940,N_3350,N_2815);
and U7941 (N_7941,N_145,N_893);
and U7942 (N_7942,N_2836,N_4069);
nand U7943 (N_7943,N_2958,N_738);
nor U7944 (N_7944,N_1736,N_4805);
or U7945 (N_7945,N_4559,N_3573);
and U7946 (N_7946,N_4954,N_2499);
nand U7947 (N_7947,N_4028,N_799);
nor U7948 (N_7948,N_368,N_2222);
nand U7949 (N_7949,N_1158,N_3048);
and U7950 (N_7950,N_1418,N_3937);
nor U7951 (N_7951,N_4618,N_523);
or U7952 (N_7952,N_1977,N_346);
or U7953 (N_7953,N_380,N_1304);
nor U7954 (N_7954,N_4987,N_4307);
nand U7955 (N_7955,N_2306,N_4691);
or U7956 (N_7956,N_4141,N_2765);
nor U7957 (N_7957,N_1413,N_3078);
nor U7958 (N_7958,N_4034,N_2300);
and U7959 (N_7959,N_1967,N_2101);
or U7960 (N_7960,N_1700,N_3895);
or U7961 (N_7961,N_1044,N_3372);
and U7962 (N_7962,N_3705,N_4382);
nor U7963 (N_7963,N_2973,N_4608);
and U7964 (N_7964,N_4713,N_3614);
xnor U7965 (N_7965,N_2119,N_131);
or U7966 (N_7966,N_1828,N_1112);
or U7967 (N_7967,N_1400,N_2596);
nor U7968 (N_7968,N_3370,N_965);
nand U7969 (N_7969,N_2598,N_1310);
nand U7970 (N_7970,N_3832,N_18);
nand U7971 (N_7971,N_1358,N_2212);
xnor U7972 (N_7972,N_1681,N_1904);
and U7973 (N_7973,N_2543,N_3056);
nand U7974 (N_7974,N_3031,N_1707);
or U7975 (N_7975,N_1195,N_982);
nor U7976 (N_7976,N_442,N_516);
nand U7977 (N_7977,N_3752,N_536);
nand U7978 (N_7978,N_3525,N_3052);
and U7979 (N_7979,N_3828,N_4895);
nand U7980 (N_7980,N_2027,N_3524);
nor U7981 (N_7981,N_1706,N_4518);
nor U7982 (N_7982,N_3746,N_3115);
and U7983 (N_7983,N_1673,N_467);
xnor U7984 (N_7984,N_4801,N_4571);
nand U7985 (N_7985,N_2083,N_2647);
nand U7986 (N_7986,N_1371,N_1555);
nor U7987 (N_7987,N_4733,N_526);
nor U7988 (N_7988,N_3742,N_707);
nand U7989 (N_7989,N_3589,N_750);
and U7990 (N_7990,N_39,N_1587);
or U7991 (N_7991,N_3065,N_3166);
or U7992 (N_7992,N_4930,N_751);
and U7993 (N_7993,N_2986,N_1055);
and U7994 (N_7994,N_1133,N_3459);
nand U7995 (N_7995,N_4580,N_3579);
and U7996 (N_7996,N_755,N_1257);
and U7997 (N_7997,N_1246,N_2495);
or U7998 (N_7998,N_4935,N_2717);
nor U7999 (N_7999,N_2861,N_540);
and U8000 (N_8000,N_2651,N_4848);
or U8001 (N_8001,N_3183,N_2678);
xnor U8002 (N_8002,N_4328,N_1344);
and U8003 (N_8003,N_1572,N_2083);
nand U8004 (N_8004,N_1420,N_2730);
or U8005 (N_8005,N_2712,N_19);
nand U8006 (N_8006,N_4167,N_890);
nor U8007 (N_8007,N_1135,N_650);
and U8008 (N_8008,N_3759,N_3860);
xor U8009 (N_8009,N_551,N_3596);
and U8010 (N_8010,N_758,N_3290);
and U8011 (N_8011,N_2516,N_3507);
and U8012 (N_8012,N_1650,N_875);
xnor U8013 (N_8013,N_2727,N_1558);
or U8014 (N_8014,N_1574,N_1447);
or U8015 (N_8015,N_2083,N_306);
and U8016 (N_8016,N_882,N_1649);
nand U8017 (N_8017,N_1897,N_1643);
or U8018 (N_8018,N_3845,N_1308);
or U8019 (N_8019,N_3350,N_1032);
and U8020 (N_8020,N_1436,N_4027);
xor U8021 (N_8021,N_4687,N_1226);
nor U8022 (N_8022,N_748,N_81);
nand U8023 (N_8023,N_3757,N_2896);
xor U8024 (N_8024,N_1764,N_4468);
and U8025 (N_8025,N_1441,N_2889);
nand U8026 (N_8026,N_4867,N_2830);
nand U8027 (N_8027,N_1992,N_1438);
nor U8028 (N_8028,N_690,N_115);
or U8029 (N_8029,N_3454,N_3987);
nor U8030 (N_8030,N_3565,N_4769);
or U8031 (N_8031,N_70,N_2753);
nand U8032 (N_8032,N_1395,N_64);
or U8033 (N_8033,N_3824,N_483);
nand U8034 (N_8034,N_3432,N_3269);
nand U8035 (N_8035,N_2924,N_4805);
and U8036 (N_8036,N_1501,N_4821);
nand U8037 (N_8037,N_2365,N_3417);
nand U8038 (N_8038,N_1822,N_4943);
or U8039 (N_8039,N_944,N_2110);
and U8040 (N_8040,N_1917,N_1096);
and U8041 (N_8041,N_993,N_2842);
nand U8042 (N_8042,N_4728,N_1316);
and U8043 (N_8043,N_1900,N_219);
nor U8044 (N_8044,N_2125,N_2269);
and U8045 (N_8045,N_1015,N_194);
nand U8046 (N_8046,N_4528,N_2504);
or U8047 (N_8047,N_3370,N_4917);
and U8048 (N_8048,N_2688,N_1937);
nand U8049 (N_8049,N_954,N_1440);
xor U8050 (N_8050,N_1623,N_544);
nor U8051 (N_8051,N_2874,N_749);
and U8052 (N_8052,N_1081,N_4281);
or U8053 (N_8053,N_3609,N_2570);
nor U8054 (N_8054,N_3325,N_4325);
nand U8055 (N_8055,N_3771,N_2591);
or U8056 (N_8056,N_2421,N_395);
nand U8057 (N_8057,N_1598,N_282);
and U8058 (N_8058,N_2077,N_2938);
nand U8059 (N_8059,N_1992,N_299);
nor U8060 (N_8060,N_992,N_4342);
nor U8061 (N_8061,N_3951,N_2736);
or U8062 (N_8062,N_1877,N_4565);
and U8063 (N_8063,N_3646,N_357);
nor U8064 (N_8064,N_427,N_3082);
and U8065 (N_8065,N_2743,N_3030);
or U8066 (N_8066,N_2323,N_3533);
or U8067 (N_8067,N_1511,N_2858);
or U8068 (N_8068,N_1589,N_3797);
nor U8069 (N_8069,N_3791,N_812);
or U8070 (N_8070,N_45,N_464);
nand U8071 (N_8071,N_3076,N_1446);
and U8072 (N_8072,N_4407,N_2898);
or U8073 (N_8073,N_4469,N_3394);
nand U8074 (N_8074,N_455,N_3338);
and U8075 (N_8075,N_3538,N_1644);
nor U8076 (N_8076,N_1553,N_783);
or U8077 (N_8077,N_237,N_2253);
or U8078 (N_8078,N_391,N_4186);
and U8079 (N_8079,N_2208,N_3214);
nor U8080 (N_8080,N_2649,N_2068);
or U8081 (N_8081,N_3251,N_3272);
or U8082 (N_8082,N_3385,N_586);
and U8083 (N_8083,N_1148,N_3395);
nor U8084 (N_8084,N_1339,N_2207);
and U8085 (N_8085,N_1408,N_4909);
and U8086 (N_8086,N_4430,N_823);
and U8087 (N_8087,N_402,N_1724);
nand U8088 (N_8088,N_1898,N_982);
nand U8089 (N_8089,N_1902,N_3556);
or U8090 (N_8090,N_3779,N_3757);
nor U8091 (N_8091,N_4354,N_3761);
nand U8092 (N_8092,N_2277,N_3275);
nand U8093 (N_8093,N_54,N_4314);
and U8094 (N_8094,N_3361,N_1174);
or U8095 (N_8095,N_969,N_971);
nor U8096 (N_8096,N_1228,N_4704);
nand U8097 (N_8097,N_464,N_2254);
or U8098 (N_8098,N_2395,N_1976);
nand U8099 (N_8099,N_2101,N_2009);
and U8100 (N_8100,N_4042,N_4732);
or U8101 (N_8101,N_1169,N_596);
nor U8102 (N_8102,N_2814,N_3433);
xnor U8103 (N_8103,N_2887,N_4964);
nor U8104 (N_8104,N_4924,N_1956);
nor U8105 (N_8105,N_4786,N_752);
nor U8106 (N_8106,N_445,N_1762);
nor U8107 (N_8107,N_4439,N_3730);
nor U8108 (N_8108,N_4431,N_2478);
nand U8109 (N_8109,N_4033,N_4204);
nor U8110 (N_8110,N_4957,N_383);
or U8111 (N_8111,N_4107,N_4173);
or U8112 (N_8112,N_2632,N_4935);
and U8113 (N_8113,N_3695,N_4499);
or U8114 (N_8114,N_165,N_3089);
xnor U8115 (N_8115,N_2989,N_1825);
and U8116 (N_8116,N_2323,N_3544);
and U8117 (N_8117,N_4311,N_3565);
nor U8118 (N_8118,N_4946,N_1936);
and U8119 (N_8119,N_374,N_1120);
and U8120 (N_8120,N_1216,N_1822);
nand U8121 (N_8121,N_482,N_78);
and U8122 (N_8122,N_3860,N_4841);
nor U8123 (N_8123,N_614,N_4954);
nand U8124 (N_8124,N_3752,N_4992);
nor U8125 (N_8125,N_12,N_4060);
nand U8126 (N_8126,N_2410,N_4241);
or U8127 (N_8127,N_4056,N_4939);
xor U8128 (N_8128,N_2425,N_4270);
nor U8129 (N_8129,N_3616,N_4210);
nand U8130 (N_8130,N_3876,N_2456);
and U8131 (N_8131,N_4585,N_1780);
or U8132 (N_8132,N_4768,N_296);
or U8133 (N_8133,N_4091,N_4984);
nand U8134 (N_8134,N_2637,N_4797);
nor U8135 (N_8135,N_3318,N_1635);
nor U8136 (N_8136,N_4533,N_1822);
nor U8137 (N_8137,N_4633,N_2486);
xnor U8138 (N_8138,N_2098,N_823);
nand U8139 (N_8139,N_1662,N_3083);
nor U8140 (N_8140,N_3019,N_2195);
or U8141 (N_8141,N_3708,N_4367);
nor U8142 (N_8142,N_1744,N_2447);
nor U8143 (N_8143,N_4913,N_2730);
nor U8144 (N_8144,N_3583,N_2633);
and U8145 (N_8145,N_317,N_605);
xor U8146 (N_8146,N_4616,N_220);
or U8147 (N_8147,N_4514,N_836);
nand U8148 (N_8148,N_1364,N_2406);
and U8149 (N_8149,N_1606,N_304);
or U8150 (N_8150,N_2191,N_3966);
nand U8151 (N_8151,N_493,N_3821);
xor U8152 (N_8152,N_2915,N_2620);
and U8153 (N_8153,N_720,N_1071);
nor U8154 (N_8154,N_4200,N_2465);
or U8155 (N_8155,N_278,N_721);
nand U8156 (N_8156,N_2740,N_3314);
nor U8157 (N_8157,N_818,N_662);
nand U8158 (N_8158,N_3851,N_2056);
or U8159 (N_8159,N_884,N_4308);
nor U8160 (N_8160,N_2538,N_3233);
xnor U8161 (N_8161,N_4812,N_616);
or U8162 (N_8162,N_4373,N_2105);
or U8163 (N_8163,N_1343,N_3633);
nor U8164 (N_8164,N_4918,N_1213);
nor U8165 (N_8165,N_1913,N_964);
nand U8166 (N_8166,N_1357,N_302);
nand U8167 (N_8167,N_3712,N_2825);
or U8168 (N_8168,N_3883,N_692);
xor U8169 (N_8169,N_4594,N_735);
or U8170 (N_8170,N_3568,N_4809);
and U8171 (N_8171,N_155,N_1536);
nand U8172 (N_8172,N_814,N_1794);
nor U8173 (N_8173,N_2880,N_2632);
and U8174 (N_8174,N_3645,N_4972);
or U8175 (N_8175,N_2431,N_1260);
xnor U8176 (N_8176,N_71,N_642);
or U8177 (N_8177,N_2344,N_3277);
nor U8178 (N_8178,N_4144,N_999);
nor U8179 (N_8179,N_4344,N_1609);
nand U8180 (N_8180,N_4071,N_761);
or U8181 (N_8181,N_4487,N_3004);
nand U8182 (N_8182,N_3943,N_880);
nor U8183 (N_8183,N_1754,N_2297);
nor U8184 (N_8184,N_3151,N_3602);
xor U8185 (N_8185,N_4873,N_3871);
nor U8186 (N_8186,N_3512,N_2665);
nand U8187 (N_8187,N_1734,N_4450);
xor U8188 (N_8188,N_4701,N_134);
xor U8189 (N_8189,N_1643,N_289);
nand U8190 (N_8190,N_20,N_1761);
or U8191 (N_8191,N_2847,N_582);
or U8192 (N_8192,N_1204,N_2457);
nor U8193 (N_8193,N_1412,N_2449);
nor U8194 (N_8194,N_4287,N_208);
and U8195 (N_8195,N_3623,N_2268);
xor U8196 (N_8196,N_364,N_3737);
nand U8197 (N_8197,N_416,N_1730);
and U8198 (N_8198,N_226,N_1678);
nand U8199 (N_8199,N_238,N_1709);
nor U8200 (N_8200,N_3650,N_1773);
and U8201 (N_8201,N_319,N_4576);
xnor U8202 (N_8202,N_3050,N_1313);
or U8203 (N_8203,N_1326,N_3675);
nor U8204 (N_8204,N_4944,N_1594);
and U8205 (N_8205,N_2833,N_2189);
nor U8206 (N_8206,N_709,N_1730);
xor U8207 (N_8207,N_3639,N_2345);
nand U8208 (N_8208,N_1784,N_482);
or U8209 (N_8209,N_3682,N_2580);
and U8210 (N_8210,N_1061,N_2765);
xnor U8211 (N_8211,N_2664,N_2909);
nor U8212 (N_8212,N_150,N_3662);
or U8213 (N_8213,N_4877,N_3841);
nand U8214 (N_8214,N_225,N_1283);
nor U8215 (N_8215,N_3575,N_3724);
or U8216 (N_8216,N_2119,N_4887);
nand U8217 (N_8217,N_482,N_2852);
xnor U8218 (N_8218,N_663,N_2316);
xor U8219 (N_8219,N_184,N_2267);
or U8220 (N_8220,N_4054,N_4723);
nand U8221 (N_8221,N_3304,N_715);
and U8222 (N_8222,N_4556,N_495);
nand U8223 (N_8223,N_2560,N_3510);
nor U8224 (N_8224,N_2714,N_1641);
or U8225 (N_8225,N_4790,N_4308);
nor U8226 (N_8226,N_574,N_3945);
nand U8227 (N_8227,N_149,N_1776);
nand U8228 (N_8228,N_2457,N_1936);
or U8229 (N_8229,N_245,N_481);
nand U8230 (N_8230,N_1305,N_2898);
xnor U8231 (N_8231,N_1243,N_182);
nor U8232 (N_8232,N_1519,N_1958);
or U8233 (N_8233,N_3226,N_504);
or U8234 (N_8234,N_2516,N_2399);
nor U8235 (N_8235,N_3294,N_3386);
nor U8236 (N_8236,N_2165,N_151);
nor U8237 (N_8237,N_3712,N_4048);
and U8238 (N_8238,N_1087,N_1937);
xnor U8239 (N_8239,N_4891,N_1546);
nand U8240 (N_8240,N_348,N_742);
or U8241 (N_8241,N_1762,N_1450);
nand U8242 (N_8242,N_1124,N_209);
nor U8243 (N_8243,N_1722,N_2074);
nor U8244 (N_8244,N_716,N_3556);
nand U8245 (N_8245,N_1594,N_4527);
nand U8246 (N_8246,N_1429,N_2376);
nand U8247 (N_8247,N_1499,N_4920);
nand U8248 (N_8248,N_4295,N_4090);
and U8249 (N_8249,N_3520,N_4807);
xor U8250 (N_8250,N_3556,N_3689);
nor U8251 (N_8251,N_1237,N_3469);
nand U8252 (N_8252,N_2363,N_3048);
xor U8253 (N_8253,N_1156,N_2827);
nor U8254 (N_8254,N_970,N_1163);
nor U8255 (N_8255,N_3702,N_1412);
nand U8256 (N_8256,N_3072,N_1910);
or U8257 (N_8257,N_2859,N_3772);
xor U8258 (N_8258,N_79,N_3238);
nor U8259 (N_8259,N_3969,N_4940);
nor U8260 (N_8260,N_415,N_357);
and U8261 (N_8261,N_1510,N_3522);
or U8262 (N_8262,N_3737,N_490);
nand U8263 (N_8263,N_3688,N_472);
and U8264 (N_8264,N_4524,N_7);
and U8265 (N_8265,N_4364,N_1703);
or U8266 (N_8266,N_3141,N_2988);
nand U8267 (N_8267,N_2463,N_521);
or U8268 (N_8268,N_2222,N_4667);
and U8269 (N_8269,N_4275,N_2605);
nor U8270 (N_8270,N_2862,N_1289);
xnor U8271 (N_8271,N_634,N_2301);
or U8272 (N_8272,N_4856,N_2423);
and U8273 (N_8273,N_559,N_2590);
nand U8274 (N_8274,N_3222,N_4504);
xnor U8275 (N_8275,N_3911,N_3058);
nand U8276 (N_8276,N_1685,N_2078);
xor U8277 (N_8277,N_2803,N_1458);
nor U8278 (N_8278,N_2474,N_1988);
nor U8279 (N_8279,N_4788,N_1179);
or U8280 (N_8280,N_1600,N_3283);
nand U8281 (N_8281,N_1661,N_1313);
and U8282 (N_8282,N_442,N_802);
and U8283 (N_8283,N_1959,N_603);
nand U8284 (N_8284,N_2553,N_467);
and U8285 (N_8285,N_2560,N_4081);
and U8286 (N_8286,N_261,N_3356);
or U8287 (N_8287,N_1848,N_3260);
nor U8288 (N_8288,N_140,N_1346);
xor U8289 (N_8289,N_844,N_1029);
and U8290 (N_8290,N_1353,N_4174);
nor U8291 (N_8291,N_4512,N_980);
nor U8292 (N_8292,N_1532,N_3560);
and U8293 (N_8293,N_4783,N_506);
nand U8294 (N_8294,N_2408,N_568);
nor U8295 (N_8295,N_4092,N_396);
or U8296 (N_8296,N_2488,N_699);
and U8297 (N_8297,N_3269,N_4689);
nor U8298 (N_8298,N_1835,N_2726);
and U8299 (N_8299,N_2243,N_3816);
or U8300 (N_8300,N_4406,N_3225);
and U8301 (N_8301,N_4959,N_1002);
nand U8302 (N_8302,N_2070,N_168);
or U8303 (N_8303,N_4551,N_1390);
or U8304 (N_8304,N_1365,N_1270);
or U8305 (N_8305,N_3227,N_2580);
and U8306 (N_8306,N_894,N_1643);
nor U8307 (N_8307,N_1949,N_478);
or U8308 (N_8308,N_1075,N_2169);
nor U8309 (N_8309,N_4311,N_65);
and U8310 (N_8310,N_820,N_2338);
and U8311 (N_8311,N_3142,N_83);
or U8312 (N_8312,N_427,N_2394);
nand U8313 (N_8313,N_3582,N_2501);
xnor U8314 (N_8314,N_491,N_4345);
nand U8315 (N_8315,N_443,N_442);
or U8316 (N_8316,N_2367,N_423);
nor U8317 (N_8317,N_3588,N_4754);
nor U8318 (N_8318,N_1536,N_936);
nand U8319 (N_8319,N_2662,N_2059);
or U8320 (N_8320,N_4842,N_3080);
xor U8321 (N_8321,N_407,N_2355);
nand U8322 (N_8322,N_4456,N_655);
xnor U8323 (N_8323,N_119,N_537);
and U8324 (N_8324,N_533,N_4056);
nand U8325 (N_8325,N_2369,N_4595);
nand U8326 (N_8326,N_161,N_2470);
nor U8327 (N_8327,N_1976,N_1493);
xnor U8328 (N_8328,N_4238,N_294);
and U8329 (N_8329,N_2466,N_1472);
nand U8330 (N_8330,N_2768,N_3025);
or U8331 (N_8331,N_1465,N_2164);
or U8332 (N_8332,N_2853,N_719);
and U8333 (N_8333,N_4732,N_3131);
nand U8334 (N_8334,N_4863,N_1779);
nand U8335 (N_8335,N_111,N_2491);
xor U8336 (N_8336,N_2287,N_3658);
nand U8337 (N_8337,N_337,N_4713);
nand U8338 (N_8338,N_1156,N_3636);
or U8339 (N_8339,N_362,N_4201);
nand U8340 (N_8340,N_1757,N_1868);
nor U8341 (N_8341,N_3814,N_520);
and U8342 (N_8342,N_343,N_297);
nand U8343 (N_8343,N_3078,N_780);
or U8344 (N_8344,N_1263,N_1728);
nor U8345 (N_8345,N_4578,N_4535);
or U8346 (N_8346,N_4658,N_768);
nor U8347 (N_8347,N_3343,N_4051);
nand U8348 (N_8348,N_2432,N_1875);
nor U8349 (N_8349,N_2494,N_3646);
nand U8350 (N_8350,N_3915,N_2418);
nor U8351 (N_8351,N_2413,N_1962);
nand U8352 (N_8352,N_428,N_3643);
nor U8353 (N_8353,N_3122,N_216);
nand U8354 (N_8354,N_4628,N_4816);
nand U8355 (N_8355,N_437,N_3987);
nor U8356 (N_8356,N_4755,N_4582);
nand U8357 (N_8357,N_1296,N_4250);
or U8358 (N_8358,N_2431,N_452);
and U8359 (N_8359,N_4701,N_2269);
nand U8360 (N_8360,N_3784,N_1624);
nand U8361 (N_8361,N_4877,N_135);
nor U8362 (N_8362,N_4930,N_3012);
nor U8363 (N_8363,N_2590,N_1348);
xnor U8364 (N_8364,N_1746,N_4951);
xnor U8365 (N_8365,N_702,N_2409);
or U8366 (N_8366,N_4879,N_391);
or U8367 (N_8367,N_2849,N_1787);
and U8368 (N_8368,N_4354,N_2810);
or U8369 (N_8369,N_3030,N_1481);
and U8370 (N_8370,N_3983,N_2051);
or U8371 (N_8371,N_2331,N_4365);
or U8372 (N_8372,N_627,N_4518);
or U8373 (N_8373,N_2310,N_273);
or U8374 (N_8374,N_4750,N_879);
xor U8375 (N_8375,N_1777,N_2910);
xnor U8376 (N_8376,N_1413,N_1801);
nand U8377 (N_8377,N_3752,N_4968);
or U8378 (N_8378,N_986,N_4996);
and U8379 (N_8379,N_1460,N_695);
nand U8380 (N_8380,N_805,N_1964);
or U8381 (N_8381,N_956,N_1883);
nor U8382 (N_8382,N_2309,N_603);
xnor U8383 (N_8383,N_479,N_532);
or U8384 (N_8384,N_3668,N_3775);
nor U8385 (N_8385,N_992,N_1494);
and U8386 (N_8386,N_772,N_1643);
or U8387 (N_8387,N_2939,N_1779);
or U8388 (N_8388,N_70,N_2308);
and U8389 (N_8389,N_3148,N_2689);
xnor U8390 (N_8390,N_2993,N_1842);
nor U8391 (N_8391,N_920,N_322);
nand U8392 (N_8392,N_1049,N_4598);
nand U8393 (N_8393,N_4763,N_4039);
and U8394 (N_8394,N_1843,N_1627);
nor U8395 (N_8395,N_1534,N_738);
xnor U8396 (N_8396,N_4816,N_1438);
and U8397 (N_8397,N_2086,N_4909);
and U8398 (N_8398,N_794,N_1970);
or U8399 (N_8399,N_636,N_2079);
xnor U8400 (N_8400,N_595,N_175);
and U8401 (N_8401,N_3405,N_1631);
and U8402 (N_8402,N_993,N_748);
nor U8403 (N_8403,N_4868,N_402);
or U8404 (N_8404,N_1065,N_3070);
and U8405 (N_8405,N_4027,N_4720);
or U8406 (N_8406,N_3197,N_4928);
or U8407 (N_8407,N_810,N_453);
xnor U8408 (N_8408,N_1966,N_4362);
and U8409 (N_8409,N_3888,N_2503);
xor U8410 (N_8410,N_2054,N_1238);
or U8411 (N_8411,N_1776,N_2425);
xnor U8412 (N_8412,N_1336,N_3118);
and U8413 (N_8413,N_184,N_4593);
nor U8414 (N_8414,N_4283,N_495);
nand U8415 (N_8415,N_3806,N_2800);
nand U8416 (N_8416,N_2833,N_1761);
or U8417 (N_8417,N_563,N_2952);
and U8418 (N_8418,N_3363,N_4714);
nor U8419 (N_8419,N_3721,N_3505);
nor U8420 (N_8420,N_256,N_507);
nand U8421 (N_8421,N_3364,N_1136);
and U8422 (N_8422,N_4785,N_2879);
and U8423 (N_8423,N_1143,N_2748);
or U8424 (N_8424,N_2685,N_1553);
and U8425 (N_8425,N_3866,N_3205);
nor U8426 (N_8426,N_669,N_3164);
and U8427 (N_8427,N_4105,N_609);
nor U8428 (N_8428,N_3917,N_3340);
xor U8429 (N_8429,N_1727,N_1152);
and U8430 (N_8430,N_2824,N_4399);
nand U8431 (N_8431,N_1549,N_2066);
or U8432 (N_8432,N_3262,N_583);
nand U8433 (N_8433,N_1343,N_3944);
nand U8434 (N_8434,N_4515,N_4379);
and U8435 (N_8435,N_1843,N_1507);
nor U8436 (N_8436,N_1880,N_1727);
xnor U8437 (N_8437,N_2641,N_924);
and U8438 (N_8438,N_4537,N_4843);
nand U8439 (N_8439,N_4754,N_22);
or U8440 (N_8440,N_3908,N_58);
xnor U8441 (N_8441,N_4465,N_3480);
nor U8442 (N_8442,N_3754,N_1680);
nand U8443 (N_8443,N_1564,N_4683);
and U8444 (N_8444,N_3519,N_552);
xor U8445 (N_8445,N_4335,N_2495);
nand U8446 (N_8446,N_2591,N_4631);
nand U8447 (N_8447,N_2681,N_4362);
or U8448 (N_8448,N_3939,N_807);
nand U8449 (N_8449,N_4557,N_2686);
and U8450 (N_8450,N_3933,N_180);
or U8451 (N_8451,N_4720,N_2307);
or U8452 (N_8452,N_3125,N_1558);
or U8453 (N_8453,N_4628,N_610);
or U8454 (N_8454,N_1338,N_4071);
xor U8455 (N_8455,N_3141,N_1786);
or U8456 (N_8456,N_4598,N_3074);
nand U8457 (N_8457,N_390,N_613);
nand U8458 (N_8458,N_4883,N_2112);
nand U8459 (N_8459,N_2933,N_4312);
and U8460 (N_8460,N_4453,N_3182);
nor U8461 (N_8461,N_2161,N_4704);
xnor U8462 (N_8462,N_2416,N_1992);
and U8463 (N_8463,N_2451,N_1471);
or U8464 (N_8464,N_2307,N_3352);
nand U8465 (N_8465,N_566,N_1384);
and U8466 (N_8466,N_1612,N_1341);
nand U8467 (N_8467,N_732,N_841);
or U8468 (N_8468,N_2435,N_4222);
xor U8469 (N_8469,N_154,N_4910);
or U8470 (N_8470,N_1434,N_1182);
nand U8471 (N_8471,N_190,N_4263);
or U8472 (N_8472,N_3725,N_2787);
nor U8473 (N_8473,N_89,N_624);
and U8474 (N_8474,N_840,N_38);
xnor U8475 (N_8475,N_2925,N_2690);
and U8476 (N_8476,N_2833,N_3439);
and U8477 (N_8477,N_218,N_4582);
nand U8478 (N_8478,N_2518,N_982);
nand U8479 (N_8479,N_1801,N_897);
or U8480 (N_8480,N_3886,N_1007);
nor U8481 (N_8481,N_1229,N_2290);
nor U8482 (N_8482,N_1825,N_4336);
and U8483 (N_8483,N_817,N_2489);
nand U8484 (N_8484,N_2995,N_1297);
and U8485 (N_8485,N_1078,N_3163);
and U8486 (N_8486,N_3013,N_198);
and U8487 (N_8487,N_3503,N_2874);
nor U8488 (N_8488,N_853,N_2108);
or U8489 (N_8489,N_1383,N_2636);
and U8490 (N_8490,N_1396,N_433);
and U8491 (N_8491,N_3643,N_3046);
nor U8492 (N_8492,N_1627,N_2918);
nor U8493 (N_8493,N_372,N_212);
nand U8494 (N_8494,N_2298,N_4474);
or U8495 (N_8495,N_709,N_3202);
and U8496 (N_8496,N_1234,N_3980);
nor U8497 (N_8497,N_4626,N_116);
xnor U8498 (N_8498,N_2202,N_2179);
and U8499 (N_8499,N_257,N_4478);
xor U8500 (N_8500,N_1483,N_1095);
xor U8501 (N_8501,N_2168,N_3271);
and U8502 (N_8502,N_3989,N_4428);
nor U8503 (N_8503,N_2420,N_2966);
and U8504 (N_8504,N_4534,N_3250);
and U8505 (N_8505,N_4460,N_1798);
nand U8506 (N_8506,N_4599,N_1414);
nor U8507 (N_8507,N_3965,N_4252);
nand U8508 (N_8508,N_2074,N_1774);
nand U8509 (N_8509,N_162,N_368);
or U8510 (N_8510,N_157,N_4030);
and U8511 (N_8511,N_3859,N_2243);
or U8512 (N_8512,N_843,N_2063);
or U8513 (N_8513,N_4090,N_2882);
nand U8514 (N_8514,N_4187,N_3622);
nor U8515 (N_8515,N_695,N_378);
nor U8516 (N_8516,N_1032,N_3559);
nand U8517 (N_8517,N_4909,N_1763);
or U8518 (N_8518,N_2627,N_1741);
or U8519 (N_8519,N_1131,N_79);
or U8520 (N_8520,N_2244,N_4001);
nor U8521 (N_8521,N_653,N_309);
and U8522 (N_8522,N_1545,N_208);
and U8523 (N_8523,N_2038,N_2850);
nand U8524 (N_8524,N_1079,N_3250);
and U8525 (N_8525,N_2355,N_333);
or U8526 (N_8526,N_151,N_4711);
or U8527 (N_8527,N_1813,N_3942);
nor U8528 (N_8528,N_961,N_415);
or U8529 (N_8529,N_4985,N_3823);
or U8530 (N_8530,N_1758,N_2428);
and U8531 (N_8531,N_820,N_110);
or U8532 (N_8532,N_484,N_472);
nand U8533 (N_8533,N_3473,N_2326);
nand U8534 (N_8534,N_617,N_4870);
and U8535 (N_8535,N_4279,N_4138);
xnor U8536 (N_8536,N_2614,N_4488);
nand U8537 (N_8537,N_4267,N_1086);
nor U8538 (N_8538,N_4410,N_859);
nand U8539 (N_8539,N_1978,N_1066);
nand U8540 (N_8540,N_1118,N_3631);
and U8541 (N_8541,N_91,N_955);
nand U8542 (N_8542,N_24,N_1970);
or U8543 (N_8543,N_3178,N_1894);
nand U8544 (N_8544,N_2740,N_4949);
and U8545 (N_8545,N_2746,N_4107);
and U8546 (N_8546,N_3069,N_2616);
and U8547 (N_8547,N_4934,N_1392);
nand U8548 (N_8548,N_2114,N_4529);
or U8549 (N_8549,N_337,N_1664);
and U8550 (N_8550,N_4813,N_3101);
and U8551 (N_8551,N_3390,N_4364);
nor U8552 (N_8552,N_1359,N_958);
or U8553 (N_8553,N_3642,N_3898);
nor U8554 (N_8554,N_256,N_2857);
nor U8555 (N_8555,N_4536,N_100);
nand U8556 (N_8556,N_1194,N_2963);
and U8557 (N_8557,N_2484,N_2826);
nor U8558 (N_8558,N_1301,N_774);
and U8559 (N_8559,N_4046,N_2084);
and U8560 (N_8560,N_236,N_4274);
and U8561 (N_8561,N_3421,N_2107);
nand U8562 (N_8562,N_1325,N_1736);
and U8563 (N_8563,N_1978,N_365);
and U8564 (N_8564,N_1200,N_1499);
and U8565 (N_8565,N_4999,N_866);
nand U8566 (N_8566,N_129,N_4655);
xor U8567 (N_8567,N_2824,N_3966);
and U8568 (N_8568,N_2255,N_1438);
and U8569 (N_8569,N_4383,N_2002);
nor U8570 (N_8570,N_4929,N_3379);
xnor U8571 (N_8571,N_1749,N_3637);
and U8572 (N_8572,N_3824,N_2105);
and U8573 (N_8573,N_2625,N_796);
nor U8574 (N_8574,N_4706,N_79);
xor U8575 (N_8575,N_1304,N_436);
nand U8576 (N_8576,N_458,N_4854);
or U8577 (N_8577,N_2291,N_1659);
nand U8578 (N_8578,N_3958,N_3138);
and U8579 (N_8579,N_1934,N_1005);
or U8580 (N_8580,N_1888,N_1275);
nor U8581 (N_8581,N_457,N_301);
nor U8582 (N_8582,N_3524,N_4626);
and U8583 (N_8583,N_1737,N_36);
nor U8584 (N_8584,N_2725,N_577);
or U8585 (N_8585,N_4510,N_4240);
and U8586 (N_8586,N_3219,N_709);
nor U8587 (N_8587,N_3235,N_1339);
and U8588 (N_8588,N_731,N_3777);
and U8589 (N_8589,N_2052,N_1924);
nand U8590 (N_8590,N_2156,N_841);
nor U8591 (N_8591,N_457,N_939);
nand U8592 (N_8592,N_3946,N_3019);
nand U8593 (N_8593,N_3156,N_748);
nand U8594 (N_8594,N_3626,N_4728);
xor U8595 (N_8595,N_3317,N_3576);
xor U8596 (N_8596,N_2168,N_285);
or U8597 (N_8597,N_1842,N_678);
nand U8598 (N_8598,N_1884,N_518);
xor U8599 (N_8599,N_3390,N_4938);
and U8600 (N_8600,N_1468,N_4325);
and U8601 (N_8601,N_708,N_3309);
nor U8602 (N_8602,N_2787,N_1980);
and U8603 (N_8603,N_909,N_4058);
or U8604 (N_8604,N_2011,N_4182);
or U8605 (N_8605,N_4586,N_4237);
and U8606 (N_8606,N_163,N_3613);
and U8607 (N_8607,N_1231,N_3007);
nor U8608 (N_8608,N_2130,N_2174);
xnor U8609 (N_8609,N_1869,N_1665);
or U8610 (N_8610,N_1152,N_4367);
nor U8611 (N_8611,N_3985,N_568);
and U8612 (N_8612,N_1342,N_2230);
nor U8613 (N_8613,N_1254,N_3573);
nand U8614 (N_8614,N_1704,N_3459);
xor U8615 (N_8615,N_4774,N_2506);
nor U8616 (N_8616,N_1143,N_3534);
or U8617 (N_8617,N_3011,N_3698);
nor U8618 (N_8618,N_3870,N_4325);
and U8619 (N_8619,N_4442,N_1015);
and U8620 (N_8620,N_3550,N_1213);
nand U8621 (N_8621,N_122,N_4981);
nand U8622 (N_8622,N_4637,N_508);
and U8623 (N_8623,N_2349,N_2491);
nand U8624 (N_8624,N_262,N_1183);
and U8625 (N_8625,N_3328,N_3459);
nor U8626 (N_8626,N_3239,N_1383);
nor U8627 (N_8627,N_4030,N_2444);
nand U8628 (N_8628,N_4325,N_3750);
xnor U8629 (N_8629,N_2083,N_1471);
xnor U8630 (N_8630,N_1355,N_2198);
or U8631 (N_8631,N_2441,N_998);
nor U8632 (N_8632,N_3733,N_563);
nor U8633 (N_8633,N_1633,N_140);
nand U8634 (N_8634,N_2931,N_1704);
xnor U8635 (N_8635,N_4027,N_317);
or U8636 (N_8636,N_1591,N_2676);
or U8637 (N_8637,N_3871,N_2474);
or U8638 (N_8638,N_4884,N_758);
xor U8639 (N_8639,N_3652,N_132);
and U8640 (N_8640,N_3546,N_465);
nor U8641 (N_8641,N_2392,N_4107);
and U8642 (N_8642,N_2394,N_2882);
or U8643 (N_8643,N_3207,N_1214);
or U8644 (N_8644,N_918,N_2130);
or U8645 (N_8645,N_1773,N_4824);
nand U8646 (N_8646,N_1449,N_1908);
or U8647 (N_8647,N_1066,N_3721);
or U8648 (N_8648,N_3311,N_3579);
nand U8649 (N_8649,N_2468,N_2346);
nand U8650 (N_8650,N_1818,N_4119);
nor U8651 (N_8651,N_4540,N_4460);
and U8652 (N_8652,N_1930,N_932);
xor U8653 (N_8653,N_4815,N_3888);
or U8654 (N_8654,N_4912,N_4139);
nand U8655 (N_8655,N_3638,N_714);
or U8656 (N_8656,N_4979,N_108);
and U8657 (N_8657,N_4865,N_2203);
nor U8658 (N_8658,N_2425,N_992);
nand U8659 (N_8659,N_3910,N_3105);
nand U8660 (N_8660,N_4497,N_2958);
xnor U8661 (N_8661,N_3284,N_3163);
nand U8662 (N_8662,N_3909,N_865);
xnor U8663 (N_8663,N_624,N_2584);
or U8664 (N_8664,N_2080,N_4487);
or U8665 (N_8665,N_2135,N_2892);
xnor U8666 (N_8666,N_756,N_1437);
and U8667 (N_8667,N_801,N_3307);
nor U8668 (N_8668,N_4316,N_2743);
nor U8669 (N_8669,N_435,N_4559);
nor U8670 (N_8670,N_4475,N_4038);
or U8671 (N_8671,N_1766,N_4214);
xor U8672 (N_8672,N_4047,N_220);
and U8673 (N_8673,N_2137,N_2224);
or U8674 (N_8674,N_3661,N_3414);
nor U8675 (N_8675,N_4339,N_3895);
nand U8676 (N_8676,N_974,N_4847);
or U8677 (N_8677,N_1902,N_2781);
nor U8678 (N_8678,N_2107,N_4369);
nand U8679 (N_8679,N_1717,N_1728);
nor U8680 (N_8680,N_4058,N_4607);
nor U8681 (N_8681,N_427,N_2980);
nand U8682 (N_8682,N_1195,N_736);
and U8683 (N_8683,N_3090,N_599);
or U8684 (N_8684,N_411,N_3081);
or U8685 (N_8685,N_1015,N_4553);
and U8686 (N_8686,N_4974,N_27);
nand U8687 (N_8687,N_469,N_2095);
or U8688 (N_8688,N_2597,N_1476);
and U8689 (N_8689,N_4138,N_2269);
and U8690 (N_8690,N_968,N_1154);
nand U8691 (N_8691,N_422,N_1360);
or U8692 (N_8692,N_1569,N_453);
or U8693 (N_8693,N_2325,N_1371);
xor U8694 (N_8694,N_2146,N_1136);
and U8695 (N_8695,N_15,N_4140);
xnor U8696 (N_8696,N_1239,N_1012);
and U8697 (N_8697,N_4182,N_405);
and U8698 (N_8698,N_4258,N_1703);
nand U8699 (N_8699,N_693,N_1275);
or U8700 (N_8700,N_4729,N_1688);
nand U8701 (N_8701,N_4019,N_698);
nor U8702 (N_8702,N_1590,N_4031);
and U8703 (N_8703,N_2625,N_3316);
or U8704 (N_8704,N_515,N_3653);
nor U8705 (N_8705,N_2865,N_1837);
nand U8706 (N_8706,N_538,N_1721);
nand U8707 (N_8707,N_2321,N_4415);
nor U8708 (N_8708,N_4452,N_457);
or U8709 (N_8709,N_1395,N_1801);
or U8710 (N_8710,N_570,N_4348);
nor U8711 (N_8711,N_1650,N_3534);
nand U8712 (N_8712,N_1975,N_4271);
or U8713 (N_8713,N_18,N_4309);
nor U8714 (N_8714,N_3414,N_3819);
and U8715 (N_8715,N_677,N_1799);
nor U8716 (N_8716,N_4372,N_1545);
and U8717 (N_8717,N_919,N_128);
or U8718 (N_8718,N_4719,N_951);
nor U8719 (N_8719,N_3237,N_1172);
nor U8720 (N_8720,N_4544,N_1812);
nor U8721 (N_8721,N_3165,N_2367);
and U8722 (N_8722,N_2185,N_535);
and U8723 (N_8723,N_4623,N_4280);
and U8724 (N_8724,N_4839,N_840);
and U8725 (N_8725,N_1443,N_4808);
nand U8726 (N_8726,N_4866,N_1331);
nor U8727 (N_8727,N_827,N_1789);
or U8728 (N_8728,N_3766,N_2530);
or U8729 (N_8729,N_3285,N_3359);
xor U8730 (N_8730,N_4638,N_4506);
and U8731 (N_8731,N_1853,N_2811);
or U8732 (N_8732,N_853,N_2258);
and U8733 (N_8733,N_1096,N_4998);
or U8734 (N_8734,N_1715,N_3123);
and U8735 (N_8735,N_2552,N_4501);
nor U8736 (N_8736,N_3304,N_1112);
nand U8737 (N_8737,N_370,N_1913);
or U8738 (N_8738,N_2437,N_4801);
and U8739 (N_8739,N_4623,N_3593);
nand U8740 (N_8740,N_4572,N_904);
and U8741 (N_8741,N_3132,N_821);
xnor U8742 (N_8742,N_225,N_4961);
xnor U8743 (N_8743,N_3007,N_676);
nand U8744 (N_8744,N_51,N_3794);
nand U8745 (N_8745,N_1508,N_1989);
and U8746 (N_8746,N_3061,N_1554);
and U8747 (N_8747,N_3640,N_1532);
nand U8748 (N_8748,N_4816,N_3924);
nand U8749 (N_8749,N_3506,N_4916);
nand U8750 (N_8750,N_3882,N_1784);
nor U8751 (N_8751,N_1254,N_4726);
and U8752 (N_8752,N_632,N_2673);
and U8753 (N_8753,N_1319,N_1413);
nand U8754 (N_8754,N_4377,N_4771);
nand U8755 (N_8755,N_4632,N_559);
nor U8756 (N_8756,N_2099,N_3448);
and U8757 (N_8757,N_4555,N_2823);
nor U8758 (N_8758,N_1454,N_1481);
xor U8759 (N_8759,N_4599,N_3161);
xor U8760 (N_8760,N_252,N_3815);
xnor U8761 (N_8761,N_73,N_2200);
nand U8762 (N_8762,N_3667,N_4337);
nand U8763 (N_8763,N_3073,N_1630);
nand U8764 (N_8764,N_2407,N_3278);
nand U8765 (N_8765,N_2334,N_1549);
nor U8766 (N_8766,N_3253,N_546);
nand U8767 (N_8767,N_1473,N_3576);
and U8768 (N_8768,N_711,N_1507);
nand U8769 (N_8769,N_1475,N_2430);
xnor U8770 (N_8770,N_1589,N_1930);
nand U8771 (N_8771,N_940,N_1121);
nand U8772 (N_8772,N_903,N_3754);
nor U8773 (N_8773,N_4735,N_3610);
nand U8774 (N_8774,N_2979,N_2906);
and U8775 (N_8775,N_366,N_1481);
nand U8776 (N_8776,N_2693,N_1009);
nand U8777 (N_8777,N_696,N_1543);
and U8778 (N_8778,N_3434,N_1244);
nand U8779 (N_8779,N_52,N_1556);
or U8780 (N_8780,N_308,N_3790);
or U8781 (N_8781,N_1656,N_4973);
or U8782 (N_8782,N_1480,N_1956);
nand U8783 (N_8783,N_922,N_2987);
or U8784 (N_8784,N_3115,N_1391);
or U8785 (N_8785,N_4810,N_3106);
or U8786 (N_8786,N_2300,N_1127);
xor U8787 (N_8787,N_1508,N_2262);
or U8788 (N_8788,N_408,N_4613);
nor U8789 (N_8789,N_376,N_2166);
and U8790 (N_8790,N_4720,N_3856);
nand U8791 (N_8791,N_1046,N_2453);
nand U8792 (N_8792,N_3965,N_4979);
nor U8793 (N_8793,N_1443,N_2348);
nand U8794 (N_8794,N_2010,N_3407);
and U8795 (N_8795,N_831,N_4112);
xnor U8796 (N_8796,N_2370,N_3899);
and U8797 (N_8797,N_1860,N_3799);
nor U8798 (N_8798,N_3530,N_589);
or U8799 (N_8799,N_109,N_600);
nand U8800 (N_8800,N_1051,N_3065);
nor U8801 (N_8801,N_861,N_2810);
nand U8802 (N_8802,N_1751,N_4321);
and U8803 (N_8803,N_4107,N_452);
or U8804 (N_8804,N_517,N_176);
and U8805 (N_8805,N_1062,N_4029);
or U8806 (N_8806,N_2684,N_4549);
or U8807 (N_8807,N_672,N_2046);
nand U8808 (N_8808,N_558,N_4058);
and U8809 (N_8809,N_1142,N_832);
xor U8810 (N_8810,N_1299,N_3923);
and U8811 (N_8811,N_323,N_4363);
nand U8812 (N_8812,N_3516,N_1335);
and U8813 (N_8813,N_4345,N_2207);
and U8814 (N_8814,N_1408,N_2466);
nor U8815 (N_8815,N_2980,N_4226);
and U8816 (N_8816,N_2086,N_208);
and U8817 (N_8817,N_135,N_2538);
or U8818 (N_8818,N_2053,N_1991);
nand U8819 (N_8819,N_1412,N_2522);
nand U8820 (N_8820,N_171,N_2560);
nand U8821 (N_8821,N_4597,N_1965);
and U8822 (N_8822,N_4238,N_3757);
xnor U8823 (N_8823,N_2195,N_782);
xnor U8824 (N_8824,N_341,N_4453);
xnor U8825 (N_8825,N_2954,N_4401);
and U8826 (N_8826,N_4372,N_1546);
or U8827 (N_8827,N_1570,N_4951);
nor U8828 (N_8828,N_163,N_4783);
nand U8829 (N_8829,N_20,N_3394);
nor U8830 (N_8830,N_4597,N_2534);
nor U8831 (N_8831,N_11,N_2053);
and U8832 (N_8832,N_4386,N_3699);
nand U8833 (N_8833,N_41,N_6);
nand U8834 (N_8834,N_4873,N_2177);
nand U8835 (N_8835,N_4985,N_413);
or U8836 (N_8836,N_1288,N_822);
and U8837 (N_8837,N_3750,N_3542);
and U8838 (N_8838,N_1405,N_1687);
xnor U8839 (N_8839,N_3007,N_3038);
or U8840 (N_8840,N_2985,N_4559);
nand U8841 (N_8841,N_4397,N_3877);
nor U8842 (N_8842,N_3148,N_253);
or U8843 (N_8843,N_4752,N_3017);
and U8844 (N_8844,N_1966,N_4441);
or U8845 (N_8845,N_1166,N_1546);
or U8846 (N_8846,N_1571,N_3460);
and U8847 (N_8847,N_4982,N_1147);
nor U8848 (N_8848,N_349,N_1384);
xor U8849 (N_8849,N_4235,N_2220);
or U8850 (N_8850,N_3797,N_3690);
and U8851 (N_8851,N_1875,N_1262);
nand U8852 (N_8852,N_2135,N_132);
nor U8853 (N_8853,N_4688,N_2663);
and U8854 (N_8854,N_3985,N_4842);
and U8855 (N_8855,N_144,N_1693);
nand U8856 (N_8856,N_1521,N_2808);
nor U8857 (N_8857,N_2624,N_681);
or U8858 (N_8858,N_3661,N_4291);
or U8859 (N_8859,N_2023,N_746);
and U8860 (N_8860,N_2650,N_2751);
and U8861 (N_8861,N_2197,N_158);
or U8862 (N_8862,N_2043,N_3946);
nand U8863 (N_8863,N_3358,N_3948);
or U8864 (N_8864,N_3250,N_4957);
or U8865 (N_8865,N_2866,N_3750);
nand U8866 (N_8866,N_3039,N_3095);
nor U8867 (N_8867,N_2081,N_3537);
nand U8868 (N_8868,N_2860,N_2526);
and U8869 (N_8869,N_4527,N_4003);
or U8870 (N_8870,N_3210,N_1238);
xor U8871 (N_8871,N_699,N_4053);
xor U8872 (N_8872,N_1913,N_3022);
and U8873 (N_8873,N_4220,N_1946);
and U8874 (N_8874,N_1146,N_1340);
nand U8875 (N_8875,N_856,N_3925);
nor U8876 (N_8876,N_2584,N_3947);
nand U8877 (N_8877,N_4862,N_3859);
and U8878 (N_8878,N_242,N_2493);
and U8879 (N_8879,N_3518,N_4972);
nor U8880 (N_8880,N_4781,N_4474);
nor U8881 (N_8881,N_3867,N_1783);
xor U8882 (N_8882,N_4047,N_2095);
xor U8883 (N_8883,N_2863,N_3714);
nor U8884 (N_8884,N_1556,N_2513);
or U8885 (N_8885,N_3793,N_844);
xnor U8886 (N_8886,N_3362,N_2461);
xor U8887 (N_8887,N_491,N_4010);
and U8888 (N_8888,N_1164,N_3717);
or U8889 (N_8889,N_2551,N_2806);
and U8890 (N_8890,N_800,N_4107);
and U8891 (N_8891,N_4629,N_4588);
nor U8892 (N_8892,N_4860,N_329);
or U8893 (N_8893,N_3058,N_1753);
nand U8894 (N_8894,N_4980,N_1135);
and U8895 (N_8895,N_2142,N_4006);
nor U8896 (N_8896,N_1367,N_3577);
and U8897 (N_8897,N_4285,N_719);
nor U8898 (N_8898,N_276,N_3201);
and U8899 (N_8899,N_294,N_930);
nand U8900 (N_8900,N_1401,N_1998);
nand U8901 (N_8901,N_2674,N_4400);
or U8902 (N_8902,N_2163,N_457);
nand U8903 (N_8903,N_240,N_2289);
nor U8904 (N_8904,N_1541,N_2043);
and U8905 (N_8905,N_40,N_4775);
nor U8906 (N_8906,N_2755,N_841);
nor U8907 (N_8907,N_676,N_1986);
nand U8908 (N_8908,N_1334,N_2982);
xnor U8909 (N_8909,N_2880,N_2425);
nand U8910 (N_8910,N_166,N_1881);
nor U8911 (N_8911,N_98,N_753);
or U8912 (N_8912,N_1031,N_960);
nor U8913 (N_8913,N_2474,N_649);
and U8914 (N_8914,N_4455,N_880);
and U8915 (N_8915,N_2353,N_54);
or U8916 (N_8916,N_1721,N_3833);
nand U8917 (N_8917,N_2454,N_1778);
and U8918 (N_8918,N_1870,N_2235);
nand U8919 (N_8919,N_4592,N_4771);
nand U8920 (N_8920,N_3417,N_279);
and U8921 (N_8921,N_1932,N_2662);
nand U8922 (N_8922,N_3587,N_17);
nor U8923 (N_8923,N_87,N_17);
nor U8924 (N_8924,N_1097,N_1027);
and U8925 (N_8925,N_1153,N_2998);
xnor U8926 (N_8926,N_4327,N_3227);
and U8927 (N_8927,N_3079,N_2792);
or U8928 (N_8928,N_238,N_3535);
and U8929 (N_8929,N_4393,N_2969);
nor U8930 (N_8930,N_2776,N_3470);
nand U8931 (N_8931,N_3067,N_3655);
and U8932 (N_8932,N_3002,N_2958);
or U8933 (N_8933,N_3658,N_4395);
nor U8934 (N_8934,N_1668,N_1373);
and U8935 (N_8935,N_4426,N_614);
xnor U8936 (N_8936,N_2700,N_3773);
or U8937 (N_8937,N_268,N_3866);
or U8938 (N_8938,N_3732,N_1267);
or U8939 (N_8939,N_1569,N_2206);
or U8940 (N_8940,N_1631,N_290);
nand U8941 (N_8941,N_2576,N_3019);
nor U8942 (N_8942,N_2621,N_2044);
nand U8943 (N_8943,N_3098,N_410);
or U8944 (N_8944,N_1847,N_178);
and U8945 (N_8945,N_670,N_4902);
and U8946 (N_8946,N_3103,N_1468);
or U8947 (N_8947,N_2309,N_3251);
nand U8948 (N_8948,N_1760,N_3697);
nand U8949 (N_8949,N_595,N_4252);
nor U8950 (N_8950,N_2256,N_4659);
and U8951 (N_8951,N_3595,N_904);
nor U8952 (N_8952,N_1684,N_3961);
and U8953 (N_8953,N_865,N_2713);
and U8954 (N_8954,N_1019,N_578);
nor U8955 (N_8955,N_2395,N_4330);
nor U8956 (N_8956,N_77,N_3768);
and U8957 (N_8957,N_3244,N_3577);
nand U8958 (N_8958,N_685,N_875);
and U8959 (N_8959,N_77,N_2806);
nand U8960 (N_8960,N_2603,N_3932);
and U8961 (N_8961,N_2181,N_557);
nand U8962 (N_8962,N_4239,N_316);
nor U8963 (N_8963,N_4707,N_3983);
xnor U8964 (N_8964,N_3510,N_458);
nand U8965 (N_8965,N_1325,N_4260);
xor U8966 (N_8966,N_3185,N_1884);
xor U8967 (N_8967,N_2460,N_1869);
and U8968 (N_8968,N_2512,N_2719);
or U8969 (N_8969,N_3953,N_4469);
or U8970 (N_8970,N_4084,N_1268);
and U8971 (N_8971,N_2243,N_2366);
nand U8972 (N_8972,N_4263,N_1658);
nand U8973 (N_8973,N_2579,N_2709);
nand U8974 (N_8974,N_580,N_1325);
nor U8975 (N_8975,N_4076,N_995);
or U8976 (N_8976,N_538,N_3346);
nor U8977 (N_8977,N_3674,N_3127);
or U8978 (N_8978,N_2878,N_137);
nor U8979 (N_8979,N_3150,N_1108);
or U8980 (N_8980,N_731,N_3357);
nand U8981 (N_8981,N_3131,N_92);
nand U8982 (N_8982,N_2006,N_732);
or U8983 (N_8983,N_226,N_1358);
xor U8984 (N_8984,N_2979,N_1444);
xor U8985 (N_8985,N_4916,N_2601);
and U8986 (N_8986,N_142,N_3064);
and U8987 (N_8987,N_1130,N_2922);
and U8988 (N_8988,N_874,N_4498);
or U8989 (N_8989,N_477,N_2105);
and U8990 (N_8990,N_1619,N_4527);
xnor U8991 (N_8991,N_2558,N_2924);
and U8992 (N_8992,N_3234,N_4898);
or U8993 (N_8993,N_410,N_4581);
nor U8994 (N_8994,N_1307,N_670);
and U8995 (N_8995,N_2405,N_4276);
or U8996 (N_8996,N_4679,N_2677);
nand U8997 (N_8997,N_3377,N_71);
or U8998 (N_8998,N_4959,N_918);
nor U8999 (N_8999,N_3990,N_2344);
or U9000 (N_9000,N_1553,N_1311);
and U9001 (N_9001,N_963,N_3789);
nand U9002 (N_9002,N_595,N_1344);
and U9003 (N_9003,N_4517,N_2938);
nand U9004 (N_9004,N_3716,N_1697);
or U9005 (N_9005,N_2790,N_994);
nand U9006 (N_9006,N_2436,N_3955);
nor U9007 (N_9007,N_3806,N_3326);
nand U9008 (N_9008,N_4728,N_1065);
and U9009 (N_9009,N_675,N_508);
xor U9010 (N_9010,N_2307,N_855);
and U9011 (N_9011,N_4752,N_3588);
and U9012 (N_9012,N_4469,N_1021);
xnor U9013 (N_9013,N_126,N_3945);
xnor U9014 (N_9014,N_4175,N_1178);
and U9015 (N_9015,N_1482,N_1705);
or U9016 (N_9016,N_4012,N_864);
nor U9017 (N_9017,N_1174,N_2375);
nor U9018 (N_9018,N_2730,N_2842);
or U9019 (N_9019,N_2513,N_2754);
or U9020 (N_9020,N_3589,N_4602);
and U9021 (N_9021,N_3277,N_101);
and U9022 (N_9022,N_3346,N_1253);
and U9023 (N_9023,N_2697,N_2164);
or U9024 (N_9024,N_1428,N_196);
and U9025 (N_9025,N_1812,N_421);
and U9026 (N_9026,N_869,N_643);
nor U9027 (N_9027,N_3393,N_4943);
or U9028 (N_9028,N_4803,N_2479);
and U9029 (N_9029,N_1208,N_4136);
nor U9030 (N_9030,N_3299,N_1557);
or U9031 (N_9031,N_3695,N_1661);
nand U9032 (N_9032,N_4904,N_1224);
or U9033 (N_9033,N_3007,N_2429);
xnor U9034 (N_9034,N_290,N_2065);
xnor U9035 (N_9035,N_3443,N_3529);
and U9036 (N_9036,N_1748,N_2514);
nand U9037 (N_9037,N_3337,N_1431);
and U9038 (N_9038,N_4911,N_4234);
xnor U9039 (N_9039,N_4108,N_450);
and U9040 (N_9040,N_2968,N_790);
xnor U9041 (N_9041,N_1002,N_1477);
nor U9042 (N_9042,N_4166,N_1393);
and U9043 (N_9043,N_3166,N_2362);
nand U9044 (N_9044,N_993,N_1467);
nor U9045 (N_9045,N_2566,N_779);
or U9046 (N_9046,N_373,N_1847);
or U9047 (N_9047,N_2952,N_2668);
nor U9048 (N_9048,N_4746,N_1721);
and U9049 (N_9049,N_3473,N_957);
nand U9050 (N_9050,N_1296,N_3580);
nor U9051 (N_9051,N_1166,N_1369);
or U9052 (N_9052,N_3905,N_3584);
nor U9053 (N_9053,N_24,N_4187);
or U9054 (N_9054,N_921,N_4003);
or U9055 (N_9055,N_111,N_3167);
nor U9056 (N_9056,N_4471,N_474);
or U9057 (N_9057,N_3333,N_3233);
and U9058 (N_9058,N_968,N_1714);
and U9059 (N_9059,N_1873,N_752);
xnor U9060 (N_9060,N_3122,N_2099);
nor U9061 (N_9061,N_2042,N_1076);
and U9062 (N_9062,N_3862,N_1179);
nand U9063 (N_9063,N_4716,N_1208);
nor U9064 (N_9064,N_3025,N_4065);
and U9065 (N_9065,N_3617,N_97);
or U9066 (N_9066,N_4664,N_3756);
nand U9067 (N_9067,N_1856,N_2700);
and U9068 (N_9068,N_3770,N_2741);
nor U9069 (N_9069,N_1422,N_3303);
nor U9070 (N_9070,N_2493,N_147);
nand U9071 (N_9071,N_3166,N_1555);
and U9072 (N_9072,N_566,N_278);
nor U9073 (N_9073,N_4297,N_4031);
nor U9074 (N_9074,N_868,N_3178);
nand U9075 (N_9075,N_1182,N_3164);
and U9076 (N_9076,N_2990,N_305);
and U9077 (N_9077,N_4064,N_958);
nor U9078 (N_9078,N_4229,N_1);
xnor U9079 (N_9079,N_1124,N_1695);
nand U9080 (N_9080,N_370,N_692);
and U9081 (N_9081,N_3250,N_2812);
or U9082 (N_9082,N_4522,N_1143);
and U9083 (N_9083,N_2951,N_3148);
and U9084 (N_9084,N_1719,N_4701);
xnor U9085 (N_9085,N_2962,N_3999);
or U9086 (N_9086,N_1940,N_1437);
xor U9087 (N_9087,N_1394,N_553);
or U9088 (N_9088,N_57,N_3077);
nand U9089 (N_9089,N_961,N_4406);
nor U9090 (N_9090,N_3497,N_2836);
nor U9091 (N_9091,N_1558,N_3171);
or U9092 (N_9092,N_3912,N_1557);
nand U9093 (N_9093,N_1864,N_3055);
xor U9094 (N_9094,N_1507,N_3310);
or U9095 (N_9095,N_3778,N_3212);
and U9096 (N_9096,N_4897,N_361);
nor U9097 (N_9097,N_152,N_3237);
nand U9098 (N_9098,N_188,N_4058);
nand U9099 (N_9099,N_3956,N_863);
nand U9100 (N_9100,N_4075,N_1499);
or U9101 (N_9101,N_1097,N_2519);
and U9102 (N_9102,N_4168,N_4915);
or U9103 (N_9103,N_4347,N_585);
and U9104 (N_9104,N_1061,N_3259);
and U9105 (N_9105,N_4781,N_4897);
nor U9106 (N_9106,N_2297,N_3790);
or U9107 (N_9107,N_2243,N_4748);
or U9108 (N_9108,N_3440,N_4398);
or U9109 (N_9109,N_3470,N_1674);
and U9110 (N_9110,N_925,N_2799);
nor U9111 (N_9111,N_4124,N_53);
and U9112 (N_9112,N_316,N_34);
nand U9113 (N_9113,N_2095,N_4116);
nand U9114 (N_9114,N_4744,N_2895);
nand U9115 (N_9115,N_2721,N_2137);
and U9116 (N_9116,N_2518,N_422);
or U9117 (N_9117,N_4477,N_183);
xnor U9118 (N_9118,N_1898,N_1807);
nand U9119 (N_9119,N_296,N_2851);
or U9120 (N_9120,N_4617,N_333);
or U9121 (N_9121,N_2819,N_4506);
nand U9122 (N_9122,N_3412,N_1092);
and U9123 (N_9123,N_1390,N_2316);
nor U9124 (N_9124,N_2329,N_2142);
and U9125 (N_9125,N_1336,N_4634);
and U9126 (N_9126,N_3505,N_1753);
nor U9127 (N_9127,N_964,N_513);
and U9128 (N_9128,N_4798,N_1221);
nand U9129 (N_9129,N_3069,N_1669);
nor U9130 (N_9130,N_4906,N_2759);
nand U9131 (N_9131,N_2324,N_4783);
nor U9132 (N_9132,N_3962,N_1005);
nand U9133 (N_9133,N_3777,N_538);
xnor U9134 (N_9134,N_3008,N_2482);
nand U9135 (N_9135,N_910,N_526);
nor U9136 (N_9136,N_1171,N_2932);
and U9137 (N_9137,N_2973,N_1668);
nor U9138 (N_9138,N_4417,N_2519);
nor U9139 (N_9139,N_1053,N_82);
xnor U9140 (N_9140,N_1737,N_1518);
xnor U9141 (N_9141,N_3874,N_1532);
or U9142 (N_9142,N_2350,N_395);
and U9143 (N_9143,N_1871,N_2817);
and U9144 (N_9144,N_1649,N_110);
nand U9145 (N_9145,N_2186,N_2885);
and U9146 (N_9146,N_2027,N_4475);
nand U9147 (N_9147,N_857,N_1012);
nand U9148 (N_9148,N_1288,N_1976);
and U9149 (N_9149,N_1820,N_841);
and U9150 (N_9150,N_1026,N_2722);
and U9151 (N_9151,N_3539,N_2472);
or U9152 (N_9152,N_1541,N_3469);
nand U9153 (N_9153,N_3290,N_1926);
and U9154 (N_9154,N_333,N_3864);
and U9155 (N_9155,N_3711,N_2930);
nand U9156 (N_9156,N_3559,N_49);
or U9157 (N_9157,N_3162,N_2444);
and U9158 (N_9158,N_3629,N_4978);
or U9159 (N_9159,N_1423,N_432);
or U9160 (N_9160,N_101,N_908);
and U9161 (N_9161,N_4141,N_4083);
xnor U9162 (N_9162,N_1367,N_1481);
nand U9163 (N_9163,N_4684,N_1521);
nor U9164 (N_9164,N_1266,N_4028);
and U9165 (N_9165,N_1894,N_1703);
nor U9166 (N_9166,N_424,N_3532);
and U9167 (N_9167,N_960,N_4416);
nor U9168 (N_9168,N_1151,N_961);
nand U9169 (N_9169,N_4362,N_4049);
nor U9170 (N_9170,N_178,N_4332);
nor U9171 (N_9171,N_1664,N_951);
nor U9172 (N_9172,N_3073,N_996);
nand U9173 (N_9173,N_2861,N_4974);
nor U9174 (N_9174,N_3656,N_1988);
nand U9175 (N_9175,N_1630,N_3192);
nand U9176 (N_9176,N_125,N_1243);
nand U9177 (N_9177,N_179,N_508);
nor U9178 (N_9178,N_674,N_101);
or U9179 (N_9179,N_1318,N_1551);
or U9180 (N_9180,N_1086,N_2409);
nor U9181 (N_9181,N_546,N_494);
or U9182 (N_9182,N_2233,N_1566);
nor U9183 (N_9183,N_3864,N_3121);
nor U9184 (N_9184,N_2431,N_2788);
or U9185 (N_9185,N_955,N_2184);
or U9186 (N_9186,N_3759,N_4406);
and U9187 (N_9187,N_2950,N_1200);
nand U9188 (N_9188,N_3216,N_3234);
xnor U9189 (N_9189,N_1442,N_1011);
xnor U9190 (N_9190,N_2142,N_4300);
and U9191 (N_9191,N_1119,N_250);
nor U9192 (N_9192,N_2682,N_2704);
nand U9193 (N_9193,N_516,N_343);
nor U9194 (N_9194,N_885,N_2621);
xnor U9195 (N_9195,N_2555,N_4636);
nand U9196 (N_9196,N_4283,N_1636);
nand U9197 (N_9197,N_3083,N_4977);
or U9198 (N_9198,N_728,N_3390);
and U9199 (N_9199,N_3289,N_3777);
or U9200 (N_9200,N_3841,N_2738);
or U9201 (N_9201,N_1502,N_2117);
xor U9202 (N_9202,N_4295,N_1311);
nand U9203 (N_9203,N_1321,N_1539);
and U9204 (N_9204,N_4624,N_3108);
or U9205 (N_9205,N_826,N_4426);
nand U9206 (N_9206,N_3320,N_4641);
and U9207 (N_9207,N_4556,N_158);
nand U9208 (N_9208,N_2506,N_340);
nand U9209 (N_9209,N_912,N_4335);
xor U9210 (N_9210,N_1011,N_849);
nor U9211 (N_9211,N_4644,N_2405);
or U9212 (N_9212,N_2666,N_3159);
or U9213 (N_9213,N_4750,N_1586);
nor U9214 (N_9214,N_329,N_4016);
nor U9215 (N_9215,N_3207,N_2715);
or U9216 (N_9216,N_2433,N_1358);
and U9217 (N_9217,N_1543,N_2495);
and U9218 (N_9218,N_1388,N_2003);
or U9219 (N_9219,N_4927,N_4059);
xor U9220 (N_9220,N_1418,N_1868);
and U9221 (N_9221,N_2395,N_2885);
or U9222 (N_9222,N_3772,N_1160);
nand U9223 (N_9223,N_3227,N_775);
xor U9224 (N_9224,N_661,N_1721);
or U9225 (N_9225,N_1965,N_2416);
nand U9226 (N_9226,N_1952,N_3211);
nand U9227 (N_9227,N_86,N_1461);
and U9228 (N_9228,N_2686,N_629);
nor U9229 (N_9229,N_1695,N_310);
and U9230 (N_9230,N_737,N_4955);
or U9231 (N_9231,N_2251,N_3755);
xor U9232 (N_9232,N_2368,N_4066);
and U9233 (N_9233,N_11,N_4172);
or U9234 (N_9234,N_3129,N_2712);
nand U9235 (N_9235,N_284,N_1108);
xor U9236 (N_9236,N_7,N_4383);
nor U9237 (N_9237,N_3263,N_792);
and U9238 (N_9238,N_4552,N_3007);
and U9239 (N_9239,N_2535,N_4073);
nor U9240 (N_9240,N_3924,N_163);
nand U9241 (N_9241,N_1312,N_127);
and U9242 (N_9242,N_1776,N_690);
and U9243 (N_9243,N_1299,N_716);
and U9244 (N_9244,N_1256,N_4816);
or U9245 (N_9245,N_4276,N_4627);
nand U9246 (N_9246,N_4529,N_4191);
nand U9247 (N_9247,N_3339,N_4927);
nor U9248 (N_9248,N_3266,N_132);
nor U9249 (N_9249,N_4780,N_1989);
and U9250 (N_9250,N_110,N_1317);
nor U9251 (N_9251,N_1058,N_4153);
or U9252 (N_9252,N_3619,N_3228);
nor U9253 (N_9253,N_1008,N_592);
and U9254 (N_9254,N_1121,N_766);
xnor U9255 (N_9255,N_4928,N_485);
nor U9256 (N_9256,N_604,N_4712);
and U9257 (N_9257,N_2785,N_3938);
nand U9258 (N_9258,N_4650,N_1266);
nand U9259 (N_9259,N_266,N_1179);
and U9260 (N_9260,N_1701,N_2580);
and U9261 (N_9261,N_2151,N_3162);
nor U9262 (N_9262,N_1834,N_2134);
nand U9263 (N_9263,N_2106,N_242);
nand U9264 (N_9264,N_1647,N_1441);
nand U9265 (N_9265,N_1306,N_404);
xnor U9266 (N_9266,N_2846,N_116);
and U9267 (N_9267,N_4419,N_1250);
and U9268 (N_9268,N_29,N_100);
and U9269 (N_9269,N_3810,N_1910);
or U9270 (N_9270,N_2919,N_3375);
nor U9271 (N_9271,N_148,N_3836);
or U9272 (N_9272,N_599,N_1476);
nand U9273 (N_9273,N_1335,N_2347);
or U9274 (N_9274,N_4944,N_1887);
nand U9275 (N_9275,N_4972,N_42);
and U9276 (N_9276,N_4989,N_529);
and U9277 (N_9277,N_117,N_914);
nand U9278 (N_9278,N_2423,N_1997);
nand U9279 (N_9279,N_978,N_4408);
nor U9280 (N_9280,N_4216,N_235);
or U9281 (N_9281,N_1343,N_531);
nand U9282 (N_9282,N_3706,N_547);
nand U9283 (N_9283,N_808,N_1744);
nor U9284 (N_9284,N_1958,N_3908);
nand U9285 (N_9285,N_2771,N_1898);
or U9286 (N_9286,N_1498,N_2558);
nor U9287 (N_9287,N_2139,N_4035);
or U9288 (N_9288,N_1476,N_2675);
or U9289 (N_9289,N_437,N_3857);
nand U9290 (N_9290,N_1568,N_2546);
nand U9291 (N_9291,N_145,N_995);
nand U9292 (N_9292,N_2297,N_1799);
and U9293 (N_9293,N_4920,N_4537);
nand U9294 (N_9294,N_2387,N_3110);
and U9295 (N_9295,N_2380,N_2191);
or U9296 (N_9296,N_3347,N_2964);
and U9297 (N_9297,N_509,N_4790);
nor U9298 (N_9298,N_1281,N_4454);
nand U9299 (N_9299,N_4712,N_3924);
nor U9300 (N_9300,N_3450,N_4280);
and U9301 (N_9301,N_1150,N_3820);
xnor U9302 (N_9302,N_4578,N_1397);
nor U9303 (N_9303,N_2458,N_2989);
or U9304 (N_9304,N_117,N_1658);
nand U9305 (N_9305,N_4239,N_2049);
nand U9306 (N_9306,N_1440,N_4600);
nand U9307 (N_9307,N_1693,N_4447);
and U9308 (N_9308,N_3128,N_2809);
and U9309 (N_9309,N_706,N_3243);
and U9310 (N_9310,N_3812,N_467);
nor U9311 (N_9311,N_2171,N_1638);
and U9312 (N_9312,N_4421,N_907);
and U9313 (N_9313,N_3976,N_1376);
nand U9314 (N_9314,N_4465,N_4376);
or U9315 (N_9315,N_1322,N_535);
or U9316 (N_9316,N_1202,N_1544);
nand U9317 (N_9317,N_1996,N_2839);
nand U9318 (N_9318,N_892,N_7);
nand U9319 (N_9319,N_4667,N_3637);
xnor U9320 (N_9320,N_2126,N_2741);
and U9321 (N_9321,N_4185,N_4072);
and U9322 (N_9322,N_2748,N_2228);
xnor U9323 (N_9323,N_4658,N_252);
and U9324 (N_9324,N_100,N_3392);
or U9325 (N_9325,N_2708,N_3057);
nand U9326 (N_9326,N_2242,N_4023);
nand U9327 (N_9327,N_4386,N_710);
nor U9328 (N_9328,N_1084,N_4419);
nand U9329 (N_9329,N_1815,N_270);
or U9330 (N_9330,N_1917,N_3909);
nor U9331 (N_9331,N_3658,N_3002);
nand U9332 (N_9332,N_895,N_3388);
nor U9333 (N_9333,N_2116,N_4799);
and U9334 (N_9334,N_1143,N_4396);
nand U9335 (N_9335,N_3106,N_211);
and U9336 (N_9336,N_1489,N_4250);
nand U9337 (N_9337,N_482,N_4606);
and U9338 (N_9338,N_1415,N_1118);
nor U9339 (N_9339,N_976,N_3410);
nor U9340 (N_9340,N_3466,N_3454);
nor U9341 (N_9341,N_3312,N_1203);
or U9342 (N_9342,N_1839,N_2005);
and U9343 (N_9343,N_1388,N_2189);
nand U9344 (N_9344,N_4183,N_342);
and U9345 (N_9345,N_2078,N_3288);
nand U9346 (N_9346,N_4243,N_9);
and U9347 (N_9347,N_155,N_4184);
and U9348 (N_9348,N_3850,N_1520);
nor U9349 (N_9349,N_3111,N_4381);
nor U9350 (N_9350,N_4865,N_4132);
nand U9351 (N_9351,N_3226,N_160);
nand U9352 (N_9352,N_210,N_3907);
nand U9353 (N_9353,N_2337,N_2569);
and U9354 (N_9354,N_1420,N_3236);
and U9355 (N_9355,N_3386,N_872);
nor U9356 (N_9356,N_2066,N_1210);
nor U9357 (N_9357,N_1500,N_3875);
and U9358 (N_9358,N_3360,N_1761);
or U9359 (N_9359,N_630,N_3342);
and U9360 (N_9360,N_864,N_4637);
nand U9361 (N_9361,N_253,N_1894);
and U9362 (N_9362,N_2560,N_1996);
and U9363 (N_9363,N_773,N_4591);
and U9364 (N_9364,N_3976,N_2016);
or U9365 (N_9365,N_2714,N_2494);
xnor U9366 (N_9366,N_4989,N_1741);
xnor U9367 (N_9367,N_2734,N_4126);
nand U9368 (N_9368,N_402,N_4893);
nand U9369 (N_9369,N_2735,N_2742);
or U9370 (N_9370,N_3188,N_3084);
nand U9371 (N_9371,N_4214,N_4835);
and U9372 (N_9372,N_967,N_3806);
and U9373 (N_9373,N_2620,N_2540);
nand U9374 (N_9374,N_1562,N_2500);
nor U9375 (N_9375,N_51,N_4271);
xnor U9376 (N_9376,N_1743,N_2461);
nor U9377 (N_9377,N_3706,N_66);
nand U9378 (N_9378,N_1789,N_824);
and U9379 (N_9379,N_478,N_42);
xor U9380 (N_9380,N_3276,N_4569);
and U9381 (N_9381,N_1465,N_4807);
nor U9382 (N_9382,N_4283,N_4068);
or U9383 (N_9383,N_2182,N_608);
nand U9384 (N_9384,N_3745,N_4544);
nand U9385 (N_9385,N_545,N_22);
or U9386 (N_9386,N_1138,N_4311);
and U9387 (N_9387,N_1204,N_4801);
nor U9388 (N_9388,N_3630,N_4739);
nor U9389 (N_9389,N_4505,N_2416);
and U9390 (N_9390,N_57,N_1262);
nand U9391 (N_9391,N_4741,N_68);
nand U9392 (N_9392,N_3849,N_3300);
nor U9393 (N_9393,N_4304,N_2824);
nand U9394 (N_9394,N_569,N_160);
or U9395 (N_9395,N_2781,N_4927);
and U9396 (N_9396,N_4475,N_1130);
nand U9397 (N_9397,N_1696,N_1971);
and U9398 (N_9398,N_288,N_884);
xnor U9399 (N_9399,N_4600,N_4012);
and U9400 (N_9400,N_1323,N_2317);
nor U9401 (N_9401,N_317,N_1620);
nand U9402 (N_9402,N_777,N_2627);
and U9403 (N_9403,N_918,N_4333);
and U9404 (N_9404,N_3475,N_2105);
nor U9405 (N_9405,N_2872,N_1205);
or U9406 (N_9406,N_3227,N_3953);
or U9407 (N_9407,N_4683,N_3729);
xor U9408 (N_9408,N_3036,N_843);
nor U9409 (N_9409,N_3179,N_2122);
and U9410 (N_9410,N_2723,N_3615);
and U9411 (N_9411,N_1772,N_986);
or U9412 (N_9412,N_4164,N_1615);
xnor U9413 (N_9413,N_4190,N_3842);
nand U9414 (N_9414,N_1547,N_2946);
xor U9415 (N_9415,N_4341,N_788);
or U9416 (N_9416,N_2877,N_3165);
or U9417 (N_9417,N_1834,N_3628);
xnor U9418 (N_9418,N_1692,N_361);
nor U9419 (N_9419,N_697,N_4269);
or U9420 (N_9420,N_490,N_234);
or U9421 (N_9421,N_1103,N_3615);
and U9422 (N_9422,N_4967,N_3618);
or U9423 (N_9423,N_487,N_2926);
nor U9424 (N_9424,N_3339,N_3095);
nand U9425 (N_9425,N_3889,N_2553);
xor U9426 (N_9426,N_2,N_3317);
nand U9427 (N_9427,N_882,N_91);
and U9428 (N_9428,N_4993,N_445);
or U9429 (N_9429,N_21,N_4708);
xor U9430 (N_9430,N_1635,N_269);
and U9431 (N_9431,N_258,N_708);
and U9432 (N_9432,N_3305,N_342);
nand U9433 (N_9433,N_1319,N_4283);
nand U9434 (N_9434,N_1238,N_1884);
nand U9435 (N_9435,N_4481,N_3143);
or U9436 (N_9436,N_4946,N_2948);
or U9437 (N_9437,N_2035,N_2461);
or U9438 (N_9438,N_3056,N_3404);
nor U9439 (N_9439,N_3267,N_2750);
nand U9440 (N_9440,N_1425,N_3741);
and U9441 (N_9441,N_3184,N_4841);
and U9442 (N_9442,N_3300,N_460);
nor U9443 (N_9443,N_1684,N_4114);
xnor U9444 (N_9444,N_4967,N_4046);
nand U9445 (N_9445,N_1217,N_1704);
nand U9446 (N_9446,N_58,N_2749);
nand U9447 (N_9447,N_4910,N_286);
or U9448 (N_9448,N_2031,N_1894);
nand U9449 (N_9449,N_3139,N_3704);
or U9450 (N_9450,N_2190,N_1864);
and U9451 (N_9451,N_216,N_2657);
nand U9452 (N_9452,N_3217,N_3376);
or U9453 (N_9453,N_4506,N_3188);
nor U9454 (N_9454,N_4599,N_1420);
xnor U9455 (N_9455,N_1483,N_3633);
nor U9456 (N_9456,N_1312,N_1037);
or U9457 (N_9457,N_2430,N_1607);
nand U9458 (N_9458,N_3001,N_3730);
nor U9459 (N_9459,N_2545,N_112);
nor U9460 (N_9460,N_2156,N_4697);
nor U9461 (N_9461,N_4427,N_208);
nand U9462 (N_9462,N_1619,N_4389);
nor U9463 (N_9463,N_1961,N_3621);
nand U9464 (N_9464,N_858,N_4060);
xnor U9465 (N_9465,N_1991,N_2839);
xnor U9466 (N_9466,N_2852,N_3216);
and U9467 (N_9467,N_2999,N_4624);
nor U9468 (N_9468,N_480,N_3856);
nand U9469 (N_9469,N_1539,N_1444);
and U9470 (N_9470,N_1634,N_1078);
nor U9471 (N_9471,N_1361,N_392);
or U9472 (N_9472,N_1621,N_4422);
and U9473 (N_9473,N_3866,N_2398);
nor U9474 (N_9474,N_2946,N_4219);
nand U9475 (N_9475,N_4259,N_2417);
xor U9476 (N_9476,N_2403,N_4109);
nor U9477 (N_9477,N_3797,N_548);
nand U9478 (N_9478,N_1967,N_3509);
and U9479 (N_9479,N_4336,N_3188);
and U9480 (N_9480,N_2392,N_965);
and U9481 (N_9481,N_2755,N_4266);
nor U9482 (N_9482,N_1135,N_3817);
or U9483 (N_9483,N_244,N_309);
or U9484 (N_9484,N_4183,N_4947);
and U9485 (N_9485,N_3866,N_848);
xor U9486 (N_9486,N_1649,N_4117);
nor U9487 (N_9487,N_4000,N_3402);
nand U9488 (N_9488,N_1307,N_3398);
nand U9489 (N_9489,N_4670,N_2859);
nor U9490 (N_9490,N_4238,N_1269);
nor U9491 (N_9491,N_730,N_3401);
and U9492 (N_9492,N_1312,N_151);
nand U9493 (N_9493,N_3135,N_853);
or U9494 (N_9494,N_1994,N_2673);
and U9495 (N_9495,N_540,N_4210);
and U9496 (N_9496,N_4473,N_2421);
nand U9497 (N_9497,N_2162,N_3459);
nand U9498 (N_9498,N_3873,N_1043);
nand U9499 (N_9499,N_1506,N_2274);
nor U9500 (N_9500,N_41,N_2061);
or U9501 (N_9501,N_162,N_1338);
or U9502 (N_9502,N_3942,N_421);
and U9503 (N_9503,N_1791,N_4044);
nand U9504 (N_9504,N_1375,N_2973);
nand U9505 (N_9505,N_642,N_4301);
and U9506 (N_9506,N_4996,N_476);
or U9507 (N_9507,N_1401,N_1280);
and U9508 (N_9508,N_219,N_4866);
nand U9509 (N_9509,N_3714,N_4292);
xnor U9510 (N_9510,N_2940,N_4955);
xor U9511 (N_9511,N_2655,N_3458);
or U9512 (N_9512,N_1219,N_3371);
xor U9513 (N_9513,N_2274,N_2202);
or U9514 (N_9514,N_76,N_1398);
xor U9515 (N_9515,N_2560,N_3371);
nand U9516 (N_9516,N_4484,N_2999);
nor U9517 (N_9517,N_3397,N_1618);
and U9518 (N_9518,N_2712,N_383);
and U9519 (N_9519,N_4897,N_4303);
nor U9520 (N_9520,N_1863,N_4682);
nor U9521 (N_9521,N_3664,N_2535);
xnor U9522 (N_9522,N_4807,N_727);
nand U9523 (N_9523,N_354,N_1779);
nand U9524 (N_9524,N_636,N_3826);
nand U9525 (N_9525,N_4715,N_4875);
and U9526 (N_9526,N_3127,N_2147);
or U9527 (N_9527,N_281,N_1531);
nand U9528 (N_9528,N_2849,N_4675);
nand U9529 (N_9529,N_4890,N_3347);
nand U9530 (N_9530,N_3656,N_4405);
nand U9531 (N_9531,N_540,N_4375);
nand U9532 (N_9532,N_1001,N_4069);
and U9533 (N_9533,N_2755,N_4308);
xor U9534 (N_9534,N_4585,N_1842);
nor U9535 (N_9535,N_1216,N_2870);
nand U9536 (N_9536,N_2658,N_2026);
nor U9537 (N_9537,N_2547,N_3529);
and U9538 (N_9538,N_2645,N_337);
nor U9539 (N_9539,N_2557,N_4802);
nor U9540 (N_9540,N_4084,N_1318);
nor U9541 (N_9541,N_4559,N_2227);
nand U9542 (N_9542,N_453,N_2888);
nand U9543 (N_9543,N_2226,N_486);
nand U9544 (N_9544,N_3362,N_1955);
xnor U9545 (N_9545,N_2499,N_4649);
nor U9546 (N_9546,N_3070,N_855);
xor U9547 (N_9547,N_477,N_3151);
nand U9548 (N_9548,N_557,N_2453);
nand U9549 (N_9549,N_3592,N_741);
or U9550 (N_9550,N_4597,N_2767);
or U9551 (N_9551,N_2634,N_323);
or U9552 (N_9552,N_341,N_3648);
and U9553 (N_9553,N_1488,N_2512);
nor U9554 (N_9554,N_3414,N_631);
and U9555 (N_9555,N_1469,N_2510);
or U9556 (N_9556,N_1257,N_2141);
nor U9557 (N_9557,N_791,N_4710);
xnor U9558 (N_9558,N_4864,N_2173);
or U9559 (N_9559,N_4851,N_2649);
and U9560 (N_9560,N_2013,N_2896);
or U9561 (N_9561,N_3958,N_4638);
or U9562 (N_9562,N_3494,N_2506);
nor U9563 (N_9563,N_4628,N_1605);
and U9564 (N_9564,N_3256,N_4113);
or U9565 (N_9565,N_2419,N_2248);
or U9566 (N_9566,N_4059,N_4474);
nor U9567 (N_9567,N_177,N_2461);
and U9568 (N_9568,N_4240,N_4037);
or U9569 (N_9569,N_1999,N_1734);
nand U9570 (N_9570,N_3674,N_600);
nor U9571 (N_9571,N_4231,N_3449);
and U9572 (N_9572,N_3799,N_299);
nand U9573 (N_9573,N_2845,N_2449);
nand U9574 (N_9574,N_809,N_1546);
nor U9575 (N_9575,N_3808,N_1909);
nand U9576 (N_9576,N_527,N_9);
nor U9577 (N_9577,N_3646,N_1764);
or U9578 (N_9578,N_4838,N_3523);
and U9579 (N_9579,N_1181,N_1799);
nand U9580 (N_9580,N_4051,N_2339);
nor U9581 (N_9581,N_2428,N_3065);
nor U9582 (N_9582,N_505,N_3703);
nor U9583 (N_9583,N_2438,N_3592);
or U9584 (N_9584,N_2492,N_4496);
xnor U9585 (N_9585,N_873,N_2666);
and U9586 (N_9586,N_3761,N_4277);
or U9587 (N_9587,N_4776,N_2881);
or U9588 (N_9588,N_881,N_2854);
or U9589 (N_9589,N_1786,N_3899);
or U9590 (N_9590,N_3025,N_353);
nor U9591 (N_9591,N_4893,N_101);
nor U9592 (N_9592,N_4101,N_1517);
nor U9593 (N_9593,N_1109,N_4689);
xor U9594 (N_9594,N_2351,N_1611);
nor U9595 (N_9595,N_2243,N_2072);
nor U9596 (N_9596,N_3723,N_1079);
nor U9597 (N_9597,N_759,N_131);
and U9598 (N_9598,N_4446,N_2573);
xnor U9599 (N_9599,N_703,N_1589);
or U9600 (N_9600,N_1394,N_451);
nor U9601 (N_9601,N_790,N_2148);
and U9602 (N_9602,N_2124,N_781);
or U9603 (N_9603,N_2358,N_1399);
or U9604 (N_9604,N_1354,N_1743);
nor U9605 (N_9605,N_3264,N_561);
or U9606 (N_9606,N_4858,N_50);
nand U9607 (N_9607,N_4428,N_2773);
or U9608 (N_9608,N_4883,N_1812);
or U9609 (N_9609,N_1334,N_3414);
xor U9610 (N_9610,N_2931,N_1240);
xor U9611 (N_9611,N_858,N_3409);
nor U9612 (N_9612,N_2104,N_4783);
or U9613 (N_9613,N_3274,N_4771);
nand U9614 (N_9614,N_1130,N_3830);
nand U9615 (N_9615,N_622,N_1382);
and U9616 (N_9616,N_1444,N_1092);
or U9617 (N_9617,N_498,N_1885);
or U9618 (N_9618,N_2313,N_1931);
nor U9619 (N_9619,N_2911,N_2102);
nor U9620 (N_9620,N_1765,N_2769);
and U9621 (N_9621,N_1353,N_3363);
or U9622 (N_9622,N_1461,N_1649);
nor U9623 (N_9623,N_3619,N_4004);
nand U9624 (N_9624,N_406,N_2683);
or U9625 (N_9625,N_4387,N_390);
or U9626 (N_9626,N_4376,N_3332);
nand U9627 (N_9627,N_2486,N_4508);
nor U9628 (N_9628,N_2122,N_4715);
nor U9629 (N_9629,N_875,N_417);
or U9630 (N_9630,N_4409,N_2652);
or U9631 (N_9631,N_3753,N_3801);
nor U9632 (N_9632,N_4003,N_1086);
and U9633 (N_9633,N_2775,N_4694);
nor U9634 (N_9634,N_2400,N_3207);
nand U9635 (N_9635,N_1543,N_4066);
nor U9636 (N_9636,N_108,N_2472);
or U9637 (N_9637,N_1040,N_2222);
nor U9638 (N_9638,N_2234,N_3549);
nor U9639 (N_9639,N_1466,N_1442);
or U9640 (N_9640,N_3536,N_4992);
and U9641 (N_9641,N_1845,N_642);
and U9642 (N_9642,N_4191,N_84);
or U9643 (N_9643,N_3367,N_700);
nor U9644 (N_9644,N_4707,N_4669);
nor U9645 (N_9645,N_1406,N_2858);
nor U9646 (N_9646,N_1002,N_1324);
nor U9647 (N_9647,N_349,N_598);
or U9648 (N_9648,N_2145,N_1699);
or U9649 (N_9649,N_371,N_3119);
nor U9650 (N_9650,N_15,N_4607);
and U9651 (N_9651,N_2646,N_277);
or U9652 (N_9652,N_2803,N_3806);
nor U9653 (N_9653,N_3761,N_3480);
or U9654 (N_9654,N_3653,N_3092);
xnor U9655 (N_9655,N_515,N_2526);
nor U9656 (N_9656,N_262,N_142);
nor U9657 (N_9657,N_371,N_2678);
and U9658 (N_9658,N_1951,N_4500);
nor U9659 (N_9659,N_4167,N_4635);
nor U9660 (N_9660,N_3057,N_88);
nand U9661 (N_9661,N_2796,N_4135);
nor U9662 (N_9662,N_1476,N_121);
xor U9663 (N_9663,N_4386,N_3163);
and U9664 (N_9664,N_226,N_4763);
nor U9665 (N_9665,N_3179,N_4013);
and U9666 (N_9666,N_4072,N_2401);
nor U9667 (N_9667,N_2589,N_441);
nand U9668 (N_9668,N_1786,N_3432);
xnor U9669 (N_9669,N_3956,N_4440);
nor U9670 (N_9670,N_2056,N_207);
or U9671 (N_9671,N_2949,N_3920);
or U9672 (N_9672,N_1427,N_3601);
nor U9673 (N_9673,N_1066,N_3320);
nor U9674 (N_9674,N_4279,N_2496);
or U9675 (N_9675,N_4175,N_4956);
or U9676 (N_9676,N_2145,N_3597);
nor U9677 (N_9677,N_3661,N_3144);
and U9678 (N_9678,N_3008,N_4327);
and U9679 (N_9679,N_4023,N_2406);
or U9680 (N_9680,N_1047,N_2229);
or U9681 (N_9681,N_156,N_2884);
or U9682 (N_9682,N_73,N_4587);
nor U9683 (N_9683,N_2344,N_2894);
and U9684 (N_9684,N_2548,N_4932);
or U9685 (N_9685,N_1765,N_364);
nor U9686 (N_9686,N_149,N_4281);
nand U9687 (N_9687,N_2451,N_4928);
and U9688 (N_9688,N_3089,N_2409);
and U9689 (N_9689,N_4974,N_880);
nand U9690 (N_9690,N_1734,N_385);
or U9691 (N_9691,N_2440,N_2672);
or U9692 (N_9692,N_3851,N_1103);
or U9693 (N_9693,N_2131,N_2559);
nor U9694 (N_9694,N_4173,N_1359);
xor U9695 (N_9695,N_313,N_4338);
nand U9696 (N_9696,N_4776,N_785);
and U9697 (N_9697,N_3204,N_2992);
and U9698 (N_9698,N_1574,N_4543);
nand U9699 (N_9699,N_3737,N_4040);
and U9700 (N_9700,N_28,N_152);
xnor U9701 (N_9701,N_2257,N_4013);
and U9702 (N_9702,N_3708,N_4228);
or U9703 (N_9703,N_413,N_884);
or U9704 (N_9704,N_2212,N_3893);
nor U9705 (N_9705,N_2533,N_3018);
and U9706 (N_9706,N_603,N_1893);
nand U9707 (N_9707,N_3853,N_2966);
xnor U9708 (N_9708,N_2064,N_1148);
and U9709 (N_9709,N_4510,N_4595);
and U9710 (N_9710,N_1484,N_4845);
nor U9711 (N_9711,N_1270,N_914);
and U9712 (N_9712,N_24,N_3224);
nand U9713 (N_9713,N_203,N_4821);
nor U9714 (N_9714,N_4446,N_2875);
nor U9715 (N_9715,N_4602,N_4454);
or U9716 (N_9716,N_492,N_1400);
and U9717 (N_9717,N_1229,N_952);
or U9718 (N_9718,N_3667,N_2136);
or U9719 (N_9719,N_3862,N_1137);
xor U9720 (N_9720,N_2622,N_1390);
and U9721 (N_9721,N_1115,N_3989);
and U9722 (N_9722,N_1227,N_2100);
and U9723 (N_9723,N_3534,N_3973);
and U9724 (N_9724,N_3738,N_2886);
xor U9725 (N_9725,N_4258,N_4333);
and U9726 (N_9726,N_2935,N_4707);
nor U9727 (N_9727,N_9,N_860);
and U9728 (N_9728,N_1117,N_4484);
and U9729 (N_9729,N_3630,N_3152);
or U9730 (N_9730,N_1752,N_3188);
and U9731 (N_9731,N_1604,N_2395);
nand U9732 (N_9732,N_1023,N_2651);
or U9733 (N_9733,N_3964,N_1338);
or U9734 (N_9734,N_8,N_2716);
or U9735 (N_9735,N_151,N_1961);
nand U9736 (N_9736,N_3946,N_3745);
nor U9737 (N_9737,N_268,N_4486);
or U9738 (N_9738,N_2232,N_3675);
nand U9739 (N_9739,N_91,N_1183);
nand U9740 (N_9740,N_775,N_2287);
or U9741 (N_9741,N_4312,N_3143);
or U9742 (N_9742,N_4542,N_4954);
nor U9743 (N_9743,N_1727,N_2749);
or U9744 (N_9744,N_136,N_1417);
nor U9745 (N_9745,N_4211,N_2880);
and U9746 (N_9746,N_1049,N_641);
and U9747 (N_9747,N_1944,N_1852);
nor U9748 (N_9748,N_4406,N_177);
nand U9749 (N_9749,N_148,N_1801);
or U9750 (N_9750,N_1962,N_208);
and U9751 (N_9751,N_3365,N_1348);
nor U9752 (N_9752,N_1039,N_4295);
and U9753 (N_9753,N_4307,N_1959);
and U9754 (N_9754,N_92,N_3032);
and U9755 (N_9755,N_804,N_477);
nor U9756 (N_9756,N_3636,N_3908);
and U9757 (N_9757,N_3151,N_1749);
nand U9758 (N_9758,N_1612,N_95);
xor U9759 (N_9759,N_1920,N_4604);
and U9760 (N_9760,N_2146,N_722);
nor U9761 (N_9761,N_4645,N_271);
nand U9762 (N_9762,N_1445,N_4345);
nor U9763 (N_9763,N_3276,N_1667);
and U9764 (N_9764,N_2177,N_2397);
nand U9765 (N_9765,N_4091,N_2315);
or U9766 (N_9766,N_1110,N_569);
or U9767 (N_9767,N_3649,N_4115);
or U9768 (N_9768,N_4912,N_1739);
or U9769 (N_9769,N_2476,N_3729);
and U9770 (N_9770,N_3403,N_4397);
and U9771 (N_9771,N_2181,N_326);
and U9772 (N_9772,N_3030,N_676);
or U9773 (N_9773,N_1554,N_4095);
nor U9774 (N_9774,N_2548,N_2960);
or U9775 (N_9775,N_2309,N_4689);
nor U9776 (N_9776,N_4689,N_3731);
nor U9777 (N_9777,N_2132,N_3107);
nand U9778 (N_9778,N_118,N_1600);
nand U9779 (N_9779,N_1199,N_3705);
nand U9780 (N_9780,N_2668,N_1824);
nor U9781 (N_9781,N_1974,N_1188);
or U9782 (N_9782,N_3638,N_4569);
and U9783 (N_9783,N_4660,N_443);
nor U9784 (N_9784,N_4842,N_1730);
and U9785 (N_9785,N_546,N_10);
xnor U9786 (N_9786,N_1293,N_1947);
nor U9787 (N_9787,N_4648,N_1781);
nand U9788 (N_9788,N_3701,N_630);
and U9789 (N_9789,N_3190,N_2030);
or U9790 (N_9790,N_1671,N_1766);
nand U9791 (N_9791,N_711,N_3540);
and U9792 (N_9792,N_4806,N_4492);
xnor U9793 (N_9793,N_555,N_481);
xor U9794 (N_9794,N_3272,N_606);
or U9795 (N_9795,N_2048,N_1252);
or U9796 (N_9796,N_3314,N_1209);
or U9797 (N_9797,N_2619,N_1175);
or U9798 (N_9798,N_762,N_4428);
or U9799 (N_9799,N_2791,N_3934);
or U9800 (N_9800,N_4101,N_3376);
nor U9801 (N_9801,N_1717,N_4204);
or U9802 (N_9802,N_1377,N_1002);
and U9803 (N_9803,N_599,N_1568);
nor U9804 (N_9804,N_1634,N_4692);
nor U9805 (N_9805,N_3466,N_3644);
nor U9806 (N_9806,N_3886,N_1411);
or U9807 (N_9807,N_1895,N_842);
nor U9808 (N_9808,N_1725,N_1099);
and U9809 (N_9809,N_1920,N_3888);
or U9810 (N_9810,N_3879,N_815);
nand U9811 (N_9811,N_2015,N_2284);
and U9812 (N_9812,N_1716,N_4807);
nor U9813 (N_9813,N_5,N_3606);
nor U9814 (N_9814,N_488,N_1211);
and U9815 (N_9815,N_1710,N_3331);
or U9816 (N_9816,N_2233,N_2131);
and U9817 (N_9817,N_765,N_2921);
or U9818 (N_9818,N_2933,N_2806);
and U9819 (N_9819,N_1971,N_956);
and U9820 (N_9820,N_263,N_4888);
nand U9821 (N_9821,N_3247,N_2576);
xnor U9822 (N_9822,N_2420,N_2199);
and U9823 (N_9823,N_662,N_3390);
or U9824 (N_9824,N_3762,N_1211);
nor U9825 (N_9825,N_4876,N_257);
nand U9826 (N_9826,N_1366,N_2476);
or U9827 (N_9827,N_3543,N_269);
nor U9828 (N_9828,N_4624,N_1269);
nor U9829 (N_9829,N_1737,N_3618);
nor U9830 (N_9830,N_3448,N_3111);
or U9831 (N_9831,N_2630,N_3060);
nand U9832 (N_9832,N_3080,N_521);
nand U9833 (N_9833,N_4736,N_4957);
nor U9834 (N_9834,N_3158,N_3829);
nor U9835 (N_9835,N_2550,N_1516);
nor U9836 (N_9836,N_2952,N_1220);
nand U9837 (N_9837,N_1107,N_4635);
nand U9838 (N_9838,N_3087,N_537);
or U9839 (N_9839,N_2702,N_4173);
nand U9840 (N_9840,N_1613,N_3039);
and U9841 (N_9841,N_2787,N_1637);
and U9842 (N_9842,N_1708,N_3276);
nand U9843 (N_9843,N_685,N_2395);
nor U9844 (N_9844,N_2505,N_1425);
or U9845 (N_9845,N_670,N_1564);
or U9846 (N_9846,N_1282,N_3083);
and U9847 (N_9847,N_804,N_1864);
or U9848 (N_9848,N_3015,N_1299);
or U9849 (N_9849,N_207,N_3512);
or U9850 (N_9850,N_1976,N_2969);
nor U9851 (N_9851,N_4067,N_4456);
nand U9852 (N_9852,N_1545,N_1765);
nor U9853 (N_9853,N_2572,N_4260);
or U9854 (N_9854,N_4722,N_155);
nand U9855 (N_9855,N_1379,N_2690);
nand U9856 (N_9856,N_3540,N_3837);
or U9857 (N_9857,N_2653,N_3551);
nand U9858 (N_9858,N_3871,N_1466);
nor U9859 (N_9859,N_2402,N_1339);
nor U9860 (N_9860,N_3922,N_4865);
nand U9861 (N_9861,N_1625,N_2711);
nor U9862 (N_9862,N_3755,N_3741);
and U9863 (N_9863,N_3225,N_2635);
nand U9864 (N_9864,N_2469,N_642);
nor U9865 (N_9865,N_61,N_4008);
and U9866 (N_9866,N_1890,N_4774);
and U9867 (N_9867,N_1059,N_505);
or U9868 (N_9868,N_4693,N_731);
or U9869 (N_9869,N_2378,N_1589);
and U9870 (N_9870,N_4866,N_3143);
or U9871 (N_9871,N_1023,N_1189);
nand U9872 (N_9872,N_4116,N_2984);
or U9873 (N_9873,N_3704,N_2440);
or U9874 (N_9874,N_4359,N_2645);
or U9875 (N_9875,N_1357,N_2350);
xnor U9876 (N_9876,N_2588,N_3217);
nor U9877 (N_9877,N_1062,N_3714);
nor U9878 (N_9878,N_192,N_4516);
or U9879 (N_9879,N_1059,N_1038);
or U9880 (N_9880,N_2746,N_1319);
nand U9881 (N_9881,N_2095,N_4729);
or U9882 (N_9882,N_3941,N_16);
xor U9883 (N_9883,N_1496,N_4074);
xor U9884 (N_9884,N_1958,N_1846);
or U9885 (N_9885,N_1156,N_4477);
and U9886 (N_9886,N_3747,N_2782);
or U9887 (N_9887,N_3746,N_3134);
nor U9888 (N_9888,N_484,N_2217);
and U9889 (N_9889,N_4505,N_2925);
nand U9890 (N_9890,N_3601,N_4985);
or U9891 (N_9891,N_2738,N_3330);
xor U9892 (N_9892,N_2080,N_1665);
xor U9893 (N_9893,N_3342,N_1383);
or U9894 (N_9894,N_1464,N_2433);
nand U9895 (N_9895,N_1657,N_4997);
nand U9896 (N_9896,N_1607,N_3417);
and U9897 (N_9897,N_2542,N_4213);
nand U9898 (N_9898,N_861,N_1086);
and U9899 (N_9899,N_4737,N_4320);
nor U9900 (N_9900,N_4945,N_2176);
nand U9901 (N_9901,N_4099,N_3311);
nand U9902 (N_9902,N_3077,N_2348);
and U9903 (N_9903,N_1505,N_3907);
nand U9904 (N_9904,N_957,N_3267);
and U9905 (N_9905,N_4680,N_597);
nand U9906 (N_9906,N_3056,N_2587);
nand U9907 (N_9907,N_4535,N_3977);
nor U9908 (N_9908,N_4035,N_3054);
nand U9909 (N_9909,N_1055,N_2848);
nand U9910 (N_9910,N_4329,N_1833);
nor U9911 (N_9911,N_1615,N_4240);
nand U9912 (N_9912,N_3330,N_2764);
or U9913 (N_9913,N_3827,N_3506);
nor U9914 (N_9914,N_4513,N_2498);
and U9915 (N_9915,N_2973,N_65);
nor U9916 (N_9916,N_4219,N_3225);
nor U9917 (N_9917,N_3339,N_4952);
and U9918 (N_9918,N_3219,N_4470);
nand U9919 (N_9919,N_4172,N_3341);
and U9920 (N_9920,N_340,N_600);
nand U9921 (N_9921,N_1707,N_4994);
and U9922 (N_9922,N_2665,N_1234);
and U9923 (N_9923,N_1498,N_905);
or U9924 (N_9924,N_3297,N_3033);
or U9925 (N_9925,N_1622,N_63);
nand U9926 (N_9926,N_1420,N_14);
and U9927 (N_9927,N_2813,N_4405);
xnor U9928 (N_9928,N_4182,N_4703);
or U9929 (N_9929,N_368,N_794);
nand U9930 (N_9930,N_3922,N_2266);
nor U9931 (N_9931,N_1134,N_319);
nor U9932 (N_9932,N_30,N_3238);
or U9933 (N_9933,N_2372,N_3262);
and U9934 (N_9934,N_1672,N_360);
nand U9935 (N_9935,N_740,N_2999);
nor U9936 (N_9936,N_2039,N_2400);
nand U9937 (N_9937,N_2425,N_4112);
or U9938 (N_9938,N_2842,N_3533);
nor U9939 (N_9939,N_115,N_1513);
nor U9940 (N_9940,N_1275,N_86);
xor U9941 (N_9941,N_4394,N_2724);
nand U9942 (N_9942,N_754,N_3174);
or U9943 (N_9943,N_2824,N_3873);
xor U9944 (N_9944,N_4417,N_419);
and U9945 (N_9945,N_3109,N_380);
and U9946 (N_9946,N_2161,N_4548);
or U9947 (N_9947,N_4295,N_685);
or U9948 (N_9948,N_1531,N_4641);
and U9949 (N_9949,N_1486,N_892);
nor U9950 (N_9950,N_808,N_3853);
or U9951 (N_9951,N_2622,N_4780);
nor U9952 (N_9952,N_4819,N_3818);
or U9953 (N_9953,N_2688,N_111);
nand U9954 (N_9954,N_4171,N_2001);
nand U9955 (N_9955,N_4592,N_3772);
nand U9956 (N_9956,N_2507,N_385);
or U9957 (N_9957,N_1761,N_2653);
and U9958 (N_9958,N_912,N_888);
or U9959 (N_9959,N_1642,N_3282);
and U9960 (N_9960,N_3866,N_54);
nand U9961 (N_9961,N_2179,N_3601);
nor U9962 (N_9962,N_1942,N_16);
and U9963 (N_9963,N_2269,N_336);
and U9964 (N_9964,N_4491,N_1427);
or U9965 (N_9965,N_2393,N_210);
nand U9966 (N_9966,N_4561,N_4411);
nor U9967 (N_9967,N_3263,N_4835);
nor U9968 (N_9968,N_704,N_2134);
nor U9969 (N_9969,N_4715,N_4869);
and U9970 (N_9970,N_4642,N_4537);
xor U9971 (N_9971,N_1932,N_1075);
and U9972 (N_9972,N_1658,N_52);
nand U9973 (N_9973,N_3726,N_1558);
and U9974 (N_9974,N_1677,N_2236);
and U9975 (N_9975,N_3807,N_3720);
nor U9976 (N_9976,N_1677,N_3703);
nor U9977 (N_9977,N_3948,N_902);
and U9978 (N_9978,N_2110,N_4593);
nor U9979 (N_9979,N_3780,N_346);
xor U9980 (N_9980,N_592,N_4733);
nand U9981 (N_9981,N_3155,N_813);
nor U9982 (N_9982,N_4040,N_4742);
or U9983 (N_9983,N_3006,N_2313);
nand U9984 (N_9984,N_2340,N_2199);
xor U9985 (N_9985,N_2654,N_2040);
or U9986 (N_9986,N_3904,N_1703);
nand U9987 (N_9987,N_498,N_4006);
and U9988 (N_9988,N_194,N_3882);
and U9989 (N_9989,N_153,N_2755);
and U9990 (N_9990,N_4864,N_2827);
and U9991 (N_9991,N_1000,N_560);
nor U9992 (N_9992,N_1270,N_2478);
or U9993 (N_9993,N_1982,N_3585);
nor U9994 (N_9994,N_3140,N_772);
xor U9995 (N_9995,N_304,N_2477);
or U9996 (N_9996,N_3685,N_520);
nand U9997 (N_9997,N_2814,N_4870);
or U9998 (N_9998,N_4221,N_2516);
xnor U9999 (N_9999,N_2845,N_69);
nor U10000 (N_10000,N_6238,N_9289);
nor U10001 (N_10001,N_7172,N_8869);
xor U10002 (N_10002,N_5409,N_9610);
nor U10003 (N_10003,N_5927,N_7175);
nand U10004 (N_10004,N_8202,N_6495);
or U10005 (N_10005,N_9735,N_7699);
nand U10006 (N_10006,N_9373,N_8461);
nand U10007 (N_10007,N_9452,N_8063);
nor U10008 (N_10008,N_8041,N_6219);
or U10009 (N_10009,N_8401,N_5147);
or U10010 (N_10010,N_5045,N_6532);
or U10011 (N_10011,N_5986,N_7994);
or U10012 (N_10012,N_9974,N_7101);
nor U10013 (N_10013,N_9739,N_5487);
nand U10014 (N_10014,N_8874,N_9169);
or U10015 (N_10015,N_9421,N_9167);
or U10016 (N_10016,N_9302,N_8757);
nand U10017 (N_10017,N_6307,N_7151);
and U10018 (N_10018,N_9328,N_9535);
and U10019 (N_10019,N_5119,N_6394);
nor U10020 (N_10020,N_8037,N_8725);
nor U10021 (N_10021,N_9769,N_6140);
nor U10022 (N_10022,N_5590,N_7763);
nor U10023 (N_10023,N_6712,N_5424);
xor U10024 (N_10024,N_9995,N_6655);
nand U10025 (N_10025,N_6041,N_6286);
or U10026 (N_10026,N_8179,N_5165);
and U10027 (N_10027,N_5386,N_5092);
or U10028 (N_10028,N_8625,N_6874);
and U10029 (N_10029,N_9187,N_8692);
nand U10030 (N_10030,N_7917,N_5219);
and U10031 (N_10031,N_6613,N_9391);
nand U10032 (N_10032,N_7906,N_5889);
nor U10033 (N_10033,N_8711,N_6296);
nand U10034 (N_10034,N_7090,N_6153);
or U10035 (N_10035,N_7998,N_7804);
or U10036 (N_10036,N_8801,N_5922);
xnor U10037 (N_10037,N_5181,N_5442);
nand U10038 (N_10038,N_6233,N_9282);
xnor U10039 (N_10039,N_6312,N_8975);
xor U10040 (N_10040,N_8512,N_7165);
and U10041 (N_10041,N_6830,N_5396);
xor U10042 (N_10042,N_5285,N_7976);
or U10043 (N_10043,N_8288,N_9372);
xnor U10044 (N_10044,N_6886,N_9012);
nand U10045 (N_10045,N_7319,N_8736);
nand U10046 (N_10046,N_7781,N_9973);
and U10047 (N_10047,N_9053,N_6323);
nor U10048 (N_10048,N_9986,N_6272);
nand U10049 (N_10049,N_7690,N_8856);
xnor U10050 (N_10050,N_9587,N_8444);
xor U10051 (N_10051,N_8132,N_9043);
nor U10052 (N_10052,N_6507,N_9180);
nand U10053 (N_10053,N_6487,N_5712);
nor U10054 (N_10054,N_9377,N_5935);
xor U10055 (N_10055,N_6134,N_6771);
nor U10056 (N_10056,N_8561,N_7695);
and U10057 (N_10057,N_8853,N_7223);
and U10058 (N_10058,N_9078,N_7208);
nand U10059 (N_10059,N_9608,N_5497);
xnor U10060 (N_10060,N_9686,N_5527);
nor U10061 (N_10061,N_5914,N_6929);
nand U10062 (N_10062,N_7078,N_6371);
and U10063 (N_10063,N_5979,N_8192);
nor U10064 (N_10064,N_8503,N_8706);
or U10065 (N_10065,N_9114,N_7145);
nand U10066 (N_10066,N_7992,N_9024);
nand U10067 (N_10067,N_6839,N_7665);
nand U10068 (N_10068,N_6401,N_5774);
or U10069 (N_10069,N_7260,N_9611);
nor U10070 (N_10070,N_7150,N_5260);
nand U10071 (N_10071,N_5582,N_7944);
or U10072 (N_10072,N_9358,N_8118);
and U10073 (N_10073,N_8435,N_6722);
xnor U10074 (N_10074,N_8618,N_5891);
and U10075 (N_10075,N_9102,N_9250);
and U10076 (N_10076,N_8762,N_5840);
and U10077 (N_10077,N_6759,N_5944);
xnor U10078 (N_10078,N_8631,N_8871);
and U10079 (N_10079,N_7147,N_5187);
nor U10080 (N_10080,N_6978,N_7636);
and U10081 (N_10081,N_7121,N_6429);
nand U10082 (N_10082,N_7915,N_7740);
xor U10083 (N_10083,N_8732,N_6321);
or U10084 (N_10084,N_6075,N_6826);
nor U10085 (N_10085,N_5311,N_6730);
nor U10086 (N_10086,N_5141,N_5003);
and U10087 (N_10087,N_7959,N_8402);
nor U10088 (N_10088,N_5539,N_6322);
or U10089 (N_10089,N_7603,N_5906);
or U10090 (N_10090,N_6498,N_9301);
nor U10091 (N_10091,N_9014,N_8659);
nor U10092 (N_10092,N_8595,N_8886);
and U10093 (N_10093,N_9305,N_8967);
nor U10094 (N_10094,N_6282,N_7266);
nand U10095 (N_10095,N_9191,N_7157);
nor U10096 (N_10096,N_8388,N_8389);
or U10097 (N_10097,N_6928,N_5619);
or U10098 (N_10098,N_7818,N_6907);
or U10099 (N_10099,N_8252,N_6751);
nor U10100 (N_10100,N_9057,N_7692);
nand U10101 (N_10101,N_6701,N_8877);
nand U10102 (N_10102,N_9704,N_5474);
nand U10103 (N_10103,N_6623,N_6943);
or U10104 (N_10104,N_5959,N_7056);
or U10105 (N_10105,N_8439,N_7517);
and U10106 (N_10106,N_7359,N_7465);
or U10107 (N_10107,N_7573,N_7632);
nor U10108 (N_10108,N_6424,N_9555);
or U10109 (N_10109,N_5751,N_8695);
nand U10110 (N_10110,N_9887,N_8948);
nor U10111 (N_10111,N_7018,N_9784);
and U10112 (N_10112,N_7766,N_6582);
nand U10113 (N_10113,N_9461,N_6392);
nor U10114 (N_10114,N_6865,N_7761);
xor U10115 (N_10115,N_6820,N_9244);
and U10116 (N_10116,N_5307,N_8870);
xor U10117 (N_10117,N_8769,N_6750);
and U10118 (N_10118,N_7430,N_7997);
nand U10119 (N_10119,N_6523,N_9834);
and U10120 (N_10120,N_8065,N_7490);
and U10121 (N_10121,N_8481,N_6368);
nor U10122 (N_10122,N_9032,N_6213);
or U10123 (N_10123,N_5061,N_7032);
xnor U10124 (N_10124,N_6629,N_5476);
or U10125 (N_10125,N_8062,N_7772);
or U10126 (N_10126,N_9891,N_9788);
nand U10127 (N_10127,N_9520,N_9726);
nor U10128 (N_10128,N_9000,N_9249);
nand U10129 (N_10129,N_6534,N_9728);
nor U10130 (N_10130,N_6504,N_8881);
or U10131 (N_10131,N_7015,N_9840);
or U10132 (N_10132,N_7424,N_7829);
and U10133 (N_10133,N_9977,N_6634);
nand U10134 (N_10134,N_8419,N_7969);
or U10135 (N_10135,N_5066,N_7231);
xnor U10136 (N_10136,N_6829,N_6210);
nor U10137 (N_10137,N_9576,N_6700);
and U10138 (N_10138,N_8153,N_9657);
or U10139 (N_10139,N_6996,N_8643);
or U10140 (N_10140,N_9117,N_6345);
xnor U10141 (N_10141,N_7434,N_6185);
or U10142 (N_10142,N_9922,N_6850);
or U10143 (N_10143,N_5067,N_6278);
nand U10144 (N_10144,N_6289,N_7350);
nor U10145 (N_10145,N_6879,N_9062);
nand U10146 (N_10146,N_6451,N_8027);
nor U10147 (N_10147,N_9936,N_9687);
and U10148 (N_10148,N_5559,N_8564);
and U10149 (N_10149,N_7155,N_7860);
nand U10150 (N_10150,N_9496,N_9400);
nor U10151 (N_10151,N_5543,N_7578);
and U10152 (N_10152,N_7677,N_5563);
xnor U10153 (N_10153,N_8640,N_6437);
nor U10154 (N_10154,N_9763,N_6559);
or U10155 (N_10155,N_5975,N_6416);
or U10156 (N_10156,N_9796,N_5659);
and U10157 (N_10157,N_8400,N_9095);
xnor U10158 (N_10158,N_5105,N_6602);
or U10159 (N_10159,N_7510,N_5835);
and U10160 (N_10160,N_8250,N_9124);
or U10161 (N_10161,N_6450,N_6260);
nand U10162 (N_10162,N_9761,N_6363);
and U10163 (N_10163,N_5286,N_6308);
nand U10164 (N_10164,N_8716,N_7331);
or U10165 (N_10165,N_6642,N_7406);
nor U10166 (N_10166,N_9134,N_6957);
and U10167 (N_10167,N_9526,N_6397);
xnor U10168 (N_10168,N_9872,N_7790);
and U10169 (N_10169,N_9516,N_9132);
and U10170 (N_10170,N_9965,N_7412);
or U10171 (N_10171,N_7956,N_8884);
nand U10172 (N_10172,N_9624,N_5369);
and U10173 (N_10173,N_6757,N_7649);
and U10174 (N_10174,N_6939,N_9151);
and U10175 (N_10175,N_7519,N_7030);
and U10176 (N_10176,N_8479,N_9446);
nor U10177 (N_10177,N_8987,N_7035);
nor U10178 (N_10178,N_9765,N_9487);
or U10179 (N_10179,N_9002,N_8607);
or U10180 (N_10180,N_8012,N_7074);
and U10181 (N_10181,N_6250,N_9190);
nor U10182 (N_10182,N_7506,N_5710);
or U10183 (N_10183,N_8827,N_9680);
nor U10184 (N_10184,N_7853,N_9578);
nand U10185 (N_10185,N_8710,N_6804);
and U10186 (N_10186,N_5454,N_5669);
and U10187 (N_10187,N_9262,N_5368);
nand U10188 (N_10188,N_5910,N_6662);
nand U10189 (N_10189,N_7285,N_6935);
or U10190 (N_10190,N_6430,N_5429);
nor U10191 (N_10191,N_8358,N_9617);
nand U10192 (N_10192,N_7064,N_5933);
or U10193 (N_10193,N_7135,N_9842);
or U10194 (N_10194,N_8768,N_7401);
nor U10195 (N_10195,N_7928,N_5724);
nor U10196 (N_10196,N_9628,N_5804);
nor U10197 (N_10197,N_8283,N_7197);
and U10198 (N_10198,N_6197,N_6959);
or U10199 (N_10199,N_8251,N_6998);
nand U10200 (N_10200,N_7258,N_7655);
nor U10201 (N_10201,N_9823,N_9110);
and U10202 (N_10202,N_7820,N_8755);
or U10203 (N_10203,N_7167,N_5276);
and U10204 (N_10204,N_6428,N_7123);
nor U10205 (N_10205,N_6702,N_6968);
nand U10206 (N_10206,N_6431,N_6986);
and U10207 (N_10207,N_6479,N_7572);
or U10208 (N_10208,N_9399,N_8740);
and U10209 (N_10209,N_5166,N_7094);
nor U10210 (N_10210,N_9904,N_8281);
xor U10211 (N_10211,N_9477,N_6654);
xnor U10212 (N_10212,N_8428,N_5788);
nand U10213 (N_10213,N_6180,N_7295);
or U10214 (N_10214,N_9017,N_7974);
nand U10215 (N_10215,N_7732,N_6896);
nand U10216 (N_10216,N_7214,N_9027);
nor U10217 (N_10217,N_8941,N_9253);
nor U10218 (N_10218,N_6698,N_8176);
nor U10219 (N_10219,N_7701,N_6169);
nor U10220 (N_10220,N_8099,N_5142);
or U10221 (N_10221,N_5170,N_7451);
or U10222 (N_10222,N_5988,N_9367);
xnor U10223 (N_10223,N_8248,N_9288);
nor U10224 (N_10224,N_6279,N_6026);
and U10225 (N_10225,N_9085,N_5213);
xnor U10226 (N_10226,N_5231,N_9813);
and U10227 (N_10227,N_5686,N_6739);
nor U10228 (N_10228,N_5981,N_5956);
and U10229 (N_10229,N_9584,N_6135);
nor U10230 (N_10230,N_8072,N_8168);
nor U10231 (N_10231,N_8704,N_8703);
xnor U10232 (N_10232,N_8605,N_7105);
and U10233 (N_10233,N_9385,N_9096);
and U10234 (N_10234,N_7536,N_9232);
xor U10235 (N_10235,N_9615,N_8983);
nor U10236 (N_10236,N_6720,N_5934);
xor U10237 (N_10237,N_5224,N_8196);
and U10238 (N_10238,N_9651,N_8112);
or U10239 (N_10239,N_8623,N_8080);
nand U10240 (N_10240,N_9721,N_7705);
nor U10241 (N_10241,N_7294,N_9456);
or U10242 (N_10242,N_5525,N_5733);
or U10243 (N_10243,N_5691,N_6492);
nand U10244 (N_10244,N_7130,N_9004);
nor U10245 (N_10245,N_9798,N_8847);
or U10246 (N_10246,N_7518,N_8669);
and U10247 (N_10247,N_7179,N_7418);
and U10248 (N_10248,N_6228,N_9465);
or U10249 (N_10249,N_7025,N_6963);
or U10250 (N_10250,N_9979,N_7270);
nand U10251 (N_10251,N_6445,N_5155);
nor U10252 (N_10252,N_8092,N_9355);
nand U10253 (N_10253,N_6987,N_6131);
and U10254 (N_10254,N_7251,N_6932);
and U10255 (N_10255,N_5829,N_6221);
or U10256 (N_10256,N_8645,N_7351);
xor U10257 (N_10257,N_8646,N_6988);
nand U10258 (N_10258,N_9410,N_6982);
or U10259 (N_10259,N_7218,N_7176);
nor U10260 (N_10260,N_9050,N_7762);
and U10261 (N_10261,N_7097,N_8174);
or U10262 (N_10262,N_9749,N_6030);
nor U10263 (N_10263,N_6717,N_7092);
xor U10264 (N_10264,N_8109,N_9360);
or U10265 (N_10265,N_8944,N_6545);
xnor U10266 (N_10266,N_8634,N_5865);
xnor U10267 (N_10267,N_9482,N_5403);
and U10268 (N_10268,N_9571,N_9895);
nor U10269 (N_10269,N_9737,N_8480);
or U10270 (N_10270,N_5360,N_9601);
or U10271 (N_10271,N_5581,N_5878);
nand U10272 (N_10272,N_5843,N_8396);
nand U10273 (N_10273,N_7799,N_6420);
or U10274 (N_10274,N_5925,N_7353);
nor U10275 (N_10275,N_5129,N_8819);
and U10276 (N_10276,N_7600,N_6673);
nor U10277 (N_10277,N_6590,N_7563);
xor U10278 (N_10278,N_9837,N_8806);
and U10279 (N_10279,N_8613,N_5658);
nor U10280 (N_10280,N_6619,N_7012);
and U10281 (N_10281,N_6005,N_5810);
nand U10282 (N_10282,N_5984,N_9406);
and U10283 (N_10283,N_6658,N_8025);
nor U10284 (N_10284,N_7069,N_6367);
xnor U10285 (N_10285,N_6348,N_9785);
nand U10286 (N_10286,N_6123,N_6078);
or U10287 (N_10287,N_7408,N_6147);
nand U10288 (N_10288,N_5894,N_7284);
nand U10289 (N_10289,N_9827,N_6137);
nor U10290 (N_10290,N_8745,N_9097);
or U10291 (N_10291,N_8050,N_8863);
and U10292 (N_10292,N_6014,N_5983);
nor U10293 (N_10293,N_6601,N_5572);
nor U10294 (N_10294,N_5085,N_8758);
and U10295 (N_10295,N_7846,N_8393);
xor U10296 (N_10296,N_7183,N_9800);
or U10297 (N_10297,N_7960,N_7849);
xor U10298 (N_10298,N_7089,N_5973);
nand U10299 (N_10299,N_8495,N_9733);
nor U10300 (N_10300,N_7300,N_7883);
nor U10301 (N_10301,N_9991,N_9336);
or U10302 (N_10302,N_7140,N_6868);
nand U10303 (N_10303,N_5776,N_5480);
nand U10304 (N_10304,N_8384,N_5179);
and U10305 (N_10305,N_7075,N_7946);
nor U10306 (N_10306,N_7831,N_5514);
and U10307 (N_10307,N_7433,N_9158);
and U10308 (N_10308,N_8053,N_6076);
or U10309 (N_10309,N_6090,N_6226);
or U10310 (N_10310,N_5701,N_6257);
nor U10311 (N_10311,N_9778,N_5486);
xor U10312 (N_10312,N_7609,N_9852);
or U10313 (N_10313,N_9600,N_6497);
or U10314 (N_10314,N_6942,N_6218);
or U10315 (N_10315,N_9646,N_5958);
or U10316 (N_10316,N_5274,N_8486);
nor U10317 (N_10317,N_7202,N_8984);
nor U10318 (N_10318,N_7845,N_9801);
xnor U10319 (N_10319,N_7232,N_9150);
or U10320 (N_10320,N_8305,N_8309);
nand U10321 (N_10321,N_9416,N_5867);
or U10322 (N_10322,N_7125,N_7927);
nor U10323 (N_10323,N_5227,N_7228);
or U10324 (N_10324,N_6708,N_6365);
or U10325 (N_10325,N_7488,N_5567);
nand U10326 (N_10326,N_7787,N_7142);
or U10327 (N_10327,N_8318,N_8748);
xor U10328 (N_10328,N_5057,N_8913);
or U10329 (N_10329,N_6885,N_6782);
nor U10330 (N_10330,N_9311,N_7267);
nor U10331 (N_10331,N_6995,N_6755);
and U10332 (N_10332,N_6519,N_9419);
and U10333 (N_10333,N_7085,N_7402);
or U10334 (N_10334,N_7065,N_8160);
nor U10335 (N_10335,N_6593,N_9942);
nor U10336 (N_10336,N_6824,N_8499);
nand U10337 (N_10337,N_9230,N_6570);
or U10338 (N_10338,N_5172,N_8530);
nand U10339 (N_10339,N_8103,N_7100);
and U10340 (N_10340,N_7411,N_7255);
and U10341 (N_10341,N_9672,N_5924);
nand U10342 (N_10342,N_5365,N_7733);
nor U10343 (N_10343,N_9016,N_6087);
and U10344 (N_10344,N_9375,N_8300);
nor U10345 (N_10345,N_9947,N_6356);
and U10346 (N_10346,N_7808,N_6084);
or U10347 (N_10347,N_5071,N_6231);
xor U10348 (N_10348,N_8619,N_9616);
nor U10349 (N_10349,N_7053,N_5535);
nor U10350 (N_10350,N_8514,N_5198);
xnor U10351 (N_10351,N_9116,N_5614);
and U10352 (N_10352,N_5591,N_7843);
and U10353 (N_10353,N_9826,N_5223);
and U10354 (N_10354,N_6423,N_9829);
and U10355 (N_10355,N_6047,N_8846);
nand U10356 (N_10356,N_5348,N_8214);
or U10357 (N_10357,N_6577,N_5941);
and U10358 (N_10358,N_8539,N_5820);
nand U10359 (N_10359,N_6889,N_5717);
nand U10360 (N_10360,N_7187,N_9722);
nor U10361 (N_10361,N_6342,N_5178);
nor U10362 (N_10362,N_6138,N_9314);
and U10363 (N_10363,N_8521,N_9604);
nand U10364 (N_10364,N_9070,N_5662);
or U10365 (N_10365,N_8074,N_6455);
and U10366 (N_10366,N_7200,N_6198);
nor U10367 (N_10367,N_8867,N_9692);
nor U10368 (N_10368,N_6129,N_7014);
or U10369 (N_10369,N_6792,N_9574);
nor U10370 (N_10370,N_9524,N_8782);
and U10371 (N_10371,N_5882,N_8259);
nand U10372 (N_10372,N_7224,N_8845);
nor U10373 (N_10373,N_8190,N_9315);
nand U10374 (N_10374,N_6639,N_7291);
or U10375 (N_10375,N_5714,N_8290);
nor U10376 (N_10376,N_8493,N_6650);
and U10377 (N_10377,N_5915,N_5901);
or U10378 (N_10378,N_7576,N_8154);
xnor U10379 (N_10379,N_9075,N_8900);
nor U10380 (N_10380,N_6770,N_9031);
xnor U10381 (N_10381,N_5097,N_6677);
nand U10382 (N_10382,N_5238,N_5855);
nor U10383 (N_10383,N_9486,N_5897);
or U10384 (N_10384,N_9300,N_9272);
nor U10385 (N_10385,N_8684,N_6491);
nand U10386 (N_10386,N_6391,N_9556);
xor U10387 (N_10387,N_9745,N_5188);
nand U10388 (N_10388,N_8651,N_5040);
or U10389 (N_10389,N_7529,N_9581);
or U10390 (N_10390,N_9590,N_9939);
or U10391 (N_10391,N_5411,N_7467);
nor U10392 (N_10392,N_8377,N_8271);
nand U10393 (N_10393,N_9005,N_8676);
and U10394 (N_10394,N_7770,N_6269);
and U10395 (N_10395,N_8432,N_8322);
or U10396 (N_10396,N_6902,N_9257);
and U10397 (N_10397,N_5090,N_7301);
and U10398 (N_10398,N_8865,N_8232);
or U10399 (N_10399,N_6678,N_7374);
nand U10400 (N_10400,N_8629,N_9656);
or U10401 (N_10401,N_9286,N_5349);
nor U10402 (N_10402,N_6983,N_9369);
nand U10403 (N_10403,N_8714,N_9649);
or U10404 (N_10404,N_7817,N_8126);
and U10405 (N_10405,N_8999,N_6288);
or U10406 (N_10406,N_7011,N_9022);
xor U10407 (N_10407,N_8991,N_6825);
xor U10408 (N_10408,N_8842,N_9488);
or U10409 (N_10409,N_6981,N_6877);
nand U10410 (N_10410,N_9658,N_7269);
or U10411 (N_10411,N_8713,N_8249);
and U10412 (N_10412,N_5235,N_8707);
xor U10413 (N_10413,N_7400,N_5971);
and U10414 (N_10414,N_6775,N_5357);
or U10415 (N_10415,N_8113,N_8262);
and U10416 (N_10416,N_7830,N_6476);
or U10417 (N_10417,N_8333,N_8737);
nand U10418 (N_10418,N_6101,N_8314);
or U10419 (N_10419,N_7582,N_8857);
and U10420 (N_10420,N_7143,N_6275);
or U10421 (N_10421,N_7264,N_9470);
nand U10422 (N_10422,N_5320,N_7347);
nand U10423 (N_10423,N_5985,N_8774);
xnor U10424 (N_10424,N_7814,N_6952);
nand U10425 (N_10425,N_6710,N_7041);
and U10426 (N_10426,N_6999,N_9126);
or U10427 (N_10427,N_5439,N_9631);
nand U10428 (N_10428,N_9238,N_9003);
nor U10429 (N_10429,N_6152,N_9504);
nand U10430 (N_10430,N_9201,N_8641);
xor U10431 (N_10431,N_5594,N_5194);
xnor U10432 (N_10432,N_7245,N_5638);
nor U10433 (N_10433,N_5383,N_6706);
nor U10434 (N_10434,N_8781,N_9933);
and U10435 (N_10435,N_9897,N_6550);
and U10436 (N_10436,N_7807,N_5404);
or U10437 (N_10437,N_7798,N_6991);
nand U10438 (N_10438,N_5435,N_6518);
or U10439 (N_10439,N_9636,N_8586);
nor U10440 (N_10440,N_8224,N_7013);
or U10441 (N_10441,N_6510,N_6227);
nand U10442 (N_10442,N_7464,N_9833);
or U10443 (N_10443,N_5026,N_6796);
or U10444 (N_10444,N_6125,N_9693);
or U10445 (N_10445,N_5881,N_6336);
and U10446 (N_10446,N_7731,N_7233);
and U10447 (N_10447,N_5420,N_7528);
nor U10448 (N_10448,N_6531,N_9293);
xor U10449 (N_10449,N_6766,N_8395);
nand U10450 (N_10450,N_8351,N_6350);
or U10451 (N_10451,N_6823,N_9724);
nor U10452 (N_10452,N_9883,N_9877);
or U10453 (N_10453,N_5158,N_8594);
nand U10454 (N_10454,N_7874,N_7082);
nor U10455 (N_10455,N_9029,N_8778);
nor U10456 (N_10456,N_9888,N_5453);
nor U10457 (N_10457,N_5737,N_6997);
nand U10458 (N_10458,N_5015,N_9677);
xor U10459 (N_10459,N_5526,N_7667);
nor U10460 (N_10460,N_6618,N_6856);
xor U10461 (N_10461,N_8341,N_5347);
and U10462 (N_10462,N_9595,N_7288);
nand U10463 (N_10463,N_8937,N_7254);
or U10464 (N_10464,N_5700,N_8600);
nor U10465 (N_10465,N_7114,N_7141);
nand U10466 (N_10466,N_8963,N_9507);
nand U10467 (N_10467,N_5589,N_5004);
nand U10468 (N_10468,N_9023,N_8054);
and U10469 (N_10469,N_5428,N_6396);
nor U10470 (N_10470,N_9094,N_5018);
and U10471 (N_10471,N_9275,N_7522);
xnor U10472 (N_10472,N_5373,N_8664);
nand U10473 (N_10473,N_8086,N_6351);
nor U10474 (N_10474,N_7635,N_8986);
and U10475 (N_10475,N_8916,N_6164);
and U10476 (N_10476,N_8134,N_6709);
nor U10477 (N_10477,N_9471,N_6054);
nor U10478 (N_10478,N_5391,N_8952);
nor U10479 (N_10479,N_7352,N_9711);
or U10480 (N_10480,N_9810,N_7570);
nand U10481 (N_10481,N_5518,N_5251);
xnor U10482 (N_10482,N_6295,N_7287);
nand U10483 (N_10483,N_9327,N_6229);
and U10484 (N_10484,N_7357,N_9948);
and U10485 (N_10485,N_9673,N_7211);
and U10486 (N_10486,N_7962,N_8279);
nand U10487 (N_10487,N_9350,N_5592);
xnor U10488 (N_10488,N_6714,N_9695);
xnor U10489 (N_10489,N_9639,N_9455);
and U10490 (N_10490,N_7730,N_6297);
nand U10491 (N_10491,N_8811,N_8136);
and U10492 (N_10492,N_9435,N_7813);
or U10493 (N_10493,N_7504,N_9679);
nand U10494 (N_10494,N_8469,N_5718);
xnor U10495 (N_10495,N_5358,N_5337);
and U10496 (N_10496,N_7937,N_6765);
nand U10497 (N_10497,N_8968,N_8839);
and U10498 (N_10498,N_6146,N_9324);
or U10499 (N_10499,N_8719,N_8497);
nor U10500 (N_10500,N_7548,N_8548);
or U10501 (N_10501,N_9824,N_8673);
and U10502 (N_10502,N_7024,N_8728);
nand U10503 (N_10503,N_8143,N_7286);
xor U10504 (N_10504,N_9753,N_9629);
and U10505 (N_10505,N_8862,N_9669);
nand U10506 (N_10506,N_7587,N_5185);
nand U10507 (N_10507,N_7334,N_7736);
nor U10508 (N_10508,N_8875,N_6086);
xnor U10509 (N_10509,N_9514,N_5586);
or U10510 (N_10510,N_9729,N_9719);
xor U10511 (N_10511,N_7745,N_6827);
nand U10512 (N_10512,N_7469,N_7055);
and U10513 (N_10513,N_9873,N_9867);
and U10514 (N_10514,N_8180,N_5886);
or U10515 (N_10515,N_8906,N_5565);
xnor U10516 (N_10516,N_5103,N_5792);
or U10517 (N_10517,N_5600,N_7895);
or U10518 (N_10518,N_7317,N_8810);
and U10519 (N_10519,N_7453,N_8108);
nor U10520 (N_10520,N_5466,N_9153);
or U10521 (N_10521,N_7163,N_5481);
or U10522 (N_10522,N_8546,N_7586);
xnor U10523 (N_10523,N_9685,N_8939);
xnor U10524 (N_10524,N_8814,N_9713);
or U10525 (N_10525,N_8560,N_6969);
nand U10526 (N_10526,N_9340,N_6888);
xor U10527 (N_10527,N_9958,N_5646);
or U10528 (N_10528,N_8285,N_9525);
and U10529 (N_10529,N_9087,N_7973);
nand U10530 (N_10530,N_7458,N_8567);
nand U10531 (N_10531,N_8317,N_5541);
xnor U10532 (N_10532,N_7002,N_9791);
nor U10533 (N_10533,N_7162,N_8922);
nor U10534 (N_10534,N_9061,N_5884);
and U10535 (N_10535,N_7484,N_6154);
or U10536 (N_10536,N_6150,N_5556);
and U10537 (N_10537,N_9540,N_9445);
nand U10538 (N_10538,N_6256,N_5107);
nor U10539 (N_10539,N_5699,N_7460);
and U10540 (N_10540,N_9285,N_9388);
nand U10541 (N_10541,N_5432,N_8630);
nand U10542 (N_10542,N_6790,N_9660);
nor U10543 (N_10543,N_7949,N_8236);
or U10544 (N_10544,N_8148,N_8721);
nand U10545 (N_10545,N_9198,N_5571);
xnor U10546 (N_10546,N_6834,N_8820);
or U10547 (N_10547,N_9381,N_5785);
and U10548 (N_10548,N_8959,N_9296);
and U10549 (N_10549,N_5024,N_6933);
and U10550 (N_10550,N_6494,N_7066);
nor U10551 (N_10551,N_5058,N_5874);
and U10552 (N_10552,N_8107,N_8043);
nor U10553 (N_10553,N_9741,N_9620);
xnor U10554 (N_10554,N_7445,N_5861);
or U10555 (N_10555,N_7207,N_9698);
nand U10556 (N_10556,N_9732,N_9530);
or U10557 (N_10557,N_8459,N_7958);
nor U10558 (N_10558,N_7466,N_6159);
nor U10559 (N_10559,N_8802,N_7702);
or U10560 (N_10560,N_7485,N_8275);
and U10561 (N_10561,N_9270,N_5968);
or U10562 (N_10562,N_9344,N_5176);
or U10563 (N_10563,N_7574,N_8783);
and U10564 (N_10564,N_6182,N_9025);
nand U10565 (N_10565,N_8079,N_9561);
nor U10566 (N_10566,N_9384,N_8312);
nand U10567 (N_10567,N_9093,N_8140);
nand U10568 (N_10568,N_7388,N_5229);
or U10569 (N_10569,N_6326,N_7858);
and U10570 (N_10570,N_5452,N_5374);
or U10571 (N_10571,N_5450,N_5131);
or U10572 (N_10572,N_7354,N_9931);
nand U10573 (N_10573,N_6632,N_8365);
nand U10574 (N_10574,N_9403,N_8151);
and U10575 (N_10575,N_8515,N_6100);
and U10576 (N_10576,N_8018,N_5501);
nand U10577 (N_10577,N_9541,N_5828);
xor U10578 (N_10578,N_7067,N_5832);
or U10579 (N_10579,N_6561,N_9582);
and U10580 (N_10580,N_9923,N_5660);
nor U10581 (N_10581,N_8956,N_8371);
or U10582 (N_10582,N_9007,N_5716);
nor U10583 (N_10583,N_9847,N_9844);
nand U10584 (N_10584,N_6779,N_7678);
xnor U10585 (N_10585,N_8907,N_8212);
nand U10586 (N_10586,N_6370,N_6974);
xnor U10587 (N_10587,N_9131,N_5864);
nor U10588 (N_10588,N_6267,N_5087);
nor U10589 (N_10589,N_7738,N_7806);
nor U10590 (N_10590,N_9474,N_9664);
or U10591 (N_10591,N_8632,N_8088);
nor U10592 (N_10592,N_9483,N_5929);
and U10593 (N_10593,N_8082,N_6028);
nor U10594 (N_10594,N_7326,N_7380);
or U10595 (N_10595,N_8429,N_7910);
nand U10596 (N_10596,N_7365,N_6199);
or U10597 (N_10597,N_8896,N_5627);
and U10598 (N_10598,N_5772,N_8780);
nand U10599 (N_10599,N_6170,N_9952);
or U10600 (N_10600,N_9981,N_7694);
nor U10601 (N_10601,N_5371,N_8293);
and U10602 (N_10602,N_8188,N_6203);
nor U10603 (N_10603,N_5536,N_9212);
and U10604 (N_10604,N_6994,N_9913);
and U10605 (N_10605,N_7021,N_8123);
nand U10606 (N_10606,N_6793,N_6273);
nand U10607 (N_10607,N_9352,N_9076);
nor U10608 (N_10608,N_9041,N_6073);
or U10609 (N_10609,N_6760,N_5351);
xnor U10610 (N_10610,N_7683,N_7339);
xnor U10611 (N_10611,N_9366,N_6626);
or U10612 (N_10612,N_5911,N_7922);
nand U10613 (N_10613,N_5296,N_8193);
nand U10614 (N_10614,N_8122,N_5551);
nand U10615 (N_10615,N_5833,N_5578);
nand U10616 (N_10616,N_9439,N_6255);
and U10617 (N_10617,N_6040,N_8552);
nor U10618 (N_10618,N_8064,N_9794);
xor U10619 (N_10619,N_9310,N_6500);
xor U10620 (N_10620,N_9259,N_5196);
nor U10621 (N_10621,N_5482,N_6093);
and U10622 (N_10622,N_7472,N_9896);
nand U10623 (N_10623,N_8349,N_7110);
and U10624 (N_10624,N_7765,N_8376);
or U10625 (N_10625,N_5610,N_8970);
nor U10626 (N_10626,N_9709,N_5756);
and U10627 (N_10627,N_7782,N_9967);
and U10628 (N_10628,N_6314,N_5082);
or U10629 (N_10629,N_9546,N_6377);
and U10630 (N_10630,N_8966,N_9740);
nor U10631 (N_10631,N_6912,N_7471);
or U10632 (N_10632,N_7450,N_7647);
and U10633 (N_10633,N_9154,N_6379);
xnor U10634 (N_10634,N_7000,N_6206);
nor U10635 (N_10635,N_5096,N_8697);
nor U10636 (N_10636,N_9192,N_9118);
or U10637 (N_10637,N_5342,N_7355);
nand U10638 (N_10638,N_6142,N_7277);
or U10639 (N_10639,N_8242,N_9982);
nand U10640 (N_10640,N_7951,N_7302);
or U10641 (N_10641,N_8045,N_5427);
nand U10642 (N_10642,N_8233,N_9589);
nor U10643 (N_10643,N_6049,N_8751);
nand U10644 (N_10644,N_7386,N_6546);
or U10645 (N_10645,N_7561,N_7703);
or U10646 (N_10646,N_6904,N_6333);
or U10647 (N_10647,N_9962,N_6950);
nor U10648 (N_10648,N_9321,N_9987);
xor U10649 (N_10649,N_6772,N_9790);
nand U10650 (N_10650,N_7366,N_6189);
nor U10651 (N_10651,N_7393,N_8849);
and U10652 (N_10652,N_5498,N_5818);
or U10653 (N_10653,N_9717,N_5455);
nand U10654 (N_10654,N_5506,N_5685);
or U10655 (N_10655,N_9978,N_8296);
and U10656 (N_10656,N_8825,N_6685);
or U10657 (N_10657,N_5345,N_5496);
nand U10658 (N_10658,N_9069,N_5458);
and U10659 (N_10659,N_9538,N_9921);
and U10660 (N_10660,N_8386,N_5749);
nor U10661 (N_10661,N_8020,N_8334);
and U10662 (N_10662,N_7646,N_7396);
nand U10663 (N_10663,N_5936,N_9989);
xor U10664 (N_10664,N_8824,N_6625);
and U10665 (N_10665,N_9060,N_8572);
and U10666 (N_10666,N_7606,N_9752);
xor U10667 (N_10667,N_6174,N_8960);
or U10668 (N_10668,N_7977,N_5588);
nand U10669 (N_10669,N_7749,N_5434);
nand U10670 (N_10670,N_8411,N_9723);
and U10671 (N_10671,N_5011,N_8215);
or U10672 (N_10672,N_7840,N_5042);
nand U10673 (N_10673,N_9049,N_8473);
and U10674 (N_10674,N_5430,N_9809);
or U10675 (N_10675,N_9671,N_9226);
nor U10676 (N_10676,N_6927,N_6205);
or U10677 (N_10677,N_7571,N_9092);
nor U10678 (N_10678,N_8830,N_9104);
or U10679 (N_10679,N_6457,N_6204);
and U10680 (N_10680,N_8243,N_7039);
and U10681 (N_10681,N_6789,N_5938);
and U10682 (N_10682,N_7063,N_6831);
nor U10683 (N_10683,N_6934,N_6120);
nand U10684 (N_10684,N_6543,N_7222);
or U10685 (N_10685,N_8919,N_5550);
or U10686 (N_10686,N_5470,N_9591);
and U10687 (N_10687,N_8124,N_5611);
nor U10688 (N_10688,N_6499,N_6908);
or U10689 (N_10689,N_5900,N_9263);
and U10690 (N_10690,N_7934,N_6989);
and U10691 (N_10691,N_9353,N_8574);
nor U10692 (N_10692,N_6372,N_8220);
nand U10693 (N_10693,N_5384,N_9512);
and U10694 (N_10694,N_8559,N_6148);
and U10695 (N_10695,N_9218,N_8273);
and U10696 (N_10696,N_9554,N_5982);
nand U10697 (N_10697,N_5264,N_7461);
nand U10698 (N_10698,N_9316,N_8369);
and U10699 (N_10699,N_7124,N_8516);
or U10700 (N_10700,N_8158,N_9892);
nand U10701 (N_10701,N_9825,N_9754);
and U10702 (N_10702,N_7675,N_7686);
nand U10703 (N_10703,N_5534,N_7653);
and U10704 (N_10704,N_5693,N_9934);
nor U10705 (N_10705,N_5798,N_7279);
or U10706 (N_10706,N_6688,N_6320);
and U10707 (N_10707,N_5350,N_9331);
or U10708 (N_10708,N_9854,N_5261);
and U10709 (N_10709,N_5634,N_5688);
nand U10710 (N_10710,N_5615,N_9028);
and U10711 (N_10711,N_9777,N_8385);
or U10712 (N_10712,N_6801,N_6327);
and U10713 (N_10713,N_6761,N_8225);
or U10714 (N_10714,N_9665,N_7562);
nor U10715 (N_10715,N_7443,N_9186);
or U10716 (N_10716,N_6664,N_9425);
nor U10717 (N_10717,N_9966,N_8680);
nor U10718 (N_10718,N_5745,N_5191);
or U10719 (N_10719,N_7882,N_7507);
xor U10720 (N_10720,N_7134,N_5327);
or U10721 (N_10721,N_8604,N_7505);
nand U10722 (N_10722,N_8321,N_7979);
or U10723 (N_10723,N_7054,N_6013);
nor U10724 (N_10724,N_8006,N_6029);
and U10725 (N_10725,N_9968,N_9542);
and U10726 (N_10726,N_8142,N_7456);
nor U10727 (N_10727,N_5996,N_8624);
or U10728 (N_10728,N_8994,N_8784);
and U10729 (N_10729,N_5932,N_8487);
nand U10730 (N_10730,N_5402,N_9281);
nand U10731 (N_10731,N_8403,N_5812);
nor U10732 (N_10732,N_7541,N_9946);
or U10733 (N_10733,N_8474,N_5043);
or U10734 (N_10734,N_8039,N_9123);
or U10735 (N_10735,N_6533,N_7391);
nand U10736 (N_10736,N_9348,N_7794);
and U10737 (N_10737,N_5294,N_6551);
or U10738 (N_10738,N_9295,N_7473);
and U10739 (N_10739,N_7212,N_6633);
and U10740 (N_10740,N_9961,N_9236);
nand U10741 (N_10741,N_9156,N_6303);
and U10742 (N_10742,N_5353,N_8023);
and U10743 (N_10743,N_9325,N_6085);
or U10744 (N_10744,N_6704,N_8807);
or U10745 (N_10745,N_8392,N_9553);
or U10746 (N_10746,N_9645,N_6251);
and U10747 (N_10747,N_7865,N_7364);
nor U10748 (N_10748,N_9183,N_9015);
nand U10749 (N_10749,N_8951,N_7892);
nor U10750 (N_10750,N_7654,N_8465);
nor U10751 (N_10751,N_7166,N_5678);
nor U10752 (N_10752,N_6385,N_8120);
or U10753 (N_10753,N_6407,N_7459);
and U10754 (N_10754,N_8301,N_6183);
nor U10755 (N_10755,N_8035,N_8822);
or U10756 (N_10756,N_5449,N_8438);
nand U10757 (N_10757,N_9137,N_8456);
nor U10758 (N_10758,N_9386,N_7957);
nor U10759 (N_10759,N_7158,N_5817);
or U10760 (N_10760,N_8667,N_8235);
nand U10761 (N_10761,N_6315,N_7335);
nor U10762 (N_10762,N_6478,N_6878);
and U10763 (N_10763,N_9609,N_5970);
xor U10764 (N_10764,N_9189,N_9997);
nand U10765 (N_10765,N_5073,N_5068);
nor U10766 (N_10766,N_5960,N_7009);
and U10767 (N_10767,N_6466,N_9181);
xor U10768 (N_10768,N_5508,N_6482);
nand U10769 (N_10769,N_7512,N_7384);
nand U10770 (N_10770,N_9146,N_7205);
or U10771 (N_10771,N_8557,N_6595);
nand U10772 (N_10772,N_5315,N_7637);
or U10773 (N_10773,N_9379,N_5495);
and U10774 (N_10774,N_8973,N_8920);
nand U10775 (N_10775,N_9056,N_5766);
and U10776 (N_10776,N_7378,N_6946);
xor U10777 (N_10777,N_6117,N_5060);
nand U10778 (N_10778,N_5744,N_6965);
nand U10779 (N_10779,N_7247,N_8754);
and U10780 (N_10780,N_7159,N_9046);
xnor U10781 (N_10781,N_7803,N_7854);
nand U10782 (N_10782,N_8742,N_5555);
and U10783 (N_10783,N_8199,N_6697);
nor U10784 (N_10784,N_9742,N_5029);
nor U10785 (N_10785,N_6594,N_5291);
nor U10786 (N_10786,N_5521,N_8085);
nand U10787 (N_10787,N_9984,N_8610);
nand U10788 (N_10788,N_7613,N_7757);
nor U10789 (N_10789,N_5545,N_8563);
nand U10790 (N_10790,N_6910,N_8046);
or U10791 (N_10791,N_7048,N_6645);
nor U10792 (N_10792,N_7113,N_9836);
or U10793 (N_10793,N_8127,N_6427);
and U10794 (N_10794,N_7871,N_6718);
or U10795 (N_10795,N_9774,N_5014);
nor U10796 (N_10796,N_7543,N_8449);
xor U10797 (N_10797,N_6922,N_8207);
nand U10798 (N_10798,N_7714,N_8462);
and U10799 (N_10799,N_7902,N_7988);
nand U10800 (N_10800,N_6188,N_9234);
and U10801 (N_10801,N_5177,N_8988);
nor U10802 (N_10802,N_9994,N_7478);
or U10803 (N_10803,N_8658,N_5576);
nand U10804 (N_10804,N_7850,N_9655);
nor U10805 (N_10805,N_7545,N_8688);
and U10806 (N_10806,N_8379,N_9570);
or U10807 (N_10807,N_7533,N_9793);
nand U10808 (N_10808,N_8570,N_6433);
nor U10809 (N_10809,N_7720,N_7515);
xor U10810 (N_10810,N_8592,N_6815);
or U10811 (N_10811,N_8145,N_5033);
and U10812 (N_10812,N_6876,N_9943);
or U10813 (N_10813,N_9472,N_9757);
nand U10814 (N_10814,N_5753,N_8921);
nand U10815 (N_10815,N_5707,N_8792);
or U10816 (N_10816,N_5821,N_7852);
and U10817 (N_10817,N_6460,N_7309);
and U10818 (N_10818,N_5005,N_7476);
xor U10819 (N_10819,N_9694,N_8933);
nor U10820 (N_10820,N_9193,N_9271);
and U10821 (N_10821,N_7639,N_6008);
or U10822 (N_10822,N_9863,N_7068);
or U10823 (N_10823,N_5811,N_8527);
nor U10824 (N_10824,N_9831,N_8150);
nand U10825 (N_10825,N_9529,N_6454);
and U10826 (N_10826,N_5708,N_7271);
and U10827 (N_10827,N_6742,N_8161);
nand U10828 (N_10828,N_5892,N_7362);
nand U10829 (N_10829,N_6721,N_6895);
xor U10830 (N_10830,N_6241,N_5719);
nand U10831 (N_10831,N_6484,N_6777);
and U10832 (N_10832,N_7426,N_9880);
nand U10833 (N_10833,N_6143,N_9307);
or U10834 (N_10834,N_5182,N_6643);
nor U10835 (N_10835,N_7879,N_9013);
and U10836 (N_10836,N_9727,N_9260);
nand U10837 (N_10837,N_9278,N_5259);
and U10838 (N_10838,N_7876,N_9111);
nor U10839 (N_10839,N_6334,N_6340);
or U10840 (N_10840,N_5604,N_9011);
or U10841 (N_10841,N_6191,N_5053);
and U10842 (N_10842,N_9767,N_8902);
xor U10843 (N_10843,N_8337,N_6465);
or U10844 (N_10844,N_5561,N_7410);
and U10845 (N_10845,N_9412,N_6924);
and U10846 (N_10846,N_8061,N_8513);
and U10847 (N_10847,N_9941,N_8209);
or U10848 (N_10848,N_7923,N_9875);
or U10849 (N_10849,N_7435,N_9105);
nand U10850 (N_10850,N_8965,N_6469);
nand U10851 (N_10851,N_6715,N_6369);
and U10852 (N_10852,N_9972,N_8683);
or U10853 (N_10853,N_7498,N_8566);
and U10854 (N_10854,N_8002,N_7281);
and U10855 (N_10855,N_6694,N_7348);
or U10856 (N_10856,N_6905,N_6338);
or U10857 (N_10857,N_7880,N_5569);
and U10858 (N_10858,N_5030,N_6690);
or U10859 (N_10859,N_5721,N_5731);
xor U10860 (N_10860,N_5244,N_8529);
xnor U10861 (N_10861,N_9937,N_5494);
nand U10862 (N_10862,N_7079,N_8191);
nand U10863 (N_10863,N_7527,N_7499);
xor U10864 (N_10864,N_8934,N_8344);
nor U10865 (N_10865,N_8976,N_9284);
nand U10866 (N_10866,N_6001,N_7729);
xor U10867 (N_10867,N_5412,N_6171);
nor U10868 (N_10868,N_6679,N_8263);
or U10869 (N_10869,N_6133,N_5609);
nand U10870 (N_10870,N_8368,N_6675);
nor U10871 (N_10871,N_9513,N_6217);
nand U10872 (N_10872,N_6558,N_9467);
or U10873 (N_10873,N_9241,N_7204);
and U10874 (N_10874,N_6657,N_6539);
nand U10875 (N_10875,N_5869,N_7131);
nand U10876 (N_10876,N_7028,N_5266);
and U10877 (N_10877,N_5920,N_7708);
nor U10878 (N_10878,N_7715,N_9362);
or U10879 (N_10879,N_8879,N_6842);
nand U10880 (N_10880,N_9605,N_7540);
or U10881 (N_10881,N_6667,N_9103);
xnor U10882 (N_10882,N_9215,N_8075);
or U10883 (N_10883,N_9975,N_8727);
xnor U10884 (N_10884,N_9434,N_9527);
and U10885 (N_10885,N_8203,N_9653);
or U10886 (N_10886,N_5281,N_9857);
or U10887 (N_10887,N_8840,N_5735);
nand U10888 (N_10888,N_5750,N_9498);
or U10889 (N_10889,N_7866,N_5355);
nand U10890 (N_10890,N_8551,N_6835);
or U10891 (N_10891,N_6425,N_9858);
nor U10892 (N_10892,N_9893,N_7967);
nor U10893 (N_10893,N_7810,N_5256);
nand U10894 (N_10894,N_5654,N_7759);
or U10895 (N_10895,N_6738,N_9756);
and U10896 (N_10896,N_9370,N_7789);
nor U10897 (N_10897,N_7640,N_6944);
nand U10898 (N_10898,N_6374,N_9030);
and U10899 (N_10899,N_7724,N_5407);
and U10900 (N_10900,N_8627,N_8001);
xnor U10901 (N_10901,N_6467,N_5715);
nor U10902 (N_10902,N_5504,N_5127);
and U10903 (N_10903,N_8356,N_8568);
or U10904 (N_10904,N_7338,N_6566);
nor U10905 (N_10905,N_7413,N_7815);
and U10906 (N_10906,N_9623,N_8638);
or U10907 (N_10907,N_5106,N_6599);
or U10908 (N_10908,N_9960,N_5484);
nand U10909 (N_10909,N_6403,N_7580);
nor U10910 (N_10910,N_7948,N_6172);
nor U10911 (N_10911,N_7491,N_5675);
nor U10912 (N_10912,N_6883,N_7325);
nand U10913 (N_10913,N_6176,N_5440);
and U10914 (N_10914,N_9720,N_9751);
or U10915 (N_10915,N_7336,N_7930);
nor U10916 (N_10916,N_9398,N_9662);
nand U10917 (N_10917,N_9442,N_7891);
nor U10918 (N_10918,N_6530,N_5195);
xnor U10919 (N_10919,N_5226,N_6016);
nand U10920 (N_10920,N_9334,N_9277);
or U10921 (N_10921,N_9894,N_8343);
nand U10922 (N_10922,N_6373,N_8304);
nor U10923 (N_10923,N_7091,N_9954);
or U10924 (N_10924,N_5942,N_9705);
and U10925 (N_10925,N_5216,N_7711);
nor U10926 (N_10926,N_8137,N_8104);
nand U10927 (N_10927,N_7422,N_6015);
or U10928 (N_10928,N_7760,N_8584);
nor U10929 (N_10929,N_7777,N_6954);
xnor U10930 (N_10930,N_7688,N_6474);
nand U10931 (N_10931,N_6270,N_6094);
nor U10932 (N_10932,N_8908,N_6287);
or U10933 (N_10933,N_9318,N_5485);
and U10934 (N_10934,N_8746,N_5138);
xor U10935 (N_10935,N_9099,N_5796);
nor U10936 (N_10936,N_9042,N_5443);
xor U10937 (N_10937,N_7192,N_9920);
or U10938 (N_10938,N_9229,N_8405);
xnor U10939 (N_10939,N_7670,N_9795);
and U10940 (N_10940,N_5262,N_5532);
and U10941 (N_10941,N_8404,N_7901);
nor U10942 (N_10942,N_8531,N_8282);
nand U10943 (N_10943,N_6592,N_7710);
nor U10944 (N_10944,N_8990,N_9363);
or U10945 (N_10945,N_5665,N_8838);
and U10946 (N_10946,N_8649,N_5573);
xnor U10947 (N_10947,N_8008,N_8331);
nand U10948 (N_10948,N_6971,N_9758);
nand U10949 (N_10949,N_5381,N_8129);
nand U10950 (N_10950,N_5672,N_5601);
nor U10951 (N_10951,N_8506,N_6800);
and U10952 (N_10952,N_6680,N_6352);
or U10953 (N_10953,N_8859,N_8187);
and U10954 (N_10954,N_8267,N_9766);
nor U10955 (N_10955,N_7120,N_8423);
and U10956 (N_10956,N_5372,N_6066);
or U10957 (N_10957,N_6707,N_9361);
xnor U10958 (N_10958,N_9932,N_6149);
nand U10959 (N_10959,N_7077,N_5465);
or U10960 (N_10960,N_5137,N_6562);
or U10961 (N_10961,N_5093,N_9688);
nand U10962 (N_10962,N_9549,N_7057);
nor U10963 (N_10963,N_5477,N_9510);
xor U10964 (N_10964,N_7462,N_7693);
nor U10965 (N_10965,N_7360,N_5243);
nor U10966 (N_10966,N_7397,N_8616);
and U10967 (N_10967,N_5217,N_8165);
nand U10968 (N_10968,N_7614,N_5304);
nor U10969 (N_10969,N_5854,N_8596);
nand U10970 (N_10970,N_8476,N_5334);
nand U10971 (N_10971,N_9308,N_9803);
or U10972 (N_10972,N_5607,N_9953);
or U10973 (N_10973,N_6970,N_6209);
or U10974 (N_10974,N_9157,N_6571);
nand U10975 (N_10975,N_5991,N_5265);
nand U10976 (N_10976,N_9929,N_8169);
or U10977 (N_10977,N_7229,N_9743);
nand U10978 (N_10978,N_5949,N_9691);
or U10979 (N_10979,N_9178,N_9115);
nor U10980 (N_10980,N_7031,N_7704);
nand U10981 (N_10981,N_5747,N_9539);
and U10982 (N_10982,N_5885,N_5628);
nand U10983 (N_10983,N_5271,N_6871);
nor U10984 (N_10984,N_9197,N_5397);
and U10985 (N_10985,N_9034,N_9663);
or U10986 (N_10986,N_6318,N_7888);
nor U10987 (N_10987,N_5425,N_8422);
nor U10988 (N_10988,N_8928,N_5282);
nor U10989 (N_10989,N_8602,N_6061);
and U10990 (N_10990,N_9394,N_7161);
and U10991 (N_10991,N_5778,N_9802);
nand U10992 (N_10992,N_9969,N_5734);
nor U10993 (N_10993,N_6025,N_7894);
or U10994 (N_10994,N_6359,N_6305);
xnor U10995 (N_10995,N_6225,N_6064);
and U10996 (N_10996,N_7802,N_5023);
nand U10997 (N_10997,N_7191,N_8759);
and U10998 (N_10998,N_8320,N_5725);
nand U10999 (N_10999,N_5171,N_8729);
nand U11000 (N_11000,N_6598,N_7836);
xnor U11001 (N_11001,N_6611,N_7785);
nor U11002 (N_11002,N_9378,N_8491);
nor U11003 (N_11003,N_6821,N_7684);
nand U11004 (N_11004,N_7535,N_6361);
nor U11005 (N_11005,N_6857,N_7748);
nand U11006 (N_11006,N_9298,N_9618);
or U11007 (N_11007,N_5978,N_5954);
or U11008 (N_11008,N_8997,N_9065);
nor U11009 (N_11009,N_6832,N_7195);
xor U11010 (N_11010,N_6873,N_7320);
nand U11011 (N_11011,N_9221,N_7523);
xor U11012 (N_11012,N_5193,N_9528);
nand U11013 (N_11013,N_5233,N_6393);
nor U11014 (N_11014,N_6132,N_8162);
nor U11015 (N_11015,N_8362,N_8898);
nor U11016 (N_11016,N_6193,N_5846);
or U11017 (N_11017,N_6786,N_5063);
nand U11018 (N_11018,N_8786,N_9380);
nor U11019 (N_11019,N_7626,N_8504);
and U11020 (N_11020,N_5145,N_9499);
nand U11021 (N_11021,N_5134,N_7431);
nor U11022 (N_11022,N_8772,N_9725);
or U11023 (N_11023,N_8526,N_5078);
and U11024 (N_11024,N_6042,N_8005);
nand U11025 (N_11025,N_9402,N_5997);
nand U11026 (N_11026,N_5801,N_6583);
nand U11027 (N_11027,N_8730,N_5445);
nand U11028 (N_11028,N_8373,N_7630);
nor U11029 (N_11029,N_6962,N_9407);
and U11030 (N_11030,N_7006,N_8244);
nor U11031 (N_11031,N_8731,N_6669);
nand U11032 (N_11032,N_9879,N_6985);
or U11033 (N_11033,N_9396,N_6727);
and U11034 (N_11034,N_6564,N_5436);
or U11035 (N_11035,N_9038,N_9476);
nor U11036 (N_11036,N_8310,N_9246);
xnor U11037 (N_11037,N_9853,N_5214);
xnor U11038 (N_11038,N_7972,N_9755);
and U11039 (N_11039,N_6635,N_8957);
nand U11040 (N_11040,N_9172,N_6417);
or U11041 (N_11041,N_9861,N_8338);
and U11042 (N_11042,N_7480,N_8034);
or U11043 (N_11043,N_8717,N_6244);
nor U11044 (N_11044,N_5617,N_6411);
and U11045 (N_11045,N_9674,N_8375);
and U11046 (N_11046,N_7797,N_5050);
nor U11047 (N_11047,N_7119,N_7070);
nand U11048 (N_11048,N_8797,N_9478);
or U11049 (N_11049,N_8313,N_9543);
or U11050 (N_11050,N_8722,N_5841);
nand U11051 (N_11051,N_7181,N_7154);
nand U11052 (N_11052,N_7755,N_6913);
nand U11053 (N_11053,N_7800,N_8346);
or U11054 (N_11054,N_5367,N_6737);
nand U11055 (N_11055,N_9613,N_7919);
nor U11056 (N_11056,N_6068,N_8914);
nand U11057 (N_11057,N_7627,N_9179);
or U11058 (N_11058,N_6095,N_7516);
nand U11059 (N_11059,N_5540,N_6442);
and U11060 (N_11060,N_6384,N_9797);
and U11061 (N_11061,N_8835,N_5275);
and U11062 (N_11062,N_8457,N_8544);
nand U11063 (N_11063,N_5711,N_7819);
nand U11064 (N_11064,N_7389,N_6268);
nor U11065 (N_11065,N_7315,N_5503);
and U11066 (N_11066,N_5741,N_9265);
nand U11067 (N_11067,N_5632,N_8945);
or U11068 (N_11068,N_8319,N_6489);
or U11069 (N_11069,N_8032,N_8642);
nor U11070 (N_11070,N_5947,N_7682);
nor U11071 (N_11071,N_8458,N_8302);
and U11072 (N_11072,N_8958,N_6398);
nor U11073 (N_11073,N_6386,N_7084);
nor U11074 (N_11074,N_6828,N_6074);
nand U11075 (N_11075,N_5184,N_6178);
nor U11076 (N_11076,N_6341,N_5215);
nand U11077 (N_11077,N_5173,N_5834);
nand U11078 (N_11078,N_8947,N_8554);
or U11079 (N_11079,N_6060,N_8776);
nand U11080 (N_11080,N_9850,N_7995);
and U11081 (N_11081,N_6743,N_6212);
or U11082 (N_11082,N_5999,N_9789);
nor U11083 (N_11083,N_6693,N_6852);
nand U11084 (N_11084,N_5793,N_8167);
nor U11085 (N_11085,N_9368,N_9862);
nand U11086 (N_11086,N_6046,N_8866);
and U11087 (N_11087,N_8222,N_8532);
xor U11088 (N_11088,N_8093,N_7554);
nand U11089 (N_11089,N_7436,N_6898);
xor U11090 (N_11090,N_7132,N_8055);
nand U11091 (N_11091,N_5401,N_5160);
or U11092 (N_11092,N_9051,N_6591);
and U11093 (N_11093,N_6328,N_7634);
nand U11094 (N_11094,N_9517,N_8935);
xnor U11095 (N_11095,N_7116,N_5413);
nor U11096 (N_11096,N_8949,N_8152);
or U11097 (N_11097,N_6733,N_9009);
and U11098 (N_11098,N_8415,N_9475);
nand U11099 (N_11099,N_7108,N_6875);
and U11100 (N_11100,N_8412,N_9196);
nor U11101 (N_11101,N_9780,N_7612);
and U11102 (N_11102,N_7848,N_8665);
or U11103 (N_11103,N_6071,N_7553);
nor U11104 (N_11104,N_7996,N_6977);
nand U11105 (N_11105,N_6052,N_7833);
or U11106 (N_11106,N_9204,N_9382);
nor U11107 (N_11107,N_7666,N_9320);
and U11108 (N_11108,N_9661,N_5019);
nand U11109 (N_11109,N_9551,N_7236);
or U11110 (N_11110,N_9506,N_8084);
nand U11111 (N_11111,N_5652,N_8894);
nand U11112 (N_11112,N_9120,N_5794);
and U11113 (N_11113,N_8077,N_5236);
nand U11114 (N_11114,N_9225,N_5272);
nor U11115 (N_11115,N_7602,N_7925);
and U11116 (N_11116,N_5779,N_9573);
and U11117 (N_11117,N_7425,N_9122);
or U11118 (N_11118,N_5248,N_7838);
or U11119 (N_11119,N_7383,N_5232);
nor U11120 (N_11120,N_5842,N_9479);
nor U11121 (N_11121,N_8226,N_5904);
and U11122 (N_11122,N_7629,N_6538);
nor U11123 (N_11123,N_6597,N_7327);
xor U11124 (N_11124,N_7337,N_6953);
or U11125 (N_11125,N_8166,N_8923);
xor U11126 (N_11126,N_7898,N_5473);
nand U11127 (N_11127,N_9998,N_7642);
xnor U11128 (N_11128,N_8326,N_7043);
or U11129 (N_11129,N_5321,N_9501);
or U11130 (N_11130,N_7982,N_6248);
nand U11131 (N_11131,N_7328,N_5657);
and U11132 (N_11132,N_5065,N_8929);
or U11133 (N_11133,N_5955,N_9444);
nor U11134 (N_11134,N_7862,N_6972);
or U11135 (N_11135,N_5845,N_5240);
nand U11136 (N_11136,N_5021,N_5948);
nand U11137 (N_11137,N_8332,N_6644);
and U11138 (N_11138,N_7081,N_9170);
and U11139 (N_11139,N_6864,N_6246);
nor U11140 (N_11140,N_5848,N_7643);
nand U11141 (N_11141,N_6605,N_9297);
nand U11142 (N_11142,N_5755,N_7743);
xor U11143 (N_11143,N_6638,N_6400);
nand U11144 (N_11144,N_5683,N_8872);
and U11145 (N_11145,N_6012,N_9764);
or U11146 (N_11146,N_8912,N_9572);
nor U11147 (N_11147,N_6293,N_7215);
xnor U11148 (N_11148,N_8698,N_5608);
nor U11149 (N_11149,N_5868,N_5300);
nand U11150 (N_11150,N_5111,N_6955);
xnor U11151 (N_11151,N_9642,N_9359);
nor U11152 (N_11152,N_9885,N_6615);
and U11153 (N_11153,N_6882,N_8739);
nand U11154 (N_11154,N_5822,N_7117);
nand U11155 (N_11155,N_5289,N_6059);
or U11156 (N_11156,N_7329,N_8416);
nor U11157 (N_11157,N_7034,N_5007);
and U11158 (N_11158,N_6812,N_5781);
and U11159 (N_11159,N_8009,N_8682);
and U11160 (N_11160,N_7532,N_6916);
and U11161 (N_11161,N_5990,N_7037);
and U11162 (N_11162,N_9219,N_8266);
nor U11163 (N_11163,N_5290,N_7173);
nand U11164 (N_11164,N_9303,N_5625);
nand U11165 (N_11165,N_5903,N_9731);
and U11166 (N_11166,N_8518,N_6869);
or U11167 (N_11167,N_6155,N_8892);
or U11168 (N_11168,N_6006,N_5513);
nor U11169 (N_11169,N_6300,N_8292);
and U11170 (N_11170,N_7341,N_6967);
nor U11171 (N_11171,N_9980,N_6022);
or U11172 (N_11172,N_5656,N_6395);
and U11173 (N_11173,N_8066,N_7728);
xnor U11174 (N_11174,N_6840,N_9869);
or U11175 (N_11175,N_6686,N_8144);
nand U11176 (N_11176,N_6647,N_8864);
nand U11177 (N_11177,N_5126,N_9577);
and U11178 (N_11178,N_7596,N_7381);
and U11179 (N_11179,N_9634,N_5993);
xnor U11180 (N_11180,N_9098,N_6567);
xor U11181 (N_11181,N_9207,N_6506);
nor U11182 (N_11182,N_6376,N_8448);
nor U11183 (N_11183,N_5757,N_6508);
and U11184 (N_11184,N_9312,N_9492);
or U11185 (N_11185,N_9547,N_7112);
nand U11186 (N_11186,N_8299,N_6362);
nor U11187 (N_11187,N_5205,N_9409);
or U11188 (N_11188,N_8685,N_5389);
or U11189 (N_11189,N_8033,N_8049);
or U11190 (N_11190,N_6736,N_8172);
and U11191 (N_11191,N_8453,N_9876);
nor U11192 (N_11192,N_7073,N_7531);
and U11193 (N_11193,N_9404,N_8622);
or U11194 (N_11194,N_5616,N_6215);
nand U11195 (N_11195,N_6656,N_8081);
or U11196 (N_11196,N_7721,N_5926);
xnor U11197 (N_11197,N_7722,N_7372);
nor U11198 (N_11198,N_5680,N_7511);
nand U11199 (N_11199,N_8489,N_8542);
or U11200 (N_11200,N_8468,N_5456);
nand U11201 (N_11201,N_9632,N_8059);
nand U11202 (N_11202,N_5790,N_8770);
nand U11203 (N_11203,N_7289,N_9493);
nand U11204 (N_11204,N_9945,N_5595);
nand U11205 (N_11205,N_7864,N_5837);
or U11206 (N_11206,N_7868,N_5907);
nor U11207 (N_11207,N_7650,N_6033);
nand U11208 (N_11208,N_6947,N_5183);
xor U11209 (N_11209,N_8443,N_6097);
nor U11210 (N_11210,N_5247,N_5118);
and U11211 (N_11211,N_7622,N_9536);
nor U11212 (N_11212,N_6990,N_7754);
or U11213 (N_11213,N_7394,N_8245);
nand U11214 (N_11214,N_6903,N_5763);
or U11215 (N_11215,N_5246,N_7457);
nor U11216 (N_11216,N_8447,N_8689);
or U11217 (N_11217,N_8340,N_5976);
nand U11218 (N_11218,N_7226,N_6649);
nor U11219 (N_11219,N_6517,N_9730);
and U11220 (N_11220,N_5062,N_8668);
and U11221 (N_11221,N_5331,N_7297);
nor U11222 (N_11222,N_6118,N_9928);
and U11223 (N_11223,N_5280,N_5128);
nand U11224 (N_11224,N_8500,N_9851);
or U11225 (N_11225,N_7071,N_8587);
nand U11226 (N_11226,N_8932,N_6665);
nand U11227 (N_11227,N_8156,N_9335);
and U11228 (N_11228,N_7102,N_6554);
and U11229 (N_11229,N_7676,N_7349);
nor U11230 (N_11230,N_8492,N_7624);
or U11231 (N_11231,N_7194,N_6113);
nor U11232 (N_11232,N_5633,N_7842);
xnor U11233 (N_11233,N_7178,N_9127);
and U11234 (N_11234,N_5000,N_6937);
or U11235 (N_11235,N_9208,N_9557);
or U11236 (N_11236,N_7373,N_6891);
and U11237 (N_11237,N_7631,N_5787);
and U11238 (N_11238,N_9356,N_9926);
xor U11239 (N_11239,N_9462,N_6513);
and U11240 (N_11240,N_8950,N_8889);
and U11241 (N_11241,N_6668,N_6388);
nand U11242 (N_11242,N_9387,N_9819);
nand U11243 (N_11243,N_5263,N_9548);
and U11244 (N_11244,N_5380,N_8723);
nor U11245 (N_11245,N_5268,N_5695);
nand U11246 (N_11246,N_8555,N_9176);
or U11247 (N_11247,N_6607,N_5905);
nand U11248 (N_11248,N_9202,N_9148);
and U11249 (N_11249,N_7897,N_5212);
nor U11250 (N_11250,N_5490,N_7559);
nor U11251 (N_11251,N_6948,N_9911);
nor U11252 (N_11252,N_9108,N_9700);
and U11253 (N_11253,N_5939,N_7713);
nand U11254 (N_11254,N_9080,N_7679);
and U11255 (N_11255,N_7878,N_7253);
xor U11256 (N_11256,N_8324,N_5965);
and U11257 (N_11257,N_8779,N_8763);
nor U11258 (N_11258,N_9365,N_6541);
nand U11259 (N_11259,N_8442,N_8924);
or U11260 (N_11260,N_8213,N_8382);
or U11261 (N_11261,N_8639,N_5702);
and U11262 (N_11262,N_9283,N_6627);
or U11263 (N_11263,N_9563,N_9864);
xnor U11264 (N_11264,N_6608,N_7608);
xor U11265 (N_11265,N_8021,N_5870);
nor U11266 (N_11266,N_9083,N_7812);
or U11267 (N_11267,N_7581,N_5875);
nand U11268 (N_11268,N_9630,N_5302);
and U11269 (N_11269,N_9565,N_6906);
and U11270 (N_11270,N_7438,N_6560);
xnor U11271 (N_11271,N_8347,N_9586);
nor U11272 (N_11272,N_7669,N_5322);
xor U11273 (N_11273,N_8195,N_5732);
xor U11274 (N_11274,N_9890,N_9792);
nand U11275 (N_11275,N_9020,N_6452);
or U11276 (N_11276,N_9287,N_7964);
and U11277 (N_11277,N_5771,N_6211);
and U11278 (N_11278,N_8971,N_8090);
and U11279 (N_11279,N_6915,N_6291);
nor U11280 (N_11280,N_8227,N_8421);
or U11281 (N_11281,N_9866,N_7244);
xnor U11282 (N_11282,N_6271,N_8992);
nor U11283 (N_11283,N_6453,N_9422);
nand U11284 (N_11284,N_5839,N_5809);
and U11285 (N_11285,N_7597,N_7723);
and U11286 (N_11286,N_8844,N_5674);
or U11287 (N_11287,N_5245,N_7968);
nor U11288 (N_11288,N_7947,N_6158);
or U11289 (N_11289,N_9018,N_7775);
nor U11290 (N_11290,N_7268,N_7346);
and U11291 (N_11291,N_5279,N_8831);
nor U11292 (N_11292,N_9063,N_8752);
and U11293 (N_11293,N_7170,N_8460);
or U11294 (N_11294,N_8381,N_7115);
nand U11295 (N_11295,N_5720,N_7872);
or U11296 (N_11296,N_7477,N_9453);
nor U11297 (N_11297,N_5577,N_5114);
or U11298 (N_11298,N_7399,N_5599);
nand U11299 (N_11299,N_6930,N_9086);
and U11300 (N_11300,N_7896,N_9633);
and U11301 (N_11301,N_7671,N_7656);
nor U11302 (N_11302,N_9210,N_6124);
nor U11303 (N_11303,N_6802,N_9008);
and U11304 (N_11304,N_9583,N_6065);
or U11305 (N_11305,N_7660,N_7932);
or U11306 (N_11306,N_8677,N_8598);
nand U11307 (N_11307,N_6062,N_8675);
nand U11308 (N_11308,N_6552,N_5305);
nor U11309 (N_11309,N_5681,N_7489);
or U11310 (N_11310,N_9676,N_9908);
nand U11311 (N_11311,N_7617,N_6671);
and U11312 (N_11312,N_6274,N_6731);
and U11313 (N_11313,N_7706,N_8451);
xor U11314 (N_11314,N_7592,N_8467);
nand U11315 (N_11315,N_6527,N_9121);
and U11316 (N_11316,N_6814,N_7298);
and U11317 (N_11317,N_6409,N_6464);
and U11318 (N_11318,N_8938,N_9222);
nor U11319 (N_11319,N_8812,N_9443);
xor U11320 (N_11320,N_6501,N_9988);
nand U11321 (N_11321,N_8115,N_9531);
nand U11322 (N_11322,N_7368,N_7776);
nor U11323 (N_11323,N_8823,N_6444);
nor U11324 (N_11324,N_6949,N_5899);
or U11325 (N_11325,N_7585,N_8930);
nor U11326 (N_11326,N_5479,N_5333);
nor U11327 (N_11327,N_9635,N_5928);
nand U11328 (N_11328,N_5469,N_5186);
and U11329 (N_11329,N_8042,N_8577);
nor U11330 (N_11330,N_9495,N_5974);
nand U11331 (N_11331,N_5008,N_5027);
nand U11332 (N_11332,N_5112,N_9351);
xor U11333 (N_11333,N_8146,N_9291);
and U11334 (N_11334,N_8363,N_9059);
nand U11335 (N_11335,N_6165,N_9637);
or U11336 (N_11336,N_8553,N_5343);
nor U11337 (N_11337,N_9427,N_5048);
or U11338 (N_11338,N_6387,N_5605);
xnor U11339 (N_11339,N_5972,N_6705);
or U11340 (N_11340,N_6925,N_6408);
nand U11341 (N_11341,N_7991,N_9413);
nand U11342 (N_11342,N_7783,N_8843);
or U11343 (N_11343,N_6031,N_7950);
or U11344 (N_11344,N_7605,N_7432);
nor U11345 (N_11345,N_5859,N_5520);
nor U11346 (N_11346,N_8230,N_9955);
nand U11347 (N_11347,N_5079,N_6088);
and U11348 (N_11348,N_9430,N_6110);
nor U11349 (N_11349,N_6992,N_7242);
and U11350 (N_11350,N_8850,N_8799);
xnor U11351 (N_11351,N_6418,N_8052);
nand U11352 (N_11352,N_8953,N_7259);
nand U11353 (N_11353,N_5507,N_8294);
and U11354 (N_11354,N_5098,N_6596);
xor U11355 (N_11355,N_7201,N_5760);
or U11356 (N_11356,N_6263,N_7376);
and U11357 (N_11357,N_9903,N_8793);
nand U11358 (N_11358,N_7217,N_5051);
nor U11359 (N_11359,N_5593,N_8571);
xor U11360 (N_11360,N_9515,N_7058);
or U11361 (N_11361,N_6672,N_5505);
and U11362 (N_11362,N_5918,N_9558);
nand U11363 (N_11363,N_5250,N_5047);
xor U11364 (N_11364,N_5764,N_5055);
nand U11365 (N_11365,N_8841,N_7796);
and U11366 (N_11366,N_5326,N_7623);
nor U11367 (N_11367,N_7036,N_6836);
nand U11368 (N_11368,N_8357,N_8575);
or U11369 (N_11369,N_6636,N_6470);
and U11370 (N_11370,N_5738,N_9625);
nor U11371 (N_11371,N_7621,N_6589);
and U11372 (N_11372,N_9648,N_9736);
or U11373 (N_11373,N_6841,N_5361);
and U11374 (N_11374,N_6794,N_8693);
and U11375 (N_11375,N_8370,N_6055);
and U11376 (N_11376,N_5940,N_6222);
and U11377 (N_11377,N_5827,N_5123);
and U11378 (N_11378,N_6111,N_7741);
nor U11379 (N_11379,N_8833,N_9855);
or U11380 (N_11380,N_5313,N_6600);
nand U11381 (N_11381,N_7520,N_8048);
or U11382 (N_11382,N_8155,N_7290);
nand U11383 (N_11383,N_9089,N_7569);
nand U11384 (N_11384,N_5366,N_8184);
nor U11385 (N_11385,N_9678,N_7227);
or U11386 (N_11386,N_9647,N_8621);
or U11387 (N_11387,N_6435,N_8940);
or U11388 (N_11388,N_9055,N_5419);
nor U11389 (N_11389,N_7641,N_6141);
or U11390 (N_11390,N_5159,N_6353);
nand U11391 (N_11391,N_8237,N_9874);
or U11392 (N_11392,N_7890,N_6104);
nand U11393 (N_11393,N_9808,N_6247);
nand U11394 (N_11394,N_5544,N_8590);
and U11395 (N_11395,N_9364,N_9491);
nand U11396 (N_11396,N_7221,N_8067);
xor U11397 (N_11397,N_6446,N_8858);
or U11398 (N_11398,N_7446,N_8734);
or U11399 (N_11399,N_5980,N_6588);
or U11400 (N_11400,N_9567,N_5574);
or U11401 (N_11401,N_6563,N_7313);
xor U11402 (N_11402,N_5961,N_8687);
and U11403 (N_11403,N_9466,N_5359);
or U11404 (N_11404,N_7137,N_8785);
and U11405 (N_11405,N_7047,N_6070);
or U11406 (N_11406,N_5762,N_9839);
nor U11407 (N_11407,N_7444,N_7087);
and U11408 (N_11408,N_7963,N_6190);
or U11409 (N_11409,N_9638,N_9433);
nand U11410 (N_11410,N_5130,N_7395);
and U11411 (N_11411,N_5560,N_7494);
nor U11412 (N_11412,N_5267,N_8096);
or U11413 (N_11413,N_9454,N_9956);
nand U11414 (N_11414,N_8173,N_6139);
nand U11415 (N_11415,N_5549,N_5524);
and U11416 (N_11416,N_5512,N_7106);
nand U11417 (N_11417,N_7945,N_5451);
nand U11418 (N_11418,N_7633,N_8891);
or U11419 (N_11419,N_6119,N_5110);
or U11420 (N_11420,N_5895,N_5568);
or U11421 (N_11421,N_7619,N_7452);
xnor U11422 (N_11422,N_8501,N_9976);
nor U11423 (N_11423,N_7744,N_7886);
nor U11424 (N_11424,N_6744,N_7918);
or U11425 (N_11425,N_8206,N_7318);
nand U11426 (N_11426,N_8327,N_6919);
nand U11427 (N_11427,N_7213,N_5410);
nand U11428 (N_11428,N_5104,N_5989);
nor U11429 (N_11429,N_9026,N_7252);
nor U11430 (N_11430,N_6163,N_6112);
nor U11431 (N_11431,N_8578,N_7575);
xor U11432 (N_11432,N_5500,N_6265);
nand U11433 (N_11433,N_7216,N_8954);
and U11434 (N_11434,N_9044,N_6056);
or U11435 (N_11435,N_7771,N_5148);
and U11436 (N_11436,N_9171,N_7022);
nor U11437 (N_11437,N_9072,N_7990);
xor U11438 (N_11438,N_6419,N_5844);
nand U11439 (N_11439,N_8420,N_5643);
nand U11440 (N_11440,N_9458,N_9502);
or U11441 (N_11441,N_6330,N_6764);
or U11442 (N_11442,N_5467,N_5220);
or U11443 (N_11443,N_6768,N_5308);
nand U11444 (N_11444,N_8359,N_6774);
or U11445 (N_11445,N_7076,N_9951);
xor U11446 (N_11446,N_6253,N_8110);
nand U11447 (N_11447,N_9480,N_7052);
nand U11448 (N_11448,N_5826,N_8743);
nand U11449 (N_11449,N_6144,N_6648);
and U11450 (N_11450,N_6441,N_8424);
or U11451 (N_11451,N_8581,N_9992);
and U11452 (N_11452,N_5696,N_9882);
nor U11453 (N_11453,N_7188,N_6846);
or U11454 (N_11454,N_6574,N_6973);
or U11455 (N_11455,N_8111,N_6186);
nor U11456 (N_11456,N_5509,N_5995);
and U11457 (N_11457,N_8955,N_5415);
and U11458 (N_11458,N_9395,N_7756);
and U11459 (N_11459,N_7390,N_8525);
nor U11460 (N_11460,N_8654,N_7940);
nand U11461 (N_11461,N_8303,N_9155);
and U11462 (N_11462,N_6381,N_5640);
nor U11463 (N_11463,N_5597,N_6909);
xor U11464 (N_11464,N_5392,N_6136);
or U11465 (N_11465,N_5211,N_7500);
and U11466 (N_11466,N_7939,N_6941);
nand U11467 (N_11467,N_5089,N_6769);
xnor U11468 (N_11468,N_6220,N_6468);
and U11469 (N_11469,N_6741,N_7040);
xnor U11470 (N_11470,N_6044,N_9907);
or U11471 (N_11471,N_6691,N_7118);
xor U11472 (N_11472,N_8980,N_9346);
or U11473 (N_11473,N_5705,N_6406);
nand U11474 (N_11474,N_8210,N_9033);
nand U11475 (N_11475,N_9100,N_9747);
nand U11476 (N_11476,N_7889,N_5957);
or U11477 (N_11477,N_7828,N_9522);
and U11478 (N_11478,N_6572,N_5395);
and U11479 (N_11479,N_8466,N_6082);
or U11480 (N_11480,N_7855,N_5324);
or U11481 (N_11481,N_7791,N_8256);
xor U11482 (N_11482,N_5252,N_6860);
and U11483 (N_11483,N_5417,N_7811);
or U11484 (N_11484,N_6780,N_8829);
or U11485 (N_11485,N_9881,N_6659);
and U11486 (N_11486,N_7827,N_5668);
and U11487 (N_11487,N_7316,N_5287);
and U11488 (N_11488,N_8636,N_7080);
and U11489 (N_11489,N_9970,N_8789);
xor U11490 (N_11490,N_9274,N_9820);
or U11491 (N_11491,N_8536,N_7503);
nor U11492 (N_11492,N_6893,N_7220);
nor U11493 (N_11493,N_8257,N_9701);
nor U11494 (N_11494,N_6745,N_9304);
or U11495 (N_11495,N_7809,N_5620);
nor U11496 (N_11496,N_7016,N_8418);
or U11497 (N_11497,N_6280,N_5726);
nor U11498 (N_11498,N_9393,N_5873);
or U11499 (N_11499,N_9165,N_6000);
and U11500 (N_11500,N_5883,N_7146);
nand U11501 (N_11501,N_7486,N_5682);
or U11502 (N_11502,N_7249,N_6811);
nor U11503 (N_11503,N_8764,N_8848);
xor U11504 (N_11504,N_6496,N_7716);
or U11505 (N_11505,N_9432,N_6299);
and U11506 (N_11506,N_7725,N_8297);
nand U11507 (N_11507,N_6128,N_8454);
xor U11508 (N_11508,N_5192,N_5623);
nand U11509 (N_11509,N_8287,N_5385);
nor U11510 (N_11510,N_7387,N_5242);
and U11511 (N_11511,N_8013,N_9776);
nand U11512 (N_11512,N_9161,N_8024);
nor U11513 (N_11513,N_6426,N_6242);
nor U11514 (N_11514,N_9322,N_8399);
or U11515 (N_11515,N_7985,N_5117);
and U11516 (N_11516,N_8943,N_7379);
nor U11517 (N_11517,N_6557,N_6514);
nor U11518 (N_11518,N_5806,N_8773);
nor U11519 (N_11519,N_7936,N_8029);
nor U11520 (N_11520,N_7825,N_7989);
xor U11521 (N_11521,N_7753,N_8430);
and U11522 (N_11522,N_5516,N_9959);
and U11523 (N_11523,N_8068,N_5713);
or U11524 (N_11524,N_5663,N_5163);
nand U11525 (N_11525,N_7909,N_5909);
and U11526 (N_11526,N_6683,N_6653);
xor U11527 (N_11527,N_7805,N_6525);
nand U11528 (N_11528,N_7311,N_9313);
xnor U11529 (N_11529,N_9138,N_9168);
xor U11530 (N_11530,N_7126,N_6838);
nand U11531 (N_11531,N_8888,N_5729);
nor U11532 (N_11532,N_9408,N_5046);
nor U11533 (N_11533,N_7107,N_9418);
nand U11534 (N_11534,N_9106,N_7638);
nand U11535 (N_11535,N_5100,N_8917);
nand U11536 (N_11536,N_7734,N_6652);
or U11537 (N_11537,N_8918,N_5122);
and U11538 (N_11538,N_7929,N_7525);
nor U11539 (N_11539,N_8808,N_6434);
or U11540 (N_11540,N_7508,N_6606);
xnor U11541 (N_11541,N_5664,N_6502);
nor U11542 (N_11542,N_9135,N_7193);
and U11543 (N_11543,N_5649,N_8767);
xnor U11544 (N_11544,N_6808,N_6569);
nor U11545 (N_11545,N_5254,N_7673);
and U11546 (N_11546,N_8804,N_5203);
xor U11547 (N_11547,N_9519,N_8060);
nor U11548 (N_11548,N_7648,N_5872);
nand U11549 (N_11549,N_9345,N_9816);
nand U11550 (N_11550,N_9545,N_8098);
nand U11551 (N_11551,N_9254,N_7385);
xor U11552 (N_11552,N_5491,N_5352);
nor U11553 (N_11553,N_7552,N_8562);
nor U11554 (N_11554,N_9748,N_6899);
nor U11555 (N_11555,N_6752,N_8164);
nand U11556 (N_11556,N_8897,N_8270);
xnor U11557 (N_11557,N_7096,N_5587);
nor U11558 (N_11558,N_6936,N_9689);
and U11559 (N_11559,N_7051,N_6019);
nor U11560 (N_11560,N_5823,N_5722);
or U11561 (N_11561,N_6252,N_8626);
nor U11562 (N_11562,N_5448,N_8240);
nor U11563 (N_11563,N_8234,N_5977);
nand U11564 (N_11564,N_7696,N_5437);
or U11565 (N_11565,N_9807,N_7210);
nor U11566 (N_11566,N_8380,N_7769);
nor U11567 (N_11567,N_8720,N_8883);
nor U11568 (N_11568,N_8125,N_9643);
nor U11569 (N_11569,N_6866,N_6360);
or U11570 (N_11570,N_8977,N_6773);
and U11571 (N_11571,N_7822,N_9592);
and U11572 (N_11572,N_5199,N_7138);
and U11573 (N_11573,N_7938,N_8308);
and U11574 (N_11574,N_9641,N_5962);
nor U11575 (N_11575,N_8942,N_7104);
and U11576 (N_11576,N_8289,N_9417);
and U11577 (N_11577,N_7700,N_5390);
xnor U11578 (N_11578,N_8608,N_9437);
or U11579 (N_11579,N_8915,N_9184);
nand U11580 (N_11580,N_6847,N_5694);
or U11581 (N_11581,N_7952,N_8962);
and U11582 (N_11582,N_5645,N_5292);
and U11583 (N_11583,N_8541,N_7534);
nor U11584 (N_11584,N_6711,N_5603);
nor U11585 (N_11585,N_9107,N_6331);
and U11586 (N_11586,N_8617,N_7881);
nor U11587 (N_11587,N_9550,N_5341);
nand U11588 (N_11588,N_7470,N_9401);
nor U11589 (N_11589,N_9696,N_5953);
or U11590 (N_11590,N_6763,N_6646);
nor U11591 (N_11591,N_5462,N_9239);
xor U11592 (N_11592,N_8163,N_7764);
or U11593 (N_11593,N_5293,N_6201);
nand U11594 (N_11594,N_9999,N_6243);
nor U11595 (N_11595,N_7439,N_7008);
nor U11596 (N_11596,N_5156,N_5153);
nor U11597 (N_11597,N_8878,N_9562);
or U11598 (N_11598,N_7547,N_9079);
and U11599 (N_11599,N_8837,N_5635);
nand U11600 (N_11600,N_7427,N_8311);
and U11601 (N_11601,N_7601,N_5471);
or U11602 (N_11602,N_6402,N_7441);
nand U11603 (N_11603,N_5221,N_6945);
nand U11604 (N_11604,N_5671,N_5006);
and U11605 (N_11605,N_5108,N_8834);
xor U11606 (N_11606,N_8455,N_8927);
nor U11607 (N_11607,N_9575,N_8718);
xnor U11608 (N_11608,N_7549,N_6858);
and U11609 (N_11609,N_8360,N_6122);
and U11610 (N_11610,N_8280,N_7539);
or U11611 (N_11611,N_6663,N_7780);
nand U11612 (N_11612,N_8265,N_7616);
nor U11613 (N_11613,N_5200,N_7544);
xnor U11614 (N_11614,N_6621,N_5298);
nor U11615 (N_11615,N_6890,N_6354);
and U11616 (N_11616,N_7345,N_6515);
nand U11617 (N_11617,N_7943,N_8477);
or U11618 (N_11618,N_6017,N_8101);
and U11619 (N_11619,N_8805,N_6586);
and U11620 (N_11620,N_8307,N_8201);
xnor U11621 (N_11621,N_6421,N_7565);
or U11622 (N_11622,N_8178,N_8316);
nor U11623 (N_11623,N_6641,N_7698);
nor U11624 (N_11624,N_8961,N_8911);
nand U11625 (N_11625,N_8339,N_7841);
and U11626 (N_11626,N_9252,N_6023);
nor U11627 (N_11627,N_7276,N_8445);
or U11628 (N_11628,N_6020,N_6848);
or U11629 (N_11629,N_9843,N_6610);
or U11630 (N_11630,N_8258,N_8777);
nand U11631 (N_11631,N_5303,N_6099);
nor U11632 (N_11632,N_7307,N_7557);
nor U11633 (N_11633,N_5777,N_6536);
or U11634 (N_11634,N_6121,N_8057);
xor U11635 (N_11635,N_7156,N_7109);
or U11636 (N_11636,N_9614,N_8593);
nor U11637 (N_11637,N_5038,N_7475);
or U11638 (N_11638,N_9220,N_9273);
and U11639 (N_11639,N_9806,N_7305);
nand U11640 (N_11640,N_5825,N_8836);
or U11641 (N_11641,N_7238,N_5687);
or U11642 (N_11642,N_8073,N_5612);
nand U11643 (N_11643,N_6214,N_6921);
xnor U11644 (N_11644,N_8905,N_8097);
nand U11645 (N_11645,N_8690,N_5382);
xnor U11646 (N_11646,N_6816,N_9566);
nand U11647 (N_11647,N_9481,N_8517);
nand U11648 (N_11648,N_8647,N_7869);
and U11649 (N_11649,N_7407,N_6349);
nand U11650 (N_11650,N_9142,N_5499);
and U11651 (N_11651,N_7483,N_5946);
and U11652 (N_11652,N_5743,N_7752);
nor U11653 (N_11653,N_9666,N_6230);
or U11654 (N_11654,N_6778,N_9559);
or U11655 (N_11655,N_6316,N_9424);
nand U11656 (N_11656,N_5438,N_5919);
nand U11657 (N_11657,N_9552,N_6236);
nor U11658 (N_11658,N_9983,N_5083);
or U11659 (N_11659,N_5606,N_8494);
nand U11660 (N_11660,N_7651,N_8100);
and U11661 (N_11661,N_9309,N_9091);
xnor U11662 (N_11662,N_7086,N_8488);
nor U11663 (N_11663,N_9935,N_8185);
nor U11664 (N_11664,N_7303,N_9856);
xnor U11665 (N_11665,N_5132,N_8925);
and U11666 (N_11666,N_7421,N_8017);
and U11667 (N_11667,N_7428,N_6051);
xor U11668 (N_11668,N_8735,N_5081);
and U11669 (N_11669,N_6443,N_8204);
or U11670 (N_11670,N_7344,N_5207);
or U11671 (N_11671,N_5241,N_6192);
nor U11672 (N_11672,N_9173,N_5952);
nand U11673 (N_11673,N_8434,N_8089);
or U11674 (N_11674,N_6493,N_6332);
or U11675 (N_11675,N_5441,N_5206);
or U11676 (N_11676,N_9195,N_8534);
or U11677 (N_11677,N_8558,N_5168);
or U11678 (N_11678,N_5653,N_8580);
nor U11679 (N_11679,N_5880,N_5377);
and U11680 (N_11680,N_9845,N_8637);
xor U11681 (N_11681,N_9924,N_6034);
nor U11682 (N_11682,N_9654,N_9783);
and U11683 (N_11683,N_5354,N_7681);
nand U11684 (N_11684,N_6719,N_7983);
or U11685 (N_11685,N_6161,N_8582);
or U11686 (N_11686,N_5598,N_8177);
nor U11687 (N_11687,N_8157,N_5056);
nor U11688 (N_11688,N_6389,N_5288);
or U11689 (N_11689,N_6783,N_6628);
or U11690 (N_11690,N_7283,N_7415);
nor U11691 (N_11691,N_5013,N_5124);
nor U11692 (N_11692,N_8410,N_8149);
and U11693 (N_11693,N_5877,N_5283);
nand U11694 (N_11694,N_5408,N_8295);
nand U11695 (N_11695,N_8031,N_6520);
nor U11696 (N_11696,N_5080,N_7577);
and U11697 (N_11697,N_8903,N_7773);
nand U11698 (N_11698,N_5621,N_9251);
xnor U11699 (N_11699,N_5075,N_5378);
nand U11700 (N_11700,N_5679,N_7414);
nor U11701 (N_11701,N_6058,N_5387);
nand U11702 (N_11702,N_5992,N_6092);
and U11703 (N_11703,N_8650,N_8277);
and U11704 (N_11704,N_7495,N_8509);
or U11705 (N_11705,N_9149,N_5768);
nor U11706 (N_11706,N_5144,N_5552);
or U11707 (N_11707,N_5388,N_7873);
nor U11708 (N_11708,N_5444,N_8753);
xor U11709 (N_11709,N_7497,N_9901);
or U11710 (N_11710,N_8121,N_8336);
nor U11711 (N_11711,N_5530,N_5463);
nor U11712 (N_11712,N_6036,N_5301);
and U11713 (N_11713,N_5022,N_6787);
and U11714 (N_11714,N_6855,N_6526);
nand U11715 (N_11715,N_5069,N_9145);
nor U11716 (N_11716,N_5888,N_5813);
or U11717 (N_11717,N_9035,N_5630);
or U11718 (N_11718,N_8298,N_5964);
and U11719 (N_11719,N_9267,N_9949);
or U11720 (N_11720,N_9159,N_6130);
and U11721 (N_11721,N_7455,N_7416);
nor U11722 (N_11722,N_8588,N_8350);
nand U11723 (N_11723,N_7098,N_8726);
nor U11724 (N_11724,N_7555,N_9707);
nand U11725 (N_11725,N_7241,N_6091);
nor U11726 (N_11726,N_5109,N_8413);
nand U11727 (N_11727,N_8007,N_7685);
nor U11728 (N_11728,N_9397,N_8200);
and U11729 (N_11729,N_8070,N_5086);
or U11730 (N_11730,N_9659,N_7225);
or U11731 (N_11731,N_5519,N_9125);
or U11732 (N_11732,N_7293,N_9129);
and U11733 (N_11733,N_8325,N_8484);
nor U11734 (N_11734,N_7709,N_5472);
nor U11735 (N_11735,N_9734,N_6887);
and U11736 (N_11736,N_8681,N_7893);
or U11737 (N_11737,N_6540,N_8425);
nand U11738 (N_11738,N_9006,N_5511);
nor U11739 (N_11739,N_9799,N_7680);
or U11740 (N_11740,N_6027,N_8817);
nand U11741 (N_11741,N_5564,N_5622);
nor U11742 (N_11742,N_8026,N_8417);
nor U11743 (N_11743,N_7899,N_9090);
nor U11744 (N_11744,N_8197,N_6920);
or U11745 (N_11745,N_6414,N_8982);
and U11746 (N_11746,N_6732,N_9830);
nor U11747 (N_11747,N_8533,N_8291);
nor U11748 (N_11748,N_7010,N_5406);
nand U11749 (N_11749,N_8472,N_5488);
and U11750 (N_11750,N_5257,N_8686);
and U11751 (N_11751,N_9047,N_8475);
and U11752 (N_11752,N_7598,N_9240);
xnor U11753 (N_11753,N_5036,N_9337);
and U11754 (N_11754,N_8181,N_6512);
and U11755 (N_11755,N_8979,N_9182);
and U11756 (N_11756,N_5838,N_5533);
nor U11757 (N_11757,N_9228,N_5856);
nand U11758 (N_11758,N_8354,N_9199);
or U11759 (N_11759,N_5963,N_5709);
nand U11760 (N_11760,N_9703,N_8182);
or U11761 (N_11761,N_6050,N_5146);
or U11762 (N_11762,N_6390,N_5169);
or U11763 (N_11763,N_7185,N_7735);
nand U11764 (N_11764,N_6239,N_9037);
nor U11765 (N_11765,N_6729,N_8091);
xnor U11766 (N_11766,N_5858,N_9185);
nand U11767 (N_11767,N_7526,N_9835);
nand U11768 (N_11768,N_9670,N_9716);
and U11769 (N_11769,N_9347,N_7993);
nand U11770 (N_11770,N_6249,N_8904);
and U11771 (N_11771,N_5034,N_7916);
and U11772 (N_11772,N_8615,N_6798);
or U11773 (N_11773,N_5299,N_6505);
xor U11774 (N_11774,N_7538,N_8427);
and U11775 (N_11775,N_6472,N_7262);
or U11776 (N_11776,N_7306,N_7625);
nor U11777 (N_11777,N_7784,N_5330);
or U11778 (N_11778,N_6818,N_6892);
nand U11779 (N_11779,N_5414,N_9036);
nand U11780 (N_11780,N_6004,N_6758);
and U11781 (N_11781,N_6784,N_6485);
and U11782 (N_11782,N_5689,N_9376);
or U11783 (N_11783,N_9684,N_7867);
nor U11784 (N_11784,N_6670,N_6762);
or U11785 (N_11785,N_7292,N_9319);
nor U11786 (N_11786,N_5548,N_5789);
and U11787 (N_11787,N_7509,N_5613);
nor U11788 (N_11788,N_5923,N_5647);
and U11789 (N_11789,N_5830,N_5876);
nand U11790 (N_11790,N_7978,N_8218);
nand U11791 (N_11791,N_6581,N_8537);
and U11792 (N_11792,N_6043,N_7986);
and U11793 (N_11793,N_9460,N_7652);
nor U11794 (N_11794,N_6412,N_5001);
xnor U11795 (N_11795,N_7367,N_9177);
or U11796 (N_11796,N_6524,N_7322);
nor U11797 (N_11797,N_7127,N_7206);
nand U11798 (N_11798,N_6240,N_7174);
nand U11799 (N_11799,N_8873,N_8816);
or U11800 (N_11800,N_5398,N_7620);
and U11801 (N_11801,N_7674,N_6157);
xor U11802 (N_11802,N_8821,N_8217);
and U11803 (N_11803,N_9211,N_9627);
or U11804 (N_11804,N_9708,N_7168);
and U11805 (N_11805,N_5916,N_8882);
or U11806 (N_11806,N_5773,N_9081);
and U11807 (N_11807,N_8520,N_8926);
nand U11808 (N_11808,N_7727,N_8342);
and U11809 (N_11809,N_7859,N_6511);
nand U11810 (N_11810,N_6926,N_7042);
and U11811 (N_11811,N_6603,N_6422);
and U11812 (N_11812,N_9216,N_5394);
nand U11813 (N_11813,N_5399,N_6103);
nor U11814 (N_11814,N_8414,N_8335);
or U11815 (N_11815,N_7847,N_8022);
nor U11816 (N_11816,N_7687,N_8851);
nor U11817 (N_11817,N_9917,N_7330);
and U11818 (N_11818,N_7718,N_8854);
or U11819 (N_11819,N_9859,N_9420);
and U11820 (N_11820,N_6355,N_5222);
nand U11821 (N_11821,N_6175,N_8995);
nor U11822 (N_11822,N_7049,N_5493);
nor U11823 (N_11823,N_6490,N_9112);
or U11824 (N_11824,N_9426,N_6660);
nor U11825 (N_11825,N_8231,N_9084);
and U11826 (N_11826,N_5651,N_5210);
nor U11827 (N_11827,N_7263,N_9532);
xor U11828 (N_11828,N_9505,N_8268);
nand U11829 (N_11829,N_5335,N_8708);
or U11830 (N_11830,N_6748,N_5797);
nand U11831 (N_11831,N_5637,N_6207);
or U11832 (N_11832,N_6089,N_8998);
nor U11833 (N_11833,N_7933,N_5805);
and U11834 (N_11834,N_5987,N_5618);
nand U11835 (N_11835,N_7152,N_6048);
and U11836 (N_11836,N_8044,N_9509);
and U11837 (N_11837,N_6817,N_6072);
nand U11838 (N_11838,N_8803,N_7604);
nand U11839 (N_11839,N_8701,N_6938);
nand U11840 (N_11840,N_9702,N_9822);
nand U11841 (N_11841,N_9268,N_7038);
nand U11842 (N_11842,N_8016,N_9828);
nand U11843 (N_11843,N_9450,N_5421);
nand U11844 (N_11844,N_7824,N_7971);
nand U11845 (N_11845,N_6325,N_5225);
nor U11846 (N_11846,N_7863,N_7198);
or U11847 (N_11847,N_9846,N_6556);
and U11848 (N_11848,N_5531,N_6799);
or U11849 (N_11849,N_6259,N_9447);
or U11850 (N_11850,N_5631,N_5851);
and U11851 (N_11851,N_6127,N_7243);
nand U11852 (N_11852,N_7591,N_9773);
nor U11853 (N_11853,N_5431,N_9343);
and U11854 (N_11854,N_7524,N_9569);
nand U11855 (N_11855,N_8969,N_7941);
or U11856 (N_11856,N_7955,N_6612);
and U11857 (N_11857,N_9341,N_6716);
and U11858 (N_11858,N_7961,N_9464);
nor U11859 (N_11859,N_6575,N_8628);
nor U11860 (N_11860,N_5850,N_6555);
and U11861 (N_11861,N_9900,N_9326);
xnor U11862 (N_11862,N_5253,N_7023);
and U11863 (N_11863,N_7189,N_9760);
nor U11864 (N_11864,N_8003,N_5930);
and U11865 (N_11865,N_9860,N_5101);
and U11866 (N_11866,N_8633,N_8433);
or U11867 (N_11867,N_7420,N_8083);
nor U11868 (N_11868,N_7668,N_5202);
nand U11869 (N_11869,N_5670,N_7502);
nor U11870 (N_11870,N_8437,N_7182);
or U11871 (N_11871,N_8620,N_9602);
xor U11872 (N_11872,N_9294,N_9868);
or U11873 (N_11873,N_7361,N_5336);
nand U11874 (N_11874,N_7296,N_7719);
or U11875 (N_11875,N_6115,N_6302);
xor U11876 (N_11876,N_8880,N_9459);
and U11877 (N_11877,N_8078,N_7835);
xor U11878 (N_11878,N_9957,N_9918);
nand U11879 (N_11879,N_8788,N_8694);
xor U11880 (N_11880,N_5016,N_5370);
nand U11881 (N_11881,N_8272,N_7513);
or U11882 (N_11882,N_8387,N_8556);
and U11883 (N_11883,N_7482,N_8868);
xor U11884 (N_11884,N_8795,N_8014);
xor U11885 (N_11885,N_8306,N_5074);
xnor U11886 (N_11886,N_6339,N_5197);
or U11887 (N_11887,N_8679,N_9805);
and U11888 (N_11888,N_9160,N_7793);
nor U11889 (N_11889,N_7924,N_9597);
or U11890 (N_11890,N_6809,N_9064);
nand U11891 (N_11891,N_8138,N_5329);
or U11892 (N_11892,N_6756,N_7398);
nand U11893 (N_11893,N_5340,N_9985);
nor U11894 (N_11894,N_9223,N_9200);
nor U11895 (N_11895,N_8221,N_8390);
and U11896 (N_11896,N_9619,N_6116);
and U11897 (N_11897,N_6168,N_6224);
and U11898 (N_11898,N_9668,N_5969);
nor U11899 (N_11899,N_6234,N_5125);
and U11900 (N_11900,N_8171,N_8662);
nor U11901 (N_11901,N_9383,N_6285);
xnor U11902 (N_11902,N_7567,N_7839);
or U11903 (N_11903,N_7885,N_5570);
nor U11904 (N_11904,N_6010,N_9484);
or U11905 (N_11905,N_7821,N_6503);
nor U11906 (N_11906,N_9280,N_5553);
nor U11907 (N_11907,N_5295,N_9256);
xor U11908 (N_11908,N_7615,N_7583);
nor U11909 (N_11909,N_8738,N_7568);
nor U11910 (N_11910,N_9349,N_7026);
or U11911 (N_11911,N_8478,N_7083);
nand U11912 (N_11912,N_5765,N_6301);
nor U11913 (N_11913,N_7987,N_8194);
nor U11914 (N_11914,N_5306,N_6399);
nor U11915 (N_11915,N_5032,N_5459);
and U11916 (N_11916,N_5218,N_7887);
and U11917 (N_11917,N_9247,N_5423);
nand U11918 (N_11918,N_8147,N_8205);
or U11919 (N_11919,N_6681,N_6661);
nand U11920 (N_11920,N_5943,N_7033);
xor U11921 (N_11921,N_8139,N_5754);
and U11922 (N_11922,N_8374,N_9697);
nand U11923 (N_11923,N_6976,N_9902);
nand U11924 (N_11924,N_8832,N_8576);
nor U11925 (N_11925,N_9759,N_6335);
and U11926 (N_11926,N_9392,N_9944);
nand U11927 (N_11927,N_8663,N_6918);
xnor U11928 (N_11928,N_5769,N_8502);
nand U11929 (N_11929,N_6807,N_9621);
nand U11930 (N_11930,N_7747,N_9905);
nand U11931 (N_11931,N_6548,N_6475);
nor U11932 (N_11932,N_9927,N_8094);
nor U11933 (N_11933,N_6975,N_6184);
nand U11934 (N_11934,N_5510,N_6961);
xnor U11935 (N_11935,N_5319,N_6181);
and U11936 (N_11936,N_6565,N_5921);
nor U11937 (N_11937,N_9389,N_6813);
or U11938 (N_11938,N_5204,N_6196);
nor U11939 (N_11939,N_7593,N_9436);
and U11940 (N_11940,N_5150,N_5759);
nand U11941 (N_11941,N_5502,N_6516);
nand U11942 (N_11942,N_7611,N_8355);
and U11943 (N_11943,N_8612,N_5012);
nor U11944 (N_11944,N_6880,N_7323);
nand U11945 (N_11945,N_6651,N_5706);
and U11946 (N_11946,N_6795,N_5784);
nand U11947 (N_11947,N_7589,N_8328);
and U11948 (N_11948,N_5704,N_8996);
and U11949 (N_11949,N_7767,N_8678);
xnor U11950 (N_11950,N_9077,N_9770);
nor U11951 (N_11951,N_9269,N_6284);
and U11952 (N_11952,N_5736,N_9224);
nand U11953 (N_11953,N_7975,N_8159);
and U11954 (N_11954,N_6960,N_5898);
xnor U11955 (N_11955,N_5492,N_5673);
nor U11956 (N_11956,N_8441,N_6703);
and U11957 (N_11957,N_7273,N_6584);
or U11958 (N_11958,N_8656,N_7610);
or U11959 (N_11959,N_5284,N_8264);
nand U11960 (N_11960,N_8826,N_9243);
nand U11961 (N_11961,N_7128,N_8585);
or U11962 (N_11962,N_7954,N_6261);
nand U11963 (N_11963,N_8229,N_9811);
xor U11964 (N_11964,N_8496,N_8771);
and U11965 (N_11965,N_6529,N_9930);
and U11966 (N_11966,N_5896,N_5422);
nor U11967 (N_11967,N_8015,N_6747);
and U11968 (N_11968,N_7160,N_7095);
xor U11969 (N_11969,N_8989,N_5375);
xor U11970 (N_11970,N_7044,N_7304);
and U11971 (N_11971,N_5596,N_6378);
or U11972 (N_11972,N_7920,N_5629);
xnor U11973 (N_11973,N_9775,N_5059);
and U11974 (N_11974,N_7661,N_8211);
and U11975 (N_11975,N_9415,N_7274);
and U11976 (N_11976,N_5044,N_8505);
xor U11977 (N_11977,N_6151,N_7750);
nor U11978 (N_11978,N_5273,N_5162);
nand U11979 (N_11979,N_9511,N_9101);
nor U11980 (N_11980,N_6382,N_8431);
and U11981 (N_11981,N_9568,N_6162);
nor U11982 (N_11982,N_6776,N_5174);
xnor U11983 (N_11983,N_9166,N_5077);
nand U11984 (N_11984,N_6438,N_7177);
nand U11985 (N_11985,N_9405,N_6614);
and U11986 (N_11986,N_8583,N_5585);
nor U11987 (N_11987,N_9109,N_6861);
nor U11988 (N_11988,N_5489,N_5994);
or U11989 (N_11989,N_5602,N_6810);
xor U11990 (N_11990,N_9203,N_7442);
and U11991 (N_11991,N_5808,N_7093);
nand U11992 (N_11992,N_6585,N_9914);
nand U11993 (N_11993,N_9235,N_7061);
and U11994 (N_11994,N_5278,N_5230);
and U11995 (N_11995,N_7657,N_7856);
or U11996 (N_11996,N_8978,N_5644);
xor U11997 (N_11997,N_8766,N_7707);
nand U11998 (N_11998,N_7375,N_9886);
xor U11999 (N_11999,N_6037,N_5228);
xnor U12000 (N_12000,N_5189,N_7664);
nor U12001 (N_12001,N_8756,N_9650);
and U12002 (N_12002,N_6684,N_8591);
xor U12003 (N_12003,N_9175,N_8239);
or U12004 (N_12004,N_9865,N_5475);
and U12005 (N_12005,N_6867,N_5234);
or U12006 (N_12006,N_8573,N_9141);
nor U12007 (N_12007,N_9718,N_6509);
and U12008 (N_12008,N_9245,N_9054);
and U12009 (N_12009,N_5538,N_6749);
xnor U12010 (N_12010,N_6145,N_5676);
or U12011 (N_12011,N_8887,N_5064);
nand U12012 (N_12012,N_7966,N_7496);
and U12013 (N_12013,N_6309,N_9681);
nand U12014 (N_12014,N_6413,N_6347);
nand U12015 (N_12015,N_9738,N_6311);
or U12016 (N_12016,N_7029,N_7246);
or U12017 (N_12017,N_9066,N_5624);
nand U12018 (N_12018,N_6258,N_5684);
and U12019 (N_12019,N_9411,N_7926);
and U12020 (N_12020,N_7658,N_8114);
nor U12021 (N_12021,N_5376,N_8744);
and U12022 (N_12022,N_6578,N_7004);
nor U12023 (N_12023,N_8809,N_8852);
nor U12024 (N_12024,N_6009,N_7111);
nand U12025 (N_12025,N_6993,N_9878);
or U12026 (N_12026,N_9996,N_7148);
or U12027 (N_12027,N_8861,N_8528);
and U12028 (N_12028,N_5690,N_9209);
nand U12029 (N_12029,N_9163,N_5393);
or U12030 (N_12030,N_6616,N_8909);
or U12031 (N_12031,N_5249,N_9001);
or U12032 (N_12032,N_8247,N_5966);
and U12033 (N_12033,N_5728,N_6797);
and U12034 (N_12034,N_8011,N_5115);
nand U12035 (N_12035,N_8398,N_8069);
and U12036 (N_12036,N_9188,N_8189);
nor U12037 (N_12037,N_6844,N_7778);
xnor U12038 (N_12038,N_6024,N_5317);
nand U12039 (N_12039,N_7377,N_8051);
or U12040 (N_12040,N_6463,N_8855);
nor U12041 (N_12041,N_8910,N_5277);
xor U12042 (N_12042,N_8601,N_5931);
nor U12043 (N_12043,N_6254,N_6114);
or U12044 (N_12044,N_8589,N_8652);
nor U12045 (N_12045,N_8087,N_8028);
and U12046 (N_12046,N_5849,N_7659);
or U12047 (N_12047,N_5041,N_9489);
xnor U12048 (N_12048,N_5483,N_9128);
and U12049 (N_12049,N_5879,N_8901);
and U12050 (N_12050,N_5786,N_8794);
nand U12051 (N_12051,N_5542,N_8936);
and U12052 (N_12052,N_7774,N_7607);
nor U12053 (N_12053,N_9715,N_9910);
or U12054 (N_12054,N_5037,N_7474);
nor U12055 (N_12055,N_5655,N_9815);
or U12056 (N_12056,N_6964,N_5816);
or U12057 (N_12057,N_9606,N_6439);
nand U12058 (N_12058,N_7492,N_9414);
or U12059 (N_12059,N_8058,N_8524);
nor U12060 (N_12060,N_5102,N_6845);
or U12061 (N_12061,N_7870,N_7122);
and U12062 (N_12062,N_6456,N_8702);
nor U12063 (N_12063,N_9667,N_5167);
xnor U12064 (N_12064,N_6216,N_5890);
xor U12065 (N_12065,N_5332,N_7001);
or U12066 (N_12066,N_5076,N_9299);
and U12067 (N_12067,N_9333,N_6695);
nand U12068 (N_12068,N_5400,N_7999);
nand U12069 (N_12069,N_6901,N_8700);
xor U12070 (N_12070,N_7537,N_5316);
or U12071 (N_12071,N_7072,N_9342);
nor U12072 (N_12072,N_9544,N_9950);
xor U12073 (N_12073,N_9762,N_5461);
or U12074 (N_12074,N_9585,N_6724);
nor U12075 (N_12075,N_7851,N_9431);
and U12076 (N_12076,N_9644,N_9323);
nand U12077 (N_12077,N_8183,N_6179);
nand U12078 (N_12078,N_6542,N_6870);
and U12079 (N_12079,N_7556,N_9071);
nor U12080 (N_12080,N_6980,N_9497);
or U12081 (N_12081,N_9537,N_5528);
or U12082 (N_12082,N_8705,N_6859);
and U12083 (N_12083,N_7449,N_9139);
or U12084 (N_12084,N_8219,N_6480);
nor U12085 (N_12085,N_8255,N_6473);
and U12086 (N_12086,N_6687,N_5799);
nor U12087 (N_12087,N_7409,N_6713);
xor U12088 (N_12088,N_9915,N_6803);
and U12089 (N_12089,N_7257,N_9494);
or U12090 (N_12090,N_8019,N_6854);
nand U12091 (N_12091,N_6083,N_8490);
nor U12092 (N_12092,N_9889,N_6357);
nand U12093 (N_12093,N_7392,N_6923);
nand U12094 (N_12094,N_5433,N_6911);
nor U12095 (N_12095,N_6753,N_8974);
nor U12096 (N_12096,N_8141,N_8260);
nor U12097 (N_12097,N_8353,N_6081);
nor U12098 (N_12098,N_8131,N_9603);
nor U12099 (N_12099,N_7237,N_7908);
nand U12100 (N_12100,N_8117,N_7834);
and U12101 (N_12101,N_5478,N_7758);
and U12102 (N_12102,N_9523,N_5028);
xor U12103 (N_12103,N_5339,N_7363);
nor U12104 (N_12104,N_8352,N_5099);
nor U12105 (N_12105,N_8791,N_8348);
nand U12106 (N_12106,N_5017,N_5661);
nand U12107 (N_12107,N_7786,N_6166);
nor U12108 (N_12108,N_9317,N_6486);
or U12109 (N_12109,N_5945,N_7884);
or U12110 (N_12110,N_6488,N_9147);
nor U12111 (N_12111,N_5270,N_6914);
nor U12112 (N_12112,N_6843,N_8378);
nor U12113 (N_12113,N_5314,N_9039);
nor U12114 (N_12114,N_5863,N_7742);
or U12115 (N_12115,N_5152,N_6849);
nand U12116 (N_12116,N_5457,N_8550);
or U12117 (N_12117,N_8547,N_7823);
nand U12118 (N_12118,N_6343,N_8800);
nor U12119 (N_12119,N_9640,N_5847);
or U12120 (N_12120,N_6038,N_7501);
nand U12121 (N_12121,N_8076,N_9599);
nand U12122 (N_12122,N_8635,N_6053);
or U12123 (N_12123,N_8655,N_6126);
nand U12124 (N_12124,N_9330,N_8813);
xor U12125 (N_12125,N_9779,N_8597);
or U12126 (N_12126,N_8611,N_5824);
xor U12127 (N_12127,N_7275,N_5133);
nand U12128 (N_12128,N_5328,N_7136);
nand U12129 (N_12129,N_8071,N_5814);
nor U12130 (N_12130,N_7196,N_9339);
and U12131 (N_12131,N_9963,N_9593);
nor U12132 (N_12132,N_8691,N_5522);
nor U12133 (N_12133,N_8899,N_5049);
or U12134 (N_12134,N_7103,N_7590);
nand U12135 (N_12135,N_9906,N_6404);
or U12136 (N_12136,N_9010,N_5136);
and U12137 (N_12137,N_8644,N_5562);
nor U12138 (N_12138,N_6692,N_7905);
nand U12139 (N_12139,N_5025,N_9580);
and U12140 (N_12140,N_8391,N_9964);
or U12141 (N_12141,N_7530,N_8440);
nand U12142 (N_12142,N_5650,N_6689);
and U12143 (N_12143,N_6018,N_7282);
and U12144 (N_12144,N_7912,N_5566);
xnor U12145 (N_12145,N_6917,N_9744);
nor U12146 (N_12146,N_8972,N_9909);
nor U12147 (N_12147,N_7046,N_5088);
or U12148 (N_12148,N_6537,N_8648);
xnor U12149 (N_12149,N_8815,N_5318);
nand U12150 (N_12150,N_5697,N_6080);
and U12151 (N_12151,N_6735,N_8119);
and U12152 (N_12152,N_8274,N_5819);
or U12153 (N_12153,N_6069,N_5807);
and U12154 (N_12154,N_9390,N_8004);
xor U12155 (N_12155,N_6579,N_6039);
nand U12156 (N_12156,N_5951,N_7921);
nor U12157 (N_12157,N_5418,N_7060);
xnor U12158 (N_12158,N_7911,N_6032);
nor U12159 (N_12159,N_7588,N_7935);
nand U12160 (N_12160,N_6366,N_7644);
and U12161 (N_12161,N_5447,N_6580);
and U12162 (N_12162,N_5648,N_6682);
nand U12163 (N_12163,N_8660,N_5752);
or U12164 (N_12164,N_8329,N_6021);
xnor U12165 (N_12165,N_8030,N_6666);
and U12166 (N_12166,N_5310,N_8666);
xnor U12167 (N_12167,N_6208,N_7788);
nor U12168 (N_12168,N_7514,N_7737);
or U12169 (N_12169,N_9068,N_9130);
and U12170 (N_12170,N_7333,N_5020);
nand U12171 (N_12171,N_6458,N_5998);
or U12172 (N_12172,N_9821,N_9045);
nor U12173 (N_12173,N_6884,N_6881);
or U12174 (N_12174,N_7184,N_9468);
nand U12175 (N_12175,N_5364,N_8485);
and U12176 (N_12176,N_6956,N_9579);
nor U12177 (N_12177,N_8482,N_7332);
nand U12178 (N_12178,N_9205,N_6304);
nand U12179 (N_12179,N_9485,N_8000);
nand U12180 (N_12180,N_8760,N_9048);
nand U12181 (N_12181,N_7340,N_9266);
and U12182 (N_12182,N_8261,N_7980);
nor U12183 (N_12183,N_7481,N_8885);
and U12184 (N_12184,N_8241,N_5363);
nor U12185 (N_12185,N_9357,N_8372);
and U12186 (N_12186,N_9500,N_9938);
and U12187 (N_12187,N_6940,N_6167);
or U12188 (N_12188,N_6822,N_5887);
nand U12189 (N_12189,N_9533,N_7153);
nor U12190 (N_12190,N_9248,N_6432);
or U12191 (N_12191,N_7584,N_8549);
nand U12192 (N_12192,N_8105,N_6461);
nor U12193 (N_12193,N_7429,N_9140);
nor U12194 (N_12194,N_8228,N_8106);
or U12195 (N_12195,N_9899,N_8796);
nand U12196 (N_12196,N_6160,N_9622);
xor U12197 (N_12197,N_5151,N_5803);
and U12198 (N_12198,N_7717,N_7566);
and U12199 (N_12199,N_8733,N_9279);
or U12200 (N_12200,N_6549,N_7816);
and U12201 (N_12201,N_5866,N_5740);
nand U12202 (N_12202,N_5426,N_8519);
xor U12203 (N_12203,N_6281,N_5836);
or U12204 (N_12204,N_6620,N_7953);
or U12205 (N_12205,N_6324,N_7914);
or U12206 (N_12206,N_7230,N_9786);
or U12207 (N_12207,N_9255,N_5190);
or U12208 (N_12208,N_9925,N_9838);
nand U12209 (N_12209,N_5937,N_6098);
or U12210 (N_12210,N_9814,N_7551);
and U12211 (N_12211,N_8284,N_8040);
and U12212 (N_12212,N_6007,N_6609);
xnor U12213 (N_12213,N_6630,N_8095);
xor U12214 (N_12214,N_6177,N_5780);
nand U12215 (N_12215,N_5094,N_7308);
nand U12216 (N_12216,N_6624,N_6900);
and U12217 (N_12217,N_5009,N_9276);
nand U12218 (N_12218,N_5579,N_7454);
nand U12219 (N_12219,N_5908,N_8538);
nand U12220 (N_12220,N_9258,N_5641);
nor U12221 (N_12221,N_8269,N_5070);
and U12222 (N_12222,N_8463,N_9898);
and U12223 (N_12223,N_6728,N_6791);
or U12224 (N_12224,N_6471,N_8522);
nand U12225 (N_12225,N_7447,N_7358);
nor U12226 (N_12226,N_5727,N_9449);
and U12227 (N_12227,N_9508,N_5730);
and U12228 (N_12228,N_6329,N_8223);
nand U12229 (N_12229,N_6109,N_5783);
and U12230 (N_12230,N_9164,N_7463);
nor U12231 (N_12231,N_9469,N_8890);
or U12232 (N_12232,N_6294,N_8345);
or U12233 (N_12233,N_9990,N_5113);
nand U12234 (N_12234,N_9596,N_8394);
nor U12235 (N_12235,N_9612,N_8715);
and U12236 (N_12236,N_6045,N_7779);
nand U12237 (N_12237,N_6734,N_8860);
nand U12238 (N_12238,N_6544,N_7027);
or U12239 (N_12239,N_8254,N_7265);
nand U12240 (N_12240,N_7050,N_5782);
or U12241 (N_12241,N_7007,N_9768);
nand U12242 (N_12242,N_6535,N_9423);
nor U12243 (N_12243,N_5639,N_6477);
and U12244 (N_12244,N_6173,N_7837);
nor U12245 (N_12245,N_6195,N_8672);
or U12246 (N_12246,N_9626,N_9534);
and U12247 (N_12247,N_8724,N_8323);
nor U12248 (N_12248,N_6674,N_5035);
xor U12249 (N_12249,N_7493,N_5703);
nor U12250 (N_12250,N_5791,N_8128);
nor U12251 (N_12251,N_5157,N_7663);
xnor U12252 (N_12252,N_5323,N_5748);
or U12253 (N_12253,N_5893,N_5312);
xor U12254 (N_12254,N_9058,N_7984);
nor U12255 (N_12255,N_9144,N_9521);
and U12256 (N_12256,N_5356,N_7312);
nand U12257 (N_12257,N_7169,N_6306);
nand U12258 (N_12258,N_6785,N_9832);
nand U12259 (N_12259,N_5739,N_7017);
nand U12260 (N_12260,N_8895,N_7579);
nor U12261 (N_12261,N_6676,N_9067);
or U12262 (N_12262,N_5135,N_7171);
or U12263 (N_12263,N_8508,N_7250);
nor U12264 (N_12264,N_8450,N_8361);
nand U12265 (N_12265,N_5580,N_8238);
and U12266 (N_12266,N_9804,N_7180);
nor U12267 (N_12267,N_7144,N_5143);
nand U12268 (N_12268,N_5950,N_9213);
or U12269 (N_12269,N_8981,N_9675);
nor U12270 (N_12270,N_5523,N_8436);
nand U12271 (N_12271,N_9473,N_9021);
and U12272 (N_12272,N_5698,N_7903);
and U12273 (N_12273,N_9371,N_9143);
nor U12274 (N_12274,N_7746,N_8198);
nor U12275 (N_12275,N_6364,N_6522);
and U12276 (N_12276,N_6631,N_6277);
and U12277 (N_12277,N_7448,N_8253);
nand U12278 (N_12278,N_9607,N_7240);
nor U12279 (N_12279,N_7278,N_9871);
and U12280 (N_12280,N_9588,N_8464);
nor U12281 (N_12281,N_5344,N_9451);
nand U12282 (N_12282,N_7792,N_5346);
nand U12283 (N_12283,N_8523,N_5297);
or U12284 (N_12284,N_7343,N_5255);
nand U12285 (N_12285,N_7801,N_6754);
xor U12286 (N_12286,N_8426,N_6283);
nor U12287 (N_12287,N_6528,N_6156);
or U12288 (N_12288,N_8383,N_7248);
nand U12289 (N_12289,N_5416,N_8507);
nor U12290 (N_12290,N_5464,N_9919);
nor U12291 (N_12291,N_6235,N_9174);
nor U12292 (N_12292,N_9019,N_8540);
nand U12293 (N_12293,N_9206,N_8946);
nor U12294 (N_12294,N_7826,N_8208);
nor U12295 (N_12295,N_6788,N_9849);
nand U12296 (N_12296,N_8741,N_9781);
or U12297 (N_12297,N_7594,N_7672);
or U12298 (N_12298,N_5446,N_7272);
nand U12299 (N_12299,N_7203,N_7256);
or U12300 (N_12300,N_8661,N_7088);
nor U12301 (N_12301,N_7099,N_5917);
xor U12302 (N_12302,N_6931,N_5802);
nor U12303 (N_12303,N_7861,N_9714);
and U12304 (N_12304,N_8116,N_9817);
and U12305 (N_12305,N_7564,N_5554);
or U12306 (N_12306,N_6449,N_7239);
nor U12307 (N_12307,N_6202,N_8102);
nor U12308 (N_12308,N_6102,N_8364);
or U12309 (N_12309,N_7487,N_9306);
and U12310 (N_12310,N_6819,N_6245);
or U12311 (N_12311,N_5853,N_9812);
or U12312 (N_12312,N_7417,N_5677);
nand U12313 (N_12313,N_8565,N_9652);
and U12314 (N_12314,N_7550,N_6746);
nor U12315 (N_12315,N_5095,N_9564);
and U12316 (N_12316,N_5140,N_5002);
nand U12317 (N_12317,N_6699,N_5913);
or U12318 (N_12318,N_6410,N_7299);
and U12319 (N_12319,N_9710,N_9699);
nand U12320 (N_12320,N_5149,N_8993);
or U12321 (N_12321,N_9040,N_8036);
nand U12322 (N_12322,N_6232,N_7371);
nand U12323 (N_12323,N_8674,N_5642);
and U12324 (N_12324,N_5761,N_6194);
nor U12325 (N_12325,N_7133,N_9073);
nand U12326 (N_12326,N_9870,N_9290);
xnor U12327 (N_12327,N_5091,N_6266);
nor U12328 (N_12328,N_5201,N_7190);
and U12329 (N_12329,N_6979,N_6481);
and U12330 (N_12330,N_8614,N_8545);
or U12331 (N_12331,N_5558,N_5857);
nand U12332 (N_12332,N_6573,N_6696);
nand U12333 (N_12333,N_5010,N_9750);
nand U12334 (N_12334,N_6521,N_5546);
nand U12335 (N_12335,N_7199,N_6894);
nand U12336 (N_12336,N_6108,N_8038);
or U12337 (N_12337,N_5517,N_8510);
and U12338 (N_12338,N_9712,N_5529);
nand U12339 (N_12339,N_8216,N_7900);
nor U12340 (N_12340,N_5239,N_8787);
or U12341 (N_12341,N_5161,N_6837);
or U12342 (N_12342,N_9884,N_6806);
or U12343 (N_12343,N_7795,N_8047);
nand U12344 (N_12344,N_6067,N_9690);
or U12345 (N_12345,N_7595,N_9772);
nand U12346 (N_12346,N_6547,N_8709);
and U12347 (N_12347,N_7662,N_9227);
and U12348 (N_12348,N_7314,N_6380);
nor U12349 (N_12349,N_6375,N_8135);
and U12350 (N_12350,N_6805,N_9438);
and U12351 (N_12351,N_7599,N_6107);
xor U12352 (N_12352,N_5325,N_7726);
and U12353 (N_12353,N_8775,N_9074);
and U12354 (N_12354,N_6459,N_9374);
and U12355 (N_12355,N_8471,N_6863);
and U12356 (N_12356,N_7628,N_8761);
nand U12357 (N_12357,N_5362,N_8985);
nor U12358 (N_12358,N_7560,N_5537);
or U12359 (N_12359,N_5815,N_7164);
nor U12360 (N_12360,N_8133,N_6862);
or U12361 (N_12361,N_5139,N_8818);
or U12362 (N_12362,N_9152,N_7149);
and U12363 (N_12363,N_9217,N_6383);
and U12364 (N_12364,N_7691,N_8470);
or U12365 (N_12365,N_6833,N_5121);
and U12366 (N_12366,N_8747,N_7219);
and U12367 (N_12367,N_7437,N_8876);
nor U12368 (N_12368,N_9940,N_7019);
nor U12369 (N_12369,N_5667,N_6767);
nand U12370 (N_12370,N_6106,N_5209);
nor U12371 (N_12371,N_8175,N_8276);
and U12372 (N_12372,N_7005,N_6310);
nand U12373 (N_12373,N_8671,N_7261);
or U12374 (N_12374,N_6966,N_6262);
and U12375 (N_12375,N_7904,N_9598);
nor U12376 (N_12376,N_5626,N_9052);
nand U12377 (N_12377,N_9782,N_7479);
nor U12378 (N_12378,N_5031,N_6346);
xnor U12379 (N_12379,N_7877,N_8446);
nand U12380 (N_12380,N_9448,N_6276);
xor U12381 (N_12381,N_7857,N_5269);
or U12382 (N_12382,N_6622,N_6079);
nor U12383 (N_12383,N_7542,N_7310);
nand U12384 (N_12384,N_7913,N_5460);
nor U12385 (N_12385,N_5692,N_5831);
or U12386 (N_12386,N_8765,N_9214);
and U12387 (N_12387,N_5871,N_9841);
or U12388 (N_12388,N_6002,N_7045);
nand U12389 (N_12389,N_7321,N_5723);
and U12390 (N_12390,N_9133,N_5309);
nor U12391 (N_12391,N_5575,N_8498);
nor U12392 (N_12392,N_5052,N_7907);
nor U12393 (N_12393,N_6723,N_6313);
nor U12394 (N_12394,N_9993,N_6011);
and U12395 (N_12395,N_7832,N_7521);
nor U12396 (N_12396,N_8653,N_6853);
and U12397 (N_12397,N_9329,N_8609);
nand U12398 (N_12398,N_6604,N_9237);
and U12399 (N_12399,N_5860,N_8893);
and U12400 (N_12400,N_6740,N_8186);
nand U12401 (N_12401,N_9912,N_8315);
or U12402 (N_12402,N_5120,N_9264);
and U12403 (N_12403,N_7618,N_5258);
or U12404 (N_12404,N_8569,N_5054);
or U12405 (N_12405,N_9787,N_9332);
or U12406 (N_12406,N_9233,N_9848);
nand U12407 (N_12407,N_8286,N_6035);
nor U12408 (N_12408,N_8606,N_9503);
and U12409 (N_12409,N_7324,N_9682);
xnor U12410 (N_12410,N_9292,N_5072);
nand U12411 (N_12411,N_5666,N_6637);
or U12412 (N_12412,N_5758,N_9440);
nor U12413 (N_12413,N_8409,N_9457);
nor U12414 (N_12414,N_9082,N_7356);
nor U12415 (N_12415,N_9231,N_6057);
or U12416 (N_12416,N_9261,N_6319);
nor U12417 (N_12417,N_7423,N_8603);
and U12418 (N_12418,N_7844,N_6298);
and U12419 (N_12419,N_6958,N_5967);
xnor U12420 (N_12420,N_8712,N_5584);
nor U12421 (N_12421,N_5547,N_8278);
or U12422 (N_12422,N_9971,N_5800);
and U12423 (N_12423,N_6553,N_9136);
xor U12424 (N_12424,N_6415,N_5468);
and U12425 (N_12425,N_5515,N_7875);
nor U12426 (N_12426,N_8828,N_9354);
and U12427 (N_12427,N_7139,N_6872);
nor U12428 (N_12428,N_6897,N_5175);
nand U12429 (N_12429,N_6617,N_7003);
nor U12430 (N_12430,N_9429,N_8749);
nand U12431 (N_12431,N_6576,N_7235);
nor U12432 (N_12432,N_8535,N_7965);
or U12433 (N_12433,N_5180,N_9771);
nand U12434 (N_12434,N_7382,N_6200);
nand U12435 (N_12435,N_5636,N_7059);
nand U12436 (N_12436,N_8330,N_9428);
nor U12437 (N_12437,N_6358,N_5767);
and U12438 (N_12438,N_8407,N_8579);
xor U12439 (N_12439,N_9916,N_7405);
and U12440 (N_12440,N_7768,N_7739);
or U12441 (N_12441,N_9706,N_8750);
xnor U12442 (N_12442,N_8543,N_8931);
and U12443 (N_12443,N_5405,N_6448);
nand U12444 (N_12444,N_9518,N_7697);
and U12445 (N_12445,N_6436,N_9594);
and U12446 (N_12446,N_5775,N_8699);
or U12447 (N_12447,N_6337,N_7020);
and U12448 (N_12448,N_9463,N_6187);
xor U12449 (N_12449,N_9441,N_9194);
nor U12450 (N_12450,N_7369,N_8798);
nor U12451 (N_12451,N_8408,N_5912);
nand U12452 (N_12452,N_9242,N_5237);
nand U12453 (N_12453,N_6640,N_9490);
nor U12454 (N_12454,N_6063,N_7209);
nand U12455 (N_12455,N_7546,N_8397);
or U12456 (N_12456,N_6462,N_5164);
xnor U12457 (N_12457,N_7234,N_9338);
or U12458 (N_12458,N_8657,N_7970);
and U12459 (N_12459,N_9119,N_5084);
or U12460 (N_12460,N_7186,N_7404);
xor U12461 (N_12461,N_7440,N_6984);
nor U12462 (N_12462,N_8246,N_7931);
or U12463 (N_12463,N_5379,N_6447);
or U12464 (N_12464,N_7689,N_7062);
and U12465 (N_12465,N_9818,N_6344);
nand U12466 (N_12466,N_9162,N_6264);
or U12467 (N_12467,N_5770,N_5116);
xor U12468 (N_12468,N_8010,N_7712);
and U12469 (N_12469,N_5852,N_6317);
or U12470 (N_12470,N_8170,N_8511);
nor U12471 (N_12471,N_5742,N_6003);
or U12472 (N_12472,N_5338,N_5154);
and U12473 (N_12473,N_7419,N_6781);
nand U12474 (N_12474,N_6440,N_5862);
nand U12475 (N_12475,N_8790,N_6568);
or U12476 (N_12476,N_8406,N_8452);
or U12477 (N_12477,N_7342,N_5208);
or U12478 (N_12478,N_5039,N_7280);
nor U12479 (N_12479,N_6223,N_6483);
nand U12480 (N_12480,N_8056,N_7370);
and U12481 (N_12481,N_6587,N_6237);
nor U12482 (N_12482,N_8130,N_9088);
nand U12483 (N_12483,N_5583,N_7751);
nor U12484 (N_12484,N_7558,N_7129);
and U12485 (N_12485,N_8366,N_7981);
nand U12486 (N_12486,N_5902,N_7468);
nor U12487 (N_12487,N_8670,N_6951);
or U12488 (N_12488,N_9746,N_6726);
or U12489 (N_12489,N_9113,N_8964);
or U12490 (N_12490,N_7942,N_6105);
and U12491 (N_12491,N_6405,N_9560);
nor U12492 (N_12492,N_8367,N_8483);
and U12493 (N_12493,N_6096,N_5557);
nor U12494 (N_12494,N_6292,N_6077);
nand U12495 (N_12495,N_9683,N_8696);
nor U12496 (N_12496,N_6851,N_5795);
nand U12497 (N_12497,N_7645,N_8599);
nand U12498 (N_12498,N_6725,N_6290);
xnor U12499 (N_12499,N_5746,N_7403);
nand U12500 (N_12500,N_7235,N_5601);
nor U12501 (N_12501,N_8928,N_8403);
and U12502 (N_12502,N_6811,N_6573);
nand U12503 (N_12503,N_9036,N_6577);
or U12504 (N_12504,N_8416,N_8338);
or U12505 (N_12505,N_7907,N_9092);
xor U12506 (N_12506,N_5664,N_5582);
or U12507 (N_12507,N_8785,N_6564);
nand U12508 (N_12508,N_8874,N_6926);
nand U12509 (N_12509,N_7474,N_7912);
nand U12510 (N_12510,N_8356,N_5404);
and U12511 (N_12511,N_9609,N_6474);
nor U12512 (N_12512,N_5055,N_7578);
nand U12513 (N_12513,N_8038,N_7462);
or U12514 (N_12514,N_7669,N_8676);
xor U12515 (N_12515,N_8633,N_9805);
nor U12516 (N_12516,N_8239,N_6666);
xnor U12517 (N_12517,N_9446,N_9422);
nor U12518 (N_12518,N_5459,N_9733);
nand U12519 (N_12519,N_5433,N_5789);
and U12520 (N_12520,N_7436,N_8923);
and U12521 (N_12521,N_5544,N_5325);
nor U12522 (N_12522,N_7998,N_6487);
xnor U12523 (N_12523,N_5117,N_8557);
nand U12524 (N_12524,N_7120,N_8251);
and U12525 (N_12525,N_6451,N_8999);
or U12526 (N_12526,N_9508,N_8874);
nor U12527 (N_12527,N_6940,N_5206);
and U12528 (N_12528,N_5125,N_7184);
xor U12529 (N_12529,N_6536,N_7785);
xor U12530 (N_12530,N_6903,N_9424);
or U12531 (N_12531,N_6594,N_5266);
or U12532 (N_12532,N_9151,N_7418);
or U12533 (N_12533,N_8201,N_8759);
nand U12534 (N_12534,N_9036,N_7724);
nor U12535 (N_12535,N_9005,N_5083);
nand U12536 (N_12536,N_7258,N_5596);
nand U12537 (N_12537,N_5238,N_5647);
and U12538 (N_12538,N_7966,N_5945);
nor U12539 (N_12539,N_8739,N_6107);
and U12540 (N_12540,N_5076,N_5271);
nand U12541 (N_12541,N_8744,N_8108);
nor U12542 (N_12542,N_8807,N_8090);
nor U12543 (N_12543,N_6096,N_9334);
or U12544 (N_12544,N_8487,N_5894);
nand U12545 (N_12545,N_8916,N_8599);
or U12546 (N_12546,N_7635,N_8587);
nor U12547 (N_12547,N_8529,N_8573);
nand U12548 (N_12548,N_5357,N_9268);
and U12549 (N_12549,N_6591,N_7997);
and U12550 (N_12550,N_6064,N_5758);
and U12551 (N_12551,N_5082,N_8639);
or U12552 (N_12552,N_7549,N_9795);
and U12553 (N_12553,N_5012,N_8920);
nor U12554 (N_12554,N_8766,N_9504);
and U12555 (N_12555,N_5090,N_6559);
xnor U12556 (N_12556,N_5125,N_9174);
or U12557 (N_12557,N_6946,N_8060);
or U12558 (N_12558,N_6720,N_5811);
and U12559 (N_12559,N_6807,N_5541);
or U12560 (N_12560,N_5246,N_9397);
nor U12561 (N_12561,N_8968,N_5664);
nand U12562 (N_12562,N_6502,N_7167);
nand U12563 (N_12563,N_6632,N_8849);
or U12564 (N_12564,N_9610,N_9715);
nor U12565 (N_12565,N_7906,N_9345);
nand U12566 (N_12566,N_9915,N_8068);
and U12567 (N_12567,N_7030,N_9220);
nor U12568 (N_12568,N_7489,N_7582);
nand U12569 (N_12569,N_6121,N_6575);
nor U12570 (N_12570,N_8000,N_5701);
or U12571 (N_12571,N_8586,N_7452);
xnor U12572 (N_12572,N_9500,N_8770);
nand U12573 (N_12573,N_7068,N_6896);
nand U12574 (N_12574,N_5609,N_6517);
or U12575 (N_12575,N_6910,N_7324);
and U12576 (N_12576,N_7700,N_5405);
and U12577 (N_12577,N_6062,N_8078);
xor U12578 (N_12578,N_7321,N_5104);
and U12579 (N_12579,N_6219,N_7070);
and U12580 (N_12580,N_6539,N_6558);
and U12581 (N_12581,N_5082,N_7281);
and U12582 (N_12582,N_5604,N_6194);
nor U12583 (N_12583,N_6376,N_5226);
nand U12584 (N_12584,N_6963,N_8981);
and U12585 (N_12585,N_5195,N_6214);
xnor U12586 (N_12586,N_7235,N_5542);
nor U12587 (N_12587,N_6736,N_8239);
xnor U12588 (N_12588,N_5108,N_9400);
and U12589 (N_12589,N_9322,N_7401);
nor U12590 (N_12590,N_8901,N_7114);
nor U12591 (N_12591,N_5802,N_8865);
and U12592 (N_12592,N_9895,N_8259);
and U12593 (N_12593,N_8883,N_6471);
and U12594 (N_12594,N_5182,N_6102);
or U12595 (N_12595,N_5915,N_7814);
and U12596 (N_12596,N_6733,N_9732);
xnor U12597 (N_12597,N_9758,N_5893);
nor U12598 (N_12598,N_5334,N_5757);
nor U12599 (N_12599,N_5374,N_8693);
nor U12600 (N_12600,N_8769,N_8248);
and U12601 (N_12601,N_9837,N_5503);
or U12602 (N_12602,N_8000,N_9187);
nor U12603 (N_12603,N_5840,N_8523);
and U12604 (N_12604,N_7248,N_8727);
nand U12605 (N_12605,N_7606,N_9258);
or U12606 (N_12606,N_6826,N_8270);
and U12607 (N_12607,N_9517,N_8070);
or U12608 (N_12608,N_6956,N_8028);
or U12609 (N_12609,N_6084,N_9696);
and U12610 (N_12610,N_7597,N_6637);
or U12611 (N_12611,N_6690,N_7572);
or U12612 (N_12612,N_8171,N_8296);
or U12613 (N_12613,N_7062,N_9063);
nor U12614 (N_12614,N_9729,N_8905);
nor U12615 (N_12615,N_7007,N_5975);
and U12616 (N_12616,N_5808,N_8937);
nand U12617 (N_12617,N_9445,N_9345);
and U12618 (N_12618,N_5494,N_5026);
or U12619 (N_12619,N_8582,N_6994);
and U12620 (N_12620,N_5458,N_7723);
nand U12621 (N_12621,N_8057,N_8680);
nand U12622 (N_12622,N_8847,N_7582);
and U12623 (N_12623,N_9590,N_8446);
nor U12624 (N_12624,N_5867,N_5341);
and U12625 (N_12625,N_7092,N_5652);
xor U12626 (N_12626,N_6990,N_9735);
nor U12627 (N_12627,N_9724,N_9010);
nor U12628 (N_12628,N_6675,N_5845);
or U12629 (N_12629,N_6296,N_7546);
nor U12630 (N_12630,N_7226,N_6906);
nor U12631 (N_12631,N_8662,N_6317);
xor U12632 (N_12632,N_5757,N_5614);
or U12633 (N_12633,N_9655,N_7281);
nor U12634 (N_12634,N_8661,N_7627);
or U12635 (N_12635,N_7198,N_6134);
nor U12636 (N_12636,N_6753,N_7402);
xnor U12637 (N_12637,N_8026,N_7942);
or U12638 (N_12638,N_9370,N_7803);
xnor U12639 (N_12639,N_9159,N_5851);
nand U12640 (N_12640,N_6532,N_7820);
or U12641 (N_12641,N_7023,N_9592);
or U12642 (N_12642,N_5204,N_5281);
nor U12643 (N_12643,N_7165,N_9489);
and U12644 (N_12644,N_5521,N_8024);
or U12645 (N_12645,N_8815,N_8363);
nor U12646 (N_12646,N_5511,N_7380);
and U12647 (N_12647,N_9979,N_5727);
or U12648 (N_12648,N_9239,N_7893);
and U12649 (N_12649,N_6642,N_9954);
nand U12650 (N_12650,N_5396,N_5744);
and U12651 (N_12651,N_8969,N_6722);
and U12652 (N_12652,N_9022,N_8099);
nor U12653 (N_12653,N_5663,N_9222);
or U12654 (N_12654,N_9576,N_8189);
and U12655 (N_12655,N_5089,N_9468);
and U12656 (N_12656,N_9314,N_6246);
and U12657 (N_12657,N_9003,N_9650);
nand U12658 (N_12658,N_8407,N_6427);
and U12659 (N_12659,N_7098,N_5208);
nand U12660 (N_12660,N_7540,N_5121);
nor U12661 (N_12661,N_5070,N_6042);
and U12662 (N_12662,N_8841,N_5399);
or U12663 (N_12663,N_7850,N_5124);
nand U12664 (N_12664,N_9580,N_8273);
nor U12665 (N_12665,N_6136,N_6189);
nor U12666 (N_12666,N_6696,N_5291);
and U12667 (N_12667,N_6273,N_8879);
nor U12668 (N_12668,N_9982,N_6607);
nor U12669 (N_12669,N_5312,N_8256);
nor U12670 (N_12670,N_6675,N_8768);
nand U12671 (N_12671,N_8555,N_5494);
and U12672 (N_12672,N_8609,N_6150);
nor U12673 (N_12673,N_6943,N_9406);
or U12674 (N_12674,N_5737,N_5998);
and U12675 (N_12675,N_8349,N_6804);
xnor U12676 (N_12676,N_6212,N_6134);
or U12677 (N_12677,N_8354,N_5614);
nand U12678 (N_12678,N_5914,N_6214);
and U12679 (N_12679,N_5173,N_9476);
nand U12680 (N_12680,N_6562,N_7573);
or U12681 (N_12681,N_9906,N_9622);
nor U12682 (N_12682,N_8059,N_5241);
or U12683 (N_12683,N_5043,N_9613);
nor U12684 (N_12684,N_7961,N_5165);
nor U12685 (N_12685,N_6076,N_6547);
nand U12686 (N_12686,N_6840,N_9501);
and U12687 (N_12687,N_9358,N_5938);
or U12688 (N_12688,N_9091,N_5962);
nor U12689 (N_12689,N_5824,N_8454);
and U12690 (N_12690,N_7853,N_7340);
nor U12691 (N_12691,N_6949,N_9346);
and U12692 (N_12692,N_8224,N_7560);
and U12693 (N_12693,N_6886,N_5020);
and U12694 (N_12694,N_7249,N_9069);
and U12695 (N_12695,N_8084,N_9612);
and U12696 (N_12696,N_6821,N_7530);
or U12697 (N_12697,N_8921,N_6519);
nor U12698 (N_12698,N_7386,N_8317);
xor U12699 (N_12699,N_6259,N_9052);
nor U12700 (N_12700,N_6060,N_7120);
and U12701 (N_12701,N_5784,N_7801);
nand U12702 (N_12702,N_6002,N_6252);
or U12703 (N_12703,N_9586,N_5423);
nand U12704 (N_12704,N_7955,N_7245);
nand U12705 (N_12705,N_7735,N_6004);
nor U12706 (N_12706,N_8099,N_9936);
or U12707 (N_12707,N_5687,N_8177);
nand U12708 (N_12708,N_8948,N_7125);
nand U12709 (N_12709,N_9323,N_7398);
xor U12710 (N_12710,N_5532,N_7165);
nor U12711 (N_12711,N_6038,N_5367);
and U12712 (N_12712,N_9603,N_9462);
and U12713 (N_12713,N_6569,N_8583);
and U12714 (N_12714,N_9825,N_8377);
xnor U12715 (N_12715,N_9875,N_8485);
and U12716 (N_12716,N_5142,N_7554);
or U12717 (N_12717,N_7124,N_5090);
and U12718 (N_12718,N_9395,N_8947);
nor U12719 (N_12719,N_8210,N_8997);
nand U12720 (N_12720,N_6674,N_9926);
nand U12721 (N_12721,N_7251,N_5815);
nand U12722 (N_12722,N_6967,N_5402);
xnor U12723 (N_12723,N_5699,N_7708);
xnor U12724 (N_12724,N_6176,N_6515);
nor U12725 (N_12725,N_9886,N_6564);
nor U12726 (N_12726,N_6152,N_5317);
and U12727 (N_12727,N_7273,N_7434);
nor U12728 (N_12728,N_7605,N_6457);
and U12729 (N_12729,N_7787,N_9781);
nand U12730 (N_12730,N_6473,N_6155);
xnor U12731 (N_12731,N_5340,N_8321);
nand U12732 (N_12732,N_5547,N_7040);
and U12733 (N_12733,N_7008,N_9010);
xnor U12734 (N_12734,N_9860,N_6140);
nand U12735 (N_12735,N_8035,N_9920);
xor U12736 (N_12736,N_7561,N_5620);
nand U12737 (N_12737,N_8262,N_6669);
xnor U12738 (N_12738,N_6241,N_5985);
nand U12739 (N_12739,N_8313,N_8356);
nand U12740 (N_12740,N_7558,N_6819);
nand U12741 (N_12741,N_5872,N_5483);
nand U12742 (N_12742,N_8273,N_9912);
nand U12743 (N_12743,N_7954,N_6049);
or U12744 (N_12744,N_6327,N_5167);
nor U12745 (N_12745,N_5857,N_8882);
or U12746 (N_12746,N_5410,N_5725);
and U12747 (N_12747,N_8398,N_7058);
or U12748 (N_12748,N_9751,N_7282);
or U12749 (N_12749,N_9398,N_7283);
or U12750 (N_12750,N_7197,N_6602);
nor U12751 (N_12751,N_5084,N_8857);
or U12752 (N_12752,N_7025,N_7702);
and U12753 (N_12753,N_5319,N_5472);
nand U12754 (N_12754,N_7502,N_8465);
nor U12755 (N_12755,N_5823,N_6997);
nand U12756 (N_12756,N_8633,N_5558);
or U12757 (N_12757,N_6512,N_5628);
and U12758 (N_12758,N_5094,N_5278);
and U12759 (N_12759,N_6429,N_7591);
nand U12760 (N_12760,N_5969,N_8591);
or U12761 (N_12761,N_8283,N_8627);
and U12762 (N_12762,N_5396,N_6357);
and U12763 (N_12763,N_7897,N_9042);
and U12764 (N_12764,N_9302,N_7213);
nand U12765 (N_12765,N_8794,N_5663);
nand U12766 (N_12766,N_9635,N_6354);
nand U12767 (N_12767,N_6497,N_7865);
or U12768 (N_12768,N_8397,N_6461);
or U12769 (N_12769,N_6464,N_7573);
nor U12770 (N_12770,N_7889,N_8862);
nor U12771 (N_12771,N_6494,N_7111);
or U12772 (N_12772,N_9735,N_9493);
nand U12773 (N_12773,N_7128,N_7028);
nor U12774 (N_12774,N_5408,N_5782);
or U12775 (N_12775,N_7396,N_7261);
and U12776 (N_12776,N_5175,N_8187);
xor U12777 (N_12777,N_9564,N_7145);
nor U12778 (N_12778,N_8101,N_9720);
or U12779 (N_12779,N_6992,N_8564);
nor U12780 (N_12780,N_9950,N_8276);
nand U12781 (N_12781,N_8835,N_6992);
xnor U12782 (N_12782,N_7284,N_8316);
nand U12783 (N_12783,N_7514,N_8890);
or U12784 (N_12784,N_9137,N_7870);
xnor U12785 (N_12785,N_7239,N_7390);
nand U12786 (N_12786,N_8824,N_7614);
or U12787 (N_12787,N_8224,N_6189);
nor U12788 (N_12788,N_5054,N_5785);
and U12789 (N_12789,N_9810,N_9116);
or U12790 (N_12790,N_5549,N_8172);
nor U12791 (N_12791,N_8958,N_5708);
nor U12792 (N_12792,N_6384,N_9436);
and U12793 (N_12793,N_5537,N_6823);
nand U12794 (N_12794,N_8176,N_9354);
nor U12795 (N_12795,N_9100,N_6911);
or U12796 (N_12796,N_8968,N_9164);
or U12797 (N_12797,N_9443,N_7811);
or U12798 (N_12798,N_8672,N_7784);
nand U12799 (N_12799,N_5245,N_6771);
nand U12800 (N_12800,N_7134,N_9280);
or U12801 (N_12801,N_6998,N_9768);
or U12802 (N_12802,N_5362,N_8203);
nand U12803 (N_12803,N_7663,N_8177);
or U12804 (N_12804,N_6474,N_6994);
nand U12805 (N_12805,N_5401,N_7798);
and U12806 (N_12806,N_9062,N_5093);
or U12807 (N_12807,N_5972,N_9269);
nand U12808 (N_12808,N_5556,N_7199);
nand U12809 (N_12809,N_7873,N_9515);
xnor U12810 (N_12810,N_7707,N_8413);
or U12811 (N_12811,N_5039,N_9941);
and U12812 (N_12812,N_7803,N_6078);
nor U12813 (N_12813,N_8200,N_5977);
or U12814 (N_12814,N_6261,N_6165);
or U12815 (N_12815,N_8026,N_6763);
and U12816 (N_12816,N_9978,N_7000);
nand U12817 (N_12817,N_7544,N_7840);
nor U12818 (N_12818,N_7995,N_5285);
and U12819 (N_12819,N_5854,N_6390);
nand U12820 (N_12820,N_9583,N_5172);
nand U12821 (N_12821,N_8908,N_6250);
nor U12822 (N_12822,N_5005,N_7148);
or U12823 (N_12823,N_9287,N_9937);
and U12824 (N_12824,N_6556,N_8206);
nor U12825 (N_12825,N_6653,N_9816);
or U12826 (N_12826,N_8309,N_9136);
nor U12827 (N_12827,N_6218,N_7131);
xnor U12828 (N_12828,N_7256,N_6782);
nand U12829 (N_12829,N_9738,N_6540);
and U12830 (N_12830,N_5079,N_6099);
or U12831 (N_12831,N_5391,N_9855);
and U12832 (N_12832,N_5851,N_7959);
nor U12833 (N_12833,N_9018,N_7236);
or U12834 (N_12834,N_8930,N_6749);
and U12835 (N_12835,N_7785,N_8124);
nor U12836 (N_12836,N_5589,N_7517);
nand U12837 (N_12837,N_6922,N_7938);
nand U12838 (N_12838,N_7399,N_9078);
or U12839 (N_12839,N_5079,N_7923);
nand U12840 (N_12840,N_6089,N_8980);
nand U12841 (N_12841,N_8522,N_5988);
or U12842 (N_12842,N_5991,N_8973);
nor U12843 (N_12843,N_6057,N_9068);
and U12844 (N_12844,N_5191,N_9272);
nand U12845 (N_12845,N_7028,N_7039);
nor U12846 (N_12846,N_9613,N_7475);
nor U12847 (N_12847,N_5149,N_6150);
nand U12848 (N_12848,N_6658,N_5778);
nor U12849 (N_12849,N_9113,N_8686);
or U12850 (N_12850,N_7949,N_7100);
or U12851 (N_12851,N_9977,N_8913);
nor U12852 (N_12852,N_7485,N_8489);
and U12853 (N_12853,N_6590,N_9513);
and U12854 (N_12854,N_7368,N_5706);
nor U12855 (N_12855,N_7480,N_8172);
or U12856 (N_12856,N_6324,N_9387);
nor U12857 (N_12857,N_7897,N_7885);
or U12858 (N_12858,N_9758,N_8430);
and U12859 (N_12859,N_6396,N_5127);
or U12860 (N_12860,N_6752,N_7927);
nand U12861 (N_12861,N_8470,N_8207);
and U12862 (N_12862,N_6621,N_7452);
or U12863 (N_12863,N_5596,N_5004);
and U12864 (N_12864,N_6300,N_8700);
nor U12865 (N_12865,N_8504,N_5473);
nand U12866 (N_12866,N_6845,N_9193);
nand U12867 (N_12867,N_8409,N_7484);
nand U12868 (N_12868,N_7417,N_9749);
nor U12869 (N_12869,N_6701,N_6341);
nor U12870 (N_12870,N_5283,N_8635);
nand U12871 (N_12871,N_8922,N_9638);
nand U12872 (N_12872,N_8963,N_5659);
nor U12873 (N_12873,N_8916,N_6781);
nand U12874 (N_12874,N_6313,N_7428);
nand U12875 (N_12875,N_7423,N_6167);
and U12876 (N_12876,N_7637,N_7689);
nand U12877 (N_12877,N_9688,N_5953);
nand U12878 (N_12878,N_5668,N_8354);
or U12879 (N_12879,N_6854,N_7536);
and U12880 (N_12880,N_7398,N_8718);
nor U12881 (N_12881,N_7976,N_8014);
nor U12882 (N_12882,N_7646,N_6292);
nand U12883 (N_12883,N_8541,N_5612);
and U12884 (N_12884,N_7978,N_8324);
or U12885 (N_12885,N_6954,N_9808);
nand U12886 (N_12886,N_7855,N_7838);
and U12887 (N_12887,N_8717,N_5730);
or U12888 (N_12888,N_7264,N_7603);
and U12889 (N_12889,N_5514,N_9285);
nor U12890 (N_12890,N_8720,N_8456);
or U12891 (N_12891,N_7905,N_6143);
and U12892 (N_12892,N_9899,N_5040);
nor U12893 (N_12893,N_7039,N_6668);
nor U12894 (N_12894,N_6554,N_5535);
and U12895 (N_12895,N_9488,N_6844);
nand U12896 (N_12896,N_6329,N_7110);
nand U12897 (N_12897,N_9603,N_8375);
nand U12898 (N_12898,N_7003,N_8981);
and U12899 (N_12899,N_6567,N_8646);
and U12900 (N_12900,N_8283,N_7858);
or U12901 (N_12901,N_8826,N_6845);
or U12902 (N_12902,N_7586,N_5252);
xor U12903 (N_12903,N_7482,N_5755);
nor U12904 (N_12904,N_6615,N_5070);
xor U12905 (N_12905,N_6542,N_9790);
or U12906 (N_12906,N_9358,N_5624);
nor U12907 (N_12907,N_8171,N_9502);
or U12908 (N_12908,N_5847,N_9688);
or U12909 (N_12909,N_8268,N_8877);
xor U12910 (N_12910,N_8082,N_5120);
nor U12911 (N_12911,N_9024,N_7286);
or U12912 (N_12912,N_7408,N_6230);
nand U12913 (N_12913,N_5160,N_8977);
xor U12914 (N_12914,N_9738,N_8508);
and U12915 (N_12915,N_6971,N_8637);
and U12916 (N_12916,N_9535,N_8735);
nor U12917 (N_12917,N_7900,N_8988);
and U12918 (N_12918,N_7403,N_5578);
nor U12919 (N_12919,N_8815,N_9201);
nand U12920 (N_12920,N_9858,N_5454);
nand U12921 (N_12921,N_7773,N_5334);
nand U12922 (N_12922,N_6706,N_5411);
and U12923 (N_12923,N_7146,N_6283);
or U12924 (N_12924,N_7040,N_9050);
and U12925 (N_12925,N_7109,N_7796);
nand U12926 (N_12926,N_8288,N_8598);
and U12927 (N_12927,N_9381,N_8981);
nand U12928 (N_12928,N_6061,N_9313);
nand U12929 (N_12929,N_8970,N_5237);
or U12930 (N_12930,N_6401,N_7333);
nand U12931 (N_12931,N_8641,N_9401);
and U12932 (N_12932,N_7491,N_7770);
or U12933 (N_12933,N_9367,N_9792);
nor U12934 (N_12934,N_8993,N_6991);
or U12935 (N_12935,N_8626,N_7717);
nand U12936 (N_12936,N_7163,N_9438);
and U12937 (N_12937,N_8548,N_8340);
or U12938 (N_12938,N_9541,N_9760);
and U12939 (N_12939,N_8001,N_9424);
nand U12940 (N_12940,N_8214,N_8753);
or U12941 (N_12941,N_6609,N_7558);
nor U12942 (N_12942,N_5035,N_6954);
and U12943 (N_12943,N_9817,N_5545);
nor U12944 (N_12944,N_9026,N_8146);
and U12945 (N_12945,N_5761,N_5161);
nor U12946 (N_12946,N_9935,N_5793);
xnor U12947 (N_12947,N_7587,N_5952);
or U12948 (N_12948,N_6829,N_9354);
or U12949 (N_12949,N_5618,N_7588);
or U12950 (N_12950,N_6143,N_9290);
nand U12951 (N_12951,N_8951,N_7677);
nand U12952 (N_12952,N_8090,N_8607);
nand U12953 (N_12953,N_5061,N_9785);
or U12954 (N_12954,N_5544,N_8818);
xor U12955 (N_12955,N_9574,N_5575);
nor U12956 (N_12956,N_9851,N_7348);
nor U12957 (N_12957,N_6336,N_9475);
and U12958 (N_12958,N_5723,N_8311);
nand U12959 (N_12959,N_6454,N_7591);
and U12960 (N_12960,N_6129,N_6330);
xor U12961 (N_12961,N_5625,N_6571);
nand U12962 (N_12962,N_7261,N_5090);
and U12963 (N_12963,N_8329,N_9644);
nor U12964 (N_12964,N_9400,N_6787);
or U12965 (N_12965,N_9719,N_8572);
xnor U12966 (N_12966,N_7269,N_6434);
or U12967 (N_12967,N_9958,N_9590);
nor U12968 (N_12968,N_9530,N_6305);
nor U12969 (N_12969,N_7950,N_7562);
or U12970 (N_12970,N_5566,N_8656);
and U12971 (N_12971,N_6308,N_5515);
xor U12972 (N_12972,N_5774,N_8204);
or U12973 (N_12973,N_9217,N_9116);
and U12974 (N_12974,N_7934,N_9406);
or U12975 (N_12975,N_6802,N_6494);
nand U12976 (N_12976,N_9700,N_9591);
and U12977 (N_12977,N_6340,N_8086);
or U12978 (N_12978,N_7224,N_7891);
nand U12979 (N_12979,N_5397,N_9751);
nor U12980 (N_12980,N_9939,N_7977);
nand U12981 (N_12981,N_5954,N_8113);
and U12982 (N_12982,N_5238,N_7924);
xnor U12983 (N_12983,N_9692,N_5875);
nor U12984 (N_12984,N_6151,N_7405);
and U12985 (N_12985,N_5649,N_5196);
or U12986 (N_12986,N_9164,N_9303);
and U12987 (N_12987,N_5715,N_5000);
nand U12988 (N_12988,N_6506,N_7972);
nand U12989 (N_12989,N_5901,N_6207);
nand U12990 (N_12990,N_8799,N_7239);
nand U12991 (N_12991,N_6678,N_5528);
nor U12992 (N_12992,N_6320,N_8213);
nor U12993 (N_12993,N_6520,N_8192);
or U12994 (N_12994,N_9781,N_5036);
nand U12995 (N_12995,N_7054,N_5392);
nor U12996 (N_12996,N_6601,N_5706);
or U12997 (N_12997,N_8582,N_6965);
and U12998 (N_12998,N_6903,N_9593);
and U12999 (N_12999,N_8755,N_8220);
nand U13000 (N_13000,N_8440,N_7282);
and U13001 (N_13001,N_5474,N_8481);
nand U13002 (N_13002,N_7402,N_5006);
nor U13003 (N_13003,N_6088,N_5812);
xor U13004 (N_13004,N_6137,N_8949);
or U13005 (N_13005,N_6213,N_8232);
and U13006 (N_13006,N_9645,N_6985);
xor U13007 (N_13007,N_7083,N_5129);
or U13008 (N_13008,N_9757,N_8194);
nor U13009 (N_13009,N_6413,N_7003);
or U13010 (N_13010,N_7445,N_7743);
and U13011 (N_13011,N_7558,N_5352);
or U13012 (N_13012,N_8680,N_7875);
or U13013 (N_13013,N_9157,N_8916);
nand U13014 (N_13014,N_6849,N_7471);
and U13015 (N_13015,N_8962,N_7159);
or U13016 (N_13016,N_8132,N_7975);
nand U13017 (N_13017,N_5714,N_8583);
or U13018 (N_13018,N_8957,N_6853);
nor U13019 (N_13019,N_5623,N_6141);
nor U13020 (N_13020,N_5867,N_7823);
xnor U13021 (N_13021,N_8921,N_8515);
or U13022 (N_13022,N_9815,N_9611);
xnor U13023 (N_13023,N_9480,N_9061);
nand U13024 (N_13024,N_7469,N_7676);
nand U13025 (N_13025,N_8657,N_8826);
nor U13026 (N_13026,N_5446,N_9437);
nand U13027 (N_13027,N_9975,N_9142);
and U13028 (N_13028,N_5367,N_5783);
nor U13029 (N_13029,N_9129,N_7233);
and U13030 (N_13030,N_8890,N_6995);
nor U13031 (N_13031,N_6552,N_5117);
nor U13032 (N_13032,N_8128,N_8874);
or U13033 (N_13033,N_7774,N_7742);
xnor U13034 (N_13034,N_6764,N_8007);
or U13035 (N_13035,N_9651,N_5395);
nor U13036 (N_13036,N_9597,N_9945);
or U13037 (N_13037,N_8214,N_6416);
nand U13038 (N_13038,N_9518,N_5271);
nand U13039 (N_13039,N_6012,N_5916);
or U13040 (N_13040,N_8772,N_9125);
nor U13041 (N_13041,N_7916,N_7694);
or U13042 (N_13042,N_6093,N_6167);
nor U13043 (N_13043,N_5041,N_9096);
or U13044 (N_13044,N_8967,N_9579);
or U13045 (N_13045,N_5042,N_9184);
nand U13046 (N_13046,N_8768,N_8916);
nor U13047 (N_13047,N_9938,N_5398);
and U13048 (N_13048,N_6555,N_5146);
and U13049 (N_13049,N_9750,N_6980);
and U13050 (N_13050,N_7953,N_9736);
nor U13051 (N_13051,N_6410,N_8017);
and U13052 (N_13052,N_9903,N_9242);
or U13053 (N_13053,N_5287,N_6324);
nand U13054 (N_13054,N_9610,N_8056);
and U13055 (N_13055,N_5743,N_8170);
and U13056 (N_13056,N_8750,N_7889);
xor U13057 (N_13057,N_9237,N_7628);
nand U13058 (N_13058,N_7148,N_9037);
and U13059 (N_13059,N_5695,N_6436);
nor U13060 (N_13060,N_9171,N_7336);
nand U13061 (N_13061,N_9363,N_9928);
nor U13062 (N_13062,N_5952,N_5473);
and U13063 (N_13063,N_9839,N_5547);
and U13064 (N_13064,N_7896,N_7707);
and U13065 (N_13065,N_7205,N_9931);
nor U13066 (N_13066,N_7276,N_5736);
nand U13067 (N_13067,N_7653,N_8544);
or U13068 (N_13068,N_8942,N_9684);
nor U13069 (N_13069,N_6041,N_9555);
or U13070 (N_13070,N_7492,N_6169);
nor U13071 (N_13071,N_9387,N_7728);
and U13072 (N_13072,N_7537,N_8291);
nor U13073 (N_13073,N_6261,N_6739);
or U13074 (N_13074,N_5829,N_5944);
or U13075 (N_13075,N_8549,N_9013);
nor U13076 (N_13076,N_6159,N_6931);
or U13077 (N_13077,N_9773,N_5625);
nor U13078 (N_13078,N_8079,N_8213);
nor U13079 (N_13079,N_8407,N_7583);
or U13080 (N_13080,N_9623,N_5010);
and U13081 (N_13081,N_5082,N_7735);
nand U13082 (N_13082,N_9580,N_6184);
and U13083 (N_13083,N_7973,N_9314);
nor U13084 (N_13084,N_5298,N_5105);
nand U13085 (N_13085,N_5592,N_8722);
nand U13086 (N_13086,N_5088,N_9447);
or U13087 (N_13087,N_8158,N_7459);
nand U13088 (N_13088,N_8639,N_7758);
nor U13089 (N_13089,N_6711,N_9582);
and U13090 (N_13090,N_9449,N_9944);
or U13091 (N_13091,N_7557,N_5988);
or U13092 (N_13092,N_5636,N_9516);
nand U13093 (N_13093,N_8921,N_6888);
xor U13094 (N_13094,N_5718,N_5967);
nor U13095 (N_13095,N_7932,N_7883);
nor U13096 (N_13096,N_9713,N_5480);
or U13097 (N_13097,N_7379,N_6900);
and U13098 (N_13098,N_5079,N_9048);
or U13099 (N_13099,N_9188,N_6029);
and U13100 (N_13100,N_6226,N_6831);
nand U13101 (N_13101,N_6471,N_6715);
xnor U13102 (N_13102,N_7658,N_9420);
or U13103 (N_13103,N_6616,N_9940);
xor U13104 (N_13104,N_5399,N_5252);
nand U13105 (N_13105,N_6738,N_5464);
and U13106 (N_13106,N_6622,N_8892);
and U13107 (N_13107,N_5592,N_9743);
nor U13108 (N_13108,N_7092,N_6902);
xor U13109 (N_13109,N_7320,N_8247);
xor U13110 (N_13110,N_5139,N_7179);
and U13111 (N_13111,N_5788,N_9860);
nor U13112 (N_13112,N_5101,N_9543);
nand U13113 (N_13113,N_7319,N_8218);
xnor U13114 (N_13114,N_9686,N_7381);
or U13115 (N_13115,N_5434,N_7498);
nor U13116 (N_13116,N_5888,N_9978);
nand U13117 (N_13117,N_9310,N_7678);
and U13118 (N_13118,N_7741,N_6380);
nand U13119 (N_13119,N_6818,N_7687);
nand U13120 (N_13120,N_9893,N_7535);
or U13121 (N_13121,N_6507,N_5765);
or U13122 (N_13122,N_7058,N_7654);
or U13123 (N_13123,N_7095,N_8065);
xnor U13124 (N_13124,N_7159,N_9644);
xor U13125 (N_13125,N_9462,N_8048);
or U13126 (N_13126,N_9097,N_5807);
nor U13127 (N_13127,N_9275,N_6764);
nand U13128 (N_13128,N_9542,N_7007);
or U13129 (N_13129,N_9219,N_7912);
or U13130 (N_13130,N_8639,N_5947);
or U13131 (N_13131,N_6220,N_5842);
nor U13132 (N_13132,N_6681,N_6939);
nor U13133 (N_13133,N_9060,N_9393);
xor U13134 (N_13134,N_8827,N_8350);
nor U13135 (N_13135,N_8622,N_8687);
nand U13136 (N_13136,N_9741,N_8742);
nand U13137 (N_13137,N_8520,N_7738);
and U13138 (N_13138,N_8207,N_5719);
nor U13139 (N_13139,N_6731,N_7704);
and U13140 (N_13140,N_6590,N_5394);
nor U13141 (N_13141,N_6482,N_8348);
nor U13142 (N_13142,N_9730,N_6383);
or U13143 (N_13143,N_6488,N_6221);
nor U13144 (N_13144,N_6264,N_7777);
nor U13145 (N_13145,N_7996,N_7574);
and U13146 (N_13146,N_5069,N_8920);
xnor U13147 (N_13147,N_5004,N_9357);
xor U13148 (N_13148,N_9999,N_6781);
or U13149 (N_13149,N_8431,N_5420);
nor U13150 (N_13150,N_7350,N_6872);
and U13151 (N_13151,N_6409,N_8090);
nor U13152 (N_13152,N_8287,N_5042);
xor U13153 (N_13153,N_7371,N_6202);
nand U13154 (N_13154,N_5520,N_9145);
nor U13155 (N_13155,N_8402,N_7013);
and U13156 (N_13156,N_6150,N_9438);
nand U13157 (N_13157,N_6657,N_5053);
and U13158 (N_13158,N_7090,N_5505);
nand U13159 (N_13159,N_5944,N_7929);
xnor U13160 (N_13160,N_6152,N_6611);
and U13161 (N_13161,N_8035,N_5540);
xor U13162 (N_13162,N_6530,N_6973);
and U13163 (N_13163,N_8240,N_7432);
or U13164 (N_13164,N_7285,N_8700);
nand U13165 (N_13165,N_8235,N_7817);
nor U13166 (N_13166,N_9471,N_7850);
and U13167 (N_13167,N_6734,N_6571);
or U13168 (N_13168,N_7998,N_7308);
or U13169 (N_13169,N_6805,N_5906);
or U13170 (N_13170,N_8152,N_6463);
xnor U13171 (N_13171,N_7730,N_5701);
and U13172 (N_13172,N_8213,N_8444);
or U13173 (N_13173,N_7052,N_5261);
nand U13174 (N_13174,N_6529,N_5823);
and U13175 (N_13175,N_8274,N_6869);
nor U13176 (N_13176,N_5631,N_5753);
nor U13177 (N_13177,N_7885,N_8347);
xor U13178 (N_13178,N_7460,N_5918);
xor U13179 (N_13179,N_6507,N_8099);
nor U13180 (N_13180,N_5713,N_6280);
nand U13181 (N_13181,N_8839,N_8659);
or U13182 (N_13182,N_5077,N_8342);
nand U13183 (N_13183,N_8619,N_6247);
and U13184 (N_13184,N_7285,N_9665);
or U13185 (N_13185,N_7539,N_7088);
and U13186 (N_13186,N_9277,N_8639);
nand U13187 (N_13187,N_8430,N_5051);
or U13188 (N_13188,N_9047,N_6415);
and U13189 (N_13189,N_8569,N_9378);
and U13190 (N_13190,N_7134,N_7807);
xor U13191 (N_13191,N_8375,N_6832);
nand U13192 (N_13192,N_7049,N_6791);
nor U13193 (N_13193,N_8678,N_9241);
and U13194 (N_13194,N_9507,N_5531);
or U13195 (N_13195,N_6119,N_8362);
or U13196 (N_13196,N_6480,N_8158);
nor U13197 (N_13197,N_8784,N_8227);
nor U13198 (N_13198,N_6042,N_5990);
or U13199 (N_13199,N_6528,N_7570);
or U13200 (N_13200,N_8144,N_9478);
or U13201 (N_13201,N_5307,N_7108);
nand U13202 (N_13202,N_9093,N_6626);
nand U13203 (N_13203,N_7289,N_8939);
nand U13204 (N_13204,N_8115,N_7957);
nor U13205 (N_13205,N_6972,N_8394);
or U13206 (N_13206,N_5133,N_7778);
nor U13207 (N_13207,N_9542,N_7418);
or U13208 (N_13208,N_7148,N_9477);
and U13209 (N_13209,N_6822,N_7913);
nor U13210 (N_13210,N_9846,N_5910);
nor U13211 (N_13211,N_9620,N_5354);
nand U13212 (N_13212,N_6521,N_8706);
nand U13213 (N_13213,N_8893,N_5121);
nor U13214 (N_13214,N_9648,N_7504);
and U13215 (N_13215,N_8407,N_9143);
and U13216 (N_13216,N_6603,N_5020);
or U13217 (N_13217,N_6676,N_6368);
nand U13218 (N_13218,N_8069,N_5826);
and U13219 (N_13219,N_8226,N_7611);
xnor U13220 (N_13220,N_9154,N_8898);
and U13221 (N_13221,N_9994,N_5087);
nor U13222 (N_13222,N_6452,N_9844);
xor U13223 (N_13223,N_5775,N_8547);
nand U13224 (N_13224,N_5581,N_6250);
nand U13225 (N_13225,N_5396,N_8939);
xnor U13226 (N_13226,N_5628,N_7720);
nand U13227 (N_13227,N_9966,N_9607);
xnor U13228 (N_13228,N_5191,N_7660);
nor U13229 (N_13229,N_6401,N_7958);
nand U13230 (N_13230,N_5855,N_7812);
and U13231 (N_13231,N_9935,N_9842);
nor U13232 (N_13232,N_9892,N_6897);
and U13233 (N_13233,N_5334,N_9675);
or U13234 (N_13234,N_7989,N_9925);
and U13235 (N_13235,N_6937,N_8235);
nor U13236 (N_13236,N_6563,N_5959);
and U13237 (N_13237,N_5908,N_8998);
nand U13238 (N_13238,N_8077,N_5277);
and U13239 (N_13239,N_6809,N_9193);
nor U13240 (N_13240,N_5785,N_9735);
nor U13241 (N_13241,N_5797,N_5280);
nor U13242 (N_13242,N_5336,N_6956);
or U13243 (N_13243,N_6125,N_6674);
and U13244 (N_13244,N_8705,N_7907);
nand U13245 (N_13245,N_5339,N_5414);
or U13246 (N_13246,N_6769,N_9473);
nor U13247 (N_13247,N_8194,N_8523);
nor U13248 (N_13248,N_7217,N_6642);
xnor U13249 (N_13249,N_6556,N_8531);
or U13250 (N_13250,N_6513,N_5118);
and U13251 (N_13251,N_7870,N_6103);
nand U13252 (N_13252,N_8284,N_8357);
xnor U13253 (N_13253,N_6425,N_6349);
nand U13254 (N_13254,N_5376,N_6451);
and U13255 (N_13255,N_5194,N_5353);
or U13256 (N_13256,N_5272,N_8416);
or U13257 (N_13257,N_8838,N_9103);
or U13258 (N_13258,N_6333,N_5939);
or U13259 (N_13259,N_8593,N_6808);
or U13260 (N_13260,N_7278,N_8917);
nand U13261 (N_13261,N_7884,N_7512);
or U13262 (N_13262,N_9089,N_9741);
nand U13263 (N_13263,N_7789,N_6328);
nand U13264 (N_13264,N_6723,N_6618);
or U13265 (N_13265,N_6504,N_9653);
or U13266 (N_13266,N_5605,N_8129);
nor U13267 (N_13267,N_9636,N_5290);
or U13268 (N_13268,N_6794,N_6283);
nand U13269 (N_13269,N_9958,N_9079);
nor U13270 (N_13270,N_9448,N_7445);
xnor U13271 (N_13271,N_5368,N_9207);
nor U13272 (N_13272,N_8391,N_5632);
xor U13273 (N_13273,N_8301,N_7974);
nor U13274 (N_13274,N_6043,N_6793);
or U13275 (N_13275,N_9030,N_7920);
and U13276 (N_13276,N_7639,N_5023);
xor U13277 (N_13277,N_9632,N_6753);
or U13278 (N_13278,N_7813,N_9532);
nor U13279 (N_13279,N_6058,N_8471);
and U13280 (N_13280,N_5193,N_9095);
nand U13281 (N_13281,N_8527,N_6581);
and U13282 (N_13282,N_6281,N_7316);
and U13283 (N_13283,N_6465,N_6639);
nand U13284 (N_13284,N_7971,N_9051);
xnor U13285 (N_13285,N_5234,N_9896);
nand U13286 (N_13286,N_9643,N_6274);
nor U13287 (N_13287,N_7046,N_9506);
nor U13288 (N_13288,N_9785,N_8750);
and U13289 (N_13289,N_5427,N_5897);
and U13290 (N_13290,N_7097,N_8771);
nand U13291 (N_13291,N_5304,N_5363);
nor U13292 (N_13292,N_5682,N_8707);
and U13293 (N_13293,N_5749,N_8245);
nor U13294 (N_13294,N_9383,N_9185);
nor U13295 (N_13295,N_7705,N_5395);
xnor U13296 (N_13296,N_5096,N_9230);
nor U13297 (N_13297,N_5095,N_9950);
or U13298 (N_13298,N_7083,N_6588);
and U13299 (N_13299,N_8440,N_9412);
nand U13300 (N_13300,N_9499,N_9891);
and U13301 (N_13301,N_8275,N_9019);
nor U13302 (N_13302,N_6523,N_9314);
or U13303 (N_13303,N_7920,N_6009);
and U13304 (N_13304,N_5185,N_5950);
and U13305 (N_13305,N_8284,N_7551);
nand U13306 (N_13306,N_9989,N_8458);
nand U13307 (N_13307,N_9192,N_9485);
nand U13308 (N_13308,N_5150,N_5019);
nand U13309 (N_13309,N_7096,N_8532);
nand U13310 (N_13310,N_8892,N_9773);
nand U13311 (N_13311,N_9553,N_5048);
nand U13312 (N_13312,N_8438,N_5911);
and U13313 (N_13313,N_7620,N_8544);
and U13314 (N_13314,N_7242,N_9596);
xor U13315 (N_13315,N_5555,N_9741);
nor U13316 (N_13316,N_9057,N_6552);
or U13317 (N_13317,N_7513,N_9729);
nor U13318 (N_13318,N_5947,N_5938);
and U13319 (N_13319,N_6901,N_6554);
and U13320 (N_13320,N_8413,N_5231);
and U13321 (N_13321,N_7131,N_6395);
xnor U13322 (N_13322,N_8899,N_5345);
nand U13323 (N_13323,N_9204,N_6722);
nor U13324 (N_13324,N_9202,N_5099);
or U13325 (N_13325,N_5737,N_5600);
nor U13326 (N_13326,N_8410,N_9289);
and U13327 (N_13327,N_6102,N_5938);
xnor U13328 (N_13328,N_8350,N_8015);
nor U13329 (N_13329,N_6906,N_6819);
nor U13330 (N_13330,N_9911,N_8653);
or U13331 (N_13331,N_5558,N_8757);
or U13332 (N_13332,N_6458,N_6283);
or U13333 (N_13333,N_5595,N_7942);
xor U13334 (N_13334,N_7989,N_7275);
and U13335 (N_13335,N_6799,N_6678);
nand U13336 (N_13336,N_7581,N_8644);
or U13337 (N_13337,N_6650,N_9319);
or U13338 (N_13338,N_8631,N_9568);
nor U13339 (N_13339,N_7605,N_9463);
nor U13340 (N_13340,N_5878,N_9619);
nand U13341 (N_13341,N_5803,N_9130);
nor U13342 (N_13342,N_5581,N_5136);
xor U13343 (N_13343,N_9944,N_7959);
nand U13344 (N_13344,N_9063,N_8163);
xor U13345 (N_13345,N_7141,N_5854);
and U13346 (N_13346,N_6451,N_8514);
or U13347 (N_13347,N_8803,N_9355);
nand U13348 (N_13348,N_8180,N_5797);
or U13349 (N_13349,N_8297,N_8432);
nand U13350 (N_13350,N_7726,N_6453);
nor U13351 (N_13351,N_5232,N_5890);
xor U13352 (N_13352,N_9246,N_6908);
nor U13353 (N_13353,N_8360,N_9897);
and U13354 (N_13354,N_6247,N_7389);
xor U13355 (N_13355,N_8002,N_8907);
or U13356 (N_13356,N_6596,N_7797);
nand U13357 (N_13357,N_7740,N_6616);
and U13358 (N_13358,N_9110,N_9551);
or U13359 (N_13359,N_5074,N_9187);
and U13360 (N_13360,N_8656,N_7622);
or U13361 (N_13361,N_9855,N_7654);
nand U13362 (N_13362,N_6759,N_5206);
nor U13363 (N_13363,N_8663,N_5125);
xor U13364 (N_13364,N_7423,N_9376);
nor U13365 (N_13365,N_7345,N_9412);
and U13366 (N_13366,N_8989,N_8824);
nand U13367 (N_13367,N_6786,N_8575);
nand U13368 (N_13368,N_7222,N_8762);
nor U13369 (N_13369,N_9782,N_5471);
nor U13370 (N_13370,N_6032,N_5067);
or U13371 (N_13371,N_9137,N_9505);
nand U13372 (N_13372,N_6142,N_6797);
nor U13373 (N_13373,N_8330,N_6504);
nor U13374 (N_13374,N_6145,N_8565);
nor U13375 (N_13375,N_6384,N_6547);
and U13376 (N_13376,N_8179,N_9811);
or U13377 (N_13377,N_9292,N_6615);
xor U13378 (N_13378,N_9274,N_9278);
xor U13379 (N_13379,N_5694,N_9077);
nor U13380 (N_13380,N_8104,N_9891);
or U13381 (N_13381,N_5426,N_8624);
or U13382 (N_13382,N_8341,N_7899);
nand U13383 (N_13383,N_5573,N_7123);
and U13384 (N_13384,N_9874,N_6831);
nand U13385 (N_13385,N_8440,N_7660);
nand U13386 (N_13386,N_8289,N_5718);
and U13387 (N_13387,N_9125,N_8800);
nor U13388 (N_13388,N_6678,N_9324);
nand U13389 (N_13389,N_9270,N_8661);
and U13390 (N_13390,N_9489,N_6119);
and U13391 (N_13391,N_9782,N_5438);
and U13392 (N_13392,N_5825,N_9646);
nor U13393 (N_13393,N_9312,N_9882);
or U13394 (N_13394,N_7888,N_9391);
or U13395 (N_13395,N_9626,N_8461);
and U13396 (N_13396,N_7902,N_7082);
xor U13397 (N_13397,N_5250,N_9966);
or U13398 (N_13398,N_6348,N_6163);
nor U13399 (N_13399,N_6788,N_6586);
or U13400 (N_13400,N_6304,N_7708);
xnor U13401 (N_13401,N_9486,N_6230);
nor U13402 (N_13402,N_5369,N_6535);
nand U13403 (N_13403,N_8840,N_7961);
or U13404 (N_13404,N_5427,N_6496);
or U13405 (N_13405,N_9650,N_8705);
and U13406 (N_13406,N_8222,N_8068);
and U13407 (N_13407,N_5519,N_5698);
or U13408 (N_13408,N_6621,N_6541);
nand U13409 (N_13409,N_6400,N_8891);
nand U13410 (N_13410,N_7593,N_7327);
and U13411 (N_13411,N_9464,N_9941);
nor U13412 (N_13412,N_8815,N_7912);
and U13413 (N_13413,N_8093,N_9279);
nor U13414 (N_13414,N_6833,N_7887);
nand U13415 (N_13415,N_9133,N_5990);
or U13416 (N_13416,N_5516,N_7487);
and U13417 (N_13417,N_6533,N_5990);
nor U13418 (N_13418,N_9162,N_5213);
nor U13419 (N_13419,N_8387,N_9078);
nand U13420 (N_13420,N_5955,N_7066);
nand U13421 (N_13421,N_8211,N_9548);
and U13422 (N_13422,N_7749,N_7161);
xor U13423 (N_13423,N_5740,N_5399);
or U13424 (N_13424,N_7793,N_5174);
or U13425 (N_13425,N_8120,N_9116);
nor U13426 (N_13426,N_6483,N_9852);
nor U13427 (N_13427,N_6030,N_7728);
or U13428 (N_13428,N_9830,N_6489);
nand U13429 (N_13429,N_9790,N_9876);
nand U13430 (N_13430,N_5632,N_7852);
nand U13431 (N_13431,N_5098,N_7899);
nor U13432 (N_13432,N_9112,N_6647);
or U13433 (N_13433,N_7578,N_5691);
nand U13434 (N_13434,N_8731,N_9605);
or U13435 (N_13435,N_5461,N_5404);
nand U13436 (N_13436,N_8772,N_8153);
nand U13437 (N_13437,N_9081,N_5072);
and U13438 (N_13438,N_8486,N_9259);
xor U13439 (N_13439,N_7867,N_8175);
nor U13440 (N_13440,N_9687,N_6498);
or U13441 (N_13441,N_6844,N_8457);
and U13442 (N_13442,N_5846,N_5209);
nor U13443 (N_13443,N_6365,N_9671);
nand U13444 (N_13444,N_9380,N_9982);
nand U13445 (N_13445,N_5438,N_5733);
and U13446 (N_13446,N_8254,N_8547);
nand U13447 (N_13447,N_9947,N_6215);
or U13448 (N_13448,N_6674,N_7937);
nand U13449 (N_13449,N_8736,N_8811);
nand U13450 (N_13450,N_8638,N_5606);
xnor U13451 (N_13451,N_6843,N_6393);
nand U13452 (N_13452,N_7977,N_6720);
nor U13453 (N_13453,N_7043,N_5564);
nand U13454 (N_13454,N_7548,N_7603);
nor U13455 (N_13455,N_7533,N_9941);
nand U13456 (N_13456,N_9496,N_5823);
or U13457 (N_13457,N_8811,N_6988);
nand U13458 (N_13458,N_8956,N_6152);
and U13459 (N_13459,N_8114,N_6372);
xor U13460 (N_13460,N_8476,N_8976);
nand U13461 (N_13461,N_5199,N_6782);
nor U13462 (N_13462,N_8644,N_9269);
nor U13463 (N_13463,N_6199,N_6483);
and U13464 (N_13464,N_6350,N_9771);
nor U13465 (N_13465,N_7028,N_9893);
nand U13466 (N_13466,N_7265,N_7620);
and U13467 (N_13467,N_6709,N_7683);
and U13468 (N_13468,N_9819,N_5705);
or U13469 (N_13469,N_6191,N_7859);
and U13470 (N_13470,N_7584,N_6547);
and U13471 (N_13471,N_8107,N_8284);
or U13472 (N_13472,N_9853,N_8962);
and U13473 (N_13473,N_8311,N_8837);
nand U13474 (N_13474,N_7518,N_8015);
or U13475 (N_13475,N_6916,N_9924);
nand U13476 (N_13476,N_8137,N_5939);
nand U13477 (N_13477,N_8078,N_8623);
or U13478 (N_13478,N_5434,N_5560);
nor U13479 (N_13479,N_9933,N_7841);
xnor U13480 (N_13480,N_7985,N_9674);
or U13481 (N_13481,N_5644,N_6943);
and U13482 (N_13482,N_7474,N_6738);
or U13483 (N_13483,N_8462,N_9296);
or U13484 (N_13484,N_9242,N_8420);
xnor U13485 (N_13485,N_5245,N_9687);
nor U13486 (N_13486,N_8552,N_7825);
xor U13487 (N_13487,N_7218,N_6355);
and U13488 (N_13488,N_6336,N_6186);
nand U13489 (N_13489,N_6147,N_5334);
and U13490 (N_13490,N_7772,N_8544);
or U13491 (N_13491,N_6177,N_5835);
xnor U13492 (N_13492,N_5886,N_7525);
nand U13493 (N_13493,N_9919,N_6098);
nand U13494 (N_13494,N_7333,N_9214);
nor U13495 (N_13495,N_6009,N_7471);
or U13496 (N_13496,N_9357,N_5898);
and U13497 (N_13497,N_5244,N_6581);
and U13498 (N_13498,N_5230,N_8566);
or U13499 (N_13499,N_8852,N_5085);
nand U13500 (N_13500,N_9987,N_5364);
nand U13501 (N_13501,N_6774,N_6175);
and U13502 (N_13502,N_5161,N_5809);
and U13503 (N_13503,N_6237,N_9434);
nand U13504 (N_13504,N_9550,N_8570);
xnor U13505 (N_13505,N_8006,N_5981);
and U13506 (N_13506,N_9951,N_9860);
nor U13507 (N_13507,N_9941,N_5934);
nand U13508 (N_13508,N_7928,N_6992);
nor U13509 (N_13509,N_9429,N_6877);
or U13510 (N_13510,N_7342,N_5442);
xnor U13511 (N_13511,N_8488,N_7580);
and U13512 (N_13512,N_8150,N_6270);
xnor U13513 (N_13513,N_8063,N_7236);
nand U13514 (N_13514,N_8282,N_8084);
nor U13515 (N_13515,N_8527,N_8468);
nor U13516 (N_13516,N_8809,N_9127);
or U13517 (N_13517,N_9454,N_5594);
nand U13518 (N_13518,N_8846,N_9947);
nand U13519 (N_13519,N_8339,N_5958);
nand U13520 (N_13520,N_9430,N_9308);
nand U13521 (N_13521,N_7506,N_9888);
and U13522 (N_13522,N_9580,N_9559);
nor U13523 (N_13523,N_8378,N_7792);
nand U13524 (N_13524,N_9711,N_6356);
nor U13525 (N_13525,N_8091,N_7242);
xnor U13526 (N_13526,N_8090,N_9511);
nand U13527 (N_13527,N_8521,N_7549);
nand U13528 (N_13528,N_6283,N_6929);
or U13529 (N_13529,N_5121,N_5522);
or U13530 (N_13530,N_5454,N_5068);
and U13531 (N_13531,N_9016,N_9992);
or U13532 (N_13532,N_5123,N_7933);
or U13533 (N_13533,N_5023,N_7959);
nor U13534 (N_13534,N_9773,N_8475);
or U13535 (N_13535,N_9667,N_6904);
or U13536 (N_13536,N_8987,N_7673);
nand U13537 (N_13537,N_9062,N_5764);
nand U13538 (N_13538,N_7230,N_6263);
and U13539 (N_13539,N_7598,N_7377);
or U13540 (N_13540,N_5806,N_6572);
nand U13541 (N_13541,N_8660,N_9592);
xnor U13542 (N_13542,N_5211,N_9306);
nor U13543 (N_13543,N_5951,N_9973);
nor U13544 (N_13544,N_5500,N_9821);
nand U13545 (N_13545,N_5398,N_9229);
or U13546 (N_13546,N_9309,N_8176);
nor U13547 (N_13547,N_8030,N_7275);
nand U13548 (N_13548,N_5124,N_6642);
xnor U13549 (N_13549,N_7688,N_9240);
and U13550 (N_13550,N_5367,N_9585);
xnor U13551 (N_13551,N_8367,N_9856);
or U13552 (N_13552,N_8534,N_8159);
or U13553 (N_13553,N_9721,N_6370);
or U13554 (N_13554,N_9230,N_8316);
nor U13555 (N_13555,N_7813,N_5291);
nand U13556 (N_13556,N_8277,N_6907);
or U13557 (N_13557,N_5180,N_5932);
and U13558 (N_13558,N_5104,N_7903);
nor U13559 (N_13559,N_9033,N_5810);
or U13560 (N_13560,N_7271,N_7354);
nand U13561 (N_13561,N_6107,N_8211);
xor U13562 (N_13562,N_7768,N_6359);
or U13563 (N_13563,N_6283,N_5058);
or U13564 (N_13564,N_8683,N_5547);
and U13565 (N_13565,N_7440,N_5286);
or U13566 (N_13566,N_7040,N_8133);
and U13567 (N_13567,N_8006,N_9998);
and U13568 (N_13568,N_8074,N_5521);
and U13569 (N_13569,N_6504,N_9912);
or U13570 (N_13570,N_5551,N_6342);
or U13571 (N_13571,N_6372,N_5263);
xnor U13572 (N_13572,N_6113,N_9412);
nor U13573 (N_13573,N_7291,N_7046);
xor U13574 (N_13574,N_6737,N_6357);
nand U13575 (N_13575,N_8680,N_7806);
or U13576 (N_13576,N_8019,N_5683);
and U13577 (N_13577,N_9785,N_6630);
nand U13578 (N_13578,N_8738,N_7830);
and U13579 (N_13579,N_9436,N_7178);
nand U13580 (N_13580,N_7389,N_5948);
nand U13581 (N_13581,N_7001,N_8174);
and U13582 (N_13582,N_6131,N_5291);
and U13583 (N_13583,N_8024,N_8243);
nor U13584 (N_13584,N_6300,N_8771);
nor U13585 (N_13585,N_7372,N_7380);
nor U13586 (N_13586,N_5518,N_7270);
nand U13587 (N_13587,N_8311,N_8685);
and U13588 (N_13588,N_8765,N_7627);
nor U13589 (N_13589,N_6607,N_6107);
nand U13590 (N_13590,N_7043,N_8473);
xnor U13591 (N_13591,N_8155,N_7386);
and U13592 (N_13592,N_9591,N_7112);
nor U13593 (N_13593,N_9009,N_8358);
nor U13594 (N_13594,N_5365,N_6664);
nand U13595 (N_13595,N_9844,N_6210);
nand U13596 (N_13596,N_6901,N_7920);
and U13597 (N_13597,N_6884,N_5898);
and U13598 (N_13598,N_7275,N_6563);
nand U13599 (N_13599,N_9056,N_6389);
and U13600 (N_13600,N_5180,N_9620);
nand U13601 (N_13601,N_8190,N_7468);
and U13602 (N_13602,N_5026,N_8670);
or U13603 (N_13603,N_9915,N_9991);
nand U13604 (N_13604,N_6728,N_8806);
and U13605 (N_13605,N_8001,N_9146);
xnor U13606 (N_13606,N_9560,N_8233);
and U13607 (N_13607,N_9419,N_5453);
and U13608 (N_13608,N_9439,N_8963);
or U13609 (N_13609,N_7773,N_8851);
nand U13610 (N_13610,N_6631,N_5637);
nand U13611 (N_13611,N_9458,N_7793);
nand U13612 (N_13612,N_9313,N_6543);
or U13613 (N_13613,N_6051,N_7404);
or U13614 (N_13614,N_8873,N_9141);
and U13615 (N_13615,N_9164,N_7139);
xor U13616 (N_13616,N_7567,N_9428);
or U13617 (N_13617,N_5498,N_7972);
or U13618 (N_13618,N_5443,N_9073);
nor U13619 (N_13619,N_8953,N_8741);
nor U13620 (N_13620,N_5144,N_6168);
and U13621 (N_13621,N_5310,N_9393);
nor U13622 (N_13622,N_5767,N_9334);
xnor U13623 (N_13623,N_9371,N_8497);
nor U13624 (N_13624,N_6755,N_8549);
and U13625 (N_13625,N_9232,N_7163);
nand U13626 (N_13626,N_8889,N_6617);
nor U13627 (N_13627,N_6514,N_8650);
or U13628 (N_13628,N_8345,N_8153);
nor U13629 (N_13629,N_5226,N_5146);
nand U13630 (N_13630,N_7199,N_6415);
or U13631 (N_13631,N_9152,N_7030);
nand U13632 (N_13632,N_7984,N_7556);
nor U13633 (N_13633,N_5703,N_6597);
or U13634 (N_13634,N_7897,N_5187);
nor U13635 (N_13635,N_7390,N_9904);
or U13636 (N_13636,N_5674,N_9123);
or U13637 (N_13637,N_6628,N_8785);
nand U13638 (N_13638,N_5146,N_8780);
nor U13639 (N_13639,N_7119,N_7237);
nand U13640 (N_13640,N_9546,N_6123);
nand U13641 (N_13641,N_6183,N_6570);
nor U13642 (N_13642,N_8295,N_5213);
or U13643 (N_13643,N_6746,N_5658);
and U13644 (N_13644,N_5824,N_6802);
and U13645 (N_13645,N_5826,N_5231);
or U13646 (N_13646,N_8963,N_6785);
nand U13647 (N_13647,N_8642,N_5924);
or U13648 (N_13648,N_7579,N_6680);
or U13649 (N_13649,N_7784,N_9904);
and U13650 (N_13650,N_6908,N_7824);
nor U13651 (N_13651,N_9297,N_6495);
nand U13652 (N_13652,N_8787,N_7969);
or U13653 (N_13653,N_9582,N_7517);
nand U13654 (N_13654,N_8228,N_7979);
nand U13655 (N_13655,N_5422,N_8156);
nand U13656 (N_13656,N_6875,N_5437);
or U13657 (N_13657,N_8196,N_7009);
nor U13658 (N_13658,N_7095,N_8259);
xor U13659 (N_13659,N_6411,N_9201);
nor U13660 (N_13660,N_8151,N_8097);
or U13661 (N_13661,N_7373,N_7495);
nor U13662 (N_13662,N_6560,N_9016);
or U13663 (N_13663,N_5532,N_7547);
nor U13664 (N_13664,N_8378,N_9669);
or U13665 (N_13665,N_6250,N_8194);
nor U13666 (N_13666,N_9936,N_8868);
nand U13667 (N_13667,N_6149,N_8490);
and U13668 (N_13668,N_8776,N_8736);
nand U13669 (N_13669,N_9305,N_7945);
and U13670 (N_13670,N_5156,N_5015);
nor U13671 (N_13671,N_6893,N_6643);
or U13672 (N_13672,N_8465,N_7613);
and U13673 (N_13673,N_5915,N_9969);
nor U13674 (N_13674,N_5362,N_7011);
and U13675 (N_13675,N_8269,N_7824);
and U13676 (N_13676,N_7906,N_9992);
or U13677 (N_13677,N_7328,N_5521);
nor U13678 (N_13678,N_5441,N_6544);
and U13679 (N_13679,N_5327,N_6738);
xor U13680 (N_13680,N_8458,N_5683);
nor U13681 (N_13681,N_9810,N_8564);
xnor U13682 (N_13682,N_5579,N_7841);
or U13683 (N_13683,N_9994,N_7641);
nand U13684 (N_13684,N_7976,N_7139);
or U13685 (N_13685,N_8092,N_7204);
nor U13686 (N_13686,N_7988,N_5811);
nand U13687 (N_13687,N_6844,N_6917);
nor U13688 (N_13688,N_6237,N_6338);
nand U13689 (N_13689,N_8391,N_9884);
or U13690 (N_13690,N_6627,N_5463);
or U13691 (N_13691,N_8047,N_8725);
nand U13692 (N_13692,N_6817,N_6222);
nor U13693 (N_13693,N_9822,N_6540);
nor U13694 (N_13694,N_8778,N_7137);
xor U13695 (N_13695,N_8214,N_7598);
and U13696 (N_13696,N_7931,N_5259);
xnor U13697 (N_13697,N_5789,N_8407);
or U13698 (N_13698,N_8201,N_6573);
nand U13699 (N_13699,N_9896,N_9895);
or U13700 (N_13700,N_6745,N_5475);
and U13701 (N_13701,N_7123,N_8886);
or U13702 (N_13702,N_5852,N_6389);
and U13703 (N_13703,N_7402,N_5901);
and U13704 (N_13704,N_8746,N_8843);
nand U13705 (N_13705,N_8782,N_9837);
nand U13706 (N_13706,N_6348,N_5010);
or U13707 (N_13707,N_8513,N_8861);
and U13708 (N_13708,N_5585,N_8284);
nand U13709 (N_13709,N_5077,N_8054);
or U13710 (N_13710,N_6763,N_5613);
or U13711 (N_13711,N_5658,N_8470);
and U13712 (N_13712,N_5238,N_6944);
or U13713 (N_13713,N_9051,N_9128);
and U13714 (N_13714,N_8308,N_6047);
nor U13715 (N_13715,N_7950,N_6003);
nor U13716 (N_13716,N_8858,N_8266);
nor U13717 (N_13717,N_8458,N_7802);
nand U13718 (N_13718,N_8493,N_5150);
xor U13719 (N_13719,N_6298,N_8213);
or U13720 (N_13720,N_7514,N_9540);
nand U13721 (N_13721,N_9902,N_5243);
and U13722 (N_13722,N_6796,N_8320);
xnor U13723 (N_13723,N_5064,N_8978);
nand U13724 (N_13724,N_9914,N_9645);
nand U13725 (N_13725,N_8008,N_8526);
xor U13726 (N_13726,N_7971,N_6543);
nor U13727 (N_13727,N_5491,N_8858);
and U13728 (N_13728,N_8631,N_5742);
xor U13729 (N_13729,N_5239,N_8866);
nor U13730 (N_13730,N_9030,N_7566);
xnor U13731 (N_13731,N_6298,N_6796);
nor U13732 (N_13732,N_8767,N_6227);
and U13733 (N_13733,N_7804,N_8192);
nand U13734 (N_13734,N_8166,N_8046);
and U13735 (N_13735,N_8475,N_9761);
nand U13736 (N_13736,N_9188,N_5750);
and U13737 (N_13737,N_8456,N_8883);
nor U13738 (N_13738,N_5144,N_5821);
and U13739 (N_13739,N_8965,N_8709);
nand U13740 (N_13740,N_6444,N_9092);
nor U13741 (N_13741,N_9976,N_5235);
and U13742 (N_13742,N_9534,N_9795);
and U13743 (N_13743,N_7326,N_7855);
nand U13744 (N_13744,N_6643,N_5590);
and U13745 (N_13745,N_8646,N_5863);
xnor U13746 (N_13746,N_9609,N_9428);
and U13747 (N_13747,N_9229,N_7574);
nand U13748 (N_13748,N_6019,N_7754);
or U13749 (N_13749,N_8413,N_7616);
xor U13750 (N_13750,N_5788,N_5398);
nand U13751 (N_13751,N_8619,N_7428);
nor U13752 (N_13752,N_9158,N_9366);
or U13753 (N_13753,N_5929,N_6614);
and U13754 (N_13754,N_9786,N_5339);
nor U13755 (N_13755,N_9029,N_5930);
nand U13756 (N_13756,N_7898,N_7000);
and U13757 (N_13757,N_7999,N_7134);
nand U13758 (N_13758,N_7678,N_9644);
nor U13759 (N_13759,N_5451,N_7403);
or U13760 (N_13760,N_7165,N_9026);
nor U13761 (N_13761,N_9764,N_6609);
and U13762 (N_13762,N_5585,N_9321);
or U13763 (N_13763,N_6749,N_8950);
nand U13764 (N_13764,N_7575,N_7082);
nand U13765 (N_13765,N_9731,N_8676);
nor U13766 (N_13766,N_5666,N_8603);
nand U13767 (N_13767,N_6475,N_9636);
and U13768 (N_13768,N_7110,N_7791);
or U13769 (N_13769,N_7555,N_5637);
or U13770 (N_13770,N_8202,N_9906);
and U13771 (N_13771,N_8462,N_9803);
nand U13772 (N_13772,N_5172,N_5800);
nor U13773 (N_13773,N_7943,N_7838);
and U13774 (N_13774,N_7852,N_9345);
nand U13775 (N_13775,N_8025,N_6017);
nor U13776 (N_13776,N_8974,N_7266);
nand U13777 (N_13777,N_9155,N_9520);
nand U13778 (N_13778,N_8609,N_5480);
xnor U13779 (N_13779,N_6779,N_9555);
xor U13780 (N_13780,N_5971,N_8239);
nor U13781 (N_13781,N_5583,N_9177);
nand U13782 (N_13782,N_6611,N_6906);
and U13783 (N_13783,N_6586,N_8741);
nand U13784 (N_13784,N_8122,N_5593);
nor U13785 (N_13785,N_9919,N_5583);
nand U13786 (N_13786,N_9830,N_9128);
and U13787 (N_13787,N_9000,N_6428);
and U13788 (N_13788,N_5627,N_7966);
xnor U13789 (N_13789,N_6325,N_8073);
or U13790 (N_13790,N_8491,N_9119);
or U13791 (N_13791,N_5022,N_8566);
nor U13792 (N_13792,N_7820,N_7849);
nand U13793 (N_13793,N_5880,N_7758);
nand U13794 (N_13794,N_7209,N_7825);
nor U13795 (N_13795,N_7964,N_9804);
nor U13796 (N_13796,N_5969,N_9049);
and U13797 (N_13797,N_5880,N_6413);
and U13798 (N_13798,N_8685,N_5305);
nor U13799 (N_13799,N_6822,N_9537);
nor U13800 (N_13800,N_9018,N_5284);
nand U13801 (N_13801,N_8395,N_7289);
or U13802 (N_13802,N_9365,N_8812);
and U13803 (N_13803,N_8030,N_5936);
nand U13804 (N_13804,N_5959,N_6358);
or U13805 (N_13805,N_5856,N_7271);
nor U13806 (N_13806,N_8550,N_8463);
or U13807 (N_13807,N_9252,N_9978);
nor U13808 (N_13808,N_7654,N_8180);
and U13809 (N_13809,N_5999,N_6342);
nand U13810 (N_13810,N_6424,N_5282);
nor U13811 (N_13811,N_6513,N_5889);
xnor U13812 (N_13812,N_5494,N_6341);
nor U13813 (N_13813,N_9960,N_7944);
or U13814 (N_13814,N_6302,N_9459);
nand U13815 (N_13815,N_7093,N_7033);
and U13816 (N_13816,N_9689,N_7116);
nor U13817 (N_13817,N_8450,N_9703);
or U13818 (N_13818,N_5574,N_7783);
nand U13819 (N_13819,N_8226,N_9849);
xnor U13820 (N_13820,N_5476,N_5744);
nand U13821 (N_13821,N_9234,N_5138);
nor U13822 (N_13822,N_8280,N_8487);
nand U13823 (N_13823,N_5823,N_7184);
or U13824 (N_13824,N_9002,N_7829);
xnor U13825 (N_13825,N_9838,N_9353);
nor U13826 (N_13826,N_8125,N_9863);
and U13827 (N_13827,N_8648,N_9757);
nand U13828 (N_13828,N_6777,N_6701);
and U13829 (N_13829,N_9009,N_9558);
and U13830 (N_13830,N_6209,N_5956);
nor U13831 (N_13831,N_6375,N_6608);
or U13832 (N_13832,N_7428,N_7073);
nand U13833 (N_13833,N_7733,N_9684);
xor U13834 (N_13834,N_7582,N_6328);
nor U13835 (N_13835,N_6527,N_5581);
and U13836 (N_13836,N_7323,N_6596);
and U13837 (N_13837,N_9365,N_5640);
and U13838 (N_13838,N_5358,N_5095);
and U13839 (N_13839,N_7591,N_7693);
and U13840 (N_13840,N_7852,N_9384);
and U13841 (N_13841,N_8491,N_5680);
nor U13842 (N_13842,N_8633,N_7564);
nand U13843 (N_13843,N_6781,N_8246);
nand U13844 (N_13844,N_9150,N_6431);
and U13845 (N_13845,N_7790,N_6586);
nor U13846 (N_13846,N_5423,N_9549);
or U13847 (N_13847,N_9335,N_6403);
nor U13848 (N_13848,N_9276,N_8397);
or U13849 (N_13849,N_8898,N_8213);
nor U13850 (N_13850,N_7067,N_6923);
and U13851 (N_13851,N_9264,N_7580);
or U13852 (N_13852,N_7158,N_7835);
nor U13853 (N_13853,N_6875,N_9262);
nor U13854 (N_13854,N_7049,N_8380);
and U13855 (N_13855,N_9891,N_5326);
nor U13856 (N_13856,N_9525,N_6268);
and U13857 (N_13857,N_8310,N_5480);
nand U13858 (N_13858,N_7066,N_6624);
xor U13859 (N_13859,N_7747,N_9856);
nor U13860 (N_13860,N_5430,N_8503);
and U13861 (N_13861,N_6744,N_5062);
nand U13862 (N_13862,N_5459,N_9342);
nor U13863 (N_13863,N_5091,N_8196);
nand U13864 (N_13864,N_6986,N_5095);
nor U13865 (N_13865,N_9761,N_7357);
and U13866 (N_13866,N_7465,N_9377);
and U13867 (N_13867,N_6435,N_5824);
xor U13868 (N_13868,N_8243,N_8525);
nand U13869 (N_13869,N_6457,N_6432);
nor U13870 (N_13870,N_5256,N_6301);
nand U13871 (N_13871,N_8752,N_5746);
xnor U13872 (N_13872,N_9475,N_7585);
nand U13873 (N_13873,N_8238,N_9379);
and U13874 (N_13874,N_8968,N_9209);
nor U13875 (N_13875,N_6852,N_6211);
nand U13876 (N_13876,N_6741,N_5384);
nand U13877 (N_13877,N_5350,N_6320);
nor U13878 (N_13878,N_8374,N_8269);
and U13879 (N_13879,N_6647,N_5705);
nor U13880 (N_13880,N_6188,N_9909);
or U13881 (N_13881,N_8937,N_7125);
and U13882 (N_13882,N_5811,N_8604);
xnor U13883 (N_13883,N_7184,N_9196);
nor U13884 (N_13884,N_5534,N_8146);
or U13885 (N_13885,N_6620,N_6844);
or U13886 (N_13886,N_9862,N_5550);
xor U13887 (N_13887,N_7794,N_9684);
nor U13888 (N_13888,N_6539,N_5450);
nand U13889 (N_13889,N_9483,N_8332);
and U13890 (N_13890,N_9140,N_8790);
xor U13891 (N_13891,N_9255,N_5416);
or U13892 (N_13892,N_5515,N_9680);
or U13893 (N_13893,N_6281,N_5861);
and U13894 (N_13894,N_6180,N_8845);
nand U13895 (N_13895,N_6554,N_6845);
nor U13896 (N_13896,N_6136,N_9859);
and U13897 (N_13897,N_9437,N_8603);
nor U13898 (N_13898,N_6043,N_6323);
xor U13899 (N_13899,N_6664,N_9596);
nor U13900 (N_13900,N_7748,N_7155);
and U13901 (N_13901,N_9258,N_7769);
and U13902 (N_13902,N_8021,N_9959);
xor U13903 (N_13903,N_6807,N_8965);
nor U13904 (N_13904,N_9924,N_9517);
nand U13905 (N_13905,N_7271,N_8688);
or U13906 (N_13906,N_6780,N_7821);
nor U13907 (N_13907,N_7173,N_5778);
nor U13908 (N_13908,N_5137,N_8841);
or U13909 (N_13909,N_6607,N_5749);
xor U13910 (N_13910,N_9266,N_8913);
nand U13911 (N_13911,N_9239,N_8509);
nor U13912 (N_13912,N_6815,N_8940);
or U13913 (N_13913,N_9204,N_7409);
nand U13914 (N_13914,N_7629,N_9080);
or U13915 (N_13915,N_8976,N_7226);
and U13916 (N_13916,N_5588,N_6790);
or U13917 (N_13917,N_9675,N_5654);
and U13918 (N_13918,N_9317,N_9445);
and U13919 (N_13919,N_7357,N_5057);
nor U13920 (N_13920,N_6029,N_5836);
or U13921 (N_13921,N_9265,N_9589);
and U13922 (N_13922,N_5708,N_9528);
nor U13923 (N_13923,N_6465,N_9517);
nand U13924 (N_13924,N_8623,N_6228);
nor U13925 (N_13925,N_5235,N_5553);
nand U13926 (N_13926,N_5374,N_7315);
nand U13927 (N_13927,N_8955,N_5781);
or U13928 (N_13928,N_6262,N_7035);
xor U13929 (N_13929,N_6007,N_7225);
or U13930 (N_13930,N_9519,N_8368);
and U13931 (N_13931,N_6137,N_6157);
nor U13932 (N_13932,N_9647,N_6093);
or U13933 (N_13933,N_5271,N_7302);
or U13934 (N_13934,N_8506,N_7308);
nand U13935 (N_13935,N_9042,N_5390);
xor U13936 (N_13936,N_6195,N_9278);
nor U13937 (N_13937,N_9108,N_8073);
nor U13938 (N_13938,N_7548,N_8027);
nand U13939 (N_13939,N_5580,N_7797);
nor U13940 (N_13940,N_9722,N_8643);
nand U13941 (N_13941,N_8122,N_5500);
or U13942 (N_13942,N_7418,N_9720);
or U13943 (N_13943,N_7452,N_5024);
or U13944 (N_13944,N_5789,N_6763);
and U13945 (N_13945,N_5953,N_8220);
nor U13946 (N_13946,N_6994,N_7541);
and U13947 (N_13947,N_5987,N_8899);
and U13948 (N_13948,N_5068,N_5325);
and U13949 (N_13949,N_7873,N_8773);
and U13950 (N_13950,N_9001,N_5161);
nand U13951 (N_13951,N_9607,N_5922);
and U13952 (N_13952,N_8812,N_9655);
or U13953 (N_13953,N_6310,N_6682);
nor U13954 (N_13954,N_8924,N_8088);
and U13955 (N_13955,N_6579,N_7239);
nand U13956 (N_13956,N_5624,N_9716);
nand U13957 (N_13957,N_5973,N_9552);
or U13958 (N_13958,N_6645,N_9351);
nor U13959 (N_13959,N_5720,N_7587);
nor U13960 (N_13960,N_8205,N_8952);
xnor U13961 (N_13961,N_7923,N_5766);
and U13962 (N_13962,N_7662,N_5291);
nand U13963 (N_13963,N_7716,N_6209);
nand U13964 (N_13964,N_6867,N_5656);
nor U13965 (N_13965,N_9081,N_9526);
nor U13966 (N_13966,N_6053,N_9693);
nor U13967 (N_13967,N_5059,N_6096);
and U13968 (N_13968,N_9471,N_7314);
nor U13969 (N_13969,N_5381,N_8474);
nand U13970 (N_13970,N_7482,N_7882);
xor U13971 (N_13971,N_6236,N_8498);
and U13972 (N_13972,N_6060,N_6212);
nand U13973 (N_13973,N_9514,N_8119);
nand U13974 (N_13974,N_8568,N_5410);
nand U13975 (N_13975,N_9099,N_7156);
or U13976 (N_13976,N_7545,N_9158);
nand U13977 (N_13977,N_5540,N_7081);
nand U13978 (N_13978,N_8465,N_6763);
and U13979 (N_13979,N_9194,N_6871);
and U13980 (N_13980,N_5748,N_5371);
nor U13981 (N_13981,N_9157,N_8761);
or U13982 (N_13982,N_6848,N_6622);
and U13983 (N_13983,N_8589,N_5565);
or U13984 (N_13984,N_5975,N_6858);
or U13985 (N_13985,N_7115,N_6582);
nand U13986 (N_13986,N_6496,N_5610);
nand U13987 (N_13987,N_6450,N_8820);
nor U13988 (N_13988,N_8418,N_8834);
nand U13989 (N_13989,N_8170,N_9345);
nand U13990 (N_13990,N_7661,N_7240);
or U13991 (N_13991,N_5479,N_5465);
nand U13992 (N_13992,N_7508,N_5285);
and U13993 (N_13993,N_8220,N_6296);
nand U13994 (N_13994,N_9730,N_5256);
and U13995 (N_13995,N_8533,N_9416);
and U13996 (N_13996,N_8237,N_5984);
or U13997 (N_13997,N_6782,N_8557);
nand U13998 (N_13998,N_8450,N_7693);
xnor U13999 (N_13999,N_8844,N_6041);
and U14000 (N_14000,N_8416,N_7153);
and U14001 (N_14001,N_8468,N_6103);
or U14002 (N_14002,N_6346,N_7978);
nand U14003 (N_14003,N_9019,N_5672);
and U14004 (N_14004,N_8215,N_8214);
nand U14005 (N_14005,N_8030,N_8047);
nor U14006 (N_14006,N_9537,N_5544);
or U14007 (N_14007,N_8487,N_9181);
or U14008 (N_14008,N_6303,N_8296);
or U14009 (N_14009,N_7894,N_9227);
or U14010 (N_14010,N_6035,N_8646);
nor U14011 (N_14011,N_7417,N_7086);
and U14012 (N_14012,N_5746,N_9492);
nor U14013 (N_14013,N_6613,N_7230);
nand U14014 (N_14014,N_7617,N_5117);
xnor U14015 (N_14015,N_9254,N_5789);
and U14016 (N_14016,N_7708,N_7674);
nand U14017 (N_14017,N_9266,N_7395);
and U14018 (N_14018,N_5261,N_7420);
or U14019 (N_14019,N_6732,N_8713);
or U14020 (N_14020,N_9083,N_9319);
nand U14021 (N_14021,N_5348,N_6081);
nand U14022 (N_14022,N_9708,N_5898);
nor U14023 (N_14023,N_8945,N_8816);
and U14024 (N_14024,N_6211,N_7513);
and U14025 (N_14025,N_8716,N_9824);
nand U14026 (N_14026,N_8094,N_5982);
nor U14027 (N_14027,N_7676,N_7841);
nand U14028 (N_14028,N_5999,N_7226);
nand U14029 (N_14029,N_7068,N_6641);
nand U14030 (N_14030,N_9306,N_8090);
nand U14031 (N_14031,N_6606,N_5913);
and U14032 (N_14032,N_7679,N_6387);
and U14033 (N_14033,N_8192,N_7316);
or U14034 (N_14034,N_7168,N_5021);
and U14035 (N_14035,N_9778,N_5191);
xnor U14036 (N_14036,N_6333,N_7737);
and U14037 (N_14037,N_9616,N_7208);
or U14038 (N_14038,N_6494,N_6370);
nand U14039 (N_14039,N_6207,N_9181);
and U14040 (N_14040,N_8936,N_8650);
xnor U14041 (N_14041,N_6366,N_6919);
nand U14042 (N_14042,N_8641,N_9151);
and U14043 (N_14043,N_6378,N_6823);
xnor U14044 (N_14044,N_5279,N_6847);
nor U14045 (N_14045,N_7559,N_6996);
and U14046 (N_14046,N_5208,N_5369);
nand U14047 (N_14047,N_9595,N_8869);
nor U14048 (N_14048,N_7877,N_7333);
nand U14049 (N_14049,N_7822,N_6772);
nand U14050 (N_14050,N_5495,N_9741);
and U14051 (N_14051,N_7322,N_6099);
nor U14052 (N_14052,N_8333,N_9047);
nand U14053 (N_14053,N_5278,N_9177);
nand U14054 (N_14054,N_5475,N_5163);
nor U14055 (N_14055,N_9225,N_8634);
nand U14056 (N_14056,N_9677,N_5045);
nand U14057 (N_14057,N_8351,N_7637);
or U14058 (N_14058,N_5962,N_6780);
nor U14059 (N_14059,N_5160,N_9863);
and U14060 (N_14060,N_7716,N_5352);
or U14061 (N_14061,N_5256,N_7397);
nand U14062 (N_14062,N_5931,N_9463);
and U14063 (N_14063,N_9526,N_6033);
nand U14064 (N_14064,N_8383,N_9124);
nand U14065 (N_14065,N_7799,N_8414);
nor U14066 (N_14066,N_9964,N_6184);
nor U14067 (N_14067,N_5945,N_8788);
or U14068 (N_14068,N_9146,N_7694);
nor U14069 (N_14069,N_7120,N_7650);
nand U14070 (N_14070,N_8567,N_8766);
nand U14071 (N_14071,N_9474,N_9030);
nor U14072 (N_14072,N_8101,N_5721);
and U14073 (N_14073,N_7739,N_6101);
nand U14074 (N_14074,N_5495,N_7890);
and U14075 (N_14075,N_5254,N_9488);
and U14076 (N_14076,N_8710,N_7198);
nand U14077 (N_14077,N_8343,N_5873);
nand U14078 (N_14078,N_5386,N_9403);
or U14079 (N_14079,N_7358,N_8756);
and U14080 (N_14080,N_5140,N_5946);
or U14081 (N_14081,N_7658,N_9957);
nor U14082 (N_14082,N_8881,N_6962);
or U14083 (N_14083,N_7381,N_7455);
or U14084 (N_14084,N_6333,N_5393);
nand U14085 (N_14085,N_5774,N_8252);
and U14086 (N_14086,N_5802,N_9902);
or U14087 (N_14087,N_8815,N_8669);
or U14088 (N_14088,N_9542,N_5251);
xnor U14089 (N_14089,N_9768,N_6872);
nand U14090 (N_14090,N_5543,N_5134);
nor U14091 (N_14091,N_9696,N_8258);
and U14092 (N_14092,N_9223,N_5264);
nor U14093 (N_14093,N_9404,N_6937);
and U14094 (N_14094,N_5232,N_9473);
and U14095 (N_14095,N_9419,N_6359);
or U14096 (N_14096,N_8650,N_7124);
or U14097 (N_14097,N_6011,N_8205);
and U14098 (N_14098,N_9203,N_5185);
and U14099 (N_14099,N_9100,N_6673);
and U14100 (N_14100,N_7776,N_9370);
xor U14101 (N_14101,N_7425,N_5792);
and U14102 (N_14102,N_8603,N_8280);
nor U14103 (N_14103,N_8574,N_5634);
and U14104 (N_14104,N_7153,N_9121);
and U14105 (N_14105,N_9232,N_7038);
nand U14106 (N_14106,N_8126,N_5167);
nor U14107 (N_14107,N_6732,N_9085);
or U14108 (N_14108,N_6087,N_5515);
or U14109 (N_14109,N_5607,N_6381);
or U14110 (N_14110,N_7721,N_5015);
and U14111 (N_14111,N_9232,N_6109);
xor U14112 (N_14112,N_8316,N_6190);
or U14113 (N_14113,N_7386,N_7464);
and U14114 (N_14114,N_8057,N_7269);
xnor U14115 (N_14115,N_5376,N_5458);
and U14116 (N_14116,N_7068,N_8497);
xnor U14117 (N_14117,N_5617,N_7248);
nor U14118 (N_14118,N_6466,N_8418);
and U14119 (N_14119,N_6210,N_6818);
nand U14120 (N_14120,N_9673,N_5691);
nor U14121 (N_14121,N_6563,N_5654);
or U14122 (N_14122,N_6576,N_6716);
or U14123 (N_14123,N_9108,N_5504);
nand U14124 (N_14124,N_7220,N_8744);
xnor U14125 (N_14125,N_8781,N_5293);
nor U14126 (N_14126,N_5310,N_6976);
nand U14127 (N_14127,N_8462,N_9154);
or U14128 (N_14128,N_5668,N_5515);
xnor U14129 (N_14129,N_9555,N_6411);
and U14130 (N_14130,N_8280,N_8955);
and U14131 (N_14131,N_9742,N_9392);
or U14132 (N_14132,N_5091,N_7566);
or U14133 (N_14133,N_5279,N_8943);
nor U14134 (N_14134,N_7753,N_9090);
or U14135 (N_14135,N_6994,N_9585);
or U14136 (N_14136,N_9263,N_8303);
nand U14137 (N_14137,N_5403,N_7763);
nor U14138 (N_14138,N_8984,N_5828);
nand U14139 (N_14139,N_9030,N_8991);
nand U14140 (N_14140,N_7883,N_8413);
or U14141 (N_14141,N_9759,N_7587);
and U14142 (N_14142,N_7678,N_8134);
and U14143 (N_14143,N_9679,N_5047);
and U14144 (N_14144,N_7011,N_6332);
and U14145 (N_14145,N_5917,N_5543);
nand U14146 (N_14146,N_5542,N_8827);
nor U14147 (N_14147,N_8243,N_9697);
nor U14148 (N_14148,N_6789,N_6045);
and U14149 (N_14149,N_5730,N_6522);
nand U14150 (N_14150,N_6448,N_8423);
xor U14151 (N_14151,N_9857,N_8810);
nor U14152 (N_14152,N_8873,N_5116);
nand U14153 (N_14153,N_9852,N_6244);
nand U14154 (N_14154,N_7736,N_8316);
or U14155 (N_14155,N_5761,N_9884);
and U14156 (N_14156,N_6549,N_5623);
and U14157 (N_14157,N_5330,N_9808);
and U14158 (N_14158,N_6780,N_8954);
or U14159 (N_14159,N_7852,N_9654);
and U14160 (N_14160,N_6472,N_9525);
nor U14161 (N_14161,N_8428,N_6249);
and U14162 (N_14162,N_6506,N_6143);
or U14163 (N_14163,N_7684,N_8708);
nand U14164 (N_14164,N_7090,N_8862);
or U14165 (N_14165,N_7381,N_9979);
or U14166 (N_14166,N_8836,N_9097);
xor U14167 (N_14167,N_7801,N_8893);
nor U14168 (N_14168,N_5337,N_6133);
or U14169 (N_14169,N_8634,N_6852);
nand U14170 (N_14170,N_8765,N_7254);
or U14171 (N_14171,N_9288,N_8240);
or U14172 (N_14172,N_6627,N_8027);
nor U14173 (N_14173,N_7529,N_6023);
and U14174 (N_14174,N_6067,N_6614);
xnor U14175 (N_14175,N_9264,N_5837);
or U14176 (N_14176,N_6006,N_7102);
or U14177 (N_14177,N_8200,N_6821);
or U14178 (N_14178,N_7147,N_6052);
nor U14179 (N_14179,N_8355,N_9527);
nand U14180 (N_14180,N_7286,N_8453);
nor U14181 (N_14181,N_7550,N_5591);
nor U14182 (N_14182,N_7770,N_5092);
nor U14183 (N_14183,N_7651,N_7626);
nor U14184 (N_14184,N_6322,N_6737);
xor U14185 (N_14185,N_6088,N_5852);
and U14186 (N_14186,N_8926,N_7335);
nor U14187 (N_14187,N_6311,N_6117);
nand U14188 (N_14188,N_6285,N_5695);
or U14189 (N_14189,N_6677,N_7545);
xnor U14190 (N_14190,N_9943,N_9169);
and U14191 (N_14191,N_7519,N_8578);
and U14192 (N_14192,N_7251,N_6106);
nor U14193 (N_14193,N_9677,N_9523);
nand U14194 (N_14194,N_9325,N_7577);
xnor U14195 (N_14195,N_5691,N_8105);
or U14196 (N_14196,N_8142,N_8736);
nand U14197 (N_14197,N_5066,N_8326);
and U14198 (N_14198,N_9763,N_7797);
or U14199 (N_14199,N_6356,N_6874);
nand U14200 (N_14200,N_7973,N_7120);
and U14201 (N_14201,N_5061,N_7180);
nor U14202 (N_14202,N_9043,N_7546);
xnor U14203 (N_14203,N_9529,N_6938);
or U14204 (N_14204,N_8329,N_8573);
or U14205 (N_14205,N_6762,N_6913);
nor U14206 (N_14206,N_6326,N_5167);
nor U14207 (N_14207,N_6843,N_7935);
nand U14208 (N_14208,N_8200,N_7127);
and U14209 (N_14209,N_9545,N_6009);
and U14210 (N_14210,N_8313,N_9267);
and U14211 (N_14211,N_5408,N_7211);
and U14212 (N_14212,N_5530,N_9990);
or U14213 (N_14213,N_5145,N_6676);
nand U14214 (N_14214,N_8889,N_5621);
nor U14215 (N_14215,N_8355,N_7559);
nor U14216 (N_14216,N_9710,N_9238);
nand U14217 (N_14217,N_7773,N_7793);
nor U14218 (N_14218,N_8120,N_5855);
nor U14219 (N_14219,N_7410,N_8794);
nor U14220 (N_14220,N_9121,N_8185);
and U14221 (N_14221,N_5751,N_9304);
nor U14222 (N_14222,N_7622,N_9608);
nand U14223 (N_14223,N_5357,N_5841);
or U14224 (N_14224,N_8524,N_9264);
nand U14225 (N_14225,N_5478,N_6588);
nand U14226 (N_14226,N_6572,N_7951);
nor U14227 (N_14227,N_9337,N_6545);
nor U14228 (N_14228,N_6637,N_6809);
and U14229 (N_14229,N_9989,N_9440);
or U14230 (N_14230,N_9822,N_6661);
nor U14231 (N_14231,N_8052,N_5512);
nand U14232 (N_14232,N_8305,N_8622);
and U14233 (N_14233,N_9416,N_9362);
xnor U14234 (N_14234,N_5727,N_5849);
or U14235 (N_14235,N_7800,N_9945);
or U14236 (N_14236,N_5797,N_5753);
nor U14237 (N_14237,N_6847,N_6294);
nor U14238 (N_14238,N_6755,N_6643);
nor U14239 (N_14239,N_6914,N_7808);
and U14240 (N_14240,N_8636,N_5279);
and U14241 (N_14241,N_5228,N_6936);
nand U14242 (N_14242,N_9869,N_6656);
xnor U14243 (N_14243,N_7219,N_9712);
nand U14244 (N_14244,N_7406,N_8065);
nand U14245 (N_14245,N_9393,N_8931);
xor U14246 (N_14246,N_8743,N_9673);
nand U14247 (N_14247,N_9125,N_7589);
and U14248 (N_14248,N_8804,N_6906);
nor U14249 (N_14249,N_6657,N_7547);
nand U14250 (N_14250,N_7333,N_7086);
or U14251 (N_14251,N_8051,N_6892);
or U14252 (N_14252,N_9031,N_8722);
nor U14253 (N_14253,N_8892,N_6088);
and U14254 (N_14254,N_7219,N_8481);
nor U14255 (N_14255,N_7439,N_7149);
and U14256 (N_14256,N_8972,N_5111);
nand U14257 (N_14257,N_5013,N_9938);
nand U14258 (N_14258,N_7471,N_9333);
or U14259 (N_14259,N_7147,N_5896);
xnor U14260 (N_14260,N_7326,N_9438);
and U14261 (N_14261,N_7212,N_7299);
nand U14262 (N_14262,N_8009,N_5941);
nand U14263 (N_14263,N_8096,N_6553);
nor U14264 (N_14264,N_6555,N_8622);
nor U14265 (N_14265,N_5055,N_8298);
nand U14266 (N_14266,N_6899,N_9170);
nand U14267 (N_14267,N_5228,N_6308);
and U14268 (N_14268,N_7983,N_9816);
and U14269 (N_14269,N_5080,N_7091);
nand U14270 (N_14270,N_5372,N_9600);
nor U14271 (N_14271,N_7160,N_8543);
xor U14272 (N_14272,N_9766,N_9253);
and U14273 (N_14273,N_7387,N_6920);
nor U14274 (N_14274,N_9266,N_8987);
and U14275 (N_14275,N_5131,N_9005);
and U14276 (N_14276,N_5110,N_6743);
nor U14277 (N_14277,N_7258,N_8642);
and U14278 (N_14278,N_8341,N_7023);
xnor U14279 (N_14279,N_8081,N_5987);
nand U14280 (N_14280,N_6943,N_6780);
and U14281 (N_14281,N_9431,N_6164);
or U14282 (N_14282,N_9238,N_9913);
nand U14283 (N_14283,N_7974,N_6697);
nor U14284 (N_14284,N_8132,N_6439);
nand U14285 (N_14285,N_9422,N_7013);
or U14286 (N_14286,N_6372,N_8626);
or U14287 (N_14287,N_9925,N_6498);
nor U14288 (N_14288,N_9196,N_7220);
nor U14289 (N_14289,N_6997,N_6238);
and U14290 (N_14290,N_7663,N_6928);
nand U14291 (N_14291,N_9137,N_6966);
or U14292 (N_14292,N_7207,N_6984);
and U14293 (N_14293,N_5345,N_5989);
xor U14294 (N_14294,N_9010,N_6552);
and U14295 (N_14295,N_8406,N_7023);
nand U14296 (N_14296,N_6838,N_7991);
nor U14297 (N_14297,N_5166,N_6678);
nand U14298 (N_14298,N_5426,N_6164);
nand U14299 (N_14299,N_7431,N_8620);
or U14300 (N_14300,N_7407,N_8398);
nor U14301 (N_14301,N_6733,N_7468);
nor U14302 (N_14302,N_6227,N_7017);
nor U14303 (N_14303,N_6571,N_6026);
nor U14304 (N_14304,N_6564,N_9674);
nand U14305 (N_14305,N_6414,N_5321);
nor U14306 (N_14306,N_6125,N_8648);
nor U14307 (N_14307,N_7064,N_5996);
or U14308 (N_14308,N_7252,N_6448);
and U14309 (N_14309,N_9014,N_5861);
or U14310 (N_14310,N_6374,N_7034);
nor U14311 (N_14311,N_7659,N_9635);
and U14312 (N_14312,N_5741,N_5327);
or U14313 (N_14313,N_5423,N_7391);
and U14314 (N_14314,N_6710,N_6678);
or U14315 (N_14315,N_6168,N_7574);
nor U14316 (N_14316,N_7222,N_6564);
nand U14317 (N_14317,N_9083,N_6846);
or U14318 (N_14318,N_8414,N_5418);
nand U14319 (N_14319,N_5677,N_6818);
xnor U14320 (N_14320,N_7868,N_6058);
xnor U14321 (N_14321,N_5815,N_6019);
nand U14322 (N_14322,N_8856,N_6656);
nor U14323 (N_14323,N_9243,N_7367);
nor U14324 (N_14324,N_8058,N_5784);
and U14325 (N_14325,N_8147,N_9706);
nor U14326 (N_14326,N_6668,N_6319);
xor U14327 (N_14327,N_9312,N_9574);
xor U14328 (N_14328,N_6216,N_5158);
nor U14329 (N_14329,N_7942,N_6712);
nor U14330 (N_14330,N_8388,N_5367);
or U14331 (N_14331,N_9936,N_5791);
nor U14332 (N_14332,N_6228,N_8921);
nand U14333 (N_14333,N_5206,N_7468);
nand U14334 (N_14334,N_9457,N_8474);
nand U14335 (N_14335,N_5903,N_6581);
nor U14336 (N_14336,N_6750,N_7199);
or U14337 (N_14337,N_9518,N_6356);
or U14338 (N_14338,N_9055,N_5939);
nor U14339 (N_14339,N_8293,N_6889);
and U14340 (N_14340,N_9363,N_6996);
nor U14341 (N_14341,N_8733,N_5128);
nor U14342 (N_14342,N_8119,N_7457);
nand U14343 (N_14343,N_7818,N_9933);
or U14344 (N_14344,N_6789,N_6320);
nand U14345 (N_14345,N_7861,N_9500);
or U14346 (N_14346,N_6607,N_9694);
and U14347 (N_14347,N_7834,N_7705);
and U14348 (N_14348,N_6066,N_8496);
or U14349 (N_14349,N_6642,N_9551);
and U14350 (N_14350,N_6728,N_7270);
nand U14351 (N_14351,N_6588,N_8397);
nand U14352 (N_14352,N_8634,N_9995);
nand U14353 (N_14353,N_5926,N_8855);
and U14354 (N_14354,N_5829,N_7062);
nor U14355 (N_14355,N_7819,N_5117);
and U14356 (N_14356,N_7506,N_8828);
nand U14357 (N_14357,N_8695,N_8477);
nor U14358 (N_14358,N_5128,N_6079);
or U14359 (N_14359,N_7561,N_8633);
or U14360 (N_14360,N_6564,N_8739);
nand U14361 (N_14361,N_8651,N_8630);
nor U14362 (N_14362,N_5221,N_5989);
and U14363 (N_14363,N_9276,N_5868);
nor U14364 (N_14364,N_8104,N_5711);
nor U14365 (N_14365,N_7581,N_6847);
nor U14366 (N_14366,N_5376,N_6104);
or U14367 (N_14367,N_5028,N_8174);
or U14368 (N_14368,N_9602,N_9311);
and U14369 (N_14369,N_6259,N_9171);
nor U14370 (N_14370,N_9932,N_7715);
and U14371 (N_14371,N_8738,N_9434);
nand U14372 (N_14372,N_8858,N_9672);
or U14373 (N_14373,N_6988,N_8723);
nor U14374 (N_14374,N_5088,N_9228);
nor U14375 (N_14375,N_8396,N_7481);
nor U14376 (N_14376,N_6709,N_7369);
or U14377 (N_14377,N_6574,N_8482);
nor U14378 (N_14378,N_8621,N_8658);
and U14379 (N_14379,N_5908,N_6260);
nand U14380 (N_14380,N_6909,N_8470);
and U14381 (N_14381,N_6435,N_8649);
and U14382 (N_14382,N_7157,N_8212);
nor U14383 (N_14383,N_7108,N_8308);
xnor U14384 (N_14384,N_7233,N_9749);
xor U14385 (N_14385,N_9050,N_8199);
nand U14386 (N_14386,N_9388,N_9424);
nand U14387 (N_14387,N_6225,N_8480);
nor U14388 (N_14388,N_8144,N_5136);
or U14389 (N_14389,N_7825,N_8736);
or U14390 (N_14390,N_6911,N_9121);
nor U14391 (N_14391,N_6972,N_6116);
nor U14392 (N_14392,N_7930,N_8726);
or U14393 (N_14393,N_6420,N_8861);
nor U14394 (N_14394,N_8850,N_6698);
and U14395 (N_14395,N_9818,N_9514);
nand U14396 (N_14396,N_9787,N_8579);
and U14397 (N_14397,N_7259,N_8575);
or U14398 (N_14398,N_7271,N_8490);
and U14399 (N_14399,N_7111,N_5841);
nor U14400 (N_14400,N_6636,N_8449);
and U14401 (N_14401,N_8506,N_9302);
nor U14402 (N_14402,N_7815,N_6005);
or U14403 (N_14403,N_5627,N_6430);
nand U14404 (N_14404,N_8751,N_9958);
or U14405 (N_14405,N_8785,N_6860);
nor U14406 (N_14406,N_8215,N_9765);
nand U14407 (N_14407,N_6152,N_7319);
or U14408 (N_14408,N_8227,N_7444);
xnor U14409 (N_14409,N_5839,N_8764);
nor U14410 (N_14410,N_5898,N_7123);
xnor U14411 (N_14411,N_8635,N_8070);
nor U14412 (N_14412,N_9189,N_8493);
or U14413 (N_14413,N_5895,N_9971);
and U14414 (N_14414,N_8287,N_5249);
nor U14415 (N_14415,N_6928,N_9383);
xnor U14416 (N_14416,N_5179,N_7222);
and U14417 (N_14417,N_6523,N_6901);
nor U14418 (N_14418,N_6029,N_9916);
or U14419 (N_14419,N_5771,N_8002);
or U14420 (N_14420,N_6194,N_9052);
or U14421 (N_14421,N_9860,N_5546);
nand U14422 (N_14422,N_6692,N_7482);
and U14423 (N_14423,N_8633,N_8590);
nor U14424 (N_14424,N_6214,N_5133);
or U14425 (N_14425,N_6571,N_9508);
or U14426 (N_14426,N_8639,N_8731);
or U14427 (N_14427,N_9508,N_6791);
nand U14428 (N_14428,N_5268,N_8554);
or U14429 (N_14429,N_6860,N_5688);
xnor U14430 (N_14430,N_6068,N_6042);
xnor U14431 (N_14431,N_5957,N_8246);
nand U14432 (N_14432,N_6852,N_5130);
nand U14433 (N_14433,N_6468,N_7441);
or U14434 (N_14434,N_8270,N_5533);
or U14435 (N_14435,N_7900,N_8955);
and U14436 (N_14436,N_6658,N_9226);
or U14437 (N_14437,N_9988,N_8234);
nor U14438 (N_14438,N_5232,N_5351);
and U14439 (N_14439,N_9718,N_8007);
or U14440 (N_14440,N_8013,N_5003);
nand U14441 (N_14441,N_8753,N_8469);
nor U14442 (N_14442,N_8819,N_5349);
or U14443 (N_14443,N_9753,N_9532);
nand U14444 (N_14444,N_8862,N_9641);
xor U14445 (N_14445,N_6684,N_6619);
nor U14446 (N_14446,N_5253,N_9540);
or U14447 (N_14447,N_6396,N_6566);
nand U14448 (N_14448,N_6363,N_8779);
and U14449 (N_14449,N_5752,N_7078);
or U14450 (N_14450,N_8939,N_8388);
and U14451 (N_14451,N_5517,N_5372);
or U14452 (N_14452,N_7034,N_9398);
nand U14453 (N_14453,N_6032,N_5859);
or U14454 (N_14454,N_7253,N_5341);
or U14455 (N_14455,N_6219,N_8386);
nand U14456 (N_14456,N_8169,N_7421);
and U14457 (N_14457,N_9192,N_6814);
and U14458 (N_14458,N_7644,N_6236);
and U14459 (N_14459,N_8113,N_9521);
nor U14460 (N_14460,N_9454,N_9003);
nand U14461 (N_14461,N_9242,N_9524);
nand U14462 (N_14462,N_5108,N_5496);
or U14463 (N_14463,N_6905,N_6669);
nor U14464 (N_14464,N_9010,N_6886);
nor U14465 (N_14465,N_7836,N_9539);
nor U14466 (N_14466,N_6488,N_6231);
and U14467 (N_14467,N_6692,N_7227);
nor U14468 (N_14468,N_9668,N_7017);
or U14469 (N_14469,N_6321,N_8761);
nand U14470 (N_14470,N_7762,N_6796);
or U14471 (N_14471,N_6121,N_5957);
nand U14472 (N_14472,N_7970,N_7908);
or U14473 (N_14473,N_9134,N_5269);
or U14474 (N_14474,N_8614,N_7971);
and U14475 (N_14475,N_5194,N_7725);
or U14476 (N_14476,N_9523,N_5540);
or U14477 (N_14477,N_6280,N_8913);
xor U14478 (N_14478,N_6098,N_9052);
and U14479 (N_14479,N_9703,N_7786);
nand U14480 (N_14480,N_8061,N_7788);
nand U14481 (N_14481,N_8808,N_5271);
or U14482 (N_14482,N_6283,N_7048);
nor U14483 (N_14483,N_9430,N_9258);
and U14484 (N_14484,N_7987,N_5803);
nor U14485 (N_14485,N_9527,N_6444);
nand U14486 (N_14486,N_8243,N_5809);
nand U14487 (N_14487,N_6865,N_7051);
nand U14488 (N_14488,N_7286,N_6493);
nand U14489 (N_14489,N_5708,N_5892);
and U14490 (N_14490,N_8039,N_6398);
nor U14491 (N_14491,N_9549,N_5825);
nand U14492 (N_14492,N_5915,N_9788);
xor U14493 (N_14493,N_9923,N_9398);
nand U14494 (N_14494,N_5525,N_8288);
and U14495 (N_14495,N_8892,N_5663);
nor U14496 (N_14496,N_9693,N_5068);
nor U14497 (N_14497,N_8625,N_8291);
nand U14498 (N_14498,N_9775,N_7368);
nand U14499 (N_14499,N_5404,N_7421);
and U14500 (N_14500,N_6941,N_8042);
nand U14501 (N_14501,N_8125,N_6472);
or U14502 (N_14502,N_9713,N_6457);
nand U14503 (N_14503,N_9560,N_7938);
xor U14504 (N_14504,N_6765,N_7547);
nand U14505 (N_14505,N_6640,N_9624);
and U14506 (N_14506,N_5734,N_9238);
nand U14507 (N_14507,N_7312,N_9610);
or U14508 (N_14508,N_5393,N_8437);
and U14509 (N_14509,N_8922,N_9504);
or U14510 (N_14510,N_6374,N_7640);
and U14511 (N_14511,N_9948,N_9560);
nor U14512 (N_14512,N_6345,N_9964);
and U14513 (N_14513,N_7748,N_9383);
nand U14514 (N_14514,N_8193,N_5429);
nor U14515 (N_14515,N_8521,N_9870);
or U14516 (N_14516,N_6650,N_6569);
nor U14517 (N_14517,N_8726,N_9811);
nand U14518 (N_14518,N_5897,N_5862);
nor U14519 (N_14519,N_9676,N_6236);
or U14520 (N_14520,N_7310,N_7372);
and U14521 (N_14521,N_8005,N_6149);
nand U14522 (N_14522,N_6253,N_7845);
or U14523 (N_14523,N_5895,N_7996);
nand U14524 (N_14524,N_8544,N_6661);
nor U14525 (N_14525,N_5917,N_8762);
nand U14526 (N_14526,N_9259,N_7771);
or U14527 (N_14527,N_7506,N_6552);
nand U14528 (N_14528,N_9828,N_7155);
nor U14529 (N_14529,N_8225,N_5580);
or U14530 (N_14530,N_6597,N_7559);
nor U14531 (N_14531,N_5936,N_9931);
nor U14532 (N_14532,N_8329,N_8291);
nand U14533 (N_14533,N_7793,N_7493);
or U14534 (N_14534,N_8177,N_8441);
xor U14535 (N_14535,N_5490,N_7905);
or U14536 (N_14536,N_7607,N_8669);
xnor U14537 (N_14537,N_8936,N_7755);
nor U14538 (N_14538,N_5085,N_6927);
and U14539 (N_14539,N_7003,N_9856);
nand U14540 (N_14540,N_7811,N_5779);
and U14541 (N_14541,N_6220,N_5323);
or U14542 (N_14542,N_5235,N_9131);
nand U14543 (N_14543,N_9780,N_6178);
or U14544 (N_14544,N_6556,N_8239);
nand U14545 (N_14545,N_6367,N_9333);
nand U14546 (N_14546,N_6948,N_9393);
nand U14547 (N_14547,N_7325,N_8904);
or U14548 (N_14548,N_7791,N_7714);
or U14549 (N_14549,N_6317,N_5171);
or U14550 (N_14550,N_7618,N_7581);
or U14551 (N_14551,N_9762,N_9108);
and U14552 (N_14552,N_5330,N_8482);
nor U14553 (N_14553,N_6489,N_6853);
xnor U14554 (N_14554,N_9411,N_7139);
nand U14555 (N_14555,N_9472,N_7937);
nor U14556 (N_14556,N_8405,N_7408);
or U14557 (N_14557,N_8556,N_5745);
nor U14558 (N_14558,N_9219,N_5780);
nand U14559 (N_14559,N_9658,N_9684);
nor U14560 (N_14560,N_7499,N_6269);
and U14561 (N_14561,N_9118,N_6375);
and U14562 (N_14562,N_8049,N_6342);
xnor U14563 (N_14563,N_7706,N_6469);
or U14564 (N_14564,N_8331,N_8719);
nor U14565 (N_14565,N_9763,N_7694);
or U14566 (N_14566,N_5711,N_9358);
and U14567 (N_14567,N_8862,N_5321);
nor U14568 (N_14568,N_8270,N_5166);
nand U14569 (N_14569,N_9236,N_6054);
xnor U14570 (N_14570,N_8633,N_5845);
nand U14571 (N_14571,N_6745,N_6523);
nand U14572 (N_14572,N_5847,N_9714);
or U14573 (N_14573,N_6348,N_6793);
and U14574 (N_14574,N_5763,N_5322);
nand U14575 (N_14575,N_5321,N_5541);
or U14576 (N_14576,N_8326,N_5217);
nand U14577 (N_14577,N_8925,N_9591);
nand U14578 (N_14578,N_8044,N_5631);
nand U14579 (N_14579,N_5046,N_5797);
and U14580 (N_14580,N_6951,N_7627);
xnor U14581 (N_14581,N_7643,N_7702);
and U14582 (N_14582,N_7340,N_9968);
nor U14583 (N_14583,N_9616,N_8545);
nor U14584 (N_14584,N_6480,N_7487);
and U14585 (N_14585,N_9482,N_6978);
or U14586 (N_14586,N_7905,N_9225);
and U14587 (N_14587,N_8718,N_7558);
nand U14588 (N_14588,N_6207,N_5789);
nand U14589 (N_14589,N_6987,N_8020);
nand U14590 (N_14590,N_8621,N_7333);
nor U14591 (N_14591,N_9987,N_8215);
nor U14592 (N_14592,N_9820,N_5256);
nand U14593 (N_14593,N_9453,N_6171);
xnor U14594 (N_14594,N_7127,N_7034);
or U14595 (N_14595,N_8195,N_7197);
or U14596 (N_14596,N_7578,N_6789);
nand U14597 (N_14597,N_5102,N_5611);
or U14598 (N_14598,N_6037,N_6912);
nor U14599 (N_14599,N_6165,N_7583);
xnor U14600 (N_14600,N_6340,N_6375);
and U14601 (N_14601,N_6739,N_5550);
nand U14602 (N_14602,N_6569,N_7806);
xor U14603 (N_14603,N_5628,N_6958);
or U14604 (N_14604,N_8184,N_6987);
and U14605 (N_14605,N_5472,N_5650);
nand U14606 (N_14606,N_7539,N_9360);
nor U14607 (N_14607,N_9585,N_7294);
nand U14608 (N_14608,N_8254,N_9642);
nand U14609 (N_14609,N_8877,N_5645);
xor U14610 (N_14610,N_7696,N_7409);
or U14611 (N_14611,N_6963,N_8161);
nand U14612 (N_14612,N_8753,N_7190);
nand U14613 (N_14613,N_7235,N_6999);
nand U14614 (N_14614,N_5160,N_8530);
and U14615 (N_14615,N_5287,N_8381);
and U14616 (N_14616,N_7863,N_9914);
nand U14617 (N_14617,N_5361,N_9930);
nand U14618 (N_14618,N_6871,N_9875);
nor U14619 (N_14619,N_8627,N_9308);
or U14620 (N_14620,N_6512,N_7740);
xor U14621 (N_14621,N_9792,N_7702);
nor U14622 (N_14622,N_5574,N_7423);
or U14623 (N_14623,N_7822,N_5073);
nand U14624 (N_14624,N_8675,N_5208);
nor U14625 (N_14625,N_6439,N_5831);
nor U14626 (N_14626,N_6542,N_6182);
and U14627 (N_14627,N_7443,N_5512);
nand U14628 (N_14628,N_5968,N_7679);
nor U14629 (N_14629,N_5356,N_6726);
nand U14630 (N_14630,N_8396,N_9467);
and U14631 (N_14631,N_7700,N_7682);
and U14632 (N_14632,N_8447,N_6211);
nor U14633 (N_14633,N_5526,N_6993);
and U14634 (N_14634,N_7066,N_8422);
or U14635 (N_14635,N_7189,N_9470);
nand U14636 (N_14636,N_8416,N_6974);
nor U14637 (N_14637,N_7978,N_9589);
xor U14638 (N_14638,N_8691,N_6193);
and U14639 (N_14639,N_6698,N_5385);
and U14640 (N_14640,N_5835,N_5687);
and U14641 (N_14641,N_8640,N_8945);
nor U14642 (N_14642,N_6321,N_7680);
or U14643 (N_14643,N_9523,N_7852);
nor U14644 (N_14644,N_5760,N_7057);
and U14645 (N_14645,N_8861,N_6591);
xor U14646 (N_14646,N_8950,N_6530);
nand U14647 (N_14647,N_7122,N_9536);
nor U14648 (N_14648,N_5302,N_5586);
nand U14649 (N_14649,N_5669,N_9058);
nor U14650 (N_14650,N_5797,N_7651);
and U14651 (N_14651,N_8148,N_9934);
nand U14652 (N_14652,N_9896,N_8725);
or U14653 (N_14653,N_5933,N_8595);
nand U14654 (N_14654,N_8805,N_5701);
or U14655 (N_14655,N_5644,N_7579);
or U14656 (N_14656,N_8223,N_8462);
and U14657 (N_14657,N_7840,N_9439);
nand U14658 (N_14658,N_6274,N_7286);
or U14659 (N_14659,N_8164,N_5244);
and U14660 (N_14660,N_8134,N_9268);
or U14661 (N_14661,N_7749,N_9276);
nand U14662 (N_14662,N_9959,N_7669);
nor U14663 (N_14663,N_5272,N_9768);
nor U14664 (N_14664,N_7943,N_6658);
nor U14665 (N_14665,N_9548,N_8318);
nand U14666 (N_14666,N_5586,N_9189);
nor U14667 (N_14667,N_9578,N_8714);
and U14668 (N_14668,N_9193,N_5855);
or U14669 (N_14669,N_9484,N_8547);
or U14670 (N_14670,N_7108,N_6348);
or U14671 (N_14671,N_7260,N_5346);
nand U14672 (N_14672,N_6781,N_8082);
and U14673 (N_14673,N_6064,N_6299);
and U14674 (N_14674,N_9994,N_9072);
and U14675 (N_14675,N_8330,N_6058);
nand U14676 (N_14676,N_5121,N_9537);
and U14677 (N_14677,N_6659,N_9313);
xnor U14678 (N_14678,N_5010,N_5911);
xor U14679 (N_14679,N_5963,N_9706);
nand U14680 (N_14680,N_7425,N_8225);
and U14681 (N_14681,N_7951,N_9829);
nand U14682 (N_14682,N_6324,N_9327);
xnor U14683 (N_14683,N_6837,N_6977);
nor U14684 (N_14684,N_6190,N_7048);
nand U14685 (N_14685,N_7384,N_7191);
xnor U14686 (N_14686,N_6433,N_5161);
and U14687 (N_14687,N_9586,N_9503);
nand U14688 (N_14688,N_6588,N_5620);
xnor U14689 (N_14689,N_9321,N_5728);
nor U14690 (N_14690,N_6361,N_8238);
nor U14691 (N_14691,N_9793,N_6875);
nand U14692 (N_14692,N_5013,N_6225);
nand U14693 (N_14693,N_6198,N_8049);
nor U14694 (N_14694,N_8005,N_9601);
nor U14695 (N_14695,N_9336,N_8737);
or U14696 (N_14696,N_5878,N_7216);
and U14697 (N_14697,N_6986,N_8026);
nor U14698 (N_14698,N_9380,N_6035);
and U14699 (N_14699,N_8610,N_6538);
nor U14700 (N_14700,N_8873,N_8391);
nand U14701 (N_14701,N_6221,N_8847);
or U14702 (N_14702,N_5070,N_7698);
or U14703 (N_14703,N_9675,N_7560);
xor U14704 (N_14704,N_8094,N_7138);
xor U14705 (N_14705,N_8846,N_9997);
nand U14706 (N_14706,N_9740,N_8681);
or U14707 (N_14707,N_8351,N_5587);
xnor U14708 (N_14708,N_7122,N_9638);
nor U14709 (N_14709,N_6027,N_8716);
nand U14710 (N_14710,N_9999,N_7855);
or U14711 (N_14711,N_8077,N_7401);
and U14712 (N_14712,N_7124,N_9628);
and U14713 (N_14713,N_6512,N_7630);
and U14714 (N_14714,N_6400,N_7547);
nand U14715 (N_14715,N_9782,N_6112);
nand U14716 (N_14716,N_7379,N_5207);
xor U14717 (N_14717,N_6420,N_6195);
and U14718 (N_14718,N_8414,N_6747);
or U14719 (N_14719,N_5877,N_7768);
nand U14720 (N_14720,N_8808,N_8501);
nand U14721 (N_14721,N_7085,N_9683);
nor U14722 (N_14722,N_8226,N_8596);
nor U14723 (N_14723,N_9791,N_6729);
nand U14724 (N_14724,N_7220,N_7516);
or U14725 (N_14725,N_8006,N_6303);
nand U14726 (N_14726,N_8004,N_7281);
nor U14727 (N_14727,N_5763,N_7697);
nor U14728 (N_14728,N_5995,N_8567);
and U14729 (N_14729,N_5619,N_7657);
nor U14730 (N_14730,N_5936,N_7056);
nand U14731 (N_14731,N_8453,N_9708);
xor U14732 (N_14732,N_7755,N_8054);
and U14733 (N_14733,N_5329,N_8593);
and U14734 (N_14734,N_5992,N_6081);
nor U14735 (N_14735,N_5576,N_6471);
nor U14736 (N_14736,N_6479,N_5795);
nand U14737 (N_14737,N_5142,N_6850);
nor U14738 (N_14738,N_7194,N_9160);
nor U14739 (N_14739,N_6491,N_9950);
nor U14740 (N_14740,N_8904,N_7968);
or U14741 (N_14741,N_7250,N_7903);
xnor U14742 (N_14742,N_9846,N_5251);
nand U14743 (N_14743,N_7689,N_8403);
or U14744 (N_14744,N_7988,N_8426);
xnor U14745 (N_14745,N_5476,N_9248);
or U14746 (N_14746,N_9568,N_9645);
nor U14747 (N_14747,N_8339,N_9689);
nor U14748 (N_14748,N_7499,N_7374);
and U14749 (N_14749,N_6896,N_7401);
nand U14750 (N_14750,N_6625,N_9501);
xor U14751 (N_14751,N_7536,N_9354);
xnor U14752 (N_14752,N_7215,N_5273);
and U14753 (N_14753,N_5529,N_9508);
and U14754 (N_14754,N_7879,N_5890);
nor U14755 (N_14755,N_8364,N_7169);
xnor U14756 (N_14756,N_6260,N_9843);
and U14757 (N_14757,N_9149,N_6095);
nor U14758 (N_14758,N_5503,N_9090);
nor U14759 (N_14759,N_7063,N_8076);
xor U14760 (N_14760,N_9975,N_6742);
nor U14761 (N_14761,N_9919,N_5669);
nor U14762 (N_14762,N_9923,N_9197);
nor U14763 (N_14763,N_7181,N_7577);
nand U14764 (N_14764,N_7801,N_8608);
nor U14765 (N_14765,N_6368,N_8878);
nor U14766 (N_14766,N_7237,N_7615);
and U14767 (N_14767,N_8376,N_5606);
nor U14768 (N_14768,N_8181,N_7954);
nand U14769 (N_14769,N_5540,N_9996);
nand U14770 (N_14770,N_9117,N_6339);
or U14771 (N_14771,N_7282,N_7946);
nand U14772 (N_14772,N_6506,N_7789);
or U14773 (N_14773,N_6977,N_7085);
nand U14774 (N_14774,N_5345,N_6394);
and U14775 (N_14775,N_8551,N_6809);
nand U14776 (N_14776,N_6456,N_7348);
or U14777 (N_14777,N_8694,N_8514);
and U14778 (N_14778,N_9326,N_8271);
or U14779 (N_14779,N_9114,N_9813);
nand U14780 (N_14780,N_9697,N_7354);
or U14781 (N_14781,N_9469,N_9637);
and U14782 (N_14782,N_6812,N_7224);
and U14783 (N_14783,N_5370,N_8828);
and U14784 (N_14784,N_6384,N_8819);
nand U14785 (N_14785,N_8304,N_7226);
nand U14786 (N_14786,N_5772,N_7405);
nand U14787 (N_14787,N_6501,N_7432);
and U14788 (N_14788,N_9404,N_5438);
nor U14789 (N_14789,N_8105,N_5088);
and U14790 (N_14790,N_5829,N_7372);
or U14791 (N_14791,N_8595,N_9648);
and U14792 (N_14792,N_9848,N_6713);
nand U14793 (N_14793,N_7366,N_7896);
or U14794 (N_14794,N_6851,N_7186);
nor U14795 (N_14795,N_6432,N_7710);
nor U14796 (N_14796,N_8743,N_8593);
nand U14797 (N_14797,N_5164,N_8052);
nand U14798 (N_14798,N_5142,N_6410);
or U14799 (N_14799,N_9882,N_6744);
or U14800 (N_14800,N_6262,N_7183);
nor U14801 (N_14801,N_8361,N_9777);
nor U14802 (N_14802,N_9854,N_5531);
nand U14803 (N_14803,N_7573,N_5390);
xor U14804 (N_14804,N_5011,N_9489);
nor U14805 (N_14805,N_7366,N_9667);
xor U14806 (N_14806,N_8541,N_5821);
nor U14807 (N_14807,N_8486,N_7040);
nand U14808 (N_14808,N_8295,N_5388);
nor U14809 (N_14809,N_8854,N_7330);
or U14810 (N_14810,N_8504,N_8313);
nand U14811 (N_14811,N_8854,N_8449);
and U14812 (N_14812,N_7357,N_5942);
or U14813 (N_14813,N_6346,N_8220);
nand U14814 (N_14814,N_7132,N_7241);
nand U14815 (N_14815,N_8984,N_8160);
nand U14816 (N_14816,N_5286,N_7605);
nor U14817 (N_14817,N_8752,N_7483);
or U14818 (N_14818,N_9870,N_7108);
nor U14819 (N_14819,N_5064,N_5426);
or U14820 (N_14820,N_8140,N_7074);
xor U14821 (N_14821,N_6753,N_8314);
and U14822 (N_14822,N_8184,N_8078);
and U14823 (N_14823,N_5307,N_7893);
xnor U14824 (N_14824,N_6562,N_8467);
or U14825 (N_14825,N_9553,N_7312);
nor U14826 (N_14826,N_8298,N_6671);
or U14827 (N_14827,N_6691,N_9060);
nand U14828 (N_14828,N_7218,N_6134);
xnor U14829 (N_14829,N_6554,N_6076);
and U14830 (N_14830,N_9127,N_8303);
or U14831 (N_14831,N_5981,N_8271);
and U14832 (N_14832,N_6878,N_6347);
or U14833 (N_14833,N_6630,N_8488);
or U14834 (N_14834,N_6208,N_8801);
and U14835 (N_14835,N_5525,N_6171);
nand U14836 (N_14836,N_8544,N_8287);
or U14837 (N_14837,N_6385,N_5157);
and U14838 (N_14838,N_7034,N_5516);
xor U14839 (N_14839,N_6339,N_8965);
nand U14840 (N_14840,N_6548,N_9935);
and U14841 (N_14841,N_7290,N_5319);
nor U14842 (N_14842,N_5272,N_9329);
and U14843 (N_14843,N_9294,N_5368);
xor U14844 (N_14844,N_9320,N_9359);
and U14845 (N_14845,N_7972,N_8943);
and U14846 (N_14846,N_5572,N_7055);
nand U14847 (N_14847,N_8078,N_6802);
nand U14848 (N_14848,N_9489,N_6770);
nor U14849 (N_14849,N_7544,N_5459);
nor U14850 (N_14850,N_6870,N_5931);
or U14851 (N_14851,N_9314,N_9204);
and U14852 (N_14852,N_6094,N_5520);
nor U14853 (N_14853,N_5132,N_6803);
nand U14854 (N_14854,N_8281,N_5565);
or U14855 (N_14855,N_5251,N_8321);
nor U14856 (N_14856,N_5136,N_8413);
and U14857 (N_14857,N_5903,N_7380);
or U14858 (N_14858,N_7266,N_6052);
xor U14859 (N_14859,N_6034,N_6245);
or U14860 (N_14860,N_5892,N_6542);
nand U14861 (N_14861,N_9345,N_9279);
xnor U14862 (N_14862,N_7099,N_9356);
nor U14863 (N_14863,N_6536,N_7318);
nand U14864 (N_14864,N_9298,N_6422);
nor U14865 (N_14865,N_9883,N_9386);
and U14866 (N_14866,N_6801,N_7369);
nor U14867 (N_14867,N_9430,N_8920);
nor U14868 (N_14868,N_8637,N_6617);
and U14869 (N_14869,N_7793,N_8193);
nand U14870 (N_14870,N_9182,N_5030);
nor U14871 (N_14871,N_9366,N_9266);
nand U14872 (N_14872,N_8985,N_9348);
xnor U14873 (N_14873,N_7635,N_8872);
and U14874 (N_14874,N_5108,N_8329);
nand U14875 (N_14875,N_7138,N_6078);
and U14876 (N_14876,N_9604,N_7595);
nor U14877 (N_14877,N_9883,N_8432);
xnor U14878 (N_14878,N_8026,N_9177);
and U14879 (N_14879,N_6567,N_6448);
and U14880 (N_14880,N_6040,N_7952);
nand U14881 (N_14881,N_9617,N_6257);
nand U14882 (N_14882,N_6841,N_5935);
or U14883 (N_14883,N_5567,N_5204);
and U14884 (N_14884,N_9827,N_9932);
nand U14885 (N_14885,N_5803,N_7054);
and U14886 (N_14886,N_6236,N_7027);
nor U14887 (N_14887,N_7208,N_7462);
and U14888 (N_14888,N_9780,N_5993);
xor U14889 (N_14889,N_7130,N_6993);
or U14890 (N_14890,N_7306,N_6910);
nand U14891 (N_14891,N_9938,N_9697);
and U14892 (N_14892,N_9637,N_9512);
nor U14893 (N_14893,N_6750,N_8357);
and U14894 (N_14894,N_5703,N_6250);
or U14895 (N_14895,N_9079,N_5828);
xnor U14896 (N_14896,N_5247,N_8380);
or U14897 (N_14897,N_6906,N_7513);
nor U14898 (N_14898,N_5072,N_9007);
nand U14899 (N_14899,N_7414,N_6711);
nor U14900 (N_14900,N_7894,N_7063);
and U14901 (N_14901,N_7742,N_8624);
nand U14902 (N_14902,N_9276,N_8174);
nor U14903 (N_14903,N_7759,N_7010);
nand U14904 (N_14904,N_7632,N_8677);
nor U14905 (N_14905,N_9147,N_7888);
nand U14906 (N_14906,N_7847,N_7313);
or U14907 (N_14907,N_9392,N_9967);
or U14908 (N_14908,N_8056,N_7839);
nor U14909 (N_14909,N_5841,N_8023);
nand U14910 (N_14910,N_8356,N_5538);
or U14911 (N_14911,N_7216,N_9075);
or U14912 (N_14912,N_9918,N_5687);
or U14913 (N_14913,N_7436,N_6629);
or U14914 (N_14914,N_9983,N_7958);
or U14915 (N_14915,N_7515,N_6644);
and U14916 (N_14916,N_5746,N_8190);
nor U14917 (N_14917,N_9348,N_8587);
nor U14918 (N_14918,N_6083,N_6312);
nand U14919 (N_14919,N_8170,N_7534);
and U14920 (N_14920,N_5359,N_8157);
and U14921 (N_14921,N_8386,N_9875);
and U14922 (N_14922,N_9418,N_7809);
and U14923 (N_14923,N_8944,N_8862);
nand U14924 (N_14924,N_8327,N_7042);
nor U14925 (N_14925,N_8016,N_8217);
nand U14926 (N_14926,N_5416,N_7313);
nand U14927 (N_14927,N_5346,N_6860);
xor U14928 (N_14928,N_5077,N_5121);
nand U14929 (N_14929,N_7717,N_9404);
nor U14930 (N_14930,N_6719,N_6369);
or U14931 (N_14931,N_6254,N_8715);
nand U14932 (N_14932,N_9301,N_6583);
and U14933 (N_14933,N_8079,N_5484);
nor U14934 (N_14934,N_5777,N_6174);
or U14935 (N_14935,N_9777,N_7156);
nand U14936 (N_14936,N_5115,N_7585);
nor U14937 (N_14937,N_7779,N_9387);
nor U14938 (N_14938,N_8982,N_5792);
or U14939 (N_14939,N_5563,N_6381);
nand U14940 (N_14940,N_9319,N_9661);
xnor U14941 (N_14941,N_8588,N_6040);
nand U14942 (N_14942,N_6500,N_9070);
xor U14943 (N_14943,N_6396,N_9119);
and U14944 (N_14944,N_7047,N_7969);
or U14945 (N_14945,N_5989,N_6527);
and U14946 (N_14946,N_7576,N_8735);
or U14947 (N_14947,N_7704,N_5156);
and U14948 (N_14948,N_9599,N_9538);
nor U14949 (N_14949,N_5448,N_5625);
and U14950 (N_14950,N_6070,N_7973);
nor U14951 (N_14951,N_7275,N_9347);
or U14952 (N_14952,N_7531,N_5191);
nand U14953 (N_14953,N_9469,N_7892);
or U14954 (N_14954,N_5363,N_6551);
or U14955 (N_14955,N_7968,N_9875);
nor U14956 (N_14956,N_9417,N_7373);
nor U14957 (N_14957,N_8728,N_7077);
or U14958 (N_14958,N_6244,N_6487);
or U14959 (N_14959,N_5689,N_5952);
nand U14960 (N_14960,N_9251,N_8066);
nand U14961 (N_14961,N_7734,N_7992);
nor U14962 (N_14962,N_6119,N_5585);
or U14963 (N_14963,N_7530,N_9061);
and U14964 (N_14964,N_6333,N_7047);
and U14965 (N_14965,N_8832,N_8611);
nand U14966 (N_14966,N_6822,N_8347);
nand U14967 (N_14967,N_9062,N_9778);
nand U14968 (N_14968,N_6664,N_9076);
xor U14969 (N_14969,N_7632,N_5950);
and U14970 (N_14970,N_8847,N_8862);
or U14971 (N_14971,N_6097,N_6336);
or U14972 (N_14972,N_6343,N_8984);
nand U14973 (N_14973,N_9658,N_7220);
or U14974 (N_14974,N_7172,N_8858);
nor U14975 (N_14975,N_6054,N_8627);
and U14976 (N_14976,N_9731,N_8227);
xor U14977 (N_14977,N_8739,N_7576);
and U14978 (N_14978,N_7187,N_8814);
or U14979 (N_14979,N_8806,N_8649);
nor U14980 (N_14980,N_6217,N_7570);
or U14981 (N_14981,N_7780,N_5778);
and U14982 (N_14982,N_6257,N_7234);
nand U14983 (N_14983,N_7686,N_7730);
and U14984 (N_14984,N_8077,N_9529);
and U14985 (N_14985,N_8467,N_7975);
nand U14986 (N_14986,N_6066,N_5375);
and U14987 (N_14987,N_7163,N_6456);
xor U14988 (N_14988,N_8030,N_8669);
nand U14989 (N_14989,N_7103,N_6393);
and U14990 (N_14990,N_6846,N_5178);
nor U14991 (N_14991,N_9503,N_8091);
nand U14992 (N_14992,N_8435,N_9745);
nor U14993 (N_14993,N_5373,N_6720);
or U14994 (N_14994,N_7582,N_6080);
and U14995 (N_14995,N_9462,N_7204);
and U14996 (N_14996,N_6838,N_7022);
and U14997 (N_14997,N_5879,N_9340);
nor U14998 (N_14998,N_8594,N_6309);
xnor U14999 (N_14999,N_9623,N_5231);
and U15000 (N_15000,N_11056,N_10086);
nor U15001 (N_15001,N_10821,N_10192);
nor U15002 (N_15002,N_10724,N_12704);
nand U15003 (N_15003,N_14532,N_10820);
xnor U15004 (N_15004,N_13425,N_10713);
nor U15005 (N_15005,N_13535,N_11923);
and U15006 (N_15006,N_14880,N_14794);
xor U15007 (N_15007,N_10774,N_12682);
and U15008 (N_15008,N_11769,N_11410);
nor U15009 (N_15009,N_12264,N_13924);
nand U15010 (N_15010,N_11831,N_10340);
or U15011 (N_15011,N_10139,N_14965);
nand U15012 (N_15012,N_10293,N_13163);
and U15013 (N_15013,N_13172,N_10051);
and U15014 (N_15014,N_10624,N_12064);
nand U15015 (N_15015,N_14859,N_10960);
xnor U15016 (N_15016,N_11797,N_10399);
or U15017 (N_15017,N_12427,N_11468);
or U15018 (N_15018,N_12449,N_13318);
nand U15019 (N_15019,N_11428,N_10559);
and U15020 (N_15020,N_11272,N_12987);
and U15021 (N_15021,N_14864,N_13586);
nand U15022 (N_15022,N_11949,N_13148);
or U15023 (N_15023,N_12342,N_14256);
and U15024 (N_15024,N_11160,N_10799);
nor U15025 (N_15025,N_13480,N_13330);
xnor U15026 (N_15026,N_13164,N_12839);
nand U15027 (N_15027,N_14206,N_11125);
or U15028 (N_15028,N_12691,N_12376);
and U15029 (N_15029,N_12948,N_14637);
or U15030 (N_15030,N_12412,N_12758);
and U15031 (N_15031,N_13388,N_10899);
and U15032 (N_15032,N_13717,N_10346);
or U15033 (N_15033,N_10874,N_11389);
and U15034 (N_15034,N_12310,N_14442);
or U15035 (N_15035,N_14839,N_11047);
nor U15036 (N_15036,N_13596,N_13809);
and U15037 (N_15037,N_13760,N_14979);
and U15038 (N_15038,N_10123,N_14426);
or U15039 (N_15039,N_14621,N_11441);
nand U15040 (N_15040,N_12651,N_10499);
xor U15041 (N_15041,N_13531,N_10373);
and U15042 (N_15042,N_10913,N_13006);
and U15043 (N_15043,N_13750,N_12582);
and U15044 (N_15044,N_10442,N_10418);
and U15045 (N_15045,N_14680,N_14054);
and U15046 (N_15046,N_13368,N_12361);
xor U15047 (N_15047,N_11878,N_14754);
or U15048 (N_15048,N_12295,N_13153);
and U15049 (N_15049,N_12410,N_12785);
nor U15050 (N_15050,N_10538,N_14057);
nand U15051 (N_15051,N_13915,N_12181);
nand U15052 (N_15052,N_11988,N_13861);
and U15053 (N_15053,N_13260,N_13081);
nand U15054 (N_15054,N_14362,N_13695);
nor U15055 (N_15055,N_12793,N_11522);
and U15056 (N_15056,N_11446,N_11614);
or U15057 (N_15057,N_13245,N_12846);
nand U15058 (N_15058,N_10746,N_13617);
or U15059 (N_15059,N_13642,N_11978);
nor U15060 (N_15060,N_13461,N_10444);
or U15061 (N_15061,N_13649,N_11263);
nor U15062 (N_15062,N_10431,N_10602);
or U15063 (N_15063,N_14263,N_10840);
or U15064 (N_15064,N_14853,N_14141);
nand U15065 (N_15065,N_12159,N_11147);
nand U15066 (N_15066,N_12912,N_11938);
nand U15067 (N_15067,N_10247,N_13893);
and U15068 (N_15068,N_12465,N_14540);
nor U15069 (N_15069,N_14456,N_12848);
nand U15070 (N_15070,N_11653,N_10339);
xnor U15071 (N_15071,N_10817,N_10710);
nand U15072 (N_15072,N_14874,N_10416);
nor U15073 (N_15073,N_10756,N_12850);
or U15074 (N_15074,N_12239,N_11453);
nor U15075 (N_15075,N_11411,N_14541);
nand U15076 (N_15076,N_10895,N_10187);
or U15077 (N_15077,N_12219,N_12795);
nor U15078 (N_15078,N_13161,N_12707);
nand U15079 (N_15079,N_10352,N_12393);
nand U15080 (N_15080,N_11423,N_14297);
nand U15081 (N_15081,N_14714,N_10301);
or U15082 (N_15082,N_12730,N_12595);
nor U15083 (N_15083,N_11964,N_13204);
nor U15084 (N_15084,N_12455,N_14108);
nor U15085 (N_15085,N_13061,N_12089);
and U15086 (N_15086,N_13125,N_12590);
or U15087 (N_15087,N_12214,N_10787);
nor U15088 (N_15088,N_12605,N_12103);
and U15089 (N_15089,N_11102,N_10269);
nor U15090 (N_15090,N_12355,N_13625);
or U15091 (N_15091,N_10026,N_13860);
and U15092 (N_15092,N_11060,N_11252);
and U15093 (N_15093,N_10833,N_12714);
and U15094 (N_15094,N_11073,N_11178);
nand U15095 (N_15095,N_11776,N_11870);
and U15096 (N_15096,N_13342,N_10462);
and U15097 (N_15097,N_12451,N_11151);
and U15098 (N_15098,N_13254,N_10590);
nand U15099 (N_15099,N_14867,N_14342);
or U15100 (N_15100,N_10395,N_14967);
nand U15101 (N_15101,N_11229,N_13089);
and U15102 (N_15102,N_12083,N_13333);
xor U15103 (N_15103,N_12504,N_12399);
and U15104 (N_15104,N_10775,N_13424);
xnor U15105 (N_15105,N_13097,N_13775);
or U15106 (N_15106,N_12980,N_13358);
and U15107 (N_15107,N_13228,N_13540);
nand U15108 (N_15108,N_12529,N_11126);
nand U15109 (N_15109,N_12278,N_14418);
or U15110 (N_15110,N_13834,N_14516);
xnor U15111 (N_15111,N_14352,N_10581);
or U15112 (N_15112,N_13502,N_12729);
and U15113 (N_15113,N_14630,N_12289);
nor U15114 (N_15114,N_10630,N_14310);
nor U15115 (N_15115,N_11367,N_13199);
and U15116 (N_15116,N_12421,N_14575);
nand U15117 (N_15117,N_12930,N_13721);
and U15118 (N_15118,N_12681,N_10058);
or U15119 (N_15119,N_10188,N_14333);
and U15120 (N_15120,N_13194,N_14629);
and U15121 (N_15121,N_13665,N_12223);
nor U15122 (N_15122,N_14649,N_10118);
and U15123 (N_15123,N_13601,N_13562);
nand U15124 (N_15124,N_14851,N_13146);
or U15125 (N_15125,N_12302,N_11068);
and U15126 (N_15126,N_14339,N_14353);
nand U15127 (N_15127,N_12572,N_10532);
nor U15128 (N_15128,N_11015,N_10699);
nor U15129 (N_15129,N_14747,N_11471);
or U15130 (N_15130,N_10831,N_13899);
or U15131 (N_15131,N_13115,N_12260);
and U15132 (N_15132,N_12722,N_12810);
nand U15133 (N_15133,N_14015,N_14602);
nor U15134 (N_15134,N_14586,N_10777);
or U15135 (N_15135,N_11830,N_12836);
nor U15136 (N_15136,N_10966,N_11117);
or U15137 (N_15137,N_12438,N_13436);
and U15138 (N_15138,N_12230,N_12804);
and U15139 (N_15139,N_13881,N_13229);
and U15140 (N_15140,N_14778,N_10637);
nand U15141 (N_15141,N_12929,N_10007);
or U15142 (N_15142,N_12444,N_11319);
nor U15143 (N_15143,N_11707,N_12114);
nand U15144 (N_15144,N_10082,N_10550);
nand U15145 (N_15145,N_10447,N_10337);
nor U15146 (N_15146,N_14706,N_14550);
nand U15147 (N_15147,N_13746,N_13608);
nor U15148 (N_15148,N_10101,N_14274);
and U15149 (N_15149,N_13565,N_10470);
or U15150 (N_15150,N_10837,N_12338);
and U15151 (N_15151,N_10454,N_14017);
or U15152 (N_15152,N_11381,N_13890);
nor U15153 (N_15153,N_12872,N_14528);
nor U15154 (N_15154,N_13396,N_11975);
nor U15155 (N_15155,N_12300,N_13246);
nand U15156 (N_15156,N_13747,N_14407);
and U15157 (N_15157,N_13118,N_14158);
and U15158 (N_15158,N_13434,N_10978);
nand U15159 (N_15159,N_11496,N_13181);
nand U15160 (N_15160,N_14558,N_13488);
nand U15161 (N_15161,N_13714,N_12461);
nand U15162 (N_15162,N_14623,N_14952);
xor U15163 (N_15163,N_11418,N_13037);
nand U15164 (N_15164,N_10389,N_14598);
and U15165 (N_15165,N_11583,N_10805);
nand U15166 (N_15166,N_11974,N_14397);
and U15167 (N_15167,N_11741,N_12928);
or U15168 (N_15168,N_14029,N_10653);
nor U15169 (N_15169,N_13939,N_13764);
and U15170 (N_15170,N_13969,N_13043);
and U15171 (N_15171,N_13618,N_12238);
nand U15172 (N_15172,N_11188,N_10488);
nor U15173 (N_15173,N_13628,N_11668);
nand U15174 (N_15174,N_12979,N_12389);
nand U15175 (N_15175,N_12241,N_14555);
nand U15176 (N_15176,N_10062,N_11807);
or U15177 (N_15177,N_13459,N_14448);
or U15178 (N_15178,N_11451,N_11306);
and U15179 (N_15179,N_13472,N_12063);
and U15180 (N_15180,N_14172,N_12129);
and U15181 (N_15181,N_14363,N_13614);
nand U15182 (N_15182,N_10839,N_12431);
or U15183 (N_15183,N_11597,N_13162);
nor U15184 (N_15184,N_10260,N_12225);
or U15185 (N_15185,N_11713,N_10726);
and U15186 (N_15186,N_14543,N_12915);
and U15187 (N_15187,N_10209,N_14790);
or U15188 (N_15188,N_13453,N_10492);
nor U15189 (N_15189,N_11899,N_11641);
nand U15190 (N_15190,N_13394,N_13656);
nor U15191 (N_15191,N_12816,N_13356);
nor U15192 (N_15192,N_11017,N_12373);
nor U15193 (N_15193,N_14007,N_12145);
and U15194 (N_15194,N_12788,N_12511);
nor U15195 (N_15195,N_14214,N_14679);
nor U15196 (N_15196,N_13561,N_12261);
xor U15197 (N_15197,N_10019,N_13982);
nand U15198 (N_15198,N_11763,N_11898);
xnor U15199 (N_15199,N_13730,N_12951);
nor U15200 (N_15200,N_11693,N_13401);
nand U15201 (N_15201,N_14593,N_11874);
or U15202 (N_15202,N_13180,N_11655);
nand U15203 (N_15203,N_14611,N_11348);
xnor U15204 (N_15204,N_14815,N_14404);
xor U15205 (N_15205,N_10725,N_13839);
or U15206 (N_15206,N_11876,N_14673);
and U15207 (N_15207,N_12500,N_13639);
and U15208 (N_15208,N_14531,N_11563);
or U15209 (N_15209,N_10932,N_14931);
or U15210 (N_15210,N_11589,N_12404);
nand U15211 (N_15211,N_13406,N_12820);
nand U15212 (N_15212,N_11948,N_14951);
nand U15213 (N_15213,N_11499,N_14733);
nor U15214 (N_15214,N_10789,N_10834);
and U15215 (N_15215,N_12199,N_11591);
nand U15216 (N_15216,N_12234,N_14605);
nand U15217 (N_15217,N_11619,N_10614);
nor U15218 (N_15218,N_12318,N_14379);
and U15219 (N_15219,N_11219,N_11660);
nand U15220 (N_15220,N_11193,N_14934);
nor U15221 (N_15221,N_14551,N_12555);
and U15222 (N_15222,N_13175,N_12016);
nand U15223 (N_15223,N_12828,N_13984);
nand U15224 (N_15224,N_14897,N_12075);
nor U15225 (N_15225,N_11625,N_11085);
nor U15226 (N_15226,N_11986,N_13374);
xnor U15227 (N_15227,N_12168,N_11430);
nor U15228 (N_15228,N_14529,N_12903);
nand U15229 (N_15229,N_12700,N_12434);
nor U15230 (N_15230,N_10857,N_12853);
or U15231 (N_15231,N_11454,N_11347);
nor U15232 (N_15232,N_12787,N_10309);
and U15233 (N_15233,N_13923,N_11857);
nor U15234 (N_15234,N_10105,N_11516);
or U15235 (N_15235,N_11795,N_12067);
xor U15236 (N_15236,N_14085,N_13227);
and U15237 (N_15237,N_13567,N_12210);
nand U15238 (N_15238,N_10999,N_12695);
nand U15239 (N_15239,N_13776,N_13782);
nor U15240 (N_15240,N_11042,N_14400);
nor U15241 (N_15241,N_11561,N_10753);
and U15242 (N_15242,N_13636,N_12671);
and U15243 (N_15243,N_12172,N_14721);
or U15244 (N_15244,N_11279,N_14760);
nor U15245 (N_15245,N_14222,N_11156);
and U15246 (N_15246,N_10589,N_13708);
nor U15247 (N_15247,N_11202,N_14360);
nand U15248 (N_15248,N_10421,N_10283);
xnor U15249 (N_15249,N_12965,N_13967);
or U15250 (N_15250,N_13755,N_10679);
or U15251 (N_15251,N_13250,N_13367);
and U15252 (N_15252,N_12432,N_12661);
nand U15253 (N_15253,N_11264,N_12437);
nand U15254 (N_15254,N_10945,N_13483);
nand U15255 (N_15255,N_14512,N_12933);
or U15256 (N_15256,N_13432,N_14066);
xnor U15257 (N_15257,N_12101,N_14654);
nand U15258 (N_15258,N_13258,N_14018);
and U15259 (N_15259,N_11150,N_12311);
nand U15260 (N_15260,N_10328,N_13290);
or U15261 (N_15261,N_12287,N_14204);
and U15262 (N_15262,N_11881,N_12351);
nand U15263 (N_15263,N_12745,N_11520);
xnor U15264 (N_15264,N_14786,N_13210);
and U15265 (N_15265,N_11474,N_11703);
or U15266 (N_15266,N_12498,N_14046);
nor U15267 (N_15267,N_11897,N_12255);
nand U15268 (N_15268,N_12509,N_11664);
xnor U15269 (N_15269,N_11801,N_11325);
nand U15270 (N_15270,N_10803,N_14603);
or U15271 (N_15271,N_13187,N_11826);
and U15272 (N_15272,N_13159,N_13033);
or U15273 (N_15273,N_11054,N_10755);
or U15274 (N_15274,N_14735,N_10429);
nand U15275 (N_15275,N_12122,N_10665);
and U15276 (N_15276,N_10361,N_12782);
nand U15277 (N_15277,N_14601,N_10060);
and U15278 (N_15278,N_10298,N_11271);
nor U15279 (N_15279,N_10354,N_10394);
nand U15280 (N_15280,N_10253,N_10696);
and U15281 (N_15281,N_13214,N_13291);
or U15282 (N_15282,N_10863,N_13121);
and U15283 (N_15283,N_12345,N_11526);
nor U15284 (N_15284,N_10761,N_14296);
nor U15285 (N_15285,N_14704,N_13598);
nor U15286 (N_15286,N_10584,N_12962);
nor U15287 (N_15287,N_13169,N_11359);
nor U15288 (N_15288,N_11911,N_13316);
or U15289 (N_15289,N_13666,N_13901);
nand U15290 (N_15290,N_14064,N_12008);
nor U15291 (N_15291,N_14372,N_11571);
and U15292 (N_15292,N_13897,N_14179);
nor U15293 (N_15293,N_10272,N_14272);
or U15294 (N_15294,N_11352,N_14135);
and U15295 (N_15295,N_12764,N_12581);
nand U15296 (N_15296,N_11221,N_10648);
nand U15297 (N_15297,N_11701,N_10281);
nor U15298 (N_15298,N_11793,N_10248);
and U15299 (N_15299,N_14666,N_11575);
nand U15300 (N_15300,N_11939,N_13437);
xor U15301 (N_15301,N_14774,N_12053);
xnor U15302 (N_15302,N_12146,N_14133);
and U15303 (N_15303,N_13541,N_10300);
or U15304 (N_15304,N_11895,N_10475);
nand U15305 (N_15305,N_12017,N_13377);
and U15306 (N_15306,N_10263,N_12685);
nor U15307 (N_15307,N_10701,N_13945);
nor U15308 (N_15308,N_14412,N_11558);
nor U15309 (N_15309,N_10638,N_13551);
nand U15310 (N_15310,N_11260,N_10672);
or U15311 (N_15311,N_14993,N_13257);
nand U15312 (N_15312,N_13460,N_14663);
and U15313 (N_15313,N_11323,N_14176);
nand U15314 (N_15314,N_13744,N_14288);
nor U15315 (N_15315,N_11327,N_14768);
or U15316 (N_15316,N_12130,N_11786);
nand U15317 (N_15317,N_11514,N_12157);
and U15318 (N_15318,N_10912,N_14157);
nand U15319 (N_15319,N_13218,N_14161);
or U15320 (N_15320,N_11353,N_10374);
or U15321 (N_15321,N_10930,N_13676);
or U15322 (N_15322,N_10592,N_14217);
nor U15323 (N_15323,N_11691,N_11543);
nand U15324 (N_15324,N_12392,N_14321);
nand U15325 (N_15325,N_12835,N_12840);
nand U15326 (N_15326,N_12757,N_10632);
nor U15327 (N_15327,N_14315,N_14656);
and U15328 (N_15328,N_10734,N_13397);
or U15329 (N_15329,N_14683,N_12815);
nor U15330 (N_15330,N_10419,N_13857);
and U15331 (N_15331,N_13120,N_14398);
and U15332 (N_15332,N_10798,N_12766);
xor U15333 (N_15333,N_14749,N_12003);
nand U15334 (N_15334,N_13289,N_12119);
nor U15335 (N_15335,N_14618,N_14791);
xor U15336 (N_15336,N_12280,N_10237);
nor U15337 (N_15337,N_13520,N_14112);
nor U15338 (N_15338,N_11431,N_10703);
nand U15339 (N_15339,N_14963,N_10401);
nand U15340 (N_15340,N_14487,N_12070);
xnor U15341 (N_15341,N_11405,N_10560);
nor U15342 (N_15342,N_10748,N_12823);
nor U15343 (N_15343,N_10047,N_12608);
nand U15344 (N_15344,N_14651,N_10119);
and U15345 (N_15345,N_14997,N_13211);
and U15346 (N_15346,N_13837,N_12967);
nor U15347 (N_15347,N_11070,N_12881);
nand U15348 (N_15348,N_11022,N_10243);
nand U15349 (N_15349,N_13370,N_14813);
or U15350 (N_15350,N_13631,N_14533);
xnor U15351 (N_15351,N_13481,N_13408);
or U15352 (N_15352,N_12161,N_12802);
and U15353 (N_15353,N_12252,N_12811);
xor U15354 (N_15354,N_11618,N_11754);
nand U15355 (N_15355,N_14882,N_11984);
nand U15356 (N_15356,N_11510,N_10513);
nand U15357 (N_15357,N_12167,N_11623);
nand U15358 (N_15358,N_11243,N_11690);
and U15359 (N_15359,N_13655,N_12880);
xnor U15360 (N_15360,N_11290,N_14798);
or U15361 (N_15361,N_13126,N_12014);
and U15362 (N_15362,N_10076,N_10125);
nand U15363 (N_15363,N_13793,N_11209);
or U15364 (N_15364,N_10471,N_10052);
or U15365 (N_15365,N_11654,N_14773);
and U15366 (N_15366,N_11470,N_13849);
xor U15367 (N_15367,N_13362,N_13339);
or U15368 (N_15368,N_13278,N_11906);
nor U15369 (N_15369,N_14674,N_13093);
nor U15370 (N_15370,N_11953,N_12152);
xor U15371 (N_15371,N_10733,N_12303);
or U15372 (N_15372,N_13456,N_11889);
nor U15373 (N_15373,N_10830,N_12968);
or U15374 (N_15374,N_11377,N_10962);
nand U15375 (N_15375,N_14136,N_14676);
or U15376 (N_15376,N_12870,N_14062);
nand U15377 (N_15377,N_13363,N_12673);
and U15378 (N_15378,N_13039,N_12217);
nor U15379 (N_15379,N_10644,N_12622);
nor U15380 (N_15380,N_10934,N_12143);
nand U15381 (N_15381,N_11071,N_11186);
nand U15382 (N_15382,N_10654,N_13584);
nand U15383 (N_15383,N_11685,N_12142);
nor U15384 (N_15384,N_12803,N_12046);
nor U15385 (N_15385,N_13983,N_12742);
nor U15386 (N_15386,N_10577,N_12667);
xnor U15387 (N_15387,N_11120,N_10880);
xnor U15388 (N_15388,N_10866,N_13390);
and U15389 (N_15389,N_11662,N_10812);
xor U15390 (N_15390,N_11236,N_10832);
nor U15391 (N_15391,N_11111,N_14509);
xor U15392 (N_15392,N_13335,N_10404);
or U15393 (N_15393,N_13269,N_10197);
and U15394 (N_15394,N_11832,N_11128);
nor U15395 (N_15395,N_10497,N_13938);
nor U15396 (N_15396,N_12925,N_14409);
and U15397 (N_15397,N_13088,N_13878);
or U15398 (N_15398,N_14995,N_12777);
nor U15399 (N_15399,N_14235,N_11745);
and U15400 (N_15400,N_13225,N_10519);
nand U15401 (N_15401,N_10040,N_11427);
nand U15402 (N_15402,N_10091,N_14285);
nor U15403 (N_15403,N_14739,N_11827);
or U15404 (N_15404,N_10074,N_10064);
xnor U15405 (N_15405,N_11821,N_14961);
and U15406 (N_15406,N_14131,N_11309);
and U15407 (N_15407,N_10694,N_11240);
and U15408 (N_15408,N_13936,N_10531);
nor U15409 (N_15409,N_14819,N_11731);
nand U15410 (N_15410,N_14536,N_11237);
nand U15411 (N_15411,N_12614,N_11550);
xor U15412 (N_15412,N_14828,N_11094);
or U15413 (N_15413,N_14566,N_10333);
or U15414 (N_15414,N_13987,N_11066);
or U15415 (N_15415,N_11037,N_11581);
and U15416 (N_15416,N_12076,N_14642);
nand U15417 (N_15417,N_14872,N_10341);
or U15418 (N_15418,N_13384,N_12124);
and U15419 (N_15419,N_13560,N_11785);
and U15420 (N_15420,N_10533,N_12821);
or U15421 (N_15421,N_10901,N_14795);
and U15422 (N_15422,N_13413,N_11644);
nand U15423 (N_15423,N_12702,N_11772);
nand U15424 (N_15424,N_11917,N_14344);
nand U15425 (N_15425,N_10898,N_12290);
and U15426 (N_15426,N_10740,N_11838);
or U15427 (N_15427,N_13308,N_12944);
xnor U15428 (N_15428,N_14019,N_14380);
or U15429 (N_15429,N_13004,N_12643);
and U15430 (N_15430,N_13787,N_13497);
and U15431 (N_15431,N_11314,N_13610);
and U15432 (N_15432,N_12994,N_13554);
nor U15433 (N_15433,N_11124,N_13034);
and U15434 (N_15434,N_13659,N_14051);
or U15435 (N_15435,N_10811,N_13765);
nand U15436 (N_15436,N_14767,N_10195);
or U15437 (N_15437,N_14446,N_14667);
nor U15438 (N_15438,N_10687,N_13174);
nand U15439 (N_15439,N_14443,N_12905);
nand U15440 (N_15440,N_10525,N_14099);
or U15441 (N_15441,N_10224,N_12890);
xnor U15442 (N_15442,N_13455,N_14591);
nor U15443 (N_15443,N_14451,N_13563);
or U15444 (N_15444,N_10652,N_14696);
nand U15445 (N_15445,N_11517,N_10478);
nor U15446 (N_15446,N_12327,N_14012);
nand U15447 (N_15447,N_14336,N_10769);
nand U15448 (N_15448,N_11119,N_11940);
nor U15449 (N_15449,N_13421,N_12633);
nand U15450 (N_15450,N_13253,N_10793);
nor U15451 (N_15451,N_14474,N_10356);
or U15452 (N_15452,N_13013,N_14570);
and U15453 (N_15453,N_11629,N_14369);
or U15454 (N_15454,N_12060,N_12332);
nor U15455 (N_15455,N_10287,N_14781);
nand U15456 (N_15456,N_11959,N_11224);
nor U15457 (N_15457,N_12380,N_10244);
nand U15458 (N_15458,N_13789,N_10069);
and U15459 (N_15459,N_11732,N_13556);
and U15460 (N_15460,N_12319,N_13552);
and U15461 (N_15461,N_13819,N_12298);
and U15462 (N_15462,N_12619,N_13446);
and U15463 (N_15463,N_13828,N_13769);
nor U15464 (N_15464,N_12022,N_13680);
and U15465 (N_15465,N_11254,N_13763);
or U15466 (N_15466,N_13411,N_14868);
nand U15467 (N_15467,N_13949,N_14756);
or U15468 (N_15468,N_13926,N_14914);
and U15469 (N_15469,N_12462,N_12895);
or U15470 (N_15470,N_14985,N_14037);
nor U15471 (N_15471,N_11605,N_11481);
nand U15472 (N_15472,N_14144,N_13021);
and U15473 (N_15473,N_14025,N_14527);
and U15474 (N_15474,N_12062,N_11683);
nand U15475 (N_15475,N_10473,N_12522);
nor U15476 (N_15476,N_11201,N_12094);
or U15477 (N_15477,N_14232,N_12160);
nand U15478 (N_15478,N_13219,N_13539);
or U15479 (N_15479,N_11168,N_10662);
nand U15480 (N_15480,N_12254,N_10169);
nor U15481 (N_15481,N_12448,N_14660);
and U15482 (N_15482,N_13448,N_12937);
or U15483 (N_15483,N_14160,N_12317);
or U15484 (N_15484,N_11256,N_13854);
or U15485 (N_15485,N_10810,N_14127);
and U15486 (N_15486,N_14361,N_11528);
and U15487 (N_15487,N_11375,N_12958);
or U15488 (N_15488,N_12887,N_12824);
nor U15489 (N_15489,N_14081,N_14137);
or U15490 (N_15490,N_10896,N_10693);
and U15491 (N_15491,N_12452,N_13048);
nor U15492 (N_15492,N_14027,N_12192);
or U15493 (N_15493,N_14999,N_14300);
nand U15494 (N_15494,N_10582,N_10961);
nor U15495 (N_15495,N_10109,N_11602);
nand U15496 (N_15496,N_12780,N_10970);
nor U15497 (N_15497,N_10189,N_14248);
nand U15498 (N_15498,N_12519,N_14640);
nor U15499 (N_15499,N_13732,N_11445);
or U15500 (N_15500,N_12270,N_10144);
nand U15501 (N_15501,N_12125,N_10965);
nand U15502 (N_15502,N_12855,N_10623);
nor U15503 (N_15503,N_12574,N_13122);
and U15504 (N_15504,N_14173,N_11737);
nand U15505 (N_15505,N_13802,N_10828);
nand U15506 (N_15506,N_14292,N_11565);
nand U15507 (N_15507,N_10979,N_12218);
nand U15508 (N_15508,N_10572,N_11513);
and U15509 (N_15509,N_10749,N_14061);
xnor U15510 (N_15510,N_13993,N_12735);
nor U15511 (N_15511,N_10975,N_14472);
xnor U15512 (N_15512,N_11058,N_11574);
nor U15513 (N_15513,N_12592,N_13671);
nand U15514 (N_15514,N_10255,N_11244);
nor U15515 (N_15515,N_14940,N_13311);
or U15516 (N_15516,N_12057,N_10093);
nand U15517 (N_15517,N_14782,N_13478);
nor U15518 (N_15518,N_14935,N_13998);
and U15519 (N_15519,N_14772,N_10607);
and U15520 (N_15520,N_14276,N_11392);
and U15521 (N_15521,N_11304,N_13593);
nand U15522 (N_15522,N_10305,N_14659);
xnor U15523 (N_15523,N_12760,N_14335);
nand U15524 (N_15524,N_14251,N_12275);
or U15525 (N_15525,N_11131,N_10849);
nand U15526 (N_15526,N_10294,N_14910);
or U15527 (N_15527,N_11180,N_10332);
nand U15528 (N_15528,N_13831,N_13473);
or U15529 (N_15529,N_14757,N_10306);
and U15530 (N_15530,N_14326,N_10608);
xor U15531 (N_15531,N_12236,N_11726);
and U15532 (N_15532,N_12868,N_11553);
or U15533 (N_15533,N_13001,N_13104);
and U15534 (N_15534,N_14294,N_11950);
xnor U15535 (N_15535,N_10203,N_10172);
nor U15536 (N_15536,N_13637,N_11919);
nor U15537 (N_15537,N_10311,N_10396);
nor U15538 (N_15538,N_13806,N_11845);
nor U15539 (N_15539,N_11095,N_10682);
or U15540 (N_15540,N_12085,N_11719);
nor U15541 (N_15541,N_14567,N_11485);
and U15542 (N_15542,N_13866,N_13025);
nand U15543 (N_15543,N_10986,N_14716);
or U15544 (N_15544,N_12208,N_13489);
xor U15545 (N_15545,N_12069,N_12784);
or U15546 (N_15546,N_14445,N_12752);
or U15547 (N_15547,N_13018,N_14182);
or U15548 (N_15548,N_12321,N_11721);
and U15549 (N_15549,N_10122,N_10021);
nand U15550 (N_15550,N_10166,N_10995);
and U15551 (N_15551,N_13203,N_11157);
or U15552 (N_15552,N_11920,N_13885);
nor U15553 (N_15553,N_11735,N_11868);
and U15554 (N_15554,N_10633,N_14959);
nor U15555 (N_15555,N_12978,N_14408);
nor U15556 (N_15556,N_10070,N_14895);
nand U15557 (N_15557,N_11842,N_10884);
and U15558 (N_15558,N_13921,N_12144);
or U15559 (N_15559,N_11135,N_13643);
nor U15560 (N_15560,N_14489,N_11996);
or U15561 (N_15561,N_10664,N_11649);
nor U15562 (N_15562,N_14134,N_12954);
nor U15563 (N_15563,N_11502,N_12276);
nor U15564 (N_15564,N_10292,N_10050);
xnor U15565 (N_15565,N_11971,N_11005);
nor U15566 (N_15566,N_12762,N_13049);
nor U15567 (N_15567,N_12718,N_14032);
nor U15568 (N_15568,N_10905,N_11551);
nor U15569 (N_15569,N_13108,N_11738);
xor U15570 (N_15570,N_14941,N_14105);
nor U15571 (N_15571,N_14507,N_14322);
and U15572 (N_15572,N_10391,N_11455);
and U15573 (N_15573,N_11001,N_13826);
or U15574 (N_15574,N_13297,N_10184);
xnor U15575 (N_15575,N_11839,N_11572);
or U15576 (N_15576,N_12191,N_14147);
nand U15577 (N_15577,N_12242,N_10134);
nor U15578 (N_15578,N_11190,N_12382);
nor U15579 (N_15579,N_10730,N_14191);
nand U15580 (N_15580,N_10400,N_13964);
nand U15581 (N_15581,N_10372,N_10520);
nor U15582 (N_15582,N_12961,N_11512);
nand U15583 (N_15583,N_14193,N_11074);
or U15584 (N_15584,N_13575,N_10336);
nor U15585 (N_15585,N_13963,N_10879);
and U15586 (N_15586,N_12805,N_12832);
nand U15587 (N_15587,N_12381,N_12406);
and U15588 (N_15588,N_10277,N_11130);
and U15589 (N_15589,N_13726,N_10526);
nor U15590 (N_15590,N_10618,N_14075);
nand U15591 (N_15591,N_14930,N_14228);
or U15592 (N_15592,N_12484,N_12982);
nor U15593 (N_15593,N_10032,N_13380);
nand U15594 (N_15594,N_10090,N_12458);
and U15595 (N_15595,N_14269,N_13249);
nor U15596 (N_15596,N_11215,N_10474);
nand U15597 (N_15597,N_13046,N_14022);
nand U15598 (N_15598,N_10523,N_12814);
or U15599 (N_15599,N_13293,N_12493);
xnor U15600 (N_15600,N_14495,N_11853);
nand U15601 (N_15601,N_11519,N_11759);
and U15602 (N_15602,N_11808,N_10017);
or U15603 (N_15603,N_12741,N_10714);
nand U15604 (N_15604,N_12911,N_12843);
and U15605 (N_15605,N_10544,N_10868);
and U15606 (N_15606,N_13581,N_11270);
nor U15607 (N_15607,N_12644,N_13155);
or U15608 (N_15608,N_10435,N_14561);
or U15609 (N_15609,N_14564,N_14424);
and U15610 (N_15610,N_14171,N_12726);
xor U15611 (N_15611,N_12783,N_12030);
nand U15612 (N_15612,N_10068,N_11903);
and U15613 (N_15613,N_10952,N_13844);
nor U15614 (N_15614,N_11504,N_13517);
nand U15615 (N_15615,N_11275,N_12174);
or U15616 (N_15616,N_10156,N_14511);
nand U15617 (N_15617,N_10455,N_12738);
or U15618 (N_15618,N_14329,N_11013);
nor U15619 (N_15619,N_14499,N_13191);
xnor U15620 (N_15620,N_14026,N_12936);
or U15621 (N_15621,N_11819,N_12447);
xnor U15622 (N_15622,N_10483,N_10212);
nand U15623 (N_15623,N_14139,N_10702);
nand U15624 (N_15624,N_11873,N_12670);
nand U15625 (N_15625,N_10627,N_10177);
and U15626 (N_15626,N_12416,N_10467);
or U15627 (N_15627,N_13523,N_14252);
and U15628 (N_15628,N_11113,N_12517);
nor U15629 (N_15629,N_14236,N_12042);
nor U15630 (N_15630,N_10451,N_11443);
and U15631 (N_15631,N_14869,N_12665);
nor U15632 (N_15632,N_13956,N_13960);
nand U15633 (N_15633,N_11204,N_12052);
nor U15634 (N_15634,N_12657,N_13230);
nor U15635 (N_15635,N_12474,N_13884);
nor U15636 (N_15636,N_13399,N_10822);
or U15637 (N_15637,N_11483,N_13068);
or U15638 (N_15638,N_10469,N_12408);
and U15639 (N_15639,N_12917,N_12133);
or U15640 (N_15640,N_14011,N_14089);
xnor U15641 (N_15641,N_11173,N_11406);
xor U15642 (N_15642,N_10299,N_10578);
and U15643 (N_15643,N_12137,N_12277);
xor U15644 (N_15644,N_11729,N_14170);
xnor U15645 (N_15645,N_13239,N_14233);
nor U15646 (N_15646,N_13661,N_12147);
xor U15647 (N_15647,N_13644,N_11321);
and U15648 (N_15648,N_11910,N_14318);
and U15649 (N_15649,N_11482,N_12372);
xnor U15650 (N_15650,N_11301,N_13758);
nand U15651 (N_15651,N_13650,N_13011);
nor U15652 (N_15652,N_13138,N_13910);
or U15653 (N_15653,N_14571,N_13604);
nand U15654 (N_15654,N_13346,N_11657);
and U15655 (N_15655,N_13052,N_10132);
or U15656 (N_15656,N_11105,N_12466);
or U15657 (N_15657,N_14168,N_12658);
or U15658 (N_15658,N_14796,N_10303);
or U15659 (N_15659,N_10222,N_14351);
nor U15660 (N_15660,N_13992,N_14331);
xnor U15661 (N_15661,N_11228,N_10851);
or U15662 (N_15662,N_11020,N_14414);
nor U15663 (N_15663,N_13952,N_11199);
nor U15664 (N_15664,N_14317,N_10973);
and U15665 (N_15665,N_12778,N_13829);
nor U15666 (N_15666,N_12158,N_13770);
nor U15667 (N_15667,N_10553,N_14454);
or U15668 (N_15668,N_13501,N_10453);
nand U15669 (N_15669,N_10402,N_10323);
xor U15670 (N_15670,N_11261,N_14280);
or U15671 (N_15671,N_11893,N_13083);
and U15672 (N_15672,N_10347,N_11886);
nor U15673 (N_15673,N_14178,N_13495);
and U15674 (N_15674,N_10661,N_13920);
or U15675 (N_15675,N_12724,N_13094);
or U15676 (N_15676,N_14042,N_14863);
and U15677 (N_15677,N_10886,N_13468);
or U15678 (N_15678,N_14625,N_10920);
nor U15679 (N_15679,N_11879,N_10179);
nand U15680 (N_15680,N_14115,N_11419);
or U15681 (N_15681,N_10819,N_11733);
nand U15682 (N_15682,N_13713,N_13814);
nand U15683 (N_15683,N_10443,N_13030);
and U15684 (N_15684,N_11981,N_11717);
or U15685 (N_15685,N_11388,N_13423);
nor U15686 (N_15686,N_14155,N_14996);
nand U15687 (N_15687,N_13326,N_13997);
or U15688 (N_15688,N_14881,N_13850);
or U15689 (N_15689,N_10161,N_12543);
or U15690 (N_15690,N_12097,N_14974);
nand U15691 (N_15691,N_14958,N_11376);
or U15692 (N_15692,N_14215,N_10691);
nor U15693 (N_15693,N_13979,N_11123);
and U15694 (N_15694,N_13267,N_14052);
nand U15695 (N_15695,N_14067,N_13648);
and U15696 (N_15696,N_12854,N_14854);
or U15697 (N_15697,N_10045,N_13606);
and U15698 (N_15698,N_10563,N_10022);
and U15699 (N_15699,N_13220,N_14687);
nor U15700 (N_15700,N_13727,N_13555);
nand U15701 (N_15701,N_10771,N_10915);
or U15702 (N_15702,N_12108,N_10823);
nand U15703 (N_15703,N_11825,N_14547);
xor U15704 (N_15704,N_10569,N_10157);
and U15705 (N_15705,N_11086,N_10668);
or U15706 (N_15706,N_13632,N_12812);
nand U15707 (N_15707,N_11506,N_13341);
and U15708 (N_15708,N_10704,N_10855);
or U15709 (N_15709,N_14635,N_14245);
and U15710 (N_15710,N_10406,N_12485);
and U15711 (N_15711,N_11777,N_10284);
nand U15712 (N_15712,N_13892,N_13752);
nor U15713 (N_15713,N_12265,N_13216);
or U15714 (N_15714,N_10368,N_11045);
and U15715 (N_15715,N_14918,N_14503);
or U15716 (N_15716,N_10273,N_11716);
nand U15717 (N_15717,N_14987,N_11761);
nand U15718 (N_15718,N_12000,N_12931);
and U15719 (N_15719,N_14537,N_14465);
and U15720 (N_15720,N_13772,N_11442);
xor U15721 (N_15721,N_10505,N_12995);
nor U15722 (N_15722,N_12841,N_12354);
and U15723 (N_15723,N_10922,N_11280);
and U15724 (N_15724,N_14109,N_11476);
nand U15725 (N_15725,N_12672,N_14492);
and U15726 (N_15726,N_14903,N_13403);
nand U15727 (N_15727,N_12353,N_12666);
and U15728 (N_15728,N_14374,N_12571);
and U15729 (N_15729,N_14468,N_11278);
and U15730 (N_15730,N_14111,N_13235);
or U15731 (N_15731,N_10432,N_14553);
xnor U15732 (N_15732,N_12395,N_14453);
or U15733 (N_15733,N_13506,N_12723);
nor U15734 (N_15734,N_10023,N_14783);
or U15735 (N_15735,N_13605,N_10194);
nor U15736 (N_15736,N_12997,N_14894);
and U15737 (N_15737,N_11635,N_12433);
and U15738 (N_15738,N_13930,N_14720);
nand U15739 (N_15739,N_10715,N_12139);
and U15740 (N_15740,N_13069,N_13711);
nand U15741 (N_15741,N_12597,N_14314);
nand U15742 (N_15742,N_13266,N_14939);
and U15743 (N_15743,N_10773,N_10458);
nand U15744 (N_15744,N_11374,N_11687);
nor U15745 (N_15745,N_12476,N_13572);
nor U15746 (N_15746,N_13595,N_11438);
and U15747 (N_15747,N_10014,N_10477);
nor U15748 (N_15748,N_14090,N_10126);
or U15749 (N_15749,N_14493,N_12445);
xnor U15750 (N_15750,N_14809,N_10918);
nand U15751 (N_15751,N_11059,N_10658);
nand U15752 (N_15752,N_14381,N_13212);
nand U15753 (N_15753,N_13469,N_12086);
and U15754 (N_15754,N_12313,N_10018);
nand U15755 (N_15755,N_14701,N_11680);
and U15756 (N_15756,N_13268,N_11404);
nand U15757 (N_15757,N_12387,N_11578);
xor U15758 (N_15758,N_13056,N_10009);
nor U15759 (N_15759,N_11225,N_14521);
nand U15760 (N_15760,N_13198,N_10674);
xor U15761 (N_15761,N_10486,N_10889);
nand U15762 (N_15762,N_12262,N_10011);
nor U15763 (N_15763,N_13778,N_13515);
nand U15764 (N_15764,N_11227,N_13183);
nor U15765 (N_15765,N_14758,N_10170);
nand U15766 (N_15766,N_12774,N_14705);
and U15767 (N_15767,N_10816,N_14595);
nor U15768 (N_15768,N_11477,N_11723);
or U15769 (N_15769,N_13740,N_14898);
nor U15770 (N_15770,N_11491,N_10776);
nand U15771 (N_15771,N_11709,N_10591);
or U15772 (N_15772,N_14340,N_10214);
nand U15773 (N_15773,N_12390,N_14645);
nand U15774 (N_15774,N_12481,N_14845);
nor U15775 (N_15775,N_11216,N_12515);
and U15776 (N_15776,N_10383,N_13487);
and U15777 (N_15777,N_12524,N_13634);
nor U15778 (N_15778,N_14394,N_12183);
or U15779 (N_15779,N_14538,N_13215);
nor U15780 (N_15780,N_10718,N_11554);
xor U15781 (N_15781,N_10987,N_12918);
or U15782 (N_15782,N_10765,N_10700);
and U15783 (N_15783,N_10910,N_14803);
or U15784 (N_15784,N_14648,N_11472);
and U15785 (N_15785,N_14530,N_10511);
and U15786 (N_15786,N_14076,N_14223);
nand U15787 (N_15787,N_11966,N_12106);
and U15788 (N_15788,N_13896,N_11656);
and U15789 (N_15789,N_12428,N_10562);
or U15790 (N_15790,N_11174,N_13516);
and U15791 (N_15791,N_14055,N_12540);
xor U15792 (N_15792,N_11566,N_11480);
nand U15793 (N_15793,N_14401,N_13462);
or U15794 (N_15794,N_14810,N_14945);
xnor U15795 (N_15795,N_13972,N_13032);
nor U15796 (N_15796,N_11646,N_13028);
nor U15797 (N_15797,N_13672,N_14937);
or U15798 (N_15798,N_10640,N_13141);
nor U15799 (N_15799,N_12884,N_13133);
nand U15800 (N_15800,N_11127,N_11907);
or U15801 (N_15801,N_10133,N_13354);
or U15802 (N_15802,N_12098,N_13729);
nand U15803 (N_15803,N_10167,N_11356);
nor U15804 (N_15804,N_12586,N_11400);
nand U15805 (N_15805,N_11901,N_12388);
and U15806 (N_15806,N_11695,N_13223);
and U15807 (N_15807,N_10546,N_14589);
nor U15808 (N_15808,N_11816,N_11265);
xnor U15809 (N_15809,N_13351,N_12488);
nand U15810 (N_15810,N_12409,N_10039);
nor U15811 (N_15811,N_13913,N_10440);
nor U15812 (N_15812,N_10900,N_10926);
and U15813 (N_15813,N_12798,N_12170);
nor U15814 (N_15814,N_12197,N_14893);
xor U15815 (N_15815,N_13853,N_11399);
and U15816 (N_15816,N_14921,N_10902);
and U15817 (N_15817,N_11500,N_13208);
or U15818 (N_15818,N_14378,N_13966);
and U15819 (N_15819,N_12584,N_11152);
nand U15820 (N_15820,N_14970,N_14906);
nand U15821 (N_15821,N_12314,N_13808);
and U15822 (N_15822,N_14102,N_12506);
or U15823 (N_15823,N_10541,N_11300);
or U15824 (N_15824,N_13526,N_10580);
nor U15825 (N_15825,N_14429,N_10906);
nand U15826 (N_15826,N_12091,N_12740);
and U15827 (N_15827,N_12576,N_11360);
nor U15828 (N_15828,N_12756,N_13441);
nor U15829 (N_15829,N_14469,N_14856);
nand U15830 (N_15830,N_13950,N_10712);
nand U15831 (N_15831,N_11595,N_11594);
and U15832 (N_15832,N_12307,N_10145);
nand U15833 (N_15833,N_14743,N_13221);
nor U15834 (N_15834,N_10048,N_11525);
or U15835 (N_15835,N_13347,N_11782);
or U15836 (N_15836,N_11136,N_10035);
or U15837 (N_15837,N_13990,N_10271);
and U15838 (N_15838,N_11495,N_10116);
xnor U15839 (N_15839,N_14988,N_11203);
and U15840 (N_15840,N_11198,N_12776);
or U15841 (N_15841,N_12007,N_14896);
xnor U15842 (N_15842,N_10760,N_14670);
nor U15843 (N_15843,N_10027,N_12209);
or U15844 (N_15844,N_13553,N_14071);
nor U15845 (N_15845,N_11678,N_13815);
nand U15846 (N_15846,N_14634,N_11748);
nand U15847 (N_15847,N_10342,N_12430);
and U15848 (N_15848,N_12011,N_11365);
or U15849 (N_15849,N_11663,N_13989);
and U15850 (N_15850,N_13014,N_12441);
and U15851 (N_15851,N_11096,N_12195);
or U15852 (N_15852,N_11538,N_13701);
nand U15853 (N_15853,N_13398,N_12617);
or U15854 (N_15854,N_12206,N_11053);
and U15855 (N_15855,N_12026,N_13428);
nand U15856 (N_15856,N_11739,N_10893);
and U15857 (N_15857,N_11055,N_13188);
nand U15858 (N_15858,N_11079,N_10721);
nand U15859 (N_15859,N_11415,N_14741);
or U15860 (N_15860,N_14647,N_13182);
xnor U15861 (N_15861,N_10928,N_10907);
nor U15862 (N_15862,N_12560,N_10639);
nand U15863 (N_15863,N_14827,N_11628);
xnor U15864 (N_15864,N_14486,N_10463);
and U15865 (N_15865,N_11820,N_13435);
nor U15866 (N_15866,N_11977,N_14391);
xor U15867 (N_15867,N_11051,N_10768);
xnor U15868 (N_15868,N_14852,N_11862);
nand U15869 (N_15869,N_14982,N_11245);
or U15870 (N_15870,N_14942,N_10741);
or U15871 (N_15871,N_14730,N_12196);
xor U15872 (N_15872,N_13470,N_11823);
or U15873 (N_15873,N_10972,N_12949);
nor U15874 (N_15874,N_12627,N_12398);
or U15875 (N_15875,N_11743,N_14962);
and U15876 (N_15876,N_10457,N_11985);
xor U15877 (N_15877,N_14968,N_11089);
xor U15878 (N_15878,N_10515,N_12501);
nor U15879 (N_15879,N_13091,N_10313);
xnor U15880 (N_15880,N_12419,N_12414);
xnor U15881 (N_15881,N_10242,N_12809);
and U15882 (N_15882,N_12680,N_11529);
nand U15883 (N_15883,N_14020,N_13607);
or U15884 (N_15884,N_11217,N_14084);
nor U15885 (N_15885,N_13580,N_11790);
nand U15886 (N_15886,N_12921,N_11110);
xor U15887 (N_15887,N_14013,N_13484);
or U15888 (N_15888,N_11814,N_10977);
nand U15889 (N_15889,N_11535,N_11802);
nand U15890 (N_15890,N_13530,N_13119);
and U15891 (N_15891,N_11585,N_12222);
and U15892 (N_15892,N_13571,N_14792);
xor U15893 (N_15893,N_13805,N_12235);
nand U15894 (N_15894,N_10137,N_14149);
or U15895 (N_15895,N_14093,N_14293);
nor U15896 (N_15896,N_13888,N_13783);
or U15897 (N_15897,N_10302,N_10615);
and U15898 (N_15898,N_10331,N_14153);
xor U15899 (N_15899,N_10846,N_14870);
or U15900 (N_15900,N_13010,N_13000);
xnor U15901 (N_15901,N_13373,N_10625);
nand U15902 (N_15902,N_10233,N_12203);
nor U15903 (N_15903,N_13935,N_10056);
and U15904 (N_15904,N_13364,N_11592);
or U15905 (N_15905,N_13674,N_13274);
nand U15906 (N_15906,N_14901,N_12221);
nor U15907 (N_15907,N_10601,N_11924);
nor U15908 (N_15908,N_14319,N_11527);
nand U15909 (N_15909,N_10521,N_14943);
nor U15910 (N_15910,N_10445,N_10288);
and U15911 (N_15911,N_14549,N_12888);
and U15912 (N_15912,N_14002,N_13040);
nor U15913 (N_15913,N_10310,N_13016);
or U15914 (N_15914,N_10770,N_11530);
nand U15915 (N_15915,N_11848,N_12789);
nand U15916 (N_15916,N_12861,N_12818);
xnor U15917 (N_15917,N_10366,N_14728);
nand U15918 (N_15918,N_11781,N_11852);
nand U15919 (N_15919,N_13431,N_14270);
nor U15920 (N_15920,N_12328,N_13931);
xnor U15921 (N_15921,N_10747,N_14606);
nand U15922 (N_15922,N_11640,N_12731);
or U15923 (N_15923,N_13623,N_13622);
and U15924 (N_15924,N_11710,N_11493);
nand U15925 (N_15925,N_11744,N_13053);
and U15926 (N_15926,N_11764,N_12541);
or U15927 (N_15927,N_13429,N_14501);
nor U15928 (N_15928,N_13999,N_11069);
or U15929 (N_15929,N_13706,N_13345);
and U15930 (N_15930,N_14655,N_11027);
nor U15931 (N_15931,N_11344,N_14626);
or U15932 (N_15932,N_10588,N_12971);
nor U15933 (N_15933,N_10386,N_12688);
or U15934 (N_15934,N_13292,N_12341);
or U15935 (N_15935,N_13780,N_12598);
or U15936 (N_15936,N_14120,N_13314);
or U15937 (N_15937,N_14096,N_13785);
nor U15938 (N_15938,N_11908,N_11159);
nand U15939 (N_15939,N_11363,N_10307);
and U15940 (N_15940,N_11185,N_13418);
xnor U15941 (N_15941,N_13682,N_13870);
nor U15942 (N_15942,N_14604,N_13591);
or U15943 (N_15943,N_13272,N_10238);
xnor U15944 (N_15944,N_14368,N_13343);
nand U15945 (N_15945,N_12249,N_11892);
xor U15946 (N_15946,N_12664,N_11184);
nand U15947 (N_15947,N_14580,N_12171);
and U15948 (N_15948,N_14695,N_11333);
nand U15949 (N_15949,N_14387,N_10046);
nor U15950 (N_15950,N_12976,N_10180);
nor U15951 (N_15951,N_13965,N_13420);
nor U15952 (N_15952,N_11232,N_14734);
xor U15953 (N_15953,N_12082,N_14608);
nand U15954 (N_15954,N_14231,N_12323);
and U15955 (N_15955,N_13492,N_12228);
and U15956 (N_15956,N_12897,N_13696);
nand U15957 (N_15957,N_12566,N_13944);
or U15958 (N_15958,N_14187,N_12825);
nand U15959 (N_15959,N_12459,N_13566);
nor U15960 (N_15960,N_11511,N_12739);
nand U15961 (N_15961,N_12165,N_14596);
xnor U15962 (N_15962,N_11414,N_11490);
nor U15963 (N_15963,N_14010,N_14578);
and U15964 (N_15964,N_11518,N_12331);
or U15965 (N_15965,N_14609,N_12792);
nor U15966 (N_15966,N_12294,N_12074);
and U15967 (N_15967,N_13360,N_10603);
or U15968 (N_15968,N_11259,N_10946);
and U15969 (N_15969,N_10149,N_13904);
nor U15970 (N_15970,N_10183,N_14259);
nor U15971 (N_15971,N_11643,N_14698);
or U15972 (N_15972,N_12397,N_12591);
xor U15973 (N_15973,N_10150,N_11396);
and U15974 (N_15974,N_14665,N_10241);
or U15975 (N_15975,N_14615,N_10360);
and U15976 (N_15976,N_14058,N_13051);
and U15977 (N_15977,N_14960,N_14712);
or U15978 (N_15978,N_10629,N_13107);
nor U15979 (N_15979,N_14713,N_13147);
nand U15980 (N_15980,N_12523,N_11932);
or U15981 (N_15981,N_12819,N_11064);
xnor U15982 (N_15982,N_14281,N_10392);
nand U15983 (N_15983,N_12226,N_12487);
and U15984 (N_15984,N_12568,N_10685);
xnor U15985 (N_15985,N_11858,N_12268);
nor U15986 (N_15986,N_13251,N_10158);
nor U15987 (N_15987,N_12283,N_13524);
nor U15988 (N_15988,N_11429,N_10847);
nand U15989 (N_15989,N_11916,N_14771);
and U15990 (N_15990,N_12366,N_12526);
or U15991 (N_15991,N_12320,N_12630);
nor U15992 (N_15992,N_13087,N_14820);
and U15993 (N_15993,N_11417,N_10185);
nand U15994 (N_15994,N_13277,N_11972);
xor U15995 (N_15995,N_10205,N_10178);
nor U15996 (N_15996,N_10675,N_10947);
xnor U15997 (N_15997,N_13568,N_13299);
nand U15998 (N_15998,N_13895,N_14932);
and U15999 (N_15999,N_12066,N_14175);
nand U16000 (N_16000,N_10646,N_13898);
nand U16001 (N_16001,N_12986,N_11548);
xnor U16002 (N_16002,N_14699,N_13626);
and U16003 (N_16003,N_14992,N_10626);
or U16004 (N_16004,N_13830,N_10282);
nor U16005 (N_16005,N_13167,N_14242);
nand U16006 (N_16006,N_14834,N_10951);
nor U16007 (N_16007,N_10098,N_14879);
xor U16008 (N_16008,N_14915,N_13452);
and U16009 (N_16009,N_11351,N_12004);
nor U16010 (N_16010,N_13285,N_10528);
or U16011 (N_16011,N_12104,N_14162);
nand U16012 (N_16012,N_13874,N_10204);
nand U16013 (N_16013,N_14582,N_14823);
or U16014 (N_16014,N_10028,N_12772);
nand U16015 (N_16015,N_14983,N_12422);
or U16016 (N_16016,N_10206,N_12530);
nor U16017 (N_16017,N_13919,N_10159);
or U16018 (N_16018,N_10496,N_14496);
or U16019 (N_16019,N_10527,N_12111);
or U16020 (N_16020,N_12048,N_11815);
nand U16021 (N_16021,N_11104,N_13873);
and U16022 (N_16022,N_10087,N_10136);
nor U16023 (N_16023,N_10289,N_14559);
nand U16024 (N_16024,N_12118,N_14899);
or U16025 (N_16025,N_11091,N_12112);
nor U16026 (N_16026,N_10985,N_10217);
xor U16027 (N_16027,N_12344,N_11426);
nor U16028 (N_16028,N_14628,N_12706);
nand U16029 (N_16029,N_11170,N_10677);
nand U16030 (N_16030,N_14257,N_13779);
nor U16031 (N_16031,N_10165,N_10666);
and U16032 (N_16032,N_14282,N_14024);
or U16033 (N_16033,N_10964,N_13583);
or U16034 (N_16034,N_14662,N_13624);
xor U16035 (N_16035,N_13005,N_12863);
xnor U16036 (N_16036,N_11024,N_12116);
nor U16037 (N_16037,N_12044,N_12990);
and U16038 (N_16038,N_11994,N_14152);
nor U16039 (N_16039,N_13232,N_10943);
and U16040 (N_16040,N_14522,N_14873);
and U16041 (N_16041,N_13574,N_10163);
or U16042 (N_16042,N_11048,N_11172);
nand U16043 (N_16043,N_13315,N_13284);
xor U16044 (N_16044,N_13286,N_14534);
and U16045 (N_16045,N_11626,N_12271);
and U16046 (N_16046,N_13959,N_11670);
or U16047 (N_16047,N_11456,N_10871);
nand U16048 (N_16048,N_13640,N_14421);
nor U16049 (N_16049,N_13669,N_13927);
nor U16050 (N_16050,N_11951,N_13042);
nand U16051 (N_16051,N_12391,N_14467);
or U16052 (N_16052,N_13355,N_12109);
and U16053 (N_16053,N_13279,N_13686);
xnor U16054 (N_16054,N_12559,N_14266);
or U16055 (N_16055,N_10692,N_12991);
or U16056 (N_16056,N_13003,N_10512);
nand U16057 (N_16057,N_10403,N_10738);
nor U16058 (N_16058,N_10579,N_13507);
nand U16059 (N_16059,N_10739,N_13331);
or U16060 (N_16060,N_11146,N_14008);
nor U16061 (N_16061,N_14239,N_13357);
nand U16062 (N_16062,N_13908,N_12308);
xnor U16063 (N_16063,N_12900,N_11798);
nor U16064 (N_16064,N_13550,N_13911);
or U16065 (N_16065,N_12535,N_12747);
or U16066 (N_16066,N_10508,N_14737);
and U16067 (N_16067,N_13876,N_10689);
and U16068 (N_16068,N_12411,N_11724);
nand U16069 (N_16069,N_14723,N_10131);
or U16070 (N_16070,N_12934,N_14386);
and U16071 (N_16071,N_11061,N_12164);
or U16072 (N_16072,N_13840,N_10762);
and U16073 (N_16073,N_14799,N_14349);
or U16074 (N_16074,N_11137,N_14227);
and U16075 (N_16075,N_11722,N_13417);
or U16076 (N_16076,N_13652,N_12149);
and U16077 (N_16077,N_10506,N_10318);
and U16078 (N_16078,N_12573,N_12827);
xor U16079 (N_16079,N_11090,N_14462);
nand U16080 (N_16080,N_10099,N_10736);
nor U16081 (N_16081,N_12077,N_11934);
nor U16082 (N_16082,N_11963,N_11728);
nand U16083 (N_16083,N_10407,N_14614);
or U16084 (N_16084,N_11667,N_11588);
nand U16085 (N_16085,N_10695,N_13718);
or U16086 (N_16086,N_11366,N_13242);
and U16087 (N_16087,N_13597,N_13641);
nor U16088 (N_16088,N_10186,N_11183);
nand U16089 (N_16089,N_14095,N_11532);
and U16090 (N_16090,N_12367,N_12306);
xor U16091 (N_16091,N_12650,N_14950);
nand U16092 (N_16092,N_13544,N_13145);
nor U16093 (N_16093,N_14078,N_14416);
and U16094 (N_16094,N_14726,N_13925);
or U16095 (N_16095,N_14348,N_14776);
or U16096 (N_16096,N_10698,N_13985);
and U16097 (N_16097,N_12198,N_12274);
and U16098 (N_16098,N_11758,N_13891);
nand U16099 (N_16099,N_11943,N_13152);
xnor U16100 (N_16100,N_11803,N_13474);
and U16101 (N_16101,N_14250,N_12496);
nand U16102 (N_16102,N_11361,N_13224);
and U16103 (N_16103,N_11034,N_10824);
and U16104 (N_16104,N_12983,N_11391);
nand U16105 (N_16105,N_14875,N_10267);
nor U16106 (N_16106,N_13735,N_10705);
nor U16107 (N_16107,N_13940,N_14836);
nor U16108 (N_16108,N_14385,N_12495);
nor U16109 (N_16109,N_12557,N_13067);
and U16110 (N_16110,N_13205,N_14917);
xnor U16111 (N_16111,N_10708,N_14234);
nor U16112 (N_16112,N_12463,N_11639);
and U16113 (N_16113,N_13055,N_14643);
nand U16114 (N_16114,N_10835,N_12992);
nor U16115 (N_16115,N_11390,N_10441);
and U16116 (N_16116,N_13736,N_13792);
nand U16117 (N_16117,N_11770,N_10199);
and U16118 (N_16118,N_14044,N_10434);
nor U16119 (N_16119,N_14545,N_11000);
and U16120 (N_16120,N_12187,N_11637);
xor U16121 (N_16121,N_10940,N_12647);
xor U16122 (N_16122,N_10936,N_10643);
or U16123 (N_16123,N_12528,N_11843);
and U16124 (N_16124,N_14306,N_13007);
or U16125 (N_16125,N_13471,N_13788);
nor U16126 (N_16126,N_14376,N_14888);
nor U16127 (N_16127,N_14764,N_10276);
nor U16128 (N_16128,N_13570,N_14261);
nand U16129 (N_16129,N_11121,N_14279);
and U16130 (N_16130,N_10683,N_13012);
and U16131 (N_16131,N_12869,N_14460);
nor U16132 (N_16132,N_11850,N_12615);
nor U16133 (N_16133,N_12385,N_10808);
nand U16134 (N_16134,N_14023,N_10315);
or U16135 (N_16135,N_11492,N_10649);
xnor U16136 (N_16136,N_13057,N_14622);
or U16137 (N_16137,N_12759,N_14599);
and U16138 (N_16138,N_12642,N_14569);
or U16139 (N_16139,N_13020,N_10516);
nor U16140 (N_16140,N_11515,N_14337);
nor U16141 (N_16141,N_11524,N_13275);
and U16142 (N_16142,N_10959,N_11730);
or U16143 (N_16143,N_12786,N_13443);
xor U16144 (N_16144,N_11276,N_11560);
xnor U16145 (N_16145,N_11546,N_14829);
nor U16146 (N_16146,N_12039,N_14504);
nor U16147 (N_16147,N_13106,N_13759);
nand U16148 (N_16148,N_14164,N_11913);
nand U16149 (N_16149,N_13703,N_11140);
and U16150 (N_16150,N_10690,N_12134);
or U16151 (N_16151,N_11302,N_12299);
nand U16152 (N_16152,N_10024,N_13334);
nand U16153 (N_16153,N_12362,N_11195);
nor U16154 (N_16154,N_14548,N_11954);
and U16155 (N_16155,N_11817,N_13393);
or U16156 (N_16156,N_10245,N_14366);
nand U16157 (N_16157,N_14969,N_13344);
and U16158 (N_16158,N_14624,N_13427);
or U16159 (N_16159,N_10164,N_14889);
nand U16160 (N_16160,N_12720,N_13588);
xor U16161 (N_16161,N_13863,N_12904);
nor U16162 (N_16162,N_14016,N_12625);
or U16163 (N_16163,N_12368,N_14437);
or U16164 (N_16164,N_12736,N_12507);
xnor U16165 (N_16165,N_11233,N_13693);
xor U16166 (N_16166,N_11274,N_11033);
nand U16167 (N_16167,N_14878,N_12284);
and U16168 (N_16168,N_14927,N_13490);
or U16169 (N_16169,N_12010,N_12710);
nand U16170 (N_16170,N_10262,N_14063);
and U16171 (N_16171,N_12705,N_13811);
or U16172 (N_16172,N_14639,N_14715);
xor U16173 (N_16173,N_12179,N_10600);
and U16174 (N_16174,N_12335,N_12212);
nor U16175 (N_16175,N_12690,N_11016);
xor U16176 (N_16176,N_12272,N_13619);
nand U16177 (N_16177,N_10885,N_13962);
or U16178 (N_16178,N_12893,N_11784);
nand U16179 (N_16179,N_12959,N_12325);
and U16180 (N_16180,N_10993,N_12497);
and U16181 (N_16181,N_14230,N_12460);
nor U16182 (N_16182,N_10290,N_13533);
nand U16183 (N_16183,N_13402,N_12383);
nand U16184 (N_16184,N_13457,N_11081);
nor U16185 (N_16185,N_13329,N_10000);
nor U16186 (N_16186,N_14031,N_11329);
nand U16187 (N_16187,N_14831,N_13044);
or U16188 (N_16188,N_11557,N_11407);
or U16189 (N_16189,N_11941,N_11435);
nor U16190 (N_16190,N_12652,N_10355);
nand U16191 (N_16191,N_14146,N_13022);
or U16192 (N_16192,N_13207,N_13941);
nand U16193 (N_16193,N_11854,N_14912);
and U16194 (N_16194,N_10456,N_13015);
or U16195 (N_16195,N_13508,N_13158);
nor U16196 (N_16196,N_12556,N_14411);
or U16197 (N_16197,N_14729,N_10616);
nor U16198 (N_16198,N_11403,N_12796);
nor U16199 (N_16199,N_12301,N_12233);
and U16200 (N_16200,N_12257,N_11882);
xor U16201 (N_16201,N_10013,N_10495);
nor U16202 (N_16202,N_10171,N_14338);
nand U16203 (N_16203,N_12599,N_10867);
nor U16204 (N_16204,N_11211,N_13189);
nor U16205 (N_16205,N_13929,N_11194);
or U16206 (N_16206,N_13476,N_10622);
or U16207 (N_16207,N_13058,N_10888);
xor U16208 (N_16208,N_11599,N_13510);
or U16209 (N_16209,N_14871,N_10929);
or U16210 (N_16210,N_11303,N_13405);
and U16211 (N_16211,N_14818,N_14587);
and U16212 (N_16212,N_13865,N_13154);
and U16213 (N_16213,N_10081,N_11976);
and U16214 (N_16214,N_12309,N_12727);
nand U16215 (N_16215,N_13968,N_12902);
nor U16216 (N_16216,N_11634,N_11171);
nor U16217 (N_16217,N_11914,N_14585);
xor U16218 (N_16218,N_12579,N_13737);
nor U16219 (N_16219,N_11650,N_14316);
nor U16220 (N_16220,N_14258,N_14719);
nand U16221 (N_16221,N_10681,N_12677);
nor U16222 (N_16222,N_12580,N_11675);
and U16223 (N_16223,N_12273,N_11615);
and U16224 (N_16224,N_10782,N_12996);
nor U16225 (N_16225,N_14989,N_11536);
nor U16226 (N_16226,N_11542,N_13348);
and U16227 (N_16227,N_11154,N_14920);
nand U16228 (N_16228,N_10264,N_14151);
or U16229 (N_16229,N_11028,N_14154);
or U16230 (N_16230,N_10631,N_11169);
or U16231 (N_16231,N_14990,N_10107);
and U16232 (N_16232,N_14425,N_10903);
and U16233 (N_16233,N_10686,N_11944);
nor U16234 (N_16234,N_14664,N_14890);
xor U16235 (N_16235,N_12213,N_11297);
or U16236 (N_16236,N_14405,N_13667);
or U16237 (N_16237,N_11145,N_10484);
nor U16238 (N_16238,N_12205,N_12749);
nand U16239 (N_16239,N_13233,N_14964);
nand U16240 (N_16240,N_12347,N_12285);
nor U16241 (N_16241,N_13678,N_13953);
nor U16242 (N_16242,N_11118,N_10409);
nand U16243 (N_16243,N_13630,N_12450);
nand U16244 (N_16244,N_12563,N_12942);
nand U16245 (N_16245,N_14434,N_13132);
or U16246 (N_16246,N_12336,N_11684);
nor U16247 (N_16247,N_10599,N_14295);
and U16248 (N_16248,N_11836,N_13864);
nor U16249 (N_16249,N_10955,N_10142);
and U16250 (N_16250,N_13651,N_11249);
or U16251 (N_16251,N_13745,N_14129);
nor U16252 (N_16252,N_10067,N_10684);
or U16253 (N_16253,N_12901,N_11771);
xnor U16254 (N_16254,N_13372,N_12761);
nor U16255 (N_16255,N_14885,N_12871);
or U16256 (N_16256,N_14262,N_10334);
and U16257 (N_16257,N_12547,N_14124);
xnor U16258 (N_16258,N_14080,N_10433);
nor U16259 (N_16259,N_10375,N_10041);
and U16260 (N_16260,N_13846,N_12015);
nand U16261 (N_16261,N_14887,N_11192);
nor U16262 (N_16262,N_12955,N_13071);
or U16263 (N_16263,N_11057,N_10079);
nand U16264 (N_16264,N_14977,N_11806);
or U16265 (N_16265,N_11181,N_10112);
or U16266 (N_16266,N_12019,N_12847);
and U16267 (N_16267,N_11718,N_10873);
and U16268 (N_16268,N_12477,N_13123);
nand U16269 (N_16269,N_10565,N_12508);
and U16270 (N_16270,N_10200,N_10948);
nand U16271 (N_16271,N_11328,N_10949);
nand U16272 (N_16272,N_11652,N_12375);
and U16273 (N_16273,N_14253,N_10892);
or U16274 (N_16274,N_10227,N_12009);
or U16275 (N_16275,N_12674,N_11004);
nor U16276 (N_16276,N_13646,N_14805);
and U16277 (N_16277,N_11734,N_11250);
nor U16278 (N_16278,N_13496,N_11720);
and U16279 (N_16279,N_14325,N_12245);
or U16280 (N_16280,N_13160,N_11230);
xnor U16281 (N_16281,N_14389,N_10193);
nand U16282 (N_16282,N_12330,N_13699);
or U16283 (N_16283,N_12346,N_11818);
and U16284 (N_16284,N_12908,N_14638);
and U16285 (N_16285,N_13171,N_11372);
nor U16286 (N_16286,N_10574,N_14954);
or U16287 (N_16287,N_11019,N_13868);
xnor U16288 (N_16288,N_12215,N_12551);
or U16289 (N_16289,N_13519,N_14583);
nor U16290 (N_16290,N_12697,N_14933);
nor U16291 (N_16291,N_11740,N_13349);
and U16292 (N_16292,N_14613,N_13629);
and U16293 (N_16293,N_10613,N_14277);
or U16294 (N_16294,N_13209,N_13685);
nand U16295 (N_16295,N_13882,N_12237);
and U16296 (N_16296,N_12851,N_10781);
nand U16297 (N_16297,N_13156,N_10143);
or U16298 (N_16298,N_14435,N_14466);
or U16299 (N_16299,N_13796,N_14264);
nor U16300 (N_16300,N_12499,N_11207);
or U16301 (N_16301,N_14816,N_12952);
and U16302 (N_16302,N_14186,N_10259);
or U16303 (N_16303,N_14991,N_10766);
nand U16304 (N_16304,N_13065,N_13532);
and U16305 (N_16305,N_12655,N_14700);
or U16306 (N_16306,N_11281,N_14021);
nand U16307 (N_16307,N_11970,N_13444);
or U16308 (N_16308,N_11268,N_12966);
and U16309 (N_16309,N_13070,N_14304);
nor U16310 (N_16310,N_10083,N_11191);
xnor U16311 (N_16311,N_14110,N_13464);
nand U16312 (N_16312,N_10536,N_11349);
nand U16313 (N_16313,N_12972,N_14074);
nand U16314 (N_16314,N_12096,N_14922);
nor U16315 (N_16315,N_11294,N_11296);
nor U16316 (N_16316,N_13244,N_14907);
nor U16317 (N_16317,N_11647,N_10751);
or U16318 (N_16318,N_13522,N_14138);
nand U16319 (N_16319,N_11143,N_10129);
nand U16320 (N_16320,N_14428,N_10826);
or U16321 (N_16321,N_13800,N_12337);
nor U16322 (N_16322,N_11083,N_12394);
nand U16323 (N_16323,N_12663,N_13404);
nand U16324 (N_16324,N_14800,N_13905);
or U16325 (N_16325,N_11837,N_10537);
nor U16326 (N_16326,N_14121,N_12189);
nand U16327 (N_16327,N_12607,N_14009);
and U16328 (N_16328,N_10461,N_12889);
and U16329 (N_16329,N_12359,N_12587);
nand U16330 (N_16330,N_12662,N_10927);
nand U16331 (N_16331,N_12371,N_14697);
or U16332 (N_16332,N_13851,N_14113);
nor U16333 (N_16333,N_10155,N_13340);
nand U16334 (N_16334,N_11935,N_10216);
or U16335 (N_16335,N_11014,N_14546);
nand U16336 (N_16336,N_14305,N_14505);
nor U16337 (N_16337,N_11179,N_11967);
or U16338 (N_16338,N_10358,N_14370);
nor U16339 (N_16339,N_10593,N_11671);
and U16340 (N_16340,N_10176,N_11078);
xnor U16341 (N_16341,N_11340,N_13902);
xor U16342 (N_16342,N_11458,N_14742);
or U16343 (N_16343,N_11487,N_11220);
or U16344 (N_16344,N_14984,N_12877);
or U16345 (N_16345,N_13409,N_11603);
and U16346 (N_16346,N_12687,N_11370);
or U16347 (N_16347,N_13150,N_10984);
xor U16348 (N_16348,N_10576,N_14515);
or U16349 (N_16349,N_11299,N_14517);
nand U16350 (N_16350,N_12604,N_14956);
and U16351 (N_16351,N_10992,N_13382);
or U16352 (N_16352,N_10783,N_12470);
or U16353 (N_16353,N_13240,N_10941);
nor U16354 (N_16354,N_11087,N_12938);
nand U16355 (N_16355,N_10115,N_11425);
nor U16356 (N_16356,N_14312,N_12924);
nor U16357 (N_16357,N_14355,N_11424);
nand U16358 (N_16358,N_11824,N_13301);
nand U16359 (N_16359,N_14787,N_13528);
and U16360 (N_16360,N_12185,N_14855);
nand U16361 (N_16361,N_13381,N_10120);
and U16362 (N_16362,N_13419,N_13248);
and U16363 (N_16363,N_10641,N_13807);
and U16364 (N_16364,N_14265,N_13324);
nor U16365 (N_16365,N_13932,N_11284);
nand U16366 (N_16366,N_13679,N_11844);
and U16367 (N_16367,N_12322,N_12763);
nor U16368 (N_16368,N_14759,N_14286);
nor U16369 (N_16369,N_13818,N_12883);
nor U16370 (N_16370,N_10950,N_11573);
nor U16371 (N_16371,N_11659,N_12227);
and U16372 (N_16372,N_11108,N_14848);
nand U16373 (N_16373,N_10270,N_11958);
nand U16374 (N_16374,N_10468,N_11805);
or U16375 (N_16375,N_14358,N_14422);
and U16376 (N_16376,N_10111,N_10657);
and U16377 (N_16377,N_13196,N_13378);
and U16378 (N_16378,N_13465,N_10938);
nor U16379 (N_16379,N_10317,N_14475);
nand U16380 (N_16380,N_10320,N_11610);
and U16381 (N_16381,N_11833,N_14196);
or U16382 (N_16382,N_14273,N_14751);
and U16383 (N_16383,N_13602,N_14694);
nor U16384 (N_16384,N_14494,N_12849);
nand U16385 (N_16385,N_10983,N_10479);
or U16386 (N_16386,N_12162,N_13416);
and U16387 (N_16387,N_12939,N_10539);
and U16388 (N_16388,N_11822,N_14483);
and U16389 (N_16389,N_12186,N_11315);
nand U16390 (N_16390,N_10858,N_14324);
and U16391 (N_16391,N_12489,N_12240);
nand U16392 (N_16392,N_12678,N_11364);
nor U16393 (N_16393,N_10422,N_14909);
nand U16394 (N_16394,N_13880,N_11642);
xor U16395 (N_16395,N_14631,N_10897);
nand U16396 (N_16396,N_12013,N_10103);
xor U16397 (N_16397,N_11962,N_10540);
and U16398 (N_16398,N_13151,N_13514);
nand U16399 (N_16399,N_11065,N_11448);
xor U16400 (N_16400,N_13795,N_11965);
or U16401 (N_16401,N_10359,N_11666);
nand U16402 (N_16402,N_10378,N_13271);
or U16403 (N_16403,N_14600,N_14116);
and U16404 (N_16404,N_12813,N_11165);
xnor U16405 (N_16405,N_10034,N_11887);
xnor U16406 (N_16406,N_14053,N_10680);
and U16407 (N_16407,N_11049,N_12797);
or U16408 (N_16408,N_14617,N_13958);
nor U16409 (N_16409,N_14825,N_14255);
and U16410 (N_16410,N_14691,N_14323);
and U16411 (N_16411,N_14769,N_14971);
nand U16412 (N_16412,N_11387,N_12637);
xnor U16413 (N_16413,N_11677,N_13073);
or U16414 (N_16414,N_11255,N_13980);
and U16415 (N_16415,N_13720,N_13479);
nor U16416 (N_16416,N_12334,N_10571);
nor U16417 (N_16417,N_14427,N_12502);
nand U16418 (N_16418,N_11469,N_10891);
or U16419 (N_16419,N_10919,N_10042);
and U16420 (N_16420,N_12001,N_11875);
nor U16421 (N_16421,N_14449,N_14260);
and U16422 (N_16422,N_10428,N_13694);
nor U16423 (N_16423,N_14438,N_14356);
and U16424 (N_16424,N_10988,N_14770);
nand U16425 (N_16425,N_14822,N_11032);
xor U16426 (N_16426,N_12636,N_14473);
xor U16427 (N_16427,N_14657,N_14123);
or U16428 (N_16428,N_11576,N_10044);
and U16429 (N_16429,N_12092,N_12800);
or U16430 (N_16430,N_11590,N_10326);
nor U16431 (N_16431,N_10376,N_11696);
or U16432 (N_16432,N_11840,N_14811);
nand U16433 (N_16433,N_13690,N_13178);
nor U16434 (N_16434,N_11035,N_14523);
or U16435 (N_16435,N_14481,N_13971);
and U16436 (N_16436,N_10006,N_12002);
or U16437 (N_16437,N_13045,N_10595);
or U16438 (N_16438,N_11241,N_14579);
or U16439 (N_16439,N_11679,N_14004);
nor U16440 (N_16440,N_14801,N_10113);
or U16441 (N_16441,N_13304,N_10957);
nand U16442 (N_16442,N_12480,N_13774);
nor U16443 (N_16443,N_14092,N_10904);
and U16444 (N_16444,N_10894,N_10364);
or U16445 (N_16445,N_14588,N_10935);
nor U16446 (N_16446,N_10232,N_10829);
and U16447 (N_16447,N_10882,N_10476);
or U16448 (N_16448,N_12844,N_12243);
or U16449 (N_16449,N_14377,N_12041);
nand U16450 (N_16450,N_11088,N_14938);
and U16451 (N_16451,N_13282,N_13467);
nand U16452 (N_16452,N_14780,N_14946);
or U16453 (N_16453,N_14005,N_14830);
xnor U16454 (N_16454,N_12423,N_12985);
nand U16455 (N_16455,N_14417,N_14563);
and U16456 (N_16456,N_12453,N_12865);
and U16457 (N_16457,N_10286,N_13136);
xnor U16458 (N_16458,N_13237,N_14762);
xor U16459 (N_16459,N_12808,N_14763);
xnor U16460 (N_16460,N_13365,N_13986);
or U16461 (N_16461,N_12369,N_14688);
xnor U16462 (N_16462,N_14430,N_10575);
nor U16463 (N_16463,N_12518,N_13757);
or U16464 (N_16464,N_14678,N_11313);
nor U16465 (N_16465,N_11624,N_10991);
nor U16466 (N_16466,N_14748,N_10610);
xor U16467 (N_16467,N_12632,N_14669);
nor U16468 (N_16468,N_12377,N_13095);
nor U16469 (N_16469,N_11672,N_13907);
nor U16470 (N_16470,N_13002,N_13482);
or U16471 (N_16471,N_13124,N_11002);
and U16472 (N_16472,N_12258,N_10731);
nand U16473 (N_16473,N_11936,N_13589);
nor U16474 (N_16474,N_14802,N_11358);
and U16475 (N_16475,N_11604,N_11009);
nor U16476 (N_16476,N_14298,N_10312);
xnor U16477 (N_16477,N_10881,N_14384);
or U16478 (N_16478,N_12711,N_12220);
and U16479 (N_16479,N_10917,N_12151);
nor U16480 (N_16480,N_11342,N_13017);
nand U16481 (N_16481,N_14107,N_13386);
or U16482 (N_16482,N_14382,N_10066);
or U16483 (N_16483,N_10911,N_13101);
and U16484 (N_16484,N_12358,N_14192);
or U16485 (N_16485,N_10518,N_10117);
and U16486 (N_16486,N_12117,N_14594);
nor U16487 (N_16487,N_10100,N_10535);
or U16488 (N_16488,N_13280,N_10969);
and U16489 (N_16489,N_10634,N_10534);
nor U16490 (N_16490,N_10937,N_10732);
and U16491 (N_16491,N_11210,N_10619);
nor U16492 (N_16492,N_11018,N_13948);
or U16493 (N_16493,N_12878,N_10030);
and U16494 (N_16494,N_11025,N_10843);
xnor U16495 (N_16495,N_10367,N_13534);
nor U16496 (N_16496,N_11398,N_10420);
nor U16497 (N_16497,N_13578,N_13127);
nand U16498 (N_16498,N_14122,N_12716);
nor U16499 (N_16499,N_12611,N_13440);
and U16500 (N_16500,N_11674,N_13310);
or U16501 (N_16501,N_14461,N_14884);
and U16502 (N_16502,N_12694,N_10583);
or U16503 (N_16503,N_10656,N_12420);
and U16504 (N_16504,N_10967,N_10073);
and U16505 (N_16505,N_12679,N_14072);
nand U16506 (N_16506,N_12469,N_10924);
and U16507 (N_16507,N_13827,N_14132);
and U16508 (N_16508,N_11999,N_11869);
or U16509 (N_16509,N_10138,N_12436);
or U16510 (N_16510,N_10551,N_11742);
xor U16511 (N_16511,N_11757,N_13144);
and U16512 (N_16512,N_11409,N_11885);
or U16513 (N_16513,N_10001,N_11326);
and U16514 (N_16514,N_12653,N_11357);
nand U16515 (N_16515,N_11196,N_13140);
xor U16516 (N_16516,N_10054,N_11098);
or U16517 (N_16517,N_10757,N_13376);
nand U16518 (N_16518,N_12216,N_10096);
or U16519 (N_16519,N_12743,N_14320);
xnor U16520 (N_16520,N_11116,N_11206);
xnor U16521 (N_16521,N_14313,N_10202);
or U16522 (N_16522,N_13350,N_14710);
xnor U16523 (N_16523,N_11692,N_11849);
xor U16524 (N_16524,N_12200,N_10723);
and U16525 (N_16525,N_11537,N_13804);
nand U16526 (N_16526,N_13691,N_11694);
nor U16527 (N_16527,N_10659,N_13715);
nand U16528 (N_16528,N_14808,N_12180);
or U16529 (N_16529,N_12999,N_11282);
nor U16530 (N_16530,N_11097,N_11401);
nor U16531 (N_16531,N_10308,N_13942);
and U16532 (N_16532,N_11556,N_12435);
and U16533 (N_16533,N_11283,N_14354);
or U16534 (N_16534,N_12250,N_11440);
nand U16535 (N_16535,N_11075,N_12926);
or U16536 (N_16536,N_13323,N_13371);
or U16537 (N_16537,N_12970,N_14065);
nand U16538 (N_16538,N_14383,N_11775);
xor U16539 (N_16539,N_13916,N_13521);
or U16540 (N_16540,N_10514,N_12606);
nand U16541 (N_16541,N_13790,N_14060);
nand U16542 (N_16542,N_10388,N_11231);
and U16543 (N_16543,N_11092,N_10852);
nor U16544 (N_16544,N_13611,N_11257);
or U16545 (N_16545,N_13322,N_13822);
nor U16546 (N_16546,N_14125,N_10280);
or U16547 (N_16547,N_12910,N_14972);
nor U16548 (N_16548,N_10670,N_13111);
or U16549 (N_16549,N_14844,N_11531);
nand U16550 (N_16550,N_13689,N_12973);
nand U16551 (N_16551,N_11385,N_12087);
or U16552 (N_16552,N_13202,N_14843);
or U16553 (N_16553,N_10786,N_11750);
nor U16554 (N_16554,N_14128,N_10015);
and U16555 (N_16555,N_11486,N_10561);
nor U16556 (N_16556,N_13270,N_10605);
or U16557 (N_16557,N_12138,N_13177);
nand U16558 (N_16558,N_11141,N_10472);
or U16559 (N_16559,N_10994,N_12998);
or U16560 (N_16560,N_12348,N_12866);
and U16561 (N_16561,N_11310,N_12343);
and U16562 (N_16562,N_14857,N_11593);
nand U16563 (N_16563,N_11567,N_10647);
or U16564 (N_16564,N_13683,N_12316);
nand U16565 (N_16565,N_13433,N_10033);
nor U16566 (N_16566,N_12960,N_11834);
and U16567 (N_16567,N_14568,N_14978);
and U16568 (N_16568,N_12356,N_11987);
nor U16569 (N_16569,N_12350,N_10807);
or U16570 (N_16570,N_10417,N_13832);
and U16571 (N_16571,N_13307,N_10635);
or U16572 (N_16572,N_13577,N_10883);
nor U16573 (N_16573,N_11856,N_12045);
or U16574 (N_16574,N_14240,N_13900);
and U16575 (N_16575,N_11632,N_13185);
nand U16576 (N_16576,N_12231,N_12402);
nand U16577 (N_16577,N_12512,N_12080);
or U16578 (N_16578,N_10878,N_13491);
nor U16579 (N_16579,N_13109,N_10660);
nor U16580 (N_16580,N_11813,N_13771);
nor U16581 (N_16581,N_12909,N_10075);
nor U16582 (N_16582,N_13134,N_11608);
and U16583 (N_16583,N_13981,N_12693);
or U16584 (N_16584,N_10841,N_10842);
nand U16585 (N_16585,N_10106,N_11979);
or U16586 (N_16586,N_13748,N_10153);
nor U16587 (N_16587,N_12953,N_11756);
nor U16588 (N_16588,N_13074,N_11164);
nand U16589 (N_16589,N_13843,N_13928);
and U16590 (N_16590,N_11109,N_14761);
nand U16591 (N_16591,N_10349,N_11606);
or U16592 (N_16592,N_12609,N_13705);
nor U16593 (N_16593,N_10745,N_14036);
nor U16594 (N_16594,N_13668,N_13259);
and U16595 (N_16595,N_13023,N_11751);
nor U16596 (N_16596,N_10997,N_12834);
or U16597 (N_16597,N_12879,N_13879);
xnor U16598 (N_16598,N_10720,N_13654);
and U16599 (N_16599,N_12531,N_11812);
and U16600 (N_16600,N_10291,N_11132);
or U16601 (N_16601,N_10487,N_11489);
xnor U16602 (N_16602,N_14949,N_13791);
xor U16603 (N_16603,N_13312,N_11700);
or U16604 (N_16604,N_13862,N_12950);
and U16605 (N_16605,N_11402,N_11189);
xor U16606 (N_16606,N_13008,N_13143);
or U16607 (N_16607,N_10201,N_11432);
nand U16608 (N_16608,N_11888,N_10875);
and U16609 (N_16609,N_14573,N_10567);
nand U16610 (N_16610,N_13692,N_11582);
or U16611 (N_16611,N_11026,N_11982);
nand U16612 (N_16612,N_10548,N_11295);
nor U16613 (N_16613,N_12490,N_13247);
nand U16614 (N_16614,N_14043,N_14750);
xor U16615 (N_16615,N_11697,N_11779);
or U16616 (N_16616,N_10043,N_14947);
and U16617 (N_16617,N_12536,N_11896);
nor U16618 (N_16618,N_14309,N_11368);
nor U16619 (N_16619,N_14684,N_14101);
or U16620 (N_16620,N_12315,N_14302);
nand U16621 (N_16621,N_10413,N_13075);
and U16622 (N_16622,N_13749,N_13062);
or U16623 (N_16623,N_14098,N_14755);
nand U16624 (N_16624,N_11350,N_11600);
xnor U16625 (N_16625,N_11139,N_14784);
nand U16626 (N_16626,N_12202,N_11457);
nor U16627 (N_16627,N_12935,N_14923);
and U16628 (N_16628,N_12028,N_13724);
nand U16629 (N_16629,N_10345,N_12974);
nor U16630 (N_16630,N_10239,N_13422);
and U16631 (N_16631,N_13391,N_12340);
xor U16632 (N_16632,N_12791,N_12401);
or U16633 (N_16633,N_11580,N_12141);
or U16634 (N_16634,N_12175,N_14557);
nor U16635 (N_16635,N_12494,N_14919);
nand U16636 (N_16636,N_10268,N_11484);
nand U16637 (N_16637,N_13321,N_10556);
or U16638 (N_16638,N_14290,N_11880);
or U16639 (N_16639,N_10501,N_10758);
nand U16640 (N_16640,N_12182,N_10351);
and U16641 (N_16641,N_12153,N_14083);
or U16642 (N_16642,N_12562,N_14006);
or U16643 (N_16643,N_14891,N_14986);
and U16644 (N_16644,N_13262,N_14519);
xnor U16645 (N_16645,N_13026,N_13389);
or U16646 (N_16646,N_14672,N_14106);
nand U16647 (N_16647,N_10568,N_12088);
or U16648 (N_16648,N_13477,N_14190);
nor U16649 (N_16649,N_10423,N_14000);
nor U16650 (N_16650,N_12031,N_10697);
or U16651 (N_16651,N_13977,N_12781);
or U16652 (N_16652,N_14040,N_14646);
nor U16653 (N_16653,N_13113,N_10503);
xnor U16654 (N_16654,N_13252,N_14722);
and U16655 (N_16655,N_14254,N_14957);
nand U16656 (N_16656,N_13739,N_11384);
nor U16657 (N_16657,N_14976,N_14390);
and U16658 (N_16658,N_12155,N_12857);
or U16659 (N_16659,N_11449,N_12312);
and U16660 (N_16660,N_11093,N_13079);
nand U16661 (N_16661,N_13883,N_13170);
or U16662 (N_16662,N_12755,N_11289);
or U16663 (N_16663,N_12072,N_14140);
or U16664 (N_16664,N_12115,N_10173);
nand U16665 (N_16665,N_14219,N_11115);
and U16666 (N_16666,N_14039,N_10594);
and U16667 (N_16667,N_12266,N_13731);
nor U16668 (N_16668,N_12396,N_12751);
xnor U16669 (N_16669,N_12475,N_11084);
and U16670 (N_16670,N_10031,N_12882);
or U16671 (N_16671,N_10628,N_13728);
nand U16672 (N_16672,N_13709,N_11040);
or U16673 (N_16673,N_10552,N_12621);
and U16674 (N_16674,N_13738,N_14216);
nand U16675 (N_16675,N_10596,N_11765);
nand U16676 (N_16676,N_10547,N_11467);
xnor U16677 (N_16677,N_13988,N_13858);
and U16678 (N_16678,N_10802,N_10152);
and U16679 (N_16679,N_10405,N_10004);
and U16680 (N_16680,N_14661,N_12456);
and U16681 (N_16681,N_11450,N_10296);
and U16682 (N_16682,N_10667,N_14221);
or U16683 (N_16683,N_11311,N_14480);
or U16684 (N_16684,N_11613,N_11107);
and U16685 (N_16685,N_11452,N_11324);
xnor U16686 (N_16686,N_13594,N_10210);
nor U16687 (N_16687,N_10933,N_12684);
nor U16688 (N_16688,N_10464,N_10877);
nand U16689 (N_16689,N_14311,N_10742);
nand U16690 (N_16690,N_10498,N_12927);
and U16691 (N_16691,N_11162,N_10053);
and U16692 (N_16692,N_14675,N_10226);
nor U16693 (N_16693,N_14341,N_12296);
and U16694 (N_16694,N_13973,N_11752);
or U16695 (N_16695,N_14156,N_14847);
and U16696 (N_16696,N_12589,N_10363);
and U16697 (N_16697,N_10012,N_11890);
xor U16698 (N_16698,N_11811,N_14535);
or U16699 (N_16699,N_14410,N_10398);
xor U16700 (N_16700,N_13072,N_13466);
nand U16701 (N_16701,N_12618,N_10385);
and U16702 (N_16702,N_12601,N_13276);
nand U16703 (N_16703,N_10140,N_10072);
nor U16704 (N_16704,N_10036,N_13096);
or U16705 (N_16705,N_13064,N_12256);
and U16706 (N_16706,N_14775,N_11269);
or U16707 (N_16707,N_13475,N_12534);
nand U16708 (N_16708,N_13579,N_14388);
and U16709 (N_16709,N_10261,N_13909);
or U16710 (N_16710,N_13078,N_11383);
nand U16711 (N_16711,N_10517,N_11318);
xnor U16712 (N_16712,N_14028,N_10976);
or U16713 (N_16713,N_12553,N_10872);
nand U16714 (N_16714,N_12748,N_11922);
nand U16715 (N_16715,N_14513,N_12649);
or U16716 (N_16716,N_12676,N_11598);
nand U16717 (N_16717,N_13313,N_14862);
nand U16718 (N_16718,N_11023,N_11702);
nand U16719 (N_16719,N_11872,N_14208);
and U16720 (N_16720,N_11043,N_14142);
and U16721 (N_16721,N_11148,N_11727);
or U16722 (N_16722,N_14357,N_13557);
or U16723 (N_16723,N_13722,N_11705);
nand U16724 (N_16724,N_11918,N_12201);
or U16725 (N_16725,N_13529,N_11099);
or U16726 (N_16726,N_12624,N_12429);
nor U16727 (N_16727,N_11248,N_10387);
or U16728 (N_16728,N_12384,N_10797);
or U16729 (N_16729,N_10864,N_14886);
nor U16730 (N_16730,N_10780,N_10297);
or U16731 (N_16731,N_10865,N_11762);
nand U16732 (N_16732,N_10716,N_10869);
nand U16733 (N_16733,N_10424,N_12478);
nor U16734 (N_16734,N_12047,N_13537);
and U16735 (N_16735,N_11791,N_11766);
or U16736 (N_16736,N_13582,N_12403);
nand U16737 (N_16737,N_12773,N_10104);
and U16738 (N_16738,N_14450,N_13086);
nand U16739 (N_16739,N_12842,N_11187);
and U16740 (N_16740,N_10231,N_14308);
or U16741 (N_16741,N_10426,N_13050);
nor U16742 (N_16742,N_10914,N_12631);
or U16743 (N_16743,N_12838,N_10168);
or U16744 (N_16744,N_11320,N_14900);
and U16745 (N_16745,N_12247,N_11463);
nand U16746 (N_16746,N_10800,N_10191);
nand U16747 (N_16747,N_10836,N_14731);
nor U16748 (N_16748,N_10408,N_13635);
and U16749 (N_16749,N_13658,N_13657);
nor U16750 (N_16750,N_12194,N_10706);
and U16751 (N_16751,N_11607,N_10438);
or U16752 (N_16752,N_12533,N_13710);
nand U16753 (N_16753,N_12754,N_10221);
nand U16754 (N_16754,N_11072,N_10549);
nand U16755 (N_16755,N_10316,N_13157);
nand U16756 (N_16756,N_13845,N_11343);
or U16757 (N_16757,N_13957,N_12339);
and U16758 (N_16758,N_10939,N_12744);
and U16759 (N_16759,N_14464,N_10678);
nand U16760 (N_16760,N_12977,N_14677);
nand U16761 (N_16761,N_12454,N_14283);
xnor U16762 (N_16762,N_11039,N_12029);
and U16763 (N_16763,N_14415,N_11167);
nand U16764 (N_16764,N_11715,N_12050);
xnor U16765 (N_16765,N_10160,N_14069);
nor U16766 (N_16766,N_13439,N_11539);
or U16767 (N_16767,N_11345,N_14038);
and U16768 (N_16768,N_12712,N_12546);
or U16769 (N_16769,N_12305,N_11725);
nor U16770 (N_16770,N_14229,N_11052);
or U16771 (N_16771,N_12975,N_11579);
nand U16772 (N_16772,N_12875,N_11507);
nand U16773 (N_16773,N_12862,N_14345);
nor U16774 (N_16774,N_12583,N_13168);
nor U16775 (N_16775,N_10655,N_14926);
or U16776 (N_16776,N_10909,N_14498);
nor U16777 (N_16777,N_14181,N_13994);
xnor U16778 (N_16778,N_13509,N_10522);
or U16779 (N_16779,N_11676,N_13263);
and U16780 (N_16780,N_13894,N_11861);
or U16781 (N_16781,N_13975,N_11768);
xnor U16782 (N_16782,N_12570,N_13499);
nand U16783 (N_16783,N_12564,N_10146);
or U16784 (N_16784,N_10729,N_11335);
nand U16785 (N_16785,N_12131,N_12668);
nor U16786 (N_16786,N_10025,N_10764);
nand U16787 (N_16787,N_11871,N_14403);
and U16788 (N_16788,N_12510,N_12229);
nor U16789 (N_16789,N_13450,N_11855);
and U16790 (N_16790,N_11464,N_14033);
and U16791 (N_16791,N_14736,N_13546);
or U16792 (N_16792,N_14616,N_14068);
nand U16793 (N_16793,N_11312,N_12034);
nor U16794 (N_16794,N_12830,N_13545);
and U16795 (N_16795,N_10564,N_11990);
or U16796 (N_16796,N_13458,N_14560);
or U16797 (N_16797,N_13359,N_14184);
xor U16798 (N_16798,N_12613,N_10809);
nor U16799 (N_16799,N_10617,N_14463);
and U16800 (N_16800,N_13951,N_11114);
nand U16801 (N_16801,N_12544,N_10671);
or U16802 (N_16802,N_10452,N_10353);
nor U16803 (N_16803,N_13946,N_10996);
or U16804 (N_16804,N_11223,N_14346);
nand U16805 (N_16805,N_13288,N_10229);
or U16806 (N_16806,N_11829,N_14188);
and U16807 (N_16807,N_14711,N_12775);
or U16808 (N_16808,N_10370,N_12503);
xnor U16809 (N_16809,N_13273,N_12940);
or U16810 (N_16810,N_14994,N_11665);
or U16811 (N_16811,N_13325,N_14865);
nor U16812 (N_16812,N_11331,N_10489);
or U16813 (N_16813,N_11835,N_14432);
nand U16814 (N_16814,N_10095,N_12552);
and U16815 (N_16815,N_10530,N_10235);
nand U16816 (N_16816,N_13887,N_10094);
or U16817 (N_16817,N_14929,N_11989);
nand U16818 (N_16818,N_11038,N_14213);
nand U16819 (N_16819,N_12090,N_11736);
and U16820 (N_16820,N_14948,N_12943);
nand U16821 (N_16821,N_12457,N_11909);
and U16822 (N_16822,N_13525,N_11658);
nor U16823 (N_16823,N_11163,N_10844);
or U16824 (N_16824,N_10870,N_11747);
nand U16825 (N_16825,N_10845,N_13543);
or U16826 (N_16826,N_14502,N_13512);
xor U16827 (N_16827,N_13449,N_14218);
and U16828 (N_16828,N_12692,N_11787);
or U16829 (N_16829,N_11420,N_12065);
nand U16830 (N_16830,N_11149,N_10555);
or U16831 (N_16831,N_12099,N_11101);
nor U16832 (N_16832,N_13493,N_12920);
and U16833 (N_16833,N_14203,N_14838);
nand U16834 (N_16834,N_14610,N_12873);
and U16835 (N_16835,N_11877,N_11494);
and U16836 (N_16836,N_12896,N_10338);
and U16837 (N_16837,N_11287,N_10314);
and U16838 (N_16838,N_12709,N_12867);
nand U16839 (N_16839,N_12721,N_13296);
and U16840 (N_16840,N_13485,N_11036);
nor U16841 (N_16841,N_10365,N_12845);
and U16842 (N_16842,N_11046,N_13217);
or U16843 (N_16843,N_14944,N_13670);
nand U16844 (N_16844,N_11497,N_12279);
and U16845 (N_16845,N_13621,N_11062);
nand U16846 (N_16846,N_12767,N_12538);
nand U16847 (N_16847,N_13590,N_12577);
nor U16848 (N_16848,N_10585,N_12988);
and U16849 (N_16849,N_13077,N_10862);
nand U16850 (N_16850,N_11421,N_11866);
nand U16851 (N_16851,N_11200,N_13633);
and U16852 (N_16852,N_14826,N_12593);
nor U16853 (N_16853,N_13047,N_13438);
and U16854 (N_16854,N_13352,N_13836);
nor U16855 (N_16855,N_11158,N_11549);
nand U16856 (N_16856,N_13991,N_13688);
and U16857 (N_16857,N_13627,N_13886);
and U16858 (N_16858,N_12527,N_12413);
nand U16859 (N_16859,N_10825,N_11501);
nand U16860 (N_16860,N_10818,N_11926);
or U16861 (N_16861,N_12056,N_10181);
xor U16862 (N_16862,N_13303,N_13504);
and U16863 (N_16863,N_12602,N_14327);
nand U16864 (N_16864,N_12400,N_12719);
and U16865 (N_16865,N_12036,N_11633);
xnor U16866 (N_16866,N_11395,N_14975);
or U16867 (N_16867,N_13265,N_11851);
and U16868 (N_16868,N_10557,N_12567);
and U16869 (N_16869,N_13918,N_14118);
or U16870 (N_16870,N_12734,N_10225);
nand U16871 (N_16871,N_13130,N_12095);
nand U16872 (N_16872,N_11636,N_13369);
nand U16873 (N_16873,N_12021,N_11212);
nand U16874 (N_16874,N_12513,N_14506);
and U16875 (N_16875,N_13100,N_14169);
or U16876 (N_16876,N_11488,N_11336);
or U16877 (N_16877,N_13741,N_14163);
and U16878 (N_16878,N_12417,N_12105);
xnor U16879 (N_16879,N_13066,N_13379);
and U16880 (N_16880,N_13599,N_12600);
nand U16881 (N_16881,N_11541,N_10688);
nor U16882 (N_16882,N_11177,N_11792);
nand U16883 (N_16883,N_14088,N_11611);
nand U16884 (N_16884,N_12696,N_13063);
or U16885 (N_16885,N_12246,N_14395);
xnor U16886 (N_16886,N_10029,N_14371);
nor U16887 (N_16887,N_12486,N_12491);
nand U16888 (N_16888,N_13609,N_13503);
or U16889 (N_16889,N_12269,N_12708);
or U16890 (N_16890,N_10989,N_10410);
or U16891 (N_16891,N_12132,N_12253);
and U16892 (N_16892,N_11859,N_12916);
nor U16893 (N_16893,N_13197,N_10213);
and U16894 (N_16894,N_14224,N_13947);
and U16895 (N_16895,N_14936,N_13569);
or U16896 (N_16896,N_13976,N_11286);
xor U16897 (N_16897,N_12023,N_10329);
xor U16898 (N_16898,N_11397,N_11379);
xnor U16899 (N_16899,N_14200,N_11788);
xor U16900 (N_16900,N_11933,N_10482);
and U16901 (N_16901,N_14837,N_12051);
or U16902 (N_16902,N_14100,N_11478);
and U16903 (N_16903,N_12177,N_12173);
nor U16904 (N_16904,N_12596,N_14641);
nand U16905 (N_16905,N_14916,N_11586);
or U16906 (N_16906,N_12858,N_10604);
or U16907 (N_16907,N_11521,N_10750);
and U16908 (N_16908,N_10182,N_13035);
nor U16909 (N_16909,N_12750,N_12492);
nand U16910 (N_16910,N_13319,N_10369);
nand U16911 (N_16911,N_12424,N_14627);
nand U16912 (N_16912,N_12864,N_10215);
and U16913 (N_16913,N_12288,N_11337);
nor U16914 (N_16914,N_10500,N_12407);
and U16915 (N_16915,N_10124,N_12806);
or U16916 (N_16916,N_13799,N_11997);
nand U16917 (N_16917,N_14876,N_11865);
and U16918 (N_16918,N_13914,N_10384);
nor U16919 (N_16919,N_11466,N_14821);
nand U16920 (N_16920,N_14452,N_11382);
nand U16921 (N_16921,N_11552,N_14689);
nand U16922 (N_16922,N_13852,N_12163);
nor U16923 (N_16923,N_12969,N_10711);
or U16924 (N_16924,N_12549,N_11540);
nand U16925 (N_16925,N_12190,N_13712);
nor U16926 (N_16926,N_11408,N_10246);
nand U16927 (N_16927,N_10545,N_12329);
or U16928 (N_16928,N_14518,N_12645);
or U16929 (N_16929,N_14644,N_12479);
and U16930 (N_16930,N_11386,N_13875);
nand U16931 (N_16931,N_12505,N_13410);
or U16932 (N_16932,N_10196,N_14436);
nand U16933 (N_16933,N_10620,N_14423);
nand U16934 (N_16934,N_12639,N_13756);
nor U16935 (N_16935,N_14211,N_12837);
or U16936 (N_16936,N_14365,N_14201);
nand U16937 (N_16937,N_10362,N_12446);
nand U16938 (N_16938,N_11946,N_12126);
and U16939 (N_16939,N_10650,N_12472);
nor U16940 (N_16940,N_10084,N_12468);
and U16941 (N_16941,N_11645,N_10728);
nor U16942 (N_16942,N_10598,N_11142);
or U16943 (N_16943,N_10065,N_10804);
and U16944 (N_16944,N_13733,N_13798);
or U16945 (N_16945,N_13412,N_11846);
or U16946 (N_16946,N_12150,N_11847);
nor U16947 (N_16947,N_12922,N_11905);
nand U16948 (N_16948,N_11749,N_13511);
and U16949 (N_16949,N_12913,N_12025);
and U16950 (N_16950,N_11437,N_13613);
xor U16951 (N_16951,N_14243,N_10249);
nand U16952 (N_16952,N_11983,N_10507);
and U16953 (N_16953,N_12703,N_13430);
and U16954 (N_16954,N_11627,N_10265);
or U16955 (N_16955,N_13281,N_12914);
and U16956 (N_16956,N_14440,N_10673);
and U16957 (N_16957,N_13723,N_11277);
and U16958 (N_16958,N_12993,N_13955);
or U16959 (N_16959,N_12251,N_13415);
nor U16960 (N_16960,N_11980,N_13725);
xor U16961 (N_16961,N_14047,N_12297);
and U16962 (N_16962,N_11577,N_11444);
xnor U16963 (N_16963,N_11021,N_14858);
nor U16964 (N_16964,N_10089,N_14373);
or U16965 (N_16965,N_13742,N_11112);
or U16966 (N_16966,N_13200,N_13794);
nand U16967 (N_16967,N_12689,N_11774);
nor U16968 (N_16968,N_11346,N_12525);
and U16969 (N_16969,N_14592,N_13784);
nor U16970 (N_16970,N_12193,N_14364);
xor U16971 (N_16971,N_12102,N_14980);
or U16972 (N_16972,N_10130,N_14119);
and U16973 (N_16973,N_13447,N_12282);
or U16974 (N_16974,N_10057,N_13486);
nand U16975 (N_16975,N_12554,N_12923);
nor U16976 (N_16976,N_11904,N_14562);
nor U16977 (N_16977,N_12886,N_13751);
or U16978 (N_16978,N_11175,N_10676);
and U16979 (N_16979,N_12058,N_12043);
nand U16980 (N_16980,N_10135,N_10102);
nor U16981 (N_16981,N_14693,N_10377);
nand U16982 (N_16982,N_13823,N_14299);
nand U16983 (N_16983,N_13186,N_13970);
nand U16984 (N_16984,N_12852,N_13917);
or U16985 (N_16985,N_12516,N_14225);
nor U16986 (N_16986,N_12352,N_13139);
nand U16987 (N_16987,N_14524,N_13704);
nand U16988 (N_16988,N_14806,N_10236);
and U16989 (N_16989,N_10779,N_11003);
and U16990 (N_16990,N_12439,N_14709);
xnor U16991 (N_16991,N_12027,N_12204);
nand U16992 (N_16992,N_13029,N_10348);
nor U16993 (N_16993,N_14807,N_12071);
nor U16994 (N_16994,N_12386,N_11298);
nand U16995 (N_16995,N_13549,N_10558);
xor U16996 (N_16996,N_12946,N_13954);
or U16997 (N_16997,N_11461,N_11753);
or U16998 (N_16998,N_14840,N_13754);
nand U16999 (N_16999,N_10460,N_13114);
or U17000 (N_17000,N_11505,N_14633);
or U17001 (N_17001,N_10923,N_13697);
and U17002 (N_17002,N_13716,N_13663);
nand U17003 (N_17003,N_13085,N_11760);
nor U17004 (N_17004,N_11968,N_13573);
or U17005 (N_17005,N_10038,N_12578);
or U17006 (N_17006,N_14620,N_13375);
nor U17007 (N_17007,N_11242,N_12989);
and U17008 (N_17008,N_11334,N_11930);
nand U17009 (N_17009,N_12093,N_13036);
nor U17010 (N_17010,N_10727,N_13076);
nor U17011 (N_17011,N_10080,N_10645);
and U17012 (N_17012,N_14928,N_10465);
and U17013 (N_17013,N_10814,N_14998);
or U17014 (N_17014,N_13353,N_12037);
or U17015 (N_17015,N_13305,N_11369);
nand U17016 (N_17016,N_10449,N_10752);
nand U17017 (N_17017,N_14332,N_12038);
or U17018 (N_17018,N_10925,N_10759);
nand U17019 (N_17019,N_14577,N_10198);
and U17020 (N_17020,N_14145,N_11509);
nor U17021 (N_17021,N_12728,N_10504);
and U17022 (N_17022,N_11942,N_12464);
and U17023 (N_17023,N_11008,N_10529);
and U17024 (N_17024,N_10154,N_11991);
and U17025 (N_17025,N_10357,N_10827);
nand U17026 (N_17026,N_11253,N_14690);
or U17027 (N_17027,N_11689,N_11262);
nor U17028 (N_17028,N_10570,N_14097);
nand U17029 (N_17029,N_12898,N_11937);
or U17030 (N_17030,N_10325,N_14301);
nand U17031 (N_17031,N_10003,N_13024);
or U17032 (N_17032,N_12733,N_12906);
nor U17033 (N_17033,N_10055,N_12683);
nor U17034 (N_17034,N_11706,N_11234);
xnor U17035 (N_17035,N_10371,N_14334);
and U17036 (N_17036,N_12020,N_13922);
and U17037 (N_17037,N_12178,N_14908);
or U17038 (N_17038,N_11462,N_11952);
xnor U17039 (N_17039,N_12281,N_12055);
and U17040 (N_17040,N_14159,N_10230);
nand U17041 (N_17041,N_10796,N_14740);
and U17042 (N_17042,N_14846,N_10266);
nor U17043 (N_17043,N_14835,N_11651);
nor U17044 (N_17044,N_12790,N_11620);
and U17045 (N_17045,N_14455,N_13824);
xor U17046 (N_17046,N_11330,N_14652);
and U17047 (N_17047,N_13392,N_11927);
nand U17048 (N_17048,N_10543,N_11213);
nand U17049 (N_17049,N_14607,N_10838);
and U17050 (N_17050,N_10110,N_11503);
nand U17051 (N_17051,N_13847,N_10005);
and U17052 (N_17052,N_10459,N_11012);
and U17053 (N_17053,N_14797,N_12860);
and U17054 (N_17054,N_12856,N_12049);
nor U17055 (N_17055,N_14636,N_10466);
nand U17056 (N_17056,N_13673,N_11864);
nand U17057 (N_17057,N_11031,N_11912);
nor U17058 (N_17058,N_10008,N_14041);
or U17059 (N_17059,N_12224,N_14817);
or U17060 (N_17060,N_12532,N_14237);
nor U17061 (N_17061,N_14544,N_12588);
xnor U17062 (N_17062,N_13974,N_12892);
nor U17063 (N_17063,N_10381,N_12176);
or U17064 (N_17064,N_10174,N_11082);
or U17065 (N_17065,N_14433,N_13426);
nor U17066 (N_17066,N_13753,N_10350);
or U17067 (N_17067,N_10794,N_13684);
nand U17068 (N_17068,N_12259,N_11928);
and U17069 (N_17069,N_10707,N_12292);
nand U17070 (N_17070,N_10092,N_14953);
or U17071 (N_17071,N_12701,N_11534);
nand U17072 (N_17072,N_12154,N_14419);
and U17073 (N_17073,N_10719,N_14195);
nor U17074 (N_17074,N_10415,N_13190);
nor U17075 (N_17075,N_12594,N_11810);
or U17076 (N_17076,N_13536,N_13912);
nand U17077 (N_17077,N_10609,N_14702);
nor U17078 (N_17078,N_13110,N_13564);
and U17079 (N_17079,N_11247,N_14581);
and U17080 (N_17080,N_11339,N_13856);
and U17081 (N_17081,N_10856,N_10801);
nand U17082 (N_17082,N_11617,N_11050);
nand U17083 (N_17083,N_14375,N_14542);
and U17084 (N_17084,N_12964,N_14150);
and U17085 (N_17085,N_14476,N_11239);
nand U17086 (N_17086,N_13295,N_10121);
nand U17087 (N_17087,N_12120,N_11686);
xnor U17088 (N_17088,N_13112,N_10737);
xor U17089 (N_17089,N_10219,N_12770);
nand U17090 (N_17090,N_14753,N_13768);
or U17091 (N_17091,N_13773,N_12442);
and U17092 (N_17092,N_14470,N_13841);
nor U17093 (N_17093,N_13766,N_12984);
nand U17094 (N_17094,N_11394,N_11931);
and U17095 (N_17095,N_11915,N_11267);
nor U17096 (N_17096,N_14048,N_11884);
nor U17097 (N_17097,N_13494,N_13173);
nor U17098 (N_17098,N_11044,N_14212);
nand U17099 (N_17099,N_14658,N_11077);
nor U17100 (N_17100,N_14904,N_10854);
xnor U17101 (N_17101,N_11011,N_11197);
nor U17102 (N_17102,N_11596,N_12575);
nand U17103 (N_17103,N_10916,N_12293);
xnor U17104 (N_17104,N_12628,N_13328);
and U17105 (N_17105,N_14185,N_10252);
nor U17106 (N_17106,N_13903,N_11341);
and U17107 (N_17107,N_12378,N_11291);
and U17108 (N_17108,N_12737,N_10077);
nor U17109 (N_17109,N_10002,N_10234);
or U17110 (N_17110,N_14396,N_10127);
and U17111 (N_17111,N_14752,N_13859);
nor U17112 (N_17112,N_14367,N_12833);
nand U17113 (N_17113,N_13867,N_11010);
xnor U17114 (N_17114,N_14556,N_12110);
or U17115 (N_17115,N_12941,N_10573);
or U17116 (N_17116,N_14892,N_10258);
nor U17117 (N_17117,N_10321,N_12248);
and U17118 (N_17118,N_10379,N_14393);
or U17119 (N_17119,N_11076,N_12957);
nor U17120 (N_17120,N_11439,N_14056);
and U17121 (N_17121,N_11612,N_14392);
or U17122 (N_17122,N_12005,N_14877);
xnor U17123 (N_17123,N_14724,N_13337);
or U17124 (N_17124,N_13192,N_13407);
and U17125 (N_17125,N_14444,N_12919);
xor U17126 (N_17126,N_10944,N_11622);
nor U17127 (N_17127,N_13995,N_14576);
nor U17128 (N_17128,N_13137,N_13638);
or U17129 (N_17129,N_13660,N_13869);
xnor U17130 (N_17130,N_13937,N_12963);
nor U17131 (N_17131,N_11925,N_11945);
nand U17132 (N_17132,N_10606,N_12801);
nand U17133 (N_17133,N_10211,N_11266);
xnor U17134 (N_17134,N_14777,N_14194);
or U17135 (N_17135,N_12550,N_13702);
and U17136 (N_17136,N_12945,N_11371);
or U17137 (N_17137,N_11523,N_10324);
or U17138 (N_17138,N_11292,N_11479);
and U17139 (N_17139,N_11960,N_11998);
or U17140 (N_17140,N_11638,N_11648);
and U17141 (N_17141,N_10380,N_10250);
nor U17142 (N_17142,N_10953,N_10437);
or U17143 (N_17143,N_11080,N_10430);
nand U17144 (N_17144,N_11961,N_14166);
nand U17145 (N_17145,N_10257,N_13662);
or U17146 (N_17146,N_13128,N_10998);
and U17147 (N_17147,N_13454,N_11100);
and U17148 (N_17148,N_13327,N_11460);
or U17149 (N_17149,N_12640,N_11688);
and U17150 (N_17150,N_14406,N_12641);
and U17151 (N_17151,N_10785,N_14925);
and U17152 (N_17152,N_11955,N_10861);
nand U17153 (N_17153,N_10071,N_11238);
xor U17154 (N_17154,N_14014,N_14328);
xnor U17155 (N_17155,N_12188,N_14238);
and U17156 (N_17156,N_11711,N_12365);
and U17157 (N_17157,N_13707,N_14247);
nor U17158 (N_17158,N_11317,N_11883);
and U17159 (N_17159,N_12467,N_13664);
nand U17160 (N_17160,N_12415,N_10722);
nor U17161 (N_17161,N_10956,N_14584);
nor U17162 (N_17162,N_10490,N_10586);
nor U17163 (N_17163,N_12603,N_10621);
nand U17164 (N_17164,N_13943,N_14793);
and U17165 (N_17165,N_12324,N_13616);
or U17166 (N_17166,N_14685,N_12620);
xor U17167 (N_17167,N_11714,N_11322);
and U17168 (N_17168,N_11041,N_13817);
nand U17169 (N_17169,N_10061,N_10078);
nor U17170 (N_17170,N_11698,N_13084);
nor U17171 (N_17171,N_14619,N_13131);
nand U17172 (N_17172,N_14526,N_14241);
or U17173 (N_17173,N_14708,N_12768);
nor U17174 (N_17174,N_14866,N_13801);
or U17175 (N_17175,N_11258,N_13099);
nor U17176 (N_17176,N_12629,N_11305);
and U17177 (N_17177,N_14148,N_14210);
or U17178 (N_17178,N_12012,N_14574);
nor U17179 (N_17179,N_13677,N_14842);
nor U17180 (N_17180,N_14458,N_14117);
or U17181 (N_17181,N_10223,N_12207);
or U17182 (N_17182,N_10275,N_13165);
nor U17183 (N_17183,N_14350,N_14727);
nand U17184 (N_17184,N_13600,N_11929);
or U17185 (N_17185,N_11841,N_10256);
nor U17186 (N_17186,N_12040,N_13855);
and U17187 (N_17187,N_14745,N_13451);
xnor U17188 (N_17188,N_11308,N_10744);
or U17189 (N_17189,N_11338,N_13193);
nand U17190 (N_17190,N_11794,N_12698);
and U17191 (N_17191,N_13261,N_10612);
nor U17192 (N_17192,N_14205,N_14091);
nor U17193 (N_17193,N_12660,N_13231);
or U17194 (N_17194,N_11712,N_13612);
nand U17195 (N_17195,N_12638,N_14246);
and U17196 (N_17196,N_14180,N_12686);
nand U17197 (N_17197,N_13848,N_10908);
nor U17198 (N_17198,N_12807,N_11433);
xnor U17199 (N_17199,N_14785,N_12054);
or U17200 (N_17200,N_14924,N_12286);
and U17201 (N_17201,N_13698,N_13176);
or U17202 (N_17202,N_10446,N_12363);
nand U17203 (N_17203,N_12612,N_12304);
and U17204 (N_17204,N_10968,N_10958);
and U17205 (N_17205,N_12521,N_14447);
nor U17206 (N_17206,N_14508,N_11891);
or U17207 (N_17207,N_10343,N_11631);
and U17208 (N_17208,N_14045,N_12113);
and U17209 (N_17209,N_13135,N_14597);
nor U17210 (N_17210,N_13842,N_11007);
xor U17211 (N_17211,N_12981,N_14905);
and U17212 (N_17212,N_14174,N_11447);
nand U17213 (N_17213,N_13031,N_13041);
nor U17214 (N_17214,N_14284,N_12765);
or U17215 (N_17215,N_10485,N_12360);
and U17216 (N_17216,N_13978,N_11669);
nand U17217 (N_17217,N_12128,N_11129);
nor U17218 (N_17218,N_12831,N_14291);
nor U17219 (N_17219,N_11285,N_13442);
and U17220 (N_17220,N_12799,N_14249);
nand U17221 (N_17221,N_13505,N_12717);
and U17222 (N_17222,N_11006,N_13797);
or U17223 (N_17223,N_14814,N_11956);
nand U17224 (N_17224,N_14500,N_12024);
or U17225 (N_17225,N_11867,N_11601);
and U17226 (N_17226,N_13105,N_12713);
or U17227 (N_17227,N_11863,N_10763);
nand U17228 (N_17228,N_10709,N_12659);
or U17229 (N_17229,N_13838,N_14788);
nand U17230 (N_17230,N_14287,N_11699);
and U17231 (N_17231,N_12548,N_10772);
nor U17232 (N_17232,N_10147,N_13587);
nand U17233 (N_17233,N_10717,N_10088);
and U17234 (N_17234,N_13338,N_10240);
or U17235 (N_17235,N_14207,N_14094);
nor U17236 (N_17236,N_10636,N_14003);
and U17237 (N_17237,N_13243,N_10278);
nor U17238 (N_17238,N_11416,N_14303);
nor U17239 (N_17239,N_11957,N_13241);
xnor U17240 (N_17240,N_11182,N_12032);
xor U17241 (N_17241,N_13019,N_12136);
nor U17242 (N_17242,N_10981,N_10010);
and U17243 (N_17243,N_14833,N_10954);
or U17244 (N_17244,N_13615,N_11947);
nor U17245 (N_17245,N_11621,N_11704);
xnor U17246 (N_17246,N_14441,N_12753);
and U17247 (N_17247,N_12135,N_13226);
nor U17248 (N_17248,N_11568,N_13332);
nand U17249 (N_17249,N_12035,N_13302);
or U17250 (N_17250,N_12675,N_11412);
nand U17251 (N_17251,N_11780,N_14860);
nor U17252 (N_17252,N_10190,N_12166);
nand U17253 (N_17253,N_11799,N_14565);
nand U17254 (N_17254,N_13812,N_12894);
or U17255 (N_17255,N_12059,N_13871);
nand U17256 (N_17256,N_12211,N_12732);
and U17257 (N_17257,N_10218,N_10502);
nand U17258 (N_17258,N_12127,N_14482);
xor U17259 (N_17259,N_14955,N_13620);
nand U17260 (N_17260,N_12829,N_14883);
and U17261 (N_17261,N_14209,N_12539);
nand U17262 (N_17262,N_11708,N_13222);
and U17263 (N_17263,N_11122,N_13933);
nor U17264 (N_17264,N_13184,N_14330);
or U17265 (N_17265,N_10251,N_14539);
nor U17266 (N_17266,N_13816,N_13777);
and U17267 (N_17267,N_12932,N_14001);
nor U17268 (N_17268,N_10279,N_13092);
or U17269 (N_17269,N_13166,N_14520);
and U17270 (N_17270,N_10108,N_14902);
nand U17271 (N_17271,N_14035,N_11465);
or U17272 (N_17272,N_12899,N_13179);
or U17273 (N_17273,N_14514,N_12473);
or U17274 (N_17274,N_14431,N_14485);
nand U17275 (N_17275,N_12699,N_12859);
and U17276 (N_17276,N_11630,N_13906);
or U17277 (N_17277,N_14177,N_10382);
and U17278 (N_17278,N_13234,N_13825);
nor U17279 (N_17279,N_14804,N_14668);
nor U17280 (N_17280,N_10791,N_14490);
nor U17281 (N_17281,N_11902,N_10208);
and U17282 (N_17282,N_11569,N_14104);
and U17283 (N_17283,N_14650,N_12817);
xnor U17284 (N_17284,N_14861,N_14202);
nor U17285 (N_17285,N_14402,N_11545);
xor U17286 (N_17286,N_14307,N_11995);
xor U17287 (N_17287,N_10319,N_14717);
xor U17288 (N_17288,N_12084,N_13700);
nand U17289 (N_17289,N_10611,N_13576);
and U17290 (N_17290,N_12357,N_13395);
or U17291 (N_17291,N_11246,N_11860);
or U17292 (N_17292,N_13719,N_10754);
nor U17293 (N_17293,N_14718,N_10778);
nand U17294 (N_17294,N_12956,N_14681);
nand U17295 (N_17295,N_13149,N_11559);
or U17296 (N_17296,N_11226,N_14197);
nand U17297 (N_17297,N_10494,N_13082);
nand U17298 (N_17298,N_14525,N_10295);
nand U17299 (N_17299,N_10148,N_13387);
or U17300 (N_17300,N_10128,N_14686);
or U17301 (N_17301,N_11029,N_11288);
and U17302 (N_17302,N_12426,N_14744);
and U17303 (N_17303,N_11992,N_10220);
and U17304 (N_17304,N_11307,N_14491);
or U17305 (N_17305,N_14497,N_10228);
and U17306 (N_17306,N_13877,N_12078);
and U17307 (N_17307,N_10322,N_12947);
nand U17308 (N_17308,N_13336,N_14114);
nor U17309 (N_17309,N_12073,N_14477);
and U17310 (N_17310,N_12794,N_10254);
and U17311 (N_17311,N_14079,N_14765);
nor U17312 (N_17312,N_11661,N_14289);
nor U17313 (N_17313,N_12635,N_12418);
or U17314 (N_17314,N_13547,N_11828);
nor U17315 (N_17315,N_10016,N_14130);
nor U17316 (N_17316,N_12443,N_11570);
or U17317 (N_17317,N_12440,N_12771);
or U17318 (N_17318,N_12107,N_10642);
nor U17319 (N_17319,N_13781,N_14653);
nor U17320 (N_17320,N_13803,N_10344);
and U17321 (N_17321,N_10663,N_12874);
nand U17322 (N_17322,N_12100,N_11778);
or U17323 (N_17323,N_10887,N_14167);
xor U17324 (N_17324,N_12148,N_10971);
and U17325 (N_17325,N_13889,N_10151);
or U17326 (N_17326,N_14732,N_11796);
and U17327 (N_17327,N_14471,N_14070);
xor U17328 (N_17328,N_13366,N_14707);
nand U17329 (N_17329,N_14484,N_10480);
nand U17330 (N_17330,N_14199,N_10921);
or U17331 (N_17331,N_14612,N_13498);
nand U17332 (N_17332,N_14343,N_13558);
and U17333 (N_17333,N_13835,N_10554);
nand U17334 (N_17334,N_12156,N_12033);
or U17335 (N_17335,N_11673,N_11973);
or U17336 (N_17336,N_14849,N_14552);
or U17337 (N_17337,N_13287,N_13038);
and U17338 (N_17338,N_11138,N_10304);
nand U17339 (N_17339,N_12079,N_12715);
and U17340 (N_17340,N_10651,N_11555);
and U17341 (N_17341,N_14973,N_14278);
or U17342 (N_17342,N_14165,N_11894);
nand U17343 (N_17343,N_11030,N_10412);
xor U17344 (N_17344,N_11362,N_14824);
or U17345 (N_17345,N_11746,N_10795);
nand U17346 (N_17346,N_14703,N_13767);
or U17347 (N_17347,N_11609,N_13206);
nor U17348 (N_17348,N_13236,N_13833);
nor U17349 (N_17349,N_10390,N_12616);
or U17350 (N_17350,N_11475,N_10425);
nand U17351 (N_17351,N_10207,N_14488);
xor U17352 (N_17352,N_12769,N_12232);
nor U17353 (N_17353,N_10436,N_10931);
nand U17354 (N_17354,N_11562,N_12068);
nor U17355 (N_17355,N_14271,N_12610);
or U17356 (N_17356,N_11208,N_12648);
nor U17357 (N_17357,N_13996,N_13500);
or U17358 (N_17358,N_10448,N_14832);
nand U17359 (N_17359,N_10848,N_11921);
nand U17360 (N_17360,N_12891,N_10890);
nand U17361 (N_17361,N_11393,N_12907);
or U17362 (N_17362,N_12482,N_10942);
and U17363 (N_17363,N_11354,N_13255);
and U17364 (N_17364,N_13645,N_11133);
or U17365 (N_17365,N_13320,N_14198);
nand U17366 (N_17366,N_14077,N_13080);
nor U17367 (N_17367,N_12514,N_11293);
nand U17368 (N_17368,N_12634,N_14841);
nand U17369 (N_17369,N_11155,N_11789);
or U17370 (N_17370,N_12545,N_10990);
or U17371 (N_17371,N_12725,N_10669);
nand U17372 (N_17372,N_13117,N_10597);
or U17373 (N_17373,N_11222,N_10815);
or U17374 (N_17374,N_12006,N_12267);
nor U17375 (N_17375,N_11067,N_12370);
or U17376 (N_17376,N_12471,N_13559);
and U17377 (N_17377,N_11547,N_11176);
and U17378 (N_17378,N_14189,N_11587);
nor U17379 (N_17379,N_10141,N_13385);
xor U17380 (N_17380,N_13400,N_10330);
nor U17381 (N_17381,N_11544,N_13743);
or U17382 (N_17382,N_10974,N_12520);
or U17383 (N_17383,N_11969,N_10037);
and U17384 (N_17384,N_13548,N_10059);
and U17385 (N_17385,N_13786,N_14457);
or U17386 (N_17386,N_11459,N_13060);
nor U17387 (N_17387,N_11436,N_13317);
nand U17388 (N_17388,N_11134,N_10743);
and U17389 (N_17389,N_14478,N_14275);
or U17390 (N_17390,N_10784,N_13518);
and U17391 (N_17391,N_14789,N_14682);
or U17392 (N_17392,N_14126,N_13810);
or U17393 (N_17393,N_10982,N_12623);
nand U17394 (N_17394,N_13961,N_13098);
or U17395 (N_17395,N_11378,N_10542);
nand U17396 (N_17396,N_10020,N_11218);
xnor U17397 (N_17397,N_12626,N_14911);
nand U17398 (N_17398,N_14226,N_13762);
and U17399 (N_17399,N_14981,N_13283);
or U17400 (N_17400,N_10509,N_13300);
or U17401 (N_17401,N_14082,N_10450);
nor U17402 (N_17402,N_11804,N_11533);
nand U17403 (N_17403,N_14554,N_13103);
nand U17404 (N_17404,N_14671,N_14459);
and U17405 (N_17405,N_12876,N_12483);
and U17406 (N_17406,N_13813,N_12669);
nand U17407 (N_17407,N_11800,N_10114);
xnor U17408 (N_17408,N_12558,N_14087);
nor U17409 (N_17409,N_12169,N_13009);
and U17410 (N_17410,N_10860,N_13256);
nor U17411 (N_17411,N_13298,N_12184);
and U17412 (N_17412,N_14510,N_14590);
and U17413 (N_17413,N_13361,N_10162);
nand U17414 (N_17414,N_13059,N_12405);
and U17415 (N_17415,N_12333,N_11809);
and U17416 (N_17416,N_13513,N_14572);
nand U17417 (N_17417,N_10806,N_10285);
xnor U17418 (N_17418,N_12018,N_14267);
xor U17419 (N_17419,N_10481,N_11681);
and U17420 (N_17420,N_10414,N_13592);
nand U17421 (N_17421,N_12537,N_11422);
nor U17422 (N_17422,N_12081,N_13195);
nand U17423 (N_17423,N_10274,N_14030);
nand U17424 (N_17424,N_10063,N_11616);
nand U17425 (N_17425,N_13238,N_11682);
nand U17426 (N_17426,N_13675,N_13872);
nor U17427 (N_17427,N_14850,N_13294);
nor U17428 (N_17428,N_11773,N_12885);
or U17429 (N_17429,N_12822,N_11205);
xnor U17430 (N_17430,N_13445,N_12646);
nand U17431 (N_17431,N_12263,N_11413);
and U17432 (N_17432,N_11063,N_11900);
or U17433 (N_17433,N_14049,N_14103);
and U17434 (N_17434,N_10085,N_11767);
or U17435 (N_17435,N_14413,N_13213);
nor U17436 (N_17436,N_10587,N_14966);
nand U17437 (N_17437,N_10792,N_14086);
nor U17438 (N_17438,N_14034,N_11434);
and U17439 (N_17439,N_14183,N_14359);
nand U17440 (N_17440,N_11355,N_11214);
or U17441 (N_17441,N_10393,N_14347);
and U17442 (N_17442,N_11783,N_10790);
nor U17443 (N_17443,N_12374,N_14746);
and U17444 (N_17444,N_11564,N_14420);
nand U17445 (N_17445,N_10767,N_13309);
nor U17446 (N_17446,N_12569,N_10850);
xor U17447 (N_17447,N_13306,N_14766);
xor U17448 (N_17448,N_10566,N_12061);
nor U17449 (N_17449,N_11166,N_13142);
nand U17450 (N_17450,N_13538,N_12326);
nand U17451 (N_17451,N_11993,N_13820);
nand U17452 (N_17452,N_12379,N_14725);
and U17453 (N_17453,N_10491,N_13527);
and U17454 (N_17454,N_11380,N_10175);
nor U17455 (N_17455,N_13653,N_13761);
nor U17456 (N_17456,N_13090,N_13934);
nor U17457 (N_17457,N_11273,N_13383);
nand U17458 (N_17458,N_11144,N_10524);
nor U17459 (N_17459,N_10963,N_14399);
or U17460 (N_17460,N_14632,N_12561);
and U17461 (N_17461,N_14738,N_13027);
and U17462 (N_17462,N_13603,N_12779);
nand U17463 (N_17463,N_10427,N_10327);
nand U17464 (N_17464,N_13681,N_13201);
or U17465 (N_17465,N_10788,N_10510);
nor U17466 (N_17466,N_13264,N_12425);
nor U17467 (N_17467,N_14812,N_10735);
or U17468 (N_17468,N_11153,N_14059);
and U17469 (N_17469,N_12244,N_12656);
and U17470 (N_17470,N_14692,N_10397);
or U17471 (N_17471,N_14220,N_13687);
nor U17472 (N_17472,N_14143,N_10335);
and U17473 (N_17473,N_12542,N_11508);
or U17474 (N_17474,N_14479,N_13102);
and U17475 (N_17475,N_13542,N_12140);
nor U17476 (N_17476,N_11755,N_10439);
nor U17477 (N_17477,N_13129,N_13734);
or U17478 (N_17478,N_10980,N_14913);
nand U17479 (N_17479,N_11251,N_10859);
or U17480 (N_17480,N_11373,N_14073);
nor U17481 (N_17481,N_11473,N_12364);
nor U17482 (N_17482,N_13116,N_12123);
and U17483 (N_17483,N_10049,N_11332);
nand U17484 (N_17484,N_11235,N_11161);
nand U17485 (N_17485,N_13585,N_13647);
or U17486 (N_17486,N_12291,N_13821);
nand U17487 (N_17487,N_10853,N_14268);
nor U17488 (N_17488,N_11103,N_11584);
or U17489 (N_17489,N_12826,N_12746);
and U17490 (N_17490,N_12654,N_12565);
or U17491 (N_17491,N_11498,N_14050);
and U17492 (N_17492,N_10411,N_10493);
nand U17493 (N_17493,N_13463,N_13414);
nor U17494 (N_17494,N_10097,N_11316);
or U17495 (N_17495,N_10876,N_12585);
and U17496 (N_17496,N_14244,N_10813);
nor U17497 (N_17497,N_14779,N_12121);
or U17498 (N_17498,N_13054,N_14439);
or U17499 (N_17499,N_12349,N_11106);
nor U17500 (N_17500,N_13901,N_11012);
xnor U17501 (N_17501,N_13561,N_13418);
or U17502 (N_17502,N_12398,N_11165);
and U17503 (N_17503,N_13080,N_10272);
nor U17504 (N_17504,N_13925,N_13555);
nor U17505 (N_17505,N_10416,N_14816);
nor U17506 (N_17506,N_14202,N_14797);
or U17507 (N_17507,N_12886,N_11748);
and U17508 (N_17508,N_14488,N_14082);
nor U17509 (N_17509,N_13261,N_10794);
nor U17510 (N_17510,N_10611,N_14213);
nand U17511 (N_17511,N_10551,N_13981);
and U17512 (N_17512,N_11356,N_13015);
nand U17513 (N_17513,N_11130,N_13488);
nand U17514 (N_17514,N_12890,N_12861);
nor U17515 (N_17515,N_14519,N_11979);
xor U17516 (N_17516,N_12773,N_13154);
and U17517 (N_17517,N_11698,N_14585);
or U17518 (N_17518,N_11644,N_13478);
and U17519 (N_17519,N_10355,N_11649);
and U17520 (N_17520,N_13567,N_12122);
or U17521 (N_17521,N_13371,N_13918);
and U17522 (N_17522,N_11004,N_13709);
nor U17523 (N_17523,N_14429,N_12979);
and U17524 (N_17524,N_10130,N_12821);
or U17525 (N_17525,N_12391,N_11865);
and U17526 (N_17526,N_14053,N_12666);
nand U17527 (N_17527,N_12341,N_11021);
nor U17528 (N_17528,N_10208,N_13120);
and U17529 (N_17529,N_13599,N_11874);
nor U17530 (N_17530,N_11125,N_12112);
and U17531 (N_17531,N_11802,N_10921);
xnor U17532 (N_17532,N_13572,N_11849);
nand U17533 (N_17533,N_13488,N_13175);
and U17534 (N_17534,N_13409,N_13908);
nand U17535 (N_17535,N_11228,N_10545);
or U17536 (N_17536,N_10115,N_13770);
or U17537 (N_17537,N_13470,N_11957);
nand U17538 (N_17538,N_14796,N_12701);
nand U17539 (N_17539,N_14016,N_13653);
nand U17540 (N_17540,N_10368,N_13874);
nand U17541 (N_17541,N_14732,N_12050);
nand U17542 (N_17542,N_12714,N_13894);
nand U17543 (N_17543,N_10620,N_12017);
or U17544 (N_17544,N_13608,N_12607);
or U17545 (N_17545,N_14929,N_11267);
nand U17546 (N_17546,N_14050,N_10890);
or U17547 (N_17547,N_10539,N_13506);
or U17548 (N_17548,N_12191,N_11840);
and U17549 (N_17549,N_10586,N_12392);
xor U17550 (N_17550,N_11423,N_14521);
nand U17551 (N_17551,N_13547,N_10540);
xor U17552 (N_17552,N_14279,N_13015);
nand U17553 (N_17553,N_10512,N_12908);
and U17554 (N_17554,N_12391,N_11143);
and U17555 (N_17555,N_13055,N_14770);
nor U17556 (N_17556,N_12956,N_11678);
or U17557 (N_17557,N_12936,N_14237);
or U17558 (N_17558,N_10703,N_12482);
nor U17559 (N_17559,N_11244,N_12828);
or U17560 (N_17560,N_10724,N_10066);
nand U17561 (N_17561,N_11961,N_14732);
or U17562 (N_17562,N_12829,N_12739);
nor U17563 (N_17563,N_10888,N_10022);
nor U17564 (N_17564,N_12320,N_11768);
nor U17565 (N_17565,N_10450,N_12986);
and U17566 (N_17566,N_14383,N_13864);
xor U17567 (N_17567,N_10815,N_13331);
nand U17568 (N_17568,N_13830,N_11444);
nand U17569 (N_17569,N_14616,N_12818);
nand U17570 (N_17570,N_11598,N_14630);
or U17571 (N_17571,N_11195,N_12461);
nor U17572 (N_17572,N_14815,N_13716);
nor U17573 (N_17573,N_14453,N_12720);
nor U17574 (N_17574,N_14673,N_11075);
and U17575 (N_17575,N_10640,N_13189);
and U17576 (N_17576,N_11359,N_11834);
and U17577 (N_17577,N_10306,N_13770);
nor U17578 (N_17578,N_14660,N_10146);
xor U17579 (N_17579,N_13568,N_11712);
nor U17580 (N_17580,N_10719,N_14890);
and U17581 (N_17581,N_11655,N_13096);
and U17582 (N_17582,N_11825,N_10090);
nor U17583 (N_17583,N_13144,N_12587);
nand U17584 (N_17584,N_11083,N_12945);
nor U17585 (N_17585,N_14870,N_11390);
and U17586 (N_17586,N_12055,N_13138);
nand U17587 (N_17587,N_13699,N_12458);
or U17588 (N_17588,N_12865,N_12062);
and U17589 (N_17589,N_10855,N_14331);
and U17590 (N_17590,N_13209,N_13233);
nor U17591 (N_17591,N_13628,N_11190);
nand U17592 (N_17592,N_11482,N_14059);
and U17593 (N_17593,N_12896,N_10232);
nor U17594 (N_17594,N_14065,N_14506);
nor U17595 (N_17595,N_14809,N_12064);
or U17596 (N_17596,N_13012,N_13427);
xnor U17597 (N_17597,N_10838,N_11952);
nor U17598 (N_17598,N_13796,N_10853);
nor U17599 (N_17599,N_11496,N_13319);
nand U17600 (N_17600,N_12346,N_12999);
nand U17601 (N_17601,N_14375,N_13491);
or U17602 (N_17602,N_10437,N_11668);
and U17603 (N_17603,N_11593,N_14132);
and U17604 (N_17604,N_14315,N_14875);
and U17605 (N_17605,N_13649,N_11461);
or U17606 (N_17606,N_11573,N_11161);
or U17607 (N_17607,N_10666,N_11949);
xnor U17608 (N_17608,N_11715,N_14949);
nand U17609 (N_17609,N_13156,N_14905);
and U17610 (N_17610,N_12562,N_14293);
or U17611 (N_17611,N_14400,N_12399);
nand U17612 (N_17612,N_13260,N_10805);
xnor U17613 (N_17613,N_12621,N_10696);
xor U17614 (N_17614,N_10137,N_13065);
nor U17615 (N_17615,N_11393,N_13431);
xnor U17616 (N_17616,N_11797,N_10160);
and U17617 (N_17617,N_14886,N_13280);
or U17618 (N_17618,N_10056,N_12813);
nor U17619 (N_17619,N_14609,N_11797);
or U17620 (N_17620,N_14608,N_10480);
or U17621 (N_17621,N_14796,N_12605);
nand U17622 (N_17622,N_14867,N_12904);
nor U17623 (N_17623,N_11641,N_11691);
nand U17624 (N_17624,N_10351,N_14117);
or U17625 (N_17625,N_13167,N_11802);
and U17626 (N_17626,N_13668,N_12096);
nor U17627 (N_17627,N_13600,N_14981);
nand U17628 (N_17628,N_11650,N_13059);
nand U17629 (N_17629,N_13993,N_10310);
and U17630 (N_17630,N_11665,N_12506);
xor U17631 (N_17631,N_12404,N_10378);
nand U17632 (N_17632,N_13476,N_13364);
xor U17633 (N_17633,N_14300,N_13915);
or U17634 (N_17634,N_10192,N_14410);
nor U17635 (N_17635,N_14444,N_10172);
nor U17636 (N_17636,N_14658,N_12759);
or U17637 (N_17637,N_11752,N_14581);
xor U17638 (N_17638,N_11103,N_13633);
nand U17639 (N_17639,N_11342,N_11385);
or U17640 (N_17640,N_13094,N_10123);
and U17641 (N_17641,N_13697,N_14652);
or U17642 (N_17642,N_13156,N_11705);
or U17643 (N_17643,N_14915,N_12264);
xnor U17644 (N_17644,N_11804,N_11108);
or U17645 (N_17645,N_13737,N_13260);
nor U17646 (N_17646,N_12152,N_13373);
or U17647 (N_17647,N_12478,N_11832);
and U17648 (N_17648,N_14701,N_10863);
xor U17649 (N_17649,N_13224,N_12245);
and U17650 (N_17650,N_11670,N_12933);
and U17651 (N_17651,N_10441,N_14305);
or U17652 (N_17652,N_12252,N_11717);
or U17653 (N_17653,N_13634,N_13812);
nor U17654 (N_17654,N_11687,N_10802);
and U17655 (N_17655,N_11790,N_13936);
and U17656 (N_17656,N_10216,N_12371);
and U17657 (N_17657,N_12039,N_13217);
xor U17658 (N_17658,N_13144,N_11160);
or U17659 (N_17659,N_12287,N_10096);
nand U17660 (N_17660,N_10774,N_12872);
and U17661 (N_17661,N_14744,N_13727);
or U17662 (N_17662,N_10229,N_13167);
and U17663 (N_17663,N_12174,N_13291);
nand U17664 (N_17664,N_14895,N_10692);
nor U17665 (N_17665,N_10558,N_14481);
xnor U17666 (N_17666,N_10600,N_12252);
nand U17667 (N_17667,N_11412,N_14683);
or U17668 (N_17668,N_12390,N_13671);
nor U17669 (N_17669,N_11292,N_13769);
and U17670 (N_17670,N_11280,N_13275);
nand U17671 (N_17671,N_10203,N_12094);
nand U17672 (N_17672,N_13629,N_12802);
nand U17673 (N_17673,N_14937,N_11268);
and U17674 (N_17674,N_12274,N_12962);
nor U17675 (N_17675,N_14735,N_12656);
or U17676 (N_17676,N_10638,N_12676);
or U17677 (N_17677,N_13921,N_11630);
or U17678 (N_17678,N_13692,N_11791);
or U17679 (N_17679,N_10118,N_10090);
nand U17680 (N_17680,N_12764,N_14646);
nor U17681 (N_17681,N_13626,N_14385);
xor U17682 (N_17682,N_11643,N_14948);
nand U17683 (N_17683,N_11915,N_13706);
nor U17684 (N_17684,N_13295,N_10880);
and U17685 (N_17685,N_14704,N_11725);
nor U17686 (N_17686,N_14958,N_10281);
xor U17687 (N_17687,N_13512,N_13043);
and U17688 (N_17688,N_10740,N_12552);
or U17689 (N_17689,N_11698,N_13215);
xnor U17690 (N_17690,N_14405,N_14943);
and U17691 (N_17691,N_11571,N_12492);
or U17692 (N_17692,N_13440,N_11113);
and U17693 (N_17693,N_12490,N_10203);
and U17694 (N_17694,N_13133,N_10422);
or U17695 (N_17695,N_12248,N_14138);
nand U17696 (N_17696,N_11806,N_13927);
nand U17697 (N_17697,N_12081,N_14273);
nand U17698 (N_17698,N_10170,N_12522);
xnor U17699 (N_17699,N_14903,N_11692);
xor U17700 (N_17700,N_12980,N_13142);
nand U17701 (N_17701,N_13028,N_14251);
nand U17702 (N_17702,N_14190,N_14363);
and U17703 (N_17703,N_10719,N_13797);
nand U17704 (N_17704,N_13870,N_12575);
xnor U17705 (N_17705,N_14427,N_14745);
nand U17706 (N_17706,N_12234,N_12995);
or U17707 (N_17707,N_11835,N_12005);
or U17708 (N_17708,N_12461,N_14213);
nand U17709 (N_17709,N_12134,N_13917);
nor U17710 (N_17710,N_14891,N_10636);
nor U17711 (N_17711,N_11602,N_14013);
and U17712 (N_17712,N_13951,N_11482);
and U17713 (N_17713,N_12026,N_12261);
or U17714 (N_17714,N_10875,N_11385);
nor U17715 (N_17715,N_12253,N_14348);
xnor U17716 (N_17716,N_11544,N_11335);
nor U17717 (N_17717,N_12310,N_11599);
or U17718 (N_17718,N_13300,N_12423);
nor U17719 (N_17719,N_12113,N_12121);
and U17720 (N_17720,N_11634,N_11657);
xnor U17721 (N_17721,N_13769,N_12639);
nand U17722 (N_17722,N_11515,N_12736);
nor U17723 (N_17723,N_10297,N_13559);
and U17724 (N_17724,N_14353,N_13872);
or U17725 (N_17725,N_11061,N_12303);
nand U17726 (N_17726,N_10495,N_10666);
nand U17727 (N_17727,N_13598,N_11971);
nand U17728 (N_17728,N_14927,N_10973);
and U17729 (N_17729,N_11505,N_12924);
and U17730 (N_17730,N_11590,N_13664);
and U17731 (N_17731,N_11126,N_12253);
and U17732 (N_17732,N_12009,N_10491);
xor U17733 (N_17733,N_12138,N_11204);
xor U17734 (N_17734,N_10973,N_14177);
or U17735 (N_17735,N_13078,N_13817);
nand U17736 (N_17736,N_13856,N_11739);
nor U17737 (N_17737,N_13228,N_13498);
and U17738 (N_17738,N_13955,N_10721);
or U17739 (N_17739,N_12149,N_10272);
and U17740 (N_17740,N_14315,N_14232);
or U17741 (N_17741,N_13151,N_11774);
and U17742 (N_17742,N_11553,N_14240);
nand U17743 (N_17743,N_11360,N_12590);
nor U17744 (N_17744,N_11097,N_10255);
nor U17745 (N_17745,N_14268,N_11181);
nand U17746 (N_17746,N_12669,N_10844);
nor U17747 (N_17747,N_11025,N_10077);
nor U17748 (N_17748,N_11285,N_12055);
and U17749 (N_17749,N_13280,N_12313);
nand U17750 (N_17750,N_14185,N_11266);
or U17751 (N_17751,N_14888,N_11798);
and U17752 (N_17752,N_12959,N_11319);
nand U17753 (N_17753,N_14695,N_11641);
nand U17754 (N_17754,N_12386,N_11448);
or U17755 (N_17755,N_13318,N_12311);
or U17756 (N_17756,N_14394,N_13956);
nor U17757 (N_17757,N_10869,N_10012);
and U17758 (N_17758,N_12823,N_12440);
nor U17759 (N_17759,N_13517,N_14793);
nand U17760 (N_17760,N_11911,N_13968);
or U17761 (N_17761,N_12107,N_14142);
nor U17762 (N_17762,N_13560,N_13285);
nor U17763 (N_17763,N_12267,N_13158);
and U17764 (N_17764,N_10024,N_11384);
nand U17765 (N_17765,N_14623,N_13819);
nor U17766 (N_17766,N_14446,N_13088);
and U17767 (N_17767,N_13479,N_11539);
nor U17768 (N_17768,N_14406,N_14821);
nor U17769 (N_17769,N_10629,N_14206);
and U17770 (N_17770,N_10678,N_14506);
nand U17771 (N_17771,N_14292,N_14511);
and U17772 (N_17772,N_14437,N_14057);
xnor U17773 (N_17773,N_11298,N_13953);
nor U17774 (N_17774,N_14458,N_12831);
nor U17775 (N_17775,N_11690,N_11596);
xnor U17776 (N_17776,N_10406,N_12481);
nand U17777 (N_17777,N_13442,N_13424);
or U17778 (N_17778,N_10818,N_10549);
xnor U17779 (N_17779,N_10417,N_12855);
nand U17780 (N_17780,N_10105,N_14026);
nor U17781 (N_17781,N_10816,N_13290);
or U17782 (N_17782,N_14565,N_14827);
nand U17783 (N_17783,N_10586,N_14248);
and U17784 (N_17784,N_11628,N_13076);
nor U17785 (N_17785,N_14271,N_10741);
and U17786 (N_17786,N_12297,N_10375);
or U17787 (N_17787,N_14831,N_14755);
nand U17788 (N_17788,N_13640,N_12198);
nand U17789 (N_17789,N_14472,N_14817);
and U17790 (N_17790,N_10217,N_13353);
or U17791 (N_17791,N_10303,N_11947);
xor U17792 (N_17792,N_14124,N_13912);
nand U17793 (N_17793,N_12862,N_10913);
nor U17794 (N_17794,N_10984,N_10784);
xnor U17795 (N_17795,N_12247,N_12060);
nor U17796 (N_17796,N_14422,N_14808);
nand U17797 (N_17797,N_14835,N_12772);
nand U17798 (N_17798,N_13053,N_11065);
nand U17799 (N_17799,N_13419,N_12916);
nand U17800 (N_17800,N_12945,N_13071);
nor U17801 (N_17801,N_13292,N_13552);
or U17802 (N_17802,N_12062,N_14842);
or U17803 (N_17803,N_11245,N_14660);
nand U17804 (N_17804,N_13549,N_11413);
and U17805 (N_17805,N_11272,N_13628);
nand U17806 (N_17806,N_13935,N_12810);
nand U17807 (N_17807,N_11326,N_10482);
or U17808 (N_17808,N_13176,N_12633);
nand U17809 (N_17809,N_12184,N_13307);
nand U17810 (N_17810,N_14775,N_10541);
nor U17811 (N_17811,N_14055,N_13361);
nor U17812 (N_17812,N_10911,N_11557);
and U17813 (N_17813,N_11113,N_13655);
and U17814 (N_17814,N_12868,N_10982);
or U17815 (N_17815,N_12291,N_12899);
nand U17816 (N_17816,N_10393,N_11731);
nor U17817 (N_17817,N_11445,N_11338);
and U17818 (N_17818,N_10955,N_12666);
or U17819 (N_17819,N_14600,N_10778);
nand U17820 (N_17820,N_12927,N_13192);
nor U17821 (N_17821,N_12841,N_12803);
or U17822 (N_17822,N_10223,N_10229);
and U17823 (N_17823,N_10723,N_11948);
xnor U17824 (N_17824,N_14909,N_14603);
or U17825 (N_17825,N_14980,N_11976);
xnor U17826 (N_17826,N_12511,N_14474);
and U17827 (N_17827,N_12361,N_13351);
nor U17828 (N_17828,N_13326,N_11252);
or U17829 (N_17829,N_11169,N_12723);
nor U17830 (N_17830,N_13147,N_14772);
nor U17831 (N_17831,N_13026,N_13452);
xor U17832 (N_17832,N_12907,N_13035);
or U17833 (N_17833,N_11885,N_11029);
nand U17834 (N_17834,N_11426,N_14914);
nor U17835 (N_17835,N_12314,N_12145);
nor U17836 (N_17836,N_11641,N_10692);
nor U17837 (N_17837,N_13939,N_10242);
nor U17838 (N_17838,N_12019,N_12905);
and U17839 (N_17839,N_10747,N_13639);
xor U17840 (N_17840,N_14199,N_11846);
and U17841 (N_17841,N_14004,N_13937);
and U17842 (N_17842,N_11965,N_12728);
nand U17843 (N_17843,N_10692,N_10376);
xnor U17844 (N_17844,N_14406,N_11303);
or U17845 (N_17845,N_13771,N_10915);
nand U17846 (N_17846,N_13756,N_10744);
nand U17847 (N_17847,N_11937,N_11651);
nand U17848 (N_17848,N_13048,N_11148);
nand U17849 (N_17849,N_12637,N_12329);
nand U17850 (N_17850,N_10578,N_10606);
and U17851 (N_17851,N_10185,N_14022);
nor U17852 (N_17852,N_11524,N_12253);
or U17853 (N_17853,N_13331,N_13595);
nor U17854 (N_17854,N_12245,N_14734);
nand U17855 (N_17855,N_12259,N_14406);
xor U17856 (N_17856,N_14744,N_14165);
and U17857 (N_17857,N_10038,N_12240);
or U17858 (N_17858,N_11940,N_13858);
or U17859 (N_17859,N_12172,N_12723);
and U17860 (N_17860,N_10100,N_11823);
and U17861 (N_17861,N_14288,N_11007);
nand U17862 (N_17862,N_13918,N_11186);
or U17863 (N_17863,N_11964,N_12340);
nor U17864 (N_17864,N_11170,N_10271);
nand U17865 (N_17865,N_13041,N_10228);
nor U17866 (N_17866,N_14815,N_14673);
xor U17867 (N_17867,N_11492,N_11739);
and U17868 (N_17868,N_14531,N_10199);
nand U17869 (N_17869,N_14706,N_13710);
and U17870 (N_17870,N_13047,N_12188);
xor U17871 (N_17871,N_12723,N_12435);
nor U17872 (N_17872,N_10885,N_11936);
and U17873 (N_17873,N_14616,N_10401);
nand U17874 (N_17874,N_10295,N_12309);
nor U17875 (N_17875,N_14493,N_11910);
nand U17876 (N_17876,N_10703,N_12825);
xnor U17877 (N_17877,N_11901,N_14676);
nor U17878 (N_17878,N_11138,N_11040);
or U17879 (N_17879,N_11503,N_14489);
nand U17880 (N_17880,N_11327,N_14880);
nor U17881 (N_17881,N_13226,N_11627);
and U17882 (N_17882,N_11316,N_11791);
nand U17883 (N_17883,N_11055,N_10191);
and U17884 (N_17884,N_10758,N_14294);
nand U17885 (N_17885,N_13113,N_12682);
and U17886 (N_17886,N_12474,N_13157);
and U17887 (N_17887,N_10637,N_12227);
nor U17888 (N_17888,N_14944,N_11218);
and U17889 (N_17889,N_11284,N_10524);
and U17890 (N_17890,N_11483,N_10351);
or U17891 (N_17891,N_13229,N_10375);
nor U17892 (N_17892,N_14409,N_12876);
and U17893 (N_17893,N_10651,N_11920);
nor U17894 (N_17894,N_13537,N_12588);
nor U17895 (N_17895,N_10027,N_13095);
nor U17896 (N_17896,N_14148,N_13143);
nand U17897 (N_17897,N_10196,N_11977);
and U17898 (N_17898,N_13875,N_12771);
or U17899 (N_17899,N_13634,N_12735);
nor U17900 (N_17900,N_14120,N_11909);
or U17901 (N_17901,N_12655,N_10349);
nand U17902 (N_17902,N_13603,N_13413);
or U17903 (N_17903,N_11388,N_10437);
or U17904 (N_17904,N_11538,N_10406);
and U17905 (N_17905,N_13769,N_12334);
nor U17906 (N_17906,N_12898,N_13824);
or U17907 (N_17907,N_12878,N_14077);
and U17908 (N_17908,N_12322,N_12225);
or U17909 (N_17909,N_14991,N_10608);
or U17910 (N_17910,N_12687,N_14416);
nand U17911 (N_17911,N_11223,N_14272);
and U17912 (N_17912,N_13516,N_11765);
xor U17913 (N_17913,N_14039,N_14736);
or U17914 (N_17914,N_12317,N_12193);
nor U17915 (N_17915,N_14016,N_12903);
or U17916 (N_17916,N_13464,N_14329);
nor U17917 (N_17917,N_13108,N_14575);
nand U17918 (N_17918,N_11154,N_12550);
or U17919 (N_17919,N_11752,N_10286);
nand U17920 (N_17920,N_10701,N_11316);
nand U17921 (N_17921,N_11572,N_12752);
or U17922 (N_17922,N_12955,N_14934);
or U17923 (N_17923,N_11634,N_11283);
nand U17924 (N_17924,N_11667,N_13357);
nand U17925 (N_17925,N_12405,N_10746);
or U17926 (N_17926,N_13252,N_14471);
nand U17927 (N_17927,N_14114,N_14867);
xor U17928 (N_17928,N_13773,N_12184);
xnor U17929 (N_17929,N_14678,N_11352);
or U17930 (N_17930,N_14037,N_12641);
nand U17931 (N_17931,N_13313,N_13622);
nor U17932 (N_17932,N_11477,N_10062);
and U17933 (N_17933,N_10915,N_14348);
nand U17934 (N_17934,N_13764,N_14528);
or U17935 (N_17935,N_14043,N_14270);
nand U17936 (N_17936,N_14957,N_10902);
nor U17937 (N_17937,N_14483,N_10836);
and U17938 (N_17938,N_14999,N_12664);
xnor U17939 (N_17939,N_10382,N_11976);
nand U17940 (N_17940,N_10132,N_14478);
and U17941 (N_17941,N_14546,N_10127);
or U17942 (N_17942,N_14690,N_10966);
or U17943 (N_17943,N_13104,N_13949);
xor U17944 (N_17944,N_10163,N_11734);
xnor U17945 (N_17945,N_12620,N_14146);
nor U17946 (N_17946,N_10252,N_10989);
and U17947 (N_17947,N_12794,N_10674);
nor U17948 (N_17948,N_10024,N_13798);
and U17949 (N_17949,N_14251,N_14753);
nor U17950 (N_17950,N_13500,N_12682);
or U17951 (N_17951,N_13922,N_12291);
or U17952 (N_17952,N_10225,N_12288);
nor U17953 (N_17953,N_14009,N_10873);
or U17954 (N_17954,N_13284,N_10030);
nor U17955 (N_17955,N_13593,N_10865);
nand U17956 (N_17956,N_13010,N_13901);
nand U17957 (N_17957,N_13823,N_14974);
nor U17958 (N_17958,N_11758,N_13414);
and U17959 (N_17959,N_13027,N_11767);
or U17960 (N_17960,N_10545,N_10774);
xnor U17961 (N_17961,N_11053,N_10216);
and U17962 (N_17962,N_14967,N_14704);
or U17963 (N_17963,N_14975,N_11748);
nand U17964 (N_17964,N_11647,N_11819);
nor U17965 (N_17965,N_12299,N_13423);
or U17966 (N_17966,N_14591,N_11168);
or U17967 (N_17967,N_11719,N_11016);
or U17968 (N_17968,N_11974,N_14681);
nand U17969 (N_17969,N_12104,N_12235);
nor U17970 (N_17970,N_10073,N_12496);
or U17971 (N_17971,N_11293,N_13934);
nor U17972 (N_17972,N_11804,N_11258);
or U17973 (N_17973,N_14687,N_12431);
nand U17974 (N_17974,N_11881,N_12076);
nor U17975 (N_17975,N_12970,N_12286);
and U17976 (N_17976,N_11390,N_11337);
nor U17977 (N_17977,N_12642,N_12662);
nand U17978 (N_17978,N_12637,N_11814);
and U17979 (N_17979,N_13330,N_11278);
and U17980 (N_17980,N_14265,N_10586);
nand U17981 (N_17981,N_11589,N_11750);
or U17982 (N_17982,N_12481,N_12763);
nand U17983 (N_17983,N_14426,N_12967);
xor U17984 (N_17984,N_11504,N_12031);
or U17985 (N_17985,N_13605,N_14721);
and U17986 (N_17986,N_11373,N_11073);
xor U17987 (N_17987,N_10464,N_13266);
nor U17988 (N_17988,N_10763,N_13827);
or U17989 (N_17989,N_10004,N_14595);
nor U17990 (N_17990,N_11151,N_12373);
xnor U17991 (N_17991,N_12842,N_14503);
nand U17992 (N_17992,N_12716,N_14342);
nor U17993 (N_17993,N_10829,N_12145);
or U17994 (N_17994,N_14556,N_11835);
and U17995 (N_17995,N_14754,N_12722);
and U17996 (N_17996,N_11331,N_11601);
nor U17997 (N_17997,N_13242,N_10838);
nand U17998 (N_17998,N_10747,N_14286);
and U17999 (N_17999,N_14342,N_12010);
xor U18000 (N_18000,N_10768,N_10435);
and U18001 (N_18001,N_10908,N_10651);
nand U18002 (N_18002,N_14099,N_13053);
nand U18003 (N_18003,N_14069,N_11029);
xor U18004 (N_18004,N_11580,N_14037);
nor U18005 (N_18005,N_14474,N_11767);
xnor U18006 (N_18006,N_11201,N_11233);
or U18007 (N_18007,N_14051,N_11475);
or U18008 (N_18008,N_12165,N_11624);
or U18009 (N_18009,N_11296,N_11014);
or U18010 (N_18010,N_14045,N_10892);
or U18011 (N_18011,N_14772,N_12823);
xnor U18012 (N_18012,N_12643,N_11680);
and U18013 (N_18013,N_12892,N_11847);
nand U18014 (N_18014,N_11510,N_13478);
or U18015 (N_18015,N_12790,N_12884);
nand U18016 (N_18016,N_13998,N_13811);
nand U18017 (N_18017,N_10929,N_11583);
and U18018 (N_18018,N_12705,N_13977);
nor U18019 (N_18019,N_13223,N_11567);
nand U18020 (N_18020,N_11995,N_14213);
or U18021 (N_18021,N_10658,N_10073);
and U18022 (N_18022,N_10168,N_13108);
xnor U18023 (N_18023,N_13614,N_13190);
and U18024 (N_18024,N_14267,N_13582);
nor U18025 (N_18025,N_12756,N_13695);
or U18026 (N_18026,N_13928,N_11518);
nand U18027 (N_18027,N_14815,N_13836);
nor U18028 (N_18028,N_13072,N_11161);
or U18029 (N_18029,N_10148,N_10194);
and U18030 (N_18030,N_13481,N_11364);
or U18031 (N_18031,N_13957,N_13147);
nor U18032 (N_18032,N_11281,N_12552);
nor U18033 (N_18033,N_11167,N_11801);
or U18034 (N_18034,N_12888,N_11853);
and U18035 (N_18035,N_13613,N_12704);
or U18036 (N_18036,N_11911,N_12456);
nand U18037 (N_18037,N_10443,N_14445);
or U18038 (N_18038,N_10786,N_13722);
xor U18039 (N_18039,N_10340,N_13656);
and U18040 (N_18040,N_10646,N_13639);
or U18041 (N_18041,N_10936,N_10403);
nand U18042 (N_18042,N_13110,N_11037);
nand U18043 (N_18043,N_12684,N_10865);
and U18044 (N_18044,N_14535,N_13250);
and U18045 (N_18045,N_13852,N_10891);
nor U18046 (N_18046,N_10952,N_13037);
xnor U18047 (N_18047,N_14031,N_12641);
and U18048 (N_18048,N_11375,N_14775);
and U18049 (N_18049,N_12227,N_11925);
or U18050 (N_18050,N_10179,N_13947);
nor U18051 (N_18051,N_14788,N_14796);
nand U18052 (N_18052,N_14750,N_12141);
nor U18053 (N_18053,N_13853,N_14746);
nor U18054 (N_18054,N_13209,N_11985);
or U18055 (N_18055,N_14191,N_11222);
nor U18056 (N_18056,N_14271,N_14227);
nor U18057 (N_18057,N_13401,N_11584);
nand U18058 (N_18058,N_12921,N_13166);
nand U18059 (N_18059,N_14549,N_10197);
nand U18060 (N_18060,N_14174,N_13732);
xnor U18061 (N_18061,N_10405,N_14913);
and U18062 (N_18062,N_10581,N_14082);
or U18063 (N_18063,N_10506,N_14679);
nor U18064 (N_18064,N_14832,N_11336);
xor U18065 (N_18065,N_10670,N_10754);
and U18066 (N_18066,N_10418,N_10165);
and U18067 (N_18067,N_13312,N_12717);
and U18068 (N_18068,N_13739,N_10633);
and U18069 (N_18069,N_11715,N_11514);
nor U18070 (N_18070,N_10379,N_10649);
nand U18071 (N_18071,N_14074,N_12966);
or U18072 (N_18072,N_12718,N_11749);
nand U18073 (N_18073,N_13209,N_10048);
nor U18074 (N_18074,N_14895,N_13813);
or U18075 (N_18075,N_13617,N_14433);
xor U18076 (N_18076,N_12034,N_11754);
xnor U18077 (N_18077,N_10942,N_14006);
and U18078 (N_18078,N_11507,N_10816);
nand U18079 (N_18079,N_10502,N_12183);
nand U18080 (N_18080,N_14997,N_11778);
nand U18081 (N_18081,N_12286,N_14488);
or U18082 (N_18082,N_13413,N_12951);
nand U18083 (N_18083,N_13071,N_13569);
or U18084 (N_18084,N_10398,N_11776);
nand U18085 (N_18085,N_14290,N_10963);
or U18086 (N_18086,N_13171,N_11321);
nand U18087 (N_18087,N_13142,N_14060);
nor U18088 (N_18088,N_12473,N_11364);
or U18089 (N_18089,N_13711,N_10712);
and U18090 (N_18090,N_14720,N_14206);
nand U18091 (N_18091,N_10998,N_13689);
nand U18092 (N_18092,N_14240,N_13530);
nor U18093 (N_18093,N_14700,N_14703);
nand U18094 (N_18094,N_10298,N_13784);
or U18095 (N_18095,N_14326,N_14272);
xor U18096 (N_18096,N_14893,N_12538);
and U18097 (N_18097,N_13944,N_10154);
xnor U18098 (N_18098,N_13102,N_14229);
xor U18099 (N_18099,N_10585,N_11201);
nand U18100 (N_18100,N_14406,N_13811);
and U18101 (N_18101,N_13724,N_12218);
and U18102 (N_18102,N_11149,N_11988);
xor U18103 (N_18103,N_14173,N_10750);
nor U18104 (N_18104,N_12251,N_13134);
or U18105 (N_18105,N_12397,N_10804);
or U18106 (N_18106,N_11376,N_14719);
nor U18107 (N_18107,N_12410,N_11735);
or U18108 (N_18108,N_11078,N_14940);
or U18109 (N_18109,N_11771,N_12698);
nor U18110 (N_18110,N_14362,N_13410);
nand U18111 (N_18111,N_12667,N_13859);
xnor U18112 (N_18112,N_11145,N_14582);
and U18113 (N_18113,N_13544,N_12047);
and U18114 (N_18114,N_10419,N_10191);
and U18115 (N_18115,N_11879,N_14522);
and U18116 (N_18116,N_11868,N_12678);
nor U18117 (N_18117,N_13394,N_12975);
nor U18118 (N_18118,N_13729,N_11279);
nor U18119 (N_18119,N_14725,N_13345);
and U18120 (N_18120,N_11137,N_10380);
and U18121 (N_18121,N_14918,N_10010);
or U18122 (N_18122,N_12100,N_14804);
or U18123 (N_18123,N_12865,N_12487);
and U18124 (N_18124,N_11480,N_11034);
or U18125 (N_18125,N_10920,N_12357);
xnor U18126 (N_18126,N_10065,N_11246);
xor U18127 (N_18127,N_14596,N_11054);
nor U18128 (N_18128,N_12451,N_12122);
nand U18129 (N_18129,N_13309,N_13613);
nand U18130 (N_18130,N_10748,N_10393);
or U18131 (N_18131,N_14369,N_10897);
or U18132 (N_18132,N_10322,N_10970);
and U18133 (N_18133,N_13492,N_10247);
or U18134 (N_18134,N_11326,N_11424);
nor U18135 (N_18135,N_13931,N_12450);
nor U18136 (N_18136,N_11040,N_12902);
nand U18137 (N_18137,N_14610,N_12496);
nor U18138 (N_18138,N_12757,N_12815);
and U18139 (N_18139,N_10518,N_12433);
or U18140 (N_18140,N_13196,N_12003);
and U18141 (N_18141,N_12414,N_14416);
and U18142 (N_18142,N_10805,N_14762);
and U18143 (N_18143,N_13432,N_11993);
nor U18144 (N_18144,N_14045,N_13693);
nand U18145 (N_18145,N_12779,N_10538);
nor U18146 (N_18146,N_10788,N_14706);
nand U18147 (N_18147,N_12653,N_14843);
or U18148 (N_18148,N_14227,N_10870);
nor U18149 (N_18149,N_12216,N_10872);
and U18150 (N_18150,N_12971,N_14455);
nor U18151 (N_18151,N_12356,N_12251);
or U18152 (N_18152,N_13658,N_10665);
or U18153 (N_18153,N_13552,N_12177);
or U18154 (N_18154,N_10338,N_14320);
xor U18155 (N_18155,N_13859,N_11178);
and U18156 (N_18156,N_13617,N_14925);
or U18157 (N_18157,N_11874,N_10800);
and U18158 (N_18158,N_11981,N_14841);
or U18159 (N_18159,N_10314,N_10194);
nor U18160 (N_18160,N_10017,N_10589);
nor U18161 (N_18161,N_14173,N_11316);
nand U18162 (N_18162,N_12134,N_13097);
and U18163 (N_18163,N_11292,N_13838);
xnor U18164 (N_18164,N_12885,N_11707);
or U18165 (N_18165,N_13586,N_12502);
and U18166 (N_18166,N_12256,N_13179);
and U18167 (N_18167,N_14580,N_12077);
nand U18168 (N_18168,N_10988,N_14794);
and U18169 (N_18169,N_11196,N_12383);
nand U18170 (N_18170,N_13116,N_11801);
nand U18171 (N_18171,N_11314,N_10833);
nand U18172 (N_18172,N_10052,N_11232);
nand U18173 (N_18173,N_12851,N_14854);
or U18174 (N_18174,N_13566,N_13633);
nor U18175 (N_18175,N_11755,N_10577);
nor U18176 (N_18176,N_14984,N_13234);
xnor U18177 (N_18177,N_10058,N_12818);
nor U18178 (N_18178,N_14768,N_12819);
nor U18179 (N_18179,N_14099,N_11496);
or U18180 (N_18180,N_12790,N_13573);
or U18181 (N_18181,N_11278,N_10572);
and U18182 (N_18182,N_11633,N_12946);
and U18183 (N_18183,N_12808,N_10537);
nand U18184 (N_18184,N_12071,N_13095);
or U18185 (N_18185,N_11190,N_10037);
xnor U18186 (N_18186,N_11257,N_14867);
nand U18187 (N_18187,N_14872,N_12007);
or U18188 (N_18188,N_13639,N_14084);
xnor U18189 (N_18189,N_13511,N_12647);
xnor U18190 (N_18190,N_11191,N_13512);
nor U18191 (N_18191,N_10296,N_14253);
nor U18192 (N_18192,N_11863,N_10179);
nor U18193 (N_18193,N_12511,N_14516);
xor U18194 (N_18194,N_11967,N_13365);
or U18195 (N_18195,N_13074,N_14633);
xor U18196 (N_18196,N_14732,N_14586);
or U18197 (N_18197,N_10597,N_10547);
or U18198 (N_18198,N_11989,N_11223);
nand U18199 (N_18199,N_14562,N_10860);
or U18200 (N_18200,N_11903,N_14039);
or U18201 (N_18201,N_13105,N_11201);
nor U18202 (N_18202,N_10053,N_14682);
or U18203 (N_18203,N_13348,N_10485);
or U18204 (N_18204,N_13312,N_12626);
nor U18205 (N_18205,N_10921,N_13906);
nor U18206 (N_18206,N_12642,N_12499);
or U18207 (N_18207,N_14324,N_10522);
nor U18208 (N_18208,N_12176,N_14125);
xor U18209 (N_18209,N_10790,N_13337);
nand U18210 (N_18210,N_12298,N_12299);
or U18211 (N_18211,N_10604,N_14126);
or U18212 (N_18212,N_13179,N_14938);
and U18213 (N_18213,N_12752,N_12376);
nor U18214 (N_18214,N_12572,N_14845);
or U18215 (N_18215,N_13916,N_13966);
or U18216 (N_18216,N_12449,N_13733);
nand U18217 (N_18217,N_12080,N_13739);
and U18218 (N_18218,N_12761,N_12063);
nor U18219 (N_18219,N_13043,N_13775);
nor U18220 (N_18220,N_11628,N_13491);
nand U18221 (N_18221,N_11771,N_12185);
and U18222 (N_18222,N_12959,N_13360);
nand U18223 (N_18223,N_13388,N_11277);
and U18224 (N_18224,N_12649,N_12765);
and U18225 (N_18225,N_12832,N_14136);
nor U18226 (N_18226,N_10362,N_10813);
or U18227 (N_18227,N_14192,N_13961);
and U18228 (N_18228,N_11673,N_11516);
nor U18229 (N_18229,N_10300,N_11434);
and U18230 (N_18230,N_14339,N_13236);
nor U18231 (N_18231,N_10192,N_13399);
or U18232 (N_18232,N_13659,N_12591);
nor U18233 (N_18233,N_10986,N_14953);
or U18234 (N_18234,N_14579,N_13113);
or U18235 (N_18235,N_12288,N_10016);
nand U18236 (N_18236,N_12099,N_11279);
or U18237 (N_18237,N_11593,N_12811);
or U18238 (N_18238,N_11983,N_12897);
or U18239 (N_18239,N_13127,N_13508);
and U18240 (N_18240,N_14599,N_10043);
or U18241 (N_18241,N_13848,N_10276);
xnor U18242 (N_18242,N_11393,N_13665);
nor U18243 (N_18243,N_14659,N_14314);
or U18244 (N_18244,N_11629,N_11010);
or U18245 (N_18245,N_10606,N_12393);
or U18246 (N_18246,N_13527,N_12061);
nand U18247 (N_18247,N_11428,N_10707);
and U18248 (N_18248,N_14568,N_12205);
nor U18249 (N_18249,N_11918,N_12332);
and U18250 (N_18250,N_12700,N_10095);
or U18251 (N_18251,N_14707,N_14854);
nand U18252 (N_18252,N_13167,N_12527);
nand U18253 (N_18253,N_10619,N_13061);
nor U18254 (N_18254,N_11727,N_10570);
or U18255 (N_18255,N_11670,N_11310);
xnor U18256 (N_18256,N_12671,N_14274);
and U18257 (N_18257,N_11111,N_12005);
nand U18258 (N_18258,N_14202,N_11302);
and U18259 (N_18259,N_11502,N_12013);
nor U18260 (N_18260,N_10390,N_13096);
nand U18261 (N_18261,N_13660,N_12697);
or U18262 (N_18262,N_14214,N_10420);
nand U18263 (N_18263,N_13143,N_11294);
nor U18264 (N_18264,N_13580,N_12563);
nand U18265 (N_18265,N_12422,N_13709);
nor U18266 (N_18266,N_14423,N_11773);
and U18267 (N_18267,N_10445,N_13022);
nand U18268 (N_18268,N_11149,N_13755);
nor U18269 (N_18269,N_12488,N_13421);
and U18270 (N_18270,N_14593,N_14158);
nand U18271 (N_18271,N_12849,N_13040);
or U18272 (N_18272,N_12352,N_13405);
nand U18273 (N_18273,N_13174,N_10889);
nor U18274 (N_18274,N_14979,N_12933);
nor U18275 (N_18275,N_12435,N_13340);
or U18276 (N_18276,N_14834,N_13792);
or U18277 (N_18277,N_11972,N_12065);
nand U18278 (N_18278,N_11183,N_13558);
xnor U18279 (N_18279,N_13323,N_12402);
xnor U18280 (N_18280,N_13598,N_12312);
nor U18281 (N_18281,N_10089,N_14852);
nand U18282 (N_18282,N_10844,N_11300);
and U18283 (N_18283,N_11676,N_12150);
or U18284 (N_18284,N_11815,N_13393);
and U18285 (N_18285,N_12665,N_12185);
or U18286 (N_18286,N_14036,N_11189);
and U18287 (N_18287,N_13509,N_11506);
nand U18288 (N_18288,N_10598,N_10627);
or U18289 (N_18289,N_10263,N_11688);
nor U18290 (N_18290,N_10631,N_10658);
or U18291 (N_18291,N_13018,N_14773);
nor U18292 (N_18292,N_10176,N_13377);
and U18293 (N_18293,N_12984,N_14349);
or U18294 (N_18294,N_13566,N_13796);
or U18295 (N_18295,N_14001,N_10275);
and U18296 (N_18296,N_13102,N_11580);
and U18297 (N_18297,N_13989,N_11925);
nand U18298 (N_18298,N_13549,N_14665);
nand U18299 (N_18299,N_10048,N_11043);
xor U18300 (N_18300,N_14468,N_13264);
nand U18301 (N_18301,N_13399,N_12156);
and U18302 (N_18302,N_14687,N_10814);
nor U18303 (N_18303,N_13614,N_12167);
nor U18304 (N_18304,N_12877,N_14158);
or U18305 (N_18305,N_14631,N_14167);
or U18306 (N_18306,N_12083,N_13487);
xor U18307 (N_18307,N_12601,N_13652);
nor U18308 (N_18308,N_10245,N_14436);
nand U18309 (N_18309,N_14275,N_11287);
xnor U18310 (N_18310,N_14189,N_10558);
nor U18311 (N_18311,N_11660,N_13462);
and U18312 (N_18312,N_14668,N_13381);
or U18313 (N_18313,N_12331,N_13548);
xnor U18314 (N_18314,N_14318,N_10074);
nand U18315 (N_18315,N_11889,N_12843);
or U18316 (N_18316,N_14192,N_14150);
nor U18317 (N_18317,N_11861,N_10724);
nand U18318 (N_18318,N_14559,N_14812);
or U18319 (N_18319,N_10193,N_14549);
or U18320 (N_18320,N_14631,N_10461);
nor U18321 (N_18321,N_10083,N_14483);
or U18322 (N_18322,N_14640,N_10574);
and U18323 (N_18323,N_11518,N_11948);
and U18324 (N_18324,N_14067,N_12268);
and U18325 (N_18325,N_14829,N_11629);
nand U18326 (N_18326,N_11831,N_12934);
xor U18327 (N_18327,N_14210,N_11844);
nand U18328 (N_18328,N_11820,N_12699);
and U18329 (N_18329,N_12014,N_12667);
nand U18330 (N_18330,N_13682,N_13415);
nor U18331 (N_18331,N_13661,N_10107);
or U18332 (N_18332,N_11268,N_13288);
and U18333 (N_18333,N_13816,N_14865);
nor U18334 (N_18334,N_10967,N_11792);
nor U18335 (N_18335,N_11478,N_11838);
nand U18336 (N_18336,N_10132,N_11369);
nand U18337 (N_18337,N_10283,N_13920);
or U18338 (N_18338,N_10612,N_12220);
xor U18339 (N_18339,N_11307,N_13550);
and U18340 (N_18340,N_13429,N_13257);
and U18341 (N_18341,N_13062,N_10545);
or U18342 (N_18342,N_13561,N_10212);
nor U18343 (N_18343,N_13165,N_10527);
nor U18344 (N_18344,N_12200,N_12577);
xnor U18345 (N_18345,N_12252,N_10376);
nor U18346 (N_18346,N_12486,N_14057);
and U18347 (N_18347,N_12722,N_12783);
and U18348 (N_18348,N_10834,N_11445);
nand U18349 (N_18349,N_10627,N_11809);
and U18350 (N_18350,N_10489,N_12315);
or U18351 (N_18351,N_13316,N_14791);
nor U18352 (N_18352,N_12563,N_13407);
or U18353 (N_18353,N_13102,N_12386);
and U18354 (N_18354,N_10693,N_14121);
nor U18355 (N_18355,N_11744,N_13245);
and U18356 (N_18356,N_14178,N_10337);
nand U18357 (N_18357,N_13140,N_10488);
or U18358 (N_18358,N_11870,N_13836);
or U18359 (N_18359,N_11748,N_13289);
and U18360 (N_18360,N_10179,N_14318);
or U18361 (N_18361,N_12355,N_13999);
xor U18362 (N_18362,N_11311,N_10623);
nor U18363 (N_18363,N_12545,N_10561);
nand U18364 (N_18364,N_11445,N_10056);
nor U18365 (N_18365,N_14812,N_10194);
and U18366 (N_18366,N_12890,N_11162);
nand U18367 (N_18367,N_10996,N_10659);
and U18368 (N_18368,N_14693,N_10502);
nor U18369 (N_18369,N_12254,N_10498);
xnor U18370 (N_18370,N_12614,N_13934);
or U18371 (N_18371,N_11183,N_12359);
or U18372 (N_18372,N_10747,N_13638);
nor U18373 (N_18373,N_12942,N_11774);
and U18374 (N_18374,N_13535,N_12699);
and U18375 (N_18375,N_13237,N_14981);
nor U18376 (N_18376,N_12854,N_11792);
xor U18377 (N_18377,N_11541,N_10784);
nor U18378 (N_18378,N_11221,N_10095);
or U18379 (N_18379,N_11843,N_10311);
nor U18380 (N_18380,N_13256,N_10198);
or U18381 (N_18381,N_10825,N_14022);
or U18382 (N_18382,N_10571,N_12125);
or U18383 (N_18383,N_11779,N_11573);
nor U18384 (N_18384,N_13147,N_14018);
nand U18385 (N_18385,N_11405,N_11034);
xnor U18386 (N_18386,N_11707,N_14673);
and U18387 (N_18387,N_13752,N_12085);
or U18388 (N_18388,N_11614,N_11383);
nand U18389 (N_18389,N_10923,N_11508);
nand U18390 (N_18390,N_11637,N_13067);
and U18391 (N_18391,N_14759,N_10644);
and U18392 (N_18392,N_10708,N_11432);
nand U18393 (N_18393,N_10807,N_13033);
nor U18394 (N_18394,N_11486,N_14036);
and U18395 (N_18395,N_10601,N_14034);
xor U18396 (N_18396,N_11464,N_13158);
and U18397 (N_18397,N_14081,N_10262);
nand U18398 (N_18398,N_10622,N_10783);
nand U18399 (N_18399,N_14801,N_14382);
nor U18400 (N_18400,N_11482,N_11681);
nand U18401 (N_18401,N_10102,N_13865);
nand U18402 (N_18402,N_13033,N_10806);
nand U18403 (N_18403,N_10589,N_12333);
or U18404 (N_18404,N_13829,N_12973);
and U18405 (N_18405,N_12543,N_11911);
and U18406 (N_18406,N_12985,N_10555);
nand U18407 (N_18407,N_12574,N_12190);
or U18408 (N_18408,N_14945,N_11575);
and U18409 (N_18409,N_11629,N_10492);
and U18410 (N_18410,N_13131,N_10099);
and U18411 (N_18411,N_10487,N_10540);
or U18412 (N_18412,N_10325,N_10611);
xor U18413 (N_18413,N_14583,N_14633);
nor U18414 (N_18414,N_14484,N_14897);
nand U18415 (N_18415,N_12248,N_11022);
and U18416 (N_18416,N_11463,N_11171);
nand U18417 (N_18417,N_10484,N_11474);
and U18418 (N_18418,N_10796,N_14577);
nor U18419 (N_18419,N_10953,N_14979);
nand U18420 (N_18420,N_13709,N_10894);
nor U18421 (N_18421,N_11404,N_14451);
nor U18422 (N_18422,N_12346,N_12343);
xor U18423 (N_18423,N_11697,N_14337);
nor U18424 (N_18424,N_14673,N_11984);
nand U18425 (N_18425,N_13531,N_14701);
nand U18426 (N_18426,N_13411,N_12298);
nor U18427 (N_18427,N_14705,N_14338);
and U18428 (N_18428,N_12516,N_12929);
nor U18429 (N_18429,N_11669,N_11901);
and U18430 (N_18430,N_12159,N_11822);
xor U18431 (N_18431,N_13735,N_11395);
nand U18432 (N_18432,N_14429,N_12782);
xor U18433 (N_18433,N_13716,N_10610);
nand U18434 (N_18434,N_11070,N_13399);
or U18435 (N_18435,N_10832,N_11359);
and U18436 (N_18436,N_14825,N_13666);
or U18437 (N_18437,N_14945,N_10744);
nor U18438 (N_18438,N_11664,N_13084);
or U18439 (N_18439,N_11209,N_10734);
xor U18440 (N_18440,N_14070,N_10731);
nand U18441 (N_18441,N_11790,N_14509);
nand U18442 (N_18442,N_13885,N_10002);
nor U18443 (N_18443,N_14649,N_11093);
nor U18444 (N_18444,N_14184,N_13832);
or U18445 (N_18445,N_14937,N_11397);
or U18446 (N_18446,N_11826,N_13410);
nand U18447 (N_18447,N_14312,N_14730);
nand U18448 (N_18448,N_14169,N_13989);
nor U18449 (N_18449,N_13638,N_12271);
nor U18450 (N_18450,N_10758,N_13345);
xor U18451 (N_18451,N_14634,N_13316);
or U18452 (N_18452,N_14724,N_10588);
nand U18453 (N_18453,N_13900,N_14184);
xnor U18454 (N_18454,N_10245,N_14525);
or U18455 (N_18455,N_12619,N_14481);
nor U18456 (N_18456,N_13549,N_14558);
and U18457 (N_18457,N_12404,N_10733);
and U18458 (N_18458,N_10076,N_13035);
nand U18459 (N_18459,N_11795,N_13223);
nand U18460 (N_18460,N_13202,N_10242);
nand U18461 (N_18461,N_10256,N_12825);
or U18462 (N_18462,N_13615,N_12803);
and U18463 (N_18463,N_11316,N_12330);
nand U18464 (N_18464,N_11368,N_13946);
xnor U18465 (N_18465,N_14921,N_12000);
nand U18466 (N_18466,N_13125,N_14807);
nand U18467 (N_18467,N_10409,N_10574);
and U18468 (N_18468,N_14890,N_12111);
nand U18469 (N_18469,N_11983,N_12887);
nor U18470 (N_18470,N_11453,N_10706);
nor U18471 (N_18471,N_10468,N_13553);
or U18472 (N_18472,N_11934,N_14329);
xor U18473 (N_18473,N_13852,N_14797);
nand U18474 (N_18474,N_11464,N_12450);
nand U18475 (N_18475,N_12495,N_10494);
nor U18476 (N_18476,N_14247,N_11962);
nor U18477 (N_18477,N_10980,N_12467);
and U18478 (N_18478,N_12638,N_14556);
and U18479 (N_18479,N_11733,N_14237);
nor U18480 (N_18480,N_13212,N_11942);
or U18481 (N_18481,N_14799,N_10819);
nor U18482 (N_18482,N_10335,N_14435);
nor U18483 (N_18483,N_14197,N_11694);
nand U18484 (N_18484,N_14319,N_10550);
and U18485 (N_18485,N_13278,N_13030);
or U18486 (N_18486,N_14840,N_10892);
nand U18487 (N_18487,N_14854,N_10125);
or U18488 (N_18488,N_13366,N_11352);
or U18489 (N_18489,N_11755,N_13163);
or U18490 (N_18490,N_11027,N_14848);
or U18491 (N_18491,N_11785,N_11130);
or U18492 (N_18492,N_14329,N_11615);
and U18493 (N_18493,N_14719,N_11246);
or U18494 (N_18494,N_13686,N_10065);
xor U18495 (N_18495,N_11502,N_14788);
and U18496 (N_18496,N_12259,N_13793);
nand U18497 (N_18497,N_12601,N_12135);
nor U18498 (N_18498,N_12208,N_14557);
and U18499 (N_18499,N_14940,N_13999);
nand U18500 (N_18500,N_12119,N_14400);
nor U18501 (N_18501,N_14128,N_14813);
nand U18502 (N_18502,N_10074,N_11735);
or U18503 (N_18503,N_11592,N_14501);
nand U18504 (N_18504,N_13132,N_12030);
nor U18505 (N_18505,N_11631,N_13713);
nand U18506 (N_18506,N_13709,N_12174);
or U18507 (N_18507,N_12797,N_11927);
xor U18508 (N_18508,N_13159,N_13371);
nand U18509 (N_18509,N_11218,N_10573);
nand U18510 (N_18510,N_13420,N_10243);
nand U18511 (N_18511,N_12967,N_11104);
nor U18512 (N_18512,N_12380,N_11998);
nand U18513 (N_18513,N_12151,N_10266);
nand U18514 (N_18514,N_10767,N_11758);
nand U18515 (N_18515,N_11074,N_10570);
and U18516 (N_18516,N_11368,N_12509);
nor U18517 (N_18517,N_13273,N_11507);
and U18518 (N_18518,N_14856,N_14900);
nand U18519 (N_18519,N_12957,N_10311);
nand U18520 (N_18520,N_12844,N_10607);
nand U18521 (N_18521,N_13248,N_14619);
nand U18522 (N_18522,N_13408,N_12743);
and U18523 (N_18523,N_12292,N_10216);
and U18524 (N_18524,N_12850,N_14481);
xor U18525 (N_18525,N_14267,N_13204);
or U18526 (N_18526,N_11405,N_10181);
nor U18527 (N_18527,N_14849,N_12312);
nand U18528 (N_18528,N_10807,N_10075);
nor U18529 (N_18529,N_13402,N_10842);
or U18530 (N_18530,N_12026,N_11061);
nand U18531 (N_18531,N_11898,N_10740);
or U18532 (N_18532,N_10774,N_11163);
xnor U18533 (N_18533,N_14670,N_10008);
nand U18534 (N_18534,N_10788,N_14028);
nand U18535 (N_18535,N_12477,N_11383);
and U18536 (N_18536,N_11202,N_14889);
and U18537 (N_18537,N_13482,N_14494);
nand U18538 (N_18538,N_11850,N_13756);
nor U18539 (N_18539,N_11861,N_14304);
or U18540 (N_18540,N_10203,N_13875);
and U18541 (N_18541,N_13834,N_12262);
and U18542 (N_18542,N_14800,N_14621);
nand U18543 (N_18543,N_11929,N_11627);
nand U18544 (N_18544,N_13268,N_11807);
and U18545 (N_18545,N_11757,N_13284);
nor U18546 (N_18546,N_14232,N_10068);
and U18547 (N_18547,N_10631,N_14748);
and U18548 (N_18548,N_12726,N_12590);
nand U18549 (N_18549,N_13881,N_12064);
and U18550 (N_18550,N_14489,N_10062);
nand U18551 (N_18551,N_14419,N_13213);
and U18552 (N_18552,N_11584,N_11651);
nand U18553 (N_18553,N_10415,N_13134);
and U18554 (N_18554,N_13658,N_11838);
nor U18555 (N_18555,N_12988,N_11387);
xnor U18556 (N_18556,N_11826,N_13429);
xnor U18557 (N_18557,N_13710,N_10560);
and U18558 (N_18558,N_10509,N_13843);
nand U18559 (N_18559,N_11946,N_12297);
and U18560 (N_18560,N_12272,N_12774);
or U18561 (N_18561,N_13210,N_12130);
nand U18562 (N_18562,N_13411,N_11415);
nor U18563 (N_18563,N_12197,N_11481);
nor U18564 (N_18564,N_13512,N_12612);
or U18565 (N_18565,N_14634,N_13963);
nor U18566 (N_18566,N_12943,N_13814);
and U18567 (N_18567,N_14558,N_13926);
xor U18568 (N_18568,N_11426,N_12773);
nand U18569 (N_18569,N_14082,N_10725);
and U18570 (N_18570,N_13770,N_11261);
nand U18571 (N_18571,N_14912,N_13235);
nand U18572 (N_18572,N_11531,N_11173);
xnor U18573 (N_18573,N_10085,N_12270);
or U18574 (N_18574,N_14226,N_12456);
nand U18575 (N_18575,N_13762,N_12990);
nand U18576 (N_18576,N_11651,N_14956);
or U18577 (N_18577,N_12134,N_12538);
and U18578 (N_18578,N_11250,N_13445);
or U18579 (N_18579,N_13290,N_11470);
nand U18580 (N_18580,N_12832,N_14030);
and U18581 (N_18581,N_14116,N_10779);
nor U18582 (N_18582,N_13065,N_13141);
and U18583 (N_18583,N_11179,N_12315);
or U18584 (N_18584,N_13221,N_10100);
nor U18585 (N_18585,N_11641,N_13351);
nand U18586 (N_18586,N_14917,N_13119);
and U18587 (N_18587,N_14555,N_11543);
nor U18588 (N_18588,N_12949,N_12945);
and U18589 (N_18589,N_10056,N_10761);
or U18590 (N_18590,N_13228,N_14389);
nor U18591 (N_18591,N_14594,N_11387);
and U18592 (N_18592,N_12179,N_14956);
nor U18593 (N_18593,N_11475,N_11828);
nand U18594 (N_18594,N_14263,N_11927);
or U18595 (N_18595,N_13178,N_10965);
nand U18596 (N_18596,N_11014,N_14574);
nand U18597 (N_18597,N_10851,N_14012);
nor U18598 (N_18598,N_14243,N_14765);
and U18599 (N_18599,N_10473,N_10140);
and U18600 (N_18600,N_14043,N_10608);
or U18601 (N_18601,N_10457,N_13507);
nand U18602 (N_18602,N_14448,N_10900);
or U18603 (N_18603,N_13095,N_10620);
nor U18604 (N_18604,N_10005,N_11443);
and U18605 (N_18605,N_13217,N_12167);
nor U18606 (N_18606,N_10072,N_12886);
nand U18607 (N_18607,N_10647,N_13997);
and U18608 (N_18608,N_11606,N_13555);
nor U18609 (N_18609,N_11223,N_14876);
nand U18610 (N_18610,N_13034,N_14533);
or U18611 (N_18611,N_14223,N_10036);
nor U18612 (N_18612,N_11063,N_10028);
nor U18613 (N_18613,N_14892,N_13770);
or U18614 (N_18614,N_14710,N_10115);
nor U18615 (N_18615,N_11542,N_12532);
nand U18616 (N_18616,N_14566,N_11873);
xor U18617 (N_18617,N_14038,N_12815);
and U18618 (N_18618,N_12060,N_12687);
or U18619 (N_18619,N_12898,N_14523);
or U18620 (N_18620,N_13719,N_12923);
and U18621 (N_18621,N_10778,N_10457);
nand U18622 (N_18622,N_10631,N_14262);
and U18623 (N_18623,N_11182,N_10881);
or U18624 (N_18624,N_11556,N_11996);
nand U18625 (N_18625,N_14080,N_10096);
nor U18626 (N_18626,N_14641,N_14665);
xor U18627 (N_18627,N_13563,N_10447);
or U18628 (N_18628,N_13647,N_13234);
nand U18629 (N_18629,N_11676,N_12528);
and U18630 (N_18630,N_12858,N_13512);
nand U18631 (N_18631,N_12562,N_13414);
nor U18632 (N_18632,N_10869,N_11290);
nor U18633 (N_18633,N_14387,N_11720);
nand U18634 (N_18634,N_10378,N_14683);
nand U18635 (N_18635,N_14950,N_10766);
or U18636 (N_18636,N_10542,N_13832);
or U18637 (N_18637,N_11156,N_14953);
or U18638 (N_18638,N_14032,N_11814);
xnor U18639 (N_18639,N_13356,N_12247);
and U18640 (N_18640,N_13272,N_13464);
nor U18641 (N_18641,N_11944,N_10102);
and U18642 (N_18642,N_14180,N_14905);
and U18643 (N_18643,N_10345,N_14135);
nand U18644 (N_18644,N_11374,N_11452);
nand U18645 (N_18645,N_12276,N_10813);
xnor U18646 (N_18646,N_13747,N_11133);
or U18647 (N_18647,N_13475,N_12561);
or U18648 (N_18648,N_11566,N_11041);
and U18649 (N_18649,N_11789,N_13568);
nand U18650 (N_18650,N_10130,N_10144);
nand U18651 (N_18651,N_11373,N_13721);
nor U18652 (N_18652,N_14451,N_11887);
and U18653 (N_18653,N_10143,N_11609);
and U18654 (N_18654,N_14485,N_12796);
nand U18655 (N_18655,N_12354,N_11860);
nor U18656 (N_18656,N_12088,N_12856);
or U18657 (N_18657,N_11984,N_13560);
xor U18658 (N_18658,N_12941,N_14731);
and U18659 (N_18659,N_10638,N_12681);
nand U18660 (N_18660,N_14410,N_11297);
xor U18661 (N_18661,N_14101,N_11321);
nand U18662 (N_18662,N_13439,N_14137);
and U18663 (N_18663,N_11579,N_10878);
nor U18664 (N_18664,N_14099,N_14392);
nor U18665 (N_18665,N_11572,N_12517);
or U18666 (N_18666,N_11935,N_12420);
and U18667 (N_18667,N_13488,N_13471);
and U18668 (N_18668,N_12773,N_14890);
and U18669 (N_18669,N_12750,N_12963);
and U18670 (N_18670,N_12583,N_10514);
or U18671 (N_18671,N_12664,N_13506);
nor U18672 (N_18672,N_12966,N_13832);
nor U18673 (N_18673,N_12785,N_12880);
xnor U18674 (N_18674,N_11505,N_12908);
or U18675 (N_18675,N_12803,N_10555);
or U18676 (N_18676,N_14724,N_11549);
xnor U18677 (N_18677,N_12004,N_11699);
or U18678 (N_18678,N_14194,N_14913);
nor U18679 (N_18679,N_14678,N_14773);
and U18680 (N_18680,N_14205,N_13746);
or U18681 (N_18681,N_12281,N_14447);
and U18682 (N_18682,N_12323,N_13226);
nor U18683 (N_18683,N_11271,N_13538);
nand U18684 (N_18684,N_12285,N_14108);
or U18685 (N_18685,N_11589,N_14600);
nand U18686 (N_18686,N_13724,N_14235);
nor U18687 (N_18687,N_14633,N_13999);
and U18688 (N_18688,N_10321,N_11227);
or U18689 (N_18689,N_11608,N_10069);
nor U18690 (N_18690,N_10899,N_12568);
nand U18691 (N_18691,N_10431,N_11286);
nor U18692 (N_18692,N_12863,N_13454);
nor U18693 (N_18693,N_12822,N_12352);
nand U18694 (N_18694,N_12218,N_12167);
xor U18695 (N_18695,N_12637,N_10375);
or U18696 (N_18696,N_11911,N_14064);
nor U18697 (N_18697,N_13241,N_14026);
and U18698 (N_18698,N_13989,N_10660);
nand U18699 (N_18699,N_14396,N_12100);
xor U18700 (N_18700,N_13966,N_12483);
xnor U18701 (N_18701,N_14654,N_11842);
or U18702 (N_18702,N_11467,N_13993);
nor U18703 (N_18703,N_10132,N_10739);
nor U18704 (N_18704,N_12204,N_13598);
nand U18705 (N_18705,N_13368,N_12177);
and U18706 (N_18706,N_14819,N_10082);
or U18707 (N_18707,N_12581,N_14226);
and U18708 (N_18708,N_12448,N_13284);
nor U18709 (N_18709,N_10766,N_10604);
xor U18710 (N_18710,N_12165,N_13615);
nand U18711 (N_18711,N_11309,N_10677);
nand U18712 (N_18712,N_10149,N_11959);
nand U18713 (N_18713,N_14355,N_11898);
nand U18714 (N_18714,N_14349,N_12505);
nor U18715 (N_18715,N_14964,N_10885);
and U18716 (N_18716,N_11896,N_11766);
xnor U18717 (N_18717,N_13760,N_14183);
and U18718 (N_18718,N_13711,N_10738);
or U18719 (N_18719,N_12590,N_14323);
and U18720 (N_18720,N_14744,N_11759);
and U18721 (N_18721,N_10828,N_12544);
nand U18722 (N_18722,N_12054,N_11428);
and U18723 (N_18723,N_14670,N_13240);
nand U18724 (N_18724,N_10126,N_10008);
or U18725 (N_18725,N_14035,N_13988);
xor U18726 (N_18726,N_10645,N_14735);
or U18727 (N_18727,N_11524,N_10017);
nor U18728 (N_18728,N_13512,N_13870);
xnor U18729 (N_18729,N_14800,N_12519);
and U18730 (N_18730,N_12620,N_12921);
nor U18731 (N_18731,N_11142,N_13246);
xor U18732 (N_18732,N_13911,N_12944);
xor U18733 (N_18733,N_13322,N_10250);
nor U18734 (N_18734,N_12015,N_11707);
or U18735 (N_18735,N_13124,N_14679);
or U18736 (N_18736,N_13592,N_10607);
nand U18737 (N_18737,N_14661,N_12711);
nand U18738 (N_18738,N_13491,N_14084);
xnor U18739 (N_18739,N_10806,N_14719);
nand U18740 (N_18740,N_13072,N_12587);
nand U18741 (N_18741,N_12335,N_11065);
nor U18742 (N_18742,N_13664,N_12402);
nand U18743 (N_18743,N_10177,N_12293);
xor U18744 (N_18744,N_14452,N_14141);
and U18745 (N_18745,N_14117,N_13322);
nor U18746 (N_18746,N_13140,N_10397);
nor U18747 (N_18747,N_10071,N_12087);
or U18748 (N_18748,N_10359,N_13347);
or U18749 (N_18749,N_11992,N_12843);
nand U18750 (N_18750,N_12476,N_14174);
or U18751 (N_18751,N_13926,N_12179);
nor U18752 (N_18752,N_12717,N_14986);
or U18753 (N_18753,N_11107,N_14849);
nor U18754 (N_18754,N_10766,N_10520);
or U18755 (N_18755,N_11587,N_12591);
nand U18756 (N_18756,N_11332,N_10933);
or U18757 (N_18757,N_11506,N_13683);
and U18758 (N_18758,N_12861,N_11961);
nor U18759 (N_18759,N_12731,N_14343);
or U18760 (N_18760,N_12679,N_14301);
or U18761 (N_18761,N_12924,N_10691);
nor U18762 (N_18762,N_10966,N_12339);
and U18763 (N_18763,N_11645,N_12619);
nand U18764 (N_18764,N_11914,N_14109);
nand U18765 (N_18765,N_12816,N_10617);
xnor U18766 (N_18766,N_11006,N_12393);
nand U18767 (N_18767,N_12380,N_11989);
and U18768 (N_18768,N_10809,N_14608);
xor U18769 (N_18769,N_12795,N_11838);
nand U18770 (N_18770,N_13581,N_11846);
and U18771 (N_18771,N_11652,N_12145);
and U18772 (N_18772,N_14289,N_14658);
and U18773 (N_18773,N_14733,N_13018);
nor U18774 (N_18774,N_12443,N_14895);
or U18775 (N_18775,N_11040,N_11385);
and U18776 (N_18776,N_12459,N_12260);
or U18777 (N_18777,N_13716,N_12625);
and U18778 (N_18778,N_10183,N_14086);
xor U18779 (N_18779,N_13620,N_12992);
nor U18780 (N_18780,N_14806,N_10302);
and U18781 (N_18781,N_13948,N_11266);
or U18782 (N_18782,N_11674,N_10509);
nor U18783 (N_18783,N_11790,N_13961);
xor U18784 (N_18784,N_12712,N_14009);
nand U18785 (N_18785,N_11300,N_11067);
and U18786 (N_18786,N_11452,N_14784);
xnor U18787 (N_18787,N_14904,N_14552);
and U18788 (N_18788,N_14413,N_11723);
nor U18789 (N_18789,N_14692,N_11076);
xnor U18790 (N_18790,N_14548,N_12825);
or U18791 (N_18791,N_11860,N_14776);
and U18792 (N_18792,N_11339,N_10994);
and U18793 (N_18793,N_14315,N_14377);
and U18794 (N_18794,N_13168,N_11332);
and U18795 (N_18795,N_11544,N_12025);
and U18796 (N_18796,N_12003,N_11413);
and U18797 (N_18797,N_12192,N_10808);
or U18798 (N_18798,N_14056,N_12650);
and U18799 (N_18799,N_10599,N_11571);
or U18800 (N_18800,N_11731,N_13750);
nor U18801 (N_18801,N_14884,N_12150);
nand U18802 (N_18802,N_11487,N_13030);
and U18803 (N_18803,N_13207,N_10314);
or U18804 (N_18804,N_12558,N_13186);
xnor U18805 (N_18805,N_12982,N_13471);
xor U18806 (N_18806,N_12102,N_14469);
nand U18807 (N_18807,N_11689,N_14705);
xnor U18808 (N_18808,N_12322,N_12487);
xor U18809 (N_18809,N_13174,N_12519);
nand U18810 (N_18810,N_11931,N_11605);
nand U18811 (N_18811,N_11029,N_14825);
xnor U18812 (N_18812,N_10200,N_13967);
nand U18813 (N_18813,N_10814,N_12632);
and U18814 (N_18814,N_13313,N_11865);
and U18815 (N_18815,N_13446,N_10057);
nor U18816 (N_18816,N_11940,N_13949);
nand U18817 (N_18817,N_12288,N_12392);
nand U18818 (N_18818,N_14508,N_13365);
or U18819 (N_18819,N_10970,N_11449);
and U18820 (N_18820,N_11001,N_10072);
nand U18821 (N_18821,N_10711,N_14023);
and U18822 (N_18822,N_13593,N_14251);
and U18823 (N_18823,N_13446,N_12011);
or U18824 (N_18824,N_12113,N_10741);
nand U18825 (N_18825,N_14105,N_14430);
or U18826 (N_18826,N_13835,N_14031);
and U18827 (N_18827,N_14063,N_12813);
nor U18828 (N_18828,N_11072,N_11867);
or U18829 (N_18829,N_13762,N_14214);
and U18830 (N_18830,N_13568,N_11077);
xor U18831 (N_18831,N_13354,N_12485);
nand U18832 (N_18832,N_11918,N_11880);
nand U18833 (N_18833,N_13504,N_14833);
nand U18834 (N_18834,N_11798,N_10716);
nand U18835 (N_18835,N_13697,N_14468);
xor U18836 (N_18836,N_10497,N_10381);
or U18837 (N_18837,N_12650,N_13706);
or U18838 (N_18838,N_13791,N_12628);
xnor U18839 (N_18839,N_11952,N_14288);
or U18840 (N_18840,N_11608,N_12709);
nand U18841 (N_18841,N_14573,N_12524);
nor U18842 (N_18842,N_10944,N_12424);
nand U18843 (N_18843,N_11856,N_12923);
and U18844 (N_18844,N_12545,N_11088);
nand U18845 (N_18845,N_13055,N_13521);
or U18846 (N_18846,N_14140,N_13425);
nor U18847 (N_18847,N_11917,N_13898);
xnor U18848 (N_18848,N_10720,N_14788);
and U18849 (N_18849,N_10441,N_11324);
and U18850 (N_18850,N_10748,N_13774);
and U18851 (N_18851,N_12658,N_14674);
or U18852 (N_18852,N_11719,N_13449);
or U18853 (N_18853,N_11244,N_13588);
and U18854 (N_18854,N_11728,N_11946);
or U18855 (N_18855,N_13725,N_12619);
or U18856 (N_18856,N_14414,N_10268);
and U18857 (N_18857,N_14036,N_11903);
nand U18858 (N_18858,N_13381,N_12818);
and U18859 (N_18859,N_14004,N_10425);
nand U18860 (N_18860,N_11988,N_13489);
and U18861 (N_18861,N_11905,N_10281);
and U18862 (N_18862,N_14895,N_12235);
nand U18863 (N_18863,N_10880,N_14289);
nand U18864 (N_18864,N_13556,N_13275);
or U18865 (N_18865,N_10556,N_13270);
nor U18866 (N_18866,N_13744,N_13652);
and U18867 (N_18867,N_13268,N_12396);
or U18868 (N_18868,N_14265,N_10948);
xor U18869 (N_18869,N_12544,N_14550);
or U18870 (N_18870,N_14786,N_11944);
nand U18871 (N_18871,N_10279,N_10712);
xnor U18872 (N_18872,N_13132,N_14726);
and U18873 (N_18873,N_14471,N_13295);
xnor U18874 (N_18874,N_10047,N_13763);
or U18875 (N_18875,N_13538,N_14999);
or U18876 (N_18876,N_11875,N_14292);
nor U18877 (N_18877,N_13041,N_12123);
or U18878 (N_18878,N_12469,N_10192);
nor U18879 (N_18879,N_11340,N_11281);
nor U18880 (N_18880,N_13928,N_13730);
xnor U18881 (N_18881,N_14538,N_10323);
or U18882 (N_18882,N_11551,N_14410);
and U18883 (N_18883,N_10792,N_11630);
nand U18884 (N_18884,N_13109,N_14526);
nor U18885 (N_18885,N_14261,N_14458);
nor U18886 (N_18886,N_13929,N_12461);
nor U18887 (N_18887,N_10725,N_13106);
nor U18888 (N_18888,N_14969,N_12271);
nor U18889 (N_18889,N_11010,N_13449);
or U18890 (N_18890,N_10258,N_11417);
nand U18891 (N_18891,N_12897,N_13916);
and U18892 (N_18892,N_14405,N_11139);
nor U18893 (N_18893,N_10578,N_12267);
and U18894 (N_18894,N_14787,N_14911);
and U18895 (N_18895,N_13720,N_11382);
and U18896 (N_18896,N_13305,N_12049);
nor U18897 (N_18897,N_14639,N_11512);
xor U18898 (N_18898,N_13098,N_12769);
and U18899 (N_18899,N_13584,N_12266);
or U18900 (N_18900,N_12287,N_13788);
or U18901 (N_18901,N_11816,N_11527);
and U18902 (N_18902,N_10610,N_10310);
or U18903 (N_18903,N_13581,N_12300);
nand U18904 (N_18904,N_11496,N_13088);
xor U18905 (N_18905,N_12953,N_10508);
nor U18906 (N_18906,N_12720,N_12016);
nand U18907 (N_18907,N_14251,N_12010);
and U18908 (N_18908,N_10863,N_11195);
nor U18909 (N_18909,N_10886,N_13464);
nand U18910 (N_18910,N_13537,N_12642);
xnor U18911 (N_18911,N_13275,N_11382);
and U18912 (N_18912,N_11836,N_10070);
nor U18913 (N_18913,N_10960,N_14526);
nand U18914 (N_18914,N_10163,N_12815);
or U18915 (N_18915,N_12420,N_10178);
and U18916 (N_18916,N_13387,N_13107);
and U18917 (N_18917,N_11137,N_13301);
nand U18918 (N_18918,N_10811,N_12678);
nor U18919 (N_18919,N_11159,N_14086);
or U18920 (N_18920,N_12891,N_10302);
nand U18921 (N_18921,N_12703,N_14702);
nand U18922 (N_18922,N_13554,N_14348);
nand U18923 (N_18923,N_10878,N_10239);
nand U18924 (N_18924,N_10106,N_11180);
xnor U18925 (N_18925,N_14389,N_11075);
nor U18926 (N_18926,N_12088,N_13894);
and U18927 (N_18927,N_14793,N_14480);
nor U18928 (N_18928,N_13441,N_14743);
or U18929 (N_18929,N_14426,N_13816);
or U18930 (N_18930,N_12930,N_12500);
nor U18931 (N_18931,N_11683,N_13080);
or U18932 (N_18932,N_13249,N_11565);
or U18933 (N_18933,N_13253,N_10286);
and U18934 (N_18934,N_14610,N_12491);
nand U18935 (N_18935,N_13995,N_13207);
and U18936 (N_18936,N_10926,N_11310);
and U18937 (N_18937,N_12426,N_10184);
and U18938 (N_18938,N_10834,N_11589);
nor U18939 (N_18939,N_13773,N_10826);
and U18940 (N_18940,N_13785,N_14031);
nor U18941 (N_18941,N_13653,N_14187);
xor U18942 (N_18942,N_10293,N_12406);
or U18943 (N_18943,N_14666,N_10376);
nor U18944 (N_18944,N_13240,N_12131);
or U18945 (N_18945,N_13311,N_13011);
nor U18946 (N_18946,N_12931,N_14020);
or U18947 (N_18947,N_14382,N_10302);
nand U18948 (N_18948,N_13302,N_10975);
or U18949 (N_18949,N_13003,N_12435);
and U18950 (N_18950,N_14247,N_13087);
nand U18951 (N_18951,N_11535,N_11464);
nor U18952 (N_18952,N_14133,N_13354);
or U18953 (N_18953,N_11635,N_14064);
nor U18954 (N_18954,N_12083,N_12971);
or U18955 (N_18955,N_12273,N_11809);
and U18956 (N_18956,N_11453,N_12048);
nor U18957 (N_18957,N_14482,N_11907);
nand U18958 (N_18958,N_10526,N_10619);
nor U18959 (N_18959,N_14938,N_14554);
nor U18960 (N_18960,N_13149,N_11232);
nand U18961 (N_18961,N_11694,N_11040);
and U18962 (N_18962,N_10872,N_13294);
or U18963 (N_18963,N_14658,N_11455);
nand U18964 (N_18964,N_10933,N_13859);
or U18965 (N_18965,N_13769,N_14986);
and U18966 (N_18966,N_12771,N_13379);
xor U18967 (N_18967,N_12675,N_14666);
and U18968 (N_18968,N_10335,N_10478);
nor U18969 (N_18969,N_11725,N_13607);
nor U18970 (N_18970,N_12749,N_10095);
and U18971 (N_18971,N_14666,N_13229);
or U18972 (N_18972,N_12078,N_10852);
nand U18973 (N_18973,N_14065,N_12755);
and U18974 (N_18974,N_12954,N_13248);
nand U18975 (N_18975,N_11074,N_11499);
and U18976 (N_18976,N_14869,N_14891);
or U18977 (N_18977,N_14701,N_12864);
nand U18978 (N_18978,N_13220,N_12758);
nand U18979 (N_18979,N_13727,N_13085);
and U18980 (N_18980,N_11312,N_12943);
or U18981 (N_18981,N_14351,N_11166);
nor U18982 (N_18982,N_11545,N_11396);
xnor U18983 (N_18983,N_11542,N_12628);
and U18984 (N_18984,N_10132,N_14123);
nor U18985 (N_18985,N_12094,N_11246);
or U18986 (N_18986,N_10493,N_11436);
and U18987 (N_18987,N_10359,N_13585);
nand U18988 (N_18988,N_12913,N_10298);
nor U18989 (N_18989,N_14153,N_14923);
nand U18990 (N_18990,N_10992,N_13672);
and U18991 (N_18991,N_12899,N_12312);
nand U18992 (N_18992,N_11199,N_14841);
nand U18993 (N_18993,N_14437,N_12524);
or U18994 (N_18994,N_11031,N_14760);
or U18995 (N_18995,N_12850,N_14673);
nand U18996 (N_18996,N_11310,N_14480);
or U18997 (N_18997,N_14965,N_10496);
nand U18998 (N_18998,N_12865,N_11602);
nand U18999 (N_18999,N_12763,N_10994);
nand U19000 (N_19000,N_11103,N_13466);
nand U19001 (N_19001,N_11761,N_13926);
or U19002 (N_19002,N_13964,N_13650);
or U19003 (N_19003,N_10006,N_12159);
nor U19004 (N_19004,N_12425,N_12492);
nor U19005 (N_19005,N_11687,N_10349);
nor U19006 (N_19006,N_14809,N_13471);
nor U19007 (N_19007,N_12390,N_13772);
or U19008 (N_19008,N_12465,N_11632);
and U19009 (N_19009,N_11432,N_14886);
nor U19010 (N_19010,N_12235,N_12904);
xor U19011 (N_19011,N_14143,N_10397);
nor U19012 (N_19012,N_10183,N_14122);
nor U19013 (N_19013,N_13346,N_14028);
and U19014 (N_19014,N_10038,N_10949);
nand U19015 (N_19015,N_11061,N_13112);
and U19016 (N_19016,N_13293,N_11684);
xor U19017 (N_19017,N_13027,N_14488);
xnor U19018 (N_19018,N_12344,N_12044);
nor U19019 (N_19019,N_12934,N_10301);
and U19020 (N_19020,N_10840,N_10481);
and U19021 (N_19021,N_14705,N_14108);
or U19022 (N_19022,N_14536,N_10379);
or U19023 (N_19023,N_12399,N_14241);
or U19024 (N_19024,N_14361,N_10321);
nor U19025 (N_19025,N_11155,N_13778);
nor U19026 (N_19026,N_12305,N_11463);
nor U19027 (N_19027,N_12569,N_13915);
or U19028 (N_19028,N_10484,N_14989);
xnor U19029 (N_19029,N_12618,N_13649);
or U19030 (N_19030,N_12795,N_10921);
nand U19031 (N_19031,N_13948,N_11884);
nand U19032 (N_19032,N_10451,N_14432);
or U19033 (N_19033,N_10954,N_12707);
or U19034 (N_19034,N_11340,N_14281);
nand U19035 (N_19035,N_10537,N_13926);
nand U19036 (N_19036,N_11418,N_10959);
nor U19037 (N_19037,N_12134,N_13943);
or U19038 (N_19038,N_10586,N_11742);
nand U19039 (N_19039,N_13712,N_13782);
and U19040 (N_19040,N_12029,N_11066);
xor U19041 (N_19041,N_14572,N_11650);
or U19042 (N_19042,N_14537,N_12695);
and U19043 (N_19043,N_10486,N_11823);
nor U19044 (N_19044,N_10182,N_11164);
nand U19045 (N_19045,N_11807,N_14348);
or U19046 (N_19046,N_11501,N_13422);
and U19047 (N_19047,N_10390,N_11767);
or U19048 (N_19048,N_13093,N_14978);
xor U19049 (N_19049,N_12183,N_12424);
nand U19050 (N_19050,N_14570,N_14750);
xnor U19051 (N_19051,N_13312,N_10597);
and U19052 (N_19052,N_14066,N_13300);
nand U19053 (N_19053,N_13327,N_11952);
nand U19054 (N_19054,N_14460,N_14721);
or U19055 (N_19055,N_14357,N_14609);
or U19056 (N_19056,N_10037,N_14491);
or U19057 (N_19057,N_12245,N_12712);
nand U19058 (N_19058,N_13490,N_12495);
nand U19059 (N_19059,N_14328,N_11058);
nand U19060 (N_19060,N_11475,N_13873);
or U19061 (N_19061,N_11875,N_10889);
xnor U19062 (N_19062,N_14658,N_10276);
nor U19063 (N_19063,N_10101,N_13471);
nand U19064 (N_19064,N_10796,N_11233);
nor U19065 (N_19065,N_10499,N_13110);
and U19066 (N_19066,N_13930,N_10428);
and U19067 (N_19067,N_12474,N_14638);
and U19068 (N_19068,N_10000,N_12205);
nand U19069 (N_19069,N_11808,N_14648);
nor U19070 (N_19070,N_11241,N_11821);
xnor U19071 (N_19071,N_14705,N_12011);
nand U19072 (N_19072,N_12954,N_12742);
or U19073 (N_19073,N_12692,N_14484);
xnor U19074 (N_19074,N_14314,N_12945);
and U19075 (N_19075,N_14712,N_12772);
and U19076 (N_19076,N_12006,N_10407);
or U19077 (N_19077,N_13480,N_10984);
nand U19078 (N_19078,N_12357,N_13389);
and U19079 (N_19079,N_13265,N_12187);
nor U19080 (N_19080,N_12009,N_10090);
nor U19081 (N_19081,N_13958,N_14478);
or U19082 (N_19082,N_12764,N_13397);
and U19083 (N_19083,N_12937,N_10229);
nor U19084 (N_19084,N_11374,N_12612);
or U19085 (N_19085,N_10935,N_11309);
nand U19086 (N_19086,N_10312,N_13178);
nand U19087 (N_19087,N_12469,N_14573);
and U19088 (N_19088,N_12705,N_13541);
nand U19089 (N_19089,N_12515,N_14259);
nand U19090 (N_19090,N_11120,N_14559);
or U19091 (N_19091,N_14914,N_11656);
or U19092 (N_19092,N_11030,N_10679);
nand U19093 (N_19093,N_13114,N_11480);
and U19094 (N_19094,N_14861,N_12281);
or U19095 (N_19095,N_11702,N_10070);
nand U19096 (N_19096,N_11505,N_12682);
and U19097 (N_19097,N_13074,N_11941);
nand U19098 (N_19098,N_12024,N_10442);
nand U19099 (N_19099,N_13054,N_12886);
nor U19100 (N_19100,N_14671,N_13497);
and U19101 (N_19101,N_12209,N_11304);
and U19102 (N_19102,N_12826,N_11251);
nor U19103 (N_19103,N_12823,N_11505);
nand U19104 (N_19104,N_14470,N_11536);
nor U19105 (N_19105,N_11819,N_12517);
and U19106 (N_19106,N_10791,N_14069);
or U19107 (N_19107,N_14789,N_10121);
or U19108 (N_19108,N_13397,N_10585);
nor U19109 (N_19109,N_10805,N_11279);
nor U19110 (N_19110,N_13506,N_14867);
nor U19111 (N_19111,N_11332,N_11974);
or U19112 (N_19112,N_14686,N_13758);
and U19113 (N_19113,N_10340,N_10703);
nand U19114 (N_19114,N_12737,N_11233);
and U19115 (N_19115,N_11097,N_10157);
or U19116 (N_19116,N_11716,N_11497);
or U19117 (N_19117,N_14953,N_12746);
nand U19118 (N_19118,N_13292,N_12426);
or U19119 (N_19119,N_14266,N_10160);
nor U19120 (N_19120,N_13462,N_13471);
nand U19121 (N_19121,N_13636,N_13645);
nand U19122 (N_19122,N_14915,N_11254);
or U19123 (N_19123,N_13817,N_13416);
nor U19124 (N_19124,N_10225,N_13593);
nor U19125 (N_19125,N_13277,N_14102);
and U19126 (N_19126,N_12623,N_11142);
nor U19127 (N_19127,N_13541,N_14810);
or U19128 (N_19128,N_10726,N_13358);
and U19129 (N_19129,N_14403,N_11388);
and U19130 (N_19130,N_11895,N_11556);
nor U19131 (N_19131,N_10804,N_11471);
nand U19132 (N_19132,N_11477,N_13283);
nand U19133 (N_19133,N_12823,N_10452);
and U19134 (N_19134,N_14974,N_11327);
xor U19135 (N_19135,N_11815,N_11122);
nand U19136 (N_19136,N_10391,N_12900);
or U19137 (N_19137,N_10560,N_11106);
nor U19138 (N_19138,N_13228,N_13008);
xnor U19139 (N_19139,N_11567,N_10156);
xnor U19140 (N_19140,N_12683,N_11900);
or U19141 (N_19141,N_12045,N_13076);
nor U19142 (N_19142,N_11395,N_11759);
or U19143 (N_19143,N_10370,N_10720);
nand U19144 (N_19144,N_12338,N_10507);
and U19145 (N_19145,N_11301,N_12562);
nor U19146 (N_19146,N_11843,N_12530);
or U19147 (N_19147,N_11965,N_14719);
nor U19148 (N_19148,N_11796,N_14403);
nor U19149 (N_19149,N_14892,N_11740);
nand U19150 (N_19150,N_10747,N_14746);
and U19151 (N_19151,N_10596,N_14118);
nor U19152 (N_19152,N_10543,N_14861);
xnor U19153 (N_19153,N_13337,N_12221);
nor U19154 (N_19154,N_10229,N_13351);
and U19155 (N_19155,N_10155,N_12143);
nand U19156 (N_19156,N_11175,N_12026);
nor U19157 (N_19157,N_10518,N_14526);
and U19158 (N_19158,N_11715,N_10537);
nor U19159 (N_19159,N_11451,N_12490);
nand U19160 (N_19160,N_11455,N_10837);
nand U19161 (N_19161,N_10570,N_14215);
and U19162 (N_19162,N_12518,N_10840);
nor U19163 (N_19163,N_14126,N_14597);
nor U19164 (N_19164,N_12748,N_11645);
nand U19165 (N_19165,N_12488,N_13615);
nor U19166 (N_19166,N_14970,N_12920);
nor U19167 (N_19167,N_11003,N_12648);
or U19168 (N_19168,N_14817,N_14310);
nor U19169 (N_19169,N_10375,N_10634);
nor U19170 (N_19170,N_14152,N_13599);
nand U19171 (N_19171,N_11438,N_12811);
nor U19172 (N_19172,N_11895,N_11637);
and U19173 (N_19173,N_12255,N_11616);
nand U19174 (N_19174,N_14349,N_11310);
nor U19175 (N_19175,N_10416,N_12195);
nand U19176 (N_19176,N_12937,N_12128);
nor U19177 (N_19177,N_13281,N_13145);
nor U19178 (N_19178,N_12062,N_11942);
nor U19179 (N_19179,N_13349,N_10955);
xor U19180 (N_19180,N_14852,N_10741);
xor U19181 (N_19181,N_10797,N_14096);
and U19182 (N_19182,N_13175,N_14655);
nor U19183 (N_19183,N_11737,N_13639);
and U19184 (N_19184,N_13311,N_14430);
nand U19185 (N_19185,N_13612,N_13724);
nor U19186 (N_19186,N_12299,N_11390);
and U19187 (N_19187,N_11147,N_12220);
nor U19188 (N_19188,N_10429,N_14916);
nor U19189 (N_19189,N_14740,N_12871);
or U19190 (N_19190,N_12523,N_12580);
and U19191 (N_19191,N_10034,N_11378);
xor U19192 (N_19192,N_13723,N_12583);
nand U19193 (N_19193,N_12903,N_11714);
xor U19194 (N_19194,N_14429,N_14192);
nand U19195 (N_19195,N_10426,N_13165);
xor U19196 (N_19196,N_13653,N_13507);
nand U19197 (N_19197,N_12934,N_14377);
nand U19198 (N_19198,N_11221,N_12186);
or U19199 (N_19199,N_14758,N_13359);
nor U19200 (N_19200,N_12559,N_12793);
nor U19201 (N_19201,N_10059,N_10303);
nand U19202 (N_19202,N_11233,N_13011);
nor U19203 (N_19203,N_10219,N_14471);
or U19204 (N_19204,N_13810,N_12573);
and U19205 (N_19205,N_10270,N_13420);
nor U19206 (N_19206,N_14284,N_13347);
or U19207 (N_19207,N_12410,N_13155);
and U19208 (N_19208,N_14383,N_10389);
nand U19209 (N_19209,N_13960,N_10932);
and U19210 (N_19210,N_11837,N_13242);
or U19211 (N_19211,N_13040,N_12514);
nor U19212 (N_19212,N_11190,N_10035);
or U19213 (N_19213,N_14848,N_11872);
xnor U19214 (N_19214,N_11870,N_10346);
and U19215 (N_19215,N_11058,N_10903);
nor U19216 (N_19216,N_14027,N_10028);
nand U19217 (N_19217,N_10568,N_13907);
nor U19218 (N_19218,N_10372,N_10028);
nand U19219 (N_19219,N_13278,N_12239);
and U19220 (N_19220,N_13610,N_10095);
xnor U19221 (N_19221,N_10391,N_10527);
nor U19222 (N_19222,N_13559,N_11718);
or U19223 (N_19223,N_13258,N_12741);
nand U19224 (N_19224,N_12186,N_12812);
nor U19225 (N_19225,N_10428,N_14074);
or U19226 (N_19226,N_12962,N_11227);
and U19227 (N_19227,N_13038,N_12537);
and U19228 (N_19228,N_13679,N_12436);
or U19229 (N_19229,N_12166,N_14293);
or U19230 (N_19230,N_14396,N_11562);
nor U19231 (N_19231,N_10836,N_11971);
or U19232 (N_19232,N_12571,N_12092);
nor U19233 (N_19233,N_14673,N_13020);
or U19234 (N_19234,N_14847,N_14914);
or U19235 (N_19235,N_12712,N_11979);
nor U19236 (N_19236,N_14967,N_14193);
and U19237 (N_19237,N_12849,N_12839);
xnor U19238 (N_19238,N_10395,N_11156);
nand U19239 (N_19239,N_10845,N_10355);
and U19240 (N_19240,N_14119,N_10142);
or U19241 (N_19241,N_12854,N_14241);
nand U19242 (N_19242,N_13579,N_14130);
nor U19243 (N_19243,N_12222,N_12078);
nor U19244 (N_19244,N_12959,N_10156);
or U19245 (N_19245,N_13629,N_13438);
or U19246 (N_19246,N_12252,N_10092);
nor U19247 (N_19247,N_14014,N_14756);
nor U19248 (N_19248,N_14604,N_12005);
nand U19249 (N_19249,N_13274,N_10041);
nand U19250 (N_19250,N_12990,N_11813);
nand U19251 (N_19251,N_11700,N_13592);
xnor U19252 (N_19252,N_13568,N_13391);
or U19253 (N_19253,N_14057,N_13322);
xor U19254 (N_19254,N_10573,N_10152);
nor U19255 (N_19255,N_11722,N_12622);
xnor U19256 (N_19256,N_12078,N_11572);
and U19257 (N_19257,N_14707,N_12408);
or U19258 (N_19258,N_11710,N_10898);
nor U19259 (N_19259,N_10446,N_13235);
xnor U19260 (N_19260,N_13566,N_14839);
or U19261 (N_19261,N_10496,N_12994);
nand U19262 (N_19262,N_13694,N_12125);
and U19263 (N_19263,N_14554,N_10389);
nand U19264 (N_19264,N_11959,N_13300);
and U19265 (N_19265,N_10428,N_10661);
xnor U19266 (N_19266,N_14748,N_13138);
nand U19267 (N_19267,N_12103,N_14416);
or U19268 (N_19268,N_11563,N_12790);
nor U19269 (N_19269,N_14458,N_11782);
or U19270 (N_19270,N_11606,N_12987);
nand U19271 (N_19271,N_13902,N_13562);
or U19272 (N_19272,N_10812,N_12025);
or U19273 (N_19273,N_14488,N_13518);
and U19274 (N_19274,N_11894,N_10508);
or U19275 (N_19275,N_10400,N_12746);
and U19276 (N_19276,N_14963,N_10810);
and U19277 (N_19277,N_14773,N_10340);
nand U19278 (N_19278,N_14943,N_14331);
and U19279 (N_19279,N_14673,N_13144);
nand U19280 (N_19280,N_12159,N_12722);
nand U19281 (N_19281,N_14434,N_11716);
and U19282 (N_19282,N_12244,N_10110);
or U19283 (N_19283,N_12854,N_12670);
and U19284 (N_19284,N_14761,N_10067);
and U19285 (N_19285,N_13619,N_13004);
or U19286 (N_19286,N_11897,N_14852);
nor U19287 (N_19287,N_14042,N_14612);
or U19288 (N_19288,N_11227,N_11884);
xnor U19289 (N_19289,N_12697,N_10402);
nand U19290 (N_19290,N_14661,N_12935);
or U19291 (N_19291,N_12913,N_12512);
nand U19292 (N_19292,N_11202,N_12994);
nor U19293 (N_19293,N_13367,N_13501);
nor U19294 (N_19294,N_10874,N_10195);
xor U19295 (N_19295,N_14642,N_14249);
and U19296 (N_19296,N_12419,N_10698);
xor U19297 (N_19297,N_11256,N_14058);
xnor U19298 (N_19298,N_13156,N_11326);
or U19299 (N_19299,N_14280,N_14240);
or U19300 (N_19300,N_14135,N_14945);
and U19301 (N_19301,N_10377,N_13486);
or U19302 (N_19302,N_14607,N_14018);
nor U19303 (N_19303,N_11052,N_11380);
xnor U19304 (N_19304,N_12588,N_11546);
nor U19305 (N_19305,N_12281,N_11315);
and U19306 (N_19306,N_14912,N_10294);
nor U19307 (N_19307,N_14671,N_11052);
nor U19308 (N_19308,N_11198,N_10907);
xnor U19309 (N_19309,N_12166,N_11096);
and U19310 (N_19310,N_10416,N_12443);
or U19311 (N_19311,N_12619,N_13772);
or U19312 (N_19312,N_10496,N_11429);
or U19313 (N_19313,N_11405,N_11173);
or U19314 (N_19314,N_12045,N_14015);
or U19315 (N_19315,N_13009,N_14535);
or U19316 (N_19316,N_10907,N_14586);
xor U19317 (N_19317,N_13170,N_14286);
or U19318 (N_19318,N_10482,N_14723);
nand U19319 (N_19319,N_13294,N_13097);
and U19320 (N_19320,N_11206,N_10424);
nand U19321 (N_19321,N_10218,N_11554);
xor U19322 (N_19322,N_14512,N_14670);
or U19323 (N_19323,N_12983,N_14485);
nand U19324 (N_19324,N_11621,N_14921);
or U19325 (N_19325,N_12456,N_11490);
nand U19326 (N_19326,N_12502,N_14271);
nor U19327 (N_19327,N_14417,N_12089);
nand U19328 (N_19328,N_10096,N_10172);
and U19329 (N_19329,N_13068,N_14745);
nand U19330 (N_19330,N_10233,N_13755);
or U19331 (N_19331,N_14213,N_11782);
nand U19332 (N_19332,N_12870,N_11803);
or U19333 (N_19333,N_11936,N_12659);
xor U19334 (N_19334,N_12266,N_13660);
and U19335 (N_19335,N_10793,N_13670);
or U19336 (N_19336,N_11933,N_13577);
and U19337 (N_19337,N_12765,N_10362);
xnor U19338 (N_19338,N_10032,N_12438);
xor U19339 (N_19339,N_12670,N_14742);
and U19340 (N_19340,N_10096,N_12503);
and U19341 (N_19341,N_11078,N_14338);
xnor U19342 (N_19342,N_14791,N_13593);
nor U19343 (N_19343,N_12027,N_11182);
or U19344 (N_19344,N_14697,N_11684);
and U19345 (N_19345,N_14357,N_13742);
nor U19346 (N_19346,N_10244,N_11491);
and U19347 (N_19347,N_14886,N_10829);
nand U19348 (N_19348,N_11752,N_13499);
xor U19349 (N_19349,N_12284,N_14616);
nor U19350 (N_19350,N_13882,N_10507);
nand U19351 (N_19351,N_12232,N_10962);
nor U19352 (N_19352,N_14752,N_12661);
nor U19353 (N_19353,N_14257,N_11762);
nor U19354 (N_19354,N_14233,N_14422);
or U19355 (N_19355,N_11528,N_11060);
or U19356 (N_19356,N_10342,N_12321);
or U19357 (N_19357,N_13476,N_14552);
nor U19358 (N_19358,N_12234,N_10524);
nand U19359 (N_19359,N_11639,N_13664);
nand U19360 (N_19360,N_10724,N_13094);
or U19361 (N_19361,N_14672,N_11629);
nor U19362 (N_19362,N_13031,N_10417);
nor U19363 (N_19363,N_10200,N_13470);
nor U19364 (N_19364,N_14098,N_13827);
xnor U19365 (N_19365,N_10661,N_10041);
xnor U19366 (N_19366,N_12716,N_14049);
or U19367 (N_19367,N_11006,N_10130);
and U19368 (N_19368,N_12851,N_10428);
nor U19369 (N_19369,N_12379,N_14700);
or U19370 (N_19370,N_13245,N_13372);
or U19371 (N_19371,N_13620,N_13179);
or U19372 (N_19372,N_12412,N_13637);
nor U19373 (N_19373,N_12044,N_13907);
nand U19374 (N_19374,N_12823,N_10623);
nand U19375 (N_19375,N_11436,N_12674);
or U19376 (N_19376,N_11765,N_12035);
nor U19377 (N_19377,N_14380,N_14541);
or U19378 (N_19378,N_13386,N_14061);
nand U19379 (N_19379,N_11452,N_12504);
xnor U19380 (N_19380,N_14446,N_12373);
or U19381 (N_19381,N_13786,N_14007);
nand U19382 (N_19382,N_10206,N_11300);
xnor U19383 (N_19383,N_14620,N_14998);
or U19384 (N_19384,N_13552,N_12370);
nand U19385 (N_19385,N_13151,N_14247);
nand U19386 (N_19386,N_10960,N_14883);
nand U19387 (N_19387,N_13105,N_12247);
and U19388 (N_19388,N_14378,N_10914);
nor U19389 (N_19389,N_11179,N_12913);
nor U19390 (N_19390,N_14190,N_11775);
nand U19391 (N_19391,N_12466,N_13054);
and U19392 (N_19392,N_14353,N_10402);
and U19393 (N_19393,N_13808,N_12723);
nor U19394 (N_19394,N_12726,N_14179);
or U19395 (N_19395,N_13882,N_10760);
nor U19396 (N_19396,N_12689,N_14917);
nand U19397 (N_19397,N_13722,N_12623);
or U19398 (N_19398,N_12155,N_13947);
nand U19399 (N_19399,N_10845,N_12081);
and U19400 (N_19400,N_13028,N_11070);
or U19401 (N_19401,N_10090,N_11668);
nor U19402 (N_19402,N_11989,N_11896);
and U19403 (N_19403,N_13180,N_11237);
or U19404 (N_19404,N_11551,N_14771);
nor U19405 (N_19405,N_12632,N_14703);
nand U19406 (N_19406,N_13159,N_12265);
nand U19407 (N_19407,N_13356,N_13512);
nor U19408 (N_19408,N_12142,N_14609);
or U19409 (N_19409,N_14419,N_14629);
and U19410 (N_19410,N_11160,N_14789);
or U19411 (N_19411,N_14307,N_13764);
or U19412 (N_19412,N_12269,N_13540);
and U19413 (N_19413,N_10047,N_13147);
or U19414 (N_19414,N_10199,N_11512);
nor U19415 (N_19415,N_12088,N_10825);
nand U19416 (N_19416,N_11184,N_11300);
and U19417 (N_19417,N_11472,N_13015);
nand U19418 (N_19418,N_14371,N_11840);
and U19419 (N_19419,N_12774,N_14483);
or U19420 (N_19420,N_13600,N_10710);
nand U19421 (N_19421,N_14063,N_12113);
nor U19422 (N_19422,N_11918,N_12185);
xor U19423 (N_19423,N_11621,N_10013);
nand U19424 (N_19424,N_14877,N_14719);
nor U19425 (N_19425,N_12400,N_13148);
xnor U19426 (N_19426,N_12725,N_11045);
nor U19427 (N_19427,N_11319,N_12286);
or U19428 (N_19428,N_14087,N_10326);
nor U19429 (N_19429,N_14899,N_12749);
nand U19430 (N_19430,N_11094,N_13100);
or U19431 (N_19431,N_13152,N_14010);
or U19432 (N_19432,N_13107,N_11219);
nand U19433 (N_19433,N_12938,N_13690);
and U19434 (N_19434,N_10328,N_12260);
nor U19435 (N_19435,N_11153,N_12122);
nor U19436 (N_19436,N_10992,N_12220);
and U19437 (N_19437,N_10294,N_11032);
or U19438 (N_19438,N_11882,N_13713);
and U19439 (N_19439,N_14302,N_14681);
and U19440 (N_19440,N_13739,N_10333);
nor U19441 (N_19441,N_14872,N_13102);
nand U19442 (N_19442,N_13457,N_11729);
nand U19443 (N_19443,N_12058,N_13297);
nor U19444 (N_19444,N_12558,N_12696);
and U19445 (N_19445,N_14843,N_11185);
and U19446 (N_19446,N_10449,N_13720);
or U19447 (N_19447,N_13718,N_11299);
nor U19448 (N_19448,N_14735,N_12713);
or U19449 (N_19449,N_13633,N_10309);
and U19450 (N_19450,N_14948,N_11833);
nor U19451 (N_19451,N_13561,N_10606);
nand U19452 (N_19452,N_12321,N_12933);
xor U19453 (N_19453,N_13081,N_13907);
and U19454 (N_19454,N_12600,N_10500);
or U19455 (N_19455,N_12038,N_14933);
or U19456 (N_19456,N_14336,N_14308);
or U19457 (N_19457,N_13428,N_11383);
nor U19458 (N_19458,N_14067,N_14246);
and U19459 (N_19459,N_10610,N_10724);
nor U19460 (N_19460,N_13021,N_13932);
and U19461 (N_19461,N_14702,N_14086);
or U19462 (N_19462,N_11500,N_14728);
and U19463 (N_19463,N_11977,N_14490);
xor U19464 (N_19464,N_12288,N_12025);
or U19465 (N_19465,N_11342,N_12039);
and U19466 (N_19466,N_14626,N_13627);
nand U19467 (N_19467,N_12145,N_13253);
nor U19468 (N_19468,N_10876,N_14176);
xor U19469 (N_19469,N_10786,N_10555);
and U19470 (N_19470,N_14348,N_14439);
xnor U19471 (N_19471,N_10850,N_12482);
nor U19472 (N_19472,N_10028,N_14855);
or U19473 (N_19473,N_12233,N_10038);
or U19474 (N_19474,N_10181,N_10537);
and U19475 (N_19475,N_10060,N_12236);
and U19476 (N_19476,N_11436,N_13721);
xnor U19477 (N_19477,N_11664,N_14392);
nand U19478 (N_19478,N_14423,N_10791);
or U19479 (N_19479,N_11330,N_12851);
and U19480 (N_19480,N_10847,N_13584);
and U19481 (N_19481,N_10894,N_11932);
or U19482 (N_19482,N_12909,N_12288);
and U19483 (N_19483,N_11043,N_10900);
nor U19484 (N_19484,N_12165,N_10588);
nor U19485 (N_19485,N_12903,N_14469);
nor U19486 (N_19486,N_11486,N_11194);
nor U19487 (N_19487,N_13512,N_14008);
nor U19488 (N_19488,N_14146,N_14950);
nor U19489 (N_19489,N_12955,N_14439);
nor U19490 (N_19490,N_11566,N_10303);
nor U19491 (N_19491,N_10107,N_13127);
or U19492 (N_19492,N_10535,N_13441);
nor U19493 (N_19493,N_13718,N_14801);
nand U19494 (N_19494,N_11205,N_10009);
nor U19495 (N_19495,N_13459,N_13685);
nor U19496 (N_19496,N_10679,N_12698);
nand U19497 (N_19497,N_13109,N_14701);
nand U19498 (N_19498,N_13907,N_14003);
and U19499 (N_19499,N_14346,N_10632);
nand U19500 (N_19500,N_13196,N_11550);
and U19501 (N_19501,N_13867,N_12798);
xnor U19502 (N_19502,N_14017,N_13539);
and U19503 (N_19503,N_13460,N_10464);
nand U19504 (N_19504,N_11792,N_13167);
and U19505 (N_19505,N_11683,N_10250);
nor U19506 (N_19506,N_10806,N_13715);
nor U19507 (N_19507,N_13720,N_11868);
nand U19508 (N_19508,N_11713,N_10371);
nor U19509 (N_19509,N_13514,N_14600);
nor U19510 (N_19510,N_10054,N_13032);
nand U19511 (N_19511,N_10806,N_12391);
nor U19512 (N_19512,N_10806,N_13463);
nor U19513 (N_19513,N_10811,N_12048);
xor U19514 (N_19514,N_14279,N_10021);
nor U19515 (N_19515,N_13117,N_11731);
or U19516 (N_19516,N_11485,N_11986);
or U19517 (N_19517,N_12641,N_14852);
or U19518 (N_19518,N_12025,N_10845);
nor U19519 (N_19519,N_10702,N_11129);
or U19520 (N_19520,N_13869,N_11146);
nor U19521 (N_19521,N_10841,N_13488);
or U19522 (N_19522,N_10691,N_13582);
nand U19523 (N_19523,N_10013,N_14141);
nand U19524 (N_19524,N_14892,N_10931);
or U19525 (N_19525,N_14642,N_14885);
nor U19526 (N_19526,N_10825,N_14260);
nor U19527 (N_19527,N_13761,N_13870);
nor U19528 (N_19528,N_11019,N_10493);
and U19529 (N_19529,N_11875,N_12715);
nand U19530 (N_19530,N_11625,N_10380);
or U19531 (N_19531,N_12970,N_14613);
or U19532 (N_19532,N_13543,N_12873);
nand U19533 (N_19533,N_12824,N_12606);
and U19534 (N_19534,N_10267,N_13903);
and U19535 (N_19535,N_13107,N_11117);
xnor U19536 (N_19536,N_12547,N_10838);
or U19537 (N_19537,N_13175,N_10797);
nor U19538 (N_19538,N_13980,N_10404);
and U19539 (N_19539,N_12796,N_12569);
nor U19540 (N_19540,N_12739,N_12882);
and U19541 (N_19541,N_14288,N_14516);
and U19542 (N_19542,N_13253,N_12364);
or U19543 (N_19543,N_10912,N_10661);
and U19544 (N_19544,N_11410,N_12168);
nor U19545 (N_19545,N_11978,N_14575);
nand U19546 (N_19546,N_10405,N_14658);
and U19547 (N_19547,N_10695,N_10754);
nor U19548 (N_19548,N_14932,N_10394);
nor U19549 (N_19549,N_11618,N_12714);
nand U19550 (N_19550,N_10297,N_11753);
and U19551 (N_19551,N_10029,N_13176);
nor U19552 (N_19552,N_14463,N_11270);
nor U19553 (N_19553,N_13938,N_12880);
or U19554 (N_19554,N_13336,N_12168);
nand U19555 (N_19555,N_10685,N_10625);
nor U19556 (N_19556,N_11165,N_12239);
and U19557 (N_19557,N_13030,N_12726);
xor U19558 (N_19558,N_11975,N_14833);
or U19559 (N_19559,N_12468,N_11411);
or U19560 (N_19560,N_13288,N_10690);
nand U19561 (N_19561,N_12045,N_14680);
or U19562 (N_19562,N_14292,N_14445);
or U19563 (N_19563,N_13029,N_13670);
or U19564 (N_19564,N_12752,N_12623);
nor U19565 (N_19565,N_10201,N_13323);
nor U19566 (N_19566,N_13673,N_13308);
and U19567 (N_19567,N_13451,N_10884);
nor U19568 (N_19568,N_13933,N_11545);
nor U19569 (N_19569,N_11983,N_13193);
nor U19570 (N_19570,N_12005,N_11434);
nor U19571 (N_19571,N_12602,N_13393);
nand U19572 (N_19572,N_11287,N_14006);
and U19573 (N_19573,N_10146,N_10212);
nand U19574 (N_19574,N_10741,N_10358);
and U19575 (N_19575,N_14014,N_13429);
nand U19576 (N_19576,N_11109,N_13072);
nand U19577 (N_19577,N_10111,N_10966);
nor U19578 (N_19578,N_11577,N_12557);
nand U19579 (N_19579,N_11079,N_11928);
or U19580 (N_19580,N_10037,N_10314);
nand U19581 (N_19581,N_10053,N_11061);
and U19582 (N_19582,N_12628,N_12368);
nor U19583 (N_19583,N_11300,N_13779);
and U19584 (N_19584,N_12330,N_10854);
and U19585 (N_19585,N_12259,N_10098);
or U19586 (N_19586,N_10991,N_10251);
nor U19587 (N_19587,N_11446,N_13978);
nand U19588 (N_19588,N_10124,N_10802);
nand U19589 (N_19589,N_12586,N_14148);
and U19590 (N_19590,N_10635,N_11462);
nor U19591 (N_19591,N_12073,N_14959);
xnor U19592 (N_19592,N_13964,N_11552);
or U19593 (N_19593,N_13954,N_14124);
nor U19594 (N_19594,N_14056,N_11291);
xnor U19595 (N_19595,N_10333,N_11695);
or U19596 (N_19596,N_14967,N_12444);
nor U19597 (N_19597,N_11965,N_12036);
and U19598 (N_19598,N_10577,N_13941);
and U19599 (N_19599,N_12120,N_11996);
and U19600 (N_19600,N_10194,N_12154);
nor U19601 (N_19601,N_14758,N_13074);
or U19602 (N_19602,N_13627,N_10338);
or U19603 (N_19603,N_10565,N_14392);
xor U19604 (N_19604,N_10431,N_13318);
nor U19605 (N_19605,N_11148,N_12190);
and U19606 (N_19606,N_10003,N_11847);
or U19607 (N_19607,N_10387,N_13354);
and U19608 (N_19608,N_12632,N_10329);
xnor U19609 (N_19609,N_13642,N_12148);
or U19610 (N_19610,N_12463,N_13068);
or U19611 (N_19611,N_14268,N_14840);
xor U19612 (N_19612,N_14649,N_13667);
and U19613 (N_19613,N_14234,N_10014);
nor U19614 (N_19614,N_13392,N_10232);
xor U19615 (N_19615,N_13296,N_12800);
xnor U19616 (N_19616,N_11085,N_10294);
and U19617 (N_19617,N_14896,N_14480);
nand U19618 (N_19618,N_14503,N_12790);
nor U19619 (N_19619,N_13928,N_12157);
nor U19620 (N_19620,N_14547,N_13894);
nand U19621 (N_19621,N_14369,N_12720);
nor U19622 (N_19622,N_10198,N_11267);
nand U19623 (N_19623,N_14413,N_11082);
nor U19624 (N_19624,N_10911,N_10721);
nand U19625 (N_19625,N_10761,N_14431);
nor U19626 (N_19626,N_10171,N_14392);
or U19627 (N_19627,N_11605,N_11959);
nand U19628 (N_19628,N_11294,N_13844);
xnor U19629 (N_19629,N_10503,N_12651);
xor U19630 (N_19630,N_12017,N_14679);
and U19631 (N_19631,N_12969,N_12757);
xnor U19632 (N_19632,N_11333,N_10353);
nand U19633 (N_19633,N_14016,N_13853);
xnor U19634 (N_19634,N_12850,N_10802);
nor U19635 (N_19635,N_14038,N_14566);
or U19636 (N_19636,N_14539,N_14024);
nor U19637 (N_19637,N_11097,N_13177);
or U19638 (N_19638,N_10511,N_13941);
and U19639 (N_19639,N_13337,N_14483);
nand U19640 (N_19640,N_10915,N_11348);
nor U19641 (N_19641,N_13066,N_10562);
nand U19642 (N_19642,N_13064,N_14238);
nor U19643 (N_19643,N_10830,N_12736);
nor U19644 (N_19644,N_11854,N_14496);
or U19645 (N_19645,N_14790,N_12158);
and U19646 (N_19646,N_10827,N_11879);
nor U19647 (N_19647,N_10119,N_10228);
xnor U19648 (N_19648,N_14170,N_12752);
nor U19649 (N_19649,N_12215,N_13621);
or U19650 (N_19650,N_11288,N_14374);
xor U19651 (N_19651,N_12573,N_14880);
or U19652 (N_19652,N_14251,N_14712);
nand U19653 (N_19653,N_11679,N_14935);
nor U19654 (N_19654,N_13348,N_10458);
or U19655 (N_19655,N_14301,N_11018);
or U19656 (N_19656,N_14043,N_10411);
nand U19657 (N_19657,N_11483,N_10238);
nand U19658 (N_19658,N_12409,N_10389);
nor U19659 (N_19659,N_11462,N_10870);
nor U19660 (N_19660,N_14547,N_12089);
nor U19661 (N_19661,N_14079,N_13897);
nor U19662 (N_19662,N_13177,N_13053);
nand U19663 (N_19663,N_13074,N_14394);
nor U19664 (N_19664,N_13837,N_10272);
nand U19665 (N_19665,N_11348,N_10924);
and U19666 (N_19666,N_13324,N_12153);
and U19667 (N_19667,N_11813,N_11978);
nand U19668 (N_19668,N_13922,N_14542);
nor U19669 (N_19669,N_13451,N_11045);
or U19670 (N_19670,N_13287,N_10810);
and U19671 (N_19671,N_11814,N_10131);
nor U19672 (N_19672,N_12115,N_11904);
nor U19673 (N_19673,N_10048,N_11673);
and U19674 (N_19674,N_11691,N_12261);
nand U19675 (N_19675,N_10282,N_13398);
or U19676 (N_19676,N_13403,N_14965);
or U19677 (N_19677,N_12641,N_11419);
or U19678 (N_19678,N_10689,N_12864);
and U19679 (N_19679,N_11467,N_14900);
nand U19680 (N_19680,N_12456,N_14989);
and U19681 (N_19681,N_13492,N_13363);
or U19682 (N_19682,N_13208,N_12515);
nand U19683 (N_19683,N_14375,N_12569);
xnor U19684 (N_19684,N_13814,N_12880);
or U19685 (N_19685,N_12017,N_10754);
and U19686 (N_19686,N_10300,N_12916);
xor U19687 (N_19687,N_10134,N_14186);
or U19688 (N_19688,N_14338,N_14274);
and U19689 (N_19689,N_12338,N_14703);
nand U19690 (N_19690,N_14397,N_11403);
and U19691 (N_19691,N_12870,N_11211);
nand U19692 (N_19692,N_10639,N_14259);
and U19693 (N_19693,N_11856,N_14749);
or U19694 (N_19694,N_12953,N_14510);
nand U19695 (N_19695,N_10115,N_11230);
nand U19696 (N_19696,N_12842,N_11113);
nor U19697 (N_19697,N_10629,N_13544);
nand U19698 (N_19698,N_11152,N_11167);
or U19699 (N_19699,N_14275,N_11998);
and U19700 (N_19700,N_11833,N_10504);
or U19701 (N_19701,N_12677,N_13720);
or U19702 (N_19702,N_14085,N_12431);
or U19703 (N_19703,N_11562,N_11188);
xnor U19704 (N_19704,N_12704,N_10741);
nor U19705 (N_19705,N_12731,N_12104);
and U19706 (N_19706,N_14083,N_14529);
and U19707 (N_19707,N_11835,N_14971);
nor U19708 (N_19708,N_11146,N_12715);
or U19709 (N_19709,N_14311,N_12838);
and U19710 (N_19710,N_14698,N_13530);
or U19711 (N_19711,N_12052,N_12502);
and U19712 (N_19712,N_10891,N_14073);
xnor U19713 (N_19713,N_11654,N_12444);
or U19714 (N_19714,N_10352,N_13691);
nand U19715 (N_19715,N_11818,N_14991);
nor U19716 (N_19716,N_12381,N_13823);
nor U19717 (N_19717,N_12254,N_14106);
or U19718 (N_19718,N_13482,N_13894);
nor U19719 (N_19719,N_14689,N_12959);
or U19720 (N_19720,N_14696,N_14959);
nand U19721 (N_19721,N_12137,N_11019);
nor U19722 (N_19722,N_13075,N_10620);
nand U19723 (N_19723,N_10036,N_14131);
nor U19724 (N_19724,N_12969,N_10477);
nor U19725 (N_19725,N_12823,N_13672);
or U19726 (N_19726,N_13803,N_13836);
and U19727 (N_19727,N_11471,N_11290);
or U19728 (N_19728,N_13783,N_11625);
or U19729 (N_19729,N_10228,N_10569);
or U19730 (N_19730,N_13294,N_10863);
or U19731 (N_19731,N_12639,N_13930);
and U19732 (N_19732,N_14365,N_13914);
nor U19733 (N_19733,N_13433,N_14490);
or U19734 (N_19734,N_12378,N_14692);
nand U19735 (N_19735,N_10314,N_11257);
or U19736 (N_19736,N_14548,N_14124);
nor U19737 (N_19737,N_14110,N_10161);
or U19738 (N_19738,N_10425,N_12105);
or U19739 (N_19739,N_13796,N_10616);
and U19740 (N_19740,N_12603,N_11963);
xor U19741 (N_19741,N_12340,N_14255);
nor U19742 (N_19742,N_13318,N_11641);
nand U19743 (N_19743,N_11401,N_10068);
and U19744 (N_19744,N_14801,N_14661);
xor U19745 (N_19745,N_13292,N_12109);
or U19746 (N_19746,N_11367,N_14890);
or U19747 (N_19747,N_12707,N_13038);
and U19748 (N_19748,N_14689,N_14425);
nand U19749 (N_19749,N_12924,N_14953);
or U19750 (N_19750,N_11741,N_10445);
nand U19751 (N_19751,N_14644,N_12144);
nor U19752 (N_19752,N_12018,N_13352);
nand U19753 (N_19753,N_10022,N_14262);
xor U19754 (N_19754,N_13601,N_14062);
or U19755 (N_19755,N_11964,N_13255);
nand U19756 (N_19756,N_11690,N_14886);
or U19757 (N_19757,N_12871,N_11489);
or U19758 (N_19758,N_11122,N_11710);
or U19759 (N_19759,N_14716,N_11263);
nor U19760 (N_19760,N_12417,N_10690);
nor U19761 (N_19761,N_14116,N_14342);
nor U19762 (N_19762,N_14308,N_13310);
or U19763 (N_19763,N_10261,N_10659);
nand U19764 (N_19764,N_13516,N_13387);
nor U19765 (N_19765,N_11108,N_13626);
and U19766 (N_19766,N_10405,N_14513);
nor U19767 (N_19767,N_12960,N_11064);
or U19768 (N_19768,N_14516,N_12696);
nor U19769 (N_19769,N_10088,N_14578);
nor U19770 (N_19770,N_13360,N_11696);
xor U19771 (N_19771,N_10842,N_11959);
nand U19772 (N_19772,N_11925,N_11873);
or U19773 (N_19773,N_10754,N_12645);
or U19774 (N_19774,N_14934,N_10261);
nor U19775 (N_19775,N_14458,N_13157);
and U19776 (N_19776,N_12226,N_11187);
or U19777 (N_19777,N_11242,N_12821);
nand U19778 (N_19778,N_12835,N_11788);
nand U19779 (N_19779,N_14171,N_14963);
nand U19780 (N_19780,N_12981,N_13694);
nand U19781 (N_19781,N_12121,N_13840);
nand U19782 (N_19782,N_14123,N_10991);
nor U19783 (N_19783,N_13093,N_11973);
nand U19784 (N_19784,N_11535,N_13703);
nor U19785 (N_19785,N_14183,N_14878);
or U19786 (N_19786,N_10593,N_14609);
nand U19787 (N_19787,N_13437,N_12424);
or U19788 (N_19788,N_11480,N_12783);
xor U19789 (N_19789,N_11154,N_12505);
or U19790 (N_19790,N_12063,N_14881);
nor U19791 (N_19791,N_13856,N_11806);
nor U19792 (N_19792,N_11251,N_13981);
nor U19793 (N_19793,N_10743,N_10232);
xnor U19794 (N_19794,N_13115,N_12921);
nor U19795 (N_19795,N_14648,N_14186);
nand U19796 (N_19796,N_13797,N_12339);
nor U19797 (N_19797,N_13635,N_14439);
nor U19798 (N_19798,N_11188,N_14840);
nor U19799 (N_19799,N_14434,N_11368);
xnor U19800 (N_19800,N_13749,N_14445);
nor U19801 (N_19801,N_10568,N_12167);
or U19802 (N_19802,N_13352,N_11196);
nand U19803 (N_19803,N_10793,N_14807);
and U19804 (N_19804,N_11050,N_12583);
xor U19805 (N_19805,N_13344,N_14864);
or U19806 (N_19806,N_12307,N_12465);
or U19807 (N_19807,N_14624,N_13996);
and U19808 (N_19808,N_12597,N_14034);
or U19809 (N_19809,N_12594,N_14281);
nand U19810 (N_19810,N_11559,N_10255);
or U19811 (N_19811,N_11018,N_14601);
or U19812 (N_19812,N_11162,N_11661);
nand U19813 (N_19813,N_13975,N_12551);
and U19814 (N_19814,N_11634,N_13839);
nor U19815 (N_19815,N_11689,N_14382);
and U19816 (N_19816,N_11704,N_14690);
nand U19817 (N_19817,N_14542,N_13790);
or U19818 (N_19818,N_11348,N_10826);
and U19819 (N_19819,N_10593,N_14026);
or U19820 (N_19820,N_12640,N_11627);
xor U19821 (N_19821,N_14838,N_10785);
nand U19822 (N_19822,N_11876,N_13185);
nand U19823 (N_19823,N_11496,N_10477);
nor U19824 (N_19824,N_14592,N_13906);
or U19825 (N_19825,N_12426,N_13721);
or U19826 (N_19826,N_14596,N_13903);
nor U19827 (N_19827,N_11059,N_12746);
or U19828 (N_19828,N_13872,N_12670);
or U19829 (N_19829,N_10133,N_10268);
xor U19830 (N_19830,N_12449,N_13597);
or U19831 (N_19831,N_10242,N_11263);
nand U19832 (N_19832,N_13716,N_12812);
and U19833 (N_19833,N_12570,N_13632);
nand U19834 (N_19834,N_12685,N_10637);
or U19835 (N_19835,N_14484,N_12315);
or U19836 (N_19836,N_13821,N_10297);
nand U19837 (N_19837,N_11380,N_12479);
nand U19838 (N_19838,N_11993,N_13307);
or U19839 (N_19839,N_11923,N_14369);
nand U19840 (N_19840,N_14961,N_13861);
nand U19841 (N_19841,N_14438,N_11643);
nand U19842 (N_19842,N_13955,N_11304);
xor U19843 (N_19843,N_12258,N_14407);
or U19844 (N_19844,N_10793,N_10192);
and U19845 (N_19845,N_10330,N_11681);
nand U19846 (N_19846,N_11383,N_12611);
nor U19847 (N_19847,N_11698,N_13936);
or U19848 (N_19848,N_12960,N_13093);
or U19849 (N_19849,N_11817,N_11317);
or U19850 (N_19850,N_12219,N_13495);
nor U19851 (N_19851,N_13020,N_11635);
nand U19852 (N_19852,N_14508,N_11325);
nand U19853 (N_19853,N_12734,N_13857);
or U19854 (N_19854,N_11174,N_10532);
and U19855 (N_19855,N_10620,N_12323);
nand U19856 (N_19856,N_12509,N_13791);
nand U19857 (N_19857,N_14226,N_10828);
nand U19858 (N_19858,N_12430,N_12197);
nand U19859 (N_19859,N_12775,N_13304);
nor U19860 (N_19860,N_11383,N_11745);
and U19861 (N_19861,N_12998,N_12060);
and U19862 (N_19862,N_11758,N_10026);
xnor U19863 (N_19863,N_12909,N_11408);
xor U19864 (N_19864,N_12672,N_13584);
nand U19865 (N_19865,N_10256,N_14637);
xnor U19866 (N_19866,N_10105,N_13743);
and U19867 (N_19867,N_14486,N_14359);
nand U19868 (N_19868,N_12666,N_13995);
or U19869 (N_19869,N_14014,N_12590);
nor U19870 (N_19870,N_11715,N_12449);
nand U19871 (N_19871,N_13000,N_13270);
nor U19872 (N_19872,N_10740,N_13486);
or U19873 (N_19873,N_13784,N_13478);
or U19874 (N_19874,N_11198,N_10087);
xor U19875 (N_19875,N_12774,N_14242);
nor U19876 (N_19876,N_12083,N_11224);
and U19877 (N_19877,N_13499,N_14762);
nor U19878 (N_19878,N_12513,N_13006);
xnor U19879 (N_19879,N_12677,N_12391);
nor U19880 (N_19880,N_12269,N_14650);
or U19881 (N_19881,N_14488,N_13126);
or U19882 (N_19882,N_11807,N_13848);
nand U19883 (N_19883,N_11006,N_12908);
nand U19884 (N_19884,N_13848,N_12354);
nor U19885 (N_19885,N_11411,N_10083);
nand U19886 (N_19886,N_13798,N_11302);
and U19887 (N_19887,N_11611,N_13565);
nand U19888 (N_19888,N_10088,N_13397);
xnor U19889 (N_19889,N_11078,N_12981);
nor U19890 (N_19890,N_10576,N_13793);
or U19891 (N_19891,N_13731,N_14052);
nand U19892 (N_19892,N_10252,N_11162);
nor U19893 (N_19893,N_10403,N_14358);
nor U19894 (N_19894,N_10320,N_10231);
nor U19895 (N_19895,N_14466,N_14813);
xor U19896 (N_19896,N_10188,N_11745);
nand U19897 (N_19897,N_10540,N_10387);
or U19898 (N_19898,N_12205,N_10377);
nand U19899 (N_19899,N_11101,N_14601);
and U19900 (N_19900,N_10757,N_11973);
nand U19901 (N_19901,N_12523,N_13012);
and U19902 (N_19902,N_13381,N_13645);
or U19903 (N_19903,N_12009,N_12116);
nor U19904 (N_19904,N_12220,N_13443);
nor U19905 (N_19905,N_12691,N_11078);
nor U19906 (N_19906,N_10204,N_13351);
nand U19907 (N_19907,N_11945,N_14374);
nor U19908 (N_19908,N_13910,N_14269);
nand U19909 (N_19909,N_13297,N_14516);
and U19910 (N_19910,N_14594,N_14586);
and U19911 (N_19911,N_13646,N_12812);
and U19912 (N_19912,N_11225,N_14332);
or U19913 (N_19913,N_13881,N_13328);
and U19914 (N_19914,N_10068,N_12232);
nand U19915 (N_19915,N_12126,N_13560);
nor U19916 (N_19916,N_13884,N_13808);
or U19917 (N_19917,N_12524,N_10457);
or U19918 (N_19918,N_13759,N_12733);
and U19919 (N_19919,N_10293,N_13755);
and U19920 (N_19920,N_14783,N_13220);
or U19921 (N_19921,N_10462,N_12563);
or U19922 (N_19922,N_13542,N_14338);
nand U19923 (N_19923,N_14536,N_14626);
xnor U19924 (N_19924,N_12507,N_12264);
and U19925 (N_19925,N_12265,N_13939);
nor U19926 (N_19926,N_10530,N_11821);
xnor U19927 (N_19927,N_12751,N_13996);
xnor U19928 (N_19928,N_13089,N_13844);
nand U19929 (N_19929,N_10240,N_14803);
or U19930 (N_19930,N_12082,N_10039);
nor U19931 (N_19931,N_11360,N_14219);
nand U19932 (N_19932,N_12277,N_11209);
and U19933 (N_19933,N_11564,N_14906);
or U19934 (N_19934,N_11570,N_10954);
and U19935 (N_19935,N_14476,N_14249);
nand U19936 (N_19936,N_13110,N_13703);
nand U19937 (N_19937,N_12270,N_12950);
nor U19938 (N_19938,N_13292,N_14892);
and U19939 (N_19939,N_13489,N_14778);
nand U19940 (N_19940,N_12198,N_13418);
nor U19941 (N_19941,N_12268,N_10861);
nand U19942 (N_19942,N_14563,N_12905);
and U19943 (N_19943,N_13175,N_14203);
nand U19944 (N_19944,N_11234,N_14016);
nand U19945 (N_19945,N_13857,N_12167);
or U19946 (N_19946,N_13086,N_14699);
and U19947 (N_19947,N_14329,N_14199);
or U19948 (N_19948,N_11173,N_13009);
or U19949 (N_19949,N_12045,N_12155);
or U19950 (N_19950,N_13109,N_11264);
or U19951 (N_19951,N_11886,N_13700);
nand U19952 (N_19952,N_10732,N_13928);
nor U19953 (N_19953,N_11670,N_10375);
and U19954 (N_19954,N_11460,N_12325);
nand U19955 (N_19955,N_10865,N_12843);
xnor U19956 (N_19956,N_14611,N_11666);
and U19957 (N_19957,N_12553,N_10113);
nand U19958 (N_19958,N_11336,N_10870);
or U19959 (N_19959,N_10126,N_13377);
or U19960 (N_19960,N_12373,N_12646);
xnor U19961 (N_19961,N_13220,N_12065);
nand U19962 (N_19962,N_14105,N_14033);
or U19963 (N_19963,N_11747,N_14352);
or U19964 (N_19964,N_12261,N_14284);
xor U19965 (N_19965,N_12529,N_10292);
or U19966 (N_19966,N_11254,N_12972);
and U19967 (N_19967,N_10151,N_10262);
nor U19968 (N_19968,N_11584,N_11404);
or U19969 (N_19969,N_13405,N_10592);
and U19970 (N_19970,N_11604,N_13721);
or U19971 (N_19971,N_13336,N_13502);
nand U19972 (N_19972,N_12803,N_10873);
and U19973 (N_19973,N_12185,N_14858);
nand U19974 (N_19974,N_13375,N_10306);
xnor U19975 (N_19975,N_10750,N_12122);
nor U19976 (N_19976,N_14321,N_13442);
nand U19977 (N_19977,N_10993,N_12480);
or U19978 (N_19978,N_14245,N_10448);
nor U19979 (N_19979,N_10697,N_14672);
nand U19980 (N_19980,N_11117,N_12591);
nor U19981 (N_19981,N_11758,N_10522);
nor U19982 (N_19982,N_11148,N_14425);
and U19983 (N_19983,N_13362,N_13467);
nor U19984 (N_19984,N_12809,N_14929);
or U19985 (N_19985,N_12855,N_14453);
xor U19986 (N_19986,N_14396,N_13361);
nor U19987 (N_19987,N_11696,N_12071);
or U19988 (N_19988,N_10427,N_10810);
nor U19989 (N_19989,N_14252,N_13254);
and U19990 (N_19990,N_10449,N_10968);
nor U19991 (N_19991,N_13782,N_11901);
or U19992 (N_19992,N_14339,N_11285);
xor U19993 (N_19993,N_12894,N_13179);
and U19994 (N_19994,N_11399,N_12300);
and U19995 (N_19995,N_13338,N_12303);
nand U19996 (N_19996,N_14521,N_12676);
nand U19997 (N_19997,N_13977,N_11064);
nor U19998 (N_19998,N_14663,N_12521);
nor U19999 (N_19999,N_12601,N_14788);
and U20000 (N_20000,N_15007,N_19830);
nand U20001 (N_20001,N_18791,N_16611);
and U20002 (N_20002,N_18639,N_19489);
nor U20003 (N_20003,N_17394,N_15482);
nand U20004 (N_20004,N_15361,N_18321);
nor U20005 (N_20005,N_17777,N_19661);
or U20006 (N_20006,N_15789,N_16787);
or U20007 (N_20007,N_15676,N_15593);
and U20008 (N_20008,N_17971,N_18705);
or U20009 (N_20009,N_16833,N_16510);
or U20010 (N_20010,N_18613,N_17736);
and U20011 (N_20011,N_15063,N_18974);
and U20012 (N_20012,N_17733,N_19110);
xnor U20013 (N_20013,N_16556,N_15832);
nand U20014 (N_20014,N_15264,N_16478);
and U20015 (N_20015,N_19935,N_17170);
nor U20016 (N_20016,N_15380,N_18760);
and U20017 (N_20017,N_18361,N_19914);
nand U20018 (N_20018,N_17022,N_18826);
nand U20019 (N_20019,N_17493,N_17140);
nor U20020 (N_20020,N_16421,N_15826);
nand U20021 (N_20021,N_19207,N_19820);
nand U20022 (N_20022,N_17849,N_16260);
or U20023 (N_20023,N_17972,N_18388);
nor U20024 (N_20024,N_19541,N_18762);
and U20025 (N_20025,N_18013,N_19642);
nor U20026 (N_20026,N_17905,N_19486);
and U20027 (N_20027,N_18953,N_18294);
nand U20028 (N_20028,N_15364,N_19390);
or U20029 (N_20029,N_16706,N_18818);
nor U20030 (N_20030,N_18028,N_18015);
or U20031 (N_20031,N_16668,N_15130);
nor U20032 (N_20032,N_15575,N_18592);
nand U20033 (N_20033,N_15247,N_18101);
nor U20034 (N_20034,N_19503,N_19129);
nor U20035 (N_20035,N_19009,N_18147);
or U20036 (N_20036,N_15419,N_16158);
or U20037 (N_20037,N_15615,N_18664);
nand U20038 (N_20038,N_19366,N_16786);
nor U20039 (N_20039,N_19946,N_19299);
nor U20040 (N_20040,N_16133,N_17573);
and U20041 (N_20041,N_18443,N_17551);
xor U20042 (N_20042,N_15988,N_16892);
and U20043 (N_20043,N_16065,N_16696);
nor U20044 (N_20044,N_18773,N_15469);
xor U20045 (N_20045,N_16800,N_19610);
or U20046 (N_20046,N_19768,N_19499);
and U20047 (N_20047,N_15002,N_18091);
or U20048 (N_20048,N_18344,N_17669);
or U20049 (N_20049,N_16533,N_17771);
nand U20050 (N_20050,N_16921,N_19670);
or U20051 (N_20051,N_15520,N_18097);
xor U20052 (N_20052,N_15874,N_18132);
and U20053 (N_20053,N_15853,N_19296);
or U20054 (N_20054,N_15598,N_17680);
or U20055 (N_20055,N_17640,N_15460);
nand U20056 (N_20056,N_15235,N_16350);
nand U20057 (N_20057,N_16915,N_15812);
or U20058 (N_20058,N_15310,N_19248);
or U20059 (N_20059,N_18650,N_16855);
xnor U20060 (N_20060,N_16048,N_17162);
or U20061 (N_20061,N_16626,N_19064);
or U20062 (N_20062,N_19228,N_18909);
nor U20063 (N_20063,N_17619,N_16842);
xor U20064 (N_20064,N_19374,N_16845);
or U20065 (N_20065,N_18307,N_16130);
and U20066 (N_20066,N_16295,N_18385);
nor U20067 (N_20067,N_17480,N_18700);
xor U20068 (N_20068,N_16363,N_19423);
nand U20069 (N_20069,N_18230,N_15614);
and U20070 (N_20070,N_19648,N_15725);
xnor U20071 (N_20071,N_19303,N_17179);
and U20072 (N_20072,N_15560,N_18858);
and U20073 (N_20073,N_18290,N_17692);
and U20074 (N_20074,N_19241,N_16730);
nand U20075 (N_20075,N_17045,N_19221);
and U20076 (N_20076,N_16671,N_19346);
nor U20077 (N_20077,N_16838,N_19536);
nor U20078 (N_20078,N_17996,N_16022);
nand U20079 (N_20079,N_15195,N_15878);
nor U20080 (N_20080,N_18469,N_19966);
nand U20081 (N_20081,N_16986,N_19615);
and U20082 (N_20082,N_17446,N_17537);
xor U20083 (N_20083,N_15496,N_15014);
nand U20084 (N_20084,N_15508,N_15766);
nand U20085 (N_20085,N_17699,N_18681);
and U20086 (N_20086,N_19348,N_17413);
and U20087 (N_20087,N_15761,N_18426);
or U20088 (N_20088,N_15576,N_16506);
nor U20089 (N_20089,N_18991,N_15799);
and U20090 (N_20090,N_18536,N_15523);
or U20091 (N_20091,N_19023,N_16781);
or U20092 (N_20092,N_17357,N_18158);
nor U20093 (N_20093,N_19012,N_19492);
nor U20094 (N_20094,N_17033,N_15749);
and U20095 (N_20095,N_16285,N_19787);
nor U20096 (N_20096,N_17097,N_18604);
and U20097 (N_20097,N_19904,N_18124);
and U20098 (N_20098,N_18244,N_15578);
and U20099 (N_20099,N_16791,N_17693);
xor U20100 (N_20100,N_18561,N_19159);
or U20101 (N_20101,N_17521,N_18793);
nor U20102 (N_20102,N_17448,N_19101);
nand U20103 (N_20103,N_15120,N_17508);
nand U20104 (N_20104,N_16316,N_16287);
nand U20105 (N_20105,N_18300,N_16358);
nand U20106 (N_20106,N_17268,N_19947);
nand U20107 (N_20107,N_16354,N_19744);
nor U20108 (N_20108,N_19294,N_18636);
and U20109 (N_20109,N_19087,N_16340);
xor U20110 (N_20110,N_18513,N_17922);
nand U20111 (N_20111,N_18541,N_19184);
and U20112 (N_20112,N_15744,N_19581);
nor U20113 (N_20113,N_17578,N_15968);
and U20114 (N_20114,N_19361,N_15328);
nand U20115 (N_20115,N_15088,N_16828);
nor U20116 (N_20116,N_17438,N_18658);
or U20117 (N_20117,N_17893,N_19688);
nor U20118 (N_20118,N_19630,N_15640);
and U20119 (N_20119,N_17564,N_15904);
and U20120 (N_20120,N_16456,N_16970);
xor U20121 (N_20121,N_15250,N_18391);
nand U20122 (N_20122,N_15180,N_17759);
xor U20123 (N_20123,N_18106,N_15727);
and U20124 (N_20124,N_19644,N_17904);
nand U20125 (N_20125,N_19852,N_18607);
and U20126 (N_20126,N_15147,N_19031);
or U20127 (N_20127,N_17721,N_17317);
nand U20128 (N_20128,N_18449,N_15820);
and U20129 (N_20129,N_19652,N_18528);
or U20130 (N_20130,N_18935,N_15896);
nand U20131 (N_20131,N_19984,N_19141);
or U20132 (N_20132,N_16508,N_18089);
nand U20133 (N_20133,N_15930,N_19730);
nor U20134 (N_20134,N_18911,N_15651);
xor U20135 (N_20135,N_16744,N_16121);
nand U20136 (N_20136,N_15022,N_15975);
nand U20137 (N_20137,N_15141,N_16330);
nand U20138 (N_20138,N_17200,N_18503);
nand U20139 (N_20139,N_17629,N_18895);
and U20140 (N_20140,N_19048,N_15753);
nand U20141 (N_20141,N_17304,N_15641);
or U20142 (N_20142,N_18008,N_17247);
nand U20143 (N_20143,N_17660,N_19238);
nand U20144 (N_20144,N_19515,N_17318);
nor U20145 (N_20145,N_19326,N_17093);
or U20146 (N_20146,N_18992,N_19573);
nor U20147 (N_20147,N_19324,N_16965);
nand U20148 (N_20148,N_15245,N_19643);
nand U20149 (N_20149,N_19538,N_18427);
and U20150 (N_20150,N_18660,N_17729);
or U20151 (N_20151,N_17032,N_15374);
xnor U20152 (N_20152,N_18638,N_15588);
nand U20153 (N_20153,N_15684,N_16712);
or U20154 (N_20154,N_17772,N_16607);
and U20155 (N_20155,N_19888,N_16951);
or U20156 (N_20156,N_17909,N_18823);
nor U20157 (N_20157,N_17159,N_15025);
or U20158 (N_20158,N_15758,N_15675);
nand U20159 (N_20159,N_15471,N_15755);
and U20160 (N_20160,N_15113,N_18123);
nor U20161 (N_20161,N_19060,N_15731);
and U20162 (N_20162,N_17152,N_17244);
nand U20163 (N_20163,N_17419,N_17106);
nor U20164 (N_20164,N_18320,N_18215);
nand U20165 (N_20165,N_15917,N_15307);
and U20166 (N_20166,N_18218,N_17555);
nor U20167 (N_20167,N_15526,N_18269);
nor U20168 (N_20168,N_19265,N_17344);
or U20169 (N_20169,N_17500,N_15194);
nand U20170 (N_20170,N_19484,N_17677);
nor U20171 (N_20171,N_19963,N_15670);
nand U20172 (N_20172,N_17435,N_18574);
nand U20173 (N_20173,N_16788,N_17254);
nand U20174 (N_20174,N_19759,N_15177);
nor U20175 (N_20175,N_16688,N_19934);
nor U20176 (N_20176,N_16038,N_19349);
or U20177 (N_20177,N_17087,N_15230);
or U20178 (N_20178,N_15237,N_15047);
nor U20179 (N_20179,N_16444,N_18640);
xor U20180 (N_20180,N_18759,N_15840);
or U20181 (N_20181,N_15199,N_16351);
xnor U20182 (N_20182,N_16715,N_16372);
nand U20183 (N_20183,N_19118,N_18862);
nand U20184 (N_20184,N_19494,N_17816);
or U20185 (N_20185,N_16032,N_15379);
nor U20186 (N_20186,N_17667,N_16063);
or U20187 (N_20187,N_18212,N_18077);
nor U20188 (N_20188,N_19080,N_18708);
xnor U20189 (N_20189,N_18422,N_17658);
nor U20190 (N_20190,N_15898,N_17248);
or U20191 (N_20191,N_19135,N_16064);
and U20192 (N_20192,N_18901,N_17334);
nand U20193 (N_20193,N_17325,N_18349);
nor U20194 (N_20194,N_18783,N_18144);
xor U20195 (N_20195,N_19473,N_18398);
or U20196 (N_20196,N_15269,N_17307);
xor U20197 (N_20197,N_16090,N_17236);
nor U20198 (N_20198,N_18839,N_17186);
and U20199 (N_20199,N_15101,N_15131);
and U20200 (N_20200,N_19126,N_19796);
or U20201 (N_20201,N_18113,N_17719);
xor U20202 (N_20202,N_19949,N_16020);
xnor U20203 (N_20203,N_19441,N_18359);
nor U20204 (N_20204,N_17786,N_17017);
nand U20205 (N_20205,N_16959,N_16750);
nor U20206 (N_20206,N_18110,N_19165);
nor U20207 (N_20207,N_18971,N_17018);
nor U20208 (N_20208,N_17841,N_16628);
nor U20209 (N_20209,N_17977,N_17063);
or U20210 (N_20210,N_18332,N_17321);
xnor U20211 (N_20211,N_17644,N_16957);
and U20212 (N_20212,N_15591,N_18169);
nor U20213 (N_20213,N_19464,N_17682);
and U20214 (N_20214,N_15791,N_17588);
or U20215 (N_20215,N_18985,N_16036);
or U20216 (N_20216,N_17223,N_19175);
or U20217 (N_20217,N_17034,N_18393);
nand U20218 (N_20218,N_15991,N_18173);
nor U20219 (N_20219,N_17826,N_15308);
nand U20220 (N_20220,N_18573,N_18632);
and U20221 (N_20221,N_18381,N_16622);
nand U20222 (N_20222,N_18583,N_18448);
nor U20223 (N_20223,N_17259,N_16543);
nor U20224 (N_20224,N_19014,N_16033);
nor U20225 (N_20225,N_15492,N_17218);
or U20226 (N_20226,N_18570,N_16699);
nor U20227 (N_20227,N_17994,N_17531);
nand U20228 (N_20228,N_15870,N_19943);
and U20229 (N_20229,N_16602,N_18776);
and U20230 (N_20230,N_18735,N_19213);
nor U20231 (N_20231,N_17476,N_15106);
nor U20232 (N_20232,N_17062,N_17890);
nor U20233 (N_20233,N_15255,N_16106);
xor U20234 (N_20234,N_16034,N_17620);
or U20235 (N_20235,N_18219,N_16975);
and U20236 (N_20236,N_19861,N_17665);
xor U20237 (N_20237,N_17896,N_17782);
and U20238 (N_20238,N_16873,N_16546);
nand U20239 (N_20239,N_19163,N_19485);
xnor U20240 (N_20240,N_19150,N_16558);
or U20241 (N_20241,N_15259,N_18825);
nand U20242 (N_20242,N_15054,N_15375);
nand U20243 (N_20243,N_16452,N_15892);
nor U20244 (N_20244,N_18420,N_17566);
and U20245 (N_20245,N_19084,N_16882);
or U20246 (N_20246,N_19574,N_19872);
nor U20247 (N_20247,N_19779,N_16512);
nor U20248 (N_20248,N_18037,N_19438);
nor U20249 (N_20249,N_17921,N_18993);
nor U20250 (N_20250,N_15564,N_15330);
nor U20251 (N_20251,N_16872,N_17160);
nor U20252 (N_20252,N_19322,N_19682);
and U20253 (N_20253,N_15290,N_18808);
or U20254 (N_20254,N_19392,N_16680);
and U20255 (N_20255,N_19773,N_19179);
nand U20256 (N_20256,N_16190,N_18897);
or U20257 (N_20257,N_19886,N_16994);
nand U20258 (N_20258,N_16905,N_18552);
and U20259 (N_20259,N_18553,N_16521);
nand U20260 (N_20260,N_15772,N_18472);
and U20261 (N_20261,N_17926,N_19646);
nand U20262 (N_20262,N_15700,N_15871);
xor U20263 (N_20263,N_17138,N_17392);
and U20264 (N_20264,N_15931,N_16958);
nor U20265 (N_20265,N_18680,N_18384);
or U20266 (N_20266,N_19425,N_15646);
and U20267 (N_20267,N_16312,N_17083);
and U20268 (N_20268,N_19289,N_15100);
and U20269 (N_20269,N_16700,N_17120);
nand U20270 (N_20270,N_15809,N_15274);
nand U20271 (N_20271,N_17421,N_18688);
or U20272 (N_20272,N_19433,N_15706);
nand U20273 (N_20273,N_16961,N_19173);
nor U20274 (N_20274,N_18237,N_19359);
xor U20275 (N_20275,N_17384,N_17336);
xor U20276 (N_20276,N_18079,N_18864);
or U20277 (N_20277,N_18525,N_16269);
nand U20278 (N_20278,N_16585,N_15343);
nand U20279 (N_20279,N_17403,N_15995);
or U20280 (N_20280,N_19414,N_16608);
and U20281 (N_20281,N_16613,N_18698);
nor U20282 (N_20282,N_15152,N_15253);
nor U20283 (N_20283,N_15779,N_19837);
and U20284 (N_20284,N_15146,N_17597);
xor U20285 (N_20285,N_18020,N_19846);
or U20286 (N_20286,N_18947,N_15422);
nor U20287 (N_20287,N_18622,N_16540);
and U20288 (N_20288,N_16014,N_16139);
nand U20289 (N_20289,N_16485,N_16297);
or U20290 (N_20290,N_17420,N_18342);
nor U20291 (N_20291,N_17608,N_19867);
and U20292 (N_20292,N_18382,N_19552);
nand U20293 (N_20293,N_18339,N_18334);
or U20294 (N_20294,N_16684,N_17800);
or U20295 (N_20295,N_15524,N_16465);
nor U20296 (N_20296,N_18521,N_16343);
nor U20297 (N_20297,N_15171,N_19936);
nor U20298 (N_20298,N_17346,N_15179);
xnor U20299 (N_20299,N_19666,N_15481);
or U20300 (N_20300,N_16814,N_16291);
and U20301 (N_20301,N_19436,N_17598);
and U20302 (N_20302,N_16311,N_19409);
nor U20303 (N_20303,N_15949,N_19605);
nand U20304 (N_20304,N_15618,N_15915);
nor U20305 (N_20305,N_18516,N_17602);
nand U20306 (N_20306,N_17023,N_16764);
or U20307 (N_20307,N_18143,N_18691);
nor U20308 (N_20308,N_15395,N_19649);
or U20309 (N_20309,N_16275,N_19338);
nor U20310 (N_20310,N_18686,N_18239);
nand U20311 (N_20311,N_16797,N_17422);
or U20312 (N_20312,N_18830,N_19956);
nor U20313 (N_20313,N_15568,N_16601);
and U20314 (N_20314,N_16366,N_15140);
xor U20315 (N_20315,N_15544,N_17916);
and U20316 (N_20316,N_15409,N_18441);
or U20317 (N_20317,N_19223,N_18271);
or U20318 (N_20318,N_17709,N_19116);
or U20319 (N_20319,N_18096,N_15213);
and U20320 (N_20320,N_18714,N_15294);
or U20321 (N_20321,N_19273,N_16498);
nand U20322 (N_20322,N_17155,N_17024);
and U20323 (N_20323,N_18980,N_17520);
and U20324 (N_20324,N_17559,N_18672);
nand U20325 (N_20325,N_19683,N_16220);
nand U20326 (N_20326,N_15719,N_18586);
nor U20327 (N_20327,N_17123,N_15090);
nor U20328 (N_20328,N_17132,N_15542);
nand U20329 (N_20329,N_15236,N_18498);
nand U20330 (N_20330,N_15355,N_16303);
xnor U20331 (N_20331,N_15792,N_15887);
and U20332 (N_20332,N_17609,N_15004);
xnor U20333 (N_20333,N_18526,N_18763);
nand U20334 (N_20334,N_17324,N_18724);
or U20335 (N_20335,N_17220,N_17740);
or U20336 (N_20336,N_18276,N_18531);
nand U20337 (N_20337,N_16457,N_15233);
nand U20338 (N_20338,N_18298,N_16829);
nand U20339 (N_20339,N_18363,N_15024);
and U20340 (N_20340,N_16049,N_19339);
nor U20341 (N_20341,N_17262,N_18118);
and U20342 (N_20342,N_19544,N_16035);
nor U20343 (N_20343,N_19099,N_16298);
and U20344 (N_20344,N_18390,N_17381);
nand U20345 (N_20345,N_19193,N_18407);
nor U20346 (N_20346,N_19725,N_15376);
nor U20347 (N_20347,N_19131,N_16194);
and U20348 (N_20348,N_19229,N_18273);
nor U20349 (N_20349,N_18183,N_17488);
nand U20350 (N_20350,N_16826,N_16093);
xor U20351 (N_20351,N_15351,N_15225);
and U20352 (N_20352,N_15559,N_18984);
nor U20353 (N_20353,N_15008,N_15982);
or U20354 (N_20354,N_16805,N_18341);
and U20355 (N_20355,N_16414,N_19836);
and U20356 (N_20356,N_15293,N_17860);
nand U20357 (N_20357,N_16239,N_19996);
nor U20358 (N_20358,N_15852,N_16904);
or U20359 (N_20359,N_19382,N_18975);
or U20360 (N_20360,N_17178,N_17028);
and U20361 (N_20361,N_17802,N_18233);
nor U20362 (N_20362,N_17172,N_15932);
and U20363 (N_20363,N_18497,N_16932);
and U20364 (N_20364,N_17058,N_17272);
or U20365 (N_20365,N_18822,N_19240);
xor U20366 (N_20366,N_16563,N_19188);
and U20367 (N_20367,N_15393,N_18706);
and U20368 (N_20368,N_15413,N_18353);
or U20369 (N_20369,N_15252,N_19106);
nand U20370 (N_20370,N_16132,N_19909);
or U20371 (N_20371,N_15954,N_17335);
nand U20372 (N_20372,N_17612,N_15306);
nand U20373 (N_20373,N_17936,N_16610);
nor U20374 (N_20374,N_16113,N_15649);
nor U20375 (N_20375,N_15331,N_19819);
and U20376 (N_20376,N_18876,N_19268);
nor U20377 (N_20377,N_17434,N_18151);
nor U20378 (N_20378,N_15743,N_19288);
or U20379 (N_20379,N_18507,N_17400);
nand U20380 (N_20380,N_18696,N_19893);
and U20381 (N_20381,N_18309,N_17151);
nor U20382 (N_20382,N_19637,N_19829);
or U20383 (N_20383,N_19266,N_19983);
nor U20384 (N_20384,N_15223,N_18865);
or U20385 (N_20385,N_19572,N_16703);
or U20386 (N_20386,N_15831,N_19810);
nor U20387 (N_20387,N_16851,N_15622);
or U20388 (N_20388,N_18241,N_17315);
nand U20389 (N_20389,N_15573,N_15861);
and U20390 (N_20390,N_15044,N_18288);
or U20391 (N_20391,N_19907,N_18164);
and U20392 (N_20392,N_15964,N_16548);
nand U20393 (N_20393,N_18090,N_17014);
or U20394 (N_20394,N_17757,N_16822);
and U20395 (N_20395,N_15965,N_16462);
xor U20396 (N_20396,N_19993,N_18149);
nand U20397 (N_20397,N_18192,N_15893);
nor U20398 (N_20398,N_18646,N_15390);
or U20399 (N_20399,N_19809,N_17576);
or U20400 (N_20400,N_16662,N_17039);
nand U20401 (N_20401,N_19148,N_15543);
or U20402 (N_20402,N_15570,N_17803);
and U20403 (N_20403,N_17923,N_15862);
or U20404 (N_20404,N_19220,N_18024);
and U20405 (N_20405,N_16169,N_18820);
nor U20406 (N_20406,N_15295,N_15934);
or U20407 (N_20407,N_16542,N_17930);
nand U20408 (N_20408,N_15768,N_19052);
nand U20409 (N_20409,N_17844,N_17397);
or U20410 (N_20410,N_19431,N_15202);
xnor U20411 (N_20411,N_18973,N_18452);
nand U20412 (N_20412,N_19334,N_19576);
nand U20413 (N_20413,N_18806,N_18589);
nand U20414 (N_20414,N_19913,N_18465);
nor U20415 (N_20415,N_15627,N_19198);
nor U20416 (N_20416,N_18730,N_18293);
nor U20417 (N_20417,N_15609,N_18414);
nor U20418 (N_20418,N_17593,N_16323);
xor U20419 (N_20419,N_17582,N_17053);
and U20420 (N_20420,N_17760,N_16434);
nand U20421 (N_20421,N_17662,N_15166);
xnor U20422 (N_20422,N_17020,N_16261);
and U20423 (N_20423,N_16742,N_16078);
or U20424 (N_20424,N_19282,N_16549);
nand U20425 (N_20425,N_19561,N_15260);
nand U20426 (N_20426,N_15270,N_17374);
nor U20427 (N_20427,N_16367,N_18761);
and U20428 (N_20428,N_15780,N_17217);
nand U20429 (N_20429,N_17457,N_18600);
nor U20430 (N_20430,N_19291,N_19524);
nor U20431 (N_20431,N_18304,N_15183);
or U20432 (N_20432,N_19741,N_16187);
nand U20433 (N_20433,N_16109,N_18889);
or U20434 (N_20434,N_17857,N_17393);
or U20435 (N_20435,N_19781,N_15845);
nor U20436 (N_20436,N_16501,N_15324);
nor U20437 (N_20437,N_15606,N_17687);
or U20438 (N_20438,N_18579,N_18948);
nand U20439 (N_20439,N_19699,N_18289);
and U20440 (N_20440,N_16483,N_15633);
or U20441 (N_20441,N_17941,N_18485);
nand U20442 (N_20442,N_16514,N_15771);
nand U20443 (N_20443,N_15312,N_19875);
nand U20444 (N_20444,N_16251,N_19007);
and U20445 (N_20445,N_15082,N_19045);
nor U20446 (N_20446,N_17797,N_16317);
nand U20447 (N_20447,N_19557,N_15629);
nor U20448 (N_20448,N_19219,N_19032);
xor U20449 (N_20449,N_18501,N_18193);
or U20450 (N_20450,N_18095,N_18804);
and U20451 (N_20451,N_17678,N_19603);
or U20452 (N_20452,N_15586,N_18796);
nor U20453 (N_20453,N_17464,N_18651);
and U20454 (N_20454,N_17169,N_18253);
nor U20455 (N_20455,N_15961,N_15696);
or U20456 (N_20456,N_18802,N_17451);
nor U20457 (N_20457,N_16524,N_18610);
and U20458 (N_20458,N_18291,N_18576);
and U20459 (N_20459,N_17925,N_16108);
nor U20460 (N_20460,N_16253,N_19216);
xor U20461 (N_20461,N_15064,N_17275);
nand U20462 (N_20462,N_19824,N_19008);
xor U20463 (N_20463,N_17267,N_16497);
nor U20464 (N_20464,N_18733,N_15071);
or U20465 (N_20465,N_17517,N_16356);
or U20466 (N_20466,N_18429,N_15770);
and U20467 (N_20467,N_16647,N_19177);
nand U20468 (N_20468,N_19332,N_15254);
nand U20469 (N_20469,N_18050,N_15455);
nor U20470 (N_20470,N_17993,N_18323);
nor U20471 (N_20471,N_16880,N_19916);
nand U20472 (N_20472,N_15026,N_19067);
nand U20473 (N_20473,N_18585,N_16355);
or U20474 (N_20474,N_16931,N_17050);
or U20475 (N_20475,N_16537,N_16545);
and U20476 (N_20476,N_18468,N_15275);
nand U20477 (N_20477,N_15685,N_17884);
and U20478 (N_20478,N_15143,N_17741);
or U20479 (N_20479,N_16609,N_19170);
nor U20480 (N_20480,N_18072,N_18296);
nand U20481 (N_20481,N_16189,N_15005);
nor U20482 (N_20482,N_15415,N_17743);
or U20483 (N_20483,N_19355,N_15738);
and U20484 (N_20484,N_16467,N_17811);
and U20485 (N_20485,N_16007,N_17758);
and U20486 (N_20486,N_18069,N_17080);
nand U20487 (N_20487,N_19261,N_18805);
nand U20488 (N_20488,N_15210,N_18251);
nand U20489 (N_20489,N_18167,N_19564);
xnor U20490 (N_20490,N_15353,N_16119);
nand U20491 (N_20491,N_19675,N_18799);
nor U20492 (N_20492,N_18972,N_15383);
nand U20493 (N_20493,N_18615,N_15052);
nand U20494 (N_20494,N_19667,N_19280);
or U20495 (N_20495,N_17214,N_18564);
nand U20496 (N_20496,N_15857,N_15894);
nand U20497 (N_20497,N_18040,N_18051);
or U20498 (N_20498,N_16687,N_19986);
and U20499 (N_20499,N_17285,N_18915);
and U20500 (N_20500,N_18861,N_19747);
and U20501 (N_20501,N_18542,N_17762);
xnor U20502 (N_20502,N_15370,N_16114);
xnor U20503 (N_20503,N_17842,N_15406);
nand U20504 (N_20504,N_19070,N_19720);
or U20505 (N_20505,N_19209,N_16762);
or U20506 (N_20506,N_18959,N_16067);
nand U20507 (N_20507,N_15730,N_16648);
nor U20508 (N_20508,N_16055,N_19145);
xnor U20509 (N_20509,N_16346,N_15597);
nand U20510 (N_20510,N_18731,N_19446);
and U20511 (N_20511,N_15282,N_19941);
nand U20512 (N_20512,N_18707,N_19608);
nor U20513 (N_20513,N_18868,N_19244);
and U20514 (N_20514,N_15139,N_16583);
nand U20515 (N_20515,N_15222,N_15813);
nor U20516 (N_20516,N_16659,N_16438);
and U20517 (N_20517,N_16041,N_17115);
xnor U20518 (N_20518,N_15883,N_15834);
nor U20519 (N_20519,N_16370,N_15807);
nor U20520 (N_20520,N_15648,N_19587);
xor U20521 (N_20521,N_16267,N_17661);
nand U20522 (N_20522,N_18004,N_15848);
nand U20523 (N_20523,N_19957,N_15592);
nand U20524 (N_20524,N_19871,N_15732);
or U20525 (N_20525,N_16653,N_19130);
and U20526 (N_20526,N_16581,N_16686);
xor U20527 (N_20527,N_19352,N_16460);
or U20528 (N_20528,N_18534,N_16751);
nand U20529 (N_20529,N_19604,N_17527);
or U20530 (N_20530,N_16695,N_17130);
xnor U20531 (N_20531,N_15504,N_17376);
or U20532 (N_20532,N_16188,N_16216);
and U20533 (N_20533,N_17156,N_15137);
xnor U20534 (N_20534,N_18517,N_15468);
or U20535 (N_20535,N_19138,N_15391);
nor U20536 (N_20536,N_16024,N_18931);
nor U20537 (N_20537,N_18612,N_15373);
nor U20538 (N_20538,N_15590,N_18652);
xor U20539 (N_20539,N_15326,N_19337);
nand U20540 (N_20540,N_18685,N_16279);
nand U20541 (N_20541,N_17042,N_19804);
nand U20542 (N_20542,N_18933,N_15548);
nor U20543 (N_20543,N_16218,N_15604);
and U20544 (N_20544,N_17369,N_15172);
nand U20545 (N_20545,N_18884,N_16985);
xor U20546 (N_20546,N_19786,N_16000);
or U20547 (N_20547,N_15271,N_17664);
nor U20548 (N_20548,N_17747,N_19236);
nor U20549 (N_20549,N_17467,N_15487);
nor U20550 (N_20550,N_19459,N_15918);
nor U20551 (N_20551,N_15824,N_19647);
and U20552 (N_20552,N_16407,N_17703);
nand U20553 (N_20553,N_19413,N_18745);
nor U20554 (N_20554,N_16205,N_18435);
and U20555 (N_20555,N_15365,N_15035);
nor U20556 (N_20556,N_15876,N_15516);
or U20557 (N_20557,N_17373,N_18140);
nor U20558 (N_20558,N_15860,N_16329);
and U20559 (N_20559,N_17180,N_16266);
and U20560 (N_20560,N_18489,N_18845);
or U20561 (N_20561,N_15742,N_17183);
nor U20562 (N_20562,N_15479,N_18105);
nand U20563 (N_20563,N_15859,N_17303);
nand U20564 (N_20564,N_19420,N_19119);
nand U20565 (N_20565,N_17366,N_17173);
nand U20566 (N_20566,N_17171,N_15754);
and U20567 (N_20567,N_16623,N_19166);
and U20568 (N_20568,N_16154,N_16231);
nand U20569 (N_20569,N_16660,N_17074);
or U20570 (N_20570,N_15133,N_19292);
and U20571 (N_20571,N_16023,N_16237);
nand U20572 (N_20572,N_15450,N_16028);
nor U20573 (N_20573,N_18080,N_19911);
xnor U20574 (N_20574,N_16940,N_19693);
or U20575 (N_20575,N_15821,N_17750);
nand U20576 (N_20576,N_17301,N_15924);
nand U20577 (N_20577,N_19923,N_17144);
nand U20578 (N_20578,N_17202,N_19921);
and U20579 (N_20579,N_18891,N_18955);
nand U20580 (N_20580,N_16541,N_17683);
nor U20581 (N_20581,N_17051,N_17888);
or U20582 (N_20582,N_15987,N_18495);
or U20583 (N_20583,N_16804,N_17892);
nand U20584 (N_20584,N_17836,N_19063);
nand U20585 (N_20585,N_18314,N_15056);
or U20586 (N_20586,N_18946,N_16678);
nor U20587 (N_20587,N_16159,N_17141);
nor U20588 (N_20588,N_16163,N_17474);
or U20589 (N_20589,N_16137,N_18721);
nand U20590 (N_20590,N_16755,N_19061);
nand U20591 (N_20591,N_18139,N_16406);
nor U20592 (N_20592,N_16990,N_17418);
or U20593 (N_20593,N_16413,N_17249);
or U20594 (N_20594,N_15811,N_17266);
xnor U20595 (N_20595,N_19117,N_19582);
or U20596 (N_20596,N_17992,N_19657);
nand U20597 (N_20597,N_16555,N_15452);
xnor U20598 (N_20598,N_19532,N_17191);
and U20599 (N_20599,N_18405,N_15369);
xor U20600 (N_20600,N_16996,N_17813);
nand U20601 (N_20601,N_15912,N_18409);
xnor U20602 (N_20602,N_16071,N_17206);
and U20603 (N_20603,N_16852,N_15950);
and U20604 (N_20604,N_19072,N_15841);
and U20605 (N_20605,N_19488,N_17444);
nand U20606 (N_20606,N_19883,N_16906);
nand U20607 (N_20607,N_17131,N_18466);
nand U20608 (N_20608,N_15473,N_19187);
nor U20609 (N_20609,N_17961,N_15790);
nor U20610 (N_20610,N_18042,N_18684);
and U20611 (N_20611,N_15491,N_17030);
nand U20612 (N_20612,N_17201,N_19152);
and U20613 (N_20613,N_15880,N_15303);
and U20614 (N_20614,N_19171,N_17825);
nor U20615 (N_20615,N_17468,N_18625);
or U20616 (N_20616,N_16375,N_19471);
and U20617 (N_20617,N_16238,N_15866);
nand U20618 (N_20618,N_18875,N_16592);
and U20619 (N_20619,N_18068,N_16480);
and U20620 (N_20620,N_17913,N_17799);
and U20621 (N_20621,N_19400,N_16449);
and U20622 (N_20622,N_16547,N_18922);
nand U20623 (N_20623,N_19487,N_17350);
and U20624 (N_20624,N_19037,N_18634);
or U20625 (N_20625,N_15666,N_17756);
and U20626 (N_20626,N_15188,N_15459);
nor U20627 (N_20627,N_16252,N_15385);
and U20628 (N_20628,N_18054,N_15302);
nor U20629 (N_20629,N_18411,N_15577);
nand U20630 (N_20630,N_15602,N_18923);
and U20631 (N_20631,N_15182,N_17250);
and U20632 (N_20632,N_18200,N_19258);
and U20633 (N_20633,N_18220,N_19718);
or U20634 (N_20634,N_17681,N_17428);
nor U20635 (N_20635,N_19569,N_18725);
xor U20636 (N_20636,N_17623,N_17095);
or U20637 (N_20637,N_18964,N_17308);
and U20638 (N_20638,N_16734,N_17895);
and U20639 (N_20639,N_19466,N_19547);
nand U20640 (N_20640,N_17118,N_17506);
or U20641 (N_20641,N_15801,N_17684);
and U20642 (N_20642,N_15956,N_18007);
and U20643 (N_20643,N_17791,N_15359);
and U20644 (N_20644,N_15914,N_15751);
nand U20645 (N_20645,N_19971,N_16993);
or U20646 (N_20646,N_17049,N_17713);
or U20647 (N_20647,N_15736,N_16318);
and U20648 (N_20648,N_18703,N_19516);
and U20649 (N_20649,N_19297,N_16361);
nand U20650 (N_20650,N_18047,N_18076);
nor U20651 (N_20651,N_16395,N_15246);
nor U20652 (N_20652,N_16887,N_18904);
and U20653 (N_20653,N_16215,N_16195);
or U20654 (N_20654,N_17071,N_19997);
nand U20655 (N_20655,N_19645,N_18111);
xnor U20656 (N_20656,N_17490,N_15048);
nand U20657 (N_20657,N_18053,N_15344);
and U20658 (N_20658,N_16857,N_19395);
nor U20659 (N_20659,N_19539,N_18775);
or U20660 (N_20660,N_17707,N_18438);
nand U20661 (N_20661,N_15802,N_19703);
nand U20662 (N_20662,N_16625,N_17773);
or U20663 (N_20663,N_15721,N_16461);
nand U20664 (N_20664,N_17554,N_18960);
and U20665 (N_20665,N_16384,N_16584);
and U20666 (N_20666,N_15619,N_15974);
or U20667 (N_20667,N_19001,N_15728);
xnor U20668 (N_20668,N_18228,N_17242);
xor U20669 (N_20669,N_15740,N_19437);
and U20670 (N_20670,N_15248,N_17470);
or U20671 (N_20671,N_16870,N_19312);
nor U20672 (N_20672,N_17878,N_18851);
nand U20673 (N_20673,N_15976,N_15318);
or U20674 (N_20674,N_19987,N_17689);
and U20675 (N_20675,N_19784,N_18044);
nor U20676 (N_20676,N_16219,N_17145);
and U20677 (N_20677,N_18565,N_16221);
and U20678 (N_20678,N_17360,N_19847);
nand U20679 (N_20679,N_16576,N_15679);
nand U20680 (N_20680,N_16614,N_17987);
or U20681 (N_20681,N_17980,N_17929);
nand U20682 (N_20682,N_15617,N_16489);
nand U20683 (N_20683,N_16247,N_15432);
xor U20684 (N_20684,N_17371,N_19103);
nand U20685 (N_20685,N_16573,N_19262);
and U20686 (N_20686,N_18356,N_15994);
or U20687 (N_20687,N_17867,N_15085);
and U20688 (N_20688,N_19202,N_16332);
nand U20689 (N_20689,N_18029,N_19300);
and U20690 (N_20690,N_17714,N_16564);
nor U20691 (N_20691,N_15557,N_15998);
nand U20692 (N_20692,N_18121,N_16271);
and U20693 (N_20693,N_18197,N_17542);
and U20694 (N_20694,N_16447,N_18368);
and U20695 (N_20695,N_19930,N_15833);
nand U20696 (N_20696,N_19447,N_19107);
and U20697 (N_20697,N_19233,N_17255);
nand U20698 (N_20698,N_15220,N_18277);
xnor U20699 (N_20699,N_18643,N_19991);
nor U20700 (N_20700,N_15613,N_19686);
nand U20701 (N_20701,N_19687,N_15436);
or U20702 (N_20702,N_18185,N_16333);
and U20703 (N_20703,N_18189,N_18620);
and U20704 (N_20704,N_19985,N_19157);
nor U20705 (N_20705,N_15156,N_17211);
or U20706 (N_20706,N_16536,N_19892);
and U20707 (N_20707,N_17319,N_16526);
xnor U20708 (N_20708,N_15350,N_16728);
and U20709 (N_20709,N_19472,N_19782);
or U20710 (N_20710,N_19685,N_18413);
or U20711 (N_20711,N_16973,N_17379);
and U20712 (N_20712,N_17801,N_15046);
nor U20713 (N_20713,N_17339,N_18318);
xor U20714 (N_20714,N_17341,N_18175);
nand U20715 (N_20715,N_17001,N_17208);
nor U20716 (N_20716,N_16017,N_16319);
xnor U20717 (N_20717,N_17853,N_15599);
and U20718 (N_20718,N_18509,N_18071);
or U20719 (N_20719,N_19897,N_16910);
nand U20720 (N_20720,N_18177,N_18981);
and U20721 (N_20721,N_15623,N_18821);
nor U20722 (N_20722,N_16198,N_16763);
nand U20723 (N_20723,N_19734,N_17387);
or U20724 (N_20724,N_18209,N_17440);
nand U20725 (N_20725,N_17712,N_18621);
xor U20726 (N_20726,N_19813,N_17225);
and U20727 (N_20727,N_18394,N_17808);
and U20728 (N_20728,N_17563,N_16605);
and U20729 (N_20729,N_19519,N_16021);
nand U20730 (N_20730,N_16691,N_18440);
nand U20731 (N_20731,N_16393,N_19039);
xor U20732 (N_20732,N_19509,N_19384);
and U20733 (N_20733,N_18306,N_18930);
or U20734 (N_20734,N_17763,N_19662);
nand U20735 (N_20735,N_17872,N_19508);
nand U20736 (N_20736,N_17368,N_18295);
nor U20737 (N_20737,N_18447,N_19479);
nor U20738 (N_20738,N_17625,N_16008);
and U20739 (N_20739,N_16365,N_15249);
or U20740 (N_20740,N_19056,N_19321);
nor U20741 (N_20741,N_17632,N_19614);
nand U20742 (N_20742,N_17090,N_17436);
nand U20743 (N_20743,N_15506,N_16840);
or U20744 (N_20744,N_16019,N_17497);
nor U20745 (N_20745,N_19938,N_17455);
nand U20746 (N_20746,N_19375,N_17101);
or U20747 (N_20747,N_18676,N_16116);
nor U20748 (N_20748,N_17973,N_19651);
and U20749 (N_20749,N_18601,N_18430);
nor U20750 (N_20750,N_17607,N_16848);
and U20751 (N_20751,N_19636,N_17694);
or U20752 (N_20752,N_16226,N_19870);
and U20753 (N_20753,N_15842,N_16559);
nand U20754 (N_20754,N_17656,N_15124);
or U20755 (N_20755,N_18756,N_17367);
nor U20756 (N_20756,N_16806,N_15773);
nor U20757 (N_20757,N_16637,N_19673);
nand U20758 (N_20758,N_17273,N_17008);
nor U20759 (N_20759,N_18162,N_18715);
nor U20760 (N_20760,N_17119,N_19098);
xnor U20761 (N_20761,N_15611,N_16103);
or U20762 (N_20762,N_17863,N_18979);
nand U20763 (N_20763,N_16339,N_16553);
nand U20764 (N_20764,N_19036,N_19158);
nor U20765 (N_20765,N_18653,N_19680);
or U20766 (N_20766,N_17950,N_16309);
or U20767 (N_20767,N_15013,N_18198);
and U20768 (N_20768,N_18112,N_17469);
nand U20769 (N_20769,N_18732,N_16745);
or U20770 (N_20770,N_15856,N_18360);
nand U20771 (N_20771,N_16336,N_17294);
or U20772 (N_20772,N_19674,N_19190);
or U20773 (N_20773,N_19827,N_19245);
and U20774 (N_20774,N_17984,N_15142);
xor U20775 (N_20775,N_16667,N_19588);
nand U20776 (N_20776,N_17544,N_17343);
and U20777 (N_20777,N_19323,N_15683);
and U20778 (N_20778,N_17601,N_18267);
or U20779 (N_20779,N_16843,N_15338);
and U20780 (N_20780,N_16850,N_18927);
xnor U20781 (N_20781,N_18754,N_18027);
xnor U20782 (N_20782,N_17540,N_19362);
nor U20783 (N_20783,N_17263,N_17955);
or U20784 (N_20784,N_19559,N_16338);
nor U20785 (N_20785,N_16293,N_17781);
and U20786 (N_20786,N_19372,N_18872);
nor U20787 (N_20787,N_18174,N_15039);
nand U20788 (N_20788,N_19942,N_16798);
and U20789 (N_20789,N_15538,N_15985);
nor U20790 (N_20790,N_17805,N_15693);
and U20791 (N_20791,N_17907,N_16759);
nand U20792 (N_20792,N_19593,N_16726);
nand U20793 (N_20793,N_16560,N_16732);
nor U20794 (N_20794,N_18246,N_18770);
and U20795 (N_20795,N_19195,N_15963);
nor U20796 (N_20796,N_15381,N_17840);
nor U20797 (N_20797,N_18560,N_19419);
and U20798 (N_20798,N_15774,N_16263);
nand U20799 (N_20799,N_19424,N_19426);
and U20800 (N_20800,N_16527,N_18750);
nor U20801 (N_20801,N_19351,N_17834);
and U20802 (N_20802,N_19520,N_15660);
or U20803 (N_20803,N_19405,N_16782);
nand U20804 (N_20804,N_17976,N_18729);
nand U20805 (N_20805,N_19343,N_18550);
or U20806 (N_20806,N_18631,N_16949);
or U20807 (N_20807,N_19427,N_19252);
nand U20808 (N_20808,N_17292,N_16308);
xor U20809 (N_20809,N_17584,N_17839);
and U20810 (N_20810,N_17483,N_17818);
and U20811 (N_20811,N_17117,N_16938);
xnor U20812 (N_20812,N_17738,N_18346);
nor U20813 (N_20813,N_19286,N_18742);
nand U20814 (N_20814,N_16903,N_18064);
or U20815 (N_20815,N_19728,N_19671);
xor U20816 (N_20816,N_18637,N_15116);
nor U20817 (N_20817,N_16262,N_17102);
xnor U20818 (N_20818,N_19164,N_16274);
nand U20819 (N_20819,N_17523,N_19855);
nor U20820 (N_20820,N_18103,N_15212);
and U20821 (N_20821,N_15796,N_17568);
nor U20822 (N_20822,N_19011,N_18879);
and U20823 (N_20823,N_16399,N_15989);
nor U20824 (N_20824,N_18833,N_18061);
and U20825 (N_20825,N_19612,N_16122);
xor U20826 (N_20826,N_17603,N_18626);
nor U20827 (N_20827,N_16084,N_18969);
and U20828 (N_20828,N_19199,N_16152);
nor U20829 (N_20829,N_17512,N_15572);
and U20830 (N_20830,N_19567,N_19483);
xor U20831 (N_20831,N_17060,N_15036);
and U20832 (N_20832,N_17154,N_19558);
and U20833 (N_20833,N_17641,N_17937);
nand U20834 (N_20834,N_17847,N_15499);
and U20835 (N_20835,N_18988,N_15261);
and U20836 (N_20836,N_19096,N_18421);
and U20837 (N_20837,N_17964,N_19690);
or U20838 (N_20838,N_17489,N_16196);
or U20839 (N_20839,N_18201,N_15939);
nor U20840 (N_20840,N_15978,N_15688);
nor U20841 (N_20841,N_19828,N_16520);
or U20842 (N_20842,N_16076,N_16928);
nand U20843 (N_20843,N_16208,N_16654);
or U20844 (N_20844,N_19811,N_15815);
nor U20845 (N_20845,N_15643,N_15081);
or U20846 (N_20846,N_17442,N_16801);
nor U20847 (N_20847,N_15787,N_16493);
xnor U20848 (N_20848,N_15537,N_19713);
nand U20849 (N_20849,N_18878,N_16492);
and U20850 (N_20850,N_15872,N_18486);
nand U20851 (N_20851,N_18446,N_15838);
nor U20852 (N_20852,N_18591,N_16532);
nand U20853 (N_20853,N_18787,N_15867);
and U20854 (N_20854,N_17443,N_19873);
nor U20855 (N_20855,N_15352,N_19899);
or U20856 (N_20856,N_17622,N_16379);
or U20857 (N_20857,N_16072,N_15503);
nor U20858 (N_20858,N_15958,N_18918);
nor U20859 (N_20859,N_19481,N_17663);
xor U20860 (N_20860,N_17163,N_15164);
nand U20861 (N_20861,N_17185,N_17526);
or U20862 (N_20862,N_16286,N_16246);
nand U20863 (N_20863,N_18231,N_15911);
nand U20864 (N_20864,N_17706,N_17427);
xnor U20865 (N_20865,N_18073,N_15201);
xor U20866 (N_20866,N_18723,N_17494);
xnor U20867 (N_20867,N_16313,N_19881);
nand U20868 (N_20868,N_16096,N_15942);
xor U20869 (N_20869,N_19439,N_16893);
and U20870 (N_20870,N_16835,N_16265);
nor U20871 (N_20871,N_15970,N_18738);
nor U20872 (N_20872,N_19449,N_17402);
and U20873 (N_20873,N_18910,N_17595);
and U20874 (N_20874,N_16378,N_18493);
nand U20875 (N_20875,N_19595,N_17157);
or U20876 (N_20876,N_15186,N_15513);
nand U20877 (N_20877,N_18350,N_16858);
nor U20878 (N_20878,N_16129,N_15363);
nor U20879 (N_20879,N_16201,N_19865);
xor U20880 (N_20880,N_15674,N_16162);
and U20881 (N_20881,N_19698,N_18657);
nor U20882 (N_20882,N_19176,N_18119);
nand U20883 (N_20883,N_15910,N_16440);
and U20884 (N_20884,N_15847,N_15726);
nand U20885 (N_20885,N_15399,N_17557);
nand U20886 (N_20886,N_16634,N_19663);
and U20887 (N_20887,N_18694,N_15890);
or U20888 (N_20888,N_16013,N_17019);
or U20889 (N_20889,N_18913,N_17866);
or U20890 (N_20890,N_19369,N_17960);
nand U20891 (N_20891,N_15009,N_15579);
and U20892 (N_20892,N_18377,N_15992);
or U20893 (N_20893,N_19858,N_16404);
or U20894 (N_20894,N_16214,N_16998);
and U20895 (N_20895,N_18788,N_16867);
nand U20896 (N_20896,N_19739,N_15451);
or U20897 (N_20897,N_19180,N_16565);
and U20898 (N_20898,N_17260,N_18457);
and U20899 (N_20899,N_17722,N_16575);
nor U20900 (N_20900,N_15979,N_18058);
and U20901 (N_20901,N_15733,N_15161);
nor U20902 (N_20902,N_16753,N_19994);
nand U20903 (N_20903,N_18547,N_17821);
nor U20904 (N_20904,N_19311,N_19416);
nand U20905 (N_20905,N_17746,N_17912);
nor U20906 (N_20906,N_15285,N_15118);
nor U20907 (N_20907,N_15664,N_19331);
nand U20908 (N_20908,N_18479,N_17459);
nor U20909 (N_20909,N_15102,N_15704);
and U20910 (N_20910,N_18527,N_17081);
nand U20911 (N_20911,N_17092,N_16244);
nor U20912 (N_20912,N_15521,N_15386);
and U20913 (N_20913,N_19434,N_16945);
and U20914 (N_20914,N_18854,N_16971);
and U20915 (N_20915,N_15818,N_18476);
nand U20916 (N_20916,N_19788,N_15268);
nor U20917 (N_20917,N_19333,N_16775);
nand U20918 (N_20918,N_18125,N_17845);
and U20919 (N_20919,N_16802,N_19835);
nor U20920 (N_20920,N_15806,N_17096);
xor U20921 (N_20921,N_16635,N_17449);
nand U20922 (N_20922,N_15529,N_16980);
or U20923 (N_20923,N_18258,N_19969);
nor U20924 (N_20924,N_18208,N_15717);
nor U20925 (N_20925,N_18870,N_19792);
and U20926 (N_20926,N_18081,N_19298);
nand U20927 (N_20927,N_17659,N_15644);
nor U20928 (N_20928,N_18188,N_16046);
nand U20929 (N_20929,N_18675,N_15447);
or U20930 (N_20930,N_19749,N_15018);
or U20931 (N_20931,N_18389,N_18171);
nor U20932 (N_20932,N_16043,N_18736);
and U20933 (N_20933,N_16768,N_19526);
nor U20934 (N_20934,N_15256,N_19094);
nand U20935 (N_20935,N_15204,N_17048);
xor U20936 (N_20936,N_15418,N_19443);
nor U20937 (N_20937,N_19656,N_18108);
or U20938 (N_20938,N_18855,N_19988);
nand U20939 (N_20939,N_16052,N_17851);
or U20940 (N_20940,N_15240,N_17135);
nor U20941 (N_20941,N_15323,N_19363);
or U20942 (N_20942,N_16636,N_18951);
nand U20943 (N_20943,N_15935,N_15489);
nand U20944 (N_20944,N_19769,N_17415);
nand U20945 (N_20945,N_19742,N_19856);
or U20946 (N_20946,N_19046,N_15967);
or U20947 (N_20947,N_18011,N_17947);
nand U20948 (N_20948,N_18046,N_17704);
nand U20949 (N_20949,N_15686,N_17647);
and U20950 (N_20950,N_15757,N_16989);
xnor U20951 (N_20951,N_16817,N_16594);
and U20952 (N_20952,N_15589,N_17804);
nand U20953 (N_20953,N_18532,N_15827);
or U20954 (N_20954,N_16716,N_18842);
xor U20955 (N_20955,N_15287,N_17133);
or U20956 (N_20956,N_19122,N_18926);
or U20957 (N_20957,N_15402,N_17134);
xnor U20958 (N_20958,N_16769,N_17822);
nand U20959 (N_20959,N_15132,N_16439);
or U20960 (N_20960,N_17806,N_15043);
and U20961 (N_20961,N_17269,N_15122);
xnor U20962 (N_20962,N_15155,N_18264);
nor U20963 (N_20963,N_19185,N_15825);
or U20964 (N_20964,N_17952,N_16101);
nor U20965 (N_20965,N_18480,N_19181);
xnor U20966 (N_20966,N_18136,N_15456);
nand U20967 (N_20967,N_18687,N_17575);
nand U20968 (N_20968,N_17970,N_15567);
nand U20969 (N_20969,N_16290,N_18156);
nor U20970 (N_20970,N_16002,N_17900);
and U20971 (N_20971,N_18311,N_18023);
nor U20972 (N_20972,N_17002,N_19295);
or U20973 (N_20973,N_16345,N_15517);
or U20974 (N_20974,N_15681,N_15829);
or U20975 (N_20975,N_15836,N_17166);
or U20976 (N_20976,N_17831,N_16310);
nand U20977 (N_20977,N_15625,N_16778);
or U20978 (N_20978,N_18801,N_17503);
or U20979 (N_20979,N_18365,N_19373);
or U20980 (N_20980,N_17395,N_15030);
nor U20981 (N_20981,N_17463,N_18943);
xnor U20982 (N_20982,N_17286,N_17340);
nand U20983 (N_20983,N_16083,N_18338);
nor U20984 (N_20984,N_17965,N_17137);
or U20985 (N_20985,N_15835,N_16603);
nor U20986 (N_20986,N_17187,N_16448);
nor U20987 (N_20987,N_19496,N_17627);
xor U20988 (N_20988,N_17278,N_16897);
nor U20989 (N_20989,N_18211,N_15341);
nand U20990 (N_20990,N_19327,N_17282);
nand U20991 (N_20991,N_19534,N_19833);
and U20992 (N_20992,N_15536,N_15808);
nor U20993 (N_20993,N_16725,N_16018);
nand U20994 (N_20994,N_16983,N_18403);
and U20995 (N_20995,N_19085,N_17000);
nor U20996 (N_20996,N_16978,N_15041);
nor U20997 (N_20997,N_18674,N_18824);
or U20998 (N_20998,N_15283,N_19745);
and U20999 (N_20999,N_17125,N_18580);
or U21000 (N_21000,N_17614,N_16566);
nor U21001 (N_21001,N_17475,N_15218);
nand U21002 (N_21002,N_19344,N_15697);
nor U21003 (N_21003,N_17954,N_15017);
nand U21004 (N_21004,N_15865,N_17698);
or U21005 (N_21005,N_17518,N_17858);
or U21006 (N_21006,N_17548,N_18885);
nor U21007 (N_21007,N_16128,N_18695);
and U21008 (N_21008,N_18917,N_17882);
xnor U21009 (N_21009,N_19168,N_18582);
nor U21010 (N_21010,N_17889,N_19053);
and U21011 (N_21011,N_16740,N_16930);
nor U21012 (N_21012,N_19961,N_16599);
nor U21013 (N_21013,N_15554,N_17809);
nand U21014 (N_21014,N_18539,N_16324);
nand U21015 (N_21015,N_16920,N_17399);
and U21016 (N_21016,N_18450,N_19571);
and U21017 (N_21017,N_16488,N_19684);
nand U21018 (N_21018,N_19869,N_19205);
or U21019 (N_21019,N_18203,N_16479);
nand U21020 (N_21020,N_19965,N_15162);
nand U21021 (N_21021,N_15437,N_19347);
nand U21022 (N_21022,N_15165,N_15110);
nor U21023 (N_21023,N_17290,N_17538);
xor U21024 (N_21024,N_16453,N_19255);
nand U21025 (N_21025,N_18608,N_15238);
nand U21026 (N_21026,N_16210,N_17807);
xnor U21027 (N_21027,N_19444,N_16964);
and U21028 (N_21028,N_19660,N_19250);
xnor U21029 (N_21029,N_19777,N_15292);
nand U21030 (N_21030,N_19404,N_17432);
or U21031 (N_21031,N_18345,N_19284);
or U21032 (N_21032,N_17215,N_19752);
nand U21033 (N_21033,N_15362,N_19533);
or U21034 (N_21034,N_18605,N_15051);
xor U21035 (N_21035,N_16982,N_16277);
nand U21036 (N_21036,N_15457,N_19896);
nand U21037 (N_21037,N_16281,N_15073);
nand U21038 (N_21038,N_15033,N_18263);
nand U21039 (N_21039,N_19890,N_15084);
nor U21040 (N_21040,N_16618,N_19407);
nor U21041 (N_21041,N_15634,N_16665);
nand U21042 (N_21042,N_15630,N_18084);
nand U21043 (N_21043,N_16515,N_19108);
nand U21044 (N_21044,N_16127,N_16861);
and U21045 (N_21045,N_16649,N_17146);
and U21046 (N_21046,N_19016,N_16661);
nand U21047 (N_21047,N_16292,N_16185);
xnor U21048 (N_21048,N_16424,N_15555);
and U21049 (N_21049,N_16200,N_17491);
or U21050 (N_21050,N_17380,N_19021);
nand U21051 (N_21051,N_17868,N_18569);
and U21052 (N_21052,N_15061,N_17975);
nand U21053 (N_21053,N_15902,N_19848);
or U21054 (N_21054,N_18588,N_15654);
and U21055 (N_21055,N_18057,N_16353);
nand U21056 (N_21056,N_16156,N_15401);
and U21057 (N_21057,N_19555,N_15160);
or U21058 (N_21058,N_15315,N_18002);
nand U21059 (N_21059,N_18970,N_15028);
xnor U21060 (N_21060,N_17968,N_19212);
or U21061 (N_21061,N_17291,N_15661);
nand U21062 (N_21062,N_19247,N_15221);
or U21063 (N_21063,N_19717,N_15276);
nor U21064 (N_21064,N_18795,N_19766);
or U21065 (N_21065,N_16144,N_17927);
nor U21066 (N_21066,N_19931,N_18460);
and U21067 (N_21067,N_16037,N_15854);
nand U21068 (N_21068,N_18297,N_19922);
xor U21069 (N_21069,N_17461,N_17710);
nand U21070 (N_21070,N_18252,N_17038);
or U21071 (N_21071,N_19866,N_18704);
and U21072 (N_21072,N_18986,N_15125);
or U21073 (N_21073,N_16051,N_15741);
and U21074 (N_21074,N_18272,N_17643);
nand U21075 (N_21075,N_19402,N_17978);
xnor U21076 (N_21076,N_19689,N_16675);
nor U21077 (N_21077,N_16593,N_17553);
and U21078 (N_21078,N_17754,N_17730);
and U21079 (N_21079,N_18978,N_16813);
and U21080 (N_21080,N_17477,N_15916);
nor U21081 (N_21081,N_17599,N_15541);
xnor U21082 (N_21082,N_18997,N_15277);
or U21083 (N_21083,N_19104,N_17783);
or U21084 (N_21084,N_17309,N_19201);
nor U21085 (N_21085,N_19951,N_17165);
or U21086 (N_21086,N_17514,N_16722);
nor U21087 (N_21087,N_16886,N_15077);
or U21088 (N_21088,N_19664,N_17906);
nand U21089 (N_21089,N_19458,N_19553);
xnor U21090 (N_21090,N_19277,N_18803);
xnor U21091 (N_21091,N_17635,N_18157);
or U21092 (N_21092,N_17605,N_17561);
or U21093 (N_21093,N_19194,N_15067);
nor U21094 (N_21094,N_19243,N_17207);
or U21095 (N_21095,N_17989,N_15969);
or U21096 (N_21096,N_19665,N_15031);
and U21097 (N_21097,N_15111,N_18163);
or U21098 (N_21098,N_19628,N_16847);
nand U21099 (N_21099,N_18161,N_18629);
nor U21100 (N_21100,N_17453,N_17586);
or U21101 (N_21101,N_18571,N_16619);
nand U21102 (N_21102,N_15421,N_19597);
nand U21103 (N_21103,N_16080,N_17143);
nor U21104 (N_21104,N_16026,N_19075);
or U21105 (N_21105,N_18487,N_18568);
nor U21106 (N_21106,N_16315,N_18925);
nand U21107 (N_21107,N_19381,N_16941);
or U21108 (N_21108,N_16522,N_16844);
xor U21109 (N_21109,N_17552,N_19876);
or U21110 (N_21110,N_16758,N_15029);
and U21111 (N_21111,N_19270,N_17798);
and U21112 (N_21112,N_18614,N_18827);
xor U21113 (N_21113,N_15279,N_16079);
nand U21114 (N_21114,N_18045,N_19939);
nor U21115 (N_21115,N_18423,N_17820);
or U21116 (N_21116,N_15423,N_19336);
and U21117 (N_21117,N_18557,N_16981);
xnor U21118 (N_21118,N_16268,N_19066);
nor U21119 (N_21119,N_18720,N_16944);
nand U21120 (N_21120,N_15673,N_19891);
and U21121 (N_21121,N_18214,N_17957);
or U21122 (N_21122,N_17865,N_17241);
nand U21123 (N_21123,N_18835,N_18410);
or U21124 (N_21124,N_17270,N_17856);
nand U21125 (N_21125,N_18711,N_18549);
xnor U21126 (N_21126,N_18018,N_19537);
or U21127 (N_21127,N_19480,N_15925);
nor U21128 (N_21128,N_17861,N_19360);
nor U21129 (N_21129,N_16443,N_15000);
nor U21130 (N_21130,N_18882,N_19839);
and U21131 (N_21131,N_19560,N_18937);
and U21132 (N_21132,N_19264,N_19495);
nand U21133 (N_21133,N_15596,N_18807);
nor U21134 (N_21134,N_19548,N_15265);
nor U21135 (N_21135,N_19740,N_18012);
or U21136 (N_21136,N_16748,N_19015);
and U21137 (N_21137,N_18102,N_15384);
or U21138 (N_21138,N_17671,N_17370);
xnor U21139 (N_21139,N_17939,N_16562);
and U21140 (N_21140,N_17864,N_19903);
nand U21141 (N_21141,N_17195,N_17348);
xnor U21142 (N_21142,N_16849,N_19995);
nor U21143 (N_21143,N_19128,N_16685);
nand U21144 (N_21144,N_16131,N_15300);
nor U21145 (N_21145,N_19354,N_19365);
or U21146 (N_21146,N_19340,N_18814);
nor U21147 (N_21147,N_17755,N_15669);
nand U21148 (N_21148,N_18316,N_17528);
and U21149 (N_21149,N_19156,N_17938);
and U21150 (N_21150,N_18372,N_17931);
nor U21151 (N_21151,N_15475,N_15901);
or U21152 (N_21152,N_18555,N_17986);
or U21153 (N_21153,N_16752,N_17297);
and U21154 (N_21154,N_19112,N_18087);
and U21155 (N_21155,N_19621,N_19976);
or U21156 (N_21156,N_16304,N_15411);
or U21157 (N_21157,N_18168,N_18616);
xnor U21158 (N_21158,N_15624,N_19783);
nor U21159 (N_21159,N_15467,N_19998);
nor U21160 (N_21160,N_18618,N_17702);
nor U21161 (N_21161,N_15527,N_17761);
or U21162 (N_21162,N_16386,N_16357);
or U21163 (N_21163,N_16227,N_17945);
and U21164 (N_21164,N_17843,N_15145);
nor U21165 (N_21165,N_18274,N_18713);
or U21166 (N_21166,N_16907,N_16876);
nor U21167 (N_21167,N_18343,N_15196);
xor U21168 (N_21168,N_18928,N_18221);
and U21169 (N_21169,N_18494,N_16772);
xnor U21170 (N_21170,N_18032,N_15777);
nor U21171 (N_21171,N_15231,N_19868);
nor U21172 (N_21172,N_19235,N_17136);
or U21173 (N_21173,N_16283,N_16098);
or U21174 (N_21174,N_15972,N_16392);
nor U21175 (N_21175,N_19111,N_17124);
nand U21176 (N_21176,N_16568,N_16669);
xor U21177 (N_21177,N_18914,N_16473);
or U21178 (N_21178,N_16554,N_17610);
xnor U21179 (N_21179,N_17792,N_19627);
and U21180 (N_21180,N_17484,N_18941);
or U21181 (N_21181,N_15803,N_16092);
nor U21182 (N_21182,N_16348,N_18520);
xnor U21183 (N_21183,N_18641,N_18437);
or U21184 (N_21184,N_18075,N_15434);
or U21185 (N_21185,N_16832,N_16203);
xnor U21186 (N_21186,N_15076,N_18899);
or U21187 (N_21187,N_16943,N_18790);
nand U21188 (N_21188,N_15687,N_19491);
nor U21189 (N_21189,N_18968,N_19758);
nor U21190 (N_21190,N_15546,N_19109);
and U21191 (N_21191,N_16066,N_15417);
nor U21192 (N_21192,N_18575,N_17630);
nor U21193 (N_21193,N_17766,N_16234);
or U21194 (N_21194,N_16516,N_17668);
nand U21195 (N_21195,N_17711,N_15864);
nor U21196 (N_21196,N_15462,N_18286);
or U21197 (N_21197,N_17109,N_19079);
nor U21198 (N_21198,N_17894,N_16125);
nor U21199 (N_21199,N_18160,N_19874);
xnor U21200 (N_21200,N_18892,N_19764);
or U21201 (N_21201,N_17084,N_19368);
nor U21202 (N_21202,N_16770,N_15628);
and U21203 (N_21203,N_18165,N_17107);
or U21204 (N_21204,N_16165,N_17425);
nor U21205 (N_21205,N_15941,N_17121);
and U21206 (N_21206,N_16376,N_15722);
nand U21207 (N_21207,N_15907,N_15797);
nor U21208 (N_21208,N_19778,N_18726);
and U21209 (N_21209,N_18940,N_15272);
nand U21210 (N_21210,N_18116,N_17204);
and U21211 (N_21211,N_16081,N_16597);
nor U21212 (N_21212,N_15478,N_15334);
and U21213 (N_21213,N_16147,N_16773);
or U21214 (N_21214,N_19013,N_19010);
nor U21215 (N_21215,N_16865,N_18749);
xnor U21216 (N_21216,N_19583,N_18335);
nand U21217 (N_21217,N_19528,N_19626);
nor U21218 (N_21218,N_19316,N_19341);
and U21219 (N_21219,N_17010,N_18034);
and U21220 (N_21220,N_16299,N_17100);
and U21221 (N_21221,N_18544,N_17969);
nor U21222 (N_21222,N_18074,N_19655);
or U21223 (N_21223,N_18100,N_17252);
xnor U21224 (N_21224,N_19790,N_17158);
and U21225 (N_21225,N_19050,N_19191);
xnor U21226 (N_21226,N_17624,N_18225);
and U21227 (N_21227,N_18248,N_19501);
nand U21228 (N_21228,N_19027,N_16426);
nor U21229 (N_21229,N_19821,N_17306);
nand U21230 (N_21230,N_15486,N_19467);
nand U21231 (N_21231,N_17085,N_15342);
and U21232 (N_21232,N_17076,N_17072);
and U21233 (N_21233,N_19805,N_19411);
or U21234 (N_21234,N_18523,N_19208);
xor U21235 (N_21235,N_15001,N_16739);
or U21236 (N_21236,N_18512,N_17626);
nand U21237 (N_21237,N_19038,N_19401);
and U21238 (N_21238,N_18962,N_16809);
nor U21239 (N_21239,N_19082,N_15091);
nor U21240 (N_21240,N_17696,N_15600);
and U21241 (N_21241,N_18172,N_15466);
nor U21242 (N_21242,N_17883,N_17852);
and U21243 (N_21243,N_17784,N_19716);
xnor U21244 (N_21244,N_19953,N_18041);
xor U21245 (N_21245,N_18995,N_18056);
and U21246 (N_21246,N_18758,N_17323);
xor U21247 (N_21247,N_19033,N_15197);
and U21248 (N_21248,N_19134,N_17454);
nand U21249 (N_21249,N_18021,N_16352);
and U21250 (N_21250,N_19465,N_17209);
or U21251 (N_21251,N_18138,N_16507);
and U21252 (N_21252,N_15647,N_15093);
and U21253 (N_21253,N_18949,N_18482);
and U21254 (N_21254,N_15151,N_19808);
and U21255 (N_21255,N_18982,N_17998);
or U21256 (N_21256,N_16871,N_15926);
nand U21257 (N_21257,N_15129,N_19851);
nand U21258 (N_21258,N_17168,N_16470);
and U21259 (N_21259,N_17150,N_18392);
or U21260 (N_21260,N_15414,N_18506);
nand U21261 (N_21261,N_18998,N_17091);
and U21262 (N_21262,N_16380,N_16391);
nand U21263 (N_21263,N_18148,N_16561);
or U21264 (N_21264,N_18850,N_17086);
or U21265 (N_21265,N_15484,N_18049);
and U21266 (N_21266,N_17723,N_19862);
and U21267 (N_21267,N_19253,N_19964);
nor U21268 (N_21268,N_15658,N_18844);
or U21269 (N_21269,N_18595,N_17650);
and U21270 (N_21270,N_18170,N_19403);
nor U21271 (N_21271,N_18352,N_17688);
nand U21272 (N_21272,N_16068,N_15863);
xor U21273 (N_21273,N_16400,N_17785);
nor U21274 (N_21274,N_18719,N_15923);
xor U21275 (N_21275,N_17949,N_18816);
or U21276 (N_21276,N_15435,N_18115);
nor U21277 (N_21277,N_16402,N_17316);
or U21278 (N_21278,N_16664,N_16241);
and U21279 (N_21279,N_17219,N_15069);
and U21280 (N_21280,N_17560,N_17547);
nor U21281 (N_21281,N_18967,N_15525);
nor U21282 (N_21282,N_19029,N_16523);
nand U21283 (N_21283,N_16754,N_17047);
nand U21284 (N_21284,N_18976,N_19114);
nand U21285 (N_21285,N_15511,N_18958);
nand U21286 (N_21286,N_15438,N_15128);
and U21287 (N_21287,N_19222,N_18587);
nand U21288 (N_21288,N_17256,N_19511);
nand U21289 (N_21289,N_19469,N_17328);
or U21290 (N_21290,N_19293,N_18533);
nor U21291 (N_21291,N_15356,N_19543);
nor U21292 (N_21292,N_16582,N_18285);
nand U21293 (N_21293,N_17621,N_18217);
or U21294 (N_21294,N_19462,N_16557);
and U21295 (N_21295,N_19701,N_15823);
xnor U21296 (N_21296,N_19845,N_18603);
or U21297 (N_21297,N_19169,N_15095);
and U21298 (N_21298,N_17676,N_18401);
or U21299 (N_21299,N_17342,N_15205);
or U21300 (N_21300,N_18066,N_18348);
and U21301 (N_21301,N_18994,N_18453);
nand U21302 (N_21302,N_19771,N_16126);
nand U21303 (N_21303,N_18780,N_16360);
and U21304 (N_21304,N_17524,N_18303);
nor U21305 (N_21305,N_17651,N_17789);
nor U21306 (N_21306,N_15458,N_18524);
nor U21307 (N_21307,N_16877,N_15445);
and U21308 (N_21308,N_18275,N_17485);
xor U21309 (N_21309,N_18094,N_17276);
and U21310 (N_21310,N_17899,N_17240);
nand U21311 (N_21311,N_15531,N_16097);
and U21312 (N_21312,N_19714,N_17983);
nor U21313 (N_21313,N_17932,N_19970);
or U21314 (N_21314,N_15470,N_19601);
nor U21315 (N_21315,N_17389,N_15662);
and U21316 (N_21316,N_18522,N_19518);
nand U21317 (N_21317,N_17066,N_15678);
nor U21318 (N_21318,N_18819,N_17386);
nand U21319 (N_21319,N_19283,N_15215);
xnor U21320 (N_21320,N_15144,N_16631);
nand U21321 (N_21321,N_18781,N_19616);
and U21322 (N_21322,N_19018,N_16956);
nor U21323 (N_21323,N_16118,N_19756);
nand U21324 (N_21324,N_17375,N_17833);
and U21325 (N_21325,N_15720,N_18083);
nand U21326 (N_21326,N_15291,N_16766);
nor U21327 (N_21327,N_15065,N_16587);
and U21328 (N_21328,N_17007,N_16248);
and U21329 (N_21329,N_16620,N_15810);
xnor U21330 (N_21330,N_15587,N_17305);
nand U21331 (N_21331,N_17951,N_18030);
and U21332 (N_21332,N_15108,N_16300);
nor U21333 (N_21333,N_19672,N_15943);
nand U21334 (N_21334,N_18659,N_15298);
and U21335 (N_21335,N_17876,N_15642);
nand U21336 (N_21336,N_18755,N_17590);
nor U21337 (N_21337,N_19724,N_19978);
nor U21338 (N_21338,N_19606,N_19189);
nor U21339 (N_21339,N_18572,N_15109);
nor U21340 (N_21340,N_19451,N_16276);
xnor U21341 (N_21341,N_19497,N_17355);
and U21342 (N_21342,N_19958,N_15297);
nor U21343 (N_21343,N_15920,N_16334);
nand U21344 (N_21344,N_17251,N_17748);
nand U21345 (N_21345,N_19259,N_15891);
or U21346 (N_21346,N_15817,N_16646);
xor U21347 (N_21347,N_19807,N_18769);
nor U21348 (N_21348,N_18697,N_19926);
xor U21349 (N_21349,N_19669,N_16598);
xnor U21350 (N_21350,N_16795,N_15477);
and U21351 (N_21351,N_15667,N_16645);
nand U21352 (N_21352,N_15278,N_18033);
xor U21353 (N_21353,N_15335,N_15510);
nor U21354 (N_21354,N_16184,N_16225);
or U21355 (N_21355,N_15289,N_16012);
and U21356 (N_21356,N_16616,N_15420);
and U21357 (N_21357,N_18340,N_17919);
or U21358 (N_21358,N_18067,N_18060);
or U21359 (N_21359,N_18647,N_17113);
or U21360 (N_21360,N_18206,N_16322);
or U21361 (N_21361,N_17690,N_19224);
nand U21362 (N_21362,N_17823,N_17108);
nand U21363 (N_21363,N_15316,N_17167);
or U21364 (N_21364,N_17727,N_19948);
and U21365 (N_21365,N_16580,N_19271);
or U21366 (N_21366,N_16325,N_15798);
nand U21367 (N_21367,N_17274,N_19918);
and U21368 (N_21368,N_16422,N_17353);
nor U21369 (N_21369,N_19850,N_19430);
nand U21370 (N_21370,N_15371,N_15193);
nand U21371 (N_21371,N_16771,N_17174);
nor U21372 (N_21372,N_19154,N_16672);
or U21373 (N_21373,N_15159,N_18367);
and U21374 (N_21374,N_19121,N_15690);
nand U21375 (N_21375,N_16229,N_16111);
nor U21376 (N_21376,N_18504,N_19639);
or U21377 (N_21377,N_16420,N_15049);
or U21378 (N_21378,N_18154,N_18190);
or U21379 (N_21379,N_15313,N_16604);
or U21380 (N_21380,N_16059,N_19863);
xor U21381 (N_21381,N_15042,N_15449);
xor U21382 (N_21382,N_18812,N_16425);
or U21383 (N_21383,N_17466,N_15097);
xor U21384 (N_21384,N_18919,N_17127);
and U21385 (N_21385,N_17716,N_15971);
and U21386 (N_21386,N_18832,N_16571);
nor U21387 (N_21387,N_18408,N_17615);
nand U21388 (N_21388,N_18400,N_18939);
or U21389 (N_21389,N_16916,N_16146);
and U21390 (N_21390,N_18137,N_18834);
and U21391 (N_21391,N_17981,N_17385);
or U21392 (N_21392,N_16746,N_15500);
or U21393 (N_21393,N_16779,N_17021);
nor U21394 (N_21394,N_18654,N_17596);
xnor U21395 (N_21395,N_16320,N_16997);
nor U21396 (N_21396,N_16342,N_16282);
and U21397 (N_21397,N_16082,N_17243);
or U21398 (N_21398,N_16666,N_19482);
or U21399 (N_21399,N_16073,N_15837);
nor U21400 (N_21400,N_16572,N_18038);
nand U21401 (N_21401,N_18847,N_16011);
nor U21402 (N_21402,N_17013,N_19617);
xor U21403 (N_21403,N_16123,N_16389);
nor U21404 (N_21404,N_18475,N_18134);
nor U21405 (N_21405,N_18461,N_17765);
and U21406 (N_21406,N_19765,N_16638);
and U21407 (N_21407,N_18977,N_17065);
and U21408 (N_21408,N_16658,N_15966);
nor U21409 (N_21409,N_18260,N_15104);
xnor U21410 (N_21410,N_17314,N_18890);
and U21411 (N_21411,N_17005,N_18354);
nor U21412 (N_21412,N_17887,N_15345);
and U21413 (N_21413,N_19452,N_15610);
and U21414 (N_21414,N_17638,N_19074);
nand U21415 (N_21415,N_18387,N_17401);
nor U21416 (N_21416,N_15922,N_15226);
xnor U21417 (N_21417,N_16808,N_18860);
nand U21418 (N_21418,N_16767,N_18464);
nand U21419 (N_21419,N_15626,N_15227);
nor U21420 (N_21420,N_16472,N_16176);
nor U21421 (N_21421,N_16181,N_17322);
and U21422 (N_21422,N_17233,N_15737);
nand U21423 (N_21423,N_15734,N_15134);
xor U21424 (N_21424,N_17423,N_19172);
nor U21425 (N_21425,N_18256,N_17070);
nand U21426 (N_21426,N_18938,N_18483);
nand U21427 (N_21427,N_16259,N_15431);
or U21428 (N_21428,N_18282,N_16505);
nand U21429 (N_21429,N_19967,N_16242);
and U21430 (N_21430,N_17430,N_15203);
xnor U21431 (N_21431,N_17556,N_16388);
and U21432 (N_21432,N_15960,N_19376);
nor U21433 (N_21433,N_16698,N_16368);
and U21434 (N_21434,N_19030,N_17832);
and U21435 (N_21435,N_15873,N_18710);
or U21436 (N_21436,N_17697,N_18481);
and U21437 (N_21437,N_19474,N_17210);
nor U21438 (N_21438,N_15173,N_18772);
or U21439 (N_21439,N_19445,N_17177);
xnor U21440 (N_21440,N_19358,N_16175);
and U21441 (N_21441,N_17142,N_16359);
nor U21442 (N_21442,N_15089,N_15360);
nand U21443 (N_21443,N_17611,N_17333);
or U21444 (N_21444,N_15945,N_16890);
xor U21445 (N_21445,N_15735,N_16466);
xor U21446 (N_21446,N_19267,N_19088);
nand U21447 (N_21447,N_19197,N_19410);
nor U21448 (N_21448,N_19513,N_16217);
or U21449 (N_21449,N_17982,N_19817);
and U21450 (N_21450,N_17492,N_17279);
nand U21451 (N_21451,N_15410,N_17616);
and U21452 (N_21452,N_17235,N_16307);
nand U21453 (N_21453,N_19535,N_17999);
or U21454 (N_21454,N_15844,N_16206);
nand U21455 (N_21455,N_15776,N_15322);
nand U21456 (N_21456,N_19383,N_16161);
nand U21457 (N_21457,N_16517,N_17911);
and U21458 (N_21458,N_19755,N_17405);
nand U21459 (N_21459,N_19754,N_19806);
nand U21460 (N_21460,N_15126,N_15190);
xnor U21461 (N_21461,N_18229,N_17409);
or U21462 (N_21462,N_18474,N_18386);
xor U21463 (N_21463,N_17959,N_15957);
or U21464 (N_21464,N_16853,N_19147);
xor U21465 (N_21465,N_15739,N_16120);
nor U21466 (N_21466,N_19776,N_19317);
or U21467 (N_21467,N_18863,N_15098);
nand U21468 (N_21468,N_16883,N_15148);
nor U21469 (N_21469,N_18329,N_16578);
nand U21470 (N_21470,N_19952,N_15534);
nor U21471 (N_21471,N_16278,N_16984);
xor U21472 (N_21472,N_18514,N_16966);
nand U21473 (N_21473,N_18141,N_19226);
or U21474 (N_21474,N_18665,N_18417);
nand U21475 (N_21475,N_17372,N_18266);
xor U21476 (N_21476,N_18247,N_17261);
nor U21477 (N_21477,N_17345,N_15333);
or U21478 (N_21478,N_18669,N_16816);
and U21479 (N_21479,N_19530,N_18331);
nand U21480 (N_21480,N_19767,N_19276);
and U21481 (N_21481,N_16639,N_19521);
and U21482 (N_21482,N_16509,N_18036);
and U21483 (N_21483,N_18308,N_16673);
nand U21484 (N_21484,N_19620,N_19658);
or U21485 (N_21485,N_18333,N_16948);
nor U21486 (N_21486,N_15535,N_16642);
and U21487 (N_21487,N_19493,N_19218);
and U21488 (N_21488,N_16991,N_17196);
or U21489 (N_21489,N_16600,N_19314);
or U21490 (N_21490,N_17725,N_17636);
nand U21491 (N_21491,N_17426,N_16390);
nand U21492 (N_21492,N_15263,N_18624);
nor U21493 (N_21493,N_18667,N_19618);
nor U21494 (N_21494,N_19263,N_19320);
or U21495 (N_21495,N_17006,N_15304);
and U21496 (N_21496,N_17460,N_15206);
xor U21497 (N_21497,N_18499,N_19895);
and U21498 (N_21498,N_18319,N_15224);
nor U21499 (N_21499,N_15072,N_18194);
nand U21500 (N_21500,N_17920,N_19798);
nand U21501 (N_21501,N_16803,N_17149);
nand U21502 (N_21502,N_17753,N_18357);
nor U21503 (N_21503,N_16364,N_15074);
nand U21504 (N_21504,N_16044,N_15509);
nand U21505 (N_21505,N_18902,N_17848);
and U21506 (N_21506,N_18431,N_19379);
or U21507 (N_21507,N_16100,N_15407);
or U21508 (N_21508,N_16410,N_17088);
and U21509 (N_21509,N_16929,N_15243);
nand U21510 (N_21510,N_18961,N_15136);
nor U21511 (N_21511,N_15565,N_16701);
nor U21512 (N_21512,N_16530,N_18379);
nand U21513 (N_21513,N_19624,N_19309);
and U21514 (N_21514,N_19380,N_19894);
nand U21515 (N_21515,N_16484,N_15795);
or U21516 (N_21516,N_18127,N_15794);
or U21517 (N_21517,N_19026,N_15050);
nand U21518 (N_21518,N_16192,N_19417);
nor U21519 (N_21519,N_17295,N_17946);
nor U21520 (N_21520,N_17094,N_17824);
or U21521 (N_21521,N_18954,N_18176);
and U21522 (N_21522,N_19780,N_15340);
and U21523 (N_21523,N_18085,N_17505);
xnor U21524 (N_21524,N_18778,N_17472);
nor U21525 (N_21525,N_19055,N_16707);
and U21526 (N_21526,N_16284,N_16710);
nand U21527 (N_21527,N_18328,N_16836);
and U21528 (N_21528,N_15480,N_16255);
nor U21529 (N_21529,N_17666,N_18886);
or U21530 (N_21530,N_19719,N_16924);
or U21531 (N_21531,N_15404,N_19596);
and U21532 (N_21532,N_17031,N_18912);
nor U21533 (N_21533,N_15191,N_16846);
nand U21534 (N_21534,N_17767,N_17918);
nor U21535 (N_21535,N_18983,N_18810);
or U21536 (N_21536,N_19735,N_15828);
or U21537 (N_21537,N_18957,N_15403);
nor U21538 (N_21538,N_19989,N_17891);
xnor U21539 (N_21539,N_17700,N_15066);
xor U21540 (N_21540,N_17914,N_17377);
xor U21541 (N_21541,N_19328,N_15493);
and U21542 (N_21542,N_18893,N_15549);
and U21543 (N_21543,N_17908,N_18717);
nor U21544 (N_21544,N_15850,N_19391);
nand U21545 (N_21545,N_16976,N_17587);
nor U21546 (N_21546,N_18841,N_19105);
nor U21547 (N_21547,N_15948,N_15105);
nand U21548 (N_21548,N_16617,N_17499);
nor U21549 (N_21549,N_17570,N_19068);
or U21550 (N_21550,N_17618,N_19584);
and U21551 (N_21551,N_15620,N_17358);
and U21552 (N_21552,N_15955,N_18538);
nand U21553 (N_21553,N_17535,N_16039);
nor U21554 (N_21554,N_17110,N_18945);
and U21555 (N_21555,N_15382,N_16629);
and U21556 (N_21556,N_18003,N_15488);
and U21557 (N_21557,N_17212,N_17827);
nand U21558 (N_21558,N_15216,N_18785);
nor U21559 (N_21559,N_15454,N_15119);
or U21560 (N_21560,N_15886,N_17691);
xor U21561 (N_21561,N_15185,N_15711);
xnor U21562 (N_21562,N_17277,N_18837);
nor U21563 (N_21563,N_19278,N_19902);
nand U21564 (N_21564,N_17974,N_19428);
nor U21565 (N_21565,N_15011,N_16841);
nor U21566 (N_21566,N_18578,N_19507);
nor U21567 (N_21567,N_15490,N_15885);
or U21568 (N_21568,N_15839,N_19527);
nand U21569 (N_21569,N_18179,N_17188);
and U21570 (N_21570,N_19982,N_16860);
nor U21571 (N_21571,N_19775,N_18740);
or U21572 (N_21572,N_16070,N_16539);
and U21573 (N_21573,N_18467,N_16197);
and U21574 (N_21574,N_18871,N_15601);
or U21575 (N_21575,N_17057,N_19183);
and U21576 (N_21576,N_18471,N_15507);
and U21577 (N_21577,N_18210,N_17046);
and U21578 (N_21578,N_15412,N_16435);
xor U21579 (N_21579,N_17495,N_17445);
or U21580 (N_21580,N_19598,N_17897);
or U21581 (N_21581,N_18932,N_16149);
nand U21582 (N_21582,N_17221,N_19017);
nand U21583 (N_21583,N_15027,N_16179);
and U21584 (N_21584,N_15314,N_15745);
nor U21585 (N_21585,N_17293,N_17465);
nand U21586 (N_21586,N_16682,N_17591);
nand U21587 (N_21587,N_19900,N_16494);
nor U21588 (N_21588,N_15115,N_17433);
and U21589 (N_21589,N_19132,N_17281);
and U21590 (N_21590,N_15192,N_17606);
or U21591 (N_21591,N_19944,N_19707);
or U21592 (N_21592,N_16881,N_17631);
and U21593 (N_21593,N_15540,N_18505);
nor U21594 (N_21594,N_18518,N_18055);
nand U21595 (N_21595,N_16415,N_17814);
and U21596 (N_21596,N_18894,N_17237);
and U21597 (N_21597,N_15900,N_15668);
and U21598 (N_21598,N_15657,N_15580);
and U21599 (N_21599,N_18813,N_15962);
nor U21600 (N_21600,N_15522,N_16153);
nor U21601 (N_21601,N_19065,N_19551);
nand U21602 (N_21602,N_16140,N_18404);
and U21603 (N_21603,N_16199,N_15498);
nor U21604 (N_21604,N_16481,N_16528);
and U21605 (N_21605,N_15881,N_17056);
xnor U21606 (N_21606,N_15616,N_17197);
nand U21607 (N_21607,N_16535,N_17966);
and U21608 (N_21608,N_18419,N_16475);
or U21609 (N_21609,N_19529,N_17347);
nand U21610 (N_21610,N_15368,N_18843);
or U21611 (N_21611,N_15075,N_18747);
nor U21612 (N_21612,N_15121,N_19315);
nor U21613 (N_21613,N_16009,N_19979);
or U21614 (N_21614,N_15299,N_15320);
xnor U21615 (N_21615,N_17569,N_16471);
nand U21616 (N_21616,N_16025,N_19632);
or U21617 (N_21617,N_15078,N_15671);
nor U21618 (N_21618,N_18130,N_15715);
or U21619 (N_21619,N_15695,N_15428);
or U21620 (N_21620,N_18299,N_19631);
nor U21621 (N_21621,N_19506,N_15607);
or U21622 (N_21622,N_19826,N_16331);
and U21623 (N_21623,N_15021,N_18602);
and U21624 (N_21624,N_19880,N_15346);
nor U21625 (N_21625,N_18846,N_18741);
or U21626 (N_21626,N_15723,N_19812);
or U21627 (N_21627,N_17351,N_17910);
nand U21628 (N_21628,N_16615,N_19206);
or U21629 (N_21629,N_19854,N_16430);
and U21630 (N_21630,N_16644,N_15094);
or U21631 (N_21631,N_16202,N_16918);
nor U21632 (N_21632,N_17238,N_19937);
and U21633 (N_21633,N_16513,N_18903);
xnor U21634 (N_21634,N_17652,N_17073);
nor U21635 (N_21635,N_17654,N_19857);
nor U21636 (N_21636,N_17153,N_17064);
nor U21637 (N_21637,N_18767,N_16621);
or U21638 (N_21638,N_15087,N_18609);
or U21639 (N_21639,N_17510,N_16733);
nand U21640 (N_21640,N_19490,N_19399);
and U21641 (N_21641,N_18470,N_15305);
nor U21642 (N_21642,N_16972,N_18666);
nor U21643 (N_21643,N_15267,N_17541);
and U21644 (N_21644,N_15677,N_18545);
and U21645 (N_21645,N_16085,N_15427);
or U21646 (N_21646,N_17320,N_19818);
or U21647 (N_21647,N_18562,N_16280);
xor U21648 (N_21648,N_18548,N_18022);
or U21649 (N_21649,N_17450,N_18370);
and U21650 (N_21650,N_15694,N_15080);
nand U21651 (N_21651,N_18488,N_15153);
or U21652 (N_21652,N_15217,N_16633);
and U21653 (N_21653,N_18852,N_17390);
nor U21654 (N_21654,N_17943,N_15632);
nor U21655 (N_21655,N_15756,N_17364);
nand U21656 (N_21656,N_17829,N_18358);
nand U21657 (N_21657,N_19668,N_17349);
xor U21658 (N_21658,N_16894,N_16719);
nor U21659 (N_21659,N_19525,N_17504);
or U21660 (N_21660,N_19843,N_15636);
nor U21661 (N_21661,N_19549,N_17794);
nand U21662 (N_21662,N_18442,N_19841);
or U21663 (N_21663,N_19968,N_15239);
and U21664 (N_21664,N_17213,N_15980);
xnor U21665 (N_21665,N_15729,N_19622);
xnor U21666 (N_21666,N_16589,N_15659);
and U21667 (N_21667,N_15167,N_17089);
or U21668 (N_21668,N_15103,N_15515);
xor U21669 (N_21669,N_17462,N_19051);
nand U21670 (N_21670,N_17192,N_18701);
nor U21671 (N_21671,N_19308,N_16878);
and U21672 (N_21672,N_19834,N_19901);
or U21673 (N_21673,N_18152,N_17299);
nor U21674 (N_21674,N_18599,N_18001);
or U21675 (N_21675,N_15631,N_18673);
or U21676 (N_21676,N_18888,N_17313);
or U21677 (N_21677,N_16859,N_17838);
or U21678 (N_21678,N_15181,N_18671);
nor U21679 (N_21679,N_16640,N_16663);
nand U21680 (N_21680,N_19700,N_17410);
or U21681 (N_21681,N_16288,N_19086);
nand U21682 (N_21682,N_16567,N_19081);
xnor U21683 (N_21683,N_19058,N_15547);
nor U21684 (N_21684,N_17227,N_18500);
and U21685 (N_21685,N_18347,N_19062);
nor U21686 (N_21686,N_16099,N_19731);
or U21687 (N_21687,N_17416,N_15107);
or U21688 (N_21688,N_16823,N_19210);
xor U21689 (N_21689,N_15003,N_19125);
and U21690 (N_21690,N_18232,N_19815);
xnor U21691 (N_21691,N_15015,N_15284);
nand U21692 (N_21692,N_19476,N_16441);
nor U21693 (N_21693,N_16937,N_18920);
nor U21694 (N_21694,N_17956,N_18473);
and U21695 (N_21695,N_18606,N_18996);
or U21696 (N_21696,N_16167,N_15996);
or U21697 (N_21697,N_19546,N_19394);
nor U21698 (N_21698,N_15389,N_15135);
or U21699 (N_21699,N_16463,N_19704);
or U21700 (N_21700,N_17004,N_18679);
or U21701 (N_21701,N_15977,N_19450);
xnor U21702 (N_21702,N_19750,N_17234);
and U21703 (N_21703,N_18445,N_16193);
xnor U21704 (N_21704,N_15319,N_18434);
and U21705 (N_21705,N_16942,N_18456);
nor U21706 (N_21706,N_17649,N_19192);
or U21707 (N_21707,N_16427,N_16445);
nand U21708 (N_21708,N_19020,N_18744);
nor U21709 (N_21709,N_18035,N_15933);
nand U21710 (N_21710,N_19697,N_15763);
nand U21711 (N_21711,N_18771,N_16186);
nand U21712 (N_21712,N_19448,N_18063);
xnor U21713 (N_21713,N_17513,N_17732);
or U21714 (N_21714,N_18305,N_16180);
nor U21715 (N_21715,N_17549,N_19609);
or U21716 (N_21716,N_15426,N_17715);
or U21717 (N_21717,N_15068,N_16164);
or U21718 (N_21718,N_16511,N_16714);
nor U21719 (N_21719,N_16062,N_15198);
nand U21720 (N_21720,N_19762,N_16442);
nor U21721 (N_21721,N_16045,N_19940);
nand U21722 (N_21722,N_16676,N_18543);
and U21723 (N_21723,N_16050,N_15767);
xor U21724 (N_21724,N_16142,N_18567);
or U21725 (N_21725,N_16612,N_19456);
and U21726 (N_21726,N_17793,N_19301);
or U21727 (N_21727,N_18722,N_17003);
nand U21728 (N_21728,N_19089,N_15286);
and U21729 (N_21729,N_16213,N_17830);
nor U21730 (N_21730,N_15764,N_19640);
xnor U21731 (N_21731,N_18867,N_18596);
nor U21732 (N_21732,N_15251,N_16783);
nand U21733 (N_21733,N_16674,N_16837);
nand U21734 (N_21734,N_19746,N_17726);
and U21735 (N_21735,N_17035,N_15702);
or U21736 (N_21736,N_18375,N_18881);
and U21737 (N_21737,N_18131,N_15595);
or U21738 (N_21738,N_19422,N_19432);
xnor U21739 (N_21739,N_16273,N_16060);
or U21740 (N_21740,N_19973,N_18828);
nor U21741 (N_21741,N_16995,N_17810);
nor U21742 (N_21742,N_16749,N_19024);
or U21743 (N_21743,N_18859,N_16643);
or U21744 (N_21744,N_17283,N_17067);
nor U21745 (N_21745,N_17934,N_17795);
or U21746 (N_21746,N_16236,N_16010);
and U21747 (N_21747,N_17398,N_17877);
nand U21748 (N_21748,N_18428,N_18683);
nand U21749 (N_21749,N_17103,N_19463);
and U21750 (N_21750,N_19565,N_18093);
or U21751 (N_21751,N_17128,N_18963);
nor U21752 (N_21752,N_16027,N_15325);
nand U21753 (N_21753,N_19929,N_18581);
or U21754 (N_21754,N_15442,N_18142);
nand U21755 (N_21755,N_15855,N_15849);
and U21756 (N_21756,N_15937,N_19100);
nor U21757 (N_21757,N_17648,N_17479);
nand U21758 (N_21758,N_18284,N_19594);
and U21759 (N_21759,N_15710,N_17522);
and U21760 (N_21760,N_16863,N_18628);
nand U21761 (N_21761,N_16168,N_16030);
or U21762 (N_21762,N_17903,N_18598);
or U21763 (N_21763,N_18213,N_15485);
and U21764 (N_21764,N_18222,N_16790);
and U21765 (N_21765,N_15869,N_17216);
or U21766 (N_21766,N_17447,N_19325);
or U21767 (N_21767,N_18187,N_15769);
nor U21768 (N_21768,N_19794,N_16979);
and U21769 (N_21769,N_17414,N_16909);
or U21770 (N_21770,N_16856,N_15070);
nand U21771 (N_21771,N_18186,N_16655);
xor U21772 (N_21772,N_19679,N_17082);
nor U21773 (N_21773,N_19954,N_18829);
and U21774 (N_21774,N_18751,N_16819);
nand U21775 (N_21775,N_17222,N_18432);
nand U21776 (N_21776,N_17406,N_18025);
nand U21777 (N_21777,N_16335,N_19043);
nor U21778 (N_21778,N_19692,N_18107);
and U21779 (N_21779,N_15708,N_18092);
xor U21780 (N_21780,N_18317,N_19440);
or U21781 (N_21781,N_19182,N_16708);
and U21782 (N_21782,N_17029,N_18786);
or U21783 (N_21783,N_19257,N_17059);
and U21784 (N_21784,N_18202,N_19955);
nor U21785 (N_21785,N_18459,N_17724);
nand U21786 (N_21786,N_15266,N_15884);
nand U21787 (N_21787,N_16004,N_17431);
nand U21788 (N_21788,N_17287,N_15689);
or U21789 (N_21789,N_15908,N_15747);
and U21790 (N_21790,N_16151,N_15929);
and U21791 (N_21791,N_15040,N_19136);
or U21792 (N_21792,N_15034,N_16160);
nand U21793 (N_21793,N_17078,N_16624);
or U21794 (N_21794,N_16731,N_17869);
nand U21795 (N_21795,N_19006,N_15349);
nand U21796 (N_21796,N_18838,N_16875);
xor U21797 (N_21797,N_15785,N_16191);
and U21798 (N_21798,N_17567,N_19153);
nor U21799 (N_21799,N_16374,N_16411);
and U21800 (N_21800,N_18444,N_18942);
xor U21801 (N_21801,N_18039,N_18315);
and U21802 (N_21802,N_15416,N_15425);
nand U21803 (N_21803,N_19879,N_18330);
and U21804 (N_21804,N_16812,N_16398);
or U21805 (N_21805,N_19215,N_18259);
or U21806 (N_21806,N_16232,N_16552);
xnor U21807 (N_21807,N_17592,N_19625);
xor U21808 (N_21808,N_16387,N_18204);
and U21809 (N_21809,N_19586,N_19069);
nand U21810 (N_21810,N_19972,N_18502);
and U21811 (N_21811,N_19461,N_15229);
nor U21812 (N_21812,N_17701,N_19269);
nor U21813 (N_21813,N_15746,N_17300);
or U21814 (N_21814,N_18546,N_17354);
or U21815 (N_21815,N_18633,N_19353);
xor U21816 (N_21816,N_18965,N_17871);
nand U21817 (N_21817,N_15372,N_18916);
xor U21818 (N_21818,N_19706,N_16656);
nand U21819 (N_21819,N_18924,N_18644);
and U21820 (N_21820,N_16477,N_15037);
or U21821 (N_21821,N_18594,N_16428);
xnor U21822 (N_21822,N_19306,N_17408);
nor U21823 (N_21823,N_19120,N_17613);
and U21824 (N_21824,N_15158,N_16110);
nor U21825 (N_21825,N_19041,N_19330);
or U21826 (N_21826,N_17902,N_16394);
or U21827 (N_21827,N_19864,N_18261);
and U21828 (N_21828,N_19460,N_15879);
nor U21829 (N_21829,N_19357,N_15377);
nor U21830 (N_21830,N_19146,N_18278);
or U21831 (N_21831,N_17111,N_16705);
nand U21832 (N_21832,N_16446,N_19721);
nand U21833 (N_21833,N_16382,N_17886);
xor U21834 (N_21834,N_15086,N_18126);
nor U21835 (N_21835,N_15530,N_15750);
nor U21836 (N_21836,N_17742,N_19980);
nor U21837 (N_21837,N_16135,N_18921);
or U21838 (N_21838,N_16810,N_15099);
or U21839 (N_21839,N_18752,N_16761);
nor U21840 (N_21840,N_15532,N_19095);
and U21841 (N_21841,N_19733,N_15200);
nor U21842 (N_21842,N_18597,N_15149);
or U21843 (N_21843,N_19960,N_15585);
or U21844 (N_21844,N_19803,N_16105);
or U21845 (N_21845,N_18166,N_17012);
nand U21846 (N_21846,N_19517,N_19715);
xnor U21847 (N_21847,N_16171,N_17388);
and U21848 (N_21848,N_18989,N_17653);
and U21849 (N_21849,N_18374,N_17529);
or U21850 (N_21850,N_18129,N_18734);
nor U21851 (N_21851,N_18336,N_18371);
and U21852 (N_21852,N_16988,N_19789);
and U21853 (N_21853,N_16228,N_19200);
nor U21854 (N_21854,N_19004,N_17600);
nand U21855 (N_21855,N_15984,N_15830);
xor U21856 (N_21856,N_17271,N_17944);
nor U21857 (N_21857,N_19242,N_16115);
or U21858 (N_21858,N_18966,N_16936);
xnor U21859 (N_21859,N_16760,N_18026);
or U21860 (N_21860,N_16950,N_19113);
and U21861 (N_21861,N_16960,N_19028);
and U21862 (N_21862,N_16211,N_15748);
nand U21863 (N_21863,N_19196,N_17768);
nor U21864 (N_21864,N_17337,N_17739);
or U21865 (N_21865,N_16264,N_19599);
xor U21866 (N_21866,N_15973,N_16895);
nand U21867 (N_21867,N_15981,N_18268);
nand U21868 (N_21868,N_17105,N_16736);
nand U21869 (N_21869,N_16889,N_16727);
or U21870 (N_21870,N_19950,N_15698);
and U21871 (N_21871,N_18809,N_15184);
nand U21872 (N_21872,N_19034,N_17873);
or U21873 (N_21873,N_15214,N_17203);
nor U21874 (N_21874,N_17637,N_16074);
xor U21875 (N_21875,N_16258,N_16015);
nand U21876 (N_21876,N_19785,N_17312);
or U21877 (N_21877,N_19470,N_16588);
nand U21878 (N_21878,N_18869,N_19822);
nand U21879 (N_21879,N_16898,N_16913);
nand U21880 (N_21880,N_18898,N_16824);
nand U21881 (N_21881,N_16117,N_16270);
nor U21882 (N_21882,N_19623,N_16172);
xnor U21883 (N_21883,N_16150,N_18856);
xor U21884 (N_21884,N_15986,N_15990);
nor U21885 (N_21885,N_15396,N_15178);
nor U21886 (N_21886,N_19217,N_17253);
nor U21887 (N_21887,N_19711,N_18234);
nor U21888 (N_21888,N_18310,N_16955);
nand U21889 (N_21889,N_19770,N_19925);
nor U21890 (N_21890,N_16305,N_18283);
nor U21891 (N_21891,N_17298,N_15175);
and U21892 (N_21892,N_16102,N_18478);
nor U21893 (N_21893,N_17673,N_19797);
nand U21894 (N_21894,N_16818,N_15533);
nand U21895 (N_21895,N_17507,N_17288);
nand U21896 (N_21896,N_19005,N_18366);
nor U21897 (N_21897,N_19722,N_15123);
and U21898 (N_21898,N_18784,N_19710);
and U21899 (N_21899,N_15899,N_16057);
nor U21900 (N_21900,N_17604,N_16486);
xor U21901 (N_21901,N_18065,N_19279);
or U21902 (N_21902,N_15691,N_16091);
nand U21903 (N_21903,N_15760,N_18896);
and U21904 (N_21904,N_18153,N_17441);
or U21905 (N_21905,N_17835,N_18078);
or U21906 (N_21906,N_19144,N_18584);
or U21907 (N_21907,N_18952,N_17452);
nand U21908 (N_21908,N_16212,N_17147);
and U21909 (N_21909,N_16408,N_15639);
nand U21910 (N_21910,N_16416,N_19681);
nor U21911 (N_21911,N_16919,N_18712);
and U21912 (N_21912,N_16383,N_18817);
and U21913 (N_21913,N_17770,N_19178);
or U21914 (N_21914,N_17511,N_15332);
nor U21915 (N_21915,N_15858,N_17481);
and U21916 (N_21916,N_17391,N_17311);
nor U21917 (N_21917,N_18491,N_15819);
nand U21918 (N_21918,N_19962,N_16595);
xor U21919 (N_21919,N_16927,N_15262);
xnor U21920 (N_21920,N_16087,N_15497);
nand U21921 (N_21921,N_17352,N_15032);
nand U21922 (N_21922,N_15762,N_19435);
xnor U21923 (N_21923,N_15707,N_19691);
nor U21924 (N_21924,N_19137,N_19919);
xnor U21925 (N_21925,N_16902,N_17061);
and U21926 (N_21926,N_18199,N_16525);
nand U21927 (N_21927,N_18905,N_16807);
and U21928 (N_21928,N_16721,N_18692);
nor U21929 (N_21929,N_18766,N_16458);
or U21930 (N_21930,N_19607,N_18455);
nand U21931 (N_21931,N_19281,N_16502);
or U21932 (N_21932,N_15045,N_17879);
nor U21933 (N_21933,N_16031,N_17478);
nor U21934 (N_21934,N_16952,N_19498);
nor U21935 (N_21935,N_16001,N_16005);
nand U21936 (N_21936,N_16104,N_15336);
nand U21937 (N_21937,N_18746,N_15558);
nor U21938 (N_21938,N_18798,N_18312);
and U21939 (N_21939,N_18383,N_18240);
nand U21940 (N_21940,N_15288,N_15621);
nor U21941 (N_21941,N_16431,N_16095);
nor U21942 (N_21942,N_16689,N_15339);
and U21943 (N_21943,N_18774,N_19580);
nor U21944 (N_21944,N_19889,N_15059);
nor U21945 (N_21945,N_17545,N_15605);
nand U21946 (N_21946,N_18180,N_17901);
and U21947 (N_21947,N_19531,N_16627);
nand U21948 (N_21948,N_17985,N_18563);
nor U21949 (N_21949,N_19696,N_18207);
xnor U21950 (N_21950,N_19204,N_16693);
nor U21951 (N_21951,N_18324,N_19585);
nand U21952 (N_21952,N_17332,N_19256);
or U21953 (N_21953,N_16006,N_17009);
and U21954 (N_21954,N_16436,N_18236);
nor U21955 (N_21955,N_15443,N_18412);
or U21956 (N_21956,N_17194,N_16272);
nor U21957 (N_21957,N_19999,N_19468);
nand U21958 (N_21958,N_18789,N_17189);
or U21959 (N_21959,N_18262,N_16409);
nor U21960 (N_21960,N_19418,N_18181);
nor U21961 (N_21961,N_19167,N_19709);
nand U21962 (N_21962,N_19367,N_16529);
and U21963 (N_21963,N_19677,N_18655);
or U21964 (N_21964,N_15653,N_15583);
and U21965 (N_21965,N_18439,N_19040);
nand U21966 (N_21966,N_16774,N_19761);
or U21967 (N_21967,N_15550,N_16397);
nand U21968 (N_21968,N_18743,N_18496);
nor U21969 (N_21969,N_17995,N_15495);
or U21970 (N_21970,N_16630,N_19877);
nand U21971 (N_21971,N_16134,N_17338);
nand U21972 (N_21972,N_18811,N_16632);
or U21973 (N_21973,N_17075,N_15889);
nor U21974 (N_21974,N_17365,N_16469);
nor U21975 (N_21975,N_19729,N_16652);
nor U21976 (N_21976,N_15211,N_19478);
nand U21977 (N_21977,N_17193,N_15999);
and U21978 (N_21978,N_18373,N_18593);
xnor U21979 (N_21979,N_18477,N_18009);
nand U21980 (N_21980,N_16884,N_18397);
or U21981 (N_21981,N_19908,N_15940);
and U21982 (N_21982,N_17228,N_18191);
and U21983 (N_21983,N_19678,N_15232);
nand U21984 (N_21984,N_19378,N_17363);
or U21985 (N_21985,N_19254,N_17533);
nor U21986 (N_21986,N_18114,N_18944);
or U21987 (N_21987,N_17580,N_19753);
nand U21988 (N_21988,N_16821,N_18510);
and U21989 (N_21989,N_18292,N_17229);
nor U21990 (N_21990,N_18617,N_19454);
or U21991 (N_21991,N_17657,N_16183);
or U21992 (N_21992,N_19246,N_17190);
and U21993 (N_21993,N_19453,N_18302);
nor U21994 (N_21994,N_17898,N_16429);
nor U21995 (N_21995,N_16450,N_16432);
or U21996 (N_21996,N_19385,N_16403);
or U21997 (N_21997,N_15699,N_17516);
nor U21998 (N_21998,N_16679,N_16953);
and U21999 (N_21999,N_15897,N_19161);
nor U22000 (N_22000,N_15465,N_19800);
nand U22001 (N_22001,N_16780,N_18378);
nand U22002 (N_22002,N_19078,N_15928);
nand U22003 (N_22003,N_18159,N_16799);
and U22004 (N_22004,N_19840,N_18554);
nand U22005 (N_22005,N_18178,N_16223);
nand U22006 (N_22006,N_17633,N_18556);
nand U22007 (N_22007,N_16717,N_16946);
and U22008 (N_22008,N_18627,N_15127);
nand U22009 (N_22009,N_18369,N_15594);
or U22010 (N_22010,N_18019,N_16257);
xnor U22011 (N_22011,N_15258,N_17915);
nand U22012 (N_22012,N_17735,N_16651);
and U22013 (N_22013,N_19751,N_17068);
nor U22014 (N_22014,N_18558,N_18727);
nor U22015 (N_22015,N_18436,N_17928);
or U22016 (N_22016,N_15502,N_18146);
xnor U22017 (N_22017,N_18728,N_17530);
and U22018 (N_22018,N_15608,N_15709);
or U22019 (N_22019,N_18425,N_15430);
xnor U22020 (N_22020,N_16347,N_15545);
nand U22021 (N_22021,N_17302,N_16157);
or U22022 (N_22022,N_17979,N_19859);
nor U22023 (N_22023,N_19802,N_15682);
nand U22024 (N_22024,N_18950,N_17963);
nand U22025 (N_22025,N_16912,N_15905);
nand U22026 (N_22026,N_15053,N_15092);
and U22027 (N_22027,N_15366,N_18014);
and U22028 (N_22028,N_15814,N_16969);
nand U22029 (N_22029,N_16240,N_16182);
nor U22030 (N_22030,N_18117,N_15822);
nand U22031 (N_22031,N_18907,N_16885);
and U22032 (N_22032,N_16124,N_16891);
nor U22033 (N_22033,N_17487,N_17796);
and U22034 (N_22034,N_19406,N_15672);
or U22035 (N_22035,N_16088,N_16741);
nand U22036 (N_22036,N_17828,N_15528);
or U22037 (N_22037,N_16496,N_16518);
or U22038 (N_22038,N_16455,N_15016);
or U22039 (N_22039,N_17558,N_18668);
or U22040 (N_22040,N_16784,N_19611);
and U22041 (N_22041,N_15057,N_16694);
nand U22042 (N_22042,N_17396,N_15163);
and U22043 (N_22043,N_15936,N_19629);
nand U22044 (N_22044,N_15472,N_19475);
and U22045 (N_22045,N_15424,N_15244);
or U22046 (N_22046,N_18836,N_17383);
or U22047 (N_22047,N_18396,N_18216);
nor U22048 (N_22048,N_19654,N_19990);
and U22049 (N_22049,N_19214,N_15843);
xnor U22050 (N_22050,N_19577,N_16173);
or U22051 (N_22051,N_19816,N_17226);
and U22052 (N_22052,N_19387,N_17967);
and U22053 (N_22053,N_17546,N_18709);
or U22054 (N_22054,N_16294,N_19882);
and U22055 (N_22055,N_17953,N_17502);
nand U22056 (N_22056,N_18062,N_16341);
and U22057 (N_22057,N_18630,N_17634);
xnor U22058 (N_22058,N_18399,N_17628);
and U22059 (N_22059,N_19702,N_16834);
nor U22060 (N_22060,N_16235,N_18900);
xor U22061 (N_22061,N_15083,N_16935);
and U22062 (N_22062,N_16369,N_16992);
nor U22063 (N_22063,N_19002,N_19726);
nand U22064 (N_22064,N_19602,N_18133);
nand U22065 (N_22065,N_19676,N_17515);
or U22066 (N_22066,N_15079,N_15868);
nor U22067 (N_22067,N_16401,N_19231);
nor U22068 (N_22068,N_17536,N_19388);
and U22069 (N_22069,N_19932,N_15571);
and U22070 (N_22070,N_19225,N_19774);
xnor U22071 (N_22071,N_15800,N_18535);
or U22072 (N_22072,N_19162,N_16143);
xnor U22073 (N_22073,N_17812,N_19653);
nor U22074 (N_22074,N_19319,N_15518);
and U22075 (N_22075,N_16888,N_15463);
nor U22076 (N_22076,N_16933,N_16704);
or U22077 (N_22077,N_17239,N_18670);
nand U22078 (N_22078,N_19500,N_19408);
nand U22079 (N_22079,N_18458,N_16574);
or U22080 (N_22080,N_18999,N_19910);
nor U22081 (N_22081,N_19575,N_16720);
nor U22082 (N_22082,N_16417,N_18255);
nor U22083 (N_22083,N_18748,N_15429);
or U22084 (N_22084,N_19650,N_19477);
or U22085 (N_22085,N_15951,N_17924);
or U22086 (N_22086,N_19562,N_18059);
xor U22087 (N_22087,N_18848,N_17040);
or U22088 (N_22088,N_19591,N_17917);
or U22089 (N_22089,N_17940,N_18195);
nand U22090 (N_22090,N_19227,N_19307);
or U22091 (N_22091,N_16490,N_15257);
and U22092 (N_22092,N_17583,N_18853);
nor U22093 (N_22093,N_15444,N_18301);
or U22094 (N_22094,N_16896,N_15242);
xor U22095 (N_22095,N_17539,N_18590);
and U22096 (N_22096,N_16349,N_19345);
and U22097 (N_22097,N_18537,N_16968);
nor U22098 (N_22098,N_18279,N_17498);
or U22099 (N_22099,N_19878,N_19290);
and U22100 (N_22100,N_15718,N_19842);
nand U22101 (N_22101,N_17642,N_17429);
xnor U22102 (N_22102,N_19142,N_17382);
nor U22103 (N_22103,N_19723,N_18326);
and U22104 (N_22104,N_17990,N_17855);
nor U22105 (N_22105,N_16939,N_15584);
xor U22106 (N_22106,N_16174,N_17778);
xnor U22107 (N_22107,N_17126,N_15337);
nor U22108 (N_22108,N_17139,N_18462);
xor U22109 (N_22109,N_18254,N_16811);
nand U22110 (N_22110,N_16396,N_19239);
nor U22111 (N_22111,N_16040,N_18800);
nand U22112 (N_22112,N_19342,N_16831);
and U22113 (N_22113,N_18070,N_16177);
or U22114 (N_22114,N_16362,N_19743);
or U22115 (N_22115,N_17935,N_16569);
nor U22116 (N_22116,N_15938,N_15650);
nor U22117 (N_22117,N_15441,N_15117);
and U22118 (N_22118,N_16934,N_17686);
nor U22119 (N_22119,N_17054,N_16094);
nand U22120 (N_22120,N_17362,N_18678);
nor U22121 (N_22121,N_16371,N_17942);
nand U22122 (N_22122,N_18281,N_18128);
nor U22123 (N_22123,N_17571,N_18355);
or U22124 (N_22124,N_19133,N_16337);
and U22125 (N_22125,N_15329,N_17685);
or U22126 (N_22126,N_15882,N_19550);
or U22127 (N_22127,N_15906,N_19000);
xor U22128 (N_22128,N_19945,N_18322);
and U22129 (N_22129,N_17645,N_15638);
nand U22130 (N_22130,N_17246,N_17329);
xnor U22131 (N_22131,N_15953,N_19310);
and U22132 (N_22132,N_17043,N_16249);
or U22133 (N_22133,N_19860,N_19975);
xnor U22134 (N_22134,N_17176,N_17015);
xor U22135 (N_22135,N_19981,N_17752);
xor U22136 (N_22136,N_17534,N_16454);
or U22137 (N_22137,N_15494,N_16459);
or U22138 (N_22138,N_19959,N_15635);
and U22139 (N_22139,N_15023,N_15574);
nor U22140 (N_22140,N_17245,N_15012);
nor U22141 (N_22141,N_19044,N_18242);
nand U22142 (N_22142,N_18006,N_16815);
nand U22143 (N_22143,N_16254,N_17988);
nor U22144 (N_22144,N_19151,N_17205);
xnor U22145 (N_22145,N_17473,N_15476);
nor U22146 (N_22146,N_19457,N_16702);
or U22147 (N_22147,N_17044,N_19397);
and U22148 (N_22148,N_18224,N_16586);
or U22149 (N_22149,N_18849,N_15038);
nand U22150 (N_22150,N_19556,N_16606);
nor U22151 (N_22151,N_16825,N_15501);
nand U22152 (N_22152,N_16690,N_17532);
xnor U22153 (N_22153,N_19736,N_19933);
and U22154 (N_22154,N_17257,N_18642);
nor U22155 (N_22155,N_16003,N_17776);
or U22156 (N_22156,N_15461,N_15169);
nor U22157 (N_22157,N_17731,N_18484);
xnor U22158 (N_22158,N_17198,N_18017);
nor U22159 (N_22159,N_17501,N_16306);
and U22160 (N_22160,N_16405,N_18313);
xor U22161 (N_22161,N_16962,N_19504);
and U22162 (N_22162,N_18906,N_19920);
nand U22163 (N_22163,N_18887,N_19705);
or U22164 (N_22164,N_17025,N_17411);
nor U22165 (N_22165,N_17874,N_19849);
or U22166 (N_22166,N_19760,N_19124);
and U22167 (N_22167,N_15927,N_19442);
or U22168 (N_22168,N_17717,N_15512);
nand U22169 (N_22169,N_16451,N_19748);
or U22170 (N_22170,N_15062,N_19566);
nand U22171 (N_22171,N_15519,N_18196);
nand U22172 (N_22172,N_17519,N_19429);
and U22173 (N_22173,N_15388,N_19832);
or U22174 (N_22174,N_17788,N_18792);
and U22175 (N_22175,N_16069,N_19613);
and U22176 (N_22176,N_19523,N_17769);
nand U22177 (N_22177,N_18577,N_16207);
nor U22178 (N_22178,N_19097,N_17232);
nand U22179 (N_22179,N_16289,N_16075);
nand U22180 (N_22180,N_18362,N_17116);
or U22181 (N_22181,N_17550,N_17161);
nand U22182 (N_22182,N_19386,N_15556);
xor U22183 (N_22183,N_15219,N_15311);
or U22184 (N_22184,N_18779,N_17734);
nor U22185 (N_22185,N_15552,N_16709);
nand U22186 (N_22186,N_16724,N_19727);
nor U22187 (N_22187,N_17052,N_15448);
and U22188 (N_22188,N_19659,N_15656);
nand U22189 (N_22189,N_18043,N_17846);
or U22190 (N_22190,N_18987,N_15913);
nand U22191 (N_22191,N_18415,N_16178);
nand U22192 (N_22192,N_18223,N_19335);
or U22193 (N_22193,N_16503,N_17674);
nor U22194 (N_22194,N_15348,N_16570);
nand U22195 (N_22195,N_16551,N_17672);
nor U22196 (N_22196,N_17181,N_18511);
nor U22197 (N_22197,N_19641,N_16776);
nor U22198 (N_22198,N_16504,N_16827);
or U22199 (N_22199,N_19059,N_16437);
nor U22200 (N_22200,N_15793,N_19502);
or U22201 (N_22201,N_17098,N_16735);
or U22202 (N_22202,N_18184,N_17695);
or U22203 (N_22203,N_19003,N_16737);
or U22204 (N_22204,N_15321,N_19732);
and U22205 (N_22205,N_19695,N_15612);
or U22206 (N_22206,N_19047,N_17456);
and U22207 (N_22207,N_18645,N_17310);
or U22208 (N_22208,N_18929,N_15096);
and U22209 (N_22209,N_19589,N_15228);
and U22210 (N_22210,N_19285,N_16926);
nor U22211 (N_22211,N_18956,N_16923);
and U22212 (N_22212,N_18016,N_16344);
nand U22213 (N_22213,N_19415,N_19272);
xor U22214 (N_22214,N_19455,N_15138);
or U22215 (N_22215,N_15716,N_18416);
or U22216 (N_22216,N_16641,N_16723);
and U22217 (N_22217,N_19825,N_17675);
and U22218 (N_22218,N_19885,N_15150);
or U22219 (N_22219,N_15474,N_19977);
nand U22220 (N_22220,N_16681,N_15439);
and U22221 (N_22221,N_17679,N_15301);
and U22222 (N_22222,N_19174,N_17509);
and U22223 (N_22223,N_17437,N_16302);
xnor U22224 (N_22224,N_19370,N_19592);
nor U22225 (N_22225,N_17815,N_19313);
nand U22226 (N_22226,N_16433,N_18782);
and U22227 (N_22227,N_15154,N_19396);
nor U22228 (N_22228,N_19140,N_15551);
and U22229 (N_22229,N_18874,N_18619);
and U22230 (N_22230,N_15783,N_17751);
and U22231 (N_22231,N_19076,N_18048);
and U22232 (N_22232,N_18765,N_17862);
nor U22233 (N_22233,N_19838,N_16381);
and U22234 (N_22234,N_15397,N_17184);
nor U22235 (N_22235,N_15895,N_18327);
or U22236 (N_22236,N_17036,N_17330);
or U22237 (N_22237,N_19545,N_15788);
nand U22238 (N_22238,N_18463,N_19203);
xor U22239 (N_22239,N_16879,N_17458);
nand U22240 (N_22240,N_16854,N_19853);
and U22241 (N_22241,N_17412,N_15405);
and U22242 (N_22242,N_19127,N_18270);
xor U22243 (N_22243,N_17775,N_16692);
and U22244 (N_22244,N_16499,N_16963);
nand U22245 (N_22245,N_19738,N_19772);
or U22246 (N_22246,N_15703,N_17258);
and U22247 (N_22247,N_16107,N_18433);
or U22248 (N_22248,N_16321,N_15775);
xor U22249 (N_22249,N_18227,N_18351);
nor U22250 (N_22250,N_15603,N_19823);
nor U22251 (N_22251,N_19542,N_19694);
and U22252 (N_22252,N_18265,N_16418);
xnor U22253 (N_22253,N_15637,N_17885);
nand U22254 (N_22254,N_18702,N_18098);
nor U22255 (N_22255,N_16538,N_17284);
or U22256 (N_22256,N_15993,N_18250);
and U22257 (N_22257,N_16765,N_19510);
and U22258 (N_22258,N_16697,N_17655);
xnor U22259 (N_22259,N_19260,N_18257);
or U22260 (N_22260,N_17817,N_16579);
nor U22261 (N_22261,N_17069,N_19590);
or U22262 (N_22262,N_19563,N_16677);
and U22263 (N_22263,N_17948,N_16141);
and U22264 (N_22264,N_15019,N_19708);
nor U22265 (N_22265,N_15273,N_18699);
or U22266 (N_22266,N_17175,N_18764);
or U22267 (N_22267,N_18551,N_17326);
nor U22268 (N_22268,N_17880,N_19025);
nor U22269 (N_22269,N_19019,N_15453);
or U22270 (N_22270,N_15168,N_15309);
or U22271 (N_22271,N_17327,N_18082);
or U22272 (N_22272,N_16058,N_15781);
nor U22273 (N_22273,N_16785,N_16086);
or U22274 (N_22274,N_18990,N_16999);
or U22275 (N_22275,N_19579,N_17011);
nor U22276 (N_22276,N_15357,N_19302);
or U22277 (N_22277,N_17424,N_16487);
nand U22278 (N_22278,N_15663,N_17933);
nor U22279 (N_22279,N_17037,N_18109);
and U22280 (N_22280,N_16373,N_19049);
and U22281 (N_22281,N_16862,N_19634);
and U22282 (N_22282,N_18757,N_16138);
xor U22283 (N_22283,N_18150,N_16230);
nand U22284 (N_22284,N_19035,N_17378);
nand U22285 (N_22285,N_15440,N_16756);
nand U22286 (N_22286,N_18635,N_16412);
or U22287 (N_22287,N_17041,N_19793);
nor U22288 (N_22288,N_15505,N_19633);
and U22289 (N_22289,N_19389,N_18120);
nand U22290 (N_22290,N_15060,N_17079);
xor U22291 (N_22291,N_16577,N_18280);
nor U22292 (N_22292,N_16145,N_16056);
nor U22293 (N_22293,N_17562,N_17104);
or U22294 (N_22294,N_19795,N_17016);
nand U22295 (N_22295,N_16793,N_19801);
and U22296 (N_22296,N_19143,N_16650);
or U22297 (N_22297,N_17744,N_16482);
or U22298 (N_22298,N_15582,N_19083);
nand U22299 (N_22299,N_18739,N_18005);
or U22300 (N_22300,N_15581,N_18566);
or U22301 (N_22301,N_19356,N_17356);
and U22302 (N_22302,N_16590,N_17439);
and U22303 (N_22303,N_18831,N_16550);
nor U22304 (N_22304,N_16954,N_15174);
nand U22305 (N_22305,N_19093,N_15058);
nand U22306 (N_22306,N_19927,N_16591);
nand U22307 (N_22307,N_16047,N_15483);
xnor U22308 (N_22308,N_15877,N_17745);
or U22309 (N_22309,N_15875,N_15392);
nand U22310 (N_22310,N_17617,N_16796);
or U22311 (N_22311,N_16729,N_17870);
or U22312 (N_22312,N_18540,N_18226);
and U22313 (N_22313,N_17718,N_17854);
and U22314 (N_22314,N_18088,N_19139);
or U22315 (N_22315,N_15112,N_18794);
and U22316 (N_22316,N_15903,N_17859);
or U22317 (N_22317,N_19814,N_16491);
nand U22318 (N_22318,N_15209,N_15358);
and U22319 (N_22319,N_16089,N_17790);
nand U22320 (N_22320,N_19568,N_17787);
or U22321 (N_22321,N_15241,N_17577);
and U22322 (N_22322,N_18418,N_19364);
nand U22323 (N_22323,N_18325,N_18492);
or U22324 (N_22324,N_19022,N_15712);
nor U22325 (N_22325,N_17589,N_19237);
nor U22326 (N_22326,N_17361,N_15752);
nand U22327 (N_22327,N_17471,N_18052);
and U22328 (N_22328,N_16054,N_17199);
and U22329 (N_22329,N_19635,N_16869);
nand U22330 (N_22330,N_19757,N_16112);
nand U22331 (N_22331,N_18908,N_18768);
or U22332 (N_22332,N_19371,N_15946);
xnor U22333 (N_22333,N_17230,N_16016);
nand U22334 (N_22334,N_17749,N_17114);
or U22335 (N_22335,N_16170,N_19393);
or U22336 (N_22336,N_17112,N_15921);
or U22337 (N_22337,N_17129,N_16657);
nor U22338 (N_22338,N_16922,N_17958);
and U22339 (N_22339,N_17027,N_19928);
or U22340 (N_22340,N_18873,N_15705);
or U22341 (N_22341,N_19924,N_18648);
nand U22342 (N_22342,N_17359,N_16947);
nor U22343 (N_22343,N_19274,N_19350);
and U22344 (N_22344,N_18490,N_18689);
nand U22345 (N_22345,N_16250,N_19638);
xnor U22346 (N_22346,N_19077,N_16053);
or U22347 (N_22347,N_19712,N_16328);
or U22348 (N_22348,N_15208,N_18559);
nand U22349 (N_22349,N_15655,N_16245);
nor U22350 (N_22350,N_18031,N_17148);
and U22351 (N_22351,N_18519,N_18135);
xnor U22352 (N_22352,N_16596,N_19540);
or U22353 (N_22353,N_19737,N_15189);
and U22354 (N_22354,N_19898,N_15400);
or U22355 (N_22355,N_17646,N_16874);
nor U22356 (N_22356,N_17720,N_17264);
nor U22357 (N_22357,N_18737,N_16711);
nor U22358 (N_22358,N_16042,N_17779);
nor U22359 (N_22359,N_19799,N_18380);
xor U22360 (N_22360,N_16792,N_17280);
nor U22361 (N_22361,N_17670,N_19123);
and U22362 (N_22362,N_17525,N_17055);
nand U22363 (N_22363,N_19554,N_15816);
and U22364 (N_22364,N_19329,N_16683);
or U22365 (N_22365,N_16531,N_15759);
xor U22366 (N_22366,N_17164,N_15170);
nand U22367 (N_22367,N_17962,N_15561);
xor U22368 (N_22368,N_16243,N_15378);
nand U22369 (N_22369,N_17837,N_19232);
and U22370 (N_22370,N_19992,N_19522);
and U22371 (N_22371,N_15553,N_15804);
nand U22372 (N_22372,N_16377,N_16911);
nor U22373 (N_22373,N_19791,N_15782);
and U22374 (N_22374,N_15207,N_18243);
nand U22375 (N_22375,N_18451,N_18682);
and U22376 (N_22376,N_18099,N_15562);
nand U22377 (N_22377,N_15888,N_19057);
nand U22378 (N_22378,N_17881,N_18086);
or U22379 (N_22379,N_18104,N_19905);
and U22380 (N_22380,N_15805,N_18693);
nand U22381 (N_22381,N_16296,N_15680);
xor U22382 (N_22382,N_18718,N_18402);
and U22383 (N_22383,N_15701,N_15157);
nand U22384 (N_22384,N_19512,N_15983);
or U22385 (N_22385,N_15959,N_18753);
or U22386 (N_22386,N_16224,N_16794);
nand U22387 (N_22387,N_17764,N_18000);
xnor U22388 (N_22388,N_19844,N_19505);
nor U22389 (N_22389,N_19514,N_16908);
and U22390 (N_22390,N_16155,N_19398);
nand U22391 (N_22391,N_17991,N_16925);
xor U22392 (N_22392,N_19071,N_15566);
nor U22393 (N_22393,N_17774,N_16204);
nand U22394 (N_22394,N_15398,N_16839);
nor U22395 (N_22395,N_15784,N_15020);
or U22396 (N_22396,N_19091,N_17296);
xor U22397 (N_22397,N_16544,N_16419);
nand U22398 (N_22398,N_17579,N_18656);
or U22399 (N_22399,N_18840,N_19160);
nor U22400 (N_22400,N_19054,N_16977);
nand U22401 (N_22401,N_16718,N_19412);
and U22402 (N_22402,N_17026,N_15909);
and U22403 (N_22403,N_15280,N_15569);
xnor U22404 (N_22404,N_15692,N_15846);
and U22405 (N_22405,N_15778,N_15433);
and U22406 (N_22406,N_17875,N_17417);
or U22407 (N_22407,N_15652,N_18424);
xor U22408 (N_22408,N_19042,N_15317);
or U22409 (N_22409,N_15394,N_17585);
or U22410 (N_22410,N_16900,N_17407);
xor U22411 (N_22411,N_16899,N_15563);
and U22412 (N_22412,N_18815,N_19578);
or U22413 (N_22413,N_15464,N_18661);
and U22414 (N_22414,N_17997,N_17543);
and U22415 (N_22415,N_15851,N_18364);
and U22416 (N_22416,N_15724,N_18777);
nor U22417 (N_22417,N_19915,N_19090);
nor U22418 (N_22418,N_16519,N_17404);
nor U22419 (N_22419,N_16868,N_19619);
nand U22420 (N_22420,N_16757,N_18649);
or U22421 (N_22421,N_19092,N_18662);
and U22422 (N_22422,N_15114,N_18690);
and U22423 (N_22423,N_18716,N_16866);
nand U22424 (N_22424,N_17728,N_18515);
nand U22425 (N_22425,N_16987,N_18623);
and U22426 (N_22426,N_19906,N_19763);
xor U22427 (N_22427,N_19887,N_17565);
nand U22428 (N_22428,N_15713,N_18454);
or U22429 (N_22429,N_16914,N_18182);
nand U22430 (N_22430,N_19115,N_16209);
or U22431 (N_22431,N_15234,N_18677);
nand U22432 (N_22432,N_16464,N_15947);
nor U22433 (N_22433,N_15446,N_19230);
nor U22434 (N_22434,N_18508,N_18530);
nor U22435 (N_22435,N_17639,N_18883);
and U22436 (N_22436,N_19149,N_18249);
nand U22437 (N_22437,N_15952,N_18155);
nor U22438 (N_22438,N_15281,N_16495);
xor U22439 (N_22439,N_19974,N_19155);
xor U22440 (N_22440,N_19102,N_16500);
or U22441 (N_22441,N_15387,N_19073);
or U22442 (N_22442,N_18857,N_18934);
nor U22443 (N_22443,N_15055,N_19304);
and U22444 (N_22444,N_16743,N_16468);
and U22445 (N_22445,N_19234,N_17581);
and U22446 (N_22446,N_16233,N_16901);
and U22447 (N_22447,N_19831,N_15347);
and U22448 (N_22448,N_18337,N_16476);
and U22449 (N_22449,N_15176,N_17077);
and U22450 (N_22450,N_17231,N_18877);
nand U22451 (N_22451,N_15665,N_16148);
nor U22452 (N_22452,N_19318,N_16423);
xor U22453 (N_22453,N_16029,N_16967);
nand U22454 (N_22454,N_16917,N_17265);
nand U22455 (N_22455,N_16738,N_18880);
nor U22456 (N_22456,N_19570,N_16327);
nor U22457 (N_22457,N_18245,N_18287);
and U22458 (N_22458,N_19377,N_18145);
nand U22459 (N_22459,N_19251,N_17496);
nand U22460 (N_22460,N_17708,N_18122);
or U22461 (N_22461,N_19884,N_18235);
or U22462 (N_22462,N_16166,N_15944);
and U22463 (N_22463,N_15367,N_18406);
nand U22464 (N_22464,N_15765,N_16974);
nor U22465 (N_22465,N_16789,N_17594);
nor U22466 (N_22466,N_17780,N_17486);
nand U22467 (N_22467,N_15187,N_17331);
xnor U22468 (N_22468,N_16256,N_16474);
and U22469 (N_22469,N_16864,N_16713);
nor U22470 (N_22470,N_18663,N_15645);
xor U22471 (N_22471,N_15006,N_16830);
nor U22472 (N_22472,N_16301,N_15408);
nor U22473 (N_22473,N_19186,N_18529);
and U22474 (N_22474,N_19249,N_19211);
xor U22475 (N_22475,N_16820,N_19275);
nand U22476 (N_22476,N_18376,N_15514);
or U22477 (N_22477,N_15714,N_18395);
and U22478 (N_22478,N_15997,N_17572);
or U22479 (N_22479,N_16077,N_16314);
nor U22480 (N_22480,N_19917,N_16747);
nor U22481 (N_22481,N_17182,N_17819);
and U22482 (N_22482,N_19600,N_16136);
nor U22483 (N_22483,N_15010,N_16534);
nand U22484 (N_22484,N_17122,N_18010);
nor U22485 (N_22485,N_17850,N_19421);
nor U22486 (N_22486,N_17574,N_15539);
and U22487 (N_22487,N_17705,N_16061);
nor U22488 (N_22488,N_17482,N_18238);
nor U22489 (N_22489,N_19287,N_18936);
or U22490 (N_22490,N_15327,N_16222);
and U22491 (N_22491,N_18866,N_16385);
or U22492 (N_22492,N_18205,N_17289);
or U22493 (N_22493,N_15296,N_18611);
nand U22494 (N_22494,N_19305,N_16670);
nor U22495 (N_22495,N_19912,N_15354);
and U22496 (N_22496,N_15786,N_16777);
or U22497 (N_22497,N_17099,N_15919);
nor U22498 (N_22498,N_16326,N_17737);
nand U22499 (N_22499,N_17224,N_18797);
or U22500 (N_22500,N_18150,N_16958);
and U22501 (N_22501,N_18029,N_19407);
nor U22502 (N_22502,N_18589,N_19726);
and U22503 (N_22503,N_16428,N_18343);
or U22504 (N_22504,N_15237,N_16171);
and U22505 (N_22505,N_19983,N_19212);
and U22506 (N_22506,N_16251,N_19024);
or U22507 (N_22507,N_18805,N_17676);
nand U22508 (N_22508,N_19227,N_19555);
nor U22509 (N_22509,N_16070,N_17430);
nor U22510 (N_22510,N_18711,N_17812);
and U22511 (N_22511,N_15708,N_17503);
nand U22512 (N_22512,N_18088,N_15752);
nand U22513 (N_22513,N_17672,N_16650);
and U22514 (N_22514,N_18049,N_16440);
nand U22515 (N_22515,N_18910,N_17364);
xnor U22516 (N_22516,N_18542,N_18804);
nand U22517 (N_22517,N_15606,N_15385);
or U22518 (N_22518,N_15816,N_18401);
or U22519 (N_22519,N_17042,N_18526);
nor U22520 (N_22520,N_16785,N_18478);
or U22521 (N_22521,N_17988,N_19131);
and U22522 (N_22522,N_17430,N_19682);
or U22523 (N_22523,N_19924,N_19888);
nand U22524 (N_22524,N_18180,N_16733);
nor U22525 (N_22525,N_15784,N_16567);
xnor U22526 (N_22526,N_15361,N_18358);
nor U22527 (N_22527,N_17050,N_16401);
nand U22528 (N_22528,N_17791,N_17426);
nor U22529 (N_22529,N_18259,N_19518);
or U22530 (N_22530,N_18589,N_17279);
nand U22531 (N_22531,N_19059,N_19553);
or U22532 (N_22532,N_17794,N_18961);
nand U22533 (N_22533,N_18356,N_17754);
or U22534 (N_22534,N_16016,N_15637);
nand U22535 (N_22535,N_15722,N_16221);
nand U22536 (N_22536,N_15949,N_15422);
nand U22537 (N_22537,N_18847,N_17980);
or U22538 (N_22538,N_17784,N_17162);
nand U22539 (N_22539,N_16294,N_15402);
or U22540 (N_22540,N_19482,N_17316);
nor U22541 (N_22541,N_18189,N_17221);
xnor U22542 (N_22542,N_17723,N_19270);
xnor U22543 (N_22543,N_17712,N_16937);
nor U22544 (N_22544,N_16195,N_16998);
or U22545 (N_22545,N_15943,N_19150);
and U22546 (N_22546,N_18549,N_15568);
and U22547 (N_22547,N_17747,N_19681);
nor U22548 (N_22548,N_17104,N_17419);
or U22549 (N_22549,N_19281,N_18911);
and U22550 (N_22550,N_17873,N_19083);
nor U22551 (N_22551,N_17470,N_16616);
nor U22552 (N_22552,N_17038,N_19830);
or U22553 (N_22553,N_15250,N_17275);
or U22554 (N_22554,N_18679,N_19539);
nand U22555 (N_22555,N_18990,N_16229);
nand U22556 (N_22556,N_18879,N_18000);
nor U22557 (N_22557,N_18093,N_18187);
or U22558 (N_22558,N_18417,N_15954);
nor U22559 (N_22559,N_16720,N_18834);
or U22560 (N_22560,N_19174,N_15602);
and U22561 (N_22561,N_16969,N_15899);
and U22562 (N_22562,N_16319,N_17030);
nor U22563 (N_22563,N_16241,N_17031);
nand U22564 (N_22564,N_17712,N_16044);
xnor U22565 (N_22565,N_19503,N_19237);
nand U22566 (N_22566,N_18323,N_18310);
nand U22567 (N_22567,N_18810,N_18600);
nand U22568 (N_22568,N_16940,N_17367);
nor U22569 (N_22569,N_16989,N_15091);
nand U22570 (N_22570,N_18522,N_16607);
and U22571 (N_22571,N_16098,N_18659);
nor U22572 (N_22572,N_16631,N_17207);
and U22573 (N_22573,N_18554,N_16942);
or U22574 (N_22574,N_15654,N_16922);
nand U22575 (N_22575,N_18187,N_19335);
or U22576 (N_22576,N_19895,N_19408);
xnor U22577 (N_22577,N_15016,N_18105);
and U22578 (N_22578,N_15749,N_19240);
xor U22579 (N_22579,N_18092,N_16157);
nor U22580 (N_22580,N_19867,N_19495);
nand U22581 (N_22581,N_19858,N_18378);
and U22582 (N_22582,N_18265,N_19677);
or U22583 (N_22583,N_17492,N_16168);
or U22584 (N_22584,N_16156,N_17960);
or U22585 (N_22585,N_18961,N_15601);
xnor U22586 (N_22586,N_16934,N_18542);
and U22587 (N_22587,N_17340,N_17783);
and U22588 (N_22588,N_16176,N_15645);
or U22589 (N_22589,N_19370,N_15198);
nor U22590 (N_22590,N_17444,N_15290);
nand U22591 (N_22591,N_17656,N_16705);
nand U22592 (N_22592,N_16693,N_17964);
nor U22593 (N_22593,N_19056,N_19042);
nor U22594 (N_22594,N_15156,N_18808);
or U22595 (N_22595,N_15108,N_18966);
or U22596 (N_22596,N_18441,N_17790);
nand U22597 (N_22597,N_16656,N_17217);
nor U22598 (N_22598,N_17453,N_17744);
nand U22599 (N_22599,N_19941,N_16445);
nor U22600 (N_22600,N_15486,N_18203);
nor U22601 (N_22601,N_19274,N_15122);
or U22602 (N_22602,N_17822,N_18620);
nand U22603 (N_22603,N_17762,N_16103);
nand U22604 (N_22604,N_19844,N_18177);
nand U22605 (N_22605,N_18102,N_18822);
or U22606 (N_22606,N_18530,N_15199);
and U22607 (N_22607,N_17111,N_15663);
and U22608 (N_22608,N_19398,N_19716);
and U22609 (N_22609,N_16801,N_16511);
and U22610 (N_22610,N_15157,N_16110);
or U22611 (N_22611,N_15342,N_16368);
or U22612 (N_22612,N_16198,N_19633);
or U22613 (N_22613,N_15695,N_16339);
nand U22614 (N_22614,N_18117,N_15418);
nor U22615 (N_22615,N_19016,N_15178);
nor U22616 (N_22616,N_18387,N_15445);
nand U22617 (N_22617,N_16059,N_16046);
nand U22618 (N_22618,N_17872,N_15140);
nor U22619 (N_22619,N_15938,N_17008);
nand U22620 (N_22620,N_15194,N_17411);
nor U22621 (N_22621,N_16087,N_17843);
nor U22622 (N_22622,N_19589,N_16883);
nor U22623 (N_22623,N_15719,N_16883);
nand U22624 (N_22624,N_15510,N_15275);
or U22625 (N_22625,N_19774,N_15067);
nor U22626 (N_22626,N_17352,N_19299);
nor U22627 (N_22627,N_18573,N_19080);
and U22628 (N_22628,N_17375,N_18863);
and U22629 (N_22629,N_17080,N_19988);
nand U22630 (N_22630,N_18199,N_19422);
nand U22631 (N_22631,N_16052,N_18775);
xor U22632 (N_22632,N_17532,N_15972);
nand U22633 (N_22633,N_18130,N_18525);
nor U22634 (N_22634,N_19359,N_16119);
or U22635 (N_22635,N_16139,N_17867);
nand U22636 (N_22636,N_16914,N_17786);
or U22637 (N_22637,N_16728,N_19395);
and U22638 (N_22638,N_17383,N_18269);
and U22639 (N_22639,N_16804,N_15746);
or U22640 (N_22640,N_18304,N_16142);
or U22641 (N_22641,N_18464,N_15981);
or U22642 (N_22642,N_18151,N_15392);
xnor U22643 (N_22643,N_18592,N_19045);
nand U22644 (N_22644,N_15343,N_15536);
nand U22645 (N_22645,N_15525,N_15297);
nand U22646 (N_22646,N_16909,N_17372);
and U22647 (N_22647,N_19325,N_18559);
nor U22648 (N_22648,N_16107,N_19915);
and U22649 (N_22649,N_19279,N_16305);
and U22650 (N_22650,N_17792,N_15862);
nand U22651 (N_22651,N_15721,N_18533);
or U22652 (N_22652,N_19225,N_19476);
or U22653 (N_22653,N_17159,N_18417);
or U22654 (N_22654,N_19504,N_15564);
or U22655 (N_22655,N_18905,N_18616);
and U22656 (N_22656,N_19420,N_16626);
nor U22657 (N_22657,N_18093,N_18520);
xnor U22658 (N_22658,N_17111,N_19529);
or U22659 (N_22659,N_15972,N_18148);
and U22660 (N_22660,N_16506,N_19014);
and U22661 (N_22661,N_17611,N_17125);
or U22662 (N_22662,N_16806,N_16372);
nor U22663 (N_22663,N_15730,N_17490);
nor U22664 (N_22664,N_15840,N_17845);
or U22665 (N_22665,N_15589,N_16687);
nor U22666 (N_22666,N_17938,N_17742);
nor U22667 (N_22667,N_15543,N_17580);
and U22668 (N_22668,N_17683,N_17668);
nor U22669 (N_22669,N_18451,N_16630);
nand U22670 (N_22670,N_17214,N_15545);
nand U22671 (N_22671,N_16283,N_19798);
and U22672 (N_22672,N_17901,N_18203);
nand U22673 (N_22673,N_18047,N_17193);
and U22674 (N_22674,N_17394,N_16324);
or U22675 (N_22675,N_18925,N_15105);
or U22676 (N_22676,N_19034,N_19965);
nor U22677 (N_22677,N_15592,N_18005);
xnor U22678 (N_22678,N_18984,N_18737);
and U22679 (N_22679,N_15082,N_17159);
and U22680 (N_22680,N_17988,N_16240);
and U22681 (N_22681,N_17126,N_16076);
nand U22682 (N_22682,N_15821,N_15465);
or U22683 (N_22683,N_18512,N_18918);
nor U22684 (N_22684,N_18837,N_16659);
nand U22685 (N_22685,N_18936,N_16421);
and U22686 (N_22686,N_16959,N_18779);
or U22687 (N_22687,N_19573,N_16826);
or U22688 (N_22688,N_18880,N_18512);
or U22689 (N_22689,N_17924,N_17913);
or U22690 (N_22690,N_19601,N_18395);
and U22691 (N_22691,N_17908,N_17164);
or U22692 (N_22692,N_19054,N_17269);
nor U22693 (N_22693,N_18026,N_16227);
nand U22694 (N_22694,N_19711,N_15399);
or U22695 (N_22695,N_18146,N_17669);
and U22696 (N_22696,N_19613,N_16772);
or U22697 (N_22697,N_15192,N_16712);
nand U22698 (N_22698,N_19232,N_17508);
and U22699 (N_22699,N_16821,N_18777);
and U22700 (N_22700,N_15377,N_18335);
and U22701 (N_22701,N_19905,N_16728);
nand U22702 (N_22702,N_19580,N_18386);
or U22703 (N_22703,N_16765,N_19221);
nor U22704 (N_22704,N_18423,N_16969);
or U22705 (N_22705,N_17044,N_19682);
and U22706 (N_22706,N_16185,N_17782);
xnor U22707 (N_22707,N_17016,N_17969);
nor U22708 (N_22708,N_19959,N_18588);
nand U22709 (N_22709,N_16836,N_19569);
and U22710 (N_22710,N_17306,N_15594);
nand U22711 (N_22711,N_18731,N_16166);
nor U22712 (N_22712,N_17557,N_17606);
or U22713 (N_22713,N_16630,N_16552);
and U22714 (N_22714,N_19027,N_18242);
and U22715 (N_22715,N_16760,N_15092);
or U22716 (N_22716,N_17911,N_16088);
and U22717 (N_22717,N_15498,N_16535);
and U22718 (N_22718,N_15904,N_19128);
nand U22719 (N_22719,N_18073,N_18364);
nor U22720 (N_22720,N_18995,N_18112);
nor U22721 (N_22721,N_16503,N_15070);
nor U22722 (N_22722,N_15445,N_16966);
nor U22723 (N_22723,N_18132,N_19069);
nor U22724 (N_22724,N_19622,N_19823);
or U22725 (N_22725,N_19489,N_17650);
and U22726 (N_22726,N_17725,N_15761);
and U22727 (N_22727,N_15590,N_15077);
or U22728 (N_22728,N_19676,N_16883);
or U22729 (N_22729,N_18868,N_18707);
and U22730 (N_22730,N_16465,N_19177);
and U22731 (N_22731,N_17226,N_15699);
and U22732 (N_22732,N_19222,N_18988);
or U22733 (N_22733,N_17077,N_16955);
xnor U22734 (N_22734,N_15493,N_16623);
and U22735 (N_22735,N_19189,N_19529);
and U22736 (N_22736,N_17440,N_18158);
xor U22737 (N_22737,N_18192,N_18743);
or U22738 (N_22738,N_18672,N_17617);
nand U22739 (N_22739,N_19211,N_18817);
nand U22740 (N_22740,N_15523,N_19603);
or U22741 (N_22741,N_18988,N_19392);
nor U22742 (N_22742,N_18705,N_16090);
or U22743 (N_22743,N_19456,N_18449);
nor U22744 (N_22744,N_18421,N_18691);
nor U22745 (N_22745,N_17395,N_19415);
nand U22746 (N_22746,N_15067,N_15372);
or U22747 (N_22747,N_19545,N_19829);
nor U22748 (N_22748,N_17728,N_18374);
nor U22749 (N_22749,N_17755,N_19076);
and U22750 (N_22750,N_16334,N_19194);
or U22751 (N_22751,N_19434,N_19904);
xnor U22752 (N_22752,N_15475,N_15946);
nor U22753 (N_22753,N_15886,N_16052);
nor U22754 (N_22754,N_18355,N_17508);
nor U22755 (N_22755,N_15382,N_18991);
or U22756 (N_22756,N_19146,N_18949);
nand U22757 (N_22757,N_19910,N_15721);
nor U22758 (N_22758,N_18204,N_19119);
nand U22759 (N_22759,N_19409,N_18126);
and U22760 (N_22760,N_19356,N_15319);
or U22761 (N_22761,N_15620,N_15141);
nand U22762 (N_22762,N_17949,N_19354);
and U22763 (N_22763,N_18273,N_19510);
or U22764 (N_22764,N_15483,N_15534);
and U22765 (N_22765,N_18792,N_19391);
or U22766 (N_22766,N_15690,N_19462);
and U22767 (N_22767,N_16482,N_19266);
xor U22768 (N_22768,N_17712,N_17526);
nand U22769 (N_22769,N_15002,N_17969);
nand U22770 (N_22770,N_17000,N_19650);
nor U22771 (N_22771,N_19407,N_19576);
nand U22772 (N_22772,N_15400,N_17139);
and U22773 (N_22773,N_18800,N_17865);
nand U22774 (N_22774,N_19751,N_18217);
or U22775 (N_22775,N_19563,N_18409);
or U22776 (N_22776,N_17652,N_17318);
nand U22777 (N_22777,N_17842,N_18336);
or U22778 (N_22778,N_19361,N_19051);
nor U22779 (N_22779,N_17068,N_16236);
nand U22780 (N_22780,N_17587,N_18182);
nand U22781 (N_22781,N_19350,N_19277);
nor U22782 (N_22782,N_19873,N_17559);
and U22783 (N_22783,N_17821,N_15695);
and U22784 (N_22784,N_15746,N_17756);
and U22785 (N_22785,N_19509,N_15955);
nor U22786 (N_22786,N_19872,N_16388);
or U22787 (N_22787,N_15149,N_19652);
or U22788 (N_22788,N_19159,N_19500);
xor U22789 (N_22789,N_16164,N_15746);
or U22790 (N_22790,N_16879,N_17244);
and U22791 (N_22791,N_17847,N_19636);
and U22792 (N_22792,N_19957,N_18885);
or U22793 (N_22793,N_19905,N_19254);
or U22794 (N_22794,N_15164,N_16619);
nor U22795 (N_22795,N_17683,N_19185);
and U22796 (N_22796,N_17081,N_18005);
or U22797 (N_22797,N_18612,N_15696);
or U22798 (N_22798,N_18913,N_19455);
or U22799 (N_22799,N_19678,N_18848);
nand U22800 (N_22800,N_18384,N_17146);
nand U22801 (N_22801,N_16289,N_19501);
xor U22802 (N_22802,N_16806,N_19198);
nor U22803 (N_22803,N_17017,N_18920);
nand U22804 (N_22804,N_15976,N_17984);
nand U22805 (N_22805,N_15914,N_16087);
or U22806 (N_22806,N_19853,N_15929);
nor U22807 (N_22807,N_19552,N_15534);
nand U22808 (N_22808,N_15442,N_15894);
nand U22809 (N_22809,N_16540,N_18322);
and U22810 (N_22810,N_15022,N_17239);
or U22811 (N_22811,N_19532,N_19602);
or U22812 (N_22812,N_18113,N_15665);
nand U22813 (N_22813,N_16994,N_16153);
nand U22814 (N_22814,N_15880,N_17650);
nand U22815 (N_22815,N_15153,N_16798);
nand U22816 (N_22816,N_16477,N_18253);
xnor U22817 (N_22817,N_15129,N_15048);
nand U22818 (N_22818,N_19275,N_18946);
and U22819 (N_22819,N_18954,N_19405);
nor U22820 (N_22820,N_19549,N_16937);
or U22821 (N_22821,N_17881,N_18527);
nand U22822 (N_22822,N_17626,N_18823);
and U22823 (N_22823,N_16437,N_17442);
and U22824 (N_22824,N_17517,N_17776);
xnor U22825 (N_22825,N_16644,N_15661);
nand U22826 (N_22826,N_19003,N_16986);
and U22827 (N_22827,N_15521,N_18081);
nor U22828 (N_22828,N_15102,N_15728);
nor U22829 (N_22829,N_16189,N_16657);
or U22830 (N_22830,N_17903,N_19580);
nor U22831 (N_22831,N_16979,N_16915);
nor U22832 (N_22832,N_15327,N_16688);
or U22833 (N_22833,N_15006,N_17118);
nand U22834 (N_22834,N_18263,N_17914);
and U22835 (N_22835,N_19425,N_16645);
and U22836 (N_22836,N_19870,N_16724);
and U22837 (N_22837,N_15077,N_16890);
nand U22838 (N_22838,N_18760,N_15199);
or U22839 (N_22839,N_16058,N_18034);
or U22840 (N_22840,N_17004,N_17782);
nor U22841 (N_22841,N_17984,N_19576);
or U22842 (N_22842,N_19534,N_18952);
nor U22843 (N_22843,N_15760,N_19641);
nor U22844 (N_22844,N_19119,N_17916);
or U22845 (N_22845,N_16080,N_16450);
nor U22846 (N_22846,N_16812,N_19568);
nand U22847 (N_22847,N_17692,N_15512);
or U22848 (N_22848,N_15592,N_18334);
nand U22849 (N_22849,N_15177,N_18306);
and U22850 (N_22850,N_17448,N_15951);
and U22851 (N_22851,N_17631,N_18818);
nand U22852 (N_22852,N_17182,N_19629);
xnor U22853 (N_22853,N_15604,N_15866);
xnor U22854 (N_22854,N_19037,N_19764);
or U22855 (N_22855,N_15617,N_15285);
and U22856 (N_22856,N_17569,N_19314);
nand U22857 (N_22857,N_18946,N_17350);
nand U22858 (N_22858,N_17096,N_19621);
and U22859 (N_22859,N_16645,N_15160);
xnor U22860 (N_22860,N_17542,N_19584);
nand U22861 (N_22861,N_17103,N_17005);
or U22862 (N_22862,N_17022,N_19907);
and U22863 (N_22863,N_17269,N_18022);
and U22864 (N_22864,N_19035,N_15659);
xor U22865 (N_22865,N_19163,N_15867);
and U22866 (N_22866,N_16842,N_16328);
or U22867 (N_22867,N_17968,N_18309);
nand U22868 (N_22868,N_15313,N_18010);
nor U22869 (N_22869,N_16772,N_17594);
and U22870 (N_22870,N_18153,N_16393);
nor U22871 (N_22871,N_17831,N_18190);
nor U22872 (N_22872,N_15416,N_17216);
or U22873 (N_22873,N_17418,N_16710);
nor U22874 (N_22874,N_18274,N_18390);
xor U22875 (N_22875,N_18243,N_19708);
xor U22876 (N_22876,N_19501,N_17157);
or U22877 (N_22877,N_18173,N_16486);
and U22878 (N_22878,N_15251,N_15546);
nand U22879 (N_22879,N_19709,N_16522);
or U22880 (N_22880,N_15327,N_18122);
nand U22881 (N_22881,N_18462,N_18901);
nand U22882 (N_22882,N_19528,N_17074);
nand U22883 (N_22883,N_17071,N_19067);
nor U22884 (N_22884,N_19925,N_16384);
or U22885 (N_22885,N_15036,N_16389);
or U22886 (N_22886,N_19424,N_16358);
xnor U22887 (N_22887,N_15729,N_15096);
xnor U22888 (N_22888,N_18156,N_16398);
or U22889 (N_22889,N_16260,N_18481);
and U22890 (N_22890,N_16826,N_15754);
nor U22891 (N_22891,N_16564,N_18060);
nor U22892 (N_22892,N_16212,N_15855);
xor U22893 (N_22893,N_17258,N_18792);
or U22894 (N_22894,N_18031,N_16000);
nor U22895 (N_22895,N_17196,N_17148);
nand U22896 (N_22896,N_18521,N_16405);
and U22897 (N_22897,N_15651,N_18327);
and U22898 (N_22898,N_17219,N_16308);
nand U22899 (N_22899,N_19437,N_19553);
nand U22900 (N_22900,N_18354,N_18269);
or U22901 (N_22901,N_17709,N_19507);
or U22902 (N_22902,N_17763,N_18811);
nor U22903 (N_22903,N_15008,N_17580);
nand U22904 (N_22904,N_15489,N_16558);
or U22905 (N_22905,N_19477,N_15166);
or U22906 (N_22906,N_17403,N_15894);
and U22907 (N_22907,N_16373,N_15046);
nand U22908 (N_22908,N_15681,N_18382);
nand U22909 (N_22909,N_15338,N_18398);
or U22910 (N_22910,N_18390,N_19115);
and U22911 (N_22911,N_17357,N_15578);
nand U22912 (N_22912,N_18382,N_19875);
and U22913 (N_22913,N_19577,N_18859);
nand U22914 (N_22914,N_19414,N_17432);
nor U22915 (N_22915,N_18465,N_15119);
nor U22916 (N_22916,N_18084,N_17834);
and U22917 (N_22917,N_15509,N_18672);
and U22918 (N_22918,N_15297,N_17935);
xnor U22919 (N_22919,N_18459,N_18139);
nor U22920 (N_22920,N_18330,N_19278);
nor U22921 (N_22921,N_16520,N_15251);
nor U22922 (N_22922,N_17824,N_19526);
or U22923 (N_22923,N_18399,N_16234);
nand U22924 (N_22924,N_16746,N_16901);
or U22925 (N_22925,N_16550,N_18704);
nor U22926 (N_22926,N_19277,N_17243);
or U22927 (N_22927,N_15479,N_18510);
nor U22928 (N_22928,N_18339,N_19480);
nor U22929 (N_22929,N_16693,N_17831);
nor U22930 (N_22930,N_16757,N_16928);
nor U22931 (N_22931,N_19721,N_15845);
nand U22932 (N_22932,N_17315,N_17238);
and U22933 (N_22933,N_15895,N_16457);
and U22934 (N_22934,N_17857,N_19740);
or U22935 (N_22935,N_15602,N_15133);
xnor U22936 (N_22936,N_16263,N_18912);
and U22937 (N_22937,N_17880,N_19885);
xnor U22938 (N_22938,N_16807,N_15455);
nor U22939 (N_22939,N_15115,N_18363);
nor U22940 (N_22940,N_16927,N_16560);
or U22941 (N_22941,N_17171,N_17713);
nor U22942 (N_22942,N_15407,N_15776);
nor U22943 (N_22943,N_17996,N_17042);
or U22944 (N_22944,N_15477,N_18588);
nand U22945 (N_22945,N_17383,N_19444);
nand U22946 (N_22946,N_16933,N_15890);
nor U22947 (N_22947,N_17825,N_16207);
nand U22948 (N_22948,N_18066,N_19253);
nand U22949 (N_22949,N_19045,N_16088);
xor U22950 (N_22950,N_18935,N_17321);
nor U22951 (N_22951,N_18489,N_19749);
nor U22952 (N_22952,N_17666,N_18295);
or U22953 (N_22953,N_18422,N_17601);
nand U22954 (N_22954,N_15025,N_18350);
or U22955 (N_22955,N_18708,N_18177);
nor U22956 (N_22956,N_16001,N_19300);
or U22957 (N_22957,N_19990,N_15139);
nor U22958 (N_22958,N_19821,N_18527);
nor U22959 (N_22959,N_15177,N_16488);
or U22960 (N_22960,N_15807,N_18150);
and U22961 (N_22961,N_18954,N_17300);
nor U22962 (N_22962,N_17257,N_15275);
and U22963 (N_22963,N_18892,N_16663);
nand U22964 (N_22964,N_18015,N_19453);
or U22965 (N_22965,N_18689,N_17348);
nor U22966 (N_22966,N_18263,N_18840);
xor U22967 (N_22967,N_16499,N_16918);
xor U22968 (N_22968,N_16473,N_16998);
or U22969 (N_22969,N_16244,N_19578);
xor U22970 (N_22970,N_18378,N_17688);
or U22971 (N_22971,N_18771,N_17396);
or U22972 (N_22972,N_18618,N_15384);
nand U22973 (N_22973,N_16312,N_18758);
and U22974 (N_22974,N_18349,N_16548);
nand U22975 (N_22975,N_17383,N_16255);
nor U22976 (N_22976,N_16052,N_15638);
nand U22977 (N_22977,N_15699,N_18248);
nand U22978 (N_22978,N_15070,N_15944);
or U22979 (N_22979,N_19745,N_16687);
nand U22980 (N_22980,N_16619,N_16854);
nand U22981 (N_22981,N_15173,N_17956);
or U22982 (N_22982,N_17238,N_16285);
or U22983 (N_22983,N_15288,N_17781);
or U22984 (N_22984,N_18400,N_15870);
or U22985 (N_22985,N_19003,N_17668);
and U22986 (N_22986,N_15560,N_18940);
xor U22987 (N_22987,N_18032,N_15687);
or U22988 (N_22988,N_17659,N_19668);
nand U22989 (N_22989,N_18155,N_16150);
nor U22990 (N_22990,N_16558,N_16262);
or U22991 (N_22991,N_19642,N_15212);
or U22992 (N_22992,N_15035,N_15949);
nor U22993 (N_22993,N_17070,N_18943);
and U22994 (N_22994,N_18068,N_18818);
or U22995 (N_22995,N_18452,N_16943);
nand U22996 (N_22996,N_18150,N_15692);
or U22997 (N_22997,N_17404,N_15435);
or U22998 (N_22998,N_18892,N_19785);
and U22999 (N_22999,N_18399,N_15779);
or U23000 (N_23000,N_19656,N_18834);
xor U23001 (N_23001,N_18475,N_16509);
xnor U23002 (N_23002,N_19244,N_17231);
or U23003 (N_23003,N_15914,N_17907);
or U23004 (N_23004,N_15501,N_19515);
xor U23005 (N_23005,N_17318,N_17587);
nand U23006 (N_23006,N_16704,N_16808);
and U23007 (N_23007,N_16539,N_19309);
and U23008 (N_23008,N_18305,N_16797);
or U23009 (N_23009,N_18349,N_16203);
or U23010 (N_23010,N_17725,N_17601);
nor U23011 (N_23011,N_16397,N_19507);
nor U23012 (N_23012,N_18355,N_17800);
nand U23013 (N_23013,N_17358,N_18215);
nor U23014 (N_23014,N_15585,N_17384);
or U23015 (N_23015,N_15037,N_15343);
and U23016 (N_23016,N_18185,N_15851);
nor U23017 (N_23017,N_19138,N_19476);
nand U23018 (N_23018,N_16425,N_18976);
and U23019 (N_23019,N_15363,N_18514);
or U23020 (N_23020,N_16987,N_15950);
xnor U23021 (N_23021,N_17122,N_15324);
xnor U23022 (N_23022,N_18490,N_17935);
nand U23023 (N_23023,N_18392,N_16799);
and U23024 (N_23024,N_15726,N_16069);
or U23025 (N_23025,N_18361,N_15024);
nand U23026 (N_23026,N_15737,N_16308);
and U23027 (N_23027,N_19835,N_19911);
nor U23028 (N_23028,N_16310,N_15903);
nand U23029 (N_23029,N_19525,N_18160);
nand U23030 (N_23030,N_15301,N_18467);
and U23031 (N_23031,N_15059,N_19448);
or U23032 (N_23032,N_19846,N_18190);
xnor U23033 (N_23033,N_16203,N_17051);
nand U23034 (N_23034,N_18667,N_18573);
and U23035 (N_23035,N_19984,N_17513);
and U23036 (N_23036,N_19258,N_15468);
and U23037 (N_23037,N_19762,N_15537);
and U23038 (N_23038,N_15742,N_16664);
or U23039 (N_23039,N_16971,N_16418);
or U23040 (N_23040,N_19684,N_19617);
and U23041 (N_23041,N_16119,N_18893);
nand U23042 (N_23042,N_19527,N_17069);
nand U23043 (N_23043,N_15732,N_17260);
and U23044 (N_23044,N_16055,N_15862);
and U23045 (N_23045,N_18726,N_19511);
nor U23046 (N_23046,N_19413,N_19708);
and U23047 (N_23047,N_16879,N_19627);
or U23048 (N_23048,N_18022,N_19888);
and U23049 (N_23049,N_18038,N_19319);
nand U23050 (N_23050,N_17555,N_16969);
nand U23051 (N_23051,N_19556,N_18439);
or U23052 (N_23052,N_18314,N_16208);
and U23053 (N_23053,N_17104,N_19138);
nand U23054 (N_23054,N_16999,N_18051);
and U23055 (N_23055,N_16373,N_18331);
and U23056 (N_23056,N_19368,N_18523);
or U23057 (N_23057,N_19939,N_16899);
nand U23058 (N_23058,N_19388,N_19187);
or U23059 (N_23059,N_16620,N_17618);
and U23060 (N_23060,N_17686,N_19780);
nand U23061 (N_23061,N_16220,N_16063);
xor U23062 (N_23062,N_18867,N_15242);
and U23063 (N_23063,N_18846,N_16789);
nand U23064 (N_23064,N_19163,N_19246);
and U23065 (N_23065,N_16815,N_17177);
nor U23066 (N_23066,N_15929,N_15868);
and U23067 (N_23067,N_16620,N_19022);
or U23068 (N_23068,N_17604,N_15819);
or U23069 (N_23069,N_15312,N_15038);
and U23070 (N_23070,N_15869,N_19620);
and U23071 (N_23071,N_15363,N_18732);
nand U23072 (N_23072,N_19694,N_15504);
nand U23073 (N_23073,N_17166,N_17906);
nor U23074 (N_23074,N_16085,N_18541);
nand U23075 (N_23075,N_15672,N_19449);
and U23076 (N_23076,N_19051,N_15397);
nand U23077 (N_23077,N_15402,N_16345);
nand U23078 (N_23078,N_15635,N_16472);
or U23079 (N_23079,N_17505,N_15296);
or U23080 (N_23080,N_17955,N_17885);
and U23081 (N_23081,N_17796,N_15763);
nand U23082 (N_23082,N_16134,N_19960);
nor U23083 (N_23083,N_18899,N_18593);
xnor U23084 (N_23084,N_16902,N_16889);
and U23085 (N_23085,N_15250,N_15003);
or U23086 (N_23086,N_17267,N_17159);
or U23087 (N_23087,N_18098,N_15682);
nand U23088 (N_23088,N_16757,N_18604);
nand U23089 (N_23089,N_15230,N_17645);
or U23090 (N_23090,N_16308,N_19734);
nand U23091 (N_23091,N_16942,N_19105);
and U23092 (N_23092,N_18062,N_17316);
nor U23093 (N_23093,N_18725,N_15292);
nand U23094 (N_23094,N_19458,N_15427);
nor U23095 (N_23095,N_18522,N_19095);
nor U23096 (N_23096,N_17913,N_15321);
nor U23097 (N_23097,N_18311,N_18548);
or U23098 (N_23098,N_18087,N_19253);
nor U23099 (N_23099,N_15685,N_16488);
nor U23100 (N_23100,N_15286,N_16562);
or U23101 (N_23101,N_16362,N_16509);
nor U23102 (N_23102,N_18636,N_16904);
xor U23103 (N_23103,N_17294,N_19355);
nor U23104 (N_23104,N_16093,N_18972);
nor U23105 (N_23105,N_18832,N_15980);
or U23106 (N_23106,N_18229,N_16472);
and U23107 (N_23107,N_17678,N_18725);
and U23108 (N_23108,N_19690,N_18282);
or U23109 (N_23109,N_16965,N_15099);
nor U23110 (N_23110,N_19783,N_19817);
nand U23111 (N_23111,N_19902,N_15974);
xor U23112 (N_23112,N_17338,N_19573);
nor U23113 (N_23113,N_19641,N_19724);
xor U23114 (N_23114,N_18106,N_17170);
xor U23115 (N_23115,N_19047,N_18064);
and U23116 (N_23116,N_17874,N_18924);
or U23117 (N_23117,N_19354,N_16735);
and U23118 (N_23118,N_17969,N_19029);
or U23119 (N_23119,N_17511,N_15938);
nor U23120 (N_23120,N_15970,N_17508);
nor U23121 (N_23121,N_19773,N_18362);
nand U23122 (N_23122,N_19447,N_19699);
and U23123 (N_23123,N_19645,N_16770);
nand U23124 (N_23124,N_17882,N_16624);
or U23125 (N_23125,N_15577,N_19301);
and U23126 (N_23126,N_15586,N_16577);
nor U23127 (N_23127,N_18610,N_17438);
and U23128 (N_23128,N_16662,N_16027);
xnor U23129 (N_23129,N_15106,N_18902);
or U23130 (N_23130,N_17111,N_18078);
xor U23131 (N_23131,N_19088,N_16271);
or U23132 (N_23132,N_17374,N_17362);
and U23133 (N_23133,N_18351,N_16818);
xor U23134 (N_23134,N_17303,N_16628);
or U23135 (N_23135,N_18825,N_19788);
and U23136 (N_23136,N_18471,N_18536);
and U23137 (N_23137,N_16312,N_17916);
xor U23138 (N_23138,N_18752,N_18617);
xor U23139 (N_23139,N_16351,N_17667);
and U23140 (N_23140,N_15694,N_18975);
and U23141 (N_23141,N_17715,N_15487);
nand U23142 (N_23142,N_18703,N_16117);
nand U23143 (N_23143,N_15388,N_15233);
nor U23144 (N_23144,N_15859,N_19885);
or U23145 (N_23145,N_18684,N_18769);
or U23146 (N_23146,N_18232,N_19163);
or U23147 (N_23147,N_16288,N_16350);
and U23148 (N_23148,N_17941,N_15617);
and U23149 (N_23149,N_17666,N_15325);
and U23150 (N_23150,N_19880,N_18967);
and U23151 (N_23151,N_16104,N_15097);
xnor U23152 (N_23152,N_17972,N_18754);
or U23153 (N_23153,N_17678,N_17080);
nand U23154 (N_23154,N_16983,N_18558);
or U23155 (N_23155,N_18102,N_16368);
or U23156 (N_23156,N_19586,N_15534);
nor U23157 (N_23157,N_16497,N_18535);
and U23158 (N_23158,N_19804,N_18098);
and U23159 (N_23159,N_15458,N_18590);
nor U23160 (N_23160,N_16747,N_17764);
nor U23161 (N_23161,N_16668,N_19874);
xnor U23162 (N_23162,N_19525,N_19945);
xor U23163 (N_23163,N_18535,N_17446);
nand U23164 (N_23164,N_19912,N_15676);
and U23165 (N_23165,N_18113,N_17321);
or U23166 (N_23166,N_15008,N_18777);
nand U23167 (N_23167,N_16469,N_16377);
xnor U23168 (N_23168,N_19215,N_19114);
nor U23169 (N_23169,N_17671,N_15738);
xor U23170 (N_23170,N_17859,N_17425);
or U23171 (N_23171,N_18726,N_17649);
nand U23172 (N_23172,N_16282,N_17503);
nor U23173 (N_23173,N_17916,N_16295);
or U23174 (N_23174,N_18561,N_16494);
nor U23175 (N_23175,N_15064,N_17147);
and U23176 (N_23176,N_15721,N_19512);
nand U23177 (N_23177,N_15024,N_17970);
and U23178 (N_23178,N_16015,N_18479);
or U23179 (N_23179,N_18134,N_19093);
nor U23180 (N_23180,N_16725,N_15505);
and U23181 (N_23181,N_17535,N_18486);
xnor U23182 (N_23182,N_17769,N_19651);
nor U23183 (N_23183,N_15053,N_16439);
xor U23184 (N_23184,N_17315,N_19852);
nor U23185 (N_23185,N_19280,N_18989);
or U23186 (N_23186,N_17281,N_19681);
xnor U23187 (N_23187,N_16110,N_18781);
xor U23188 (N_23188,N_18931,N_15076);
nor U23189 (N_23189,N_17593,N_19758);
and U23190 (N_23190,N_17558,N_19980);
and U23191 (N_23191,N_15104,N_16080);
xnor U23192 (N_23192,N_19393,N_17210);
nor U23193 (N_23193,N_19300,N_19543);
or U23194 (N_23194,N_15303,N_16466);
nand U23195 (N_23195,N_16063,N_19267);
and U23196 (N_23196,N_17302,N_16120);
nor U23197 (N_23197,N_15911,N_18950);
xor U23198 (N_23198,N_19635,N_17309);
nand U23199 (N_23199,N_16910,N_19405);
nor U23200 (N_23200,N_16521,N_15142);
nor U23201 (N_23201,N_16616,N_19022);
and U23202 (N_23202,N_18606,N_16215);
nor U23203 (N_23203,N_15117,N_16771);
xor U23204 (N_23204,N_17210,N_19729);
and U23205 (N_23205,N_16750,N_18425);
and U23206 (N_23206,N_19894,N_16918);
and U23207 (N_23207,N_17129,N_15949);
nand U23208 (N_23208,N_17899,N_15435);
and U23209 (N_23209,N_19112,N_15316);
xor U23210 (N_23210,N_16739,N_18821);
nor U23211 (N_23211,N_15677,N_18117);
nor U23212 (N_23212,N_15074,N_18521);
or U23213 (N_23213,N_19153,N_15525);
nor U23214 (N_23214,N_16554,N_17796);
nand U23215 (N_23215,N_19253,N_18861);
or U23216 (N_23216,N_19845,N_18528);
or U23217 (N_23217,N_16264,N_15334);
nand U23218 (N_23218,N_17446,N_17687);
xor U23219 (N_23219,N_19244,N_18551);
nor U23220 (N_23220,N_17336,N_15841);
or U23221 (N_23221,N_19253,N_16799);
or U23222 (N_23222,N_18469,N_18693);
nand U23223 (N_23223,N_17140,N_16278);
and U23224 (N_23224,N_17921,N_19061);
nor U23225 (N_23225,N_17185,N_15243);
nand U23226 (N_23226,N_15401,N_15867);
nand U23227 (N_23227,N_18620,N_17471);
xor U23228 (N_23228,N_18405,N_16948);
and U23229 (N_23229,N_17695,N_19728);
xnor U23230 (N_23230,N_18861,N_15249);
nor U23231 (N_23231,N_16878,N_19538);
or U23232 (N_23232,N_19834,N_16849);
nand U23233 (N_23233,N_17521,N_18903);
and U23234 (N_23234,N_18869,N_16939);
nand U23235 (N_23235,N_16119,N_19196);
and U23236 (N_23236,N_17534,N_17566);
nand U23237 (N_23237,N_15361,N_17919);
nor U23238 (N_23238,N_18807,N_19787);
and U23239 (N_23239,N_16006,N_19115);
or U23240 (N_23240,N_17281,N_18163);
xnor U23241 (N_23241,N_17181,N_17627);
and U23242 (N_23242,N_18243,N_19832);
nand U23243 (N_23243,N_15594,N_16996);
or U23244 (N_23244,N_17827,N_15951);
nor U23245 (N_23245,N_18521,N_15909);
or U23246 (N_23246,N_17440,N_17452);
and U23247 (N_23247,N_15416,N_18922);
and U23248 (N_23248,N_17207,N_16862);
or U23249 (N_23249,N_15832,N_15458);
nor U23250 (N_23250,N_17152,N_15459);
nor U23251 (N_23251,N_19921,N_15690);
nand U23252 (N_23252,N_15349,N_19489);
nand U23253 (N_23253,N_18626,N_17526);
and U23254 (N_23254,N_18080,N_15947);
nor U23255 (N_23255,N_15842,N_16965);
or U23256 (N_23256,N_15596,N_16484);
and U23257 (N_23257,N_16495,N_17735);
and U23258 (N_23258,N_16260,N_15431);
or U23259 (N_23259,N_15673,N_18591);
nor U23260 (N_23260,N_19760,N_15394);
nor U23261 (N_23261,N_17279,N_17249);
xor U23262 (N_23262,N_18814,N_15310);
nand U23263 (N_23263,N_18800,N_15782);
xnor U23264 (N_23264,N_15222,N_16252);
nand U23265 (N_23265,N_16353,N_17017);
nor U23266 (N_23266,N_18777,N_19700);
nand U23267 (N_23267,N_16421,N_19311);
nor U23268 (N_23268,N_19034,N_15261);
and U23269 (N_23269,N_16871,N_17690);
nand U23270 (N_23270,N_15950,N_19749);
or U23271 (N_23271,N_15254,N_15704);
xnor U23272 (N_23272,N_19342,N_19057);
nand U23273 (N_23273,N_19624,N_17999);
and U23274 (N_23274,N_15855,N_17081);
nor U23275 (N_23275,N_17033,N_16855);
nor U23276 (N_23276,N_18834,N_18615);
nand U23277 (N_23277,N_17041,N_15802);
xor U23278 (N_23278,N_18280,N_19680);
and U23279 (N_23279,N_19929,N_17860);
nand U23280 (N_23280,N_17201,N_19486);
or U23281 (N_23281,N_15160,N_19869);
or U23282 (N_23282,N_16416,N_16301);
nor U23283 (N_23283,N_19656,N_17175);
nand U23284 (N_23284,N_16587,N_17907);
or U23285 (N_23285,N_18559,N_16301);
nand U23286 (N_23286,N_16763,N_15474);
nor U23287 (N_23287,N_15415,N_19970);
nand U23288 (N_23288,N_16420,N_15917);
and U23289 (N_23289,N_15303,N_19359);
nand U23290 (N_23290,N_16914,N_16876);
nor U23291 (N_23291,N_19643,N_15286);
or U23292 (N_23292,N_16364,N_17732);
nand U23293 (N_23293,N_15075,N_18603);
or U23294 (N_23294,N_15945,N_16797);
and U23295 (N_23295,N_15618,N_15381);
nor U23296 (N_23296,N_18579,N_16308);
or U23297 (N_23297,N_19718,N_18769);
and U23298 (N_23298,N_16286,N_17803);
nand U23299 (N_23299,N_16242,N_19054);
xnor U23300 (N_23300,N_18636,N_16689);
or U23301 (N_23301,N_19754,N_17983);
nor U23302 (N_23302,N_15414,N_17508);
xor U23303 (N_23303,N_15618,N_19422);
nand U23304 (N_23304,N_16497,N_16853);
nand U23305 (N_23305,N_17218,N_19224);
or U23306 (N_23306,N_16633,N_18923);
nor U23307 (N_23307,N_16950,N_16410);
nand U23308 (N_23308,N_15428,N_15682);
nand U23309 (N_23309,N_17441,N_17082);
and U23310 (N_23310,N_15807,N_17436);
or U23311 (N_23311,N_15014,N_17107);
nand U23312 (N_23312,N_16138,N_18054);
and U23313 (N_23313,N_17184,N_16954);
and U23314 (N_23314,N_16561,N_16188);
or U23315 (N_23315,N_15585,N_15246);
or U23316 (N_23316,N_16005,N_15475);
or U23317 (N_23317,N_17603,N_18722);
nor U23318 (N_23318,N_16968,N_17867);
or U23319 (N_23319,N_16698,N_18859);
nand U23320 (N_23320,N_18261,N_19481);
nor U23321 (N_23321,N_19279,N_16637);
nand U23322 (N_23322,N_16121,N_15654);
nor U23323 (N_23323,N_19041,N_18580);
nor U23324 (N_23324,N_18435,N_18552);
nand U23325 (N_23325,N_18955,N_15284);
or U23326 (N_23326,N_19871,N_16746);
nor U23327 (N_23327,N_16678,N_17428);
or U23328 (N_23328,N_17124,N_15250);
or U23329 (N_23329,N_15709,N_19027);
and U23330 (N_23330,N_15567,N_16101);
or U23331 (N_23331,N_16225,N_19647);
nand U23332 (N_23332,N_17244,N_16283);
nand U23333 (N_23333,N_19051,N_17005);
xnor U23334 (N_23334,N_17071,N_17477);
nand U23335 (N_23335,N_17275,N_16341);
nor U23336 (N_23336,N_18445,N_18507);
xor U23337 (N_23337,N_15513,N_19418);
and U23338 (N_23338,N_17198,N_19438);
xnor U23339 (N_23339,N_18022,N_19027);
and U23340 (N_23340,N_17271,N_15916);
nor U23341 (N_23341,N_17731,N_15932);
nor U23342 (N_23342,N_18131,N_18564);
or U23343 (N_23343,N_19736,N_15841);
and U23344 (N_23344,N_18848,N_19721);
and U23345 (N_23345,N_19953,N_15990);
and U23346 (N_23346,N_17486,N_18719);
nand U23347 (N_23347,N_15859,N_17315);
nor U23348 (N_23348,N_17449,N_16051);
nand U23349 (N_23349,N_16042,N_15495);
nand U23350 (N_23350,N_17610,N_18072);
nor U23351 (N_23351,N_15384,N_18363);
nand U23352 (N_23352,N_17854,N_16615);
nor U23353 (N_23353,N_16272,N_15024);
nand U23354 (N_23354,N_15329,N_15020);
nand U23355 (N_23355,N_18761,N_17325);
nand U23356 (N_23356,N_16600,N_18332);
nor U23357 (N_23357,N_15863,N_16046);
or U23358 (N_23358,N_18395,N_17452);
xnor U23359 (N_23359,N_17564,N_16253);
and U23360 (N_23360,N_16147,N_15749);
nand U23361 (N_23361,N_16679,N_16615);
and U23362 (N_23362,N_19830,N_18488);
nand U23363 (N_23363,N_15568,N_17659);
or U23364 (N_23364,N_16453,N_15850);
nor U23365 (N_23365,N_18906,N_17738);
or U23366 (N_23366,N_17692,N_15175);
nor U23367 (N_23367,N_16209,N_18143);
or U23368 (N_23368,N_19586,N_18191);
xnor U23369 (N_23369,N_18320,N_18549);
nor U23370 (N_23370,N_17808,N_16909);
nand U23371 (N_23371,N_16965,N_19172);
or U23372 (N_23372,N_18589,N_18864);
or U23373 (N_23373,N_19215,N_17691);
nand U23374 (N_23374,N_15452,N_15721);
nor U23375 (N_23375,N_18644,N_18116);
nor U23376 (N_23376,N_17487,N_15345);
nor U23377 (N_23377,N_15241,N_15026);
or U23378 (N_23378,N_18631,N_15734);
nor U23379 (N_23379,N_15586,N_16893);
nand U23380 (N_23380,N_18470,N_17792);
or U23381 (N_23381,N_19340,N_19505);
nand U23382 (N_23382,N_16006,N_17543);
or U23383 (N_23383,N_19871,N_17989);
or U23384 (N_23384,N_19245,N_15461);
nand U23385 (N_23385,N_18332,N_19166);
and U23386 (N_23386,N_18261,N_16069);
and U23387 (N_23387,N_17841,N_16125);
nand U23388 (N_23388,N_15691,N_18532);
nand U23389 (N_23389,N_18252,N_16055);
and U23390 (N_23390,N_19418,N_18414);
nand U23391 (N_23391,N_15637,N_16986);
nor U23392 (N_23392,N_17594,N_16781);
xnor U23393 (N_23393,N_19782,N_16668);
or U23394 (N_23394,N_19299,N_15666);
nor U23395 (N_23395,N_18235,N_18901);
nor U23396 (N_23396,N_16773,N_17705);
nor U23397 (N_23397,N_19998,N_18652);
xor U23398 (N_23398,N_18180,N_17207);
or U23399 (N_23399,N_18663,N_19928);
nor U23400 (N_23400,N_17359,N_15204);
or U23401 (N_23401,N_15250,N_18470);
and U23402 (N_23402,N_17791,N_17662);
and U23403 (N_23403,N_16599,N_18201);
nand U23404 (N_23404,N_16249,N_17502);
nand U23405 (N_23405,N_16335,N_15131);
nor U23406 (N_23406,N_15120,N_19008);
xnor U23407 (N_23407,N_15429,N_16936);
nand U23408 (N_23408,N_19157,N_15362);
or U23409 (N_23409,N_16879,N_16477);
nand U23410 (N_23410,N_16167,N_18374);
or U23411 (N_23411,N_19209,N_16536);
xor U23412 (N_23412,N_17018,N_16380);
nor U23413 (N_23413,N_18568,N_17265);
xnor U23414 (N_23414,N_17020,N_17104);
nor U23415 (N_23415,N_18804,N_16965);
and U23416 (N_23416,N_16200,N_16213);
nand U23417 (N_23417,N_18965,N_17019);
nand U23418 (N_23418,N_16844,N_17243);
or U23419 (N_23419,N_19663,N_17016);
or U23420 (N_23420,N_15538,N_16132);
and U23421 (N_23421,N_18405,N_15522);
or U23422 (N_23422,N_18900,N_19916);
and U23423 (N_23423,N_16839,N_19383);
nor U23424 (N_23424,N_19118,N_15989);
and U23425 (N_23425,N_19768,N_17481);
or U23426 (N_23426,N_17288,N_19594);
or U23427 (N_23427,N_15122,N_16328);
nor U23428 (N_23428,N_18095,N_16048);
and U23429 (N_23429,N_19190,N_17928);
nor U23430 (N_23430,N_15425,N_17285);
nand U23431 (N_23431,N_19740,N_18344);
and U23432 (N_23432,N_16155,N_18900);
xnor U23433 (N_23433,N_19632,N_19031);
nand U23434 (N_23434,N_15706,N_18159);
or U23435 (N_23435,N_15155,N_17304);
or U23436 (N_23436,N_18058,N_15764);
nor U23437 (N_23437,N_17182,N_15675);
or U23438 (N_23438,N_19961,N_18026);
nand U23439 (N_23439,N_19328,N_16790);
nand U23440 (N_23440,N_16929,N_17243);
nor U23441 (N_23441,N_16709,N_17040);
and U23442 (N_23442,N_17982,N_19947);
or U23443 (N_23443,N_15354,N_17609);
and U23444 (N_23444,N_16754,N_16748);
nand U23445 (N_23445,N_15616,N_17716);
and U23446 (N_23446,N_17894,N_19246);
nand U23447 (N_23447,N_16289,N_19883);
xnor U23448 (N_23448,N_19593,N_19915);
nand U23449 (N_23449,N_17503,N_19913);
nand U23450 (N_23450,N_19497,N_17483);
nand U23451 (N_23451,N_19120,N_17922);
and U23452 (N_23452,N_18336,N_15365);
nand U23453 (N_23453,N_16546,N_16775);
nand U23454 (N_23454,N_16017,N_18366);
nor U23455 (N_23455,N_15344,N_15994);
nand U23456 (N_23456,N_18969,N_19258);
and U23457 (N_23457,N_17719,N_15082);
and U23458 (N_23458,N_15041,N_15754);
or U23459 (N_23459,N_17175,N_17036);
or U23460 (N_23460,N_19077,N_15059);
nor U23461 (N_23461,N_18851,N_17613);
and U23462 (N_23462,N_15389,N_17482);
and U23463 (N_23463,N_15656,N_19497);
nand U23464 (N_23464,N_17541,N_16680);
or U23465 (N_23465,N_16242,N_19215);
and U23466 (N_23466,N_16122,N_19327);
and U23467 (N_23467,N_15987,N_19770);
and U23468 (N_23468,N_15059,N_15884);
nor U23469 (N_23469,N_18631,N_17099);
or U23470 (N_23470,N_17288,N_19417);
or U23471 (N_23471,N_16854,N_18144);
xnor U23472 (N_23472,N_19911,N_16996);
xnor U23473 (N_23473,N_17117,N_15390);
nand U23474 (N_23474,N_15206,N_16899);
nand U23475 (N_23475,N_18920,N_15265);
and U23476 (N_23476,N_19967,N_18243);
nor U23477 (N_23477,N_19665,N_18838);
nor U23478 (N_23478,N_19307,N_18563);
or U23479 (N_23479,N_17426,N_19214);
and U23480 (N_23480,N_19659,N_19066);
nor U23481 (N_23481,N_18855,N_17716);
or U23482 (N_23482,N_19144,N_19207);
nor U23483 (N_23483,N_18580,N_19280);
nand U23484 (N_23484,N_19150,N_16570);
and U23485 (N_23485,N_19144,N_17488);
and U23486 (N_23486,N_16847,N_17076);
or U23487 (N_23487,N_17352,N_18739);
and U23488 (N_23488,N_19919,N_16316);
xnor U23489 (N_23489,N_17842,N_16440);
nor U23490 (N_23490,N_19658,N_18135);
xor U23491 (N_23491,N_15971,N_18396);
or U23492 (N_23492,N_19136,N_17693);
nor U23493 (N_23493,N_16770,N_16828);
nor U23494 (N_23494,N_16336,N_17232);
nor U23495 (N_23495,N_15149,N_16804);
nor U23496 (N_23496,N_19042,N_16627);
xnor U23497 (N_23497,N_19283,N_17904);
and U23498 (N_23498,N_17684,N_16250);
and U23499 (N_23499,N_19755,N_19046);
xor U23500 (N_23500,N_18223,N_15663);
nand U23501 (N_23501,N_16437,N_17765);
and U23502 (N_23502,N_15903,N_17520);
xor U23503 (N_23503,N_18303,N_19054);
xnor U23504 (N_23504,N_18774,N_17513);
nor U23505 (N_23505,N_19812,N_18129);
nor U23506 (N_23506,N_15907,N_15593);
or U23507 (N_23507,N_17503,N_16263);
nor U23508 (N_23508,N_19939,N_15436);
nor U23509 (N_23509,N_16752,N_15056);
or U23510 (N_23510,N_17141,N_18172);
nand U23511 (N_23511,N_16156,N_19554);
or U23512 (N_23512,N_16098,N_17385);
and U23513 (N_23513,N_15369,N_19727);
xnor U23514 (N_23514,N_19331,N_16210);
nand U23515 (N_23515,N_16977,N_16062);
nand U23516 (N_23516,N_16971,N_19692);
nand U23517 (N_23517,N_15997,N_19022);
or U23518 (N_23518,N_15432,N_16129);
or U23519 (N_23519,N_15092,N_16598);
or U23520 (N_23520,N_16885,N_15541);
nor U23521 (N_23521,N_17430,N_19288);
nor U23522 (N_23522,N_19445,N_16882);
nand U23523 (N_23523,N_19830,N_16904);
or U23524 (N_23524,N_17839,N_15361);
nor U23525 (N_23525,N_19959,N_18272);
nor U23526 (N_23526,N_16803,N_16105);
or U23527 (N_23527,N_15292,N_16670);
and U23528 (N_23528,N_16869,N_16549);
nor U23529 (N_23529,N_16180,N_19201);
or U23530 (N_23530,N_19840,N_17531);
or U23531 (N_23531,N_17085,N_15032);
or U23532 (N_23532,N_18612,N_18972);
nor U23533 (N_23533,N_15188,N_19864);
and U23534 (N_23534,N_18012,N_15041);
nor U23535 (N_23535,N_15076,N_17600);
xor U23536 (N_23536,N_17060,N_18568);
or U23537 (N_23537,N_18757,N_19133);
nor U23538 (N_23538,N_19538,N_19021);
and U23539 (N_23539,N_17622,N_15108);
xor U23540 (N_23540,N_19373,N_16755);
nand U23541 (N_23541,N_18394,N_15169);
nand U23542 (N_23542,N_15358,N_15896);
xor U23543 (N_23543,N_16743,N_19621);
nor U23544 (N_23544,N_15480,N_18611);
nand U23545 (N_23545,N_19226,N_19083);
and U23546 (N_23546,N_19427,N_17621);
or U23547 (N_23547,N_15883,N_16250);
or U23548 (N_23548,N_17485,N_15263);
or U23549 (N_23549,N_17185,N_18262);
or U23550 (N_23550,N_17248,N_17622);
nor U23551 (N_23551,N_19416,N_15132);
nor U23552 (N_23552,N_15772,N_15010);
and U23553 (N_23553,N_17526,N_15620);
xnor U23554 (N_23554,N_16350,N_17966);
or U23555 (N_23555,N_18798,N_18861);
or U23556 (N_23556,N_15115,N_15166);
and U23557 (N_23557,N_16368,N_16976);
or U23558 (N_23558,N_16585,N_19146);
nor U23559 (N_23559,N_15845,N_17959);
or U23560 (N_23560,N_19682,N_18809);
and U23561 (N_23561,N_16190,N_18339);
nand U23562 (N_23562,N_15999,N_16295);
and U23563 (N_23563,N_17008,N_19262);
or U23564 (N_23564,N_17286,N_19527);
nand U23565 (N_23565,N_18430,N_17710);
or U23566 (N_23566,N_19727,N_16913);
nor U23567 (N_23567,N_19514,N_18190);
or U23568 (N_23568,N_17339,N_19194);
nand U23569 (N_23569,N_17866,N_19236);
or U23570 (N_23570,N_17958,N_17480);
or U23571 (N_23571,N_18913,N_16290);
or U23572 (N_23572,N_19825,N_15831);
and U23573 (N_23573,N_19116,N_16448);
nor U23574 (N_23574,N_16800,N_19752);
nor U23575 (N_23575,N_17654,N_15324);
and U23576 (N_23576,N_15745,N_17579);
nand U23577 (N_23577,N_15847,N_16056);
or U23578 (N_23578,N_17659,N_19353);
nor U23579 (N_23579,N_16679,N_17610);
nand U23580 (N_23580,N_18334,N_15979);
nor U23581 (N_23581,N_17685,N_15724);
nor U23582 (N_23582,N_15772,N_17721);
and U23583 (N_23583,N_16931,N_15213);
nor U23584 (N_23584,N_18021,N_17313);
nor U23585 (N_23585,N_15599,N_17558);
nand U23586 (N_23586,N_17900,N_16096);
nand U23587 (N_23587,N_18987,N_19926);
nor U23588 (N_23588,N_18318,N_16361);
and U23589 (N_23589,N_15286,N_15345);
nand U23590 (N_23590,N_19043,N_15871);
nand U23591 (N_23591,N_17236,N_16767);
nand U23592 (N_23592,N_15231,N_15335);
or U23593 (N_23593,N_15810,N_16128);
nor U23594 (N_23594,N_19035,N_19533);
or U23595 (N_23595,N_17223,N_17501);
nor U23596 (N_23596,N_18971,N_15105);
nand U23597 (N_23597,N_17895,N_19973);
or U23598 (N_23598,N_18688,N_15547);
nor U23599 (N_23599,N_17387,N_15832);
nand U23600 (N_23600,N_16801,N_17735);
or U23601 (N_23601,N_17891,N_16674);
xor U23602 (N_23602,N_18328,N_17149);
and U23603 (N_23603,N_16247,N_19721);
nand U23604 (N_23604,N_16208,N_17568);
nand U23605 (N_23605,N_18464,N_15616);
and U23606 (N_23606,N_16238,N_16598);
xor U23607 (N_23607,N_19032,N_15785);
or U23608 (N_23608,N_18595,N_17981);
and U23609 (N_23609,N_15362,N_17305);
and U23610 (N_23610,N_17948,N_18361);
xor U23611 (N_23611,N_19621,N_17477);
nand U23612 (N_23612,N_19344,N_15743);
nor U23613 (N_23613,N_15859,N_18537);
nand U23614 (N_23614,N_18158,N_18425);
nand U23615 (N_23615,N_15375,N_17954);
nor U23616 (N_23616,N_17942,N_17794);
nand U23617 (N_23617,N_17150,N_17544);
nor U23618 (N_23618,N_18322,N_15011);
nor U23619 (N_23619,N_15254,N_16828);
and U23620 (N_23620,N_19480,N_15180);
or U23621 (N_23621,N_18411,N_18124);
nor U23622 (N_23622,N_19441,N_17689);
xnor U23623 (N_23623,N_17318,N_19129);
nor U23624 (N_23624,N_15174,N_15935);
or U23625 (N_23625,N_16272,N_16999);
and U23626 (N_23626,N_18050,N_15313);
or U23627 (N_23627,N_17462,N_17787);
or U23628 (N_23628,N_15711,N_19028);
xor U23629 (N_23629,N_16218,N_15078);
or U23630 (N_23630,N_15315,N_17739);
and U23631 (N_23631,N_17216,N_18923);
and U23632 (N_23632,N_15205,N_15025);
and U23633 (N_23633,N_18261,N_16681);
nor U23634 (N_23634,N_17478,N_18053);
nor U23635 (N_23635,N_18437,N_15615);
nor U23636 (N_23636,N_15394,N_16545);
nand U23637 (N_23637,N_18418,N_16504);
nand U23638 (N_23638,N_19310,N_15392);
xor U23639 (N_23639,N_17445,N_16790);
nand U23640 (N_23640,N_15187,N_15625);
or U23641 (N_23641,N_17937,N_19284);
xor U23642 (N_23642,N_19859,N_18557);
or U23643 (N_23643,N_15196,N_16934);
nand U23644 (N_23644,N_16407,N_16339);
nor U23645 (N_23645,N_16821,N_19147);
and U23646 (N_23646,N_18279,N_18132);
and U23647 (N_23647,N_18046,N_16517);
nand U23648 (N_23648,N_15762,N_16709);
nor U23649 (N_23649,N_19563,N_18785);
nand U23650 (N_23650,N_15730,N_15798);
and U23651 (N_23651,N_16768,N_17569);
nand U23652 (N_23652,N_15475,N_16968);
nand U23653 (N_23653,N_15254,N_15948);
or U23654 (N_23654,N_16310,N_18899);
nor U23655 (N_23655,N_18869,N_19306);
and U23656 (N_23656,N_17300,N_16653);
or U23657 (N_23657,N_16562,N_17310);
nor U23658 (N_23658,N_16372,N_19500);
nor U23659 (N_23659,N_19451,N_15993);
and U23660 (N_23660,N_16257,N_18709);
nor U23661 (N_23661,N_16193,N_15821);
nand U23662 (N_23662,N_17225,N_16083);
nor U23663 (N_23663,N_19159,N_18264);
nor U23664 (N_23664,N_15898,N_16832);
or U23665 (N_23665,N_16812,N_16959);
xnor U23666 (N_23666,N_15531,N_16017);
nand U23667 (N_23667,N_15384,N_18945);
and U23668 (N_23668,N_15102,N_18385);
or U23669 (N_23669,N_16080,N_15178);
and U23670 (N_23670,N_19904,N_15075);
nor U23671 (N_23671,N_17376,N_19983);
nand U23672 (N_23672,N_17560,N_15018);
xor U23673 (N_23673,N_19293,N_18744);
and U23674 (N_23674,N_17668,N_17791);
nor U23675 (N_23675,N_18565,N_19199);
and U23676 (N_23676,N_18896,N_18323);
xnor U23677 (N_23677,N_15585,N_16086);
nor U23678 (N_23678,N_18934,N_17803);
nor U23679 (N_23679,N_19529,N_15151);
or U23680 (N_23680,N_17915,N_18384);
xor U23681 (N_23681,N_15292,N_19466);
or U23682 (N_23682,N_19902,N_15130);
or U23683 (N_23683,N_18941,N_16929);
nor U23684 (N_23684,N_16887,N_18576);
or U23685 (N_23685,N_15152,N_16360);
or U23686 (N_23686,N_19782,N_19013);
nor U23687 (N_23687,N_16068,N_18189);
nor U23688 (N_23688,N_15429,N_18307);
xnor U23689 (N_23689,N_17693,N_17843);
nor U23690 (N_23690,N_18070,N_15579);
nand U23691 (N_23691,N_16028,N_17878);
nor U23692 (N_23692,N_16603,N_17816);
nand U23693 (N_23693,N_18360,N_19672);
nand U23694 (N_23694,N_15912,N_16992);
nor U23695 (N_23695,N_19560,N_15826);
or U23696 (N_23696,N_18287,N_15458);
or U23697 (N_23697,N_16309,N_19566);
or U23698 (N_23698,N_19557,N_17065);
nand U23699 (N_23699,N_16687,N_16106);
or U23700 (N_23700,N_19755,N_17446);
or U23701 (N_23701,N_15191,N_15565);
nand U23702 (N_23702,N_15588,N_15010);
nand U23703 (N_23703,N_17835,N_16046);
nand U23704 (N_23704,N_19632,N_17459);
or U23705 (N_23705,N_18841,N_18272);
or U23706 (N_23706,N_16955,N_15989);
nand U23707 (N_23707,N_18433,N_19666);
nand U23708 (N_23708,N_18790,N_19310);
nor U23709 (N_23709,N_18535,N_16090);
nand U23710 (N_23710,N_17308,N_17711);
and U23711 (N_23711,N_17174,N_17287);
nand U23712 (N_23712,N_19728,N_19384);
and U23713 (N_23713,N_15300,N_16432);
and U23714 (N_23714,N_15725,N_15401);
and U23715 (N_23715,N_18242,N_15975);
xor U23716 (N_23716,N_18890,N_15842);
xor U23717 (N_23717,N_18362,N_15943);
and U23718 (N_23718,N_16150,N_16955);
and U23719 (N_23719,N_16697,N_15476);
nor U23720 (N_23720,N_18076,N_17972);
nor U23721 (N_23721,N_15679,N_18985);
or U23722 (N_23722,N_19516,N_15756);
and U23723 (N_23723,N_17035,N_19202);
nor U23724 (N_23724,N_15703,N_16801);
or U23725 (N_23725,N_18955,N_18827);
xor U23726 (N_23726,N_15956,N_16615);
or U23727 (N_23727,N_17066,N_16295);
xnor U23728 (N_23728,N_15939,N_16474);
nor U23729 (N_23729,N_15455,N_16153);
and U23730 (N_23730,N_15143,N_18890);
xnor U23731 (N_23731,N_16468,N_17812);
and U23732 (N_23732,N_16284,N_17125);
nor U23733 (N_23733,N_15139,N_18658);
or U23734 (N_23734,N_18324,N_16121);
or U23735 (N_23735,N_16841,N_15440);
xor U23736 (N_23736,N_19893,N_17772);
nand U23737 (N_23737,N_18472,N_18085);
or U23738 (N_23738,N_17987,N_19511);
and U23739 (N_23739,N_16255,N_18600);
nand U23740 (N_23740,N_19447,N_15282);
xor U23741 (N_23741,N_17411,N_17482);
nor U23742 (N_23742,N_15773,N_19325);
nor U23743 (N_23743,N_18691,N_15091);
nand U23744 (N_23744,N_17206,N_16038);
or U23745 (N_23745,N_17678,N_19068);
nor U23746 (N_23746,N_17741,N_16423);
or U23747 (N_23747,N_17302,N_16143);
or U23748 (N_23748,N_16620,N_16003);
nand U23749 (N_23749,N_17716,N_17337);
and U23750 (N_23750,N_16913,N_19236);
xnor U23751 (N_23751,N_19675,N_15391);
or U23752 (N_23752,N_16361,N_17847);
nor U23753 (N_23753,N_17895,N_18969);
nand U23754 (N_23754,N_15913,N_15044);
nor U23755 (N_23755,N_15558,N_17206);
nand U23756 (N_23756,N_15946,N_16502);
nor U23757 (N_23757,N_19412,N_19568);
nand U23758 (N_23758,N_15084,N_16278);
nand U23759 (N_23759,N_19855,N_17541);
and U23760 (N_23760,N_19106,N_16576);
nor U23761 (N_23761,N_16564,N_19433);
nand U23762 (N_23762,N_19309,N_18492);
and U23763 (N_23763,N_18468,N_18377);
nand U23764 (N_23764,N_17201,N_18232);
or U23765 (N_23765,N_18019,N_15690);
and U23766 (N_23766,N_19388,N_15153);
xnor U23767 (N_23767,N_16423,N_15879);
nor U23768 (N_23768,N_16370,N_16740);
or U23769 (N_23769,N_16408,N_16587);
xor U23770 (N_23770,N_18185,N_18559);
or U23771 (N_23771,N_16348,N_16771);
nor U23772 (N_23772,N_19402,N_16241);
and U23773 (N_23773,N_15924,N_17428);
or U23774 (N_23774,N_15508,N_16405);
nor U23775 (N_23775,N_19093,N_18618);
nand U23776 (N_23776,N_17907,N_18416);
nand U23777 (N_23777,N_19417,N_17974);
and U23778 (N_23778,N_16505,N_19715);
nand U23779 (N_23779,N_17563,N_16709);
or U23780 (N_23780,N_15012,N_15101);
and U23781 (N_23781,N_18310,N_18055);
nor U23782 (N_23782,N_17645,N_16872);
and U23783 (N_23783,N_19544,N_19641);
nand U23784 (N_23784,N_15325,N_16986);
nor U23785 (N_23785,N_19391,N_18818);
or U23786 (N_23786,N_16830,N_15914);
nand U23787 (N_23787,N_15705,N_15087);
nand U23788 (N_23788,N_17322,N_17221);
nand U23789 (N_23789,N_18288,N_15867);
and U23790 (N_23790,N_16680,N_15771);
xor U23791 (N_23791,N_18356,N_15584);
and U23792 (N_23792,N_19539,N_19542);
or U23793 (N_23793,N_15360,N_16275);
and U23794 (N_23794,N_17669,N_19001);
nor U23795 (N_23795,N_17605,N_18684);
nor U23796 (N_23796,N_17097,N_17264);
xor U23797 (N_23797,N_18137,N_16086);
nand U23798 (N_23798,N_18623,N_19722);
nand U23799 (N_23799,N_18703,N_18012);
xor U23800 (N_23800,N_17025,N_17850);
or U23801 (N_23801,N_18189,N_17234);
and U23802 (N_23802,N_17902,N_19732);
nand U23803 (N_23803,N_17573,N_17547);
xor U23804 (N_23804,N_16240,N_15915);
and U23805 (N_23805,N_15492,N_16230);
or U23806 (N_23806,N_16077,N_16579);
nor U23807 (N_23807,N_15006,N_19466);
or U23808 (N_23808,N_18040,N_19071);
nand U23809 (N_23809,N_16456,N_19436);
nor U23810 (N_23810,N_19472,N_19701);
nand U23811 (N_23811,N_18726,N_16543);
nand U23812 (N_23812,N_16170,N_15915);
and U23813 (N_23813,N_17948,N_17753);
nor U23814 (N_23814,N_16296,N_18819);
or U23815 (N_23815,N_17491,N_18031);
or U23816 (N_23816,N_16586,N_15837);
nand U23817 (N_23817,N_15700,N_17482);
nor U23818 (N_23818,N_18120,N_18040);
nor U23819 (N_23819,N_15020,N_17527);
or U23820 (N_23820,N_18756,N_19056);
nor U23821 (N_23821,N_17468,N_17271);
nand U23822 (N_23822,N_15406,N_19895);
or U23823 (N_23823,N_18174,N_16944);
and U23824 (N_23824,N_18423,N_15366);
nor U23825 (N_23825,N_18469,N_19886);
or U23826 (N_23826,N_18551,N_16389);
nor U23827 (N_23827,N_16322,N_19709);
or U23828 (N_23828,N_16421,N_19784);
nor U23829 (N_23829,N_18530,N_17768);
and U23830 (N_23830,N_18567,N_19992);
and U23831 (N_23831,N_16328,N_15221);
xor U23832 (N_23832,N_16030,N_17044);
and U23833 (N_23833,N_18706,N_16704);
nor U23834 (N_23834,N_15297,N_19226);
nor U23835 (N_23835,N_19400,N_16697);
and U23836 (N_23836,N_19258,N_19929);
xor U23837 (N_23837,N_17161,N_16939);
and U23838 (N_23838,N_17439,N_15448);
nor U23839 (N_23839,N_19036,N_15905);
nand U23840 (N_23840,N_18165,N_16887);
nand U23841 (N_23841,N_19953,N_16988);
and U23842 (N_23842,N_19531,N_19315);
or U23843 (N_23843,N_15863,N_18385);
nor U23844 (N_23844,N_17149,N_18236);
nand U23845 (N_23845,N_19895,N_17763);
and U23846 (N_23846,N_15934,N_15482);
or U23847 (N_23847,N_16902,N_17526);
nand U23848 (N_23848,N_18750,N_18625);
and U23849 (N_23849,N_18898,N_17484);
or U23850 (N_23850,N_15482,N_15444);
nand U23851 (N_23851,N_15418,N_18011);
nor U23852 (N_23852,N_17106,N_15220);
nand U23853 (N_23853,N_16210,N_18781);
nor U23854 (N_23854,N_15059,N_17614);
and U23855 (N_23855,N_18433,N_19391);
and U23856 (N_23856,N_17368,N_18488);
and U23857 (N_23857,N_19496,N_19455);
nand U23858 (N_23858,N_17285,N_18550);
and U23859 (N_23859,N_16372,N_19235);
and U23860 (N_23860,N_17866,N_19366);
nand U23861 (N_23861,N_19926,N_15462);
and U23862 (N_23862,N_17558,N_19726);
nor U23863 (N_23863,N_16760,N_16419);
nand U23864 (N_23864,N_16518,N_16905);
or U23865 (N_23865,N_18643,N_17256);
or U23866 (N_23866,N_19015,N_15457);
xor U23867 (N_23867,N_17358,N_17080);
nand U23868 (N_23868,N_17358,N_18816);
and U23869 (N_23869,N_19787,N_18766);
or U23870 (N_23870,N_15386,N_15591);
and U23871 (N_23871,N_16979,N_19146);
and U23872 (N_23872,N_19471,N_19229);
and U23873 (N_23873,N_15020,N_19540);
nand U23874 (N_23874,N_16106,N_15897);
nand U23875 (N_23875,N_16894,N_16114);
and U23876 (N_23876,N_18024,N_19650);
and U23877 (N_23877,N_15899,N_17014);
nand U23878 (N_23878,N_15673,N_16521);
and U23879 (N_23879,N_16699,N_19936);
and U23880 (N_23880,N_16291,N_18353);
or U23881 (N_23881,N_19694,N_15342);
or U23882 (N_23882,N_17879,N_17800);
nor U23883 (N_23883,N_18981,N_15865);
or U23884 (N_23884,N_16041,N_19827);
and U23885 (N_23885,N_18472,N_18894);
nor U23886 (N_23886,N_17919,N_19022);
nand U23887 (N_23887,N_18276,N_17207);
nand U23888 (N_23888,N_16615,N_17438);
and U23889 (N_23889,N_17757,N_18343);
or U23890 (N_23890,N_15979,N_16057);
nand U23891 (N_23891,N_15896,N_17645);
nor U23892 (N_23892,N_18026,N_17438);
nand U23893 (N_23893,N_18953,N_19086);
and U23894 (N_23894,N_16184,N_18033);
or U23895 (N_23895,N_17017,N_19107);
nand U23896 (N_23896,N_19346,N_18098);
or U23897 (N_23897,N_16421,N_16456);
or U23898 (N_23898,N_17778,N_19725);
nand U23899 (N_23899,N_17387,N_17124);
nor U23900 (N_23900,N_15834,N_15480);
and U23901 (N_23901,N_19088,N_16900);
nor U23902 (N_23902,N_18481,N_19753);
nand U23903 (N_23903,N_16419,N_17758);
and U23904 (N_23904,N_15104,N_16128);
nand U23905 (N_23905,N_16716,N_16967);
nor U23906 (N_23906,N_15409,N_17347);
and U23907 (N_23907,N_18083,N_16731);
nand U23908 (N_23908,N_15240,N_18501);
or U23909 (N_23909,N_16456,N_19426);
and U23910 (N_23910,N_18812,N_16156);
xor U23911 (N_23911,N_18567,N_17548);
nand U23912 (N_23912,N_18783,N_18223);
or U23913 (N_23913,N_17903,N_19528);
and U23914 (N_23914,N_16761,N_16497);
nand U23915 (N_23915,N_18101,N_19780);
nor U23916 (N_23916,N_17052,N_17122);
nor U23917 (N_23917,N_19051,N_17416);
nor U23918 (N_23918,N_19377,N_19131);
and U23919 (N_23919,N_18644,N_16063);
and U23920 (N_23920,N_16081,N_19183);
or U23921 (N_23921,N_17567,N_17401);
nor U23922 (N_23922,N_16890,N_15121);
xor U23923 (N_23923,N_17008,N_16590);
or U23924 (N_23924,N_16928,N_16850);
nor U23925 (N_23925,N_19628,N_19456);
and U23926 (N_23926,N_16507,N_18505);
nor U23927 (N_23927,N_18324,N_19487);
and U23928 (N_23928,N_15157,N_15341);
nor U23929 (N_23929,N_19695,N_16019);
and U23930 (N_23930,N_18701,N_15090);
xor U23931 (N_23931,N_15337,N_17150);
and U23932 (N_23932,N_19610,N_15302);
and U23933 (N_23933,N_19724,N_18831);
nand U23934 (N_23934,N_15561,N_17765);
xor U23935 (N_23935,N_17097,N_15786);
nand U23936 (N_23936,N_18724,N_17790);
nor U23937 (N_23937,N_16414,N_19273);
and U23938 (N_23938,N_18434,N_16634);
nand U23939 (N_23939,N_16209,N_17017);
nor U23940 (N_23940,N_17251,N_17738);
nor U23941 (N_23941,N_18054,N_15048);
or U23942 (N_23942,N_19299,N_18697);
nor U23943 (N_23943,N_19416,N_15312);
and U23944 (N_23944,N_18716,N_16147);
or U23945 (N_23945,N_15556,N_19631);
nand U23946 (N_23946,N_15232,N_19586);
xor U23947 (N_23947,N_17876,N_17316);
and U23948 (N_23948,N_19418,N_18170);
nor U23949 (N_23949,N_15413,N_17298);
nor U23950 (N_23950,N_19995,N_16072);
or U23951 (N_23951,N_16508,N_17134);
nor U23952 (N_23952,N_18726,N_19479);
or U23953 (N_23953,N_17137,N_17453);
and U23954 (N_23954,N_16116,N_19325);
nand U23955 (N_23955,N_15978,N_18348);
nand U23956 (N_23956,N_17280,N_17790);
or U23957 (N_23957,N_16467,N_19766);
nor U23958 (N_23958,N_19247,N_18851);
nand U23959 (N_23959,N_15127,N_17021);
or U23960 (N_23960,N_15812,N_18568);
xor U23961 (N_23961,N_15959,N_16414);
and U23962 (N_23962,N_15779,N_18486);
and U23963 (N_23963,N_16943,N_19284);
nand U23964 (N_23964,N_18463,N_18121);
nor U23965 (N_23965,N_17083,N_16982);
xor U23966 (N_23966,N_16509,N_17096);
nor U23967 (N_23967,N_17255,N_15735);
xor U23968 (N_23968,N_16847,N_18898);
nand U23969 (N_23969,N_15014,N_16140);
xor U23970 (N_23970,N_18215,N_15708);
and U23971 (N_23971,N_17426,N_19127);
or U23972 (N_23972,N_18132,N_17909);
xor U23973 (N_23973,N_15469,N_16070);
or U23974 (N_23974,N_16515,N_15344);
and U23975 (N_23975,N_18481,N_18492);
or U23976 (N_23976,N_16870,N_15485);
and U23977 (N_23977,N_19597,N_15451);
nand U23978 (N_23978,N_19658,N_17402);
and U23979 (N_23979,N_19657,N_16594);
nand U23980 (N_23980,N_17235,N_15516);
and U23981 (N_23981,N_18972,N_18091);
or U23982 (N_23982,N_17319,N_16199);
and U23983 (N_23983,N_17544,N_19968);
nand U23984 (N_23984,N_15743,N_15343);
nor U23985 (N_23985,N_15062,N_16851);
nand U23986 (N_23986,N_18546,N_16230);
and U23987 (N_23987,N_17719,N_19798);
or U23988 (N_23988,N_15667,N_17779);
and U23989 (N_23989,N_18554,N_15320);
nor U23990 (N_23990,N_16109,N_18896);
and U23991 (N_23991,N_16880,N_16151);
or U23992 (N_23992,N_16059,N_15496);
nand U23993 (N_23993,N_19861,N_19725);
and U23994 (N_23994,N_15379,N_17309);
nand U23995 (N_23995,N_15891,N_17041);
nor U23996 (N_23996,N_18740,N_15664);
and U23997 (N_23997,N_18060,N_19328);
and U23998 (N_23998,N_16607,N_18687);
nor U23999 (N_23999,N_19001,N_17643);
nor U24000 (N_24000,N_18003,N_17708);
and U24001 (N_24001,N_16684,N_17301);
nand U24002 (N_24002,N_17295,N_19382);
nand U24003 (N_24003,N_18141,N_18441);
and U24004 (N_24004,N_17972,N_15228);
nand U24005 (N_24005,N_17905,N_15296);
or U24006 (N_24006,N_19683,N_19179);
and U24007 (N_24007,N_16109,N_18172);
or U24008 (N_24008,N_15613,N_17990);
xnor U24009 (N_24009,N_18663,N_19049);
and U24010 (N_24010,N_19565,N_18120);
and U24011 (N_24011,N_19774,N_16011);
nand U24012 (N_24012,N_16124,N_15853);
and U24013 (N_24013,N_19351,N_19532);
nor U24014 (N_24014,N_16533,N_17489);
or U24015 (N_24015,N_15845,N_18847);
or U24016 (N_24016,N_17325,N_16710);
nand U24017 (N_24017,N_19368,N_16688);
or U24018 (N_24018,N_19074,N_15548);
and U24019 (N_24019,N_15764,N_16953);
and U24020 (N_24020,N_16394,N_19420);
and U24021 (N_24021,N_16890,N_18889);
nor U24022 (N_24022,N_16672,N_18803);
nand U24023 (N_24023,N_17432,N_18324);
and U24024 (N_24024,N_19542,N_15757);
nand U24025 (N_24025,N_18566,N_15177);
xnor U24026 (N_24026,N_19777,N_18077);
nor U24027 (N_24027,N_18088,N_16387);
nand U24028 (N_24028,N_19732,N_19209);
nor U24029 (N_24029,N_18775,N_19871);
nor U24030 (N_24030,N_18592,N_18297);
nand U24031 (N_24031,N_16355,N_17174);
nor U24032 (N_24032,N_18753,N_18788);
nand U24033 (N_24033,N_17584,N_19308);
xor U24034 (N_24034,N_19264,N_17544);
nand U24035 (N_24035,N_17514,N_15011);
nor U24036 (N_24036,N_17043,N_18566);
and U24037 (N_24037,N_16041,N_19685);
nand U24038 (N_24038,N_16134,N_15075);
xnor U24039 (N_24039,N_16437,N_17812);
nand U24040 (N_24040,N_17228,N_16331);
nand U24041 (N_24041,N_16639,N_16882);
nand U24042 (N_24042,N_19508,N_17902);
and U24043 (N_24043,N_18251,N_16115);
and U24044 (N_24044,N_15973,N_17011);
nor U24045 (N_24045,N_18790,N_15370);
nand U24046 (N_24046,N_17273,N_16520);
and U24047 (N_24047,N_15557,N_17586);
or U24048 (N_24048,N_15034,N_16061);
xor U24049 (N_24049,N_17023,N_18657);
nand U24050 (N_24050,N_18834,N_16886);
and U24051 (N_24051,N_16062,N_19682);
or U24052 (N_24052,N_17690,N_16173);
nor U24053 (N_24053,N_15186,N_15970);
nor U24054 (N_24054,N_17428,N_15446);
and U24055 (N_24055,N_19459,N_15435);
nand U24056 (N_24056,N_17167,N_18653);
nand U24057 (N_24057,N_17561,N_16041);
and U24058 (N_24058,N_18485,N_18747);
nor U24059 (N_24059,N_19382,N_18814);
or U24060 (N_24060,N_17707,N_16622);
and U24061 (N_24061,N_16903,N_19470);
nor U24062 (N_24062,N_17319,N_19410);
and U24063 (N_24063,N_18635,N_17361);
or U24064 (N_24064,N_15674,N_18206);
nor U24065 (N_24065,N_19536,N_16836);
nor U24066 (N_24066,N_18802,N_15355);
nor U24067 (N_24067,N_15661,N_15672);
or U24068 (N_24068,N_16231,N_17241);
nor U24069 (N_24069,N_15139,N_18053);
and U24070 (N_24070,N_19778,N_17508);
or U24071 (N_24071,N_19107,N_16139);
nor U24072 (N_24072,N_17638,N_15007);
and U24073 (N_24073,N_16994,N_19432);
nand U24074 (N_24074,N_16001,N_15439);
nand U24075 (N_24075,N_16776,N_15544);
and U24076 (N_24076,N_15063,N_16100);
nand U24077 (N_24077,N_16937,N_19337);
or U24078 (N_24078,N_16424,N_19798);
and U24079 (N_24079,N_19093,N_16903);
and U24080 (N_24080,N_16948,N_15443);
nand U24081 (N_24081,N_19630,N_17929);
nor U24082 (N_24082,N_19544,N_16801);
and U24083 (N_24083,N_18120,N_17046);
xor U24084 (N_24084,N_17109,N_16042);
and U24085 (N_24085,N_18466,N_15893);
and U24086 (N_24086,N_17594,N_18143);
or U24087 (N_24087,N_16484,N_15423);
nor U24088 (N_24088,N_19520,N_17819);
or U24089 (N_24089,N_16444,N_18960);
nand U24090 (N_24090,N_16871,N_15775);
nand U24091 (N_24091,N_15741,N_16675);
or U24092 (N_24092,N_15052,N_19546);
or U24093 (N_24093,N_15932,N_16807);
and U24094 (N_24094,N_17616,N_18228);
nand U24095 (N_24095,N_18920,N_16321);
and U24096 (N_24096,N_18256,N_15183);
and U24097 (N_24097,N_16312,N_16898);
nor U24098 (N_24098,N_15834,N_17365);
nand U24099 (N_24099,N_15623,N_19202);
nor U24100 (N_24100,N_17113,N_16221);
nor U24101 (N_24101,N_16152,N_15004);
or U24102 (N_24102,N_15002,N_16473);
xor U24103 (N_24103,N_16960,N_17254);
nor U24104 (N_24104,N_19749,N_19743);
nor U24105 (N_24105,N_18501,N_15454);
xor U24106 (N_24106,N_15720,N_18183);
or U24107 (N_24107,N_17359,N_15363);
or U24108 (N_24108,N_15722,N_15958);
nand U24109 (N_24109,N_19953,N_17319);
nand U24110 (N_24110,N_19843,N_17274);
nor U24111 (N_24111,N_19970,N_15908);
and U24112 (N_24112,N_17053,N_16697);
or U24113 (N_24113,N_16542,N_17589);
and U24114 (N_24114,N_17422,N_19500);
xor U24115 (N_24115,N_18851,N_17531);
or U24116 (N_24116,N_16221,N_17979);
nor U24117 (N_24117,N_16962,N_16543);
nand U24118 (N_24118,N_15876,N_17230);
or U24119 (N_24119,N_16137,N_18884);
and U24120 (N_24120,N_15846,N_17738);
and U24121 (N_24121,N_19379,N_16408);
nor U24122 (N_24122,N_17419,N_16300);
or U24123 (N_24123,N_19118,N_16614);
nand U24124 (N_24124,N_17158,N_18754);
and U24125 (N_24125,N_16178,N_17007);
or U24126 (N_24126,N_16679,N_19760);
or U24127 (N_24127,N_17376,N_15937);
nand U24128 (N_24128,N_17888,N_15549);
nand U24129 (N_24129,N_18101,N_19448);
or U24130 (N_24130,N_16519,N_15261);
and U24131 (N_24131,N_16711,N_18513);
nor U24132 (N_24132,N_17196,N_15943);
nor U24133 (N_24133,N_16341,N_16045);
nor U24134 (N_24134,N_18199,N_16662);
or U24135 (N_24135,N_19638,N_16233);
nor U24136 (N_24136,N_15687,N_17544);
and U24137 (N_24137,N_18709,N_17123);
nor U24138 (N_24138,N_19080,N_15775);
nor U24139 (N_24139,N_18192,N_18541);
nand U24140 (N_24140,N_18239,N_19172);
and U24141 (N_24141,N_18993,N_17725);
nor U24142 (N_24142,N_15690,N_19301);
or U24143 (N_24143,N_15441,N_15377);
nor U24144 (N_24144,N_19055,N_17604);
or U24145 (N_24145,N_17497,N_16028);
nor U24146 (N_24146,N_18468,N_18080);
and U24147 (N_24147,N_15723,N_18519);
or U24148 (N_24148,N_15476,N_17814);
nand U24149 (N_24149,N_16348,N_17331);
nor U24150 (N_24150,N_15913,N_17958);
or U24151 (N_24151,N_15265,N_16190);
nand U24152 (N_24152,N_17518,N_16550);
nand U24153 (N_24153,N_16080,N_16372);
and U24154 (N_24154,N_16742,N_17440);
or U24155 (N_24155,N_19718,N_18922);
and U24156 (N_24156,N_15906,N_18626);
and U24157 (N_24157,N_15339,N_19737);
nor U24158 (N_24158,N_15137,N_17125);
nor U24159 (N_24159,N_15603,N_16909);
nand U24160 (N_24160,N_17003,N_17546);
or U24161 (N_24161,N_15850,N_18853);
and U24162 (N_24162,N_16627,N_18398);
or U24163 (N_24163,N_19438,N_15091);
nor U24164 (N_24164,N_19019,N_17458);
nor U24165 (N_24165,N_17030,N_18604);
nor U24166 (N_24166,N_15315,N_15323);
nor U24167 (N_24167,N_15349,N_17306);
and U24168 (N_24168,N_19912,N_16956);
or U24169 (N_24169,N_19243,N_18389);
and U24170 (N_24170,N_19756,N_15093);
or U24171 (N_24171,N_18883,N_17887);
nor U24172 (N_24172,N_17567,N_15627);
nor U24173 (N_24173,N_18074,N_17606);
nand U24174 (N_24174,N_15242,N_16264);
or U24175 (N_24175,N_15020,N_15380);
and U24176 (N_24176,N_18710,N_16884);
nand U24177 (N_24177,N_17101,N_15204);
xnor U24178 (N_24178,N_17498,N_19721);
nand U24179 (N_24179,N_16730,N_15661);
or U24180 (N_24180,N_17041,N_15356);
nor U24181 (N_24181,N_19182,N_15312);
nand U24182 (N_24182,N_18542,N_16096);
nand U24183 (N_24183,N_17441,N_18619);
or U24184 (N_24184,N_18406,N_19572);
or U24185 (N_24185,N_18711,N_17724);
xor U24186 (N_24186,N_17053,N_17587);
or U24187 (N_24187,N_19551,N_19559);
and U24188 (N_24188,N_19646,N_19614);
and U24189 (N_24189,N_18753,N_18968);
or U24190 (N_24190,N_16390,N_18203);
or U24191 (N_24191,N_16218,N_19465);
nand U24192 (N_24192,N_15731,N_18786);
or U24193 (N_24193,N_19625,N_18487);
xnor U24194 (N_24194,N_19105,N_16488);
xnor U24195 (N_24195,N_15997,N_17553);
and U24196 (N_24196,N_16332,N_19637);
and U24197 (N_24197,N_16972,N_15310);
xnor U24198 (N_24198,N_18427,N_16570);
and U24199 (N_24199,N_18877,N_15660);
and U24200 (N_24200,N_18484,N_17453);
nor U24201 (N_24201,N_17478,N_17396);
nor U24202 (N_24202,N_16591,N_19939);
nand U24203 (N_24203,N_18935,N_16976);
nand U24204 (N_24204,N_16429,N_15660);
nor U24205 (N_24205,N_18247,N_15192);
xor U24206 (N_24206,N_15712,N_15176);
and U24207 (N_24207,N_16477,N_19611);
nor U24208 (N_24208,N_19739,N_18830);
and U24209 (N_24209,N_16899,N_19837);
nor U24210 (N_24210,N_19266,N_17709);
nand U24211 (N_24211,N_18127,N_17171);
and U24212 (N_24212,N_15630,N_15791);
nand U24213 (N_24213,N_19600,N_15606);
nor U24214 (N_24214,N_16232,N_19774);
and U24215 (N_24215,N_19110,N_19398);
or U24216 (N_24216,N_18623,N_15442);
and U24217 (N_24217,N_19603,N_17408);
nor U24218 (N_24218,N_17333,N_15485);
nand U24219 (N_24219,N_18780,N_19559);
xor U24220 (N_24220,N_18543,N_17354);
nor U24221 (N_24221,N_17796,N_15750);
xnor U24222 (N_24222,N_18404,N_17134);
or U24223 (N_24223,N_16239,N_19140);
or U24224 (N_24224,N_15698,N_19859);
nor U24225 (N_24225,N_17772,N_16514);
xnor U24226 (N_24226,N_19266,N_18001);
or U24227 (N_24227,N_15937,N_17789);
or U24228 (N_24228,N_18256,N_17636);
nand U24229 (N_24229,N_15081,N_19803);
nor U24230 (N_24230,N_18914,N_18395);
nor U24231 (N_24231,N_17362,N_15508);
nand U24232 (N_24232,N_17249,N_16799);
and U24233 (N_24233,N_17152,N_17870);
and U24234 (N_24234,N_15575,N_17808);
nor U24235 (N_24235,N_18680,N_16725);
nand U24236 (N_24236,N_15355,N_15094);
and U24237 (N_24237,N_18250,N_15024);
or U24238 (N_24238,N_16129,N_19653);
or U24239 (N_24239,N_16390,N_15892);
or U24240 (N_24240,N_16998,N_15272);
and U24241 (N_24241,N_16809,N_16600);
or U24242 (N_24242,N_15216,N_16171);
nand U24243 (N_24243,N_17328,N_16549);
nor U24244 (N_24244,N_17545,N_17061);
or U24245 (N_24245,N_17288,N_15908);
nand U24246 (N_24246,N_15145,N_15639);
nand U24247 (N_24247,N_18512,N_15114);
or U24248 (N_24248,N_18809,N_18332);
nor U24249 (N_24249,N_17056,N_17856);
and U24250 (N_24250,N_17568,N_16353);
nand U24251 (N_24251,N_16093,N_17136);
or U24252 (N_24252,N_15897,N_15006);
nand U24253 (N_24253,N_19964,N_17078);
or U24254 (N_24254,N_18010,N_16533);
nor U24255 (N_24255,N_16783,N_16316);
or U24256 (N_24256,N_16646,N_18328);
or U24257 (N_24257,N_17109,N_15808);
xor U24258 (N_24258,N_18375,N_19845);
nor U24259 (N_24259,N_19234,N_17852);
and U24260 (N_24260,N_16758,N_17187);
xnor U24261 (N_24261,N_18580,N_16447);
xor U24262 (N_24262,N_17597,N_17716);
or U24263 (N_24263,N_17075,N_19417);
or U24264 (N_24264,N_17740,N_19520);
nor U24265 (N_24265,N_18584,N_18716);
xnor U24266 (N_24266,N_15201,N_16384);
and U24267 (N_24267,N_17744,N_18268);
and U24268 (N_24268,N_17445,N_19614);
or U24269 (N_24269,N_18663,N_18611);
nand U24270 (N_24270,N_15521,N_15589);
xnor U24271 (N_24271,N_16103,N_16533);
and U24272 (N_24272,N_16940,N_16902);
or U24273 (N_24273,N_16254,N_18867);
or U24274 (N_24274,N_18417,N_16728);
nand U24275 (N_24275,N_15853,N_19808);
or U24276 (N_24276,N_17839,N_18529);
or U24277 (N_24277,N_18653,N_17414);
nor U24278 (N_24278,N_19689,N_19082);
and U24279 (N_24279,N_19458,N_19286);
nor U24280 (N_24280,N_16844,N_19235);
nand U24281 (N_24281,N_19655,N_19583);
nand U24282 (N_24282,N_18945,N_16798);
nor U24283 (N_24283,N_18403,N_16251);
or U24284 (N_24284,N_16089,N_16944);
or U24285 (N_24285,N_18162,N_18720);
or U24286 (N_24286,N_16118,N_19333);
nor U24287 (N_24287,N_16565,N_15610);
xor U24288 (N_24288,N_17368,N_17938);
and U24289 (N_24289,N_15450,N_15062);
xnor U24290 (N_24290,N_18050,N_16790);
and U24291 (N_24291,N_19207,N_15671);
and U24292 (N_24292,N_17888,N_16340);
nor U24293 (N_24293,N_19911,N_19847);
or U24294 (N_24294,N_19398,N_19010);
nor U24295 (N_24295,N_18113,N_17279);
nand U24296 (N_24296,N_19389,N_16249);
xor U24297 (N_24297,N_16408,N_19667);
or U24298 (N_24298,N_18025,N_16125);
or U24299 (N_24299,N_17943,N_18235);
or U24300 (N_24300,N_16729,N_18092);
nor U24301 (N_24301,N_19316,N_16449);
nand U24302 (N_24302,N_16573,N_15726);
or U24303 (N_24303,N_17926,N_18906);
and U24304 (N_24304,N_15825,N_15637);
nand U24305 (N_24305,N_19639,N_19715);
nand U24306 (N_24306,N_18714,N_17049);
and U24307 (N_24307,N_19456,N_19153);
and U24308 (N_24308,N_18583,N_19707);
nand U24309 (N_24309,N_15171,N_17516);
or U24310 (N_24310,N_19064,N_17107);
nand U24311 (N_24311,N_18214,N_16296);
nand U24312 (N_24312,N_18920,N_16964);
nor U24313 (N_24313,N_16562,N_16138);
nand U24314 (N_24314,N_15275,N_15272);
nand U24315 (N_24315,N_17646,N_19863);
or U24316 (N_24316,N_15668,N_16671);
nor U24317 (N_24317,N_16733,N_15908);
or U24318 (N_24318,N_16550,N_17018);
and U24319 (N_24319,N_17211,N_15121);
nor U24320 (N_24320,N_18120,N_16885);
and U24321 (N_24321,N_18628,N_17156);
or U24322 (N_24322,N_16497,N_18096);
and U24323 (N_24323,N_16103,N_15206);
nand U24324 (N_24324,N_15209,N_16285);
or U24325 (N_24325,N_19815,N_15194);
or U24326 (N_24326,N_17072,N_19643);
and U24327 (N_24327,N_17321,N_17843);
nor U24328 (N_24328,N_19857,N_18505);
xnor U24329 (N_24329,N_15761,N_18008);
nand U24330 (N_24330,N_16072,N_19021);
or U24331 (N_24331,N_16115,N_15618);
and U24332 (N_24332,N_16226,N_15658);
or U24333 (N_24333,N_17857,N_18858);
or U24334 (N_24334,N_19987,N_17990);
nand U24335 (N_24335,N_16943,N_17782);
nor U24336 (N_24336,N_15958,N_15079);
nor U24337 (N_24337,N_19262,N_18704);
nand U24338 (N_24338,N_17556,N_16099);
and U24339 (N_24339,N_19956,N_17666);
or U24340 (N_24340,N_16420,N_19030);
nand U24341 (N_24341,N_16091,N_15265);
nor U24342 (N_24342,N_17952,N_15187);
nand U24343 (N_24343,N_17947,N_15178);
nor U24344 (N_24344,N_18104,N_18440);
and U24345 (N_24345,N_19939,N_15421);
or U24346 (N_24346,N_18410,N_18309);
nand U24347 (N_24347,N_19782,N_15419);
and U24348 (N_24348,N_18992,N_15018);
and U24349 (N_24349,N_19838,N_18710);
nand U24350 (N_24350,N_16296,N_19830);
nand U24351 (N_24351,N_18720,N_15542);
or U24352 (N_24352,N_15816,N_18477);
xnor U24353 (N_24353,N_16331,N_16475);
or U24354 (N_24354,N_17926,N_16729);
xor U24355 (N_24355,N_18953,N_15465);
nand U24356 (N_24356,N_17988,N_19755);
nor U24357 (N_24357,N_19693,N_19969);
and U24358 (N_24358,N_16822,N_19049);
nor U24359 (N_24359,N_19100,N_18776);
nand U24360 (N_24360,N_18661,N_16299);
nor U24361 (N_24361,N_18988,N_19621);
or U24362 (N_24362,N_15489,N_15647);
or U24363 (N_24363,N_17594,N_19506);
nor U24364 (N_24364,N_17073,N_19915);
nand U24365 (N_24365,N_18429,N_19234);
or U24366 (N_24366,N_15615,N_17024);
nand U24367 (N_24367,N_15582,N_15924);
or U24368 (N_24368,N_18624,N_15335);
nand U24369 (N_24369,N_16199,N_19641);
nand U24370 (N_24370,N_15120,N_18328);
nor U24371 (N_24371,N_17369,N_15202);
xor U24372 (N_24372,N_18707,N_15657);
nor U24373 (N_24373,N_17185,N_15967);
or U24374 (N_24374,N_15990,N_19664);
nor U24375 (N_24375,N_17578,N_16976);
nand U24376 (N_24376,N_19570,N_19842);
and U24377 (N_24377,N_19778,N_17325);
nand U24378 (N_24378,N_19064,N_16426);
and U24379 (N_24379,N_19225,N_18031);
and U24380 (N_24380,N_17618,N_16193);
or U24381 (N_24381,N_19638,N_18008);
nor U24382 (N_24382,N_15503,N_19508);
nand U24383 (N_24383,N_18969,N_17414);
and U24384 (N_24384,N_19069,N_18295);
nor U24385 (N_24385,N_15117,N_16690);
and U24386 (N_24386,N_18432,N_15286);
nor U24387 (N_24387,N_19148,N_19249);
nand U24388 (N_24388,N_19716,N_15418);
nand U24389 (N_24389,N_19262,N_17437);
or U24390 (N_24390,N_19644,N_17715);
nor U24391 (N_24391,N_15457,N_16184);
and U24392 (N_24392,N_19426,N_19978);
and U24393 (N_24393,N_16875,N_18354);
xnor U24394 (N_24394,N_17052,N_17266);
nand U24395 (N_24395,N_15501,N_17467);
nand U24396 (N_24396,N_16061,N_19570);
nor U24397 (N_24397,N_17624,N_19788);
or U24398 (N_24398,N_19623,N_17774);
nor U24399 (N_24399,N_18610,N_18447);
or U24400 (N_24400,N_18614,N_15596);
nand U24401 (N_24401,N_18753,N_19477);
or U24402 (N_24402,N_16808,N_19158);
or U24403 (N_24403,N_15108,N_18098);
nor U24404 (N_24404,N_17337,N_17808);
nor U24405 (N_24405,N_19737,N_17859);
or U24406 (N_24406,N_19064,N_17256);
or U24407 (N_24407,N_15439,N_19630);
and U24408 (N_24408,N_17009,N_16678);
nor U24409 (N_24409,N_19421,N_17839);
or U24410 (N_24410,N_19556,N_18289);
or U24411 (N_24411,N_18968,N_17500);
nand U24412 (N_24412,N_16658,N_17985);
or U24413 (N_24413,N_15816,N_18270);
or U24414 (N_24414,N_17379,N_18435);
and U24415 (N_24415,N_19828,N_17302);
or U24416 (N_24416,N_18484,N_15209);
and U24417 (N_24417,N_16612,N_19389);
nor U24418 (N_24418,N_18281,N_19913);
xor U24419 (N_24419,N_18930,N_19327);
and U24420 (N_24420,N_15138,N_18575);
xnor U24421 (N_24421,N_16411,N_15829);
nor U24422 (N_24422,N_19217,N_19089);
nor U24423 (N_24423,N_15339,N_18295);
nand U24424 (N_24424,N_16363,N_18263);
and U24425 (N_24425,N_15226,N_16085);
or U24426 (N_24426,N_15712,N_17701);
and U24427 (N_24427,N_17277,N_17833);
and U24428 (N_24428,N_18712,N_17917);
and U24429 (N_24429,N_16719,N_16154);
nand U24430 (N_24430,N_18034,N_16483);
or U24431 (N_24431,N_15998,N_17024);
nor U24432 (N_24432,N_19346,N_15955);
nand U24433 (N_24433,N_16054,N_17176);
or U24434 (N_24434,N_19872,N_17521);
nor U24435 (N_24435,N_18655,N_15446);
nor U24436 (N_24436,N_16147,N_16994);
nor U24437 (N_24437,N_15989,N_16589);
nor U24438 (N_24438,N_18480,N_16759);
and U24439 (N_24439,N_15564,N_17975);
nand U24440 (N_24440,N_19077,N_19425);
nand U24441 (N_24441,N_18976,N_19759);
nand U24442 (N_24442,N_17296,N_19977);
nand U24443 (N_24443,N_15732,N_17043);
nand U24444 (N_24444,N_19012,N_19022);
xor U24445 (N_24445,N_18743,N_18088);
or U24446 (N_24446,N_15229,N_19703);
or U24447 (N_24447,N_17352,N_17527);
nor U24448 (N_24448,N_17804,N_18415);
nand U24449 (N_24449,N_17490,N_16522);
and U24450 (N_24450,N_18213,N_16702);
nor U24451 (N_24451,N_17303,N_16771);
or U24452 (N_24452,N_19555,N_17894);
nor U24453 (N_24453,N_16194,N_15181);
nor U24454 (N_24454,N_19781,N_16487);
or U24455 (N_24455,N_15945,N_16648);
nand U24456 (N_24456,N_19642,N_15513);
nand U24457 (N_24457,N_16471,N_15108);
and U24458 (N_24458,N_17005,N_19664);
or U24459 (N_24459,N_18705,N_15957);
and U24460 (N_24460,N_15914,N_18343);
or U24461 (N_24461,N_15208,N_19223);
nor U24462 (N_24462,N_19736,N_17478);
or U24463 (N_24463,N_17846,N_19167);
nand U24464 (N_24464,N_15724,N_18221);
nor U24465 (N_24465,N_17265,N_17807);
nand U24466 (N_24466,N_17320,N_16445);
or U24467 (N_24467,N_17204,N_17920);
nand U24468 (N_24468,N_19997,N_16197);
nand U24469 (N_24469,N_19566,N_17255);
or U24470 (N_24470,N_15000,N_15041);
and U24471 (N_24471,N_15867,N_18513);
xnor U24472 (N_24472,N_17896,N_17927);
xnor U24473 (N_24473,N_17823,N_16980);
nand U24474 (N_24474,N_18001,N_15550);
xor U24475 (N_24475,N_18179,N_17352);
or U24476 (N_24476,N_17085,N_19475);
or U24477 (N_24477,N_17698,N_17634);
or U24478 (N_24478,N_15018,N_16588);
nor U24479 (N_24479,N_18743,N_19834);
nor U24480 (N_24480,N_18369,N_15015);
xnor U24481 (N_24481,N_16054,N_18642);
nor U24482 (N_24482,N_15353,N_17476);
nand U24483 (N_24483,N_15462,N_18359);
or U24484 (N_24484,N_15410,N_17279);
nand U24485 (N_24485,N_17615,N_15452);
or U24486 (N_24486,N_16489,N_18977);
nor U24487 (N_24487,N_16577,N_19202);
and U24488 (N_24488,N_18955,N_18835);
nand U24489 (N_24489,N_18817,N_17435);
and U24490 (N_24490,N_19587,N_15078);
nor U24491 (N_24491,N_19893,N_17876);
or U24492 (N_24492,N_15438,N_15800);
nand U24493 (N_24493,N_15315,N_19768);
nor U24494 (N_24494,N_15425,N_19603);
or U24495 (N_24495,N_17961,N_18225);
and U24496 (N_24496,N_15745,N_15601);
nor U24497 (N_24497,N_15551,N_16253);
or U24498 (N_24498,N_15497,N_16905);
nand U24499 (N_24499,N_19107,N_17606);
and U24500 (N_24500,N_15748,N_18288);
or U24501 (N_24501,N_17667,N_15889);
and U24502 (N_24502,N_16667,N_16075);
nor U24503 (N_24503,N_17809,N_15818);
or U24504 (N_24504,N_18844,N_15278);
nand U24505 (N_24505,N_16594,N_17242);
nand U24506 (N_24506,N_18219,N_18180);
or U24507 (N_24507,N_15661,N_19157);
xnor U24508 (N_24508,N_18242,N_15875);
and U24509 (N_24509,N_18243,N_17360);
and U24510 (N_24510,N_16973,N_17738);
and U24511 (N_24511,N_18284,N_18938);
nor U24512 (N_24512,N_18522,N_17160);
or U24513 (N_24513,N_19337,N_18029);
nand U24514 (N_24514,N_15615,N_19649);
or U24515 (N_24515,N_18634,N_16791);
nor U24516 (N_24516,N_15357,N_19301);
or U24517 (N_24517,N_17218,N_17611);
nor U24518 (N_24518,N_17407,N_18455);
and U24519 (N_24519,N_19965,N_15652);
or U24520 (N_24520,N_15920,N_15784);
and U24521 (N_24521,N_19027,N_19119);
and U24522 (N_24522,N_17986,N_16947);
nand U24523 (N_24523,N_16723,N_18799);
nand U24524 (N_24524,N_16909,N_16103);
nand U24525 (N_24525,N_18200,N_15156);
or U24526 (N_24526,N_17526,N_16505);
nand U24527 (N_24527,N_15209,N_15336);
nor U24528 (N_24528,N_19384,N_18858);
and U24529 (N_24529,N_17769,N_19721);
and U24530 (N_24530,N_17089,N_18837);
and U24531 (N_24531,N_15941,N_18272);
nor U24532 (N_24532,N_15539,N_15581);
and U24533 (N_24533,N_18384,N_15309);
xor U24534 (N_24534,N_15666,N_17127);
nand U24535 (N_24535,N_18314,N_15019);
and U24536 (N_24536,N_19865,N_15718);
and U24537 (N_24537,N_19545,N_16049);
nor U24538 (N_24538,N_19721,N_19841);
and U24539 (N_24539,N_18249,N_18312);
or U24540 (N_24540,N_16047,N_17235);
or U24541 (N_24541,N_17293,N_18097);
nor U24542 (N_24542,N_15401,N_17499);
nand U24543 (N_24543,N_17487,N_18535);
or U24544 (N_24544,N_18237,N_15477);
or U24545 (N_24545,N_16006,N_18813);
nand U24546 (N_24546,N_16001,N_19266);
or U24547 (N_24547,N_16370,N_17320);
nand U24548 (N_24548,N_17331,N_15172);
nand U24549 (N_24549,N_18282,N_19325);
nand U24550 (N_24550,N_18517,N_16773);
or U24551 (N_24551,N_17774,N_17704);
xor U24552 (N_24552,N_16681,N_16601);
nand U24553 (N_24553,N_16195,N_18671);
or U24554 (N_24554,N_18797,N_15469);
nor U24555 (N_24555,N_18811,N_19186);
or U24556 (N_24556,N_17969,N_18921);
or U24557 (N_24557,N_17653,N_19245);
xnor U24558 (N_24558,N_17565,N_17343);
nor U24559 (N_24559,N_16945,N_19166);
or U24560 (N_24560,N_15406,N_19970);
nor U24561 (N_24561,N_16198,N_15117);
nor U24562 (N_24562,N_15233,N_15892);
nor U24563 (N_24563,N_17853,N_19877);
and U24564 (N_24564,N_17473,N_19026);
nor U24565 (N_24565,N_19505,N_15473);
and U24566 (N_24566,N_19026,N_15656);
nand U24567 (N_24567,N_17924,N_18152);
and U24568 (N_24568,N_19633,N_18522);
or U24569 (N_24569,N_18180,N_19696);
and U24570 (N_24570,N_19368,N_17443);
nand U24571 (N_24571,N_19461,N_18954);
or U24572 (N_24572,N_16710,N_16679);
and U24573 (N_24573,N_19867,N_16268);
and U24574 (N_24574,N_15460,N_17921);
or U24575 (N_24575,N_15605,N_17174);
xor U24576 (N_24576,N_17480,N_18474);
nand U24577 (N_24577,N_15061,N_17075);
or U24578 (N_24578,N_15451,N_19742);
or U24579 (N_24579,N_19965,N_16300);
or U24580 (N_24580,N_15455,N_17728);
or U24581 (N_24581,N_18994,N_17237);
nand U24582 (N_24582,N_16860,N_16093);
and U24583 (N_24583,N_18619,N_16509);
and U24584 (N_24584,N_15249,N_19740);
or U24585 (N_24585,N_18885,N_18388);
nor U24586 (N_24586,N_19023,N_18250);
nand U24587 (N_24587,N_17363,N_15382);
nor U24588 (N_24588,N_15927,N_16208);
xnor U24589 (N_24589,N_16083,N_18697);
xnor U24590 (N_24590,N_17854,N_17644);
or U24591 (N_24591,N_17163,N_16184);
nand U24592 (N_24592,N_18095,N_18189);
or U24593 (N_24593,N_19922,N_17410);
or U24594 (N_24594,N_15637,N_19225);
nor U24595 (N_24595,N_17661,N_18853);
nand U24596 (N_24596,N_17394,N_15337);
nor U24597 (N_24597,N_15524,N_18762);
and U24598 (N_24598,N_15743,N_15787);
or U24599 (N_24599,N_16648,N_18893);
nor U24600 (N_24600,N_17814,N_16778);
xor U24601 (N_24601,N_19816,N_19636);
or U24602 (N_24602,N_15132,N_16017);
nand U24603 (N_24603,N_15801,N_18921);
xnor U24604 (N_24604,N_18324,N_18830);
or U24605 (N_24605,N_15476,N_17711);
and U24606 (N_24606,N_17147,N_15306);
or U24607 (N_24607,N_18544,N_17257);
xnor U24608 (N_24608,N_19885,N_19737);
nor U24609 (N_24609,N_19356,N_15025);
or U24610 (N_24610,N_19935,N_19453);
nand U24611 (N_24611,N_16543,N_19814);
nand U24612 (N_24612,N_18069,N_16804);
nor U24613 (N_24613,N_16652,N_18994);
and U24614 (N_24614,N_17117,N_19227);
or U24615 (N_24615,N_18694,N_16881);
nand U24616 (N_24616,N_15309,N_18609);
nand U24617 (N_24617,N_18360,N_18797);
and U24618 (N_24618,N_16473,N_18893);
nor U24619 (N_24619,N_15292,N_17135);
nand U24620 (N_24620,N_19340,N_18893);
nor U24621 (N_24621,N_16330,N_16172);
nor U24622 (N_24622,N_16765,N_19034);
nand U24623 (N_24623,N_15580,N_18586);
or U24624 (N_24624,N_16716,N_17965);
nand U24625 (N_24625,N_16902,N_15150);
nand U24626 (N_24626,N_19015,N_18948);
nor U24627 (N_24627,N_19457,N_16971);
nor U24628 (N_24628,N_19489,N_15686);
and U24629 (N_24629,N_17599,N_15830);
nand U24630 (N_24630,N_18822,N_19232);
or U24631 (N_24631,N_18157,N_17580);
and U24632 (N_24632,N_15649,N_16347);
or U24633 (N_24633,N_16932,N_16878);
nand U24634 (N_24634,N_17973,N_16452);
nand U24635 (N_24635,N_15349,N_19189);
nand U24636 (N_24636,N_19907,N_16808);
or U24637 (N_24637,N_18105,N_15850);
and U24638 (N_24638,N_19754,N_18842);
nor U24639 (N_24639,N_18006,N_16702);
and U24640 (N_24640,N_16352,N_17814);
nor U24641 (N_24641,N_17880,N_18266);
nor U24642 (N_24642,N_18267,N_16535);
and U24643 (N_24643,N_16986,N_15048);
nand U24644 (N_24644,N_15798,N_18371);
nor U24645 (N_24645,N_18124,N_17053);
nor U24646 (N_24646,N_18407,N_17463);
nand U24647 (N_24647,N_17399,N_16641);
nand U24648 (N_24648,N_19150,N_15398);
nand U24649 (N_24649,N_19489,N_17034);
nand U24650 (N_24650,N_18308,N_18866);
and U24651 (N_24651,N_18192,N_16853);
nand U24652 (N_24652,N_17700,N_16806);
or U24653 (N_24653,N_16714,N_16674);
or U24654 (N_24654,N_15958,N_16166);
and U24655 (N_24655,N_15240,N_19766);
or U24656 (N_24656,N_17670,N_15796);
or U24657 (N_24657,N_16571,N_18463);
and U24658 (N_24658,N_15028,N_16581);
nand U24659 (N_24659,N_15608,N_19371);
or U24660 (N_24660,N_18836,N_16671);
or U24661 (N_24661,N_18263,N_18471);
nor U24662 (N_24662,N_15360,N_16095);
or U24663 (N_24663,N_16757,N_19237);
and U24664 (N_24664,N_16036,N_15862);
nand U24665 (N_24665,N_17804,N_19440);
xor U24666 (N_24666,N_19469,N_15976);
nand U24667 (N_24667,N_19313,N_17750);
or U24668 (N_24668,N_17637,N_16603);
xnor U24669 (N_24669,N_17750,N_17153);
nand U24670 (N_24670,N_19681,N_16193);
and U24671 (N_24671,N_19891,N_17891);
nor U24672 (N_24672,N_18736,N_16384);
nand U24673 (N_24673,N_18010,N_19049);
xor U24674 (N_24674,N_15801,N_16076);
and U24675 (N_24675,N_16235,N_15995);
and U24676 (N_24676,N_15043,N_18946);
nand U24677 (N_24677,N_16090,N_18164);
or U24678 (N_24678,N_17259,N_19442);
and U24679 (N_24679,N_19580,N_15154);
and U24680 (N_24680,N_19290,N_16434);
nor U24681 (N_24681,N_16836,N_18162);
nor U24682 (N_24682,N_17918,N_19197);
xor U24683 (N_24683,N_18616,N_16211);
nor U24684 (N_24684,N_16981,N_19887);
nand U24685 (N_24685,N_18645,N_15074);
xor U24686 (N_24686,N_16507,N_18523);
and U24687 (N_24687,N_17126,N_19121);
nand U24688 (N_24688,N_16091,N_18167);
nand U24689 (N_24689,N_18656,N_17050);
or U24690 (N_24690,N_17147,N_19527);
nor U24691 (N_24691,N_15006,N_19240);
or U24692 (N_24692,N_15759,N_15401);
and U24693 (N_24693,N_19859,N_18778);
and U24694 (N_24694,N_15291,N_17533);
and U24695 (N_24695,N_15670,N_17624);
or U24696 (N_24696,N_18484,N_18853);
and U24697 (N_24697,N_19556,N_18669);
xnor U24698 (N_24698,N_17730,N_16077);
nand U24699 (N_24699,N_19384,N_16855);
and U24700 (N_24700,N_18540,N_16214);
and U24701 (N_24701,N_18432,N_19772);
or U24702 (N_24702,N_17815,N_18430);
nor U24703 (N_24703,N_16731,N_19171);
or U24704 (N_24704,N_17727,N_16997);
and U24705 (N_24705,N_16573,N_17853);
nand U24706 (N_24706,N_19513,N_18370);
nand U24707 (N_24707,N_16294,N_16121);
xor U24708 (N_24708,N_15523,N_16041);
nand U24709 (N_24709,N_18338,N_17693);
or U24710 (N_24710,N_17067,N_18211);
nor U24711 (N_24711,N_18395,N_19114);
or U24712 (N_24712,N_15948,N_15332);
nand U24713 (N_24713,N_16887,N_18091);
and U24714 (N_24714,N_15494,N_16304);
or U24715 (N_24715,N_15385,N_16926);
and U24716 (N_24716,N_18483,N_17231);
and U24717 (N_24717,N_15620,N_18247);
or U24718 (N_24718,N_15385,N_19811);
nor U24719 (N_24719,N_16746,N_17943);
and U24720 (N_24720,N_18632,N_19174);
and U24721 (N_24721,N_16423,N_16842);
and U24722 (N_24722,N_16184,N_17318);
and U24723 (N_24723,N_15844,N_17713);
nor U24724 (N_24724,N_16345,N_17067);
nor U24725 (N_24725,N_16423,N_17906);
and U24726 (N_24726,N_18762,N_18148);
nand U24727 (N_24727,N_15527,N_17269);
nand U24728 (N_24728,N_17637,N_19708);
nand U24729 (N_24729,N_18130,N_19863);
xnor U24730 (N_24730,N_17829,N_19399);
nand U24731 (N_24731,N_19406,N_19367);
nand U24732 (N_24732,N_17881,N_16512);
or U24733 (N_24733,N_16172,N_18742);
nand U24734 (N_24734,N_17862,N_15536);
and U24735 (N_24735,N_19424,N_15484);
and U24736 (N_24736,N_19141,N_19839);
or U24737 (N_24737,N_19985,N_16510);
or U24738 (N_24738,N_16487,N_18730);
and U24739 (N_24739,N_19443,N_17356);
or U24740 (N_24740,N_16758,N_17831);
nand U24741 (N_24741,N_19277,N_17662);
and U24742 (N_24742,N_18378,N_19328);
nor U24743 (N_24743,N_15877,N_18018);
or U24744 (N_24744,N_15206,N_16626);
or U24745 (N_24745,N_17327,N_15550);
and U24746 (N_24746,N_15367,N_17985);
nor U24747 (N_24747,N_15967,N_17222);
xor U24748 (N_24748,N_18803,N_16123);
nor U24749 (N_24749,N_17400,N_19313);
xor U24750 (N_24750,N_19226,N_16585);
nor U24751 (N_24751,N_16705,N_19834);
or U24752 (N_24752,N_15836,N_15833);
nor U24753 (N_24753,N_18633,N_15475);
nor U24754 (N_24754,N_16680,N_17657);
xnor U24755 (N_24755,N_18222,N_15410);
or U24756 (N_24756,N_15061,N_15514);
and U24757 (N_24757,N_18914,N_16306);
or U24758 (N_24758,N_17154,N_16872);
nand U24759 (N_24759,N_15103,N_17450);
or U24760 (N_24760,N_18207,N_15092);
and U24761 (N_24761,N_18649,N_17565);
or U24762 (N_24762,N_18956,N_17736);
and U24763 (N_24763,N_18832,N_15137);
nor U24764 (N_24764,N_19088,N_15036);
or U24765 (N_24765,N_19323,N_18764);
and U24766 (N_24766,N_18959,N_19127);
nor U24767 (N_24767,N_16362,N_17165);
and U24768 (N_24768,N_17125,N_19054);
and U24769 (N_24769,N_18496,N_16636);
xor U24770 (N_24770,N_17144,N_16415);
nand U24771 (N_24771,N_17456,N_17558);
and U24772 (N_24772,N_15845,N_16657);
nor U24773 (N_24773,N_16260,N_19115);
and U24774 (N_24774,N_18137,N_18416);
nor U24775 (N_24775,N_17761,N_18569);
nor U24776 (N_24776,N_19190,N_16789);
nand U24777 (N_24777,N_19834,N_18521);
or U24778 (N_24778,N_19246,N_17001);
xnor U24779 (N_24779,N_16031,N_17713);
xor U24780 (N_24780,N_16285,N_17557);
xor U24781 (N_24781,N_16632,N_15255);
and U24782 (N_24782,N_19486,N_16888);
nor U24783 (N_24783,N_15136,N_19688);
or U24784 (N_24784,N_19131,N_17797);
nor U24785 (N_24785,N_17616,N_19008);
or U24786 (N_24786,N_18283,N_19248);
nor U24787 (N_24787,N_15522,N_15575);
and U24788 (N_24788,N_19382,N_16288);
nor U24789 (N_24789,N_17759,N_18190);
or U24790 (N_24790,N_16407,N_17472);
or U24791 (N_24791,N_15591,N_15773);
nor U24792 (N_24792,N_19585,N_17205);
or U24793 (N_24793,N_19710,N_15473);
nand U24794 (N_24794,N_16087,N_18574);
nand U24795 (N_24795,N_16753,N_18061);
nand U24796 (N_24796,N_19125,N_16288);
or U24797 (N_24797,N_17134,N_15705);
nor U24798 (N_24798,N_19827,N_16446);
or U24799 (N_24799,N_17721,N_16859);
and U24800 (N_24800,N_15472,N_17415);
nor U24801 (N_24801,N_17189,N_17070);
nand U24802 (N_24802,N_19597,N_17897);
or U24803 (N_24803,N_15698,N_18513);
nor U24804 (N_24804,N_15210,N_16971);
nor U24805 (N_24805,N_19487,N_16241);
xor U24806 (N_24806,N_19443,N_16684);
nor U24807 (N_24807,N_15304,N_19035);
nand U24808 (N_24808,N_17968,N_19416);
nor U24809 (N_24809,N_15258,N_15236);
nand U24810 (N_24810,N_17729,N_15675);
and U24811 (N_24811,N_17797,N_17304);
nor U24812 (N_24812,N_16041,N_16347);
nor U24813 (N_24813,N_17468,N_17765);
nand U24814 (N_24814,N_15848,N_18961);
and U24815 (N_24815,N_17357,N_15477);
and U24816 (N_24816,N_15419,N_16792);
or U24817 (N_24817,N_19693,N_15912);
nor U24818 (N_24818,N_17351,N_16879);
and U24819 (N_24819,N_18362,N_19655);
xnor U24820 (N_24820,N_15030,N_18273);
nand U24821 (N_24821,N_17697,N_19667);
nor U24822 (N_24822,N_16177,N_18192);
or U24823 (N_24823,N_17572,N_15174);
and U24824 (N_24824,N_16886,N_15302);
nor U24825 (N_24825,N_15361,N_19827);
nand U24826 (N_24826,N_19930,N_19500);
nor U24827 (N_24827,N_15434,N_17086);
and U24828 (N_24828,N_19230,N_18719);
nand U24829 (N_24829,N_18022,N_16156);
or U24830 (N_24830,N_16120,N_15971);
or U24831 (N_24831,N_15574,N_16842);
xor U24832 (N_24832,N_17372,N_16569);
nor U24833 (N_24833,N_17255,N_17862);
or U24834 (N_24834,N_17434,N_17909);
nor U24835 (N_24835,N_18489,N_15281);
nand U24836 (N_24836,N_18171,N_19427);
or U24837 (N_24837,N_17300,N_15976);
and U24838 (N_24838,N_15364,N_18258);
or U24839 (N_24839,N_15984,N_16744);
and U24840 (N_24840,N_17580,N_18213);
and U24841 (N_24841,N_18077,N_16876);
or U24842 (N_24842,N_19828,N_17531);
nand U24843 (N_24843,N_18201,N_18627);
and U24844 (N_24844,N_15822,N_17121);
and U24845 (N_24845,N_18085,N_15966);
nand U24846 (N_24846,N_18820,N_16028);
and U24847 (N_24847,N_17002,N_18404);
or U24848 (N_24848,N_19617,N_19846);
and U24849 (N_24849,N_16038,N_15555);
nand U24850 (N_24850,N_17264,N_16333);
or U24851 (N_24851,N_18332,N_15314);
nand U24852 (N_24852,N_19771,N_15369);
nand U24853 (N_24853,N_19288,N_19079);
nand U24854 (N_24854,N_18124,N_19124);
nor U24855 (N_24855,N_17021,N_19876);
nand U24856 (N_24856,N_17542,N_15867);
and U24857 (N_24857,N_15763,N_15202);
and U24858 (N_24858,N_18026,N_17195);
nand U24859 (N_24859,N_19682,N_17683);
and U24860 (N_24860,N_17365,N_15860);
and U24861 (N_24861,N_16916,N_19504);
or U24862 (N_24862,N_17058,N_15318);
and U24863 (N_24863,N_16970,N_19916);
or U24864 (N_24864,N_16257,N_18470);
or U24865 (N_24865,N_15562,N_19283);
nor U24866 (N_24866,N_19759,N_18394);
nor U24867 (N_24867,N_15034,N_17789);
nor U24868 (N_24868,N_18632,N_18049);
or U24869 (N_24869,N_19502,N_19595);
nor U24870 (N_24870,N_17255,N_17423);
nand U24871 (N_24871,N_15279,N_18615);
nand U24872 (N_24872,N_15735,N_15775);
or U24873 (N_24873,N_16262,N_16972);
and U24874 (N_24874,N_16139,N_16645);
nor U24875 (N_24875,N_18627,N_17284);
and U24876 (N_24876,N_17984,N_16313);
and U24877 (N_24877,N_15929,N_15983);
nor U24878 (N_24878,N_15428,N_16674);
nand U24879 (N_24879,N_19555,N_16533);
nor U24880 (N_24880,N_19305,N_17293);
or U24881 (N_24881,N_17924,N_18457);
xor U24882 (N_24882,N_17592,N_18078);
and U24883 (N_24883,N_15120,N_15130);
nor U24884 (N_24884,N_15529,N_16731);
nor U24885 (N_24885,N_19104,N_19247);
and U24886 (N_24886,N_18493,N_18996);
or U24887 (N_24887,N_17559,N_19675);
nor U24888 (N_24888,N_15034,N_15734);
nor U24889 (N_24889,N_16203,N_19443);
nand U24890 (N_24890,N_19470,N_15690);
nor U24891 (N_24891,N_16934,N_16051);
xor U24892 (N_24892,N_18205,N_17351);
nand U24893 (N_24893,N_17356,N_18381);
and U24894 (N_24894,N_18508,N_16890);
or U24895 (N_24895,N_16170,N_18384);
or U24896 (N_24896,N_16706,N_18842);
xor U24897 (N_24897,N_16353,N_18286);
nor U24898 (N_24898,N_17313,N_15175);
nor U24899 (N_24899,N_16119,N_16797);
nor U24900 (N_24900,N_15624,N_17802);
nand U24901 (N_24901,N_19762,N_18911);
nor U24902 (N_24902,N_16218,N_15332);
or U24903 (N_24903,N_18976,N_17812);
and U24904 (N_24904,N_17513,N_18043);
nand U24905 (N_24905,N_17501,N_17571);
or U24906 (N_24906,N_15555,N_18629);
or U24907 (N_24907,N_17021,N_17136);
nand U24908 (N_24908,N_16567,N_15574);
and U24909 (N_24909,N_19645,N_16043);
nor U24910 (N_24910,N_17547,N_16763);
xnor U24911 (N_24911,N_16843,N_17002);
nand U24912 (N_24912,N_18665,N_19457);
nand U24913 (N_24913,N_18869,N_19662);
or U24914 (N_24914,N_16500,N_19216);
or U24915 (N_24915,N_17656,N_18507);
nor U24916 (N_24916,N_15433,N_17677);
xnor U24917 (N_24917,N_19320,N_19257);
nor U24918 (N_24918,N_16908,N_19462);
nand U24919 (N_24919,N_15928,N_17921);
nand U24920 (N_24920,N_18501,N_16510);
xor U24921 (N_24921,N_19412,N_19330);
nor U24922 (N_24922,N_16163,N_16023);
nor U24923 (N_24923,N_15566,N_19672);
nand U24924 (N_24924,N_17218,N_19547);
nor U24925 (N_24925,N_17222,N_19998);
nor U24926 (N_24926,N_17891,N_19095);
or U24927 (N_24927,N_15648,N_17494);
nand U24928 (N_24928,N_17039,N_15018);
nand U24929 (N_24929,N_17878,N_17048);
nor U24930 (N_24930,N_19083,N_15165);
nand U24931 (N_24931,N_17793,N_18311);
or U24932 (N_24932,N_16718,N_17651);
and U24933 (N_24933,N_16726,N_17633);
or U24934 (N_24934,N_17514,N_19712);
or U24935 (N_24935,N_18680,N_15060);
xor U24936 (N_24936,N_16626,N_15853);
or U24937 (N_24937,N_16948,N_16034);
nor U24938 (N_24938,N_15839,N_18495);
nor U24939 (N_24939,N_19656,N_18617);
nor U24940 (N_24940,N_18627,N_19142);
and U24941 (N_24941,N_18861,N_15910);
and U24942 (N_24942,N_16265,N_18297);
or U24943 (N_24943,N_19087,N_18402);
or U24944 (N_24944,N_16408,N_19566);
and U24945 (N_24945,N_18141,N_18937);
and U24946 (N_24946,N_18696,N_16308);
or U24947 (N_24947,N_15705,N_16592);
nor U24948 (N_24948,N_15469,N_15135);
nand U24949 (N_24949,N_17270,N_18164);
nor U24950 (N_24950,N_18881,N_16232);
or U24951 (N_24951,N_17154,N_16507);
and U24952 (N_24952,N_19426,N_15550);
and U24953 (N_24953,N_19589,N_18263);
and U24954 (N_24954,N_18210,N_16255);
nand U24955 (N_24955,N_19233,N_17216);
and U24956 (N_24956,N_16016,N_17285);
and U24957 (N_24957,N_17908,N_19796);
nand U24958 (N_24958,N_16910,N_17385);
nor U24959 (N_24959,N_17235,N_15314);
or U24960 (N_24960,N_19480,N_19886);
nand U24961 (N_24961,N_15316,N_19834);
nand U24962 (N_24962,N_19381,N_17380);
and U24963 (N_24963,N_17376,N_16632);
and U24964 (N_24964,N_17067,N_17463);
nor U24965 (N_24965,N_16769,N_18471);
nor U24966 (N_24966,N_18377,N_15761);
and U24967 (N_24967,N_19224,N_19911);
and U24968 (N_24968,N_18476,N_19804);
nand U24969 (N_24969,N_17684,N_17542);
or U24970 (N_24970,N_18645,N_15886);
nand U24971 (N_24971,N_18902,N_19216);
and U24972 (N_24972,N_17276,N_17198);
and U24973 (N_24973,N_18342,N_17456);
nor U24974 (N_24974,N_17050,N_18715);
nand U24975 (N_24975,N_19791,N_17862);
or U24976 (N_24976,N_17740,N_17225);
xnor U24977 (N_24977,N_18411,N_15412);
nor U24978 (N_24978,N_19907,N_17722);
and U24979 (N_24979,N_17947,N_15840);
nand U24980 (N_24980,N_19883,N_17076);
nand U24981 (N_24981,N_19238,N_16243);
and U24982 (N_24982,N_18442,N_15963);
nor U24983 (N_24983,N_16791,N_16257);
nor U24984 (N_24984,N_15197,N_18188);
nor U24985 (N_24985,N_18322,N_15108);
or U24986 (N_24986,N_19300,N_16762);
and U24987 (N_24987,N_15277,N_19759);
xor U24988 (N_24988,N_18882,N_17976);
nand U24989 (N_24989,N_16092,N_17956);
nand U24990 (N_24990,N_16674,N_18408);
nand U24991 (N_24991,N_16804,N_15928);
or U24992 (N_24992,N_15535,N_19592);
and U24993 (N_24993,N_15621,N_16250);
nor U24994 (N_24994,N_18916,N_17867);
or U24995 (N_24995,N_16467,N_16424);
nand U24996 (N_24996,N_16925,N_19147);
and U24997 (N_24997,N_17774,N_16728);
nand U24998 (N_24998,N_15514,N_16912);
nand U24999 (N_24999,N_16033,N_16953);
or U25000 (N_25000,N_23324,N_20796);
and U25001 (N_25001,N_23506,N_24404);
nor U25002 (N_25002,N_24806,N_21691);
nor U25003 (N_25003,N_24565,N_20846);
or U25004 (N_25004,N_21720,N_22726);
and U25005 (N_25005,N_20953,N_22751);
nand U25006 (N_25006,N_23206,N_24031);
nand U25007 (N_25007,N_20842,N_23195);
nor U25008 (N_25008,N_20476,N_21052);
and U25009 (N_25009,N_22311,N_24725);
nand U25010 (N_25010,N_20705,N_21296);
and U25011 (N_25011,N_21257,N_22058);
xnor U25012 (N_25012,N_20664,N_20871);
nand U25013 (N_25013,N_20960,N_20653);
nand U25014 (N_25014,N_23732,N_22964);
xor U25015 (N_25015,N_22625,N_24350);
or U25016 (N_25016,N_20732,N_20429);
nand U25017 (N_25017,N_22144,N_23948);
and U25018 (N_25018,N_24080,N_22739);
or U25019 (N_25019,N_24804,N_21463);
nor U25020 (N_25020,N_21405,N_20722);
nand U25021 (N_25021,N_21186,N_22712);
nand U25022 (N_25022,N_20752,N_21306);
nand U25023 (N_25023,N_20158,N_24466);
or U25024 (N_25024,N_21890,N_23331);
or U25025 (N_25025,N_20764,N_22330);
or U25026 (N_25026,N_23704,N_20630);
and U25027 (N_25027,N_20516,N_21985);
and U25028 (N_25028,N_24816,N_23281);
and U25029 (N_25029,N_24023,N_22850);
nand U25030 (N_25030,N_24034,N_24390);
nand U25031 (N_25031,N_24107,N_22286);
or U25032 (N_25032,N_20514,N_22025);
or U25033 (N_25033,N_21141,N_23252);
nand U25034 (N_25034,N_22766,N_24194);
or U25035 (N_25035,N_20982,N_23373);
xnor U25036 (N_25036,N_21277,N_24388);
or U25037 (N_25037,N_21718,N_22041);
nor U25038 (N_25038,N_22655,N_21849);
nand U25039 (N_25039,N_20600,N_23313);
and U25040 (N_25040,N_20777,N_20954);
or U25041 (N_25041,N_21017,N_20091);
or U25042 (N_25042,N_20466,N_21444);
nand U25043 (N_25043,N_22489,N_20591);
nor U25044 (N_25044,N_22646,N_23973);
nand U25045 (N_25045,N_24637,N_24342);
or U25046 (N_25046,N_22167,N_23580);
nor U25047 (N_25047,N_23045,N_22693);
or U25048 (N_25048,N_21863,N_24656);
xnor U25049 (N_25049,N_24065,N_20730);
nand U25050 (N_25050,N_24789,N_23679);
nand U25051 (N_25051,N_23882,N_23077);
and U25052 (N_25052,N_22702,N_23770);
nor U25053 (N_25053,N_21504,N_23174);
or U25054 (N_25054,N_24675,N_24621);
nand U25055 (N_25055,N_21152,N_23030);
or U25056 (N_25056,N_24612,N_23242);
nor U25057 (N_25057,N_22852,N_22876);
and U25058 (N_25058,N_22152,N_24484);
nor U25059 (N_25059,N_21800,N_22658);
and U25060 (N_25060,N_23895,N_23773);
nand U25061 (N_25061,N_23286,N_20488);
or U25062 (N_25062,N_21478,N_22432);
or U25063 (N_25063,N_23249,N_22187);
and U25064 (N_25064,N_21422,N_24084);
xor U25065 (N_25065,N_21237,N_23917);
and U25066 (N_25066,N_24918,N_22734);
nor U25067 (N_25067,N_23156,N_22699);
or U25068 (N_25068,N_21181,N_20017);
nand U25069 (N_25069,N_22283,N_24636);
nand U25070 (N_25070,N_21406,N_21270);
nor U25071 (N_25071,N_21710,N_21189);
and U25072 (N_25072,N_22153,N_24204);
nor U25073 (N_25073,N_20082,N_23122);
or U25074 (N_25074,N_22138,N_20596);
nand U25075 (N_25075,N_21951,N_20532);
nand U25076 (N_25076,N_21185,N_20166);
and U25077 (N_25077,N_24146,N_21906);
nand U25078 (N_25078,N_20921,N_22263);
or U25079 (N_25079,N_24116,N_23932);
xor U25080 (N_25080,N_20186,N_22907);
or U25081 (N_25081,N_20909,N_21260);
xor U25082 (N_25082,N_21748,N_23926);
nor U25083 (N_25083,N_20922,N_23504);
or U25084 (N_25084,N_23959,N_22372);
nor U25085 (N_25085,N_22870,N_23043);
or U25086 (N_25086,N_24000,N_24276);
xor U25087 (N_25087,N_24371,N_24154);
nor U25088 (N_25088,N_20447,N_20864);
nor U25089 (N_25089,N_24422,N_23050);
xnor U25090 (N_25090,N_24890,N_20381);
nand U25091 (N_25091,N_21211,N_20760);
nand U25092 (N_25092,N_23335,N_24938);
nor U25093 (N_25093,N_20622,N_24591);
and U25094 (N_25094,N_21283,N_24764);
or U25095 (N_25095,N_21591,N_24797);
and U25096 (N_25096,N_24483,N_23055);
and U25097 (N_25097,N_22410,N_21001);
xor U25098 (N_25098,N_20357,N_20207);
nand U25099 (N_25099,N_22287,N_21379);
and U25100 (N_25100,N_22196,N_24909);
and U25101 (N_25101,N_20182,N_21923);
nor U25102 (N_25102,N_22357,N_23906);
xor U25103 (N_25103,N_20999,N_23755);
xor U25104 (N_25104,N_22672,N_23224);
nand U25105 (N_25105,N_24322,N_20165);
nor U25106 (N_25106,N_22468,N_21394);
and U25107 (N_25107,N_21264,N_20229);
nand U25108 (N_25108,N_24115,N_23471);
nor U25109 (N_25109,N_20251,N_20454);
and U25110 (N_25110,N_23312,N_20432);
or U25111 (N_25111,N_22742,N_22441);
nor U25112 (N_25112,N_22791,N_24281);
nor U25113 (N_25113,N_21135,N_23622);
nand U25114 (N_25114,N_23523,N_22760);
nor U25115 (N_25115,N_24171,N_23179);
and U25116 (N_25116,N_22096,N_24622);
xor U25117 (N_25117,N_21614,N_20575);
and U25118 (N_25118,N_22368,N_22900);
nand U25119 (N_25119,N_20333,N_21819);
and U25120 (N_25120,N_24510,N_22926);
nor U25121 (N_25121,N_23134,N_24410);
or U25122 (N_25122,N_23595,N_23269);
or U25123 (N_25123,N_21663,N_21558);
nor U25124 (N_25124,N_23792,N_20947);
nand U25125 (N_25125,N_23391,N_22957);
or U25126 (N_25126,N_20606,N_23138);
or U25127 (N_25127,N_20160,N_23176);
and U25128 (N_25128,N_23094,N_22610);
nor U25129 (N_25129,N_23494,N_23382);
nor U25130 (N_25130,N_21364,N_20433);
nand U25131 (N_25131,N_22984,N_21274);
nor U25132 (N_25132,N_22979,N_24412);
nand U25133 (N_25133,N_23688,N_22384);
nor U25134 (N_25134,N_21959,N_24375);
nor U25135 (N_25135,N_24958,N_24288);
and U25136 (N_25136,N_24187,N_24572);
or U25137 (N_25137,N_23485,N_21292);
and U25138 (N_25138,N_22696,N_22663);
or U25139 (N_25139,N_21240,N_20098);
xnor U25140 (N_25140,N_24777,N_22986);
nor U25141 (N_25141,N_20128,N_24181);
or U25142 (N_25142,N_21688,N_20066);
or U25143 (N_25143,N_21332,N_22838);
nor U25144 (N_25144,N_24454,N_23983);
nand U25145 (N_25145,N_21242,N_21142);
or U25146 (N_25146,N_23996,N_23302);
or U25147 (N_25147,N_22199,N_23237);
xnor U25148 (N_25148,N_22763,N_23609);
nand U25149 (N_25149,N_24880,N_21085);
or U25150 (N_25150,N_22163,N_22700);
xor U25151 (N_25151,N_23818,N_21241);
nor U25152 (N_25152,N_24189,N_20255);
nand U25153 (N_25153,N_24014,N_21266);
and U25154 (N_25154,N_23939,N_21537);
or U25155 (N_25155,N_24178,N_20254);
and U25156 (N_25156,N_23082,N_24044);
and U25157 (N_25157,N_20267,N_21054);
xor U25158 (N_25158,N_21158,N_23785);
nor U25159 (N_25159,N_20713,N_24402);
nor U25160 (N_25160,N_21037,N_23786);
or U25161 (N_25161,N_24653,N_22054);
xnor U25162 (N_25162,N_21459,N_23899);
xor U25163 (N_25163,N_23475,N_24716);
or U25164 (N_25164,N_23949,N_23910);
nand U25165 (N_25165,N_20812,N_20996);
nor U25166 (N_25166,N_20015,N_21335);
xor U25167 (N_25167,N_21940,N_21759);
and U25168 (N_25168,N_21816,N_24294);
nor U25169 (N_25169,N_21757,N_22030);
xor U25170 (N_25170,N_21029,N_20721);
xor U25171 (N_25171,N_24134,N_24141);
nand U25172 (N_25172,N_20348,N_23934);
and U25173 (N_25173,N_23665,N_21942);
and U25174 (N_25174,N_24383,N_22029);
nor U25175 (N_25175,N_22430,N_21131);
nand U25176 (N_25176,N_24507,N_24824);
or U25177 (N_25177,N_21225,N_22397);
or U25178 (N_25178,N_22936,N_22776);
nand U25179 (N_25179,N_21174,N_24345);
and U25180 (N_25180,N_20441,N_23065);
nor U25181 (N_25181,N_23225,N_21899);
and U25182 (N_25182,N_24741,N_23809);
and U25183 (N_25183,N_20057,N_21999);
nor U25184 (N_25184,N_24196,N_23482);
and U25185 (N_25185,N_24587,N_24334);
nor U25186 (N_25186,N_21170,N_24414);
or U25187 (N_25187,N_22858,N_24083);
xor U25188 (N_25188,N_24831,N_22222);
nand U25189 (N_25189,N_22818,N_21293);
nand U25190 (N_25190,N_21018,N_20481);
nor U25191 (N_25191,N_24710,N_23651);
and U25192 (N_25192,N_24761,N_22393);
nand U25193 (N_25193,N_24177,N_21986);
or U25194 (N_25194,N_24911,N_22248);
nand U25195 (N_25195,N_20840,N_21735);
and U25196 (N_25196,N_23650,N_23446);
xnor U25197 (N_25197,N_20944,N_24057);
or U25198 (N_25198,N_22094,N_24151);
and U25199 (N_25199,N_20997,N_24287);
or U25200 (N_25200,N_20416,N_24629);
and U25201 (N_25201,N_23112,N_23396);
and U25202 (N_25202,N_21953,N_21763);
nand U25203 (N_25203,N_24211,N_23301);
and U25204 (N_25204,N_20647,N_22069);
nor U25205 (N_25205,N_22374,N_24376);
and U25206 (N_25206,N_23834,N_23379);
nand U25207 (N_25207,N_20623,N_20314);
and U25208 (N_25208,N_20436,N_24055);
nand U25209 (N_25209,N_23291,N_21374);
nand U25210 (N_25210,N_24222,N_24331);
xnor U25211 (N_25211,N_24139,N_20442);
nor U25212 (N_25212,N_21072,N_23952);
nor U25213 (N_25213,N_21705,N_23991);
or U25214 (N_25214,N_20230,N_20593);
or U25215 (N_25215,N_21214,N_23885);
or U25216 (N_25216,N_23388,N_20099);
and U25217 (N_25217,N_24238,N_22972);
nor U25218 (N_25218,N_23553,N_22772);
and U25219 (N_25219,N_24513,N_23576);
nor U25220 (N_25220,N_22262,N_23178);
nor U25221 (N_25221,N_24459,N_23722);
and U25222 (N_25222,N_21419,N_24954);
nor U25223 (N_25223,N_24093,N_23524);
and U25224 (N_25224,N_24967,N_21752);
nand U25225 (N_25225,N_22569,N_24188);
and U25226 (N_25226,N_22684,N_24185);
and U25227 (N_25227,N_21822,N_21132);
nand U25228 (N_25228,N_24326,N_20265);
and U25229 (N_25229,N_23984,N_21471);
or U25230 (N_25230,N_23276,N_21902);
nand U25231 (N_25231,N_22648,N_23240);
nand U25232 (N_25232,N_21082,N_22583);
nor U25233 (N_25233,N_21627,N_22131);
nand U25234 (N_25234,N_20109,N_20523);
and U25235 (N_25235,N_22185,N_20284);
nand U25236 (N_25236,N_21998,N_20029);
nand U25237 (N_25237,N_23871,N_24048);
xor U25238 (N_25238,N_20312,N_21570);
nor U25239 (N_25239,N_20949,N_23491);
or U25240 (N_25240,N_22724,N_22182);
or U25241 (N_25241,N_23498,N_20769);
nand U25242 (N_25242,N_23526,N_23878);
nand U25243 (N_25243,N_21445,N_21144);
nor U25244 (N_25244,N_20761,N_22747);
or U25245 (N_25245,N_23921,N_20998);
or U25246 (N_25246,N_20150,N_20748);
nor U25247 (N_25247,N_21039,N_23493);
nor U25248 (N_25248,N_24360,N_23978);
nand U25249 (N_25249,N_22600,N_20878);
nand U25250 (N_25250,N_24498,N_23909);
or U25251 (N_25251,N_22165,N_21716);
or U25252 (N_25252,N_24776,N_22965);
and U25253 (N_25253,N_24427,N_24872);
or U25254 (N_25254,N_22879,N_23574);
nor U25255 (N_25255,N_20594,N_24198);
and U25256 (N_25256,N_21889,N_22976);
xnor U25257 (N_25257,N_23795,N_22922);
or U25258 (N_25258,N_22433,N_23459);
xnor U25259 (N_25259,N_22156,N_22834);
nand U25260 (N_25260,N_21799,N_24436);
and U25261 (N_25261,N_21555,N_24500);
or U25262 (N_25262,N_24193,N_22890);
xnor U25263 (N_25263,N_23404,N_23121);
nand U25264 (N_25264,N_21818,N_21113);
or U25265 (N_25265,N_24482,N_22950);
xnor U25266 (N_25266,N_24556,N_23708);
nor U25267 (N_25267,N_21060,N_22299);
or U25268 (N_25268,N_22055,N_24730);
and U25269 (N_25269,N_23069,N_24689);
nand U25270 (N_25270,N_21137,N_24791);
nand U25271 (N_25271,N_23659,N_24253);
nor U25272 (N_25272,N_22321,N_20065);
or U25273 (N_25273,N_24568,N_24015);
xor U25274 (N_25274,N_21695,N_20978);
nand U25275 (N_25275,N_24236,N_20520);
nand U25276 (N_25276,N_22475,N_23480);
xor U25277 (N_25277,N_21620,N_20400);
nand U25278 (N_25278,N_21316,N_23836);
nor U25279 (N_25279,N_21837,N_24298);
nand U25280 (N_25280,N_24428,N_22703);
nor U25281 (N_25281,N_21969,N_24532);
nor U25282 (N_25282,N_23115,N_21623);
or U25283 (N_25283,N_22981,N_21308);
or U25284 (N_25284,N_24680,N_23189);
and U25285 (N_25285,N_20503,N_21340);
or U25286 (N_25286,N_22920,N_20360);
or U25287 (N_25287,N_24392,N_21817);
nor U25288 (N_25288,N_21057,N_20686);
and U25289 (N_25289,N_22395,N_23900);
nand U25290 (N_25290,N_22008,N_24129);
nor U25291 (N_25291,N_24038,N_20053);
xor U25292 (N_25292,N_21605,N_24990);
nor U25293 (N_25293,N_20782,N_24068);
nand U25294 (N_25294,N_24813,N_22183);
nand U25295 (N_25295,N_24752,N_22644);
and U25296 (N_25296,N_20773,N_20731);
nor U25297 (N_25297,N_21217,N_23344);
nand U25298 (N_25298,N_22908,N_23469);
or U25299 (N_25299,N_24947,N_24856);
or U25300 (N_25300,N_21284,N_20948);
nand U25301 (N_25301,N_24301,N_22992);
and U25302 (N_25302,N_24553,N_22051);
nor U25303 (N_25303,N_23368,N_21207);
and U25304 (N_25304,N_23215,N_23613);
and U25305 (N_25305,N_21871,N_24695);
or U25306 (N_25306,N_22252,N_24757);
xor U25307 (N_25307,N_23505,N_21034);
xnor U25308 (N_25308,N_21746,N_23245);
nor U25309 (N_25309,N_23430,N_23071);
and U25310 (N_25310,N_24317,N_21832);
nand U25311 (N_25311,N_22186,N_20327);
xnor U25312 (N_25312,N_22867,N_23590);
nand U25313 (N_25313,N_23527,N_23720);
xnor U25314 (N_25314,N_23913,N_23440);
nor U25315 (N_25315,N_20200,N_20618);
or U25316 (N_25316,N_21988,N_21913);
xor U25317 (N_25317,N_22011,N_23953);
nor U25318 (N_25318,N_21930,N_24170);
or U25319 (N_25319,N_23777,N_22994);
nand U25320 (N_25320,N_20311,N_20894);
and U25321 (N_25321,N_22429,N_23719);
nand U25322 (N_25322,N_24095,N_23886);
nor U25323 (N_25323,N_22933,N_20924);
or U25324 (N_25324,N_20231,N_20278);
xnor U25325 (N_25325,N_23352,N_21904);
nand U25326 (N_25326,N_23966,N_21051);
or U25327 (N_25327,N_23337,N_21202);
nand U25328 (N_25328,N_24693,N_22497);
and U25329 (N_25329,N_20859,N_21631);
nor U25330 (N_25330,N_23700,N_20479);
nand U25331 (N_25331,N_21080,N_20887);
and U25332 (N_25332,N_24249,N_21835);
nor U25333 (N_25333,N_22948,N_24597);
nor U25334 (N_25334,N_20869,N_24417);
nor U25335 (N_25335,N_23671,N_24605);
nor U25336 (N_25336,N_24105,N_21288);
nor U25337 (N_25337,N_20174,N_23967);
nand U25338 (N_25338,N_22151,N_23113);
nand U25339 (N_25339,N_21852,N_21020);
xnor U25340 (N_25340,N_23167,N_21071);
or U25341 (N_25341,N_20681,N_21022);
and U25342 (N_25342,N_21026,N_24949);
nand U25343 (N_25343,N_20958,N_22579);
xor U25344 (N_25344,N_23848,N_24818);
and U25345 (N_25345,N_23799,N_22173);
nor U25346 (N_25346,N_24986,N_20990);
and U25347 (N_25347,N_22479,N_24843);
xnor U25348 (N_25348,N_23188,N_21924);
and U25349 (N_25349,N_24749,N_21190);
nor U25350 (N_25350,N_21616,N_23323);
xor U25351 (N_25351,N_23976,N_24913);
or U25352 (N_25352,N_21858,N_22520);
nor U25353 (N_25353,N_22768,N_20486);
nor U25354 (N_25354,N_22954,N_21511);
and U25355 (N_25355,N_23147,N_21253);
nand U25356 (N_25356,N_20295,N_22371);
nor U25357 (N_25357,N_23296,N_22634);
nand U25358 (N_25358,N_24114,N_23308);
or U25359 (N_25359,N_23101,N_21676);
and U25360 (N_25360,N_22603,N_24098);
xnor U25361 (N_25361,N_21854,N_20347);
nor U25362 (N_25362,N_21823,N_21291);
or U25363 (N_25363,N_24155,N_23262);
or U25364 (N_25364,N_22504,N_21365);
nor U25365 (N_25365,N_20562,N_22709);
nand U25366 (N_25366,N_20236,N_22670);
nor U25367 (N_25367,N_21510,N_24150);
or U25368 (N_25368,N_21880,N_24252);
or U25369 (N_25369,N_24664,N_23640);
nand U25370 (N_25370,N_20077,N_21154);
xor U25371 (N_25371,N_23304,N_21128);
nor U25372 (N_25372,N_20838,N_20192);
or U25373 (N_25373,N_22340,N_22974);
nand U25374 (N_25374,N_24758,N_21140);
and U25375 (N_25375,N_23782,N_23803);
or U25376 (N_25376,N_22808,N_22329);
nor U25377 (N_25377,N_23017,N_24729);
or U25378 (N_25378,N_24324,N_22581);
or U25379 (N_25379,N_24128,N_22750);
or U25380 (N_25380,N_20468,N_23058);
nor U25381 (N_25381,N_22271,N_24200);
and U25382 (N_25382,N_23319,N_21779);
and U25383 (N_25383,N_21680,N_23295);
and U25384 (N_25384,N_20807,N_24078);
and U25385 (N_25385,N_24579,N_24224);
nor U25386 (N_25386,N_22009,N_23938);
nand U25387 (N_25387,N_24453,N_23813);
xnor U25388 (N_25388,N_21625,N_24923);
or U25389 (N_25389,N_22293,N_20215);
nor U25390 (N_25390,N_21715,N_24275);
nor U25391 (N_25391,N_22109,N_24739);
nor U25392 (N_25392,N_21758,N_21641);
xnor U25393 (N_25393,N_24104,N_21441);
or U25394 (N_25394,N_20781,N_21220);
xor U25395 (N_25395,N_21978,N_23843);
or U25396 (N_25396,N_24993,N_24610);
and U25397 (N_25397,N_20176,N_22949);
and U25398 (N_25398,N_24136,N_22927);
nand U25399 (N_25399,N_22324,N_21601);
and U25400 (N_25400,N_23383,N_23032);
xor U25401 (N_25401,N_20984,N_24047);
or U25402 (N_25402,N_23078,N_21084);
nand U25403 (N_25403,N_20072,N_21066);
nor U25404 (N_25404,N_24348,N_22653);
and U25405 (N_25405,N_23145,N_21329);
nand U25406 (N_25406,N_23963,N_24346);
or U25407 (N_25407,N_20185,N_24940);
and U25408 (N_25408,N_24291,N_22480);
nand U25409 (N_25409,N_21370,N_23729);
nor U25410 (N_25410,N_20242,N_24602);
nor U25411 (N_25411,N_22595,N_20007);
nor U25412 (N_25412,N_20202,N_20256);
and U25413 (N_25413,N_20844,N_23946);
xnor U25414 (N_25414,N_20492,N_23100);
nand U25415 (N_25415,N_20977,N_24506);
or U25416 (N_25416,N_22465,N_22202);
and U25417 (N_25417,N_20213,N_24691);
xnor U25418 (N_25418,N_21059,N_23555);
and U25419 (N_25419,N_21783,N_22692);
nand U25420 (N_25420,N_22515,N_21133);
xor U25421 (N_25421,N_24679,N_20405);
and U25422 (N_25422,N_20518,N_20536);
and U25423 (N_25423,N_23087,N_20526);
and U25424 (N_25424,N_23823,N_20786);
or U25425 (N_25425,N_22066,N_23995);
nor U25426 (N_25426,N_20271,N_22540);
and U25427 (N_25427,N_22110,N_22020);
nor U25428 (N_25428,N_21315,N_24829);
xnor U25429 (N_25429,N_24518,N_23896);
nor U25430 (N_25430,N_24678,N_22975);
nor U25431 (N_25431,N_20170,N_23644);
nor U25432 (N_25432,N_23194,N_24477);
or U25433 (N_25433,N_24216,N_23131);
and U25434 (N_25434,N_20701,N_22048);
and U25435 (N_25435,N_22416,N_21247);
and U25436 (N_25436,N_23582,N_20275);
or U25437 (N_25437,N_23608,N_21653);
or U25438 (N_25438,N_21110,N_22973);
nor U25439 (N_25439,N_23479,N_23979);
or U25440 (N_25440,N_23033,N_22690);
or U25441 (N_25441,N_22115,N_24707);
nand U25442 (N_25442,N_24335,N_23841);
nand U25443 (N_25443,N_24369,N_21425);
nand U25444 (N_25444,N_20024,N_22748);
or U25445 (N_25445,N_22661,N_22740);
nor U25446 (N_25446,N_20349,N_21377);
nand U25447 (N_25447,N_23250,N_23024);
and U25448 (N_25448,N_20819,N_24669);
or U25449 (N_25449,N_20666,N_23117);
or U25450 (N_25450,N_22951,N_24700);
or U25451 (N_25451,N_22854,N_24479);
or U25452 (N_25452,N_24961,N_24087);
or U25453 (N_25453,N_22026,N_24895);
or U25454 (N_25454,N_21290,N_23051);
nand U25455 (N_25455,N_24836,N_21661);
and U25456 (N_25456,N_23175,N_20167);
nand U25457 (N_25457,N_22608,N_21032);
and U25458 (N_25458,N_20813,N_20407);
xor U25459 (N_25459,N_21023,N_24751);
or U25460 (N_25460,N_22729,N_24305);
or U25461 (N_25461,N_22458,N_22963);
nand U25462 (N_25462,N_20232,N_24391);
and U25463 (N_25463,N_22626,N_23762);
or U25464 (N_25464,N_23894,N_20248);
nor U25465 (N_25465,N_24606,N_21624);
nor U25466 (N_25466,N_22320,N_24699);
and U25467 (N_25467,N_23954,N_20219);
and U25468 (N_25468,N_20849,N_24473);
nand U25469 (N_25469,N_22356,N_24340);
or U25470 (N_25470,N_23827,N_20391);
xnor U25471 (N_25471,N_21903,N_21326);
nand U25472 (N_25472,N_23484,N_20413);
or U25473 (N_25473,N_20801,N_22237);
nand U25474 (N_25474,N_22212,N_20803);
nand U25475 (N_25475,N_20541,N_21884);
nor U25476 (N_25476,N_23342,N_22560);
nand U25477 (N_25477,N_22482,N_24060);
nand U25478 (N_25478,N_23448,N_20788);
or U25479 (N_25479,N_24694,N_22180);
xnor U25480 (N_25480,N_23897,N_24997);
nand U25481 (N_25481,N_20943,N_24685);
or U25482 (N_25482,N_20089,N_22457);
or U25483 (N_25483,N_22073,N_21865);
and U25484 (N_25484,N_21442,N_22304);
nand U25485 (N_25485,N_22921,N_24991);
and U25486 (N_25486,N_20854,N_21106);
nor U25487 (N_25487,N_22488,N_20553);
xor U25488 (N_25488,N_21475,N_24912);
nand U25489 (N_25489,N_24163,N_24732);
nand U25490 (N_25490,N_23341,N_24557);
nor U25491 (N_25491,N_20190,N_21188);
and U25492 (N_25492,N_24663,N_20865);
xor U25493 (N_25493,N_20249,N_21950);
nor U25494 (N_25494,N_20445,N_23683);
xnor U25495 (N_25495,N_21921,N_21428);
xor U25496 (N_25496,N_22354,N_24564);
or U25497 (N_25497,N_21790,N_20003);
nor U25498 (N_25498,N_22998,N_21298);
nor U25499 (N_25499,N_21512,N_20790);
xnor U25500 (N_25500,N_24359,N_24365);
or U25501 (N_25501,N_24205,N_21399);
and U25502 (N_25502,N_22238,N_24930);
or U25503 (N_25503,N_24355,N_23974);
or U25504 (N_25504,N_21311,N_20464);
and U25505 (N_25505,N_22911,N_20086);
nand U25506 (N_25506,N_23763,N_20610);
or U25507 (N_25507,N_24312,N_22942);
or U25508 (N_25508,N_24600,N_23208);
nor U25509 (N_25509,N_22099,N_24493);
and U25510 (N_25510,N_24952,N_21393);
or U25511 (N_25511,N_23549,N_22122);
xnor U25512 (N_25512,N_21747,N_21829);
nand U25513 (N_25513,N_24344,N_21717);
nand U25514 (N_25514,N_21908,N_21476);
nand U25515 (N_25515,N_22197,N_24212);
nand U25516 (N_25516,N_23380,N_23703);
and U25517 (N_25517,N_24096,N_21856);
or U25518 (N_25518,N_24648,N_23346);
nand U25519 (N_25519,N_24618,N_22300);
or U25520 (N_25520,N_20968,N_20315);
or U25521 (N_25521,N_22327,N_22511);
nor U25522 (N_25522,N_24394,N_23309);
nor U25523 (N_25523,N_21030,N_21159);
or U25524 (N_25524,N_21431,N_24601);
and U25525 (N_25525,N_20749,N_23793);
nand U25526 (N_25526,N_22711,N_22568);
or U25527 (N_25527,N_24463,N_21500);
and U25528 (N_25528,N_24633,N_22208);
nand U25529 (N_25529,N_20321,N_20453);
nand U25530 (N_25530,N_22141,N_22087);
and U25531 (N_25531,N_24906,N_21496);
xnor U25532 (N_25532,N_22977,N_22015);
or U25533 (N_25533,N_23663,N_22542);
nand U25534 (N_25534,N_23349,N_22514);
nor U25535 (N_25535,N_22561,N_21990);
xnor U25536 (N_25536,N_20475,N_24873);
nand U25537 (N_25537,N_23544,N_20026);
nor U25538 (N_25538,N_23359,N_20477);
nor U25539 (N_25539,N_24647,N_23940);
and U25540 (N_25540,N_21786,N_23985);
and U25541 (N_25541,N_20364,N_20995);
nand U25542 (N_25542,N_21321,N_22413);
or U25543 (N_25543,N_24118,N_20884);
or U25544 (N_25544,N_21839,N_21369);
nor U25545 (N_25545,N_22848,N_22334);
or U25546 (N_25546,N_22464,N_21304);
nand U25547 (N_25547,N_23472,N_22898);
and U25548 (N_25548,N_23496,N_22469);
nor U25549 (N_25549,N_23508,N_22070);
nor U25550 (N_25550,N_24984,N_23883);
nand U25551 (N_25551,N_24852,N_23833);
nor U25552 (N_25552,N_22481,N_20292);
nand U25553 (N_25553,N_24541,N_20642);
and U25554 (N_25554,N_21646,N_23787);
nand U25555 (N_25555,N_20123,N_24070);
and U25556 (N_25556,N_20474,N_23560);
nor U25557 (N_25557,N_20142,N_22917);
or U25558 (N_25558,N_22004,N_20262);
xnor U25559 (N_25559,N_20724,N_20266);
and U25560 (N_25560,N_24972,N_24218);
nor U25561 (N_25561,N_23829,N_20935);
or U25562 (N_25562,N_23003,N_23705);
or U25563 (N_25563,N_21499,N_21983);
or U25564 (N_25564,N_21384,N_24955);
nor U25565 (N_25565,N_22744,N_20741);
nand U25566 (N_25566,N_22798,N_21677);
nor U25567 (N_25567,N_22851,N_21019);
or U25568 (N_25568,N_21935,N_23365);
or U25569 (N_25569,N_20480,N_22820);
xnor U25570 (N_25570,N_20635,N_24882);
and U25571 (N_25571,N_22459,N_24870);
and U25572 (N_25572,N_22507,N_23764);
nand U25573 (N_25573,N_22585,N_20750);
nor U25574 (N_25574,N_20798,N_24119);
nor U25575 (N_25575,N_23625,N_24546);
or U25576 (N_25576,N_23196,N_24674);
and U25577 (N_25577,N_21898,N_23274);
nor U25578 (N_25578,N_22335,N_22874);
and U25579 (N_25579,N_24814,N_22909);
nand U25580 (N_25580,N_22767,N_20395);
xor U25581 (N_25581,N_20472,N_24891);
nor U25582 (N_25582,N_20665,N_24295);
nand U25583 (N_25583,N_24595,N_24770);
nor U25584 (N_25584,N_20209,N_23318);
and U25585 (N_25585,N_20950,N_20143);
xnor U25586 (N_25586,N_20028,N_24377);
and U25587 (N_25587,N_23903,N_21645);
or U25588 (N_25588,N_22717,N_22407);
xnor U25589 (N_25589,N_20052,N_24140);
and U25590 (N_25590,N_23586,N_23059);
and U25591 (N_25591,N_23858,N_24424);
and U25592 (N_25592,N_23137,N_21003);
nor U25593 (N_25593,N_22945,N_21657);
xor U25594 (N_25594,N_20012,N_22524);
and U25595 (N_25595,N_20130,N_23627);
nand U25596 (N_25596,N_22343,N_22349);
xor U25597 (N_25597,N_24123,N_21485);
or U25598 (N_25598,N_21285,N_24736);
nand U25599 (N_25599,N_23745,N_21138);
and U25600 (N_25600,N_22731,N_21010);
or U25601 (N_25601,N_21878,N_20671);
nand U25602 (N_25602,N_22040,N_20509);
and U25603 (N_25603,N_24667,N_20323);
nor U25604 (N_25604,N_24438,N_22529);
nor U25605 (N_25605,N_22150,N_24373);
nor U25606 (N_25606,N_22573,N_21409);
and U25607 (N_25607,N_22273,N_21972);
nand U25608 (N_25608,N_21363,N_24016);
or U25609 (N_25609,N_22219,N_20155);
or U25610 (N_25610,N_23105,N_21012);
or U25611 (N_25611,N_24109,N_21473);
nand U25612 (N_25612,N_24001,N_23605);
and U25613 (N_25613,N_24871,N_22784);
nand U25614 (N_25614,N_20547,N_22398);
nor U25615 (N_25615,N_23497,N_24508);
xnor U25616 (N_25616,N_23172,N_24248);
or U25617 (N_25617,N_24303,N_23754);
or U25618 (N_25618,N_24166,N_22841);
and U25619 (N_25619,N_23148,N_21666);
and U25620 (N_25620,N_24135,N_22934);
nand U25621 (N_25621,N_22039,N_22506);
or U25622 (N_25622,N_20394,N_22012);
xnor U25623 (N_25623,N_20451,N_20951);
or U25624 (N_25624,N_21047,N_22752);
nand U25625 (N_25625,N_20450,N_22113);
nor U25626 (N_25626,N_24615,N_24755);
or U25627 (N_25627,N_23311,N_23880);
nor U25628 (N_25628,N_20524,N_21464);
nor U25629 (N_25629,N_21078,N_20319);
or U25630 (N_25630,N_21098,N_24783);
or U25631 (N_25631,N_24026,N_20279);
nor U25632 (N_25632,N_23876,N_21539);
nand U25633 (N_25633,N_21469,N_21045);
nand U25634 (N_25634,N_21104,N_24687);
and U25635 (N_25635,N_23091,N_20156);
nand U25636 (N_25636,N_21233,N_20885);
and U25637 (N_25637,N_21014,N_24889);
xor U25638 (N_25638,N_20994,N_20818);
and U25639 (N_25639,N_23686,N_20409);
xor U25640 (N_25640,N_24468,N_22946);
and U25641 (N_25641,N_22582,N_22623);
and U25642 (N_25642,N_23102,N_22759);
nor U25643 (N_25643,N_21299,N_20237);
or U25644 (N_25644,N_24754,N_21774);
nand U25645 (N_25645,N_22000,N_22057);
nor U25646 (N_25646,N_21659,N_21724);
nor U25647 (N_25647,N_23861,N_23185);
or U25648 (N_25648,N_21491,N_23125);
or U25649 (N_25649,N_22154,N_23092);
and U25650 (N_25650,N_22652,N_24948);
or U25651 (N_25651,N_22741,N_22336);
or U25652 (N_25652,N_20328,N_21089);
nor U25653 (N_25653,N_21789,N_20191);
or U25654 (N_25654,N_21427,N_24946);
or U25655 (N_25655,N_20038,N_21212);
or U25656 (N_25656,N_22842,N_22875);
xor U25657 (N_25657,N_22082,N_22386);
or U25658 (N_25658,N_22135,N_21704);
and U25659 (N_25659,N_22332,N_21305);
nor U25660 (N_25660,N_21434,N_22725);
nand U25661 (N_25661,N_20023,N_23390);
nand U25662 (N_25662,N_21551,N_21147);
or U25663 (N_25663,N_20855,N_20351);
or U25664 (N_25664,N_22801,N_20976);
nand U25665 (N_25665,N_24826,N_23411);
and U25666 (N_25666,N_24443,N_21199);
nand U25667 (N_25667,N_24266,N_20302);
nor U25668 (N_25668,N_20907,N_21203);
and U25669 (N_25669,N_21862,N_21901);
nor U25670 (N_25670,N_23830,N_22859);
nor U25671 (N_25671,N_20178,N_22785);
nand U25672 (N_25672,N_24063,N_24869);
or U25673 (N_25673,N_22987,N_24030);
and U25674 (N_25674,N_24432,N_20542);
nand U25675 (N_25675,N_22315,N_23466);
nor U25676 (N_25676,N_24067,N_22679);
nor U25677 (N_25677,N_24709,N_21834);
nor U25678 (N_25678,N_22415,N_24378);
xor U25679 (N_25679,N_21338,N_20690);
and U25680 (N_25680,N_20538,N_23007);
nand U25681 (N_25681,N_21224,N_22580);
or U25682 (N_25682,N_21655,N_21672);
nand U25683 (N_25683,N_22268,N_21325);
nor U25684 (N_25684,N_24530,N_22421);
nand U25685 (N_25685,N_23419,N_23718);
or U25686 (N_25686,N_21262,N_20212);
nor U25687 (N_25687,N_20181,N_22201);
and U25688 (N_25688,N_22816,N_22538);
nand U25689 (N_25689,N_22795,N_21629);
nor U25690 (N_25690,N_24481,N_20148);
nand U25691 (N_25691,N_22997,N_20793);
nor U25692 (N_25692,N_22490,N_23387);
nand U25693 (N_25693,N_23692,N_21693);
and U25694 (N_25694,N_23643,N_23402);
and U25695 (N_25695,N_23744,N_22651);
and U25696 (N_25696,N_20964,N_23442);
nor U25697 (N_25697,N_22125,N_24441);
nand U25698 (N_25698,N_24718,N_23213);
nor U25699 (N_25699,N_22414,N_24296);
nor U25700 (N_25700,N_21300,N_23588);
nor U25701 (N_25701,N_20329,N_21557);
and U25702 (N_25702,N_21125,N_23399);
nor U25703 (N_25703,N_21836,N_20927);
nand U25704 (N_25704,N_23698,N_24850);
and U25705 (N_25705,N_21286,N_24926);
or U25706 (N_25706,N_24698,N_21801);
or U25707 (N_25707,N_23293,N_22189);
xor U25708 (N_25708,N_23461,N_22824);
or U25709 (N_25709,N_21341,N_20051);
nand U25710 (N_25710,N_23120,N_20320);
or U25711 (N_25711,N_24142,N_24274);
nor U25712 (N_25712,N_23397,N_20078);
and U25713 (N_25713,N_20205,N_20899);
nor U25714 (N_25714,N_23816,N_24284);
or U25715 (N_25715,N_23751,N_20092);
and U25716 (N_25716,N_23982,N_24165);
nand U25717 (N_25717,N_22800,N_23048);
nand U25718 (N_25718,N_21637,N_20422);
nand U25719 (N_25719,N_24386,N_22272);
or U25720 (N_25720,N_23254,N_20605);
and U25721 (N_25721,N_21579,N_24802);
xor U25722 (N_25722,N_23476,N_22778);
or U25723 (N_25723,N_21302,N_23290);
nor U25724 (N_25724,N_24963,N_23824);
nand U25725 (N_25725,N_24077,N_23420);
or U25726 (N_25726,N_21230,N_22993);
and U25727 (N_25727,N_20355,N_23695);
and U25728 (N_25728,N_20800,N_24830);
nand U25729 (N_25729,N_24233,N_22172);
and U25730 (N_25730,N_23186,N_24769);
or U25731 (N_25731,N_22269,N_24992);
nor U25732 (N_25732,N_23021,N_24032);
xor U25733 (N_25733,N_21375,N_20804);
nor U25734 (N_25734,N_23925,N_21974);
or U25735 (N_25735,N_23587,N_24713);
or U25736 (N_25736,N_22826,N_21991);
nor U25737 (N_25737,N_20380,N_21725);
nand U25738 (N_25738,N_21900,N_23656);
nor U25739 (N_25739,N_21977,N_22517);
xor U25740 (N_25740,N_23398,N_20224);
and U25741 (N_25741,N_21702,N_22140);
xnor U25742 (N_25742,N_23628,N_22732);
and U25743 (N_25743,N_24120,N_21313);
and U25744 (N_25744,N_24632,N_21421);
and U25745 (N_25745,N_22380,N_21401);
nand U25746 (N_25746,N_22621,N_22302);
nor U25747 (N_25747,N_24537,N_24846);
nand U25748 (N_25748,N_23096,N_23619);
nor U25749 (N_25749,N_24550,N_22442);
and U25750 (N_25750,N_22807,N_20244);
xor U25751 (N_25751,N_20264,N_20289);
nand U25752 (N_25752,N_21802,N_24258);
or U25753 (N_25753,N_20382,N_20611);
or U25754 (N_25754,N_22342,N_21494);
or U25755 (N_25755,N_20134,N_23918);
and U25756 (N_25756,N_20602,N_24599);
and U25757 (N_25757,N_23429,N_20404);
or U25758 (N_25758,N_24863,N_24859);
or U25759 (N_25759,N_20316,N_20636);
and U25760 (N_25760,N_21671,N_20709);
nor U25761 (N_25761,N_22243,N_20408);
and U25762 (N_25762,N_23778,N_24103);
and U25763 (N_25763,N_22347,N_22373);
nor U25764 (N_25764,N_21073,N_21261);
nor U25765 (N_25765,N_20246,N_22467);
or U25766 (N_25766,N_24786,N_24671);
xnor U25767 (N_25767,N_22285,N_21634);
nand U25768 (N_25768,N_24130,N_24184);
or U25769 (N_25769,N_22227,N_23328);
nand U25770 (N_25770,N_23289,N_22101);
or U25771 (N_25771,N_20079,N_24138);
or U25772 (N_25772,N_24666,N_21454);
nor U25773 (N_25773,N_22194,N_23875);
nand U25774 (N_25774,N_24692,N_23532);
nor U25775 (N_25775,N_22193,N_22510);
nand U25776 (N_25776,N_22487,N_20897);
xor U25777 (N_25777,N_24668,N_22387);
and U25778 (N_25778,N_24381,N_22891);
nand U25779 (N_25779,N_21893,N_20490);
nand U25780 (N_25780,N_20966,N_24677);
nand U25781 (N_25781,N_24478,N_22642);
and U25782 (N_25782,N_23728,N_21568);
nand U25783 (N_25783,N_23641,N_21895);
or U25784 (N_25784,N_22117,N_24174);
nand U25785 (N_25785,N_21446,N_20847);
xor U25786 (N_25786,N_23013,N_21544);
and U25787 (N_25787,N_24714,N_20423);
or U25788 (N_25788,N_23676,N_23298);
nor U25789 (N_25789,N_20214,N_21883);
nand U25790 (N_25790,N_21443,N_24019);
and U25791 (N_25791,N_22590,N_22897);
nand U25792 (N_25792,N_24515,N_23811);
nor U25793 (N_25793,N_21997,N_20568);
or U25794 (N_25794,N_21967,N_24328);
nand U25795 (N_25795,N_20707,N_22567);
and U25796 (N_25796,N_24620,N_24835);
and U25797 (N_25797,N_24090,N_24996);
and U25798 (N_25798,N_21611,N_20062);
xor U25799 (N_25799,N_22355,N_20698);
and U25800 (N_25800,N_23283,N_20728);
and U25801 (N_25801,N_21356,N_24405);
xor U25802 (N_25802,N_21006,N_21946);
or U25803 (N_25803,N_20607,N_22005);
xnor U25804 (N_25804,N_22390,N_21420);
xor U25805 (N_25805,N_24649,N_24919);
or U25806 (N_25806,N_24400,N_24214);
nor U25807 (N_25807,N_23322,N_23866);
and U25808 (N_25808,N_21867,N_21038);
or U25809 (N_25809,N_24226,N_22074);
and U25810 (N_25810,N_23181,N_22278);
nor U25811 (N_25811,N_23143,N_20992);
or U25812 (N_25812,N_22547,N_23579);
or U25813 (N_25813,N_24720,N_24995);
nor U25814 (N_25814,N_21008,N_22123);
and U25815 (N_25815,N_23951,N_20608);
nand U25816 (N_25816,N_23334,N_20448);
and U25817 (N_25817,N_24594,N_20833);
nand U25818 (N_25818,N_20579,N_20008);
xnor U25819 (N_25819,N_24033,N_21542);
nor U25820 (N_25820,N_20794,N_20088);
or U25821 (N_25821,N_21339,N_23768);
or U25822 (N_25822,N_24505,N_21255);
nor U25823 (N_25823,N_24723,N_24753);
nand U25824 (N_25824,N_23986,N_22006);
and U25825 (N_25825,N_21065,N_23749);
nand U25826 (N_25826,N_20826,N_24313);
and U25827 (N_25827,N_21915,N_23060);
nand U25828 (N_25828,N_21712,N_20649);
or U25829 (N_25829,N_22112,N_20034);
nand U25830 (N_25830,N_24857,N_20745);
nor U25831 (N_25831,N_24511,N_20934);
or U25832 (N_25832,N_23486,N_21228);
or U25833 (N_25833,N_23336,N_24061);
nor U25834 (N_25834,N_23604,N_23944);
or U25835 (N_25835,N_23759,N_24273);
and U25836 (N_25836,N_21575,N_22982);
xnor U25837 (N_25837,N_24382,N_20621);
and U25838 (N_25838,N_24583,N_23244);
and U25839 (N_25839,N_23950,N_21108);
nor U25840 (N_25840,N_22129,N_21656);
and U25841 (N_25841,N_22425,N_24903);
nor U25842 (N_25842,N_23847,N_20019);
or U25843 (N_25843,N_23093,N_22284);
nand U25844 (N_25844,N_21886,N_22217);
xor U25845 (N_25845,N_20048,N_21102);
nand U25846 (N_25846,N_22225,N_24172);
xor U25847 (N_25847,N_23488,N_24379);
nor U25848 (N_25848,N_21536,N_20720);
nand U25849 (N_25849,N_21124,N_21552);
nor U25850 (N_25850,N_21766,N_20900);
nor U25851 (N_25851,N_20739,N_23106);
nor U25852 (N_25852,N_22594,N_23908);
nand U25853 (N_25853,N_23081,N_22525);
or U25854 (N_25854,N_20263,N_22297);
and U25855 (N_25855,N_24041,N_24853);
nand U25856 (N_25856,N_20904,N_22147);
and U25857 (N_25857,N_22961,N_21885);
nor U25858 (N_25858,N_22647,N_24028);
nand U25859 (N_25859,N_24091,N_24197);
nand U25860 (N_25860,N_23839,N_22830);
and U25861 (N_25861,N_24861,N_22901);
and U25862 (N_25862,N_23920,N_20776);
xor U25863 (N_25863,N_22587,N_21777);
nand U25864 (N_25864,N_20983,N_23168);
nor U25865 (N_25865,N_21429,N_24354);
or U25866 (N_25866,N_21600,N_23351);
nand U25867 (N_25867,N_24179,N_20696);
or U25868 (N_25868,N_24356,N_20862);
and U25869 (N_25869,N_20159,N_21821);
or U25870 (N_25870,N_24766,N_23812);
or U25871 (N_25871,N_20268,N_21843);
or U25872 (N_25872,N_22512,N_20563);
nand U25873 (N_25873,N_21840,N_20070);
and U25874 (N_25874,N_23804,N_21456);
nand U25875 (N_25875,N_23463,N_21391);
or U25876 (N_25876,N_20716,N_23104);
nand U25877 (N_25877,N_24064,N_22723);
nand U25878 (N_25878,N_22176,N_20513);
and U25879 (N_25879,N_23273,N_24147);
and U25880 (N_25880,N_22501,N_23546);
xnor U25881 (N_25881,N_21227,N_24514);
nor U25882 (N_25882,N_20689,N_20358);
xnor U25883 (N_25883,N_22839,N_23035);
nand U25884 (N_25884,N_20482,N_22177);
nand U25885 (N_25885,N_22853,N_20458);
nor U25886 (N_25886,N_20870,N_23265);
or U25887 (N_25887,N_22913,N_20094);
nand U25888 (N_25888,N_24796,N_20435);
nor U25889 (N_25889,N_20645,N_24966);
or U25890 (N_25890,N_24635,N_21449);
and U25891 (N_25891,N_24223,N_23023);
nor U25892 (N_25892,N_21268,N_24418);
and U25893 (N_25893,N_21971,N_20586);
xor U25894 (N_25894,N_20714,N_22735);
or U25895 (N_25895,N_21083,N_22381);
and U25896 (N_25896,N_20925,N_21626);
nand U25897 (N_25897,N_23253,N_20457);
and U25898 (N_25898,N_22686,N_20428);
and U25899 (N_25899,N_22519,N_22714);
nor U25900 (N_25900,N_24801,N_21015);
nor U25901 (N_25901,N_23474,N_21642);
nor U25902 (N_25902,N_23356,N_24158);
and U25903 (N_25903,N_24229,N_22067);
nand U25904 (N_25904,N_22978,N_23251);
nor U25905 (N_25905,N_23614,N_24848);
nor U25906 (N_25906,N_20455,N_24800);
nand U25907 (N_25907,N_22523,N_22799);
and U25908 (N_25908,N_22046,N_22781);
nand U25909 (N_25909,N_23901,N_24894);
nand U25910 (N_25910,N_23173,N_23109);
or U25911 (N_25911,N_20569,N_23052);
nand U25912 (N_25912,N_22584,N_24458);
or U25913 (N_25913,N_20036,N_20340);
xnor U25914 (N_25914,N_23757,N_21684);
nand U25915 (N_25915,N_22181,N_20067);
nand U25916 (N_25916,N_23533,N_20857);
or U25917 (N_25917,N_21120,N_23232);
and U25918 (N_25918,N_20733,N_20961);
nor U25919 (N_25919,N_24838,N_24884);
nand U25920 (N_25920,N_24696,N_24520);
nor U25921 (N_25921,N_22052,N_21675);
nand U25922 (N_25922,N_22204,N_23080);
or U25923 (N_25923,N_22382,N_20203);
nand U25924 (N_25924,N_21027,N_20784);
nor U25925 (N_25925,N_20054,N_24673);
xnor U25926 (N_25926,N_24785,N_23715);
nand U25927 (N_25927,N_21498,N_20867);
or U25928 (N_25928,N_20440,N_20059);
nand U25929 (N_25929,N_21169,N_23453);
nand U25930 (N_25930,N_21529,N_20478);
and U25931 (N_25931,N_20699,N_20548);
or U25932 (N_25932,N_24533,N_20969);
nand U25933 (N_25933,N_22969,N_23507);
and U25934 (N_25934,N_20712,N_23489);
nor U25935 (N_25935,N_22555,N_21244);
nor U25936 (N_25936,N_20661,N_21352);
nor U25937 (N_25937,N_21093,N_20106);
nand U25938 (N_25938,N_22084,N_20866);
or U25939 (N_25939,N_21973,N_24787);
nand U25940 (N_25940,N_21079,N_21432);
nor U25941 (N_25941,N_24247,N_23303);
or U25942 (N_25942,N_20303,N_22691);
nor U25943 (N_25943,N_20324,N_20359);
nor U25944 (N_25944,N_22379,N_21455);
and U25945 (N_25945,N_21859,N_21366);
and U25946 (N_25946,N_24536,N_20525);
or U25947 (N_25947,N_21385,N_23259);
or U25948 (N_25948,N_20704,N_24230);
nand U25949 (N_25949,N_24024,N_23706);
or U25950 (N_25950,N_22783,N_22924);
and U25951 (N_25951,N_22366,N_24464);
nand U25952 (N_25952,N_24245,N_24168);
or U25953 (N_25953,N_21162,N_24936);
and U25954 (N_25954,N_20115,N_24998);
and U25955 (N_25955,N_20912,N_22565);
nand U25956 (N_25956,N_24585,N_21619);
or U25957 (N_25957,N_23110,N_22541);
nand U25958 (N_25958,N_24195,N_23428);
xnor U25959 (N_25959,N_20858,N_21919);
and U25960 (N_25960,N_20388,N_23307);
nor U25961 (N_25961,N_22313,N_23702);
nor U25962 (N_25962,N_22127,N_24657);
nor U25963 (N_25963,N_23801,N_21532);
or U25964 (N_25964,N_23905,N_22435);
nand U25965 (N_25965,N_20585,N_23366);
nor U25966 (N_25966,N_23638,N_22613);
and U25967 (N_25967,N_23750,N_23922);
and U25968 (N_25968,N_22836,N_24099);
nand U25969 (N_25969,N_20726,N_22531);
or U25970 (N_25970,N_20941,N_21282);
nand U25971 (N_25971,N_20633,N_21788);
or U25972 (N_25972,N_22279,N_24496);
nor U25973 (N_25973,N_23165,N_21148);
nand U25974 (N_25974,N_20470,N_23070);
nor U25975 (N_25975,N_24029,N_23654);
or U25976 (N_25976,N_23450,N_22364);
and U25977 (N_25977,N_22521,N_20797);
xor U25978 (N_25978,N_22078,N_20828);
xor U25979 (N_25979,N_23723,N_23135);
xor U25980 (N_25980,N_22632,N_22736);
and U25981 (N_25981,N_24688,N_23828);
nor U25982 (N_25982,N_22023,N_20581);
and U25983 (N_25983,N_24357,N_23470);
and U25984 (N_25984,N_24208,N_22774);
nand U25985 (N_25985,N_21956,N_22536);
or U25986 (N_25986,N_20742,N_20427);
xnor U25987 (N_25987,N_20715,N_22925);
nand U25988 (N_25988,N_24112,N_24372);
nand U25989 (N_25989,N_21187,N_23849);
nand U25990 (N_25990,N_21507,N_22681);
nor U25991 (N_25991,N_22532,N_20506);
nand U25992 (N_25992,N_21395,N_23040);
or U25993 (N_25993,N_23837,N_24708);
xnor U25994 (N_25994,N_21355,N_20325);
nand U25995 (N_25995,N_24661,N_21639);
nand U25996 (N_25996,N_20154,N_23297);
and U25997 (N_25997,N_24914,N_21825);
nand U25998 (N_25998,N_22124,N_23567);
nor U25999 (N_25999,N_24343,N_21122);
nand U26000 (N_26000,N_23914,N_21869);
or U26001 (N_26001,N_20043,N_22602);
nand U26002 (N_26002,N_24217,N_24430);
nor U26003 (N_26003,N_22139,N_23713);
nor U26004 (N_26004,N_23547,N_22021);
and U26005 (N_26005,N_21402,N_23272);
and U26006 (N_26006,N_23981,N_22809);
and U26007 (N_26007,N_22991,N_24327);
and U26008 (N_26008,N_21344,N_24329);
and U26009 (N_26009,N_23872,N_21468);
nor U26010 (N_26010,N_22246,N_23814);
or U26011 (N_26011,N_21042,N_23369);
nor U26012 (N_26012,N_20060,N_22086);
nand U26013 (N_26013,N_24442,N_22439);
or U26014 (N_26014,N_22493,N_20888);
and U26015 (N_26015,N_21398,N_22033);
and U26016 (N_26016,N_20942,N_24977);
nor U26017 (N_26017,N_22314,N_22338);
and U26018 (N_26018,N_22616,N_23740);
nand U26019 (N_26019,N_24058,N_20438);
nand U26020 (N_26020,N_20496,N_22659);
nand U26021 (N_26021,N_20247,N_22718);
nor U26022 (N_26022,N_21891,N_24614);
nor U26023 (N_26023,N_24316,N_20313);
nor U26024 (N_26024,N_24262,N_21803);
nor U26025 (N_26025,N_21526,N_21678);
xor U26026 (N_26026,N_23282,N_22420);
nand U26027 (N_26027,N_21172,N_21697);
xor U26028 (N_26028,N_20939,N_23075);
and U26029 (N_26029,N_23540,N_23381);
or U26030 (N_26030,N_20133,N_23856);
nor U26031 (N_26031,N_20389,N_24336);
and U26032 (N_26032,N_23645,N_24837);
or U26033 (N_26033,N_21234,N_20643);
nor U26034 (N_26034,N_21649,N_24237);
or U26035 (N_26035,N_21873,N_20180);
nand U26036 (N_26036,N_22705,N_23062);
or U26037 (N_26037,N_22044,N_23340);
or U26038 (N_26038,N_23263,N_22098);
nand U26039 (N_26039,N_20345,N_20093);
and U26040 (N_26040,N_22952,N_24529);
or U26041 (N_26041,N_24578,N_22966);
nand U26042 (N_26042,N_24781,N_24137);
nor U26043 (N_26043,N_24489,N_21743);
nor U26044 (N_26044,N_21598,N_24828);
nor U26045 (N_26045,N_22796,N_20640);
nand U26046 (N_26046,N_20533,N_23675);
or U26047 (N_26047,N_21297,N_21278);
or U26048 (N_26048,N_22016,N_24917);
nand U26049 (N_26049,N_21272,N_23364);
nor U26050 (N_26050,N_20018,N_23191);
or U26051 (N_26051,N_23733,N_24018);
or U26052 (N_26052,N_24571,N_20765);
xor U26053 (N_26053,N_21481,N_22592);
or U26054 (N_26054,N_22120,N_22106);
nand U26055 (N_26055,N_22537,N_20930);
xor U26056 (N_26056,N_24982,N_23144);
xnor U26057 (N_26057,N_21372,N_20758);
nand U26058 (N_26058,N_22378,N_20317);
nand U26059 (N_26059,N_23923,N_21949);
nor U26060 (N_26060,N_22446,N_23970);
or U26061 (N_26061,N_24243,N_22409);
nor U26062 (N_26062,N_24492,N_23806);
nor U26063 (N_26063,N_21975,N_22968);
nor U26064 (N_26064,N_20197,N_20193);
or U26065 (N_26065,N_23039,N_23029);
nor U26066 (N_26066,N_23530,N_21879);
nor U26067 (N_26067,N_22629,N_20022);
and U26068 (N_26068,N_20332,N_22369);
nor U26069 (N_26069,N_21404,N_20157);
nand U26070 (N_26070,N_21756,N_24547);
or U26071 (N_26071,N_23620,N_20095);
xnor U26072 (N_26072,N_23431,N_20512);
or U26073 (N_26073,N_23377,N_22601);
or U26074 (N_26074,N_20550,N_23947);
nor U26075 (N_26075,N_22451,N_24985);
xnor U26076 (N_26076,N_22881,N_24756);
nor U26077 (N_26077,N_20010,N_24619);
xnor U26078 (N_26078,N_23556,N_21928);
or U26079 (N_26079,N_22815,N_23305);
and U26080 (N_26080,N_21380,N_24809);
or U26081 (N_26081,N_24586,N_23935);
or U26082 (N_26082,N_24364,N_21251);
and U26083 (N_26083,N_24059,N_22229);
nand U26084 (N_26084,N_21827,N_21192);
nor U26085 (N_26085,N_23701,N_22032);
nor U26086 (N_26086,N_22024,N_21952);
nor U26087 (N_26087,N_21736,N_20570);
xor U26088 (N_26088,N_24403,N_20895);
nor U26089 (N_26089,N_20162,N_24461);
or U26090 (N_26090,N_20889,N_22245);
nor U26091 (N_26091,N_23158,N_24173);
or U26092 (N_26092,N_21905,N_22322);
or U26093 (N_26093,N_21171,N_22892);
xor U26094 (N_26094,N_23807,N_22462);
or U26095 (N_26095,N_23881,N_23204);
xor U26096 (N_26096,N_21221,N_22463);
and U26097 (N_26097,N_20047,N_22038);
nor U26098 (N_26098,N_20368,N_23846);
nand U26099 (N_26099,N_23779,N_24054);
xnor U26100 (N_26100,N_23136,N_24975);
or U26101 (N_26101,N_21615,N_22289);
and U26102 (N_26102,N_24944,N_20946);
nor U26103 (N_26103,N_23343,N_20738);
nor U26104 (N_26104,N_21173,N_21543);
or U26105 (N_26105,N_21772,N_23127);
and U26106 (N_26106,N_21563,N_23854);
nand U26107 (N_26107,N_24011,N_21160);
and U26108 (N_26108,N_24397,N_21167);
or U26109 (N_26109,N_20031,N_20049);
and U26110 (N_26110,N_23422,N_21651);
or U26111 (N_26111,N_23079,N_24706);
and U26112 (N_26112,N_23015,N_23819);
or U26113 (N_26113,N_22450,N_24086);
nor U26114 (N_26114,N_24157,N_22251);
nand U26115 (N_26115,N_21472,N_23667);
or U26116 (N_26116,N_24960,N_22939);
or U26117 (N_26117,N_22175,N_23154);
and U26118 (N_26118,N_24176,N_22720);
nor U26119 (N_26119,N_21565,N_22226);
nand U26120 (N_26120,N_23357,N_21191);
xor U26121 (N_26121,N_22280,N_21265);
nor U26122 (N_26122,N_24598,N_23943);
nor U26123 (N_26123,N_22914,N_22214);
nor U26124 (N_26124,N_21327,N_21636);
and U26125 (N_26125,N_22609,N_23888);
nand U26126 (N_26126,N_20336,N_23255);
nand U26127 (N_26127,N_24411,N_20396);
nand U26128 (N_26128,N_22494,N_24455);
and U26129 (N_26129,N_22277,N_24082);
nor U26130 (N_26130,N_20754,N_23277);
nor U26131 (N_26131,N_24815,N_23503);
and U26132 (N_26132,N_21954,N_23292);
and U26133 (N_26133,N_22904,N_20877);
xnor U26134 (N_26134,N_24607,N_23054);
or U26135 (N_26135,N_21795,N_23193);
nand U26136 (N_26136,N_22402,N_20283);
nand U26137 (N_26137,N_22806,N_22308);
xor U26138 (N_26138,N_23612,N_21493);
and U26139 (N_26139,N_24330,N_20725);
xor U26140 (N_26140,N_21773,N_20543);
and U26141 (N_26141,N_22035,N_21457);
and U26142 (N_26142,N_23820,N_21944);
nand U26143 (N_26143,N_22857,N_20915);
and U26144 (N_26144,N_20963,N_20920);
nor U26145 (N_26145,N_22618,N_22823);
nor U26146 (N_26146,N_20564,N_23817);
and U26147 (N_26147,N_24672,N_23212);
or U26148 (N_26148,N_20565,N_20814);
nand U26149 (N_26149,N_20161,N_21633);
nand U26150 (N_26150,N_22427,N_22886);
or U26151 (N_26151,N_20851,N_22149);
and U26152 (N_26152,N_20495,N_23797);
xor U26153 (N_26153,N_23001,N_21465);
nand U26154 (N_26154,N_21256,N_24321);
and U26155 (N_26155,N_20668,N_22404);
or U26156 (N_26156,N_20753,N_21711);
xnor U26157 (N_26157,N_20799,N_20113);
and U26158 (N_26158,N_22548,N_20080);
nand U26159 (N_26159,N_24069,N_21955);
and U26160 (N_26160,N_21337,N_20693);
nand U26161 (N_26161,N_21964,N_21156);
and U26162 (N_26162,N_23473,N_24887);
nor U26163 (N_26163,N_21194,N_21564);
xor U26164 (N_26164,N_21602,N_21830);
nor U26165 (N_26165,N_22132,N_20439);
xor U26166 (N_26166,N_22376,N_24231);
and U26167 (N_26167,N_22793,N_24419);
nor U26168 (N_26168,N_20650,N_21489);
and U26169 (N_26169,N_21005,N_24325);
nor U26170 (N_26170,N_20199,N_23639);
nand U26171 (N_26171,N_24429,N_20974);
nand U26172 (N_26172,N_23672,N_21841);
nand U26173 (N_26173,N_23439,N_21201);
and U26174 (N_26174,N_20825,N_20483);
and U26175 (N_26175,N_21271,N_21094);
and U26176 (N_26176,N_22526,N_24201);
and U26177 (N_26177,N_22111,N_22169);
and U26178 (N_26178,N_20228,N_24445);
nand U26179 (N_26179,N_21161,N_24652);
or U26180 (N_26180,N_20644,N_24651);
nor U26181 (N_26181,N_23076,N_21936);
nand U26182 (N_26182,N_23652,N_23571);
nor U26183 (N_26183,N_20882,N_20687);
and U26184 (N_26184,N_20415,N_22146);
xor U26185 (N_26185,N_20126,N_23395);
nand U26186 (N_26186,N_24617,N_21572);
nand U26187 (N_26187,N_21870,N_23942);
or U26188 (N_26188,N_20535,N_21145);
or U26189 (N_26189,N_23758,N_20484);
nand U26190 (N_26190,N_23958,N_23583);
nor U26191 (N_26191,N_21887,N_22034);
or U26192 (N_26192,N_23791,N_21289);
nand U26193 (N_26193,N_20537,N_23229);
nand U26194 (N_26194,N_24626,N_24811);
nand U26195 (N_26195,N_22764,N_23537);
or U26196 (N_26196,N_24160,N_20376);
nand U26197 (N_26197,N_20437,N_22910);
and U26198 (N_26198,N_23107,N_22527);
and U26199 (N_26199,N_24246,N_22223);
nor U26200 (N_26200,N_22637,N_22476);
nand U26201 (N_26201,N_24722,N_21603);
nor U26202 (N_26202,N_24874,N_22118);
or U26203 (N_26203,N_20085,N_24867);
xor U26204 (N_26204,N_20110,N_21239);
and U26205 (N_26205,N_21490,N_22780);
or U26206 (N_26206,N_23499,N_24819);
and U26207 (N_26207,N_22352,N_23657);
nor U26208 (N_26208,N_22589,N_22456);
nand U26209 (N_26209,N_23371,N_23631);
nand U26210 (N_26210,N_24260,N_23038);
or U26211 (N_26211,N_23707,N_20676);
or U26212 (N_26212,N_22697,N_22802);
nor U26213 (N_26213,N_22860,N_23712);
or U26214 (N_26214,N_24304,N_24440);
and U26215 (N_26215,N_21002,N_20471);
nor U26216 (N_26216,N_20589,N_21826);
or U26217 (N_26217,N_20414,N_20393);
xor U26218 (N_26218,N_22967,N_23629);
nor U26219 (N_26219,N_20558,N_22787);
xnor U26220 (N_26220,N_22331,N_22255);
or U26221 (N_26221,N_22037,N_24899);
or U26222 (N_26222,N_22665,N_24474);
nor U26223 (N_26223,N_20868,N_22650);
or U26224 (N_26224,N_21548,N_21458);
nor U26225 (N_26225,N_23633,N_23975);
nor U26226 (N_26226,N_22789,N_23406);
and U26227 (N_26227,N_21714,N_23246);
nand U26228 (N_26228,N_20805,N_24558);
nor U26229 (N_26229,N_24548,N_21046);
nor U26230 (N_26230,N_22856,N_24517);
and U26231 (N_26231,N_21541,N_24040);
and U26232 (N_26232,N_21477,N_23591);
nor U26233 (N_26233,N_22466,N_20789);
and U26234 (N_26234,N_22546,N_20374);
nand U26235 (N_26235,N_22923,N_21580);
xor U26236 (N_26236,N_20597,N_23714);
or U26237 (N_26237,N_21828,N_22184);
xnor U26238 (N_26238,N_20298,N_23018);
nand U26239 (N_26239,N_23610,N_24215);
or U26240 (N_26240,N_23004,N_23578);
nand U26241 (N_26241,N_23095,N_24644);
and U26242 (N_26242,N_21857,N_21294);
nor U26243 (N_26243,N_21314,N_21848);
nor U26244 (N_26244,N_21961,N_20221);
and U26245 (N_26245,N_23150,N_23306);
or U26246 (N_26246,N_20529,N_21833);
or U26247 (N_26247,N_24132,N_21099);
nor U26248 (N_26248,N_24841,N_22989);
nor U26249 (N_26249,N_22400,N_24825);
and U26250 (N_26250,N_24590,N_20766);
and U26251 (N_26251,N_21389,N_20970);
nand U26252 (N_26252,N_23680,N_21086);
or U26253 (N_26253,N_21943,N_24790);
xnor U26254 (N_26254,N_23569,N_22574);
and U26255 (N_26255,N_24865,N_24408);
or U26256 (N_26256,N_24319,N_20291);
nor U26257 (N_26257,N_24133,N_22203);
nand U26258 (N_26258,N_20955,N_20832);
nor U26259 (N_26259,N_23201,N_23647);
xor U26260 (N_26260,N_23884,N_21709);
and U26261 (N_26261,N_24182,N_21524);
nand U26262 (N_26262,N_21729,N_22291);
and U26263 (N_26263,N_24592,N_21390);
or U26264 (N_26264,N_24005,N_21116);
nor U26265 (N_26265,N_22218,N_21696);
xor U26266 (N_26266,N_24462,N_20831);
nand U26267 (N_26267,N_20848,N_23455);
xnor U26268 (N_26268,N_22788,N_23968);
or U26269 (N_26269,N_20624,N_20574);
nand U26270 (N_26270,N_20411,N_20544);
nor U26271 (N_26271,N_22179,N_22840);
and U26272 (N_26272,N_23648,N_21703);
nand U26273 (N_26273,N_24039,N_23210);
and U26274 (N_26274,N_24169,N_24261);
nand U26275 (N_26275,N_21415,N_20434);
or U26276 (N_26276,N_22042,N_23661);
and U26277 (N_26277,N_21168,N_24502);
nor U26278 (N_26278,N_20890,N_22383);
or U26279 (N_26279,N_23765,N_22256);
or U26280 (N_26280,N_20566,N_23490);
nor U26281 (N_26281,N_23529,N_24976);
or U26282 (N_26282,N_24989,N_24750);
nand U26283 (N_26283,N_22220,N_21470);
and U26284 (N_26284,N_23731,N_22662);
and U26285 (N_26285,N_22606,N_20280);
and U26286 (N_26286,N_21810,N_22701);
nor U26287 (N_26287,N_21719,N_23684);
xnor U26288 (N_26288,N_23456,N_21303);
or U26289 (N_26289,N_22564,N_24686);
and U26290 (N_26290,N_23649,N_23682);
and U26291 (N_26291,N_23867,N_23236);
and U26292 (N_26292,N_23378,N_24973);
nand U26293 (N_26293,N_22444,N_22361);
and U26294 (N_26294,N_20163,N_20164);
or U26295 (N_26295,N_22571,N_24265);
nor U26296 (N_26296,N_23243,N_22999);
nand U26297 (N_26297,N_21860,N_20403);
or U26298 (N_26298,N_24097,N_20456);
nor U26299 (N_26299,N_22365,N_24102);
nand U26300 (N_26300,N_21206,N_24728);
or U26301 (N_26301,N_24289,N_20184);
nand U26302 (N_26302,N_21738,N_23288);
and U26303 (N_26303,N_23437,N_20580);
xnor U26304 (N_26304,N_21966,N_22061);
and U26305 (N_26305,N_22837,N_20829);
xor U26306 (N_26306,N_23315,N_21958);
or U26307 (N_26307,N_20204,N_22633);
nor U26308 (N_26308,N_21595,N_20297);
nand U26309 (N_26309,N_22443,N_23022);
or U26310 (N_26310,N_23026,N_23200);
and U26311 (N_26311,N_22756,N_24075);
xnor U26312 (N_26312,N_20683,N_20539);
xnor U26313 (N_26313,N_23960,N_23717);
xor U26314 (N_26314,N_23677,N_23842);
xor U26315 (N_26315,N_21868,N_24563);
nand U26316 (N_26316,N_21064,N_23531);
nor U26317 (N_26317,N_22988,N_22090);
nor U26318 (N_26318,N_22103,N_21989);
nand U26319 (N_26319,N_20670,N_24056);
xor U26320 (N_26320,N_20114,N_24263);
nor U26321 (N_26321,N_21538,N_21196);
nor U26322 (N_26322,N_22797,N_23589);
or U26323 (N_26323,N_24465,N_21577);
xor U26324 (N_26324,N_21129,N_21213);
nor U26325 (N_26325,N_21216,N_20874);
nand U26326 (N_26326,N_20515,N_22454);
or U26327 (N_26327,N_24488,N_24624);
or U26328 (N_26328,N_23562,N_22880);
and U26329 (N_26329,N_23678,N_24153);
nand U26330 (N_26330,N_23893,N_23694);
xor U26331 (N_26331,N_24608,N_24864);
nor U26332 (N_26332,N_21984,N_20037);
nand U26333 (N_26333,N_24711,N_23403);
nand U26334 (N_26334,N_21530,N_20144);
nand U26335 (N_26335,N_21096,N_22377);
and U26336 (N_26336,N_24747,N_22905);
or U26337 (N_26337,N_22894,N_21948);
nor U26338 (N_26338,N_23031,N_21246);
or U26339 (N_26339,N_22492,N_21590);
or U26340 (N_26340,N_20919,N_20845);
nand U26341 (N_26341,N_24987,N_23360);
or U26342 (N_26342,N_20223,N_21583);
or U26343 (N_26343,N_21679,N_21197);
and U26344 (N_26344,N_21360,N_23161);
or U26345 (N_26345,N_24037,N_23084);
xor U26346 (N_26346,N_20620,N_23767);
and U26347 (N_26347,N_20734,N_20373);
and U26348 (N_26348,N_24036,N_21087);
nand U26349 (N_26349,N_20583,N_23690);
and U26350 (N_26350,N_20588,N_22166);
nand U26351 (N_26351,N_20337,N_23139);
nor U26352 (N_26352,N_21518,N_23927);
or U26353 (N_26353,N_20910,N_24475);
nor U26354 (N_26354,N_21178,N_22664);
or U26355 (N_26355,N_23915,N_21593);
nand U26356 (N_26356,N_23221,N_24306);
or U26357 (N_26357,N_23088,N_23575);
or U26358 (N_26358,N_24953,N_23353);
xnor U26359 (N_26359,N_20551,N_22641);
nand U26360 (N_26360,N_21820,N_22210);
xor U26361 (N_26361,N_21183,N_24731);
nor U26362 (N_26362,N_23155,N_21762);
nand U26363 (N_26363,N_21778,N_22872);
and U26364 (N_26364,N_21077,N_20658);
nor U26365 (N_26365,N_22097,N_23129);
and U26366 (N_26366,N_24540,N_24832);
nor U26367 (N_26367,N_23044,N_21630);
or U26368 (N_26368,N_20421,N_23157);
nor U26369 (N_26369,N_23933,N_23697);
xnor U26370 (N_26370,N_23594,N_24487);
nor U26371 (N_26371,N_22471,N_23216);
nor U26372 (N_26372,N_22811,N_23228);
nand U26373 (N_26373,N_24311,N_24358);
and U26374 (N_26374,N_23501,N_24207);
nor U26375 (N_26375,N_21222,N_20430);
xor U26376 (N_26376,N_20425,N_21114);
nand U26377 (N_26377,N_21876,N_21075);
xnor U26378 (N_26378,N_21381,N_24062);
or U26379 (N_26379,N_24308,N_23572);
nand U26380 (N_26380,N_24892,N_21408);
and U26381 (N_26381,N_22628,N_20631);
nand U26382 (N_26382,N_23634,N_22518);
nand U26383 (N_26383,N_21699,N_22733);
or U26384 (N_26384,N_23123,N_20592);
nor U26385 (N_26385,N_22773,N_22762);
or U26386 (N_26386,N_20075,N_24257);
nor U26387 (N_26387,N_21797,N_20703);
nor U26388 (N_26388,N_22678,N_23868);
nor U26389 (N_26389,N_20188,N_24904);
and U26390 (N_26390,N_24631,N_20498);
and U26391 (N_26391,N_20914,N_21749);
and U26392 (N_26392,N_22031,N_21439);
and U26393 (N_26393,N_21838,N_24682);
nand U26394 (N_26394,N_21533,N_23049);
nor U26395 (N_26395,N_23367,N_21238);
nor U26396 (N_26396,N_20129,N_21644);
nor U26397 (N_26397,N_24727,N_22017);
xor U26398 (N_26398,N_21388,N_20876);
or U26399 (N_26399,N_20346,N_22906);
nor U26400 (N_26400,N_20680,N_21448);
nand U26401 (N_26401,N_24042,N_20140);
or U26402 (N_26402,N_20932,N_21508);
nand U26403 (N_26403,N_24315,N_23410);
nor U26404 (N_26404,N_21134,N_24469);
or U26405 (N_26405,N_23559,N_20775);
nor U26406 (N_26406,N_20141,N_21371);
nor U26407 (N_26407,N_23911,N_22206);
xor U26408 (N_26408,N_21753,N_20918);
nor U26409 (N_26409,N_20187,N_20702);
nor U26410 (N_26410,N_23234,N_24407);
nor U26411 (N_26411,N_23209,N_24285);
and U26412 (N_26412,N_20770,N_22323);
nand U26413 (N_26413,N_23316,N_23573);
and U26414 (N_26414,N_24535,N_23260);
or U26415 (N_26415,N_21976,N_24684);
xor U26416 (N_26416,N_24642,N_21855);
nor U26417 (N_26417,N_23203,N_24765);
or U26418 (N_26418,N_22522,N_24593);
nor U26419 (N_26419,N_23153,N_20601);
or U26420 (N_26420,N_20747,N_22221);
xor U26421 (N_26421,N_24113,N_23670);
nand U26422 (N_26422,N_23891,N_21912);
nor U26423 (N_26423,N_23214,N_20736);
nand U26424 (N_26424,N_24100,N_23223);
and U26425 (N_26425,N_22375,N_22405);
and U26426 (N_26426,N_23716,N_24660);
or U26427 (N_26427,N_23794,N_24250);
or U26428 (N_26428,N_23857,N_20118);
and U26429 (N_26429,N_21150,N_21994);
or U26430 (N_26430,N_21535,N_23465);
nand U26431 (N_26431,N_20127,N_21872);
nor U26432 (N_26432,N_21263,N_23256);
xor U26433 (N_26433,N_20646,N_22351);
and U26434 (N_26434,N_22440,N_22846);
or U26435 (N_26435,N_21917,N_20195);
nor U26436 (N_26436,N_24927,N_21254);
nor U26437 (N_26437,N_20108,N_23761);
and U26438 (N_26438,N_21198,N_24613);
and U26439 (N_26439,N_22612,N_24858);
nand U26440 (N_26440,N_24733,N_24471);
nand U26441 (N_26441,N_20791,N_20913);
nor U26442 (N_26442,N_22640,N_24339);
xnor U26443 (N_26443,N_23528,N_20841);
nand U26444 (N_26444,N_23616,N_22370);
nor U26445 (N_26445,N_24413,N_21024);
nor U26446 (N_26446,N_20856,N_22200);
and U26447 (N_26447,N_24228,N_22599);
and U26448 (N_26448,N_23936,N_23892);
or U26449 (N_26449,N_22232,N_21574);
nor U26450 (N_26450,N_21479,N_24941);
xnor U26451 (N_26451,N_22918,N_20227);
and U26452 (N_26452,N_23957,N_23990);
nand U26453 (N_26453,N_20967,N_20241);
nand U26454 (N_26454,N_21981,N_22882);
nand U26455 (N_26455,N_20582,N_20238);
or U26456 (N_26456,N_20519,N_22673);
nand U26457 (N_26457,N_24738,N_20194);
and U26458 (N_26458,N_20011,N_22028);
or U26459 (N_26459,N_20522,N_22597);
nor U26460 (N_26460,N_23551,N_24003);
or U26461 (N_26461,N_21892,N_24117);
or U26462 (N_26462,N_22871,N_22319);
and U26463 (N_26463,N_21275,N_24320);
nand U26464 (N_26464,N_21165,N_23036);
or U26465 (N_26465,N_22247,N_23073);
or U26466 (N_26466,N_20901,N_23602);
nand U26467 (N_26467,N_24221,N_24337);
or U26468 (N_26468,N_22171,N_20626);
or U26469 (N_26469,N_24808,N_21775);
nand U26470 (N_26470,N_23338,N_23980);
and U26471 (N_26471,N_21127,N_22190);
nand U26472 (N_26472,N_21812,N_22270);
nor U26473 (N_26473,N_24916,N_24562);
nand U26474 (N_26474,N_24883,N_21569);
or U26475 (N_26475,N_24338,N_24942);
nor U26476 (N_26476,N_21845,N_20559);
nor U26477 (N_26477,N_24444,N_20045);
and U26478 (N_26478,N_23329,N_23681);
nand U26479 (N_26479,N_21652,N_21210);
and U26480 (N_26480,N_22960,N_20240);
nand U26481 (N_26481,N_20743,N_24349);
nor U26482 (N_26482,N_24734,N_24902);
nand U26483 (N_26483,N_22915,N_23230);
xnor U26484 (N_26484,N_21462,N_24962);
nand U26485 (N_26485,N_24542,N_20663);
nand U26486 (N_26486,N_22161,N_20648);
and U26487 (N_26487,N_21596,N_23000);
or U26488 (N_26488,N_24374,N_23217);
nor U26489 (N_26489,N_22045,N_22687);
nor U26490 (N_26490,N_21243,N_24332);
or U26491 (N_26491,N_20446,N_20767);
nor U26492 (N_26492,N_23630,N_23637);
xnor U26493 (N_26493,N_23310,N_23098);
or U26494 (N_26494,N_21608,N_22604);
nor U26495 (N_26495,N_20896,N_24833);
nor U26496 (N_26496,N_22242,N_20273);
or U26497 (N_26497,N_20660,N_24191);
nor U26498 (N_26498,N_24156,N_20282);
nor U26499 (N_26499,N_20517,N_23802);
or U26500 (N_26500,N_22666,N_21740);
or U26501 (N_26501,N_23969,N_23772);
xor U26502 (N_26502,N_21175,N_24820);
nand U26503 (N_26503,N_24844,N_20083);
nand U26504 (N_26504,N_24006,N_24234);
or U26505 (N_26505,N_20824,N_21025);
or U26506 (N_26506,N_22849,N_23780);
and U26507 (N_26507,N_20196,N_24435);
nor U26508 (N_26508,N_20820,N_23615);
nand U26509 (N_26509,N_20835,N_21317);
xor U26510 (N_26510,N_21987,N_22081);
and U26511 (N_26511,N_20121,N_21358);
xnor U26512 (N_26512,N_20981,N_24206);
nor U26513 (N_26513,N_21588,N_24971);
and U26514 (N_26514,N_21897,N_21931);
and U26515 (N_26515,N_23266,N_24555);
or U26516 (N_26516,N_20117,N_24092);
nand U26517 (N_26517,N_22264,N_24922);
or U26518 (N_26518,N_20285,N_22362);
or U26519 (N_26519,N_24771,N_21909);
nor U26520 (N_26520,N_24845,N_23887);
and U26521 (N_26521,N_24920,N_22213);
xnor U26522 (N_26522,N_20258,N_22985);
or U26523 (N_26523,N_20729,N_23405);
or U26524 (N_26524,N_22276,N_21992);
nor U26525 (N_26525,N_21760,N_20153);
xor U26526 (N_26526,N_22235,N_23600);
xnor U26527 (N_26527,N_21318,N_23961);
and U26528 (N_26528,N_22423,N_21628);
or U26529 (N_26529,N_21519,N_24951);
nor U26530 (N_26530,N_22660,N_23994);
nand U26531 (N_26531,N_24051,N_20372);
and U26532 (N_26532,N_20808,N_22043);
nor U26533 (N_26533,N_20718,N_20613);
and U26534 (N_26534,N_20104,N_22133);
nand U26535 (N_26535,N_23339,N_23879);
nand U26536 (N_26536,N_24823,N_21578);
and U26537 (N_26537,N_22134,N_23421);
nand U26538 (N_26538,N_21396,N_24705);
nor U26539 (N_26539,N_24560,N_20277);
and U26540 (N_26540,N_24676,N_20746);
nand U26541 (N_26541,N_24021,N_24202);
or U26542 (N_26542,N_23014,N_22014);
nor U26543 (N_26543,N_23515,N_21785);
or U26544 (N_26544,N_23238,N_20629);
and U26545 (N_26545,N_23844,N_20096);
nor U26546 (N_26546,N_24341,N_23815);
nor U26547 (N_26547,N_21621,N_21707);
and U26548 (N_26548,N_24264,N_21640);
or U26549 (N_26549,N_21692,N_24516);
or U26550 (N_26550,N_23997,N_21926);
nand U26551 (N_26551,N_21245,N_22677);
nor U26552 (N_26552,N_20290,N_23458);
or U26553 (N_26553,N_20823,N_22396);
nand U26554 (N_26554,N_20300,N_22615);
nand U26555 (N_26555,N_21382,N_23725);
and U26556 (N_26556,N_23180,N_23151);
nor U26557 (N_26557,N_21796,N_20723);
nor U26558 (N_26558,N_20296,N_20571);
nand U26559 (N_26559,N_20383,N_22543);
nand U26560 (N_26560,N_22500,N_21765);
nand U26561 (N_26561,N_23607,N_20929);
nor U26562 (N_26562,N_23103,N_24645);
nor U26563 (N_26563,N_22348,N_24910);
xnor U26564 (N_26564,N_20354,N_20119);
nand U26565 (N_26565,N_21320,N_24368);
xor U26566 (N_26566,N_23775,N_20177);
nor U26567 (N_26567,N_22737,N_22170);
nor U26568 (N_26568,N_23863,N_22786);
and U26569 (N_26569,N_24567,N_22325);
nor U26570 (N_26570,N_22298,N_24127);
and U26571 (N_26571,N_20444,N_22657);
or U26572 (N_26572,N_23183,N_21368);
and U26573 (N_26573,N_20993,N_21146);
or U26574 (N_26574,N_21613,N_22930);
nor U26575 (N_26575,N_21324,N_21585);
nor U26576 (N_26576,N_21349,N_23222);
xnor U26577 (N_26577,N_22064,N_20810);
or U26578 (N_26578,N_20891,N_21407);
or U26579 (N_26579,N_22126,N_22996);
and U26580 (N_26580,N_20875,N_21417);
or U26581 (N_26581,N_23902,N_21549);
nand U26582 (N_26582,N_22344,N_21957);
or U26583 (N_26583,N_24697,N_23089);
nand U26584 (N_26584,N_20326,N_20168);
or U26585 (N_26585,N_20304,N_21685);
nor U26586 (N_26586,N_22473,N_22060);
nand U26587 (N_26587,N_24020,N_24175);
or U26588 (N_26588,N_21831,N_20226);
nor U26589 (N_26589,N_20612,N_24994);
or U26590 (N_26590,N_20033,N_24269);
or U26591 (N_26591,N_23870,N_22575);
nor U26592 (N_26592,N_21123,N_24881);
nor U26593 (N_26593,N_23207,N_21095);
nand U26594 (N_26594,N_20489,N_21483);
nand U26595 (N_26595,N_20342,N_22903);
nand U26596 (N_26596,N_20632,N_20287);
and U26597 (N_26597,N_23988,N_21698);
or U26598 (N_26598,N_20853,N_21007);
nand U26599 (N_26599,N_24658,N_23083);
nor U26600 (N_26600,N_22873,N_22855);
nand U26601 (N_26601,N_20727,N_23090);
xor U26602 (N_26602,N_22513,N_21520);
xnor U26603 (N_26603,N_21103,N_22056);
nand U26604 (N_26604,N_23006,N_22698);
nand U26605 (N_26605,N_24690,N_20398);
or U26606 (N_26606,N_24744,N_21784);
and U26607 (N_26607,N_21013,N_20936);
nor U26608 (N_26608,N_21606,N_20988);
nand U26609 (N_26609,N_22588,N_22363);
nand U26610 (N_26610,N_22254,N_24760);
nor U26611 (N_26611,N_21635,N_20299);
and U26612 (N_26612,N_20973,N_21281);
and U26613 (N_26613,N_23053,N_22944);
nand U26614 (N_26614,N_22114,N_23916);
nand U26615 (N_26615,N_20898,N_20040);
and U26616 (N_26616,N_23673,N_24641);
xor U26617 (N_26617,N_21359,N_22828);
nand U26618 (N_26618,N_23739,N_24486);
or U26619 (N_26619,N_24293,N_24817);
xnor U26620 (N_26620,N_24979,N_24943);
nor U26621 (N_26621,N_23279,N_21768);
xor U26622 (N_26622,N_21176,N_20768);
or U26623 (N_26623,N_21560,N_21609);
nand U26624 (N_26624,N_22233,N_22539);
and U26625 (N_26625,N_24634,N_20412);
or U26626 (N_26626,N_23810,N_24423);
nor U26627 (N_26627,N_20253,N_24449);
nor U26628 (N_26628,N_22350,N_24868);
and U26629 (N_26629,N_24584,N_22491);
nor U26630 (N_26630,N_22829,N_20493);
or U26631 (N_26631,N_21467,N_22715);
nor U26632 (N_26632,N_22496,N_24066);
or U26633 (N_26633,N_23955,N_21937);
xnor U26634 (N_26634,N_22437,N_21258);
xor U26635 (N_26635,N_22775,N_22883);
or U26636 (N_26636,N_24209,N_22810);
or U26637 (N_26637,N_23993,N_21528);
nor U26638 (N_26638,N_20816,N_21741);
nor U26639 (N_26639,N_22639,N_24240);
xnor U26640 (N_26640,N_22895,N_21236);
or U26641 (N_26641,N_23511,N_20281);
nor U26642 (N_26642,N_22188,N_24235);
xnor U26643 (N_26643,N_24183,N_24839);
xor U26644 (N_26644,N_22813,N_24745);
or U26645 (N_26645,N_23130,N_24580);
or U26646 (N_26646,N_23796,N_21668);
or U26647 (N_26647,N_24398,N_20700);
nor U26648 (N_26648,N_20027,N_24232);
and U26649 (N_26649,N_21566,N_22312);
nor U26650 (N_26650,N_23756,N_22743);
nand U26651 (N_26651,N_23721,N_23776);
nor U26652 (N_26652,N_20917,N_22453);
or U26653 (N_26653,N_22065,N_21416);
and U26654 (N_26654,N_21058,N_20567);
and U26655 (N_26655,N_24978,N_20418);
nand U26656 (N_26656,N_23691,N_21330);
nor U26657 (N_26657,N_24439,N_21063);
nand U26658 (N_26658,N_24522,N_22777);
nor U26659 (N_26659,N_20971,N_20505);
and U26660 (N_26660,N_23904,N_21276);
or U26661 (N_26661,N_22157,N_22142);
or U26662 (N_26662,N_23418,N_24361);
nand U26663 (N_26663,N_22216,N_20903);
nor U26664 (N_26664,N_23432,N_21350);
or U26665 (N_26665,N_23227,N_23284);
and U26666 (N_26666,N_23865,N_23862);
nor U26667 (N_26667,N_20449,N_20064);
xnor U26668 (N_26668,N_21713,N_24362);
nor U26669 (N_26669,N_24387,N_24655);
xor U26670 (N_26670,N_23517,N_20985);
nand U26671 (N_26671,N_21177,N_23425);
nor U26672 (N_26672,N_24292,N_22049);
or U26673 (N_26673,N_22085,N_20604);
or U26674 (N_26674,N_24267,N_24773);
and U26675 (N_26675,N_24519,N_23687);
nor U26676 (N_26676,N_21215,N_20250);
and U26677 (N_26677,N_22695,N_20902);
or U26678 (N_26678,N_24074,N_24393);
xnor U26679 (N_26679,N_22794,N_24395);
nor U26680 (N_26680,N_22819,N_24782);
nor U26681 (N_26681,N_22477,N_20385);
nor U26682 (N_26682,N_23063,N_22649);
nor U26683 (N_26683,N_22108,N_21682);
nand U26684 (N_26684,N_24670,N_22105);
and U26685 (N_26685,N_20674,N_20962);
nand U26686 (N_26686,N_23187,N_20534);
nand U26687 (N_26687,N_22281,N_24485);
nor U26688 (N_26688,N_21055,N_24384);
or U26689 (N_26689,N_21734,N_21049);
and U26690 (N_26690,N_23538,N_24543);
xor U26691 (N_26691,N_20039,N_23826);
xor U26692 (N_26692,N_23581,N_21686);
xnor U26693 (N_26693,N_21523,N_23163);
or U26694 (N_26694,N_22317,N_22484);
nand U26695 (N_26695,N_23774,N_21781);
nor U26696 (N_26696,N_22757,N_20837);
or U26697 (N_26697,N_24616,N_23964);
nand U26698 (N_26698,N_22889,N_22424);
and U26699 (N_26699,N_21599,N_24778);
nand U26700 (N_26700,N_22448,N_20576);
nand U26701 (N_26701,N_23116,N_23699);
nor U26702 (N_26702,N_23565,N_22654);
nor U26703 (N_26703,N_24149,N_21279);
and U26704 (N_26704,N_23361,N_24190);
nor U26705 (N_26705,N_20206,N_23325);
nand U26706 (N_26706,N_20834,N_23321);
nor U26707 (N_26707,N_22865,N_21513);
or U26708 (N_26708,N_24121,N_20691);
or U26709 (N_26709,N_21048,N_22095);
xor U26710 (N_26710,N_21068,N_21287);
or U26711 (N_26711,N_20619,N_22558);
nor U26712 (N_26712,N_22228,N_22645);
or U26713 (N_26713,N_21516,N_20557);
nor U26714 (N_26714,N_22572,N_24347);
and U26715 (N_26715,N_20852,N_22563);
or U26716 (N_26716,N_20511,N_23160);
and U26717 (N_26717,N_24851,N_23326);
or U26718 (N_26718,N_23520,N_22116);
nor U26719 (N_26719,N_23294,N_23025);
or U26720 (N_26720,N_20387,N_21121);
and U26721 (N_26721,N_21307,N_23132);
and U26722 (N_26722,N_21793,N_23376);
or U26723 (N_26723,N_24539,N_22495);
nand U26724 (N_26724,N_21361,N_22258);
nor U26725 (N_26725,N_24526,N_24122);
xor U26726 (N_26726,N_24425,N_23400);
xor U26727 (N_26727,N_21650,N_21960);
or U26728 (N_26728,N_23414,N_20463);
nor U26729 (N_26729,N_24774,N_24822);
nand U26730 (N_26730,N_24022,N_24049);
or U26731 (N_26731,N_20309,N_22130);
nor U26732 (N_26732,N_22885,N_23114);
and U26733 (N_26733,N_20111,N_20737);
xnor U26734 (N_26734,N_22088,N_22333);
or U26735 (N_26735,N_24370,N_21727);
nand U26736 (N_26736,N_23085,N_20641);
nor U26737 (N_26737,N_24467,N_22935);
nand U26738 (N_26738,N_24241,N_20735);
or U26739 (N_26739,N_24574,N_24225);
nor U26740 (N_26740,N_24534,N_21488);
nor U26741 (N_26741,N_22022,N_22399);
or U26742 (N_26742,N_20679,N_23041);
or U26743 (N_26743,N_21232,N_23937);
and U26744 (N_26744,N_22007,N_22516);
and U26745 (N_26745,N_21347,N_20906);
or U26746 (N_26746,N_21700,N_20171);
and U26747 (N_26747,N_24495,N_20087);
nor U26748 (N_26748,N_22557,N_22158);
and U26749 (N_26749,N_22159,N_23931);
nand U26750 (N_26750,N_20069,N_23449);
and U26751 (N_26751,N_22624,N_23642);
nor U26752 (N_26752,N_24866,N_22461);
nor U26753 (N_26753,N_23592,N_20778);
nand U26754 (N_26754,N_23971,N_23548);
nand U26755 (N_26755,N_24283,N_22792);
nand U26756 (N_26756,N_22337,N_22452);
and U26757 (N_26757,N_22716,N_24551);
nor U26758 (N_26758,N_24420,N_20120);
xnor U26759 (N_26759,N_21525,N_22326);
nand U26760 (N_26760,N_22937,N_22071);
xor U26761 (N_26761,N_20980,N_21963);
or U26762 (N_26762,N_23554,N_22980);
nor U26763 (N_26763,N_20473,N_20673);
xor U26764 (N_26764,N_21149,N_23299);
nand U26765 (N_26765,N_22428,N_24854);
xor U26766 (N_26766,N_22241,N_23869);
nand U26767 (N_26767,N_24180,N_24759);
or U26768 (N_26768,N_21486,N_24719);
and U26769 (N_26769,N_21815,N_24862);
nor U26770 (N_26770,N_21888,N_24876);
and U26771 (N_26771,N_20584,N_24569);
and U26772 (N_26772,N_20370,N_22445);
or U26773 (N_26773,N_22290,N_21556);
nand U26774 (N_26774,N_22758,N_21965);
nand U26775 (N_26775,N_20774,N_23064);
and U26776 (N_26776,N_21674,N_21041);
nor U26777 (N_26777,N_22821,N_23487);
xnor U26778 (N_26778,N_22770,N_20350);
or U26779 (N_26779,N_20572,N_20684);
or U26780 (N_26780,N_21118,N_21184);
nor U26781 (N_26781,N_23037,N_23005);
nand U26782 (N_26782,N_20390,N_21435);
nand U26783 (N_26783,N_22552,N_21881);
or U26784 (N_26784,N_22835,N_24905);
or U26785 (N_26785,N_21505,N_24472);
nand U26786 (N_26786,N_22630,N_21319);
nand U26787 (N_26787,N_22092,N_23907);
nand U26788 (N_26788,N_23197,N_23736);
nand U26789 (N_26789,N_20485,N_23374);
nand U26790 (N_26790,N_20105,N_20549);
nand U26791 (N_26791,N_20074,N_24167);
nor U26792 (N_26792,N_23257,N_23258);
nor U26793 (N_26793,N_22119,N_24043);
nor U26794 (N_26794,N_22680,N_21400);
xnor U26795 (N_26795,N_20462,N_22545);
nand U26796 (N_26796,N_22619,N_21223);
xor U26797 (N_26797,N_21939,N_23192);
nor U26798 (N_26798,N_22869,N_21480);
and U26799 (N_26799,N_22578,N_21681);
nor U26800 (N_26800,N_23874,N_23275);
and U26801 (N_26801,N_22535,N_23545);
and U26802 (N_26802,N_21667,N_23460);
and U26803 (N_26803,N_22983,N_21755);
or U26804 (N_26804,N_23541,N_21844);
nor U26805 (N_26805,N_20261,N_24108);
and U26806 (N_26806,N_23510,N_24715);
or U26807 (N_26807,N_24531,N_23664);
or U26808 (N_26808,N_21706,N_20006);
nor U26809 (N_26809,N_20061,N_21907);
nand U26810 (N_26810,N_20361,N_23962);
xor U26811 (N_26811,N_22128,N_21665);
and U26812 (N_26812,N_20318,N_24089);
and U26813 (N_26813,N_23247,N_20063);
or U26814 (N_26814,N_23696,N_23685);
xnor U26815 (N_26815,N_22075,N_20286);
nand U26816 (N_26816,N_21331,N_22706);
nand U26817 (N_26817,N_22551,N_20507);
and U26818 (N_26818,N_24628,N_24352);
or U26819 (N_26819,N_20183,N_20879);
and U26820 (N_26820,N_23231,N_23415);
or U26821 (N_26821,N_22019,N_23798);
or U26822 (N_26822,N_23825,N_24561);
nor U26823 (N_26823,N_22803,N_23853);
nand U26824 (N_26824,N_23626,N_22401);
or U26825 (N_26825,N_24426,N_21545);
and U26826 (N_26826,N_24849,N_24925);
and U26827 (N_26827,N_23423,N_22877);
nand U26828 (N_26828,N_23618,N_21882);
nand U26829 (N_26829,N_23598,N_21153);
and U26830 (N_26830,N_20931,N_21824);
xnor U26831 (N_26831,N_22305,N_20836);
xor U26832 (N_26832,N_22509,N_24073);
and U26833 (N_26833,N_22919,N_22505);
nand U26834 (N_26834,N_21180,N_20175);
and U26835 (N_26835,N_22995,N_21461);
or U26836 (N_26836,N_21383,N_21028);
or U26837 (N_26837,N_21561,N_20886);
nor U26838 (N_26838,N_24793,N_20269);
or U26839 (N_26839,N_23118,N_21938);
nor U26840 (N_26840,N_23481,N_21896);
nand U26841 (N_26841,N_22896,N_22422);
nor U26842 (N_26842,N_22790,N_23621);
or U26843 (N_26843,N_24827,N_21155);
nor U26844 (N_26844,N_24447,N_22143);
nand U26845 (N_26845,N_20614,N_23956);
nor U26846 (N_26846,N_20772,N_22868);
or U26847 (N_26847,N_21208,N_20363);
or U26848 (N_26848,N_21273,N_20556);
nand U26849 (N_26849,N_21249,N_23945);
xnor U26850 (N_26850,N_20628,N_24898);
and U26851 (N_26851,N_23514,N_24434);
xnor U26852 (N_26852,N_22261,N_20872);
nor U26853 (N_26853,N_24076,N_24549);
nand U26854 (N_26854,N_24351,N_24017);
xor U26855 (N_26855,N_23097,N_22003);
nor U26856 (N_26856,N_23769,N_22083);
nor U26857 (N_26857,N_23478,N_20669);
nand U26858 (N_26858,N_20459,N_22192);
or U26859 (N_26859,N_23570,N_21660);
xnor U26860 (N_26860,N_20004,N_21664);
or U26861 (N_26861,N_24639,N_22825);
nand U26862 (N_26862,N_24282,N_20375);
xor U26863 (N_26863,N_20787,N_23438);
and U26864 (N_26864,N_21571,N_20627);
nand U26865 (N_26865,N_23742,N_21301);
or U26866 (N_26866,N_23239,N_20817);
nand U26867 (N_26867,N_20892,N_22812);
and U26868 (N_26868,N_21195,N_24101);
nor U26869 (N_26869,N_20410,N_23108);
nor U26870 (N_26870,N_21151,N_20991);
nor U26871 (N_26871,N_23965,N_24665);
or U26872 (N_26872,N_23159,N_23653);
nor U26873 (N_26873,N_20322,N_23747);
nor U26874 (N_26874,N_23385,N_24406);
nor U26875 (N_26875,N_21527,N_24763);
and U26876 (N_26876,N_21119,N_24875);
and U26877 (N_26877,N_24855,N_23563);
nor U26878 (N_26878,N_21492,N_24545);
or U26879 (N_26879,N_22001,N_24552);
xnor U26880 (N_26880,N_24271,N_21466);
and U26881 (N_26881,N_20839,N_24988);
nand U26882 (N_26882,N_23427,N_24528);
nand U26883 (N_26883,N_20139,N_22310);
nand U26884 (N_26884,N_22817,N_21387);
nand U26885 (N_26885,N_23550,N_20234);
or U26886 (N_26886,N_23056,N_22107);
nor U26887 (N_26887,N_21562,N_20843);
nand U26888 (N_26888,N_24965,N_22394);
or U26889 (N_26889,N_24409,N_21547);
nor U26890 (N_26890,N_20599,N_24244);
nand U26891 (N_26891,N_20625,N_20863);
or U26892 (N_26892,N_22534,N_23198);
and U26893 (N_26893,N_20009,N_20933);
xor U26894 (N_26894,N_20975,N_23435);
and U26895 (N_26895,N_21143,N_22814);
and U26896 (N_26896,N_20419,N_23999);
nor U26897 (N_26897,N_20122,N_24050);
nand U26898 (N_26898,N_20508,N_22683);
xnor U26899 (N_26899,N_22533,N_22047);
or U26900 (N_26900,N_21204,N_24010);
nor U26901 (N_26901,N_20211,N_22275);
nor U26902 (N_26902,N_24199,N_23805);
nand U26903 (N_26903,N_21982,N_24389);
nor U26904 (N_26904,N_24983,N_21618);
or U26905 (N_26905,N_22137,N_21043);
or U26906 (N_26906,N_24297,N_21808);
nand U26907 (N_26907,N_24460,N_21451);
and U26908 (N_26908,N_23019,N_21814);
and U26909 (N_26909,N_23412,N_21861);
nand U26910 (N_26910,N_20397,N_21916);
nand U26911 (N_26911,N_22887,N_22593);
xnor U26912 (N_26912,N_20655,N_23355);
nand U26913 (N_26913,N_23890,N_20189);
or U26914 (N_26914,N_22753,N_23611);
nor U26915 (N_26915,N_21744,N_21179);
xor U26916 (N_26916,N_20861,N_23864);
or U26917 (N_26917,N_22878,N_20744);
or U26918 (N_26918,N_22316,N_21109);
and U26919 (N_26919,N_20331,N_22947);
nand U26920 (N_26920,N_21235,N_23509);
nor U26921 (N_26921,N_24081,N_22656);
nor U26922 (N_26922,N_20695,N_22607);
nor U26923 (N_26923,N_22845,N_23535);
and U26924 (N_26924,N_21546,N_22053);
or U26925 (N_26925,N_24286,N_22474);
nor U26926 (N_26926,N_20384,N_24366);
nand U26927 (N_26927,N_20795,N_21348);
xor U26928 (N_26928,N_21495,N_24950);
and U26929 (N_26929,N_20694,N_23330);
nor U26930 (N_26930,N_21040,N_22928);
and U26931 (N_26931,N_23468,N_21554);
or U26932 (N_26932,N_20152,N_22240);
and U26933 (N_26933,N_23433,N_20338);
nor U26934 (N_26934,N_22211,N_22406);
or U26935 (N_26935,N_21328,N_23119);
nor U26936 (N_26936,N_20578,N_21864);
and U26937 (N_26937,N_20528,N_21414);
nor U26938 (N_26938,N_21076,N_24203);
nor U26939 (N_26939,N_20046,N_20013);
and U26940 (N_26940,N_22155,N_24812);
nor U26941 (N_26941,N_21750,N_20873);
nand U26942 (N_26942,N_21226,N_23268);
nand U26943 (N_26943,N_20546,N_22694);
or U26944 (N_26944,N_22010,N_21769);
nand U26945 (N_26945,N_23362,N_23467);
and U26946 (N_26946,N_20100,N_22301);
nand U26947 (N_26947,N_21922,N_24491);
xnor U26948 (N_26948,N_22938,N_22207);
nor U26949 (N_26949,N_23002,N_24280);
nand U26950 (N_26950,N_22267,N_20252);
or U26951 (N_26951,N_23417,N_23808);
or U26952 (N_26952,N_22392,N_20654);
nand U26953 (N_26953,N_21947,N_24921);
and U26954 (N_26954,N_24242,N_22931);
nor U26955 (N_26955,N_22614,N_21920);
nor U26956 (N_26956,N_20081,N_23771);
nand U26957 (N_26957,N_23126,N_21487);
and U26958 (N_26958,N_24002,N_24780);
or U26959 (N_26959,N_23711,N_24627);
or U26960 (N_26960,N_23972,N_22559);
and U26961 (N_26961,N_22888,N_21506);
and U26962 (N_26962,N_20545,N_20216);
and U26963 (N_26963,N_20050,N_22168);
and U26964 (N_26964,N_20504,N_22746);
xnor U26965 (N_26965,N_22929,N_24503);
or U26966 (N_26966,N_21708,N_22804);
and U26967 (N_26967,N_21874,N_23790);
xor U26968 (N_26968,N_23669,N_23171);
nand U26969 (N_26969,N_22174,N_24717);
or U26970 (N_26970,N_20595,N_20527);
nand U26971 (N_26971,N_23502,N_23646);
or U26972 (N_26972,N_20617,N_22191);
nor U26973 (N_26973,N_22861,N_20779);
or U26974 (N_26974,N_22478,N_23317);
xnor U26975 (N_26975,N_20785,N_23066);
or U26976 (N_26976,N_20335,N_20132);
nor U26977 (N_26977,N_21447,N_23666);
xnor U26978 (N_26978,N_22755,N_22339);
nand U26979 (N_26979,N_23424,N_23008);
nand U26980 (N_26980,N_24433,N_21163);
and U26981 (N_26981,N_23566,N_24932);
and U26982 (N_26982,N_22345,N_21061);
nor U26983 (N_26983,N_23597,N_21918);
nor U26984 (N_26984,N_20827,N_23992);
or U26985 (N_26985,N_22685,N_22556);
nor U26986 (N_26986,N_22971,N_23358);
and U26987 (N_26987,N_21687,N_23998);
or U26988 (N_26988,N_24908,N_24333);
and U26989 (N_26989,N_21567,N_21576);
and U26990 (N_26990,N_21742,N_24053);
nand U26991 (N_26991,N_24842,N_24934);
or U26992 (N_26992,N_20697,N_20220);
and U26993 (N_26993,N_23832,N_20272);
or U26994 (N_26994,N_20014,N_24277);
nand U26995 (N_26995,N_20379,N_21000);
xor U26996 (N_26996,N_20677,N_21910);
nand U26997 (N_26997,N_21853,N_23987);
nand U26998 (N_26998,N_24309,N_22164);
and U26999 (N_26999,N_24821,N_22231);
and U27000 (N_27000,N_23061,N_23441);
and U27001 (N_27001,N_21610,N_23889);
nor U27002 (N_27002,N_24227,N_23636);
nand U27003 (N_27003,N_21927,N_24788);
nor U27004 (N_27004,N_23218,N_20002);
xor U27005 (N_27005,N_20131,N_22093);
or U27006 (N_27006,N_20771,N_22749);
and U27007 (N_27007,N_20402,N_21334);
xnor U27008 (N_27008,N_23451,N_20362);
or U27009 (N_27009,N_24703,N_21126);
or U27010 (N_27010,N_24538,N_20656);
or U27011 (N_27011,N_21410,N_22622);
and U27012 (N_27012,N_23941,N_20334);
or U27013 (N_27013,N_23416,N_23409);
nor U27014 (N_27014,N_21418,N_23838);
and U27015 (N_27015,N_21980,N_24144);
nand U27016 (N_27016,N_24643,N_21632);
or U27017 (N_27017,N_22710,N_20639);
nand U27018 (N_27018,N_24840,N_24805);
xor U27019 (N_27019,N_23354,N_21540);
or U27020 (N_27020,N_20937,N_24968);
and U27021 (N_27021,N_22408,N_24126);
nand U27022 (N_27022,N_20420,N_20598);
xor U27023 (N_27023,N_23525,N_24772);
and U27024 (N_27024,N_23384,N_22544);
nor U27025 (N_27025,N_21745,N_23662);
nor U27026 (N_27026,N_23345,N_24929);
nand U27027 (N_27027,N_22530,N_21056);
nand U27028 (N_27028,N_23542,N_24743);
nor U27029 (N_27029,N_24148,N_23534);
and U27030 (N_27030,N_22391,N_21097);
nand U27031 (N_27031,N_23930,N_20145);
or U27032 (N_27032,N_21460,N_24630);
nand U27033 (N_27033,N_23748,N_23898);
or U27034 (N_27034,N_24885,N_23727);
and U27035 (N_27035,N_21101,N_22831);
nand U27036 (N_27036,N_20561,N_21842);
or U27037 (N_27037,N_24577,N_21597);
xor U27038 (N_27038,N_24886,N_24494);
nor U27039 (N_27039,N_21911,N_20378);
xnor U27040 (N_27040,N_23599,N_20016);
nand U27041 (N_27041,N_21996,N_21962);
nand U27042 (N_27042,N_21804,N_23086);
and U27043 (N_27043,N_21941,N_23577);
nand U27044 (N_27044,N_24959,N_23443);
and U27045 (N_27045,N_22306,N_23457);
nor U27046 (N_27046,N_22827,N_22417);
nor U27047 (N_27047,N_20880,N_22091);
and U27048 (N_27048,N_20659,N_20233);
nand U27049 (N_27049,N_24213,N_24490);
and U27050 (N_27050,N_22916,N_21267);
or U27051 (N_27051,N_21521,N_22089);
nor U27052 (N_27052,N_24310,N_20343);
nor U27053 (N_27053,N_23845,N_21792);
and U27054 (N_27054,N_23512,N_24900);
nor U27055 (N_27055,N_22195,N_20112);
nor U27056 (N_27056,N_20706,N_24609);
xnor U27057 (N_27057,N_24470,N_20881);
nand U27058 (N_27058,N_23784,N_21515);
nand U27059 (N_27059,N_23852,N_23821);
and U27060 (N_27060,N_20952,N_21648);
or U27061 (N_27061,N_20001,N_21689);
and U27062 (N_27062,N_21412,N_24762);
or U27063 (N_27063,N_21115,N_22805);
nor U27064 (N_27064,N_22485,N_24803);
nand U27065 (N_27065,N_21430,N_23363);
xnor U27066 (N_27066,N_23202,N_20657);
nand U27067 (N_27067,N_22643,N_21426);
xnor U27068 (N_27068,N_21604,N_22761);
nor U27069 (N_27069,N_24589,N_24007);
nand U27070 (N_27070,N_20500,N_20956);
nor U27071 (N_27071,N_20365,N_24625);
nor U27072 (N_27072,N_21280,N_20667);
xnor U27073 (N_27073,N_21805,N_23072);
and U27074 (N_27074,N_24110,N_22449);
or U27075 (N_27075,N_22771,N_20201);
and U27076 (N_27076,N_24004,N_23822);
nand U27077 (N_27077,N_24437,N_23464);
or U27078 (N_27078,N_22941,N_20367);
and U27079 (N_27079,N_21424,N_21004);
and U27080 (N_27080,N_21231,N_23047);
and U27081 (N_27081,N_22586,N_23226);
and U27082 (N_27082,N_23519,N_22765);
and U27083 (N_27083,N_20035,N_24094);
nand U27084 (N_27084,N_21850,N_21813);
xnor U27085 (N_27085,N_20763,N_24523);
nor U27086 (N_27086,N_21309,N_21182);
nand U27087 (N_27087,N_24106,N_21452);
and U27088 (N_27088,N_21074,N_24045);
and U27089 (N_27089,N_24220,N_22689);
or U27090 (N_27090,N_21694,N_22779);
or U27091 (N_27091,N_20989,N_24300);
nor U27092 (N_27092,N_23220,N_23492);
xnor U27093 (N_27093,N_21754,N_22570);
and U27094 (N_27094,N_24450,N_23375);
nor U27095 (N_27095,N_23182,N_24611);
nand U27096 (N_27096,N_23743,N_20386);
nand U27097 (N_27097,N_20257,N_24575);
and U27098 (N_27098,N_23585,N_24251);
nor U27099 (N_27099,N_23753,N_20210);
nor U27100 (N_27100,N_24775,N_22274);
xor U27101 (N_27101,N_21643,N_23408);
nor U27102 (N_27102,N_21690,N_24452);
or U27103 (N_27103,N_20759,N_23434);
and U27104 (N_27104,N_20560,N_21346);
xnor U27105 (N_27105,N_24416,N_22638);
nor U27106 (N_27106,N_22062,N_24662);
nor U27107 (N_27107,N_22470,N_23781);
xor U27108 (N_27108,N_20308,N_22068);
nand U27109 (N_27109,N_20460,N_21250);
nor U27110 (N_27110,N_23617,N_22224);
or U27111 (N_27111,N_22367,N_23012);
nor U27112 (N_27112,N_24970,N_23593);
nand U27113 (N_27113,N_22843,N_22863);
and U27114 (N_27114,N_23177,N_22104);
and U27115 (N_27115,N_21009,N_23516);
xor U27116 (N_27116,N_20151,N_21794);
or U27117 (N_27117,N_20443,N_20102);
or U27118 (N_27118,N_22447,N_20926);
and U27119 (N_27119,N_21011,N_23057);
nor U27120 (N_27120,N_22472,N_23009);
or U27121 (N_27121,N_21100,N_24239);
xnor U27122 (N_27122,N_24650,N_24659);
and U27123 (N_27123,N_20531,N_21771);
nor U27124 (N_27124,N_24521,N_22360);
or U27125 (N_27125,N_21322,N_20987);
and U27126 (N_27126,N_23539,N_24186);
or U27127 (N_27127,N_20330,N_24742);
and U27128 (N_27128,N_22434,N_22953);
and U27129 (N_27129,N_21035,N_22822);
nor U27130 (N_27130,N_22059,N_23264);
or U27131 (N_27131,N_22566,N_24554);
nand U27132 (N_27132,N_20469,N_22674);
nor U27133 (N_27133,N_24219,N_21807);
or U27134 (N_27134,N_23477,N_24701);
nor U27135 (N_27135,N_20467,N_24254);
nand U27136 (N_27136,N_24726,N_20235);
nand U27137 (N_27137,N_24746,N_21345);
and U27138 (N_27138,N_24125,N_24164);
nand U27139 (N_27139,N_20259,N_21164);
nand U27140 (N_27140,N_21914,N_20809);
and U27141 (N_27141,N_23738,N_20076);
xor U27142 (N_27142,N_23693,N_23452);
or U27143 (N_27143,N_20554,N_24131);
nor U27144 (N_27144,N_23500,N_22912);
nand U27145 (N_27145,N_22389,N_20071);
and U27146 (N_27146,N_24646,N_23860);
nor U27147 (N_27147,N_24888,N_20751);
and U27148 (N_27148,N_24544,N_21353);
and U27149 (N_27149,N_20055,N_23248);
or U27150 (N_27150,N_22627,N_24559);
or U27151 (N_27151,N_21392,N_23241);
nand U27152 (N_27152,N_20957,N_21323);
xnor U27153 (N_27153,N_23042,N_23016);
nor U27154 (N_27154,N_21310,N_22050);
nand U27155 (N_27155,N_20762,N_23011);
or U27156 (N_27156,N_21438,N_22436);
or U27157 (N_27157,N_24421,N_22160);
and U27158 (N_27158,N_20073,N_20811);
nand U27159 (N_27159,N_21582,N_24712);
nor U27160 (N_27160,N_22596,N_24318);
nor U27161 (N_27161,N_21673,N_22722);
nand U27162 (N_27162,N_23674,N_22077);
and U27163 (N_27163,N_21336,N_20755);
nand U27164 (N_27164,N_21929,N_23850);
xnor U27165 (N_27165,N_22554,N_21722);
nand U27166 (N_27166,N_22598,N_24877);
or U27167 (N_27167,N_24497,N_20288);
or U27168 (N_27168,N_21514,N_24278);
nand U27169 (N_27169,N_24931,N_21343);
or U27170 (N_27170,N_23350,N_21229);
and U27171 (N_27171,N_24737,N_20424);
nand U27172 (N_27172,N_23348,N_24964);
and U27173 (N_27173,N_20135,N_21589);
and U27174 (N_27174,N_20173,N_24210);
nor U27175 (N_27175,N_21312,N_21654);
xor U27176 (N_27176,N_23462,N_21112);
nand U27177 (N_27177,N_23169,N_22617);
and U27178 (N_27178,N_20307,N_21044);
nor U27179 (N_27179,N_23635,N_23199);
nor U27180 (N_27180,N_22076,N_20783);
or U27181 (N_27181,N_21739,N_22265);
nor U27182 (N_27182,N_23658,N_24702);
nand U27183 (N_27183,N_24603,N_22940);
nor U27184 (N_27184,N_20573,N_24640);
and U27185 (N_27185,N_23184,N_22027);
or U27186 (N_27186,N_22738,N_23219);
nor U27187 (N_27187,N_21219,N_21993);
nand U27188 (N_27188,N_22296,N_23141);
and U27189 (N_27189,N_21497,N_20616);
nor U27190 (N_27190,N_23447,N_24768);
and U27191 (N_27191,N_22072,N_20137);
nor U27192 (N_27192,N_21846,N_24152);
and U27193 (N_27193,N_23020,N_22577);
or U27194 (N_27194,N_23873,N_20103);
xnor U27195 (N_27195,N_23521,N_21531);
and U27196 (N_27196,N_20530,N_20239);
and U27197 (N_27197,N_23445,N_22431);
nand U27198 (N_27198,N_21534,N_22002);
and U27199 (N_27199,N_20306,N_22676);
nor U27200 (N_27200,N_20494,N_22230);
xor U27201 (N_27201,N_20107,N_22295);
nor U27202 (N_27202,N_20940,N_24897);
nand U27203 (N_27203,N_23287,N_23413);
nor U27204 (N_27204,N_24937,N_22318);
xor U27205 (N_27205,N_24807,N_20692);
or U27206 (N_27206,N_20682,N_22635);
nor U27207 (N_27207,N_21105,N_24367);
or U27208 (N_27208,N_23444,N_21397);
nor U27209 (N_27209,N_23142,N_21933);
or U27210 (N_27210,N_20501,N_22605);
nand U27211 (N_27211,N_22257,N_22249);
nand U27212 (N_27212,N_24999,N_23632);
and U27213 (N_27213,N_24893,N_22754);
or U27214 (N_27214,N_22388,N_20301);
and U27215 (N_27215,N_22288,N_20217);
and U27216 (N_27216,N_24798,N_20041);
or U27217 (N_27217,N_23034,N_20021);
nand U27218 (N_27218,N_21403,N_23370);
or U27219 (N_27219,N_23235,N_24124);
nand U27220 (N_27220,N_21200,N_23668);
or U27221 (N_27221,N_20208,N_22418);
and U27222 (N_27222,N_21770,N_22018);
and U27223 (N_27223,N_23067,N_24162);
and U27224 (N_27224,N_20276,N_21594);
nand U27225 (N_27225,N_21157,N_22178);
nand U27226 (N_27226,N_23561,N_22611);
nor U27227 (N_27227,N_23552,N_21517);
nand U27228 (N_27228,N_20169,N_20025);
nand U27229 (N_27229,N_21218,N_24457);
nor U27230 (N_27230,N_24272,N_24795);
nand U27231 (N_27231,N_23536,N_22932);
and U27232 (N_27232,N_24935,N_23709);
xnor U27233 (N_27233,N_22704,N_24527);
nand U27234 (N_27234,N_24307,N_22080);
nand U27235 (N_27235,N_21550,N_23584);
and U27236 (N_27236,N_21091,N_22866);
and U27237 (N_27237,N_20923,N_24476);
or U27238 (N_27238,N_23454,N_24299);
and U27239 (N_27239,N_22079,N_22864);
and U27240 (N_27240,N_24401,N_24385);
and U27241 (N_27241,N_24928,N_20587);
or U27242 (N_27242,N_20806,N_23912);
xor U27243 (N_27243,N_22259,N_20138);
and U27244 (N_27244,N_21453,N_21662);
and U27245 (N_27245,N_22209,N_20688);
or U27246 (N_27246,N_23327,N_22631);
nor U27247 (N_27247,N_23601,N_22844);
or U27248 (N_27248,N_21669,N_23735);
xnor U27249 (N_27249,N_22455,N_22136);
xnor U27250 (N_27250,N_24008,N_21776);
or U27251 (N_27251,N_21378,N_22550);
xor U27252 (N_27252,N_23261,N_21107);
nand U27253 (N_27253,N_21436,N_22832);
nor U27254 (N_27254,N_21894,N_24380);
nor U27255 (N_27255,N_20651,N_23152);
nor U27256 (N_27256,N_21701,N_20147);
nand U27257 (N_27257,N_20146,N_24604);
nor U27258 (N_27258,N_20615,N_23099);
nor U27259 (N_27259,N_21450,N_21979);
nand U27260 (N_27260,N_21440,N_22667);
nand U27261 (N_27261,N_24779,N_20609);
and U27262 (N_27262,N_20965,N_23205);
nand U27263 (N_27263,N_20032,N_24683);
nand U27264 (N_27264,N_21117,N_24279);
xor U27265 (N_27265,N_22502,N_21376);
xnor U27266 (N_27266,N_21995,N_23877);
or U27267 (N_27267,N_21252,N_23623);
nor U27268 (N_27268,N_23140,N_20116);
or U27269 (N_27269,N_21209,N_22893);
nor U27270 (N_27270,N_23924,N_21413);
and U27271 (N_27271,N_20979,N_22576);
and U27272 (N_27272,N_22412,N_24860);
or U27273 (N_27273,N_21050,N_24085);
nand U27274 (N_27274,N_23372,N_21728);
and U27275 (N_27275,N_22307,N_20850);
and U27276 (N_27276,N_21070,N_23495);
and U27277 (N_27277,N_23270,N_23267);
or U27278 (N_27278,N_24192,N_22013);
and U27279 (N_27279,N_24363,N_20802);
and U27280 (N_27280,N_20172,N_21925);
xor U27281 (N_27281,N_20637,N_21333);
and U27282 (N_27282,N_21932,N_21764);
nand U27283 (N_27283,N_23278,N_22328);
xor U27284 (N_27284,N_22719,N_21342);
or U27285 (N_27285,N_21780,N_20678);
nand U27286 (N_27286,N_24013,N_24524);
and U27287 (N_27287,N_23746,N_23730);
or U27288 (N_27288,N_20499,N_20540);
nand U27289 (N_27289,N_20883,N_21423);
nor U27290 (N_27290,N_21573,N_21733);
nand U27291 (N_27291,N_22958,N_24724);
nand U27292 (N_27292,N_20822,N_24794);
xor U27293 (N_27293,N_20000,N_20044);
or U27294 (N_27294,N_23164,N_23074);
and U27295 (N_27295,N_24270,N_22121);
and U27296 (N_27296,N_22102,N_20860);
and U27297 (N_27297,N_21354,N_20030);
nor U27298 (N_27298,N_21411,N_20502);
or U27299 (N_27299,N_22688,N_22962);
or U27300 (N_27300,N_21877,N_22990);
and U27301 (N_27301,N_20972,N_24924);
or U27302 (N_27302,N_21945,N_24581);
nor U27303 (N_27303,N_22145,N_21248);
nand U27304 (N_27304,N_23564,N_22215);
nor U27305 (N_27305,N_21031,N_23407);
nor U27306 (N_27306,N_20399,N_20792);
nand U27307 (N_27307,N_24448,N_21139);
nand U27308 (N_27308,N_23929,N_21269);
nand U27309 (N_27309,N_21090,N_24799);
or U27310 (N_27310,N_20406,N_22943);
nand U27311 (N_27311,N_20821,N_21559);
or U27312 (N_27312,N_23211,N_22708);
nand U27313 (N_27313,N_20417,N_20101);
xor U27314 (N_27314,N_24810,N_23606);
nor U27315 (N_27315,N_24079,N_23401);
nand U27316 (N_27316,N_24980,N_23800);
and U27317 (N_27317,N_21617,N_22669);
and U27318 (N_27318,N_21581,N_23027);
nor U27319 (N_27319,N_20401,N_23726);
and U27320 (N_27320,N_21782,N_22862);
nor U27321 (N_27321,N_24945,N_20260);
or U27322 (N_27322,N_21723,N_20056);
and U27323 (N_27323,N_23783,N_20908);
nand U27324 (N_27324,N_23170,N_21970);
xnor U27325 (N_27325,N_24957,N_22727);
xnor U27326 (N_27326,N_21053,N_24784);
and U27327 (N_27327,N_22668,N_21509);
or U27328 (N_27328,N_23392,N_24792);
or U27329 (N_27329,N_23624,N_21798);
and U27330 (N_27330,N_21638,N_22562);
or U27331 (N_27331,N_21067,N_23831);
and U27332 (N_27332,N_24740,N_23660);
and U27333 (N_27333,N_24576,N_20005);
and U27334 (N_27334,N_21553,N_20356);
and U27335 (N_27335,N_21767,N_22236);
xor U27336 (N_27336,N_22198,N_21934);
or U27337 (N_27337,N_24035,N_23689);
or U27338 (N_27338,N_23788,N_21502);
nand U27339 (N_27339,N_22460,N_21016);
and U27340 (N_27340,N_24654,N_24956);
nor U27341 (N_27341,N_20719,N_21259);
or U27342 (N_27342,N_22528,N_24159);
and U27343 (N_27343,N_20431,N_21503);
nor U27344 (N_27344,N_24145,N_23426);
or U27345 (N_27345,N_20830,N_22341);
nand U27346 (N_27346,N_22508,N_22884);
or U27347 (N_27347,N_24290,N_20672);
nor U27348 (N_27348,N_24834,N_21751);
nor U27349 (N_27349,N_21670,N_24025);
nand U27350 (N_27350,N_20274,N_20928);
nor U27351 (N_27351,N_21136,N_21787);
xnor U27352 (N_27352,N_24570,N_21658);
nand U27353 (N_27353,N_23386,N_21351);
nor U27354 (N_27354,N_21726,N_24939);
nand U27355 (N_27355,N_24596,N_20959);
nand U27356 (N_27356,N_21482,N_24072);
or U27357 (N_27357,N_22959,N_22847);
nand U27358 (N_27358,N_21484,N_22899);
xor U27359 (N_27359,N_23752,N_24256);
nand U27360 (N_27360,N_23989,N_24399);
nand U27361 (N_27361,N_20986,N_20352);
or U27362 (N_27362,N_23133,N_21295);
nand U27363 (N_27363,N_21586,N_24009);
nand U27364 (N_27364,N_21092,N_22063);
nand U27365 (N_27365,N_20708,N_23128);
nor U27366 (N_27366,N_24111,N_20097);
or U27367 (N_27367,N_22782,N_21088);
or U27368 (N_27368,N_24504,N_23859);
xnor U27369 (N_27369,N_21522,N_21062);
or U27370 (N_27370,N_20590,N_21607);
or U27371 (N_27371,N_22745,N_23603);
or U27372 (N_27372,N_24396,N_23271);
nor U27373 (N_27373,N_21474,N_23760);
xnor U27374 (N_27374,N_21647,N_20938);
nor U27375 (N_27375,N_20497,N_24681);
nor U27376 (N_27376,N_20366,N_23111);
nor U27377 (N_27377,N_22411,N_21731);
xnor U27378 (N_27378,N_20893,N_21033);
nand U27379 (N_27379,N_22956,N_24456);
or U27380 (N_27380,N_21081,N_21968);
and U27381 (N_27381,N_20577,N_23543);
or U27382 (N_27382,N_20603,N_24143);
or U27383 (N_27383,N_21166,N_24088);
nand U27384 (N_27384,N_20377,N_22359);
and U27385 (N_27385,N_20136,N_23314);
nand U27386 (N_27386,N_20634,N_23320);
xnor U27387 (N_27387,N_23789,N_22250);
and U27388 (N_27388,N_20042,N_20510);
nand U27389 (N_27389,N_20521,N_20652);
nor U27390 (N_27390,N_21791,N_20179);
nor U27391 (N_27391,N_23280,N_22728);
or U27392 (N_27392,N_24431,N_21866);
and U27393 (N_27393,N_23558,N_24012);
nor U27394 (N_27394,N_21732,N_22282);
or U27395 (N_27395,N_23436,N_22303);
nor U27396 (N_27396,N_20344,N_23655);
nor U27397 (N_27397,N_20662,N_22253);
and U27398 (N_27398,N_22730,N_22713);
nor U27399 (N_27399,N_23389,N_20125);
or U27400 (N_27400,N_20084,N_22682);
and U27401 (N_27401,N_21584,N_22549);
and U27402 (N_27402,N_20717,N_24704);
and U27403 (N_27403,N_21809,N_24071);
xor U27404 (N_27404,N_23166,N_24878);
nand U27405 (N_27405,N_24302,N_23010);
nor U27406 (N_27406,N_20124,N_20225);
nand U27407 (N_27407,N_22591,N_23734);
nor U27408 (N_27408,N_24161,N_20552);
and U27409 (N_27409,N_23149,N_20757);
and U27410 (N_27410,N_24512,N_21587);
nand U27411 (N_27411,N_23146,N_20905);
or U27412 (N_27412,N_23766,N_23046);
nor U27413 (N_27413,N_24499,N_24748);
nand U27414 (N_27414,N_24735,N_21367);
nand U27415 (N_27415,N_22205,N_22486);
xnor U27416 (N_27416,N_23596,N_22309);
nor U27417 (N_27417,N_22620,N_22499);
or U27418 (N_27418,N_20555,N_22636);
nand U27419 (N_27419,N_22403,N_22426);
and U27420 (N_27420,N_22902,N_22721);
nand U27421 (N_27421,N_24969,N_23347);
nor U27422 (N_27422,N_20710,N_24268);
nand U27423 (N_27423,N_21622,N_20149);
or U27424 (N_27424,N_21036,N_23741);
or U27425 (N_27425,N_21811,N_23710);
nor U27426 (N_27426,N_20911,N_21730);
or U27427 (N_27427,N_20711,N_20426);
and U27428 (N_27428,N_21069,N_23518);
nand U27429 (N_27429,N_20465,N_22358);
nand U27430 (N_27430,N_22675,N_22970);
nand U27431 (N_27431,N_24353,N_23737);
nand U27432 (N_27432,N_20198,N_22239);
nand U27433 (N_27433,N_23162,N_24915);
and U27434 (N_27434,N_22503,N_21357);
nand U27435 (N_27435,N_24501,N_22707);
nor U27436 (N_27436,N_20270,N_24446);
nand U27437 (N_27437,N_24582,N_20491);
nor U27438 (N_27438,N_21433,N_24879);
or U27439 (N_27439,N_20815,N_20068);
nand U27440 (N_27440,N_24573,N_20916);
or U27441 (N_27441,N_21721,N_20452);
nand U27442 (N_27442,N_24907,N_22234);
and U27443 (N_27443,N_20339,N_24314);
nand U27444 (N_27444,N_22769,N_20638);
or U27445 (N_27445,N_22036,N_21373);
and U27446 (N_27446,N_23285,N_20245);
nor U27447 (N_27447,N_22833,N_20353);
and U27448 (N_27448,N_21683,N_20371);
and U27449 (N_27449,N_20685,N_20369);
xor U27450 (N_27450,N_24901,N_20020);
nor U27451 (N_27451,N_20341,N_21130);
and U27452 (N_27452,N_22438,N_21612);
nand U27453 (N_27453,N_22292,N_24974);
or U27454 (N_27454,N_23919,N_24415);
nand U27455 (N_27455,N_23568,N_23855);
nand U27456 (N_27456,N_24933,N_20294);
or U27457 (N_27457,N_21875,N_22346);
nand U27458 (N_27458,N_22553,N_21205);
nand U27459 (N_27459,N_23835,N_22260);
nor U27460 (N_27460,N_22385,N_24509);
nor U27461 (N_27461,N_24323,N_22483);
xnor U27462 (N_27462,N_20218,N_24847);
nor U27463 (N_27463,N_23068,N_21193);
nor U27464 (N_27464,N_20222,N_20756);
nand U27465 (N_27465,N_22294,N_20675);
nor U27466 (N_27466,N_24767,N_20243);
xor U27467 (N_27467,N_21021,N_23332);
nor U27468 (N_27468,N_20740,N_24566);
nand U27469 (N_27469,N_23124,N_20058);
xor U27470 (N_27470,N_20487,N_24451);
or U27471 (N_27471,N_20780,N_23928);
nor U27472 (N_27472,N_22955,N_24480);
nor U27473 (N_27473,N_23557,N_20461);
xor U27474 (N_27474,N_21851,N_24721);
nor U27475 (N_27475,N_23513,N_21386);
or U27476 (N_27476,N_22100,N_24588);
nor U27477 (N_27477,N_23028,N_21847);
xnor U27478 (N_27478,N_22419,N_21362);
nor U27479 (N_27479,N_22162,N_23190);
and U27480 (N_27480,N_20392,N_23840);
nand U27481 (N_27481,N_22266,N_24046);
and U27482 (N_27482,N_23483,N_22148);
nand U27483 (N_27483,N_23851,N_22671);
or U27484 (N_27484,N_24525,N_20090);
or U27485 (N_27485,N_21501,N_21737);
or U27486 (N_27486,N_21111,N_24255);
or U27487 (N_27487,N_21592,N_23522);
nand U27488 (N_27488,N_24638,N_22498);
nor U27489 (N_27489,N_21806,N_23300);
nand U27490 (N_27490,N_24896,N_24981);
nand U27491 (N_27491,N_21761,N_22244);
nor U27492 (N_27492,N_24027,N_23333);
nand U27493 (N_27493,N_20293,N_24259);
or U27494 (N_27494,N_20305,N_23977);
nand U27495 (N_27495,N_23393,N_24623);
and U27496 (N_27496,N_22353,N_20310);
nand U27497 (N_27497,N_23394,N_23233);
and U27498 (N_27498,N_20945,N_21437);
and U27499 (N_27499,N_23724,N_24052);
and U27500 (N_27500,N_22855,N_20359);
and U27501 (N_27501,N_21856,N_21985);
and U27502 (N_27502,N_24928,N_20613);
or U27503 (N_27503,N_23857,N_21128);
or U27504 (N_27504,N_24549,N_24652);
or U27505 (N_27505,N_22009,N_20556);
nor U27506 (N_27506,N_23807,N_20605);
and U27507 (N_27507,N_20305,N_23611);
nand U27508 (N_27508,N_23314,N_23190);
nor U27509 (N_27509,N_21995,N_23324);
nor U27510 (N_27510,N_23070,N_22175);
nor U27511 (N_27511,N_20444,N_24370);
xnor U27512 (N_27512,N_20108,N_22119);
nand U27513 (N_27513,N_22784,N_24388);
nor U27514 (N_27514,N_21935,N_24706);
nand U27515 (N_27515,N_24780,N_21369);
nor U27516 (N_27516,N_20984,N_23935);
or U27517 (N_27517,N_23492,N_24182);
and U27518 (N_27518,N_22123,N_23471);
nor U27519 (N_27519,N_22692,N_23559);
nand U27520 (N_27520,N_23494,N_21858);
and U27521 (N_27521,N_23632,N_20136);
or U27522 (N_27522,N_23515,N_20304);
nand U27523 (N_27523,N_21149,N_20171);
xnor U27524 (N_27524,N_20277,N_21712);
nand U27525 (N_27525,N_21766,N_23437);
nand U27526 (N_27526,N_24290,N_22146);
or U27527 (N_27527,N_23689,N_22947);
and U27528 (N_27528,N_21812,N_24040);
or U27529 (N_27529,N_21265,N_20606);
and U27530 (N_27530,N_22022,N_20801);
nor U27531 (N_27531,N_20222,N_21059);
nor U27532 (N_27532,N_21606,N_21526);
nand U27533 (N_27533,N_20880,N_22916);
and U27534 (N_27534,N_23480,N_23271);
nor U27535 (N_27535,N_23014,N_22104);
or U27536 (N_27536,N_20994,N_23304);
or U27537 (N_27537,N_22449,N_24625);
nand U27538 (N_27538,N_20004,N_20629);
xnor U27539 (N_27539,N_23618,N_20094);
and U27540 (N_27540,N_24492,N_21943);
nor U27541 (N_27541,N_20029,N_22700);
or U27542 (N_27542,N_23960,N_24184);
and U27543 (N_27543,N_20954,N_21167);
nor U27544 (N_27544,N_23142,N_24329);
or U27545 (N_27545,N_24843,N_21982);
or U27546 (N_27546,N_22759,N_24009);
and U27547 (N_27547,N_24354,N_20668);
xor U27548 (N_27548,N_21383,N_20010);
nor U27549 (N_27549,N_24045,N_23491);
nor U27550 (N_27550,N_20758,N_21765);
or U27551 (N_27551,N_22923,N_21927);
or U27552 (N_27552,N_20553,N_22519);
nand U27553 (N_27553,N_23537,N_23408);
or U27554 (N_27554,N_22013,N_20112);
or U27555 (N_27555,N_23292,N_24200);
or U27556 (N_27556,N_22781,N_21487);
and U27557 (N_27557,N_22552,N_23209);
or U27558 (N_27558,N_23634,N_22956);
and U27559 (N_27559,N_21517,N_20697);
or U27560 (N_27560,N_21037,N_20215);
or U27561 (N_27561,N_21549,N_22134);
xor U27562 (N_27562,N_22877,N_24640);
or U27563 (N_27563,N_20621,N_22846);
xor U27564 (N_27564,N_21380,N_21760);
nor U27565 (N_27565,N_24729,N_20375);
and U27566 (N_27566,N_24089,N_24232);
nand U27567 (N_27567,N_22112,N_23221);
and U27568 (N_27568,N_23640,N_24270);
nor U27569 (N_27569,N_20700,N_22939);
or U27570 (N_27570,N_24586,N_24025);
or U27571 (N_27571,N_21103,N_24434);
nand U27572 (N_27572,N_22691,N_24477);
and U27573 (N_27573,N_20853,N_20641);
xor U27574 (N_27574,N_20237,N_24099);
nor U27575 (N_27575,N_22292,N_21709);
or U27576 (N_27576,N_21401,N_21995);
or U27577 (N_27577,N_21146,N_20178);
or U27578 (N_27578,N_21086,N_23111);
and U27579 (N_27579,N_23807,N_24167);
and U27580 (N_27580,N_20938,N_23040);
nor U27581 (N_27581,N_22412,N_21684);
nand U27582 (N_27582,N_23810,N_24827);
nor U27583 (N_27583,N_21046,N_23384);
and U27584 (N_27584,N_22968,N_24230);
nor U27585 (N_27585,N_24991,N_24462);
and U27586 (N_27586,N_24465,N_22784);
or U27587 (N_27587,N_22114,N_22356);
nor U27588 (N_27588,N_20759,N_22890);
nor U27589 (N_27589,N_23666,N_20698);
and U27590 (N_27590,N_23062,N_21139);
nand U27591 (N_27591,N_22198,N_22220);
and U27592 (N_27592,N_23324,N_21444);
nor U27593 (N_27593,N_23518,N_21215);
or U27594 (N_27594,N_20014,N_23766);
nand U27595 (N_27595,N_24633,N_23186);
xor U27596 (N_27596,N_20125,N_24247);
nor U27597 (N_27597,N_24294,N_23192);
nor U27598 (N_27598,N_20882,N_22629);
xor U27599 (N_27599,N_24929,N_24937);
and U27600 (N_27600,N_20447,N_24114);
nor U27601 (N_27601,N_22817,N_22408);
or U27602 (N_27602,N_20678,N_24862);
and U27603 (N_27603,N_20276,N_22693);
or U27604 (N_27604,N_20202,N_24143);
and U27605 (N_27605,N_23178,N_23712);
and U27606 (N_27606,N_20348,N_23535);
nor U27607 (N_27607,N_21269,N_23135);
and U27608 (N_27608,N_24060,N_20610);
or U27609 (N_27609,N_22738,N_22884);
nor U27610 (N_27610,N_21509,N_22810);
nor U27611 (N_27611,N_21552,N_20837);
nor U27612 (N_27612,N_21485,N_24914);
xor U27613 (N_27613,N_24870,N_24105);
or U27614 (N_27614,N_24790,N_21721);
or U27615 (N_27615,N_22144,N_20802);
nand U27616 (N_27616,N_22025,N_21336);
xor U27617 (N_27617,N_24500,N_21538);
and U27618 (N_27618,N_22274,N_22690);
and U27619 (N_27619,N_22686,N_22061);
xnor U27620 (N_27620,N_23671,N_23404);
or U27621 (N_27621,N_23589,N_24875);
and U27622 (N_27622,N_21834,N_23471);
nor U27623 (N_27623,N_21859,N_24992);
and U27624 (N_27624,N_24270,N_22372);
nand U27625 (N_27625,N_21406,N_23754);
xor U27626 (N_27626,N_24526,N_24395);
nand U27627 (N_27627,N_24204,N_21852);
or U27628 (N_27628,N_20216,N_20772);
nand U27629 (N_27629,N_20484,N_21640);
nor U27630 (N_27630,N_24609,N_21487);
and U27631 (N_27631,N_21251,N_21412);
xor U27632 (N_27632,N_23166,N_21700);
nand U27633 (N_27633,N_20995,N_24202);
nand U27634 (N_27634,N_23263,N_21643);
nand U27635 (N_27635,N_23110,N_23542);
or U27636 (N_27636,N_24816,N_21130);
nor U27637 (N_27637,N_24594,N_20010);
and U27638 (N_27638,N_22760,N_21439);
and U27639 (N_27639,N_20911,N_20914);
or U27640 (N_27640,N_23804,N_21480);
nor U27641 (N_27641,N_24115,N_21886);
nor U27642 (N_27642,N_21771,N_22480);
and U27643 (N_27643,N_23774,N_23159);
and U27644 (N_27644,N_22999,N_20148);
nand U27645 (N_27645,N_20689,N_23296);
nand U27646 (N_27646,N_21153,N_24272);
nor U27647 (N_27647,N_21498,N_21672);
nand U27648 (N_27648,N_24581,N_20228);
and U27649 (N_27649,N_20518,N_23987);
nor U27650 (N_27650,N_21233,N_23864);
and U27651 (N_27651,N_24356,N_23500);
nor U27652 (N_27652,N_20248,N_21830);
or U27653 (N_27653,N_24825,N_20055);
or U27654 (N_27654,N_20072,N_23003);
nand U27655 (N_27655,N_24669,N_23896);
nor U27656 (N_27656,N_20202,N_22393);
nor U27657 (N_27657,N_20263,N_22145);
nand U27658 (N_27658,N_24060,N_22259);
and U27659 (N_27659,N_22669,N_24415);
nand U27660 (N_27660,N_24630,N_23216);
nand U27661 (N_27661,N_20139,N_21734);
nand U27662 (N_27662,N_24208,N_23020);
nor U27663 (N_27663,N_22617,N_24291);
and U27664 (N_27664,N_22334,N_22466);
xnor U27665 (N_27665,N_21340,N_20705);
or U27666 (N_27666,N_22447,N_21990);
xnor U27667 (N_27667,N_22285,N_20693);
and U27668 (N_27668,N_22514,N_23891);
or U27669 (N_27669,N_21670,N_20762);
nor U27670 (N_27670,N_24627,N_24215);
nand U27671 (N_27671,N_20847,N_23680);
and U27672 (N_27672,N_21060,N_23414);
nor U27673 (N_27673,N_22871,N_21229);
or U27674 (N_27674,N_21882,N_22048);
or U27675 (N_27675,N_21622,N_22429);
nor U27676 (N_27676,N_22358,N_24787);
nand U27677 (N_27677,N_20671,N_23861);
or U27678 (N_27678,N_20384,N_23734);
or U27679 (N_27679,N_23115,N_22452);
and U27680 (N_27680,N_23144,N_24678);
and U27681 (N_27681,N_22991,N_22929);
nor U27682 (N_27682,N_23667,N_21415);
and U27683 (N_27683,N_24642,N_22018);
or U27684 (N_27684,N_21450,N_24985);
xnor U27685 (N_27685,N_21430,N_21926);
nor U27686 (N_27686,N_22038,N_21706);
or U27687 (N_27687,N_22039,N_23850);
or U27688 (N_27688,N_23690,N_20099);
or U27689 (N_27689,N_22729,N_22073);
xor U27690 (N_27690,N_20807,N_20743);
xor U27691 (N_27691,N_22994,N_22329);
or U27692 (N_27692,N_22559,N_21492);
nor U27693 (N_27693,N_24176,N_24687);
nor U27694 (N_27694,N_24860,N_20136);
nor U27695 (N_27695,N_22877,N_20400);
or U27696 (N_27696,N_23722,N_20670);
nand U27697 (N_27697,N_20853,N_23521);
nand U27698 (N_27698,N_22261,N_24684);
or U27699 (N_27699,N_21463,N_22156);
and U27700 (N_27700,N_23525,N_23152);
or U27701 (N_27701,N_22386,N_20154);
and U27702 (N_27702,N_23151,N_24353);
or U27703 (N_27703,N_24009,N_23323);
and U27704 (N_27704,N_23139,N_24549);
and U27705 (N_27705,N_23193,N_20423);
nor U27706 (N_27706,N_21145,N_21980);
nor U27707 (N_27707,N_21737,N_24835);
and U27708 (N_27708,N_20750,N_21876);
nand U27709 (N_27709,N_22116,N_23928);
nor U27710 (N_27710,N_22317,N_20803);
nand U27711 (N_27711,N_20682,N_24604);
or U27712 (N_27712,N_22997,N_24819);
and U27713 (N_27713,N_21300,N_21149);
and U27714 (N_27714,N_24868,N_24679);
xor U27715 (N_27715,N_24089,N_23490);
nor U27716 (N_27716,N_23097,N_23499);
and U27717 (N_27717,N_24690,N_20483);
xor U27718 (N_27718,N_21108,N_22465);
nand U27719 (N_27719,N_23137,N_22152);
or U27720 (N_27720,N_22096,N_22580);
or U27721 (N_27721,N_23999,N_23318);
or U27722 (N_27722,N_20152,N_23941);
nand U27723 (N_27723,N_20503,N_23400);
nor U27724 (N_27724,N_24652,N_22522);
nand U27725 (N_27725,N_24007,N_22244);
and U27726 (N_27726,N_20250,N_22246);
and U27727 (N_27727,N_21715,N_22683);
nor U27728 (N_27728,N_21409,N_24069);
nand U27729 (N_27729,N_21863,N_20001);
or U27730 (N_27730,N_22230,N_20764);
nand U27731 (N_27731,N_24723,N_21582);
or U27732 (N_27732,N_23543,N_23542);
or U27733 (N_27733,N_20449,N_23675);
xor U27734 (N_27734,N_23117,N_22559);
and U27735 (N_27735,N_23996,N_24497);
and U27736 (N_27736,N_23108,N_24403);
and U27737 (N_27737,N_20754,N_24738);
and U27738 (N_27738,N_24862,N_23668);
xnor U27739 (N_27739,N_22545,N_21212);
or U27740 (N_27740,N_22082,N_22180);
nor U27741 (N_27741,N_22125,N_24984);
xor U27742 (N_27742,N_21040,N_22886);
xnor U27743 (N_27743,N_23297,N_20118);
or U27744 (N_27744,N_22063,N_21724);
nand U27745 (N_27745,N_20660,N_24896);
nor U27746 (N_27746,N_24424,N_24733);
xnor U27747 (N_27747,N_20564,N_23562);
nand U27748 (N_27748,N_21087,N_20522);
nor U27749 (N_27749,N_21281,N_22603);
nand U27750 (N_27750,N_23834,N_24300);
nand U27751 (N_27751,N_22017,N_22589);
or U27752 (N_27752,N_20924,N_23762);
and U27753 (N_27753,N_20765,N_24181);
nor U27754 (N_27754,N_22233,N_23855);
nor U27755 (N_27755,N_20791,N_22435);
or U27756 (N_27756,N_23539,N_21187);
and U27757 (N_27757,N_24068,N_20972);
and U27758 (N_27758,N_24053,N_24792);
xor U27759 (N_27759,N_21571,N_23091);
nor U27760 (N_27760,N_20910,N_23860);
nor U27761 (N_27761,N_23967,N_21759);
and U27762 (N_27762,N_22645,N_23181);
or U27763 (N_27763,N_20270,N_21997);
and U27764 (N_27764,N_24600,N_21886);
xnor U27765 (N_27765,N_23961,N_22723);
and U27766 (N_27766,N_21181,N_23313);
and U27767 (N_27767,N_22937,N_21238);
or U27768 (N_27768,N_21988,N_21918);
nor U27769 (N_27769,N_20845,N_24444);
nor U27770 (N_27770,N_24481,N_23080);
nor U27771 (N_27771,N_21427,N_20708);
xor U27772 (N_27772,N_23113,N_24089);
nand U27773 (N_27773,N_24603,N_23737);
or U27774 (N_27774,N_20580,N_20413);
and U27775 (N_27775,N_24625,N_20217);
nor U27776 (N_27776,N_20964,N_21639);
or U27777 (N_27777,N_23497,N_21416);
and U27778 (N_27778,N_22472,N_22490);
nand U27779 (N_27779,N_24365,N_21684);
nand U27780 (N_27780,N_24405,N_23570);
xnor U27781 (N_27781,N_24996,N_22555);
nor U27782 (N_27782,N_20706,N_23308);
and U27783 (N_27783,N_23727,N_23184);
or U27784 (N_27784,N_21540,N_21294);
or U27785 (N_27785,N_23590,N_22068);
and U27786 (N_27786,N_20681,N_23264);
and U27787 (N_27787,N_20553,N_24412);
nor U27788 (N_27788,N_24949,N_24948);
nand U27789 (N_27789,N_21878,N_21673);
nor U27790 (N_27790,N_24345,N_20540);
or U27791 (N_27791,N_21188,N_20576);
nand U27792 (N_27792,N_20631,N_24091);
nor U27793 (N_27793,N_24251,N_23745);
nand U27794 (N_27794,N_23320,N_20508);
nand U27795 (N_27795,N_24227,N_24402);
or U27796 (N_27796,N_23358,N_20709);
and U27797 (N_27797,N_23524,N_22434);
xor U27798 (N_27798,N_24237,N_23245);
or U27799 (N_27799,N_20850,N_20544);
xor U27800 (N_27800,N_20595,N_24955);
xor U27801 (N_27801,N_22640,N_24347);
nor U27802 (N_27802,N_23194,N_23605);
nand U27803 (N_27803,N_23267,N_21058);
nand U27804 (N_27804,N_21945,N_24287);
nand U27805 (N_27805,N_22528,N_23696);
nand U27806 (N_27806,N_22567,N_20238);
nor U27807 (N_27807,N_22443,N_23349);
or U27808 (N_27808,N_20358,N_23481);
or U27809 (N_27809,N_22672,N_24263);
and U27810 (N_27810,N_24599,N_20237);
and U27811 (N_27811,N_20665,N_22610);
nor U27812 (N_27812,N_24562,N_22534);
or U27813 (N_27813,N_23436,N_23394);
and U27814 (N_27814,N_24777,N_22076);
and U27815 (N_27815,N_24403,N_21072);
nor U27816 (N_27816,N_20706,N_24695);
or U27817 (N_27817,N_22647,N_22127);
and U27818 (N_27818,N_22846,N_24647);
or U27819 (N_27819,N_23488,N_23009);
or U27820 (N_27820,N_23945,N_20914);
nor U27821 (N_27821,N_22632,N_20226);
and U27822 (N_27822,N_20065,N_23966);
nand U27823 (N_27823,N_22844,N_21035);
or U27824 (N_27824,N_24715,N_20809);
nor U27825 (N_27825,N_22876,N_21070);
xnor U27826 (N_27826,N_21319,N_24597);
nor U27827 (N_27827,N_23895,N_23925);
nand U27828 (N_27828,N_24170,N_21448);
and U27829 (N_27829,N_21437,N_22943);
nand U27830 (N_27830,N_24729,N_21860);
or U27831 (N_27831,N_20058,N_20757);
or U27832 (N_27832,N_20967,N_24443);
or U27833 (N_27833,N_20954,N_22764);
or U27834 (N_27834,N_23789,N_23124);
and U27835 (N_27835,N_23738,N_24602);
or U27836 (N_27836,N_20964,N_24599);
and U27837 (N_27837,N_21487,N_22241);
nor U27838 (N_27838,N_23023,N_20646);
nor U27839 (N_27839,N_21035,N_21515);
or U27840 (N_27840,N_22362,N_20263);
or U27841 (N_27841,N_22212,N_24390);
nor U27842 (N_27842,N_22728,N_20761);
or U27843 (N_27843,N_23556,N_23088);
xor U27844 (N_27844,N_23128,N_22292);
nand U27845 (N_27845,N_21621,N_22704);
and U27846 (N_27846,N_22299,N_22618);
or U27847 (N_27847,N_22139,N_21397);
xor U27848 (N_27848,N_24234,N_24684);
and U27849 (N_27849,N_21770,N_23173);
and U27850 (N_27850,N_20160,N_24278);
nand U27851 (N_27851,N_24804,N_21576);
and U27852 (N_27852,N_24356,N_23569);
nand U27853 (N_27853,N_24875,N_24717);
or U27854 (N_27854,N_24944,N_21629);
and U27855 (N_27855,N_23403,N_24582);
xor U27856 (N_27856,N_21188,N_24348);
or U27857 (N_27857,N_22336,N_21041);
nand U27858 (N_27858,N_21446,N_21785);
nor U27859 (N_27859,N_23113,N_20233);
xnor U27860 (N_27860,N_20249,N_20860);
xor U27861 (N_27861,N_23684,N_20577);
or U27862 (N_27862,N_21617,N_23971);
and U27863 (N_27863,N_24991,N_20633);
nand U27864 (N_27864,N_21061,N_22160);
or U27865 (N_27865,N_24753,N_20296);
xnor U27866 (N_27866,N_20573,N_22318);
nand U27867 (N_27867,N_24130,N_20402);
and U27868 (N_27868,N_22627,N_20892);
nand U27869 (N_27869,N_20096,N_22128);
or U27870 (N_27870,N_23900,N_20843);
nand U27871 (N_27871,N_20350,N_23024);
xor U27872 (N_27872,N_22885,N_21473);
or U27873 (N_27873,N_23162,N_20291);
xor U27874 (N_27874,N_21558,N_23192);
and U27875 (N_27875,N_23341,N_22561);
nand U27876 (N_27876,N_20195,N_23461);
and U27877 (N_27877,N_23988,N_22322);
xnor U27878 (N_27878,N_22039,N_24278);
and U27879 (N_27879,N_23113,N_21466);
nand U27880 (N_27880,N_24083,N_24324);
nor U27881 (N_27881,N_22958,N_22843);
nor U27882 (N_27882,N_21172,N_23257);
nor U27883 (N_27883,N_22847,N_24694);
nor U27884 (N_27884,N_23992,N_20804);
and U27885 (N_27885,N_20050,N_24122);
nand U27886 (N_27886,N_20672,N_20156);
or U27887 (N_27887,N_21740,N_22552);
xor U27888 (N_27888,N_21861,N_22847);
and U27889 (N_27889,N_23394,N_21020);
or U27890 (N_27890,N_23135,N_24632);
nand U27891 (N_27891,N_21711,N_20828);
and U27892 (N_27892,N_23967,N_21410);
or U27893 (N_27893,N_24480,N_21792);
nand U27894 (N_27894,N_22575,N_22767);
or U27895 (N_27895,N_22677,N_20172);
nor U27896 (N_27896,N_21138,N_23483);
and U27897 (N_27897,N_21058,N_20942);
nor U27898 (N_27898,N_21624,N_22231);
and U27899 (N_27899,N_20772,N_20611);
nor U27900 (N_27900,N_21363,N_22171);
nor U27901 (N_27901,N_23571,N_21478);
nand U27902 (N_27902,N_24475,N_24329);
and U27903 (N_27903,N_20320,N_22333);
or U27904 (N_27904,N_21371,N_23134);
nand U27905 (N_27905,N_23166,N_24575);
xnor U27906 (N_27906,N_24442,N_20963);
xnor U27907 (N_27907,N_21831,N_24689);
and U27908 (N_27908,N_20102,N_20095);
and U27909 (N_27909,N_21403,N_24176);
and U27910 (N_27910,N_24058,N_23872);
and U27911 (N_27911,N_20744,N_20925);
and U27912 (N_27912,N_23492,N_21991);
xnor U27913 (N_27913,N_23189,N_20396);
and U27914 (N_27914,N_21584,N_20416);
nor U27915 (N_27915,N_23967,N_22030);
nand U27916 (N_27916,N_23405,N_21724);
nor U27917 (N_27917,N_21678,N_24248);
nand U27918 (N_27918,N_22029,N_21896);
or U27919 (N_27919,N_23880,N_24034);
nor U27920 (N_27920,N_24032,N_22353);
nor U27921 (N_27921,N_20171,N_20606);
or U27922 (N_27922,N_21860,N_22090);
xor U27923 (N_27923,N_20507,N_22882);
nor U27924 (N_27924,N_21776,N_20192);
and U27925 (N_27925,N_24825,N_20164);
nor U27926 (N_27926,N_23026,N_23569);
nand U27927 (N_27927,N_24097,N_20023);
or U27928 (N_27928,N_24567,N_23101);
xor U27929 (N_27929,N_24834,N_20879);
nand U27930 (N_27930,N_21038,N_24491);
or U27931 (N_27931,N_20585,N_20551);
and U27932 (N_27932,N_22385,N_21815);
and U27933 (N_27933,N_20382,N_20710);
nor U27934 (N_27934,N_21562,N_22376);
nand U27935 (N_27935,N_20118,N_24540);
nand U27936 (N_27936,N_24585,N_20584);
or U27937 (N_27937,N_22603,N_22034);
and U27938 (N_27938,N_23039,N_21855);
or U27939 (N_27939,N_24058,N_20492);
nand U27940 (N_27940,N_22385,N_20773);
or U27941 (N_27941,N_21520,N_20880);
nor U27942 (N_27942,N_20067,N_23921);
or U27943 (N_27943,N_24406,N_23160);
nor U27944 (N_27944,N_23434,N_23459);
nand U27945 (N_27945,N_22186,N_21618);
and U27946 (N_27946,N_22333,N_23688);
nand U27947 (N_27947,N_23597,N_24861);
and U27948 (N_27948,N_24089,N_20771);
nand U27949 (N_27949,N_20197,N_22000);
nand U27950 (N_27950,N_22643,N_21629);
xor U27951 (N_27951,N_21494,N_23943);
nor U27952 (N_27952,N_22201,N_22187);
or U27953 (N_27953,N_22493,N_23181);
nand U27954 (N_27954,N_24792,N_23496);
nand U27955 (N_27955,N_22327,N_21730);
nor U27956 (N_27956,N_21770,N_23789);
nand U27957 (N_27957,N_23033,N_21420);
and U27958 (N_27958,N_23830,N_24601);
nor U27959 (N_27959,N_22467,N_20427);
and U27960 (N_27960,N_21688,N_24105);
xnor U27961 (N_27961,N_24166,N_21420);
and U27962 (N_27962,N_24274,N_22966);
nor U27963 (N_27963,N_22970,N_22787);
nand U27964 (N_27964,N_22948,N_20531);
and U27965 (N_27965,N_22293,N_24029);
nor U27966 (N_27966,N_21676,N_21552);
nor U27967 (N_27967,N_23337,N_22986);
or U27968 (N_27968,N_22785,N_24038);
and U27969 (N_27969,N_21580,N_22017);
and U27970 (N_27970,N_24251,N_21832);
nand U27971 (N_27971,N_22632,N_24165);
and U27972 (N_27972,N_22904,N_23663);
and U27973 (N_27973,N_24574,N_21226);
nor U27974 (N_27974,N_21185,N_24440);
nor U27975 (N_27975,N_23177,N_23129);
or U27976 (N_27976,N_23906,N_23587);
or U27977 (N_27977,N_22202,N_20279);
nor U27978 (N_27978,N_24674,N_20155);
xnor U27979 (N_27979,N_21547,N_22089);
nand U27980 (N_27980,N_24457,N_24482);
nor U27981 (N_27981,N_23048,N_22018);
and U27982 (N_27982,N_20577,N_23209);
and U27983 (N_27983,N_22439,N_20415);
or U27984 (N_27984,N_20590,N_24459);
nand U27985 (N_27985,N_20601,N_23928);
or U27986 (N_27986,N_23582,N_23159);
or U27987 (N_27987,N_23193,N_20081);
nor U27988 (N_27988,N_23477,N_23830);
or U27989 (N_27989,N_21161,N_22566);
nand U27990 (N_27990,N_21028,N_24921);
and U27991 (N_27991,N_21428,N_20454);
nand U27992 (N_27992,N_20985,N_20552);
nor U27993 (N_27993,N_24175,N_22721);
and U27994 (N_27994,N_22373,N_24850);
nor U27995 (N_27995,N_22256,N_22073);
and U27996 (N_27996,N_21026,N_23862);
or U27997 (N_27997,N_22952,N_22851);
and U27998 (N_27998,N_20525,N_21628);
or U27999 (N_27999,N_23825,N_22299);
and U28000 (N_28000,N_24624,N_22517);
nor U28001 (N_28001,N_21470,N_24967);
or U28002 (N_28002,N_23264,N_20448);
nor U28003 (N_28003,N_24192,N_21244);
nand U28004 (N_28004,N_23498,N_21843);
nor U28005 (N_28005,N_21054,N_21843);
nand U28006 (N_28006,N_20720,N_20270);
xor U28007 (N_28007,N_22390,N_23366);
xor U28008 (N_28008,N_21315,N_22296);
and U28009 (N_28009,N_22054,N_22406);
or U28010 (N_28010,N_24185,N_24336);
and U28011 (N_28011,N_20064,N_24139);
nor U28012 (N_28012,N_23050,N_21480);
nor U28013 (N_28013,N_20675,N_23170);
nor U28014 (N_28014,N_22031,N_23763);
nor U28015 (N_28015,N_21234,N_22623);
nand U28016 (N_28016,N_20211,N_21031);
nor U28017 (N_28017,N_21155,N_21869);
nor U28018 (N_28018,N_24898,N_21157);
or U28019 (N_28019,N_24690,N_21260);
and U28020 (N_28020,N_20743,N_20647);
nor U28021 (N_28021,N_20874,N_20824);
or U28022 (N_28022,N_21084,N_21321);
and U28023 (N_28023,N_22820,N_24496);
or U28024 (N_28024,N_24856,N_24776);
nor U28025 (N_28025,N_23742,N_20096);
or U28026 (N_28026,N_21784,N_24396);
xor U28027 (N_28027,N_24739,N_23677);
xnor U28028 (N_28028,N_23423,N_24258);
xor U28029 (N_28029,N_23423,N_22090);
and U28030 (N_28030,N_20546,N_21829);
or U28031 (N_28031,N_23835,N_20343);
and U28032 (N_28032,N_20971,N_21938);
nand U28033 (N_28033,N_23900,N_23140);
nor U28034 (N_28034,N_23501,N_22503);
and U28035 (N_28035,N_20028,N_22709);
nor U28036 (N_28036,N_20877,N_20509);
nor U28037 (N_28037,N_21249,N_22812);
nand U28038 (N_28038,N_23255,N_21124);
and U28039 (N_28039,N_23349,N_22455);
nand U28040 (N_28040,N_20557,N_21425);
or U28041 (N_28041,N_22412,N_24293);
and U28042 (N_28042,N_21359,N_24907);
and U28043 (N_28043,N_21962,N_24370);
or U28044 (N_28044,N_24858,N_21997);
nor U28045 (N_28045,N_20591,N_22626);
and U28046 (N_28046,N_20887,N_24981);
nand U28047 (N_28047,N_24441,N_24259);
or U28048 (N_28048,N_21955,N_20609);
nand U28049 (N_28049,N_20577,N_21980);
nor U28050 (N_28050,N_23100,N_21594);
nand U28051 (N_28051,N_21973,N_23124);
or U28052 (N_28052,N_23975,N_24907);
nor U28053 (N_28053,N_24808,N_23687);
or U28054 (N_28054,N_23074,N_22429);
nand U28055 (N_28055,N_21977,N_24613);
and U28056 (N_28056,N_22766,N_23865);
or U28057 (N_28057,N_21980,N_20374);
and U28058 (N_28058,N_23525,N_20693);
xor U28059 (N_28059,N_24896,N_20994);
nor U28060 (N_28060,N_21734,N_20856);
nor U28061 (N_28061,N_21182,N_20200);
nor U28062 (N_28062,N_24495,N_24510);
nand U28063 (N_28063,N_21074,N_20699);
and U28064 (N_28064,N_23351,N_22524);
or U28065 (N_28065,N_21241,N_21437);
xor U28066 (N_28066,N_23974,N_20430);
xor U28067 (N_28067,N_24828,N_20518);
nand U28068 (N_28068,N_21044,N_20678);
and U28069 (N_28069,N_23035,N_24391);
nand U28070 (N_28070,N_21669,N_24786);
and U28071 (N_28071,N_22375,N_23205);
and U28072 (N_28072,N_20000,N_21005);
or U28073 (N_28073,N_22283,N_21242);
or U28074 (N_28074,N_21302,N_20347);
or U28075 (N_28075,N_23825,N_20458);
xor U28076 (N_28076,N_23981,N_22193);
nor U28077 (N_28077,N_20931,N_22187);
nand U28078 (N_28078,N_23163,N_21114);
xnor U28079 (N_28079,N_24266,N_22050);
nand U28080 (N_28080,N_23746,N_22161);
or U28081 (N_28081,N_20738,N_20745);
and U28082 (N_28082,N_20401,N_23806);
nand U28083 (N_28083,N_21039,N_23949);
and U28084 (N_28084,N_24339,N_24048);
nand U28085 (N_28085,N_24299,N_21860);
or U28086 (N_28086,N_24178,N_21027);
xnor U28087 (N_28087,N_23428,N_20701);
and U28088 (N_28088,N_21729,N_20279);
and U28089 (N_28089,N_20123,N_23419);
nand U28090 (N_28090,N_24322,N_21505);
xnor U28091 (N_28091,N_23245,N_24488);
nand U28092 (N_28092,N_20785,N_24680);
and U28093 (N_28093,N_23277,N_21314);
and U28094 (N_28094,N_20499,N_21086);
and U28095 (N_28095,N_20357,N_22403);
or U28096 (N_28096,N_20814,N_23550);
nand U28097 (N_28097,N_21775,N_22466);
xor U28098 (N_28098,N_21880,N_22071);
nand U28099 (N_28099,N_24333,N_21635);
or U28100 (N_28100,N_24668,N_23454);
or U28101 (N_28101,N_24947,N_22091);
nor U28102 (N_28102,N_22299,N_23443);
and U28103 (N_28103,N_23705,N_21298);
nand U28104 (N_28104,N_24161,N_21172);
nor U28105 (N_28105,N_24803,N_22860);
or U28106 (N_28106,N_20866,N_23380);
nand U28107 (N_28107,N_20176,N_22576);
nand U28108 (N_28108,N_23108,N_24346);
and U28109 (N_28109,N_21633,N_23704);
or U28110 (N_28110,N_23138,N_23743);
and U28111 (N_28111,N_20243,N_23701);
xnor U28112 (N_28112,N_21220,N_21310);
nor U28113 (N_28113,N_24537,N_24129);
and U28114 (N_28114,N_21957,N_24220);
and U28115 (N_28115,N_23847,N_20440);
nand U28116 (N_28116,N_24137,N_22164);
and U28117 (N_28117,N_22909,N_23070);
nand U28118 (N_28118,N_21729,N_21378);
and U28119 (N_28119,N_21910,N_23033);
and U28120 (N_28120,N_21593,N_23008);
and U28121 (N_28121,N_21402,N_20445);
nand U28122 (N_28122,N_21429,N_22857);
and U28123 (N_28123,N_21001,N_23416);
or U28124 (N_28124,N_24520,N_23372);
or U28125 (N_28125,N_20265,N_20000);
or U28126 (N_28126,N_23723,N_23513);
and U28127 (N_28127,N_23329,N_20665);
nand U28128 (N_28128,N_22792,N_24187);
or U28129 (N_28129,N_22522,N_24194);
or U28130 (N_28130,N_20802,N_22197);
nand U28131 (N_28131,N_21350,N_21604);
nor U28132 (N_28132,N_22066,N_22866);
nand U28133 (N_28133,N_22297,N_23773);
nor U28134 (N_28134,N_21747,N_21138);
xor U28135 (N_28135,N_21293,N_24368);
nor U28136 (N_28136,N_23723,N_24412);
nor U28137 (N_28137,N_22423,N_23691);
nand U28138 (N_28138,N_24600,N_22213);
and U28139 (N_28139,N_23967,N_20025);
nor U28140 (N_28140,N_20562,N_22254);
or U28141 (N_28141,N_23538,N_24638);
nor U28142 (N_28142,N_20599,N_24081);
nor U28143 (N_28143,N_24209,N_21989);
or U28144 (N_28144,N_20909,N_23761);
nand U28145 (N_28145,N_23040,N_20759);
nor U28146 (N_28146,N_22816,N_21579);
and U28147 (N_28147,N_23087,N_24522);
and U28148 (N_28148,N_24662,N_21897);
and U28149 (N_28149,N_20915,N_24349);
or U28150 (N_28150,N_21977,N_20649);
nor U28151 (N_28151,N_21236,N_22049);
nor U28152 (N_28152,N_24143,N_24067);
nand U28153 (N_28153,N_22277,N_22027);
nor U28154 (N_28154,N_21002,N_20248);
nor U28155 (N_28155,N_21846,N_22142);
or U28156 (N_28156,N_20979,N_24934);
nor U28157 (N_28157,N_20515,N_23348);
nand U28158 (N_28158,N_24170,N_24362);
xnor U28159 (N_28159,N_23719,N_24972);
or U28160 (N_28160,N_22701,N_22375);
and U28161 (N_28161,N_24006,N_22151);
nand U28162 (N_28162,N_24569,N_21645);
and U28163 (N_28163,N_20917,N_24251);
or U28164 (N_28164,N_24496,N_24944);
nand U28165 (N_28165,N_23796,N_21430);
xnor U28166 (N_28166,N_24809,N_22837);
or U28167 (N_28167,N_20860,N_20765);
nor U28168 (N_28168,N_23733,N_21907);
or U28169 (N_28169,N_20016,N_23846);
nor U28170 (N_28170,N_23192,N_21089);
and U28171 (N_28171,N_21964,N_20829);
or U28172 (N_28172,N_23204,N_24639);
and U28173 (N_28173,N_23673,N_24566);
or U28174 (N_28174,N_23816,N_24647);
or U28175 (N_28175,N_23111,N_23628);
xor U28176 (N_28176,N_23571,N_21560);
and U28177 (N_28177,N_22360,N_20362);
nand U28178 (N_28178,N_20336,N_23590);
and U28179 (N_28179,N_24377,N_21222);
xnor U28180 (N_28180,N_21942,N_21286);
and U28181 (N_28181,N_21191,N_22316);
xor U28182 (N_28182,N_23845,N_22585);
xnor U28183 (N_28183,N_20131,N_21969);
nand U28184 (N_28184,N_23872,N_24628);
nor U28185 (N_28185,N_23614,N_24907);
and U28186 (N_28186,N_22191,N_23544);
nand U28187 (N_28187,N_20547,N_24857);
nor U28188 (N_28188,N_24412,N_24724);
xor U28189 (N_28189,N_23679,N_20256);
nand U28190 (N_28190,N_23442,N_20807);
xor U28191 (N_28191,N_23939,N_22137);
xnor U28192 (N_28192,N_21865,N_21566);
nor U28193 (N_28193,N_22067,N_22200);
nor U28194 (N_28194,N_20548,N_20767);
nand U28195 (N_28195,N_24230,N_22448);
nand U28196 (N_28196,N_21918,N_23197);
nor U28197 (N_28197,N_20137,N_24913);
nor U28198 (N_28198,N_21175,N_22969);
and U28199 (N_28199,N_21100,N_23536);
and U28200 (N_28200,N_20276,N_20185);
nor U28201 (N_28201,N_21982,N_23354);
nor U28202 (N_28202,N_21417,N_24658);
and U28203 (N_28203,N_23239,N_21947);
nand U28204 (N_28204,N_20110,N_20806);
or U28205 (N_28205,N_20484,N_21633);
nand U28206 (N_28206,N_23908,N_22856);
nand U28207 (N_28207,N_23540,N_21601);
or U28208 (N_28208,N_20750,N_22657);
nand U28209 (N_28209,N_23300,N_23453);
and U28210 (N_28210,N_23222,N_24841);
xor U28211 (N_28211,N_21393,N_20127);
and U28212 (N_28212,N_20731,N_22042);
or U28213 (N_28213,N_20184,N_23927);
nand U28214 (N_28214,N_21797,N_20312);
and U28215 (N_28215,N_22335,N_22449);
and U28216 (N_28216,N_22526,N_23573);
nand U28217 (N_28217,N_20740,N_22979);
nor U28218 (N_28218,N_23750,N_24212);
or U28219 (N_28219,N_20805,N_20142);
xor U28220 (N_28220,N_21561,N_20298);
xnor U28221 (N_28221,N_24879,N_24944);
xnor U28222 (N_28222,N_23436,N_22567);
nand U28223 (N_28223,N_23617,N_23462);
xnor U28224 (N_28224,N_22050,N_21312);
nand U28225 (N_28225,N_22512,N_22197);
nor U28226 (N_28226,N_22368,N_20968);
nand U28227 (N_28227,N_22266,N_23137);
and U28228 (N_28228,N_24288,N_21204);
xor U28229 (N_28229,N_24790,N_20935);
nand U28230 (N_28230,N_22464,N_24995);
nand U28231 (N_28231,N_20262,N_20197);
nor U28232 (N_28232,N_22467,N_22697);
or U28233 (N_28233,N_22106,N_20944);
or U28234 (N_28234,N_23400,N_21565);
and U28235 (N_28235,N_21028,N_24203);
nor U28236 (N_28236,N_21847,N_22233);
and U28237 (N_28237,N_23704,N_24745);
nand U28238 (N_28238,N_23327,N_20742);
and U28239 (N_28239,N_24342,N_20724);
and U28240 (N_28240,N_24217,N_24541);
or U28241 (N_28241,N_22469,N_21710);
and U28242 (N_28242,N_21652,N_23651);
xor U28243 (N_28243,N_23503,N_24194);
nand U28244 (N_28244,N_20871,N_23607);
xor U28245 (N_28245,N_20220,N_21293);
nand U28246 (N_28246,N_21548,N_20975);
and U28247 (N_28247,N_23978,N_21344);
or U28248 (N_28248,N_23836,N_24561);
or U28249 (N_28249,N_24070,N_22918);
nor U28250 (N_28250,N_20149,N_20012);
nor U28251 (N_28251,N_21128,N_20957);
or U28252 (N_28252,N_23346,N_22059);
nor U28253 (N_28253,N_22805,N_24375);
or U28254 (N_28254,N_20967,N_23369);
or U28255 (N_28255,N_22051,N_22812);
xor U28256 (N_28256,N_23560,N_20695);
nand U28257 (N_28257,N_24711,N_21330);
nor U28258 (N_28258,N_23566,N_24136);
nor U28259 (N_28259,N_22503,N_23701);
nand U28260 (N_28260,N_23133,N_20424);
nand U28261 (N_28261,N_23796,N_23656);
nor U28262 (N_28262,N_22367,N_23807);
nor U28263 (N_28263,N_20887,N_22436);
nand U28264 (N_28264,N_22910,N_20685);
nor U28265 (N_28265,N_24322,N_20271);
nand U28266 (N_28266,N_20096,N_21600);
nor U28267 (N_28267,N_20796,N_20776);
and U28268 (N_28268,N_22443,N_23551);
and U28269 (N_28269,N_20384,N_20986);
xor U28270 (N_28270,N_23714,N_23833);
xor U28271 (N_28271,N_23317,N_21516);
nor U28272 (N_28272,N_20509,N_23593);
and U28273 (N_28273,N_23696,N_21001);
and U28274 (N_28274,N_20681,N_23521);
or U28275 (N_28275,N_21275,N_20738);
nand U28276 (N_28276,N_23904,N_23042);
nand U28277 (N_28277,N_23631,N_23418);
nand U28278 (N_28278,N_20939,N_22731);
nor U28279 (N_28279,N_23475,N_23250);
xnor U28280 (N_28280,N_22651,N_21241);
or U28281 (N_28281,N_20681,N_21776);
or U28282 (N_28282,N_23309,N_21898);
nand U28283 (N_28283,N_24947,N_21227);
xnor U28284 (N_28284,N_23952,N_22438);
or U28285 (N_28285,N_23273,N_24016);
nor U28286 (N_28286,N_22050,N_24135);
nor U28287 (N_28287,N_24071,N_22477);
or U28288 (N_28288,N_22338,N_22412);
nand U28289 (N_28289,N_23529,N_23563);
nor U28290 (N_28290,N_24920,N_20691);
or U28291 (N_28291,N_23713,N_20438);
or U28292 (N_28292,N_22711,N_21783);
nand U28293 (N_28293,N_22821,N_22471);
xor U28294 (N_28294,N_20395,N_22599);
and U28295 (N_28295,N_24713,N_24145);
nand U28296 (N_28296,N_24586,N_20232);
nor U28297 (N_28297,N_20087,N_24129);
nand U28298 (N_28298,N_21451,N_24244);
nor U28299 (N_28299,N_24965,N_22022);
nor U28300 (N_28300,N_20918,N_22155);
and U28301 (N_28301,N_22566,N_22972);
and U28302 (N_28302,N_21808,N_22302);
xor U28303 (N_28303,N_21516,N_21140);
nand U28304 (N_28304,N_20376,N_24647);
and U28305 (N_28305,N_21332,N_20267);
or U28306 (N_28306,N_22792,N_21419);
nand U28307 (N_28307,N_23504,N_22759);
nand U28308 (N_28308,N_22840,N_24614);
nor U28309 (N_28309,N_23747,N_24678);
and U28310 (N_28310,N_20424,N_23569);
xnor U28311 (N_28311,N_20567,N_23360);
nor U28312 (N_28312,N_20683,N_22062);
or U28313 (N_28313,N_22849,N_23685);
nor U28314 (N_28314,N_24044,N_20956);
or U28315 (N_28315,N_21423,N_21213);
or U28316 (N_28316,N_24912,N_24675);
nand U28317 (N_28317,N_22252,N_24479);
nand U28318 (N_28318,N_23558,N_21822);
and U28319 (N_28319,N_20288,N_22459);
and U28320 (N_28320,N_21450,N_23778);
and U28321 (N_28321,N_20061,N_22554);
nand U28322 (N_28322,N_24945,N_22004);
xor U28323 (N_28323,N_22705,N_23195);
nor U28324 (N_28324,N_22954,N_24352);
and U28325 (N_28325,N_20706,N_22968);
or U28326 (N_28326,N_23325,N_22549);
nor U28327 (N_28327,N_22447,N_23314);
and U28328 (N_28328,N_23716,N_20449);
xnor U28329 (N_28329,N_23246,N_24378);
or U28330 (N_28330,N_22881,N_22914);
or U28331 (N_28331,N_21918,N_24740);
nor U28332 (N_28332,N_22947,N_22146);
nor U28333 (N_28333,N_20803,N_23110);
nand U28334 (N_28334,N_22730,N_22246);
or U28335 (N_28335,N_24652,N_21975);
nand U28336 (N_28336,N_23899,N_23873);
or U28337 (N_28337,N_24349,N_21255);
nand U28338 (N_28338,N_23467,N_20834);
nor U28339 (N_28339,N_23368,N_23119);
and U28340 (N_28340,N_22821,N_21830);
nor U28341 (N_28341,N_24963,N_23587);
nor U28342 (N_28342,N_24162,N_23680);
nor U28343 (N_28343,N_20487,N_24424);
and U28344 (N_28344,N_22724,N_23577);
nor U28345 (N_28345,N_22170,N_22991);
nand U28346 (N_28346,N_21394,N_22217);
nor U28347 (N_28347,N_24769,N_23180);
nor U28348 (N_28348,N_21141,N_23446);
nand U28349 (N_28349,N_23626,N_21861);
and U28350 (N_28350,N_22017,N_24505);
xnor U28351 (N_28351,N_21861,N_20175);
xor U28352 (N_28352,N_21011,N_23095);
nand U28353 (N_28353,N_24786,N_20812);
or U28354 (N_28354,N_21082,N_24545);
nor U28355 (N_28355,N_21940,N_20514);
nor U28356 (N_28356,N_20634,N_24463);
and U28357 (N_28357,N_24615,N_22375);
and U28358 (N_28358,N_22988,N_22802);
nor U28359 (N_28359,N_23231,N_23504);
nand U28360 (N_28360,N_24877,N_21754);
nand U28361 (N_28361,N_21386,N_22282);
nor U28362 (N_28362,N_20586,N_20911);
and U28363 (N_28363,N_22161,N_20647);
and U28364 (N_28364,N_21332,N_22745);
nor U28365 (N_28365,N_24372,N_21517);
nor U28366 (N_28366,N_24192,N_24206);
or U28367 (N_28367,N_23133,N_20255);
or U28368 (N_28368,N_22339,N_20886);
and U28369 (N_28369,N_23039,N_22124);
and U28370 (N_28370,N_22972,N_24410);
nor U28371 (N_28371,N_21565,N_24635);
or U28372 (N_28372,N_20457,N_24995);
nor U28373 (N_28373,N_22136,N_22651);
or U28374 (N_28374,N_22094,N_24067);
or U28375 (N_28375,N_20424,N_24028);
and U28376 (N_28376,N_23008,N_20782);
nand U28377 (N_28377,N_24876,N_23693);
xor U28378 (N_28378,N_22528,N_23465);
and U28379 (N_28379,N_24658,N_24510);
and U28380 (N_28380,N_20959,N_22414);
nor U28381 (N_28381,N_22231,N_20243);
and U28382 (N_28382,N_20459,N_20092);
or U28383 (N_28383,N_22418,N_22680);
nand U28384 (N_28384,N_23547,N_21251);
or U28385 (N_28385,N_23728,N_22857);
nand U28386 (N_28386,N_24566,N_23850);
nand U28387 (N_28387,N_21582,N_22983);
nand U28388 (N_28388,N_21004,N_21253);
or U28389 (N_28389,N_22791,N_21359);
or U28390 (N_28390,N_23434,N_20548);
xor U28391 (N_28391,N_21761,N_21919);
nor U28392 (N_28392,N_23943,N_22060);
and U28393 (N_28393,N_22769,N_20125);
and U28394 (N_28394,N_24937,N_24476);
nor U28395 (N_28395,N_20094,N_22494);
or U28396 (N_28396,N_20099,N_22075);
or U28397 (N_28397,N_23811,N_20576);
nand U28398 (N_28398,N_24498,N_22273);
nor U28399 (N_28399,N_20701,N_20625);
nand U28400 (N_28400,N_23618,N_24305);
xor U28401 (N_28401,N_23003,N_24038);
and U28402 (N_28402,N_21629,N_21279);
or U28403 (N_28403,N_20741,N_21267);
or U28404 (N_28404,N_22590,N_21577);
or U28405 (N_28405,N_24928,N_23758);
or U28406 (N_28406,N_23640,N_22335);
nand U28407 (N_28407,N_22176,N_21381);
nand U28408 (N_28408,N_21934,N_20658);
nand U28409 (N_28409,N_23279,N_20660);
and U28410 (N_28410,N_22479,N_21479);
and U28411 (N_28411,N_21923,N_22689);
nor U28412 (N_28412,N_21003,N_24316);
xor U28413 (N_28413,N_23512,N_22573);
nor U28414 (N_28414,N_24461,N_24627);
nand U28415 (N_28415,N_21248,N_23735);
xnor U28416 (N_28416,N_23025,N_22314);
or U28417 (N_28417,N_20145,N_22853);
nor U28418 (N_28418,N_24422,N_23640);
nand U28419 (N_28419,N_23130,N_20189);
nor U28420 (N_28420,N_22284,N_24777);
nor U28421 (N_28421,N_21048,N_22479);
and U28422 (N_28422,N_20440,N_21143);
or U28423 (N_28423,N_22496,N_24587);
nand U28424 (N_28424,N_20285,N_23844);
nand U28425 (N_28425,N_23477,N_20502);
and U28426 (N_28426,N_20072,N_23605);
or U28427 (N_28427,N_22202,N_22508);
and U28428 (N_28428,N_22856,N_22287);
xor U28429 (N_28429,N_24507,N_20510);
xnor U28430 (N_28430,N_22815,N_23119);
and U28431 (N_28431,N_21291,N_20106);
nor U28432 (N_28432,N_22925,N_20281);
or U28433 (N_28433,N_24560,N_24673);
nand U28434 (N_28434,N_20278,N_21211);
nand U28435 (N_28435,N_22020,N_23011);
xor U28436 (N_28436,N_20385,N_22908);
nor U28437 (N_28437,N_21189,N_20842);
or U28438 (N_28438,N_21155,N_24994);
or U28439 (N_28439,N_24169,N_24265);
or U28440 (N_28440,N_22268,N_24524);
or U28441 (N_28441,N_21768,N_23213);
nand U28442 (N_28442,N_20328,N_22705);
and U28443 (N_28443,N_21783,N_22986);
and U28444 (N_28444,N_24534,N_22568);
nand U28445 (N_28445,N_24691,N_20488);
or U28446 (N_28446,N_21146,N_22015);
nor U28447 (N_28447,N_22948,N_20511);
or U28448 (N_28448,N_24808,N_21106);
xnor U28449 (N_28449,N_22840,N_22090);
xnor U28450 (N_28450,N_24160,N_20681);
and U28451 (N_28451,N_22977,N_24775);
or U28452 (N_28452,N_24864,N_24663);
nand U28453 (N_28453,N_24681,N_24789);
nor U28454 (N_28454,N_24371,N_22666);
nor U28455 (N_28455,N_23458,N_24040);
nor U28456 (N_28456,N_24700,N_24624);
and U28457 (N_28457,N_20543,N_22583);
nor U28458 (N_28458,N_22932,N_23317);
and U28459 (N_28459,N_23632,N_22747);
nor U28460 (N_28460,N_20973,N_24729);
or U28461 (N_28461,N_23018,N_24644);
or U28462 (N_28462,N_20725,N_23646);
xnor U28463 (N_28463,N_20423,N_24377);
and U28464 (N_28464,N_21616,N_23665);
or U28465 (N_28465,N_24290,N_22526);
nor U28466 (N_28466,N_20562,N_20764);
and U28467 (N_28467,N_20941,N_23943);
nand U28468 (N_28468,N_22619,N_24536);
or U28469 (N_28469,N_24365,N_21863);
xor U28470 (N_28470,N_20662,N_22520);
or U28471 (N_28471,N_20475,N_22132);
nand U28472 (N_28472,N_22321,N_24447);
or U28473 (N_28473,N_21150,N_22347);
or U28474 (N_28474,N_23679,N_20527);
nand U28475 (N_28475,N_20505,N_24621);
xnor U28476 (N_28476,N_21712,N_21273);
nor U28477 (N_28477,N_22290,N_20423);
nand U28478 (N_28478,N_22205,N_23930);
nor U28479 (N_28479,N_21822,N_20559);
or U28480 (N_28480,N_23280,N_23544);
nand U28481 (N_28481,N_23400,N_20506);
or U28482 (N_28482,N_20773,N_23943);
nor U28483 (N_28483,N_21508,N_20618);
nand U28484 (N_28484,N_21032,N_23908);
nor U28485 (N_28485,N_20254,N_23576);
nor U28486 (N_28486,N_22637,N_22422);
nor U28487 (N_28487,N_22173,N_20845);
or U28488 (N_28488,N_23620,N_20917);
or U28489 (N_28489,N_24426,N_23551);
xor U28490 (N_28490,N_23037,N_24379);
or U28491 (N_28491,N_22498,N_24163);
nand U28492 (N_28492,N_21175,N_22057);
nand U28493 (N_28493,N_21997,N_20806);
nor U28494 (N_28494,N_21411,N_21951);
nand U28495 (N_28495,N_21332,N_23222);
or U28496 (N_28496,N_22304,N_23370);
nand U28497 (N_28497,N_22081,N_24317);
xor U28498 (N_28498,N_21504,N_21017);
nor U28499 (N_28499,N_24071,N_24106);
or U28500 (N_28500,N_20016,N_22415);
nor U28501 (N_28501,N_21053,N_23162);
nand U28502 (N_28502,N_24152,N_23951);
and U28503 (N_28503,N_23125,N_23779);
nor U28504 (N_28504,N_24283,N_24828);
and U28505 (N_28505,N_23593,N_23458);
nor U28506 (N_28506,N_22809,N_24902);
xor U28507 (N_28507,N_24430,N_21937);
and U28508 (N_28508,N_22546,N_24174);
xnor U28509 (N_28509,N_23185,N_23867);
nor U28510 (N_28510,N_21581,N_23021);
xor U28511 (N_28511,N_22083,N_23131);
xnor U28512 (N_28512,N_23255,N_22303);
nand U28513 (N_28513,N_21290,N_23665);
or U28514 (N_28514,N_23639,N_21520);
or U28515 (N_28515,N_24881,N_24713);
nand U28516 (N_28516,N_20832,N_22480);
nor U28517 (N_28517,N_20076,N_20293);
and U28518 (N_28518,N_21994,N_23458);
nor U28519 (N_28519,N_20245,N_22546);
xnor U28520 (N_28520,N_24117,N_22619);
nor U28521 (N_28521,N_22477,N_24641);
or U28522 (N_28522,N_22198,N_22787);
nand U28523 (N_28523,N_22681,N_21932);
and U28524 (N_28524,N_20573,N_23446);
xor U28525 (N_28525,N_23018,N_24654);
and U28526 (N_28526,N_20995,N_23994);
and U28527 (N_28527,N_23338,N_20655);
or U28528 (N_28528,N_23220,N_21153);
nor U28529 (N_28529,N_20132,N_24219);
nand U28530 (N_28530,N_22224,N_21129);
nor U28531 (N_28531,N_23209,N_22134);
nand U28532 (N_28532,N_24445,N_24152);
nor U28533 (N_28533,N_20183,N_22649);
nand U28534 (N_28534,N_23026,N_21792);
nor U28535 (N_28535,N_22918,N_23729);
and U28536 (N_28536,N_22025,N_22027);
xor U28537 (N_28537,N_20488,N_22541);
and U28538 (N_28538,N_22581,N_23883);
or U28539 (N_28539,N_21088,N_22009);
or U28540 (N_28540,N_20615,N_21620);
nor U28541 (N_28541,N_20923,N_24389);
or U28542 (N_28542,N_21653,N_21242);
and U28543 (N_28543,N_24213,N_22655);
or U28544 (N_28544,N_23329,N_23090);
and U28545 (N_28545,N_23811,N_20058);
and U28546 (N_28546,N_22480,N_24077);
and U28547 (N_28547,N_22154,N_21881);
nand U28548 (N_28548,N_20895,N_22127);
or U28549 (N_28549,N_24452,N_23119);
or U28550 (N_28550,N_22092,N_23606);
or U28551 (N_28551,N_21735,N_23044);
and U28552 (N_28552,N_21931,N_22693);
and U28553 (N_28553,N_21160,N_20900);
nor U28554 (N_28554,N_20474,N_24126);
nand U28555 (N_28555,N_22794,N_21648);
nand U28556 (N_28556,N_23083,N_23413);
nor U28557 (N_28557,N_24370,N_23723);
or U28558 (N_28558,N_20883,N_24558);
nand U28559 (N_28559,N_21956,N_22116);
xor U28560 (N_28560,N_23379,N_20821);
nand U28561 (N_28561,N_20635,N_21899);
nand U28562 (N_28562,N_20751,N_21590);
and U28563 (N_28563,N_24244,N_21069);
or U28564 (N_28564,N_20756,N_20173);
or U28565 (N_28565,N_23488,N_22108);
or U28566 (N_28566,N_22976,N_22096);
or U28567 (N_28567,N_20739,N_22395);
nand U28568 (N_28568,N_21212,N_24901);
xor U28569 (N_28569,N_21023,N_22434);
and U28570 (N_28570,N_21100,N_22284);
or U28571 (N_28571,N_24779,N_23672);
or U28572 (N_28572,N_21355,N_23368);
nand U28573 (N_28573,N_23739,N_20977);
nand U28574 (N_28574,N_21580,N_22967);
or U28575 (N_28575,N_24839,N_24338);
nor U28576 (N_28576,N_21388,N_21287);
xnor U28577 (N_28577,N_21857,N_23566);
or U28578 (N_28578,N_24236,N_20115);
nand U28579 (N_28579,N_23978,N_20691);
xnor U28580 (N_28580,N_23774,N_21906);
nand U28581 (N_28581,N_24487,N_20769);
nor U28582 (N_28582,N_24452,N_20568);
nor U28583 (N_28583,N_24513,N_22229);
or U28584 (N_28584,N_20142,N_21812);
and U28585 (N_28585,N_21890,N_24834);
nor U28586 (N_28586,N_23279,N_20453);
and U28587 (N_28587,N_21043,N_21882);
nand U28588 (N_28588,N_24638,N_23363);
nor U28589 (N_28589,N_22282,N_24770);
or U28590 (N_28590,N_21814,N_20843);
nor U28591 (N_28591,N_21718,N_21134);
or U28592 (N_28592,N_20448,N_21573);
or U28593 (N_28593,N_22803,N_23976);
or U28594 (N_28594,N_20337,N_20166);
nand U28595 (N_28595,N_22162,N_23315);
nand U28596 (N_28596,N_20482,N_20314);
and U28597 (N_28597,N_23728,N_20279);
nor U28598 (N_28598,N_24447,N_24297);
and U28599 (N_28599,N_22334,N_21905);
nor U28600 (N_28600,N_22251,N_21478);
or U28601 (N_28601,N_22967,N_24987);
nand U28602 (N_28602,N_24105,N_20091);
xnor U28603 (N_28603,N_23570,N_21497);
nor U28604 (N_28604,N_20749,N_21393);
nand U28605 (N_28605,N_24722,N_20652);
nand U28606 (N_28606,N_22348,N_22768);
or U28607 (N_28607,N_22962,N_24549);
nor U28608 (N_28608,N_22739,N_23504);
or U28609 (N_28609,N_20497,N_21326);
and U28610 (N_28610,N_23609,N_22005);
and U28611 (N_28611,N_23039,N_23611);
or U28612 (N_28612,N_24390,N_22375);
xnor U28613 (N_28613,N_22652,N_21871);
and U28614 (N_28614,N_21491,N_20825);
nor U28615 (N_28615,N_23851,N_22641);
or U28616 (N_28616,N_23850,N_21408);
nand U28617 (N_28617,N_22020,N_23685);
xor U28618 (N_28618,N_23136,N_20137);
and U28619 (N_28619,N_20487,N_23226);
nor U28620 (N_28620,N_22311,N_24762);
nand U28621 (N_28621,N_24409,N_23800);
nand U28622 (N_28622,N_24632,N_23031);
nand U28623 (N_28623,N_20834,N_21685);
or U28624 (N_28624,N_24540,N_20191);
and U28625 (N_28625,N_24026,N_23544);
and U28626 (N_28626,N_22682,N_22092);
and U28627 (N_28627,N_24856,N_24457);
or U28628 (N_28628,N_23474,N_23387);
nor U28629 (N_28629,N_24873,N_22295);
and U28630 (N_28630,N_24574,N_20204);
nand U28631 (N_28631,N_22385,N_24667);
or U28632 (N_28632,N_21803,N_24569);
nor U28633 (N_28633,N_24783,N_22767);
nor U28634 (N_28634,N_24369,N_20034);
nor U28635 (N_28635,N_24688,N_20236);
nand U28636 (N_28636,N_24052,N_23195);
or U28637 (N_28637,N_21081,N_21189);
and U28638 (N_28638,N_20423,N_24739);
nor U28639 (N_28639,N_23382,N_24705);
xnor U28640 (N_28640,N_24188,N_23459);
and U28641 (N_28641,N_24964,N_24228);
nand U28642 (N_28642,N_23285,N_21369);
or U28643 (N_28643,N_23079,N_24829);
nand U28644 (N_28644,N_22996,N_21439);
nor U28645 (N_28645,N_24157,N_23557);
nand U28646 (N_28646,N_24423,N_21697);
nand U28647 (N_28647,N_21201,N_24679);
and U28648 (N_28648,N_20186,N_21978);
nand U28649 (N_28649,N_24700,N_20410);
or U28650 (N_28650,N_24051,N_24475);
nand U28651 (N_28651,N_22260,N_23602);
or U28652 (N_28652,N_24265,N_22528);
xor U28653 (N_28653,N_23607,N_23810);
or U28654 (N_28654,N_24092,N_24858);
nand U28655 (N_28655,N_20726,N_20280);
nor U28656 (N_28656,N_24038,N_23191);
nand U28657 (N_28657,N_23791,N_23798);
nand U28658 (N_28658,N_20627,N_23264);
and U28659 (N_28659,N_20956,N_22903);
nand U28660 (N_28660,N_24203,N_24711);
or U28661 (N_28661,N_20179,N_22281);
nand U28662 (N_28662,N_23058,N_22431);
nor U28663 (N_28663,N_24368,N_20220);
xor U28664 (N_28664,N_21331,N_20728);
nor U28665 (N_28665,N_22721,N_20744);
nand U28666 (N_28666,N_22685,N_21539);
and U28667 (N_28667,N_21124,N_23401);
and U28668 (N_28668,N_24051,N_24748);
or U28669 (N_28669,N_24111,N_24178);
nand U28670 (N_28670,N_21154,N_21980);
nand U28671 (N_28671,N_21861,N_23641);
nor U28672 (N_28672,N_22442,N_20612);
or U28673 (N_28673,N_24366,N_21842);
nand U28674 (N_28674,N_20376,N_20726);
nand U28675 (N_28675,N_20774,N_24967);
nor U28676 (N_28676,N_20978,N_24420);
nor U28677 (N_28677,N_20802,N_21231);
nand U28678 (N_28678,N_21546,N_23255);
nor U28679 (N_28679,N_22240,N_23337);
xor U28680 (N_28680,N_24504,N_24751);
xnor U28681 (N_28681,N_22065,N_21011);
nand U28682 (N_28682,N_24919,N_24332);
nor U28683 (N_28683,N_21369,N_21968);
and U28684 (N_28684,N_23258,N_22444);
and U28685 (N_28685,N_21417,N_20139);
and U28686 (N_28686,N_22696,N_24681);
nor U28687 (N_28687,N_23033,N_23078);
and U28688 (N_28688,N_24071,N_20832);
or U28689 (N_28689,N_23183,N_24811);
nor U28690 (N_28690,N_24331,N_23480);
nand U28691 (N_28691,N_23222,N_23943);
and U28692 (N_28692,N_24233,N_24058);
and U28693 (N_28693,N_21996,N_21990);
nor U28694 (N_28694,N_22140,N_24189);
and U28695 (N_28695,N_23939,N_23715);
nand U28696 (N_28696,N_23160,N_21389);
or U28697 (N_28697,N_20118,N_21385);
or U28698 (N_28698,N_22125,N_24159);
and U28699 (N_28699,N_22645,N_22463);
or U28700 (N_28700,N_24702,N_21948);
nand U28701 (N_28701,N_22445,N_23304);
and U28702 (N_28702,N_21825,N_23468);
xor U28703 (N_28703,N_22733,N_22875);
nor U28704 (N_28704,N_23663,N_20146);
xor U28705 (N_28705,N_22725,N_20486);
nor U28706 (N_28706,N_21441,N_20154);
nor U28707 (N_28707,N_20364,N_23952);
nor U28708 (N_28708,N_21688,N_24568);
nor U28709 (N_28709,N_24931,N_24783);
xor U28710 (N_28710,N_21627,N_20226);
and U28711 (N_28711,N_22427,N_20337);
nand U28712 (N_28712,N_24784,N_21847);
or U28713 (N_28713,N_22108,N_21991);
nor U28714 (N_28714,N_21975,N_20286);
nand U28715 (N_28715,N_24429,N_22342);
nand U28716 (N_28716,N_21972,N_21030);
or U28717 (N_28717,N_24003,N_23652);
nand U28718 (N_28718,N_22214,N_24745);
nor U28719 (N_28719,N_21896,N_20285);
and U28720 (N_28720,N_23349,N_22304);
or U28721 (N_28721,N_23485,N_21807);
nor U28722 (N_28722,N_22527,N_20069);
xnor U28723 (N_28723,N_22542,N_24520);
nand U28724 (N_28724,N_21737,N_23482);
nor U28725 (N_28725,N_21604,N_22120);
or U28726 (N_28726,N_23813,N_23405);
xnor U28727 (N_28727,N_22720,N_20199);
and U28728 (N_28728,N_23105,N_20194);
xor U28729 (N_28729,N_21386,N_23871);
nor U28730 (N_28730,N_23577,N_20139);
or U28731 (N_28731,N_20990,N_24480);
nand U28732 (N_28732,N_22021,N_23634);
and U28733 (N_28733,N_20225,N_21204);
xor U28734 (N_28734,N_20160,N_21778);
and U28735 (N_28735,N_20810,N_22086);
xnor U28736 (N_28736,N_20289,N_24965);
nor U28737 (N_28737,N_23604,N_24491);
or U28738 (N_28738,N_20491,N_24740);
and U28739 (N_28739,N_23203,N_21848);
and U28740 (N_28740,N_24680,N_22808);
or U28741 (N_28741,N_21191,N_21361);
nand U28742 (N_28742,N_21601,N_20208);
or U28743 (N_28743,N_24032,N_21514);
and U28744 (N_28744,N_21133,N_23190);
nor U28745 (N_28745,N_23306,N_22466);
or U28746 (N_28746,N_24222,N_21942);
and U28747 (N_28747,N_20466,N_21317);
nor U28748 (N_28748,N_24282,N_22410);
nand U28749 (N_28749,N_20560,N_22403);
xor U28750 (N_28750,N_24978,N_21198);
xnor U28751 (N_28751,N_23225,N_23132);
and U28752 (N_28752,N_23275,N_24918);
and U28753 (N_28753,N_23245,N_23370);
nor U28754 (N_28754,N_21249,N_23741);
nor U28755 (N_28755,N_21383,N_21396);
nand U28756 (N_28756,N_23192,N_20275);
or U28757 (N_28757,N_21308,N_23601);
and U28758 (N_28758,N_21063,N_24925);
nand U28759 (N_28759,N_22240,N_20591);
nor U28760 (N_28760,N_21054,N_21829);
or U28761 (N_28761,N_23420,N_23081);
nor U28762 (N_28762,N_24520,N_21547);
nand U28763 (N_28763,N_20793,N_24005);
xor U28764 (N_28764,N_21519,N_20606);
and U28765 (N_28765,N_21975,N_24436);
nand U28766 (N_28766,N_22063,N_23597);
and U28767 (N_28767,N_24945,N_22782);
or U28768 (N_28768,N_21631,N_22960);
or U28769 (N_28769,N_22456,N_23250);
or U28770 (N_28770,N_22305,N_24815);
or U28771 (N_28771,N_20022,N_20119);
and U28772 (N_28772,N_22686,N_21013);
nor U28773 (N_28773,N_21678,N_21748);
nor U28774 (N_28774,N_22174,N_20188);
nor U28775 (N_28775,N_23631,N_23811);
and U28776 (N_28776,N_23409,N_21630);
nor U28777 (N_28777,N_24468,N_22779);
nand U28778 (N_28778,N_22052,N_23874);
nand U28779 (N_28779,N_21855,N_24820);
or U28780 (N_28780,N_21286,N_24429);
and U28781 (N_28781,N_21566,N_21240);
or U28782 (N_28782,N_21721,N_20297);
nand U28783 (N_28783,N_24983,N_24702);
nand U28784 (N_28784,N_23891,N_24842);
nand U28785 (N_28785,N_22244,N_23485);
and U28786 (N_28786,N_23196,N_21798);
nand U28787 (N_28787,N_21291,N_24404);
nand U28788 (N_28788,N_24418,N_24607);
nor U28789 (N_28789,N_24822,N_24200);
nor U28790 (N_28790,N_24322,N_21448);
nand U28791 (N_28791,N_21637,N_24692);
nand U28792 (N_28792,N_23406,N_20489);
nor U28793 (N_28793,N_23925,N_21102);
nand U28794 (N_28794,N_24264,N_24938);
nor U28795 (N_28795,N_23710,N_23658);
and U28796 (N_28796,N_20286,N_23096);
and U28797 (N_28797,N_23823,N_20999);
nand U28798 (N_28798,N_23440,N_24307);
nor U28799 (N_28799,N_24238,N_23037);
nor U28800 (N_28800,N_22364,N_24534);
xnor U28801 (N_28801,N_24674,N_20553);
or U28802 (N_28802,N_21858,N_22445);
nand U28803 (N_28803,N_20384,N_21818);
nand U28804 (N_28804,N_24193,N_21307);
xor U28805 (N_28805,N_21992,N_23892);
xor U28806 (N_28806,N_23810,N_23624);
and U28807 (N_28807,N_22947,N_22124);
or U28808 (N_28808,N_24996,N_22341);
and U28809 (N_28809,N_21482,N_24375);
nand U28810 (N_28810,N_23100,N_20906);
or U28811 (N_28811,N_24423,N_20303);
or U28812 (N_28812,N_22706,N_21772);
nand U28813 (N_28813,N_21522,N_20077);
or U28814 (N_28814,N_23803,N_21617);
or U28815 (N_28815,N_21534,N_21544);
nand U28816 (N_28816,N_20492,N_24667);
xor U28817 (N_28817,N_23717,N_21706);
nand U28818 (N_28818,N_24394,N_20959);
or U28819 (N_28819,N_21209,N_24262);
nand U28820 (N_28820,N_24335,N_24628);
or U28821 (N_28821,N_24960,N_21461);
and U28822 (N_28822,N_21407,N_23776);
nand U28823 (N_28823,N_22747,N_21210);
or U28824 (N_28824,N_22156,N_22767);
xnor U28825 (N_28825,N_23471,N_22844);
or U28826 (N_28826,N_23827,N_21053);
nand U28827 (N_28827,N_22374,N_22586);
or U28828 (N_28828,N_21536,N_20323);
or U28829 (N_28829,N_22054,N_22127);
nor U28830 (N_28830,N_21175,N_23405);
nor U28831 (N_28831,N_21166,N_21254);
nand U28832 (N_28832,N_21810,N_21922);
nand U28833 (N_28833,N_22138,N_23217);
nand U28834 (N_28834,N_21055,N_20944);
and U28835 (N_28835,N_21875,N_20389);
or U28836 (N_28836,N_20546,N_22105);
nor U28837 (N_28837,N_22794,N_24551);
xnor U28838 (N_28838,N_22212,N_24966);
nand U28839 (N_28839,N_22617,N_24800);
or U28840 (N_28840,N_23370,N_23139);
nand U28841 (N_28841,N_22865,N_22850);
xnor U28842 (N_28842,N_22502,N_21227);
or U28843 (N_28843,N_22863,N_22915);
or U28844 (N_28844,N_22263,N_22340);
nand U28845 (N_28845,N_21345,N_23754);
or U28846 (N_28846,N_20633,N_21503);
and U28847 (N_28847,N_21342,N_21103);
or U28848 (N_28848,N_24941,N_24975);
xnor U28849 (N_28849,N_21928,N_21256);
nor U28850 (N_28850,N_21211,N_24142);
nor U28851 (N_28851,N_21225,N_20954);
or U28852 (N_28852,N_24431,N_20836);
or U28853 (N_28853,N_20536,N_21130);
or U28854 (N_28854,N_23379,N_23397);
nand U28855 (N_28855,N_23799,N_22474);
or U28856 (N_28856,N_24159,N_23066);
and U28857 (N_28857,N_20421,N_24991);
nor U28858 (N_28858,N_24467,N_22288);
and U28859 (N_28859,N_24473,N_24224);
or U28860 (N_28860,N_22103,N_20244);
and U28861 (N_28861,N_22003,N_22354);
nor U28862 (N_28862,N_22745,N_23436);
and U28863 (N_28863,N_21354,N_20255);
nand U28864 (N_28864,N_21233,N_23947);
xnor U28865 (N_28865,N_24317,N_20848);
nor U28866 (N_28866,N_22580,N_22334);
xnor U28867 (N_28867,N_20842,N_22430);
and U28868 (N_28868,N_21437,N_20005);
xnor U28869 (N_28869,N_22566,N_24976);
and U28870 (N_28870,N_21718,N_24810);
nand U28871 (N_28871,N_22474,N_21282);
or U28872 (N_28872,N_23794,N_24342);
and U28873 (N_28873,N_24101,N_20181);
nor U28874 (N_28874,N_20212,N_21959);
or U28875 (N_28875,N_23090,N_21673);
or U28876 (N_28876,N_23301,N_20706);
nand U28877 (N_28877,N_23863,N_20594);
xor U28878 (N_28878,N_23567,N_24708);
nand U28879 (N_28879,N_21511,N_22820);
or U28880 (N_28880,N_21861,N_22725);
and U28881 (N_28881,N_23709,N_24273);
and U28882 (N_28882,N_22229,N_24302);
xor U28883 (N_28883,N_22511,N_20643);
and U28884 (N_28884,N_21903,N_20782);
nor U28885 (N_28885,N_24975,N_23610);
or U28886 (N_28886,N_23587,N_21292);
and U28887 (N_28887,N_20465,N_23090);
nand U28888 (N_28888,N_24130,N_23819);
and U28889 (N_28889,N_21016,N_22050);
and U28890 (N_28890,N_20086,N_23816);
nand U28891 (N_28891,N_23346,N_20778);
or U28892 (N_28892,N_23759,N_24121);
nor U28893 (N_28893,N_24975,N_23830);
nand U28894 (N_28894,N_24570,N_20574);
or U28895 (N_28895,N_21056,N_21052);
or U28896 (N_28896,N_20107,N_21402);
or U28897 (N_28897,N_21187,N_21635);
or U28898 (N_28898,N_20738,N_21302);
xnor U28899 (N_28899,N_23899,N_23013);
or U28900 (N_28900,N_24532,N_23672);
nor U28901 (N_28901,N_24017,N_22890);
nand U28902 (N_28902,N_24814,N_22512);
nor U28903 (N_28903,N_20799,N_20259);
xnor U28904 (N_28904,N_24459,N_24609);
nand U28905 (N_28905,N_22819,N_22690);
and U28906 (N_28906,N_22199,N_24493);
xor U28907 (N_28907,N_23908,N_21359);
or U28908 (N_28908,N_20224,N_24238);
nand U28909 (N_28909,N_24128,N_22645);
or U28910 (N_28910,N_22359,N_22522);
nor U28911 (N_28911,N_23165,N_20558);
and U28912 (N_28912,N_21268,N_20220);
and U28913 (N_28913,N_23441,N_24908);
nand U28914 (N_28914,N_22531,N_23820);
nor U28915 (N_28915,N_21730,N_22130);
or U28916 (N_28916,N_22931,N_22976);
nand U28917 (N_28917,N_24348,N_24162);
and U28918 (N_28918,N_20118,N_24136);
and U28919 (N_28919,N_23273,N_24701);
and U28920 (N_28920,N_20380,N_23154);
or U28921 (N_28921,N_21150,N_23812);
nor U28922 (N_28922,N_22808,N_21475);
nor U28923 (N_28923,N_21964,N_21969);
and U28924 (N_28924,N_21309,N_24925);
nor U28925 (N_28925,N_21894,N_23922);
and U28926 (N_28926,N_20065,N_23934);
or U28927 (N_28927,N_22083,N_22274);
and U28928 (N_28928,N_23436,N_22737);
nor U28929 (N_28929,N_21466,N_23814);
and U28930 (N_28930,N_24027,N_24697);
xnor U28931 (N_28931,N_24875,N_23054);
or U28932 (N_28932,N_24276,N_21200);
nor U28933 (N_28933,N_22735,N_22211);
and U28934 (N_28934,N_22959,N_24460);
or U28935 (N_28935,N_21901,N_21974);
nand U28936 (N_28936,N_20751,N_24479);
nand U28937 (N_28937,N_21691,N_21201);
and U28938 (N_28938,N_24531,N_20916);
nor U28939 (N_28939,N_23232,N_22701);
nand U28940 (N_28940,N_23598,N_20363);
nor U28941 (N_28941,N_21359,N_23119);
and U28942 (N_28942,N_23064,N_24991);
nand U28943 (N_28943,N_20548,N_22856);
nor U28944 (N_28944,N_22420,N_23946);
and U28945 (N_28945,N_20379,N_22445);
or U28946 (N_28946,N_22558,N_20641);
and U28947 (N_28947,N_23893,N_21852);
and U28948 (N_28948,N_23641,N_22100);
and U28949 (N_28949,N_22073,N_20711);
xnor U28950 (N_28950,N_23870,N_22194);
nand U28951 (N_28951,N_22842,N_21781);
nand U28952 (N_28952,N_23061,N_23492);
nor U28953 (N_28953,N_23896,N_24735);
or U28954 (N_28954,N_20814,N_20666);
and U28955 (N_28955,N_23698,N_22861);
and U28956 (N_28956,N_20843,N_20102);
nand U28957 (N_28957,N_23862,N_24366);
nor U28958 (N_28958,N_23153,N_23921);
nand U28959 (N_28959,N_23164,N_22165);
and U28960 (N_28960,N_23352,N_24116);
and U28961 (N_28961,N_20720,N_24758);
nand U28962 (N_28962,N_23402,N_20079);
and U28963 (N_28963,N_23457,N_21993);
nor U28964 (N_28964,N_21027,N_20544);
nor U28965 (N_28965,N_21736,N_23259);
nor U28966 (N_28966,N_24646,N_23919);
xnor U28967 (N_28967,N_22030,N_23323);
xnor U28968 (N_28968,N_24934,N_22755);
or U28969 (N_28969,N_23600,N_20628);
xnor U28970 (N_28970,N_20848,N_21922);
or U28971 (N_28971,N_22101,N_24333);
nand U28972 (N_28972,N_21543,N_23070);
or U28973 (N_28973,N_23803,N_22607);
xor U28974 (N_28974,N_20339,N_21892);
xnor U28975 (N_28975,N_24753,N_23468);
nand U28976 (N_28976,N_22890,N_24764);
nand U28977 (N_28977,N_22141,N_20256);
and U28978 (N_28978,N_24972,N_21142);
nor U28979 (N_28979,N_20967,N_22210);
or U28980 (N_28980,N_23556,N_22493);
nand U28981 (N_28981,N_22760,N_20631);
or U28982 (N_28982,N_20474,N_22564);
and U28983 (N_28983,N_20327,N_23691);
or U28984 (N_28984,N_24552,N_21498);
xnor U28985 (N_28985,N_22357,N_21970);
and U28986 (N_28986,N_22624,N_21646);
or U28987 (N_28987,N_20447,N_24592);
nor U28988 (N_28988,N_23044,N_24323);
or U28989 (N_28989,N_21846,N_24993);
xor U28990 (N_28990,N_20010,N_20177);
or U28991 (N_28991,N_22584,N_24072);
or U28992 (N_28992,N_21287,N_24714);
or U28993 (N_28993,N_22700,N_23542);
or U28994 (N_28994,N_21974,N_20334);
or U28995 (N_28995,N_21396,N_21502);
or U28996 (N_28996,N_21441,N_24838);
nor U28997 (N_28997,N_20615,N_20668);
or U28998 (N_28998,N_20601,N_23799);
nand U28999 (N_28999,N_20717,N_23085);
or U29000 (N_29000,N_24119,N_23789);
nand U29001 (N_29001,N_21253,N_24177);
xnor U29002 (N_29002,N_20414,N_20387);
nand U29003 (N_29003,N_20592,N_20265);
or U29004 (N_29004,N_23686,N_22795);
and U29005 (N_29005,N_23927,N_22855);
nor U29006 (N_29006,N_20337,N_22532);
nand U29007 (N_29007,N_23840,N_20226);
and U29008 (N_29008,N_22661,N_21733);
and U29009 (N_29009,N_20173,N_21035);
xor U29010 (N_29010,N_24916,N_20434);
nor U29011 (N_29011,N_20128,N_22205);
or U29012 (N_29012,N_21429,N_21870);
xnor U29013 (N_29013,N_22111,N_20638);
nor U29014 (N_29014,N_23166,N_24892);
nand U29015 (N_29015,N_21153,N_20361);
or U29016 (N_29016,N_23240,N_22463);
xor U29017 (N_29017,N_20372,N_21342);
nand U29018 (N_29018,N_23805,N_21099);
and U29019 (N_29019,N_24907,N_20458);
or U29020 (N_29020,N_21953,N_22865);
and U29021 (N_29021,N_21059,N_20597);
nand U29022 (N_29022,N_24280,N_20958);
or U29023 (N_29023,N_23988,N_20363);
nand U29024 (N_29024,N_24911,N_20938);
nor U29025 (N_29025,N_23030,N_24372);
nor U29026 (N_29026,N_20911,N_22797);
nand U29027 (N_29027,N_24073,N_22232);
or U29028 (N_29028,N_24763,N_22859);
and U29029 (N_29029,N_24743,N_20395);
nand U29030 (N_29030,N_20135,N_22278);
or U29031 (N_29031,N_21672,N_24427);
and U29032 (N_29032,N_24253,N_21284);
and U29033 (N_29033,N_23276,N_24331);
or U29034 (N_29034,N_21489,N_21093);
or U29035 (N_29035,N_24675,N_23318);
xor U29036 (N_29036,N_22261,N_24265);
nand U29037 (N_29037,N_23476,N_21077);
nor U29038 (N_29038,N_21469,N_21504);
and U29039 (N_29039,N_22704,N_24141);
or U29040 (N_29040,N_21454,N_21228);
nand U29041 (N_29041,N_23220,N_21136);
or U29042 (N_29042,N_24568,N_23585);
nand U29043 (N_29043,N_20048,N_23175);
and U29044 (N_29044,N_22817,N_23626);
xor U29045 (N_29045,N_23325,N_21878);
nor U29046 (N_29046,N_21508,N_24898);
xor U29047 (N_29047,N_23022,N_21919);
or U29048 (N_29048,N_24233,N_20446);
nand U29049 (N_29049,N_22876,N_22933);
nand U29050 (N_29050,N_21852,N_22608);
nor U29051 (N_29051,N_24730,N_22642);
nand U29052 (N_29052,N_23306,N_24600);
and U29053 (N_29053,N_20903,N_22932);
nand U29054 (N_29054,N_20651,N_22023);
nor U29055 (N_29055,N_22364,N_23048);
nand U29056 (N_29056,N_22511,N_21417);
nand U29057 (N_29057,N_20189,N_20385);
and U29058 (N_29058,N_24898,N_22021);
xor U29059 (N_29059,N_24077,N_22148);
and U29060 (N_29060,N_20255,N_22427);
nor U29061 (N_29061,N_23023,N_23270);
and U29062 (N_29062,N_22925,N_24837);
nand U29063 (N_29063,N_23604,N_24757);
xnor U29064 (N_29064,N_21050,N_24140);
nand U29065 (N_29065,N_21635,N_20305);
nor U29066 (N_29066,N_23094,N_24933);
nor U29067 (N_29067,N_24755,N_20726);
and U29068 (N_29068,N_24334,N_23861);
xor U29069 (N_29069,N_23675,N_21312);
nand U29070 (N_29070,N_20595,N_24027);
and U29071 (N_29071,N_23081,N_23389);
or U29072 (N_29072,N_20771,N_20584);
xor U29073 (N_29073,N_21726,N_24187);
nand U29074 (N_29074,N_20487,N_24392);
or U29075 (N_29075,N_24931,N_24104);
nor U29076 (N_29076,N_20400,N_23602);
nand U29077 (N_29077,N_24342,N_23063);
nand U29078 (N_29078,N_24826,N_23565);
nor U29079 (N_29079,N_22310,N_22916);
or U29080 (N_29080,N_24393,N_21241);
nand U29081 (N_29081,N_24165,N_20795);
or U29082 (N_29082,N_21819,N_20083);
or U29083 (N_29083,N_20100,N_20662);
and U29084 (N_29084,N_24905,N_22682);
or U29085 (N_29085,N_21476,N_20965);
or U29086 (N_29086,N_22603,N_23888);
and U29087 (N_29087,N_22903,N_22131);
or U29088 (N_29088,N_22496,N_22700);
or U29089 (N_29089,N_22882,N_22966);
or U29090 (N_29090,N_23578,N_22481);
nor U29091 (N_29091,N_24814,N_20408);
nand U29092 (N_29092,N_24239,N_24815);
or U29093 (N_29093,N_21711,N_21029);
nor U29094 (N_29094,N_21778,N_23958);
xnor U29095 (N_29095,N_23324,N_20804);
nand U29096 (N_29096,N_24556,N_20135);
or U29097 (N_29097,N_22452,N_21064);
nor U29098 (N_29098,N_20425,N_21798);
and U29099 (N_29099,N_22485,N_20145);
nand U29100 (N_29100,N_23680,N_23724);
nand U29101 (N_29101,N_22509,N_21388);
or U29102 (N_29102,N_24451,N_20443);
nand U29103 (N_29103,N_21965,N_20712);
and U29104 (N_29104,N_21064,N_22749);
nand U29105 (N_29105,N_23801,N_22730);
or U29106 (N_29106,N_22068,N_20250);
nor U29107 (N_29107,N_21931,N_20909);
and U29108 (N_29108,N_23950,N_23685);
or U29109 (N_29109,N_24633,N_22543);
nand U29110 (N_29110,N_23900,N_21942);
xor U29111 (N_29111,N_23414,N_22207);
or U29112 (N_29112,N_22738,N_23765);
or U29113 (N_29113,N_21210,N_23385);
nand U29114 (N_29114,N_20906,N_23427);
or U29115 (N_29115,N_22886,N_23456);
and U29116 (N_29116,N_21824,N_20578);
or U29117 (N_29117,N_23763,N_24572);
or U29118 (N_29118,N_22874,N_20244);
and U29119 (N_29119,N_23593,N_24348);
and U29120 (N_29120,N_21291,N_22590);
nor U29121 (N_29121,N_24527,N_23643);
and U29122 (N_29122,N_24972,N_23846);
or U29123 (N_29123,N_23414,N_21711);
and U29124 (N_29124,N_24735,N_22663);
nand U29125 (N_29125,N_22510,N_20430);
nand U29126 (N_29126,N_20011,N_22384);
xnor U29127 (N_29127,N_20897,N_20805);
and U29128 (N_29128,N_21772,N_22276);
nand U29129 (N_29129,N_23081,N_22092);
nand U29130 (N_29130,N_24587,N_24192);
and U29131 (N_29131,N_23271,N_20924);
and U29132 (N_29132,N_22135,N_21468);
nor U29133 (N_29133,N_23611,N_24837);
nor U29134 (N_29134,N_23866,N_21847);
and U29135 (N_29135,N_24393,N_22699);
nand U29136 (N_29136,N_21873,N_22027);
nand U29137 (N_29137,N_23557,N_21948);
or U29138 (N_29138,N_23680,N_20739);
nand U29139 (N_29139,N_21264,N_23532);
and U29140 (N_29140,N_24337,N_24201);
nor U29141 (N_29141,N_20456,N_24076);
or U29142 (N_29142,N_23502,N_23630);
and U29143 (N_29143,N_23208,N_20000);
or U29144 (N_29144,N_21228,N_21108);
and U29145 (N_29145,N_21118,N_22130);
or U29146 (N_29146,N_22272,N_21324);
or U29147 (N_29147,N_23396,N_21542);
nand U29148 (N_29148,N_20494,N_21156);
nand U29149 (N_29149,N_23724,N_22756);
xor U29150 (N_29150,N_24633,N_22420);
nand U29151 (N_29151,N_24110,N_20613);
and U29152 (N_29152,N_24497,N_20142);
xor U29153 (N_29153,N_24343,N_21088);
nand U29154 (N_29154,N_23421,N_22198);
nand U29155 (N_29155,N_22516,N_24785);
xnor U29156 (N_29156,N_22367,N_20147);
and U29157 (N_29157,N_24779,N_23409);
xor U29158 (N_29158,N_20027,N_23116);
or U29159 (N_29159,N_20550,N_20768);
nor U29160 (N_29160,N_22635,N_21293);
xnor U29161 (N_29161,N_21865,N_23007);
or U29162 (N_29162,N_24048,N_22479);
or U29163 (N_29163,N_23658,N_22058);
nor U29164 (N_29164,N_24099,N_20903);
or U29165 (N_29165,N_22121,N_21227);
and U29166 (N_29166,N_20486,N_20523);
and U29167 (N_29167,N_21655,N_22058);
or U29168 (N_29168,N_23079,N_23046);
or U29169 (N_29169,N_21347,N_23310);
nand U29170 (N_29170,N_22285,N_22217);
and U29171 (N_29171,N_21838,N_24508);
and U29172 (N_29172,N_20741,N_21129);
xnor U29173 (N_29173,N_20956,N_24310);
and U29174 (N_29174,N_20483,N_24370);
or U29175 (N_29175,N_23665,N_23441);
or U29176 (N_29176,N_21151,N_24534);
and U29177 (N_29177,N_20725,N_23520);
xor U29178 (N_29178,N_23838,N_21267);
nand U29179 (N_29179,N_22436,N_22869);
nand U29180 (N_29180,N_22357,N_22816);
nor U29181 (N_29181,N_23034,N_24213);
and U29182 (N_29182,N_21875,N_24242);
and U29183 (N_29183,N_23797,N_20354);
or U29184 (N_29184,N_21246,N_20301);
nor U29185 (N_29185,N_20399,N_23430);
or U29186 (N_29186,N_20807,N_20478);
nand U29187 (N_29187,N_23387,N_23593);
nand U29188 (N_29188,N_21609,N_21745);
nor U29189 (N_29189,N_24165,N_21990);
nand U29190 (N_29190,N_24313,N_24608);
xnor U29191 (N_29191,N_23696,N_22471);
xnor U29192 (N_29192,N_20029,N_24703);
and U29193 (N_29193,N_23276,N_24660);
and U29194 (N_29194,N_21506,N_22957);
xor U29195 (N_29195,N_23551,N_22677);
nor U29196 (N_29196,N_23103,N_23054);
or U29197 (N_29197,N_20768,N_21087);
or U29198 (N_29198,N_24197,N_20167);
nor U29199 (N_29199,N_22573,N_22337);
nor U29200 (N_29200,N_23754,N_24900);
or U29201 (N_29201,N_20147,N_22714);
or U29202 (N_29202,N_24059,N_21158);
and U29203 (N_29203,N_21925,N_24327);
and U29204 (N_29204,N_21691,N_22301);
nor U29205 (N_29205,N_20762,N_21877);
or U29206 (N_29206,N_22818,N_23811);
nor U29207 (N_29207,N_21653,N_23470);
or U29208 (N_29208,N_24083,N_24200);
and U29209 (N_29209,N_22323,N_20490);
or U29210 (N_29210,N_21700,N_22533);
xnor U29211 (N_29211,N_24818,N_20335);
nand U29212 (N_29212,N_20438,N_22739);
nand U29213 (N_29213,N_22285,N_22121);
nand U29214 (N_29214,N_21230,N_22002);
nand U29215 (N_29215,N_22774,N_21080);
and U29216 (N_29216,N_24446,N_20369);
or U29217 (N_29217,N_24233,N_21779);
or U29218 (N_29218,N_23061,N_20466);
nor U29219 (N_29219,N_23090,N_20259);
nand U29220 (N_29220,N_20184,N_20831);
or U29221 (N_29221,N_24651,N_24881);
nor U29222 (N_29222,N_20986,N_21710);
nor U29223 (N_29223,N_23281,N_20148);
and U29224 (N_29224,N_20537,N_21904);
nor U29225 (N_29225,N_21606,N_22286);
nor U29226 (N_29226,N_23919,N_22937);
nand U29227 (N_29227,N_23664,N_21706);
nand U29228 (N_29228,N_23160,N_22315);
or U29229 (N_29229,N_21947,N_22531);
nand U29230 (N_29230,N_24157,N_22435);
nor U29231 (N_29231,N_22899,N_20299);
and U29232 (N_29232,N_21647,N_22451);
nand U29233 (N_29233,N_24818,N_22328);
nor U29234 (N_29234,N_23085,N_21892);
nor U29235 (N_29235,N_24330,N_23790);
nor U29236 (N_29236,N_21832,N_22318);
nor U29237 (N_29237,N_22763,N_23767);
and U29238 (N_29238,N_23202,N_22348);
or U29239 (N_29239,N_22048,N_24449);
nand U29240 (N_29240,N_21874,N_23217);
nor U29241 (N_29241,N_23283,N_21686);
or U29242 (N_29242,N_21184,N_20722);
and U29243 (N_29243,N_20865,N_21067);
nand U29244 (N_29244,N_22139,N_22525);
nand U29245 (N_29245,N_23934,N_21998);
nand U29246 (N_29246,N_23705,N_23177);
nor U29247 (N_29247,N_21506,N_22719);
nand U29248 (N_29248,N_23721,N_24328);
and U29249 (N_29249,N_21962,N_24062);
nand U29250 (N_29250,N_21057,N_20780);
or U29251 (N_29251,N_24773,N_23044);
or U29252 (N_29252,N_21813,N_22720);
nor U29253 (N_29253,N_23768,N_22687);
or U29254 (N_29254,N_24026,N_24326);
xor U29255 (N_29255,N_24029,N_23041);
nor U29256 (N_29256,N_24035,N_20015);
nand U29257 (N_29257,N_24683,N_20582);
nor U29258 (N_29258,N_22770,N_23430);
xor U29259 (N_29259,N_20502,N_24271);
nor U29260 (N_29260,N_22189,N_21210);
and U29261 (N_29261,N_21819,N_22854);
or U29262 (N_29262,N_22715,N_20588);
or U29263 (N_29263,N_22490,N_24017);
or U29264 (N_29264,N_20488,N_21344);
and U29265 (N_29265,N_24148,N_22248);
or U29266 (N_29266,N_24023,N_20980);
nand U29267 (N_29267,N_20122,N_21208);
nor U29268 (N_29268,N_20881,N_22170);
nand U29269 (N_29269,N_24763,N_22949);
or U29270 (N_29270,N_22758,N_23991);
nor U29271 (N_29271,N_23641,N_20441);
and U29272 (N_29272,N_21353,N_20779);
nand U29273 (N_29273,N_24136,N_20111);
and U29274 (N_29274,N_20583,N_22592);
or U29275 (N_29275,N_20625,N_23894);
and U29276 (N_29276,N_23288,N_24227);
nor U29277 (N_29277,N_21907,N_23192);
nand U29278 (N_29278,N_20129,N_20475);
nor U29279 (N_29279,N_22572,N_21976);
nor U29280 (N_29280,N_20312,N_23875);
nand U29281 (N_29281,N_20425,N_20865);
and U29282 (N_29282,N_23204,N_23562);
nand U29283 (N_29283,N_22652,N_20785);
xnor U29284 (N_29284,N_20216,N_24873);
nand U29285 (N_29285,N_24530,N_21383);
or U29286 (N_29286,N_22854,N_21885);
and U29287 (N_29287,N_24534,N_20698);
and U29288 (N_29288,N_20160,N_22657);
nor U29289 (N_29289,N_21903,N_24356);
nand U29290 (N_29290,N_21357,N_24816);
nor U29291 (N_29291,N_22783,N_22719);
or U29292 (N_29292,N_24856,N_24898);
or U29293 (N_29293,N_24206,N_20590);
or U29294 (N_29294,N_23706,N_20861);
or U29295 (N_29295,N_23829,N_24132);
or U29296 (N_29296,N_24412,N_24869);
nand U29297 (N_29297,N_24302,N_21079);
nor U29298 (N_29298,N_21324,N_21650);
nand U29299 (N_29299,N_21430,N_23058);
nor U29300 (N_29300,N_22745,N_20144);
nand U29301 (N_29301,N_24116,N_21740);
nor U29302 (N_29302,N_21341,N_22180);
nor U29303 (N_29303,N_24899,N_24315);
nand U29304 (N_29304,N_23149,N_21516);
and U29305 (N_29305,N_24325,N_22223);
nand U29306 (N_29306,N_23556,N_20709);
and U29307 (N_29307,N_22740,N_22148);
nor U29308 (N_29308,N_20995,N_23258);
nor U29309 (N_29309,N_22565,N_20198);
nor U29310 (N_29310,N_21320,N_21609);
and U29311 (N_29311,N_22573,N_21063);
nor U29312 (N_29312,N_22060,N_22249);
nand U29313 (N_29313,N_24882,N_20328);
and U29314 (N_29314,N_24811,N_24500);
nand U29315 (N_29315,N_23442,N_23291);
or U29316 (N_29316,N_21284,N_22013);
xor U29317 (N_29317,N_24150,N_23517);
nand U29318 (N_29318,N_20197,N_22239);
nor U29319 (N_29319,N_24040,N_21374);
or U29320 (N_29320,N_24202,N_22774);
nand U29321 (N_29321,N_21670,N_21496);
and U29322 (N_29322,N_24068,N_20904);
nor U29323 (N_29323,N_20261,N_22501);
nand U29324 (N_29324,N_22063,N_23603);
or U29325 (N_29325,N_21107,N_23961);
nor U29326 (N_29326,N_22649,N_24377);
and U29327 (N_29327,N_22978,N_20727);
nand U29328 (N_29328,N_21596,N_24583);
or U29329 (N_29329,N_23220,N_23947);
nor U29330 (N_29330,N_23723,N_24099);
nor U29331 (N_29331,N_20210,N_22928);
nor U29332 (N_29332,N_24704,N_23682);
nor U29333 (N_29333,N_24888,N_20509);
or U29334 (N_29334,N_22204,N_20485);
or U29335 (N_29335,N_24383,N_23909);
and U29336 (N_29336,N_21079,N_20850);
nand U29337 (N_29337,N_20216,N_22408);
and U29338 (N_29338,N_21217,N_22218);
xnor U29339 (N_29339,N_22780,N_21882);
xnor U29340 (N_29340,N_21353,N_21270);
xnor U29341 (N_29341,N_21743,N_21157);
or U29342 (N_29342,N_23943,N_20220);
nor U29343 (N_29343,N_20765,N_23626);
nor U29344 (N_29344,N_20247,N_24822);
and U29345 (N_29345,N_20420,N_21586);
xnor U29346 (N_29346,N_20448,N_23843);
nor U29347 (N_29347,N_20920,N_20072);
xor U29348 (N_29348,N_21225,N_21893);
nand U29349 (N_29349,N_20159,N_22757);
nand U29350 (N_29350,N_20222,N_20871);
nand U29351 (N_29351,N_23539,N_24878);
or U29352 (N_29352,N_24123,N_21365);
nand U29353 (N_29353,N_20121,N_20171);
and U29354 (N_29354,N_24377,N_22169);
nand U29355 (N_29355,N_23199,N_21871);
nand U29356 (N_29356,N_20050,N_24116);
nand U29357 (N_29357,N_24666,N_24031);
or U29358 (N_29358,N_20035,N_22200);
and U29359 (N_29359,N_24518,N_24385);
nor U29360 (N_29360,N_24515,N_21883);
or U29361 (N_29361,N_22531,N_21533);
nand U29362 (N_29362,N_20926,N_23152);
and U29363 (N_29363,N_23483,N_21822);
nor U29364 (N_29364,N_22517,N_22843);
and U29365 (N_29365,N_24411,N_23333);
nand U29366 (N_29366,N_24197,N_20694);
nor U29367 (N_29367,N_20167,N_20562);
and U29368 (N_29368,N_20429,N_20065);
xor U29369 (N_29369,N_24131,N_20910);
nand U29370 (N_29370,N_24704,N_24074);
nand U29371 (N_29371,N_24704,N_21760);
nor U29372 (N_29372,N_24477,N_24832);
nand U29373 (N_29373,N_22882,N_23992);
nor U29374 (N_29374,N_22284,N_23523);
or U29375 (N_29375,N_20041,N_20774);
nand U29376 (N_29376,N_24220,N_21982);
nor U29377 (N_29377,N_22345,N_24163);
and U29378 (N_29378,N_22426,N_21058);
nor U29379 (N_29379,N_24349,N_24551);
nor U29380 (N_29380,N_21861,N_21325);
nand U29381 (N_29381,N_20174,N_24836);
nand U29382 (N_29382,N_23842,N_20302);
or U29383 (N_29383,N_20940,N_22936);
or U29384 (N_29384,N_23117,N_21043);
or U29385 (N_29385,N_21093,N_24169);
nand U29386 (N_29386,N_23817,N_24017);
nand U29387 (N_29387,N_23861,N_22384);
nor U29388 (N_29388,N_24114,N_22004);
or U29389 (N_29389,N_20515,N_24473);
nand U29390 (N_29390,N_23907,N_23234);
and U29391 (N_29391,N_22294,N_24059);
nand U29392 (N_29392,N_24290,N_22458);
or U29393 (N_29393,N_23023,N_22569);
or U29394 (N_29394,N_23902,N_20745);
nor U29395 (N_29395,N_23207,N_23744);
nand U29396 (N_29396,N_21008,N_21679);
nor U29397 (N_29397,N_23069,N_21604);
xor U29398 (N_29398,N_21625,N_20693);
nor U29399 (N_29399,N_21750,N_23492);
nand U29400 (N_29400,N_24572,N_24332);
nor U29401 (N_29401,N_23829,N_23924);
or U29402 (N_29402,N_22513,N_21079);
and U29403 (N_29403,N_22894,N_24298);
nand U29404 (N_29404,N_22660,N_20336);
or U29405 (N_29405,N_22755,N_24218);
nor U29406 (N_29406,N_23038,N_20839);
nand U29407 (N_29407,N_23594,N_21483);
nand U29408 (N_29408,N_24557,N_23834);
nor U29409 (N_29409,N_20410,N_23798);
xnor U29410 (N_29410,N_22809,N_21171);
nand U29411 (N_29411,N_22652,N_20897);
and U29412 (N_29412,N_22587,N_20684);
and U29413 (N_29413,N_22758,N_22595);
or U29414 (N_29414,N_21960,N_23537);
and U29415 (N_29415,N_23499,N_22749);
and U29416 (N_29416,N_23403,N_20054);
nor U29417 (N_29417,N_22813,N_21890);
nand U29418 (N_29418,N_24550,N_22495);
or U29419 (N_29419,N_20196,N_22747);
nand U29420 (N_29420,N_23063,N_22363);
nor U29421 (N_29421,N_21716,N_24378);
nand U29422 (N_29422,N_24475,N_22649);
or U29423 (N_29423,N_20570,N_20450);
or U29424 (N_29424,N_21958,N_21518);
nor U29425 (N_29425,N_22594,N_20560);
and U29426 (N_29426,N_24998,N_20937);
nor U29427 (N_29427,N_23523,N_22590);
or U29428 (N_29428,N_23361,N_20914);
and U29429 (N_29429,N_20493,N_24271);
xnor U29430 (N_29430,N_21596,N_24742);
and U29431 (N_29431,N_20021,N_21733);
and U29432 (N_29432,N_23848,N_23498);
nor U29433 (N_29433,N_23721,N_20737);
and U29434 (N_29434,N_24017,N_23035);
or U29435 (N_29435,N_21468,N_23080);
nor U29436 (N_29436,N_20561,N_22216);
nor U29437 (N_29437,N_24154,N_21029);
nor U29438 (N_29438,N_21460,N_22853);
nor U29439 (N_29439,N_22540,N_21823);
and U29440 (N_29440,N_22755,N_22624);
nor U29441 (N_29441,N_22938,N_23211);
nor U29442 (N_29442,N_21746,N_20964);
or U29443 (N_29443,N_21068,N_21427);
and U29444 (N_29444,N_21425,N_23421);
and U29445 (N_29445,N_21714,N_23860);
nor U29446 (N_29446,N_23800,N_21512);
nor U29447 (N_29447,N_21850,N_21561);
and U29448 (N_29448,N_24591,N_24629);
and U29449 (N_29449,N_21037,N_22447);
nor U29450 (N_29450,N_21382,N_24844);
xnor U29451 (N_29451,N_22919,N_21212);
nand U29452 (N_29452,N_22100,N_21992);
nor U29453 (N_29453,N_22792,N_24299);
nor U29454 (N_29454,N_20271,N_23555);
and U29455 (N_29455,N_24108,N_20922);
and U29456 (N_29456,N_24558,N_21927);
xor U29457 (N_29457,N_21156,N_21711);
nor U29458 (N_29458,N_21704,N_21613);
or U29459 (N_29459,N_22744,N_24990);
or U29460 (N_29460,N_20321,N_21152);
and U29461 (N_29461,N_24401,N_24755);
or U29462 (N_29462,N_24327,N_21641);
nand U29463 (N_29463,N_24219,N_23801);
and U29464 (N_29464,N_21321,N_20794);
and U29465 (N_29465,N_21006,N_20884);
nand U29466 (N_29466,N_24315,N_23593);
and U29467 (N_29467,N_22858,N_24173);
xor U29468 (N_29468,N_20644,N_22801);
or U29469 (N_29469,N_22389,N_22068);
and U29470 (N_29470,N_20258,N_22333);
nand U29471 (N_29471,N_24832,N_22389);
xnor U29472 (N_29472,N_20988,N_23158);
nor U29473 (N_29473,N_20010,N_24252);
and U29474 (N_29474,N_24899,N_20479);
nor U29475 (N_29475,N_21224,N_21758);
or U29476 (N_29476,N_21514,N_21521);
xnor U29477 (N_29477,N_21108,N_21936);
and U29478 (N_29478,N_22321,N_21849);
or U29479 (N_29479,N_22728,N_22152);
nand U29480 (N_29480,N_21236,N_24069);
nand U29481 (N_29481,N_22479,N_24838);
nor U29482 (N_29482,N_23879,N_20684);
xnor U29483 (N_29483,N_24191,N_20621);
nand U29484 (N_29484,N_23012,N_20603);
nor U29485 (N_29485,N_24022,N_20769);
nand U29486 (N_29486,N_24882,N_22787);
or U29487 (N_29487,N_20957,N_22513);
or U29488 (N_29488,N_24287,N_20463);
or U29489 (N_29489,N_21335,N_20708);
or U29490 (N_29490,N_23735,N_20939);
nand U29491 (N_29491,N_24696,N_22562);
nor U29492 (N_29492,N_22909,N_22547);
nor U29493 (N_29493,N_22142,N_24079);
nand U29494 (N_29494,N_22015,N_23846);
and U29495 (N_29495,N_21425,N_21314);
nor U29496 (N_29496,N_24323,N_21006);
or U29497 (N_29497,N_22401,N_20611);
or U29498 (N_29498,N_22761,N_23538);
nand U29499 (N_29499,N_20177,N_22407);
nand U29500 (N_29500,N_21533,N_24954);
and U29501 (N_29501,N_23055,N_20655);
or U29502 (N_29502,N_21353,N_20293);
xnor U29503 (N_29503,N_24605,N_21522);
xor U29504 (N_29504,N_21916,N_20012);
nor U29505 (N_29505,N_20661,N_22376);
or U29506 (N_29506,N_21567,N_23072);
nand U29507 (N_29507,N_23004,N_20738);
and U29508 (N_29508,N_20649,N_24296);
nor U29509 (N_29509,N_23120,N_20922);
nor U29510 (N_29510,N_23521,N_23608);
and U29511 (N_29511,N_24083,N_20089);
or U29512 (N_29512,N_23514,N_24068);
nand U29513 (N_29513,N_21236,N_21609);
nor U29514 (N_29514,N_22799,N_23563);
xor U29515 (N_29515,N_22320,N_20751);
nor U29516 (N_29516,N_20616,N_21678);
nand U29517 (N_29517,N_23505,N_23695);
xnor U29518 (N_29518,N_24937,N_22249);
xnor U29519 (N_29519,N_23169,N_22103);
or U29520 (N_29520,N_21098,N_23922);
nor U29521 (N_29521,N_24448,N_24787);
and U29522 (N_29522,N_23543,N_20909);
nor U29523 (N_29523,N_20357,N_22362);
nand U29524 (N_29524,N_21970,N_23236);
nor U29525 (N_29525,N_24506,N_21042);
nor U29526 (N_29526,N_24801,N_21916);
and U29527 (N_29527,N_24680,N_20603);
and U29528 (N_29528,N_23815,N_23995);
nor U29529 (N_29529,N_22775,N_24412);
or U29530 (N_29530,N_21633,N_21771);
nor U29531 (N_29531,N_24463,N_24687);
and U29532 (N_29532,N_23731,N_23790);
nor U29533 (N_29533,N_23012,N_22732);
nand U29534 (N_29534,N_23924,N_23667);
and U29535 (N_29535,N_23977,N_22920);
nor U29536 (N_29536,N_23320,N_23569);
and U29537 (N_29537,N_22374,N_22026);
or U29538 (N_29538,N_20089,N_22529);
and U29539 (N_29539,N_24117,N_24166);
and U29540 (N_29540,N_22710,N_23647);
nand U29541 (N_29541,N_22953,N_20005);
or U29542 (N_29542,N_20481,N_24400);
nand U29543 (N_29543,N_20962,N_21576);
or U29544 (N_29544,N_20242,N_20243);
and U29545 (N_29545,N_23286,N_23597);
and U29546 (N_29546,N_20574,N_20232);
or U29547 (N_29547,N_22896,N_22770);
nand U29548 (N_29548,N_20771,N_21253);
nor U29549 (N_29549,N_22026,N_23484);
and U29550 (N_29550,N_24778,N_23382);
and U29551 (N_29551,N_23455,N_24558);
or U29552 (N_29552,N_22954,N_22994);
and U29553 (N_29553,N_22021,N_22469);
or U29554 (N_29554,N_20198,N_21904);
or U29555 (N_29555,N_20848,N_23580);
nor U29556 (N_29556,N_23498,N_23967);
xnor U29557 (N_29557,N_21824,N_21901);
xnor U29558 (N_29558,N_21073,N_23326);
or U29559 (N_29559,N_24932,N_20258);
or U29560 (N_29560,N_21127,N_22918);
and U29561 (N_29561,N_20259,N_20845);
nor U29562 (N_29562,N_24818,N_22679);
or U29563 (N_29563,N_22349,N_22985);
or U29564 (N_29564,N_22731,N_21535);
nand U29565 (N_29565,N_21958,N_21080);
nor U29566 (N_29566,N_24109,N_20945);
nand U29567 (N_29567,N_21853,N_20259);
or U29568 (N_29568,N_22559,N_24318);
nor U29569 (N_29569,N_22369,N_20900);
and U29570 (N_29570,N_22731,N_21059);
nand U29571 (N_29571,N_22983,N_22211);
and U29572 (N_29572,N_23295,N_22341);
nand U29573 (N_29573,N_24883,N_23819);
nor U29574 (N_29574,N_22008,N_24742);
or U29575 (N_29575,N_24078,N_20154);
nand U29576 (N_29576,N_23293,N_22101);
and U29577 (N_29577,N_20884,N_20010);
nand U29578 (N_29578,N_21033,N_22642);
nand U29579 (N_29579,N_23464,N_24714);
or U29580 (N_29580,N_20309,N_23951);
nor U29581 (N_29581,N_20782,N_24783);
or U29582 (N_29582,N_23879,N_21436);
nand U29583 (N_29583,N_22182,N_20459);
and U29584 (N_29584,N_21998,N_21110);
or U29585 (N_29585,N_23506,N_23589);
and U29586 (N_29586,N_20567,N_24660);
or U29587 (N_29587,N_24855,N_20719);
nand U29588 (N_29588,N_23081,N_24370);
nand U29589 (N_29589,N_22603,N_23916);
nor U29590 (N_29590,N_24137,N_23012);
nand U29591 (N_29591,N_21983,N_23516);
and U29592 (N_29592,N_21231,N_23587);
or U29593 (N_29593,N_24631,N_24510);
and U29594 (N_29594,N_21400,N_23378);
nand U29595 (N_29595,N_24548,N_21766);
nand U29596 (N_29596,N_20642,N_20243);
nand U29597 (N_29597,N_21447,N_24693);
nand U29598 (N_29598,N_23705,N_24692);
or U29599 (N_29599,N_23863,N_20614);
nor U29600 (N_29600,N_23501,N_21447);
and U29601 (N_29601,N_22416,N_22707);
nand U29602 (N_29602,N_24716,N_20382);
and U29603 (N_29603,N_22999,N_23513);
or U29604 (N_29604,N_23687,N_23483);
xnor U29605 (N_29605,N_22418,N_23072);
and U29606 (N_29606,N_20517,N_24680);
xor U29607 (N_29607,N_20804,N_20934);
or U29608 (N_29608,N_22945,N_20264);
nand U29609 (N_29609,N_23294,N_21311);
and U29610 (N_29610,N_21772,N_22731);
or U29611 (N_29611,N_22690,N_20571);
or U29612 (N_29612,N_21883,N_20766);
and U29613 (N_29613,N_24832,N_21625);
xnor U29614 (N_29614,N_24914,N_22821);
or U29615 (N_29615,N_22905,N_23409);
or U29616 (N_29616,N_22582,N_21436);
nor U29617 (N_29617,N_24351,N_22141);
or U29618 (N_29618,N_23217,N_22728);
and U29619 (N_29619,N_22484,N_23094);
and U29620 (N_29620,N_21829,N_21938);
or U29621 (N_29621,N_21382,N_20020);
nor U29622 (N_29622,N_21446,N_23028);
nor U29623 (N_29623,N_20193,N_23655);
or U29624 (N_29624,N_21993,N_22441);
nand U29625 (N_29625,N_21940,N_23987);
nand U29626 (N_29626,N_20638,N_22913);
nor U29627 (N_29627,N_20569,N_22984);
and U29628 (N_29628,N_22130,N_22102);
nor U29629 (N_29629,N_21018,N_24612);
or U29630 (N_29630,N_23580,N_20040);
or U29631 (N_29631,N_21961,N_23202);
nand U29632 (N_29632,N_20437,N_23922);
and U29633 (N_29633,N_20204,N_24095);
and U29634 (N_29634,N_23431,N_20022);
nand U29635 (N_29635,N_21195,N_24694);
xnor U29636 (N_29636,N_20005,N_21350);
or U29637 (N_29637,N_24972,N_23821);
or U29638 (N_29638,N_24996,N_22325);
nor U29639 (N_29639,N_20629,N_24137);
nand U29640 (N_29640,N_21551,N_21888);
nor U29641 (N_29641,N_22357,N_21821);
and U29642 (N_29642,N_20429,N_23611);
and U29643 (N_29643,N_22096,N_20564);
nand U29644 (N_29644,N_21607,N_20756);
nor U29645 (N_29645,N_22114,N_20966);
nor U29646 (N_29646,N_24728,N_24863);
xor U29647 (N_29647,N_23887,N_21338);
and U29648 (N_29648,N_24940,N_24531);
or U29649 (N_29649,N_22979,N_22263);
nor U29650 (N_29650,N_21819,N_24438);
nand U29651 (N_29651,N_24425,N_22788);
nand U29652 (N_29652,N_22401,N_22613);
nor U29653 (N_29653,N_20336,N_24372);
and U29654 (N_29654,N_22706,N_24818);
or U29655 (N_29655,N_24668,N_23135);
or U29656 (N_29656,N_24532,N_23758);
and U29657 (N_29657,N_21891,N_21054);
xnor U29658 (N_29658,N_21577,N_21090);
and U29659 (N_29659,N_20950,N_21193);
xnor U29660 (N_29660,N_24458,N_23751);
and U29661 (N_29661,N_21065,N_21351);
or U29662 (N_29662,N_23774,N_21475);
nor U29663 (N_29663,N_21901,N_20039);
or U29664 (N_29664,N_23988,N_24033);
xnor U29665 (N_29665,N_24272,N_24858);
nor U29666 (N_29666,N_23428,N_21391);
xnor U29667 (N_29667,N_20436,N_21012);
or U29668 (N_29668,N_20706,N_21766);
and U29669 (N_29669,N_24567,N_22505);
and U29670 (N_29670,N_20334,N_23467);
or U29671 (N_29671,N_21495,N_24153);
or U29672 (N_29672,N_21524,N_24640);
or U29673 (N_29673,N_22707,N_22383);
or U29674 (N_29674,N_20192,N_22463);
nand U29675 (N_29675,N_22894,N_22649);
nor U29676 (N_29676,N_24810,N_23144);
xnor U29677 (N_29677,N_23748,N_21286);
or U29678 (N_29678,N_20632,N_20432);
and U29679 (N_29679,N_23912,N_20854);
and U29680 (N_29680,N_23164,N_23287);
nor U29681 (N_29681,N_24739,N_24833);
or U29682 (N_29682,N_24976,N_24750);
or U29683 (N_29683,N_21183,N_24555);
nand U29684 (N_29684,N_21271,N_24373);
xor U29685 (N_29685,N_22894,N_20586);
xor U29686 (N_29686,N_22469,N_20201);
and U29687 (N_29687,N_22995,N_21599);
nor U29688 (N_29688,N_23165,N_20008);
or U29689 (N_29689,N_20371,N_23605);
and U29690 (N_29690,N_21975,N_23986);
or U29691 (N_29691,N_24142,N_21498);
nand U29692 (N_29692,N_21476,N_21207);
or U29693 (N_29693,N_24346,N_23363);
and U29694 (N_29694,N_23510,N_21888);
and U29695 (N_29695,N_20383,N_23438);
and U29696 (N_29696,N_24554,N_20955);
and U29697 (N_29697,N_22418,N_22752);
and U29698 (N_29698,N_21953,N_24860);
and U29699 (N_29699,N_24302,N_21118);
or U29700 (N_29700,N_22106,N_24532);
and U29701 (N_29701,N_23815,N_21925);
nor U29702 (N_29702,N_21275,N_22046);
and U29703 (N_29703,N_24944,N_21870);
nand U29704 (N_29704,N_24119,N_22978);
nor U29705 (N_29705,N_21398,N_21920);
nor U29706 (N_29706,N_22326,N_21808);
or U29707 (N_29707,N_21604,N_24473);
nand U29708 (N_29708,N_24736,N_21487);
nor U29709 (N_29709,N_20005,N_21998);
or U29710 (N_29710,N_21715,N_24687);
nand U29711 (N_29711,N_24011,N_23674);
or U29712 (N_29712,N_23898,N_24870);
or U29713 (N_29713,N_21847,N_21468);
or U29714 (N_29714,N_21757,N_20214);
nor U29715 (N_29715,N_22033,N_22044);
nor U29716 (N_29716,N_20069,N_22212);
and U29717 (N_29717,N_20551,N_22905);
and U29718 (N_29718,N_20846,N_24204);
nor U29719 (N_29719,N_23927,N_20826);
nor U29720 (N_29720,N_20928,N_22654);
or U29721 (N_29721,N_22575,N_24798);
xor U29722 (N_29722,N_21159,N_20468);
or U29723 (N_29723,N_23030,N_20619);
nand U29724 (N_29724,N_23431,N_20361);
and U29725 (N_29725,N_21706,N_23384);
or U29726 (N_29726,N_23226,N_23124);
and U29727 (N_29727,N_21840,N_23512);
or U29728 (N_29728,N_20412,N_24109);
and U29729 (N_29729,N_21908,N_24783);
nor U29730 (N_29730,N_21071,N_24238);
xor U29731 (N_29731,N_21049,N_23515);
nand U29732 (N_29732,N_21341,N_21855);
nor U29733 (N_29733,N_24673,N_22499);
and U29734 (N_29734,N_24975,N_22115);
nand U29735 (N_29735,N_24354,N_22563);
nor U29736 (N_29736,N_21342,N_20011);
nand U29737 (N_29737,N_21121,N_24067);
nand U29738 (N_29738,N_21891,N_21075);
or U29739 (N_29739,N_24853,N_20292);
or U29740 (N_29740,N_21962,N_21506);
xnor U29741 (N_29741,N_20814,N_23412);
xnor U29742 (N_29742,N_21788,N_22687);
and U29743 (N_29743,N_21196,N_24597);
and U29744 (N_29744,N_22530,N_21025);
nor U29745 (N_29745,N_23223,N_22460);
xnor U29746 (N_29746,N_23496,N_22247);
or U29747 (N_29747,N_24309,N_20646);
xor U29748 (N_29748,N_23512,N_22187);
nor U29749 (N_29749,N_20131,N_24323);
or U29750 (N_29750,N_22328,N_24404);
nor U29751 (N_29751,N_22499,N_22494);
nand U29752 (N_29752,N_20705,N_20748);
and U29753 (N_29753,N_24881,N_23893);
xor U29754 (N_29754,N_24222,N_22649);
nand U29755 (N_29755,N_21014,N_23052);
and U29756 (N_29756,N_21304,N_20420);
nand U29757 (N_29757,N_24218,N_21328);
nor U29758 (N_29758,N_23719,N_20511);
nand U29759 (N_29759,N_23045,N_20614);
nand U29760 (N_29760,N_24994,N_23230);
or U29761 (N_29761,N_23301,N_22508);
nor U29762 (N_29762,N_23068,N_21893);
nand U29763 (N_29763,N_23597,N_23186);
and U29764 (N_29764,N_22041,N_21686);
nor U29765 (N_29765,N_24806,N_23170);
and U29766 (N_29766,N_24499,N_20867);
or U29767 (N_29767,N_21587,N_20494);
nand U29768 (N_29768,N_24033,N_22523);
nand U29769 (N_29769,N_21123,N_23245);
or U29770 (N_29770,N_20981,N_24359);
and U29771 (N_29771,N_23410,N_21237);
or U29772 (N_29772,N_21236,N_20086);
nor U29773 (N_29773,N_23852,N_21052);
or U29774 (N_29774,N_24757,N_20443);
or U29775 (N_29775,N_21990,N_20063);
nor U29776 (N_29776,N_24936,N_24257);
nor U29777 (N_29777,N_23555,N_21236);
nand U29778 (N_29778,N_21385,N_22756);
xnor U29779 (N_29779,N_23702,N_22197);
and U29780 (N_29780,N_23919,N_22192);
or U29781 (N_29781,N_24880,N_23371);
xnor U29782 (N_29782,N_23052,N_24698);
nand U29783 (N_29783,N_22754,N_21441);
nor U29784 (N_29784,N_22604,N_22593);
and U29785 (N_29785,N_21506,N_23713);
nor U29786 (N_29786,N_22298,N_22083);
or U29787 (N_29787,N_24275,N_20655);
nand U29788 (N_29788,N_21141,N_20152);
and U29789 (N_29789,N_24920,N_21382);
nor U29790 (N_29790,N_23430,N_23006);
nor U29791 (N_29791,N_24202,N_21804);
and U29792 (N_29792,N_20027,N_20567);
nand U29793 (N_29793,N_23289,N_23814);
or U29794 (N_29794,N_24586,N_22807);
or U29795 (N_29795,N_22142,N_23683);
and U29796 (N_29796,N_22483,N_24875);
nor U29797 (N_29797,N_22657,N_24364);
nor U29798 (N_29798,N_23588,N_24793);
xor U29799 (N_29799,N_23905,N_24640);
and U29800 (N_29800,N_23030,N_20538);
nor U29801 (N_29801,N_22847,N_23125);
or U29802 (N_29802,N_21746,N_22560);
and U29803 (N_29803,N_22997,N_24892);
nor U29804 (N_29804,N_22604,N_20592);
nor U29805 (N_29805,N_20696,N_22129);
xnor U29806 (N_29806,N_22384,N_24372);
and U29807 (N_29807,N_20841,N_24244);
nor U29808 (N_29808,N_23685,N_23030);
nor U29809 (N_29809,N_24660,N_23889);
nor U29810 (N_29810,N_21538,N_24584);
or U29811 (N_29811,N_21392,N_21709);
and U29812 (N_29812,N_23876,N_21285);
nor U29813 (N_29813,N_24970,N_24967);
or U29814 (N_29814,N_23440,N_24851);
and U29815 (N_29815,N_22025,N_22570);
xor U29816 (N_29816,N_20547,N_20989);
and U29817 (N_29817,N_23895,N_22758);
or U29818 (N_29818,N_24422,N_24218);
and U29819 (N_29819,N_23077,N_24426);
and U29820 (N_29820,N_23991,N_20733);
and U29821 (N_29821,N_20801,N_24666);
nor U29822 (N_29822,N_22177,N_21759);
nor U29823 (N_29823,N_20729,N_23579);
nor U29824 (N_29824,N_21033,N_22059);
nand U29825 (N_29825,N_22890,N_21566);
nor U29826 (N_29826,N_22295,N_20576);
nor U29827 (N_29827,N_24383,N_20243);
nand U29828 (N_29828,N_20766,N_22987);
or U29829 (N_29829,N_22990,N_23221);
and U29830 (N_29830,N_22843,N_21858);
and U29831 (N_29831,N_23901,N_21026);
or U29832 (N_29832,N_20896,N_24369);
nand U29833 (N_29833,N_23212,N_20201);
xor U29834 (N_29834,N_21170,N_24638);
nand U29835 (N_29835,N_20366,N_24299);
xor U29836 (N_29836,N_20412,N_20949);
or U29837 (N_29837,N_23742,N_22441);
or U29838 (N_29838,N_21123,N_21710);
or U29839 (N_29839,N_20977,N_24634);
xnor U29840 (N_29840,N_21147,N_22791);
nand U29841 (N_29841,N_21159,N_20984);
and U29842 (N_29842,N_22783,N_23601);
and U29843 (N_29843,N_24772,N_23827);
or U29844 (N_29844,N_21167,N_22022);
nand U29845 (N_29845,N_20530,N_23901);
or U29846 (N_29846,N_21766,N_24988);
nor U29847 (N_29847,N_23844,N_24479);
nand U29848 (N_29848,N_20170,N_22129);
nand U29849 (N_29849,N_24089,N_24265);
nor U29850 (N_29850,N_23530,N_22570);
or U29851 (N_29851,N_23273,N_22860);
nor U29852 (N_29852,N_24692,N_20794);
nor U29853 (N_29853,N_20945,N_22008);
or U29854 (N_29854,N_21586,N_22835);
xor U29855 (N_29855,N_22780,N_24749);
and U29856 (N_29856,N_23954,N_23902);
xor U29857 (N_29857,N_21005,N_24727);
nor U29858 (N_29858,N_23196,N_21107);
and U29859 (N_29859,N_21674,N_21528);
or U29860 (N_29860,N_23249,N_23919);
nor U29861 (N_29861,N_22031,N_24276);
nand U29862 (N_29862,N_20138,N_21630);
or U29863 (N_29863,N_22888,N_20993);
nand U29864 (N_29864,N_20954,N_21381);
nor U29865 (N_29865,N_20325,N_20707);
nor U29866 (N_29866,N_24177,N_23117);
nor U29867 (N_29867,N_21902,N_24190);
xnor U29868 (N_29868,N_23872,N_24255);
or U29869 (N_29869,N_23342,N_23474);
or U29870 (N_29870,N_24189,N_24545);
nand U29871 (N_29871,N_24662,N_23103);
nor U29872 (N_29872,N_24753,N_20321);
and U29873 (N_29873,N_24333,N_24669);
xor U29874 (N_29874,N_20749,N_23393);
and U29875 (N_29875,N_23415,N_23068);
and U29876 (N_29876,N_21147,N_24232);
or U29877 (N_29877,N_24070,N_24799);
nor U29878 (N_29878,N_23138,N_21023);
nor U29879 (N_29879,N_23635,N_21739);
nor U29880 (N_29880,N_20823,N_22963);
and U29881 (N_29881,N_21414,N_20911);
nand U29882 (N_29882,N_24822,N_20245);
nor U29883 (N_29883,N_23518,N_20946);
nand U29884 (N_29884,N_22067,N_23553);
nor U29885 (N_29885,N_21330,N_22291);
and U29886 (N_29886,N_20555,N_23294);
nand U29887 (N_29887,N_23436,N_20968);
nand U29888 (N_29888,N_22141,N_23111);
nand U29889 (N_29889,N_21849,N_24320);
xnor U29890 (N_29890,N_20208,N_22112);
nand U29891 (N_29891,N_23905,N_24343);
nor U29892 (N_29892,N_24590,N_22818);
and U29893 (N_29893,N_20311,N_24474);
nand U29894 (N_29894,N_23279,N_23201);
and U29895 (N_29895,N_21561,N_23969);
nor U29896 (N_29896,N_21141,N_21573);
or U29897 (N_29897,N_24585,N_20576);
or U29898 (N_29898,N_21826,N_23937);
xnor U29899 (N_29899,N_23190,N_20729);
nor U29900 (N_29900,N_20940,N_20703);
nand U29901 (N_29901,N_22950,N_21754);
and U29902 (N_29902,N_24767,N_23064);
or U29903 (N_29903,N_24860,N_21283);
nor U29904 (N_29904,N_24839,N_22989);
or U29905 (N_29905,N_24931,N_22537);
xnor U29906 (N_29906,N_24989,N_24386);
nor U29907 (N_29907,N_22451,N_22843);
nand U29908 (N_29908,N_20050,N_22416);
nand U29909 (N_29909,N_22260,N_22580);
nor U29910 (N_29910,N_23826,N_21093);
nand U29911 (N_29911,N_23460,N_21089);
and U29912 (N_29912,N_20986,N_24419);
or U29913 (N_29913,N_23407,N_20260);
and U29914 (N_29914,N_24587,N_23210);
and U29915 (N_29915,N_23737,N_21165);
and U29916 (N_29916,N_22840,N_22742);
or U29917 (N_29917,N_23325,N_22681);
and U29918 (N_29918,N_21471,N_21473);
and U29919 (N_29919,N_23422,N_21024);
nor U29920 (N_29920,N_22761,N_23866);
nor U29921 (N_29921,N_24243,N_22348);
nand U29922 (N_29922,N_21646,N_21417);
and U29923 (N_29923,N_24863,N_22302);
nor U29924 (N_29924,N_24964,N_24877);
or U29925 (N_29925,N_24709,N_20039);
and U29926 (N_29926,N_22824,N_23913);
xor U29927 (N_29927,N_22109,N_23316);
nand U29928 (N_29928,N_21203,N_23164);
xnor U29929 (N_29929,N_22689,N_23933);
nor U29930 (N_29930,N_20799,N_23680);
or U29931 (N_29931,N_24719,N_24177);
or U29932 (N_29932,N_23017,N_24239);
nand U29933 (N_29933,N_23099,N_20200);
and U29934 (N_29934,N_24044,N_23202);
nand U29935 (N_29935,N_24157,N_21157);
nand U29936 (N_29936,N_23218,N_20651);
and U29937 (N_29937,N_22443,N_24113);
nand U29938 (N_29938,N_24838,N_21676);
and U29939 (N_29939,N_22649,N_23526);
nand U29940 (N_29940,N_21608,N_20852);
or U29941 (N_29941,N_22524,N_20756);
or U29942 (N_29942,N_21851,N_21876);
nor U29943 (N_29943,N_22628,N_22612);
nor U29944 (N_29944,N_23672,N_24084);
or U29945 (N_29945,N_23781,N_21537);
nand U29946 (N_29946,N_20583,N_23940);
nand U29947 (N_29947,N_24256,N_21762);
and U29948 (N_29948,N_24807,N_23728);
nand U29949 (N_29949,N_24442,N_20970);
nor U29950 (N_29950,N_23892,N_22768);
xnor U29951 (N_29951,N_21433,N_21134);
nand U29952 (N_29952,N_22911,N_22529);
and U29953 (N_29953,N_21016,N_22779);
and U29954 (N_29954,N_21615,N_21941);
and U29955 (N_29955,N_22491,N_22290);
and U29956 (N_29956,N_21856,N_23408);
nor U29957 (N_29957,N_22820,N_23514);
and U29958 (N_29958,N_21922,N_21001);
or U29959 (N_29959,N_20743,N_23501);
nand U29960 (N_29960,N_24758,N_22413);
or U29961 (N_29961,N_24526,N_24229);
and U29962 (N_29962,N_23868,N_24738);
or U29963 (N_29963,N_22309,N_23296);
xor U29964 (N_29964,N_20731,N_21026);
nor U29965 (N_29965,N_24753,N_24745);
nand U29966 (N_29966,N_20388,N_24445);
or U29967 (N_29967,N_21889,N_23888);
nor U29968 (N_29968,N_23573,N_21069);
nor U29969 (N_29969,N_23571,N_24541);
or U29970 (N_29970,N_23037,N_22241);
xnor U29971 (N_29971,N_22079,N_23056);
nand U29972 (N_29972,N_24578,N_21653);
or U29973 (N_29973,N_20166,N_22749);
and U29974 (N_29974,N_24739,N_24130);
nand U29975 (N_29975,N_23851,N_21564);
or U29976 (N_29976,N_22182,N_23110);
or U29977 (N_29977,N_20704,N_23650);
and U29978 (N_29978,N_24220,N_24011);
nor U29979 (N_29979,N_22611,N_23948);
and U29980 (N_29980,N_20464,N_23663);
and U29981 (N_29981,N_21736,N_20015);
or U29982 (N_29982,N_23129,N_21172);
and U29983 (N_29983,N_20628,N_20909);
nor U29984 (N_29984,N_22675,N_22536);
or U29985 (N_29985,N_20944,N_24208);
nand U29986 (N_29986,N_23101,N_23354);
nand U29987 (N_29987,N_23898,N_20517);
and U29988 (N_29988,N_23213,N_20377);
and U29989 (N_29989,N_24489,N_22353);
nand U29990 (N_29990,N_22200,N_21339);
xnor U29991 (N_29991,N_22507,N_23502);
and U29992 (N_29992,N_20159,N_20000);
nand U29993 (N_29993,N_23867,N_23868);
or U29994 (N_29994,N_22978,N_21652);
nor U29995 (N_29995,N_20213,N_23591);
nand U29996 (N_29996,N_20589,N_22262);
nor U29997 (N_29997,N_24193,N_21544);
and U29998 (N_29998,N_20505,N_20618);
nand U29999 (N_29999,N_20097,N_20137);
and UO_0 (O_0,N_29692,N_25076);
and UO_1 (O_1,N_27404,N_26327);
and UO_2 (O_2,N_29684,N_26511);
nand UO_3 (O_3,N_28920,N_28153);
or UO_4 (O_4,N_28757,N_29112);
nand UO_5 (O_5,N_29321,N_25461);
and UO_6 (O_6,N_26861,N_26828);
or UO_7 (O_7,N_26714,N_28255);
and UO_8 (O_8,N_29824,N_29432);
nand UO_9 (O_9,N_25985,N_25987);
nor UO_10 (O_10,N_25474,N_25115);
nor UO_11 (O_11,N_29600,N_28179);
nand UO_12 (O_12,N_26660,N_26846);
nand UO_13 (O_13,N_25731,N_27299);
nand UO_14 (O_14,N_26668,N_25056);
and UO_15 (O_15,N_27427,N_28527);
nand UO_16 (O_16,N_26029,N_26051);
xor UO_17 (O_17,N_25278,N_28744);
nor UO_18 (O_18,N_28949,N_26486);
or UO_19 (O_19,N_28495,N_27514);
or UO_20 (O_20,N_27483,N_28098);
or UO_21 (O_21,N_28806,N_27978);
xor UO_22 (O_22,N_29224,N_26210);
nand UO_23 (O_23,N_26705,N_29906);
nand UO_24 (O_24,N_27668,N_29821);
nand UO_25 (O_25,N_27154,N_28501);
or UO_26 (O_26,N_27629,N_25757);
or UO_27 (O_27,N_27466,N_27983);
nor UO_28 (O_28,N_25431,N_29033);
xor UO_29 (O_29,N_28418,N_28860);
nand UO_30 (O_30,N_27546,N_25108);
or UO_31 (O_31,N_27971,N_29789);
and UO_32 (O_32,N_27111,N_27521);
and UO_33 (O_33,N_29485,N_28552);
or UO_34 (O_34,N_26479,N_25833);
nor UO_35 (O_35,N_27790,N_27573);
or UO_36 (O_36,N_29628,N_27248);
xor UO_37 (O_37,N_26424,N_29062);
and UO_38 (O_38,N_25724,N_25682);
nor UO_39 (O_39,N_27630,N_28632);
and UO_40 (O_40,N_25589,N_25995);
or UO_41 (O_41,N_25222,N_29669);
or UO_42 (O_42,N_29254,N_27879);
nand UO_43 (O_43,N_25605,N_29881);
nor UO_44 (O_44,N_25824,N_28246);
or UO_45 (O_45,N_27115,N_25162);
nand UO_46 (O_46,N_25733,N_29987);
and UO_47 (O_47,N_28162,N_28155);
xor UO_48 (O_48,N_25096,N_26840);
nand UO_49 (O_49,N_26801,N_26058);
nand UO_50 (O_50,N_25260,N_25259);
xor UO_51 (O_51,N_26164,N_25692);
nand UO_52 (O_52,N_26226,N_25738);
xnor UO_53 (O_53,N_27650,N_29914);
nand UO_54 (O_54,N_25418,N_27187);
and UO_55 (O_55,N_26987,N_29848);
nand UO_56 (O_56,N_26155,N_27534);
or UO_57 (O_57,N_27543,N_25262);
nand UO_58 (O_58,N_28511,N_27662);
nand UO_59 (O_59,N_28139,N_27909);
xor UO_60 (O_60,N_25070,N_27163);
nor UO_61 (O_61,N_25591,N_29688);
nand UO_62 (O_62,N_25652,N_28621);
or UO_63 (O_63,N_25925,N_29615);
or UO_64 (O_64,N_25338,N_28054);
and UO_65 (O_65,N_27673,N_27600);
nor UO_66 (O_66,N_25402,N_27590);
and UO_67 (O_67,N_25101,N_26826);
or UO_68 (O_68,N_25311,N_28036);
and UO_69 (O_69,N_27785,N_25825);
nor UO_70 (O_70,N_25964,N_29280);
nor UO_71 (O_71,N_28203,N_25837);
or UO_72 (O_72,N_26024,N_26417);
nand UO_73 (O_73,N_28195,N_29621);
nand UO_74 (O_74,N_25419,N_26009);
nor UO_75 (O_75,N_27621,N_27347);
or UO_76 (O_76,N_28886,N_28277);
or UO_77 (O_77,N_25221,N_29999);
nor UO_78 (O_78,N_29098,N_29808);
or UO_79 (O_79,N_27409,N_25487);
xnor UO_80 (O_80,N_27179,N_29035);
nand UO_81 (O_81,N_29758,N_29643);
and UO_82 (O_82,N_28345,N_29685);
xnor UO_83 (O_83,N_27724,N_26475);
and UO_84 (O_84,N_27817,N_28285);
and UO_85 (O_85,N_26062,N_28116);
nor UO_86 (O_86,N_25919,N_26493);
and UO_87 (O_87,N_28346,N_26719);
nor UO_88 (O_88,N_28655,N_27087);
and UO_89 (O_89,N_25239,N_25483);
xor UO_90 (O_90,N_26474,N_28704);
nor UO_91 (O_91,N_29016,N_27456);
or UO_92 (O_92,N_25729,N_26923);
and UO_93 (O_93,N_25107,N_26735);
or UO_94 (O_94,N_26976,N_27820);
nor UO_95 (O_95,N_25683,N_28395);
nand UO_96 (O_96,N_26132,N_25462);
nor UO_97 (O_97,N_25271,N_25631);
nor UO_98 (O_98,N_27905,N_26144);
nor UO_99 (O_99,N_25238,N_28338);
and UO_100 (O_100,N_25810,N_26581);
nand UO_101 (O_101,N_28944,N_26563);
and UO_102 (O_102,N_26872,N_26508);
and UO_103 (O_103,N_27839,N_26884);
or UO_104 (O_104,N_26489,N_26100);
nand UO_105 (O_105,N_25867,N_28491);
nand UO_106 (O_106,N_25646,N_29198);
and UO_107 (O_107,N_26723,N_26797);
and UO_108 (O_108,N_26050,N_28076);
and UO_109 (O_109,N_27917,N_25913);
or UO_110 (O_110,N_28065,N_26152);
or UO_111 (O_111,N_29993,N_29962);
and UO_112 (O_112,N_25320,N_25484);
and UO_113 (O_113,N_28684,N_27602);
and UO_114 (O_114,N_28990,N_26224);
nand UO_115 (O_115,N_28851,N_25007);
and UO_116 (O_116,N_27858,N_29780);
xor UO_117 (O_117,N_26598,N_25923);
or UO_118 (O_118,N_27101,N_25686);
or UO_119 (O_119,N_28661,N_25614);
nor UO_120 (O_120,N_26843,N_26295);
nor UO_121 (O_121,N_29579,N_29181);
or UO_122 (O_122,N_25073,N_25520);
or UO_123 (O_123,N_27583,N_27616);
nand UO_124 (O_124,N_27828,N_28440);
nand UO_125 (O_125,N_27228,N_27618);
and UO_126 (O_126,N_27369,N_27174);
and UO_127 (O_127,N_26388,N_27923);
or UO_128 (O_128,N_27067,N_25308);
nor UO_129 (O_129,N_25938,N_28674);
or UO_130 (O_130,N_29578,N_27829);
or UO_131 (O_131,N_29304,N_25504);
nor UO_132 (O_132,N_27282,N_27535);
or UO_133 (O_133,N_26256,N_27370);
nor UO_134 (O_134,N_29971,N_27557);
and UO_135 (O_135,N_25106,N_28653);
or UO_136 (O_136,N_29605,N_26338);
or UO_137 (O_137,N_29138,N_29361);
or UO_138 (O_138,N_27635,N_25847);
nor UO_139 (O_139,N_25679,N_27088);
nand UO_140 (O_140,N_28651,N_26766);
and UO_141 (O_141,N_27420,N_28317);
nor UO_142 (O_142,N_29195,N_29139);
xor UO_143 (O_143,N_28478,N_28064);
and UO_144 (O_144,N_28397,N_26174);
nor UO_145 (O_145,N_27939,N_28218);
nand UO_146 (O_146,N_28363,N_29590);
or UO_147 (O_147,N_25324,N_29410);
and UO_148 (O_148,N_25202,N_26115);
nor UO_149 (O_149,N_29857,N_28538);
xnor UO_150 (O_150,N_26579,N_28333);
nand UO_151 (O_151,N_26876,N_25400);
and UO_152 (O_152,N_28687,N_26216);
nand UO_153 (O_153,N_28196,N_26538);
nor UO_154 (O_154,N_29301,N_29132);
or UO_155 (O_155,N_27375,N_26985);
and UO_156 (O_156,N_25710,N_27171);
xnor UO_157 (O_157,N_28735,N_26067);
nand UO_158 (O_158,N_27993,N_28781);
and UO_159 (O_159,N_25637,N_28736);
nor UO_160 (O_160,N_28185,N_27753);
or UO_161 (O_161,N_27463,N_26955);
xor UO_162 (O_162,N_25761,N_28932);
or UO_163 (O_163,N_27515,N_29977);
xor UO_164 (O_164,N_25765,N_29858);
and UO_165 (O_165,N_28096,N_28536);
and UO_166 (O_166,N_26943,N_25636);
and UO_167 (O_167,N_25798,N_25575);
xnor UO_168 (O_168,N_29347,N_29046);
or UO_169 (O_169,N_29760,N_26408);
or UO_170 (O_170,N_26005,N_28306);
xor UO_171 (O_171,N_25454,N_26845);
nor UO_172 (O_172,N_26756,N_28312);
nor UO_173 (O_173,N_25063,N_26090);
xnor UO_174 (O_174,N_25481,N_25873);
nand UO_175 (O_175,N_29746,N_29443);
and UO_176 (O_176,N_27784,N_25282);
or UO_177 (O_177,N_27508,N_29874);
xor UO_178 (O_178,N_29441,N_28644);
xor UO_179 (O_179,N_26888,N_29551);
and UO_180 (O_180,N_27360,N_26098);
or UO_181 (O_181,N_27502,N_26034);
xnor UO_182 (O_182,N_25806,N_28942);
nand UO_183 (O_183,N_25494,N_29572);
and UO_184 (O_184,N_29735,N_28351);
and UO_185 (O_185,N_29414,N_28328);
nor UO_186 (O_186,N_25766,N_27609);
nand UO_187 (O_187,N_29500,N_28493);
and UO_188 (O_188,N_26467,N_26466);
nand UO_189 (O_189,N_27775,N_28862);
or UO_190 (O_190,N_25573,N_27361);
nor UO_191 (O_191,N_26679,N_25032);
xnor UO_192 (O_192,N_28953,N_29703);
nand UO_193 (O_193,N_28919,N_28889);
or UO_194 (O_194,N_27624,N_27918);
xnor UO_195 (O_195,N_25478,N_27712);
nor UO_196 (O_196,N_25163,N_26587);
and UO_197 (O_197,N_26434,N_25179);
or UO_198 (O_198,N_25066,N_28362);
and UO_199 (O_199,N_25788,N_28393);
nor UO_200 (O_200,N_27715,N_26425);
nor UO_201 (O_201,N_28045,N_27809);
nand UO_202 (O_202,N_25942,N_26383);
or UO_203 (O_203,N_27537,N_27302);
nor UO_204 (O_204,N_28241,N_27599);
nand UO_205 (O_205,N_26659,N_26558);
xor UO_206 (O_206,N_27530,N_25954);
and UO_207 (O_207,N_26671,N_26416);
nand UO_208 (O_208,N_26266,N_27436);
xnor UO_209 (O_209,N_27830,N_28688);
nand UO_210 (O_210,N_25304,N_25095);
nand UO_211 (O_211,N_26418,N_27938);
nand UO_212 (O_212,N_29701,N_27475);
nor UO_213 (O_213,N_28847,N_26000);
and UO_214 (O_214,N_26992,N_27131);
nand UO_215 (O_215,N_26576,N_26946);
xnor UO_216 (O_216,N_29575,N_26727);
nor UO_217 (O_217,N_29745,N_27988);
or UO_218 (O_218,N_29636,N_25362);
nand UO_219 (O_219,N_26450,N_27191);
nand UO_220 (O_220,N_28559,N_27610);
or UO_221 (O_221,N_28716,N_29083);
or UO_222 (O_222,N_26856,N_25709);
nor UO_223 (O_223,N_28398,N_28631);
and UO_224 (O_224,N_28452,N_25924);
xnor UO_225 (O_225,N_27268,N_25609);
nand UO_226 (O_226,N_26161,N_28016);
xnor UO_227 (O_227,N_28660,N_28563);
xnor UO_228 (O_228,N_27150,N_25296);
or UO_229 (O_229,N_29627,N_29331);
or UO_230 (O_230,N_25055,N_25561);
nor UO_231 (O_231,N_26770,N_26973);
xor UO_232 (O_232,N_29385,N_29922);
nor UO_233 (O_233,N_26236,N_25009);
or UO_234 (O_234,N_25287,N_26962);
nor UO_235 (O_235,N_29416,N_27844);
nor UO_236 (O_236,N_28824,N_25414);
nor UO_237 (O_237,N_29173,N_29274);
and UO_238 (O_238,N_27874,N_28239);
nor UO_239 (O_239,N_27910,N_25604);
xor UO_240 (O_240,N_28747,N_26636);
nand UO_241 (O_241,N_27104,N_27183);
and UO_242 (O_242,N_25297,N_27452);
xnor UO_243 (O_243,N_26281,N_29056);
nand UO_244 (O_244,N_27936,N_29952);
nand UO_245 (O_245,N_25728,N_29994);
nand UO_246 (O_246,N_27118,N_27506);
nand UO_247 (O_247,N_29639,N_26283);
and UO_248 (O_248,N_25983,N_28545);
and UO_249 (O_249,N_29126,N_29980);
and UO_250 (O_250,N_26672,N_27294);
nor UO_251 (O_251,N_25716,N_25970);
xor UO_252 (O_252,N_29378,N_29839);
nor UO_253 (O_253,N_27655,N_27745);
and UO_254 (O_254,N_29110,N_28857);
nand UO_255 (O_255,N_26703,N_29661);
and UO_256 (O_256,N_28720,N_26806);
and UO_257 (O_257,N_28331,N_27849);
xor UO_258 (O_258,N_28946,N_28129);
nand UO_259 (O_259,N_26673,N_26974);
or UO_260 (O_260,N_26363,N_29492);
and UO_261 (O_261,N_27134,N_25730);
and UO_262 (O_262,N_29798,N_27002);
or UO_263 (O_263,N_26481,N_29136);
nand UO_264 (O_264,N_26308,N_26299);
nand UO_265 (O_265,N_28214,N_26426);
and UO_266 (O_266,N_26421,N_28580);
nor UO_267 (O_267,N_29912,N_25687);
xor UO_268 (O_268,N_28481,N_25253);
nor UO_269 (O_269,N_28777,N_29634);
nor UO_270 (O_270,N_26428,N_27890);
or UO_271 (O_271,N_27014,N_28237);
nor UO_272 (O_272,N_29523,N_28400);
nand UO_273 (O_273,N_25545,N_28270);
nand UO_274 (O_274,N_25527,N_25118);
or UO_275 (O_275,N_29064,N_29084);
nand UO_276 (O_276,N_27687,N_27980);
nand UO_277 (O_277,N_25752,N_27872);
and UO_278 (O_278,N_27805,N_29781);
nand UO_279 (O_279,N_25469,N_29530);
nor UO_280 (O_280,N_28258,N_29719);
or UO_281 (O_281,N_25852,N_25141);
xnor UO_282 (O_282,N_29695,N_26621);
nand UO_283 (O_283,N_25799,N_28063);
and UO_284 (O_284,N_27042,N_26102);
nor UO_285 (O_285,N_27469,N_26940);
or UO_286 (O_286,N_29566,N_26699);
nand UO_287 (O_287,N_25902,N_26173);
and UO_288 (O_288,N_27676,N_25886);
and UO_289 (O_289,N_25376,N_28366);
nand UO_290 (O_290,N_26244,N_26983);
nand UO_291 (O_291,N_29955,N_29903);
nand UO_292 (O_292,N_25486,N_28034);
nor UO_293 (O_293,N_29219,N_27645);
and UO_294 (O_294,N_27903,N_27194);
nor UO_295 (O_295,N_25223,N_26465);
and UO_296 (O_296,N_28074,N_28370);
xnor UO_297 (O_297,N_29174,N_28508);
nor UO_298 (O_298,N_28087,N_28784);
and UO_299 (O_299,N_29061,N_29997);
nor UO_300 (O_300,N_28975,N_26347);
nor UO_301 (O_301,N_27921,N_28251);
or UO_302 (O_302,N_29583,N_27197);
nand UO_303 (O_303,N_25570,N_29768);
nor UO_304 (O_304,N_27560,N_27995);
nor UO_305 (O_305,N_26270,N_28112);
and UO_306 (O_306,N_27700,N_25707);
nand UO_307 (O_307,N_27093,N_25447);
nor UO_308 (O_308,N_27545,N_25663);
or UO_309 (O_309,N_29226,N_26113);
and UO_310 (O_310,N_26361,N_28826);
and UO_311 (O_311,N_27328,N_25768);
or UO_312 (O_312,N_26160,N_26045);
or UO_313 (O_313,N_29491,N_25751);
or UO_314 (O_314,N_29159,N_26191);
and UO_315 (O_315,N_26092,N_29803);
nor UO_316 (O_316,N_29613,N_29948);
nor UO_317 (O_317,N_27773,N_29853);
xor UO_318 (O_318,N_28721,N_27015);
or UO_319 (O_319,N_25755,N_26459);
nor UO_320 (O_320,N_25582,N_27140);
nor UO_321 (O_321,N_29430,N_27390);
and UO_322 (O_322,N_25309,N_28711);
nand UO_323 (O_323,N_29574,N_25890);
nor UO_324 (O_324,N_26345,N_29468);
and UO_325 (O_325,N_28009,N_28850);
nor UO_326 (O_326,N_27227,N_26397);
nand UO_327 (O_327,N_27598,N_28149);
or UO_328 (O_328,N_26810,N_25876);
and UO_329 (O_329,N_26573,N_28356);
nand UO_330 (O_330,N_25908,N_28396);
nand UO_331 (O_331,N_28590,N_25244);
and UO_332 (O_332,N_27632,N_29614);
and UO_333 (O_333,N_27143,N_29317);
nand UO_334 (O_334,N_26728,N_26264);
xnor UO_335 (O_335,N_27725,N_27453);
nor UO_336 (O_336,N_28471,N_29005);
nor UO_337 (O_337,N_27457,N_29757);
xnor UO_338 (O_338,N_27400,N_25005);
or UO_339 (O_339,N_29223,N_25741);
nor UO_340 (O_340,N_26780,N_29189);
or UO_341 (O_341,N_25937,N_29070);
nor UO_342 (O_342,N_26107,N_26292);
and UO_343 (O_343,N_29622,N_25388);
nand UO_344 (O_344,N_29705,N_25291);
xor UO_345 (O_345,N_28531,N_25148);
or UO_346 (O_346,N_28616,N_29886);
or UO_347 (O_347,N_25608,N_25611);
nand UO_348 (O_348,N_25409,N_29640);
xor UO_349 (O_349,N_29055,N_28534);
or UO_350 (O_350,N_26114,N_25784);
nor UO_351 (O_351,N_26444,N_28128);
nand UO_352 (O_352,N_26831,N_27408);
xnor UO_353 (O_353,N_26061,N_26385);
nor UO_354 (O_354,N_25129,N_28145);
or UO_355 (O_355,N_28722,N_29986);
and UO_356 (O_356,N_26232,N_26189);
and UO_357 (O_357,N_25269,N_28428);
nor UO_358 (O_358,N_27714,N_28421);
nand UO_359 (O_359,N_28766,N_27511);
nor UO_360 (O_360,N_25011,N_28458);
nor UO_361 (O_361,N_27852,N_27384);
or UO_362 (O_362,N_28275,N_28177);
nand UO_363 (O_363,N_29201,N_29733);
or UO_364 (O_364,N_26978,N_27801);
nand UO_365 (O_365,N_26557,N_26799);
and UO_366 (O_366,N_28587,N_25256);
nand UO_367 (O_367,N_29392,N_26582);
and UO_368 (O_368,N_29854,N_29398);
nor UO_369 (O_369,N_26879,N_27358);
nand UO_370 (O_370,N_29453,N_25022);
or UO_371 (O_371,N_28211,N_25412);
nor UO_372 (O_372,N_29013,N_29052);
nand UO_373 (O_373,N_25762,N_28007);
and UO_374 (O_374,N_27837,N_25003);
nor UO_375 (O_375,N_25516,N_26580);
or UO_376 (O_376,N_25025,N_28120);
nor UO_377 (O_377,N_25531,N_25109);
nor UO_378 (O_378,N_28602,N_26566);
or UO_379 (O_379,N_29532,N_29645);
nand UO_380 (O_380,N_28402,N_29076);
and UO_381 (O_381,N_28467,N_26020);
nand UO_382 (O_382,N_26147,N_28224);
and UO_383 (O_383,N_28406,N_25911);
or UO_384 (O_384,N_25422,N_26146);
xnor UO_385 (O_385,N_28760,N_27721);
nor UO_386 (O_386,N_26869,N_28518);
and UO_387 (O_387,N_28540,N_27070);
or UO_388 (O_388,N_29957,N_29704);
nand UO_389 (O_389,N_29506,N_28705);
or UO_390 (O_390,N_26346,N_29783);
or UO_391 (O_391,N_26053,N_27353);
xor UO_392 (O_392,N_29763,N_27876);
nand UO_393 (O_393,N_28530,N_29365);
nor UO_394 (O_394,N_27845,N_28437);
or UO_395 (O_395,N_29095,N_29015);
xor UO_396 (O_396,N_26852,N_27325);
and UO_397 (O_397,N_27387,N_26517);
or UO_398 (O_398,N_26004,N_29211);
nand UO_399 (O_399,N_27432,N_28487);
and UO_400 (O_400,N_28499,N_25172);
xor UO_401 (O_401,N_29377,N_26718);
and UO_402 (O_402,N_29819,N_25581);
nor UO_403 (O_403,N_27096,N_27863);
nor UO_404 (O_404,N_28035,N_26704);
and UO_405 (O_405,N_26323,N_25142);
and UO_406 (O_406,N_29842,N_27940);
nand UO_407 (O_407,N_25206,N_28698);
xnor UO_408 (O_408,N_27727,N_25796);
or UO_409 (O_409,N_27161,N_26712);
nand UO_410 (O_410,N_27717,N_27622);
nor UO_411 (O_411,N_29652,N_26919);
xor UO_412 (O_412,N_27904,N_28191);
xor UO_413 (O_413,N_28097,N_26742);
nor UO_414 (O_414,N_29360,N_29216);
nor UO_415 (O_415,N_25910,N_25535);
nand UO_416 (O_416,N_29893,N_29008);
nand UO_417 (O_417,N_25882,N_27044);
and UO_418 (O_418,N_29447,N_26953);
or UO_419 (O_419,N_25258,N_26022);
nand UO_420 (O_420,N_29477,N_25458);
nor UO_421 (O_421,N_26214,N_29721);
nor UO_422 (O_422,N_28814,N_28247);
nand UO_423 (O_423,N_28659,N_26296);
and UO_424 (O_424,N_25054,N_27544);
or UO_425 (O_425,N_25382,N_26066);
and UO_426 (O_426,N_26838,N_26084);
nand UO_427 (O_427,N_29119,N_27585);
nor UO_428 (O_428,N_29431,N_29236);
or UO_429 (O_429,N_29549,N_26824);
and UO_430 (O_430,N_29460,N_26073);
and UO_431 (O_431,N_29423,N_26003);
or UO_432 (O_432,N_28364,N_28274);
or UO_433 (O_433,N_25398,N_27608);
and UO_434 (O_434,N_25087,N_27473);
or UO_435 (O_435,N_28011,N_25057);
nor UO_436 (O_436,N_26958,N_28694);
xor UO_437 (O_437,N_29764,N_28604);
nor UO_438 (O_438,N_28005,N_27367);
and UO_439 (O_439,N_26219,N_29286);
nor UO_440 (O_440,N_29743,N_25089);
nand UO_441 (O_441,N_26841,N_26805);
nor UO_442 (O_442,N_27204,N_27311);
and UO_443 (O_443,N_25960,N_25379);
and UO_444 (O_444,N_28411,N_29755);
and UO_445 (O_445,N_29908,N_29649);
or UO_446 (O_446,N_28564,N_26651);
nor UO_447 (O_447,N_29455,N_28204);
and UO_448 (O_448,N_26626,N_26362);
nor UO_449 (O_449,N_29945,N_27192);
nand UO_450 (O_450,N_28892,N_27276);
and UO_451 (O_451,N_28319,N_28287);
or UO_452 (O_452,N_29060,N_26882);
nor UO_453 (O_453,N_28355,N_26453);
nand UO_454 (O_454,N_29723,N_27951);
and UO_455 (O_455,N_25984,N_28608);
nand UO_456 (O_456,N_29493,N_27212);
nor UO_457 (O_457,N_27716,N_28193);
nor UO_458 (O_458,N_26653,N_26101);
nor UO_459 (O_459,N_29524,N_29318);
and UO_460 (O_460,N_28947,N_26623);
nand UO_461 (O_461,N_25931,N_26063);
or UO_462 (O_462,N_27316,N_26666);
nand UO_463 (O_463,N_27338,N_26354);
and UO_464 (O_464,N_29972,N_26922);
and UO_465 (O_465,N_27245,N_28524);
nand UO_466 (O_466,N_28868,N_26647);
and UO_467 (O_467,N_27571,N_29330);
or UO_468 (O_468,N_25112,N_25992);
or UO_469 (O_469,N_27402,N_28968);
xor UO_470 (O_470,N_26082,N_27527);
nand UO_471 (O_471,N_25830,N_26850);
or UO_472 (O_472,N_25236,N_26982);
or UO_473 (O_473,N_27695,N_25941);
nor UO_474 (O_474,N_27682,N_27949);
or UO_475 (O_475,N_29959,N_26335);
nor UO_476 (O_476,N_27924,N_25329);
xnor UO_477 (O_477,N_25415,N_29873);
or UO_478 (O_478,N_29457,N_27703);
nand UO_479 (O_479,N_26044,N_26991);
xnor UO_480 (O_480,N_26056,N_26248);
or UO_481 (O_481,N_27968,N_29712);
xnor UO_482 (O_482,N_29038,N_28092);
and UO_483 (O_483,N_25353,N_25295);
or UO_484 (O_484,N_25915,N_27144);
nor UO_485 (O_485,N_28089,N_29438);
nand UO_486 (O_486,N_27326,N_28611);
nor UO_487 (O_487,N_25489,N_28554);
xor UO_488 (O_488,N_29290,N_27769);
nand UO_489 (O_489,N_29671,N_28879);
xnor UO_490 (O_490,N_26083,N_26764);
or UO_491 (O_491,N_29935,N_29635);
and UO_492 (O_492,N_26410,N_26455);
xnor UO_493 (O_493,N_27581,N_25918);
nand UO_494 (O_494,N_26588,N_29394);
and UO_495 (O_495,N_26615,N_28286);
and UO_496 (O_496,N_27634,N_27626);
and UO_497 (O_497,N_27766,N_27549);
xnor UO_498 (O_498,N_25149,N_25850);
nand UO_499 (O_499,N_25781,N_27371);
and UO_500 (O_500,N_27866,N_25292);
or UO_501 (O_501,N_26960,N_28965);
nand UO_502 (O_502,N_27643,N_28980);
or UO_503 (O_503,N_26423,N_27791);
or UO_504 (O_504,N_26237,N_25574);
and UO_505 (O_505,N_27733,N_26141);
nand UO_506 (O_506,N_27329,N_25990);
nor UO_507 (O_507,N_29264,N_26892);
nor UO_508 (O_508,N_26887,N_25613);
and UO_509 (O_509,N_25934,N_26664);
and UO_510 (O_510,N_25712,N_28809);
nand UO_511 (O_511,N_25550,N_29827);
or UO_512 (O_512,N_28436,N_29479);
nand UO_513 (O_513,N_29150,N_28972);
or UO_514 (O_514,N_26605,N_28138);
nand UO_515 (O_515,N_25072,N_28117);
or UO_516 (O_516,N_28322,N_25758);
xor UO_517 (O_517,N_25763,N_28451);
nor UO_518 (O_518,N_29775,N_27808);
nor UO_519 (O_519,N_26039,N_28813);
xor UO_520 (O_520,N_25060,N_28995);
xor UO_521 (O_521,N_29357,N_27063);
or UO_522 (O_522,N_26018,N_28184);
and UO_523 (O_523,N_26087,N_25128);
nand UO_524 (O_524,N_28130,N_25690);
or UO_525 (O_525,N_27049,N_29049);
nor UO_526 (O_526,N_29396,N_29856);
nor UO_527 (O_527,N_25615,N_28325);
nand UO_528 (O_528,N_27577,N_28151);
nor UO_529 (O_529,N_25164,N_27082);
and UO_530 (O_530,N_28885,N_28629);
and UO_531 (O_531,N_25043,N_26552);
or UO_532 (O_532,N_29260,N_27162);
nand UO_533 (O_533,N_28412,N_28100);
and UO_534 (O_534,N_27189,N_26619);
and UO_535 (O_535,N_25444,N_26537);
nand UO_536 (O_536,N_28171,N_27977);
nor UO_537 (O_537,N_29312,N_26451);
nor UO_538 (O_538,N_25452,N_28874);
nand UO_539 (O_539,N_25346,N_26959);
nand UO_540 (O_540,N_25302,N_25969);
and UO_541 (O_541,N_28125,N_29817);
nor UO_542 (O_542,N_29229,N_27831);
or UO_543 (O_543,N_26175,N_25555);
nor UO_544 (O_544,N_26686,N_26263);
and UO_545 (O_545,N_29667,N_25186);
and UO_546 (O_546,N_25365,N_27587);
nand UO_547 (O_547,N_27355,N_28625);
nand UO_548 (O_548,N_27962,N_29143);
and UO_549 (O_549,N_27776,N_29909);
nor UO_550 (O_550,N_26143,N_25879);
and UO_551 (O_551,N_29182,N_25718);
and UO_552 (O_552,N_26395,N_29884);
and UO_553 (O_553,N_26337,N_29001);
nor UO_554 (O_554,N_26844,N_26837);
or UO_555 (O_555,N_27819,N_28751);
nor UO_556 (O_556,N_29251,N_27222);
nand UO_557 (O_557,N_26166,N_27123);
and UO_558 (O_558,N_26559,N_29148);
nand UO_559 (O_559,N_27768,N_27128);
or UO_560 (O_560,N_25343,N_29168);
nand UO_561 (O_561,N_29593,N_25530);
or UO_562 (O_562,N_27350,N_27386);
xnor UO_563 (O_563,N_28380,N_25322);
or UO_564 (O_564,N_27066,N_25303);
nand UO_565 (O_565,N_28550,N_26341);
nor UO_566 (O_566,N_28877,N_29979);
or UO_567 (O_567,N_29875,N_28513);
nor UO_568 (O_568,N_27399,N_27932);
nor UO_569 (O_569,N_25887,N_25482);
and UO_570 (O_570,N_28815,N_28453);
xor UO_571 (O_571,N_28273,N_27957);
nor UO_572 (O_572,N_28209,N_27190);
or UO_573 (O_573,N_29372,N_28558);
and UO_574 (O_574,N_26663,N_29407);
nor UO_575 (O_575,N_29163,N_26560);
nor UO_576 (O_576,N_29464,N_25666);
and UO_577 (O_577,N_29458,N_29494);
nor UO_578 (O_578,N_25159,N_27416);
or UO_579 (O_579,N_27000,N_27315);
nor UO_580 (O_580,N_28354,N_28435);
and UO_581 (O_581,N_25541,N_29461);
nand UO_582 (O_582,N_29662,N_27458);
nand UO_583 (O_583,N_26015,N_28991);
or UO_584 (O_584,N_29533,N_26972);
or UO_585 (O_585,N_25146,N_26789);
nor UO_586 (O_586,N_28198,N_29976);
and UO_587 (O_587,N_28441,N_27548);
xor UO_588 (O_588,N_26855,N_27536);
and UO_589 (O_589,N_26688,N_27750);
nor UO_590 (O_590,N_25791,N_27476);
nor UO_591 (O_591,N_26725,N_29869);
nor UO_592 (O_592,N_29569,N_26187);
xnor UO_593 (O_593,N_26402,N_28940);
nand UO_594 (O_594,N_25667,N_25587);
and UO_595 (O_595,N_27045,N_26431);
and UO_596 (O_596,N_25745,N_25190);
and UO_597 (O_597,N_25044,N_29930);
or UO_598 (O_598,N_28221,N_27417);
or UO_599 (O_599,N_25801,N_25579);
or UO_600 (O_600,N_27855,N_25086);
xnor UO_601 (O_601,N_26629,N_28656);
and UO_602 (O_602,N_26730,N_26916);
nor UO_603 (O_603,N_25340,N_29655);
and UO_604 (O_604,N_27095,N_27461);
nand UO_605 (O_605,N_28585,N_25445);
nand UO_606 (O_606,N_25859,N_27448);
and UO_607 (O_607,N_26956,N_25480);
nand UO_608 (O_608,N_27763,N_29521);
nand UO_609 (O_609,N_27945,N_25396);
xnor UO_610 (O_610,N_28582,N_28283);
nand UO_611 (O_611,N_25335,N_29802);
nor UO_612 (O_612,N_26370,N_27652);
or UO_613 (O_613,N_26889,N_26145);
or UO_614 (O_614,N_25972,N_28310);
nand UO_615 (O_615,N_29849,N_29601);
or UO_616 (O_616,N_27559,N_26105);
and UO_617 (O_617,N_27398,N_25261);
or UO_618 (O_618,N_29204,N_28516);
and UO_619 (O_619,N_29011,N_28663);
and UO_620 (O_620,N_25871,N_29310);
or UO_621 (O_621,N_25927,N_25367);
or UO_622 (O_622,N_27006,N_25284);
nand UO_623 (O_623,N_29267,N_26675);
nor UO_624 (O_624,N_26693,N_26138);
or UO_625 (O_625,N_29826,N_25020);
and UO_626 (O_626,N_26698,N_25705);
and UO_627 (O_627,N_26545,N_26071);
xor UO_628 (O_628,N_25563,N_27211);
nand UO_629 (O_629,N_28334,N_29349);
xnor UO_630 (O_630,N_29063,N_25008);
nand UO_631 (O_631,N_25283,N_28101);
nand UO_632 (O_632,N_29476,N_27611);
nor UO_633 (O_633,N_29599,N_25933);
or UO_634 (O_634,N_28365,N_27658);
nand UO_635 (O_635,N_26567,N_25994);
nand UO_636 (O_636,N_29316,N_28767);
or UO_637 (O_637,N_27196,N_28768);
nor UO_638 (O_638,N_26033,N_29904);
nor UO_639 (O_639,N_27484,N_29386);
or UO_640 (O_640,N_26240,N_27468);
and UO_641 (O_641,N_29259,N_25167);
xor UO_642 (O_642,N_29983,N_27069);
and UO_643 (O_643,N_27480,N_29883);
nand UO_644 (O_644,N_26935,N_28080);
nand UO_645 (O_645,N_28158,N_28790);
nand UO_646 (O_646,N_26289,N_28392);
and UO_647 (O_647,N_29294,N_26254);
and UO_648 (O_648,N_29026,N_28374);
nor UO_649 (O_649,N_28669,N_27300);
nor UO_650 (O_650,N_26936,N_26052);
or UO_651 (O_651,N_26998,N_28152);
and UO_652 (O_652,N_25192,N_25753);
nor UO_653 (O_653,N_27933,N_27443);
and UO_654 (O_654,N_28647,N_29753);
and UO_655 (O_655,N_28867,N_29075);
nand UO_656 (O_656,N_26608,N_29877);
nand UO_657 (O_657,N_29887,N_29951);
and UO_658 (O_658,N_25831,N_27772);
or UO_659 (O_659,N_26597,N_28828);
nand UO_660 (O_660,N_25819,N_29510);
nor UO_661 (O_661,N_28603,N_27201);
and UO_662 (O_662,N_25058,N_29379);
and UO_663 (O_663,N_28808,N_26706);
xor UO_664 (O_664,N_29896,N_25477);
nand UO_665 (O_665,N_25818,N_27771);
or UO_666 (O_666,N_29050,N_26681);
nand UO_667 (O_667,N_28424,N_29560);
nand UO_668 (O_668,N_29245,N_25027);
xor UO_669 (O_669,N_29546,N_26350);
and UO_670 (O_670,N_26961,N_25015);
nor UO_671 (O_671,N_29445,N_27246);
or UO_672 (O_672,N_29689,N_29144);
and UO_673 (O_673,N_27024,N_27862);
and UO_674 (O_674,N_25529,N_26811);
nand UO_675 (O_675,N_28142,N_26534);
xnor UO_676 (O_676,N_27027,N_27956);
or UO_677 (O_677,N_26482,N_27568);
or UO_678 (O_678,N_28061,N_25453);
or UO_679 (O_679,N_26640,N_25926);
nor UO_680 (O_680,N_28628,N_25578);
or UO_681 (O_681,N_25576,N_29346);
nor UO_682 (O_682,N_28997,N_29004);
or UO_683 (O_683,N_26125,N_25413);
or UO_684 (O_684,N_29232,N_25034);
nand UO_685 (O_685,N_25473,N_28150);
and UO_686 (O_686,N_27283,N_26874);
nor UO_687 (O_687,N_28327,N_27251);
nand UO_688 (O_688,N_27130,N_27013);
nor UO_689 (O_689,N_28457,N_26432);
nor UO_690 (O_690,N_26119,N_27133);
xnor UO_691 (O_691,N_28996,N_28566);
nor UO_692 (O_692,N_28578,N_27125);
nor UO_693 (O_693,N_28115,N_29214);
xnor UO_694 (O_694,N_26736,N_28717);
and UO_695 (O_695,N_29104,N_28053);
nand UO_696 (O_696,N_26409,N_29653);
xor UO_697 (O_697,N_26783,N_25495);
and UO_698 (O_698,N_27265,N_26204);
nand UO_699 (O_699,N_27526,N_27364);
or UO_700 (O_700,N_26201,N_27915);
and UO_701 (O_701,N_26123,N_29792);
or UO_702 (O_702,N_25042,N_28732);
nor UO_703 (O_703,N_25953,N_27948);
nand UO_704 (O_704,N_27459,N_28304);
nor UO_705 (O_705,N_29452,N_26367);
xnor UO_706 (O_706,N_26895,N_26740);
and UO_707 (O_707,N_26899,N_26967);
nor UO_708 (O_708,N_29244,N_25133);
or UO_709 (O_709,N_26507,N_27865);
xor UO_710 (O_710,N_25313,N_28915);
nor UO_711 (O_711,N_27654,N_29212);
nor UO_712 (O_712,N_29810,N_26070);
nor UO_713 (O_713,N_25554,N_26530);
or UO_714 (O_714,N_25098,N_25746);
nand UO_715 (O_715,N_26150,N_27992);
or UO_716 (O_716,N_28132,N_29339);
nand UO_717 (O_717,N_26218,N_26374);
or UO_718 (O_718,N_28532,N_26633);
nand UO_719 (O_719,N_26639,N_26276);
xnor UO_720 (O_720,N_26225,N_28192);
and UO_721 (O_721,N_25851,N_26069);
nor UO_722 (O_722,N_27856,N_28292);
or UO_723 (O_723,N_25776,N_26912);
nor UO_724 (O_724,N_27318,N_29754);
nand UO_725 (O_725,N_26504,N_29535);
xnor UO_726 (O_726,N_27184,N_25317);
nor UO_727 (O_727,N_29255,N_26628);
or UO_728 (O_728,N_29953,N_25891);
or UO_729 (O_729,N_27572,N_26348);
or UO_730 (O_730,N_27942,N_26377);
nand UO_731 (O_731,N_26617,N_25227);
nand UO_732 (O_732,N_29069,N_27792);
nor UO_733 (O_733,N_26109,N_28741);
and UO_734 (O_734,N_29716,N_26340);
and UO_735 (O_735,N_28020,N_27954);
nand UO_736 (O_736,N_29870,N_28743);
or UO_737 (O_737,N_25270,N_29344);
or UO_738 (O_738,N_25393,N_27664);
and UO_739 (O_739,N_29125,N_28290);
xnor UO_740 (O_740,N_29834,N_25161);
nand UO_741 (O_741,N_29960,N_25446);
nor UO_742 (O_742,N_26258,N_29550);
or UO_743 (O_743,N_29592,N_26683);
nor UO_744 (O_744,N_29167,N_29910);
xor UO_745 (O_745,N_26172,N_26937);
or UO_746 (O_746,N_26261,N_29197);
nor UO_747 (O_747,N_28922,N_25021);
nand UO_748 (O_748,N_28352,N_25471);
nor UO_749 (O_749,N_25889,N_27147);
nor UO_750 (O_750,N_25212,N_29140);
or UO_751 (O_751,N_27965,N_25203);
xnor UO_752 (O_752,N_28379,N_26795);
or UO_753 (O_753,N_29591,N_25884);
and UO_754 (O_754,N_25677,N_28029);
and UO_755 (O_755,N_29405,N_25790);
nor UO_756 (O_756,N_28443,N_28869);
nand UO_757 (O_757,N_29288,N_26088);
and UO_758 (O_758,N_27106,N_25077);
or UO_759 (O_759,N_26952,N_26868);
nand UO_760 (O_760,N_28770,N_29362);
or UO_761 (O_761,N_29715,N_25858);
and UO_762 (O_762,N_27403,N_29256);
or UO_763 (O_763,N_25328,N_26866);
or UO_764 (O_764,N_27623,N_27116);
nand UO_765 (O_765,N_29192,N_26394);
and UO_766 (O_766,N_28535,N_29619);
xor UO_767 (O_767,N_29343,N_26834);
or UO_768 (O_768,N_28361,N_25111);
xnor UO_769 (O_769,N_25334,N_28473);
xnor UO_770 (O_770,N_25117,N_28910);
xnor UO_771 (O_771,N_29230,N_27898);
nand UO_772 (O_772,N_25364,N_26539);
and UO_773 (O_773,N_28391,N_29248);
nand UO_774 (O_774,N_26999,N_27823);
xor UO_775 (O_775,N_27195,N_29730);
xnor UO_776 (O_776,N_26313,N_29088);
or UO_777 (O_777,N_25564,N_28099);
and UO_778 (O_778,N_26328,N_25944);
nand UO_779 (O_779,N_28226,N_27007);
nor UO_780 (O_780,N_27552,N_28308);
or UO_781 (O_781,N_27026,N_29633);
nand UO_782 (O_782,N_29141,N_25280);
or UO_783 (O_783,N_26392,N_26802);
and UO_784 (O_784,N_29309,N_26014);
and UO_785 (O_785,N_26037,N_25448);
nand UO_786 (O_786,N_27802,N_26966);
or UO_787 (O_787,N_28797,N_25517);
nand UO_788 (O_788,N_26769,N_29561);
nor UO_789 (O_789,N_25213,N_29890);
nor UO_790 (O_790,N_27847,N_25792);
or UO_791 (O_791,N_25357,N_28785);
xnor UO_792 (O_792,N_25047,N_27729);
nor UO_793 (O_793,N_25820,N_25294);
or UO_794 (O_794,N_27699,N_26011);
and UO_795 (O_795,N_27807,N_25441);
and UO_796 (O_796,N_28805,N_28225);
and UO_797 (O_797,N_28533,N_25706);
and UO_798 (O_798,N_27158,N_29077);
or UO_799 (O_799,N_29419,N_27730);
nand UO_800 (O_800,N_27788,N_27704);
nand UO_801 (O_801,N_29488,N_29880);
nor UO_802 (O_802,N_29283,N_25059);
or UO_803 (O_803,N_29830,N_29998);
or UO_804 (O_804,N_25958,N_26447);
nand UO_805 (O_805,N_28413,N_25693);
nand UO_806 (O_806,N_27253,N_26180);
nand UO_807 (O_807,N_25828,N_28870);
or UO_808 (O_808,N_29275,N_29185);
xnor UO_809 (O_809,N_28164,N_29879);
nand UO_810 (O_810,N_25612,N_26412);
nor UO_811 (O_811,N_26816,N_28945);
nor UO_812 (O_812,N_26042,N_25125);
nor UO_813 (O_813,N_25814,N_27112);
and UO_814 (O_814,N_26896,N_26762);
nor UO_815 (O_815,N_29611,N_27697);
or UO_816 (O_816,N_27539,N_26803);
xor UO_817 (O_817,N_26364,N_28012);
nand UO_818 (O_818,N_26032,N_28180);
xor UO_819 (O_819,N_29122,N_27011);
xor UO_820 (O_820,N_27671,N_28254);
xnor UO_821 (O_821,N_28048,N_26583);
or UO_822 (O_822,N_25316,N_28316);
or UO_823 (O_823,N_28110,N_27958);
and UO_824 (O_824,N_25016,N_25399);
and UO_825 (O_825,N_25872,N_28840);
and UO_826 (O_826,N_26784,N_28713);
nand UO_827 (O_827,N_27306,N_29040);
or UO_828 (O_828,N_25767,N_25523);
or UO_829 (O_829,N_25134,N_29779);
and UO_830 (O_830,N_25174,N_28817);
and UO_831 (O_831,N_29442,N_26915);
or UO_832 (O_832,N_29067,N_29832);
nor UO_833 (O_833,N_26928,N_26941);
and UO_834 (O_834,N_28692,N_27119);
or UO_835 (O_835,N_29135,N_27477);
nor UO_836 (O_836,N_26731,N_28811);
or UO_837 (O_837,N_26349,N_29929);
nor UO_838 (O_838,N_28296,N_27908);
nand UO_839 (O_839,N_26190,N_25131);
nor UO_840 (O_840,N_29941,N_29631);
or UO_841 (O_841,N_29329,N_26242);
and UO_842 (O_842,N_26768,N_25907);
nor UO_843 (O_843,N_28260,N_27913);
nor UO_844 (O_844,N_26572,N_28375);
or UO_845 (O_845,N_25349,N_25821);
or UO_846 (O_846,N_27894,N_29654);
or UO_847 (O_847,N_28509,N_27359);
and UO_848 (O_848,N_25209,N_29106);
or UO_849 (O_849,N_29336,N_28685);
nand UO_850 (O_850,N_29608,N_29044);
and UO_851 (O_851,N_26533,N_25932);
or UO_852 (O_852,N_27439,N_28299);
xnor UO_853 (O_853,N_28483,N_29381);
xnor UO_854 (O_854,N_25041,N_26749);
nand UO_855 (O_855,N_28935,N_27381);
or UO_856 (O_856,N_25662,N_25694);
or UO_857 (O_857,N_26275,N_28381);
and UO_858 (O_858,N_25298,N_26165);
xnor UO_859 (O_859,N_26169,N_25996);
nand UO_860 (O_860,N_29923,N_25102);
and UO_861 (O_861,N_25275,N_26188);
nor UO_862 (O_862,N_28622,N_26311);
nor UO_863 (O_863,N_28165,N_27815);
and UO_864 (O_864,N_28734,N_29732);
xor UO_865 (O_865,N_25084,N_25000);
nand UO_866 (O_866,N_25305,N_26336);
nand UO_867 (O_867,N_29502,N_27225);
nor UO_868 (O_868,N_26914,N_26381);
and UO_869 (O_869,N_29162,N_28978);
or UO_870 (O_870,N_29371,N_29925);
and UO_871 (O_871,N_29587,N_26905);
and UO_872 (O_872,N_28780,N_27550);
nor UO_873 (O_873,N_27906,N_26304);
and UO_874 (O_874,N_27892,N_28888);
xor UO_875 (O_875,N_27250,N_27796);
or UO_876 (O_876,N_29668,N_26076);
nor UO_877 (O_877,N_28321,N_27028);
xor UO_878 (O_878,N_25732,N_25896);
or UO_879 (O_879,N_29632,N_26771);
nor UO_880 (O_880,N_29595,N_28737);
and UO_881 (O_881,N_29436,N_28557);
and UO_882 (O_882,N_26965,N_26049);
or UO_883 (O_883,N_28610,N_28598);
nand UO_884 (O_884,N_28433,N_25534);
nand UO_885 (O_885,N_29152,N_29609);
or UO_886 (O_886,N_29686,N_27561);
nor UO_887 (O_887,N_25961,N_28448);
and UO_888 (O_888,N_28866,N_28238);
or UO_889 (O_889,N_27762,N_29072);
or UO_890 (O_890,N_27238,N_26532);
and UO_891 (O_891,N_28594,N_25750);
or UO_892 (O_892,N_27237,N_25120);
and UO_893 (O_893,N_29171,N_29678);
nand UO_894 (O_894,N_25391,N_27893);
nand UO_895 (O_895,N_28326,N_27025);
nand UO_896 (O_896,N_29323,N_28027);
or UO_897 (O_897,N_25878,N_26827);
nand UO_898 (O_898,N_26790,N_26565);
nor UO_899 (O_899,N_27744,N_25749);
nor UO_900 (O_900,N_27944,N_26678);
or UO_901 (O_901,N_28618,N_28405);
or UO_902 (O_902,N_28070,N_27922);
nand UO_903 (O_903,N_25426,N_25491);
xor UO_904 (O_904,N_29094,N_25082);
nor UO_905 (O_905,N_25711,N_28748);
and UO_906 (O_906,N_28245,N_28044);
and UO_907 (O_907,N_28078,N_28753);
or UO_908 (O_908,N_25080,N_26871);
and UO_909 (O_909,N_26355,N_27339);
nor UO_910 (O_910,N_29202,N_28541);
nor UO_911 (O_911,N_27129,N_27239);
and UO_912 (O_912,N_25544,N_27777);
and UO_913 (O_913,N_27077,N_27324);
or UO_914 (O_914,N_28505,N_28205);
or UO_915 (O_915,N_26413,N_26751);
nor UO_916 (O_916,N_27354,N_27152);
nor UO_917 (O_917,N_26217,N_27202);
and UO_918 (O_918,N_27896,N_25525);
nand UO_919 (O_919,N_27696,N_28023);
and UO_920 (O_920,N_27051,N_26947);
xor UO_921 (O_921,N_25100,N_27199);
nand UO_922 (O_922,N_27596,N_27926);
nor UO_923 (O_923,N_25945,N_26930);
nand UO_924 (O_924,N_25638,N_28109);
or UO_925 (O_925,N_28896,N_26944);
and UO_926 (O_926,N_27365,N_27665);
nand UO_927 (O_927,N_28654,N_28055);
xor UO_928 (O_928,N_29429,N_26980);
and UO_929 (O_929,N_27649,N_26885);
and UO_930 (O_930,N_26932,N_25397);
and UO_931 (O_931,N_28459,N_27198);
and UO_932 (O_932,N_27575,N_29670);
and UO_933 (O_933,N_26792,N_28108);
or UO_934 (O_934,N_29456,N_28854);
nand UO_935 (O_935,N_29559,N_29913);
nand UO_936 (O_936,N_28037,N_26642);
and UO_937 (O_937,N_25366,N_28105);
and UO_938 (O_938,N_29415,N_28252);
or UO_939 (O_939,N_26707,N_25250);
xnor UO_940 (O_940,N_29607,N_28820);
or UO_941 (O_941,N_29841,N_25565);
and UO_942 (O_942,N_26196,N_29543);
nor UO_943 (O_943,N_26195,N_26696);
xor UO_944 (O_944,N_25623,N_28126);
or UO_945 (O_945,N_28507,N_25210);
xnor UO_946 (O_946,N_27694,N_25017);
nor UO_947 (O_947,N_28071,N_27970);
or UO_948 (O_948,N_27236,N_25130);
nor UO_949 (O_949,N_26198,N_25228);
or UO_950 (O_950,N_26124,N_27787);
and UO_951 (O_951,N_29271,N_27235);
or UO_952 (O_952,N_25583,N_25464);
nand UO_953 (O_953,N_29938,N_26010);
nor UO_954 (O_954,N_29121,N_26521);
nor UO_955 (O_955,N_25672,N_26078);
nor UO_956 (O_956,N_29556,N_26494);
and UO_957 (O_957,N_26765,N_26464);
xor UO_958 (O_958,N_27705,N_28015);
nand UO_959 (O_959,N_29175,N_29739);
or UO_960 (O_960,N_25476,N_27068);
nor UO_961 (O_961,N_26531,N_27058);
or UO_962 (O_962,N_29526,N_26060);
and UO_963 (O_963,N_28371,N_28049);
nand UO_964 (O_964,N_27838,N_29233);
or UO_965 (O_965,N_29969,N_28776);
nor UO_966 (O_966,N_25394,N_27220);
nand UO_967 (O_967,N_28954,N_27646);
or UO_968 (O_968,N_29885,N_25702);
nor UO_969 (O_969,N_27720,N_27751);
nand UO_970 (O_970,N_25390,N_25355);
nand UO_971 (O_971,N_27160,N_28763);
nand UO_972 (O_972,N_27604,N_28742);
and UO_973 (O_973,N_27994,N_26215);
nand UO_974 (O_974,N_29988,N_25438);
or UO_975 (O_975,N_25597,N_25507);
nand UO_976 (O_976,N_27351,N_29474);
and UO_977 (O_977,N_26542,N_28271);
or UO_978 (O_978,N_28342,N_28030);
or UO_979 (O_979,N_25675,N_25053);
or UO_980 (O_980,N_29105,N_28293);
nand UO_981 (O_981,N_26891,N_28232);
or UO_982 (O_982,N_26815,N_28340);
nor UO_983 (O_983,N_28739,N_28841);
nand UO_984 (O_984,N_29580,N_29536);
nor UO_985 (O_985,N_25656,N_26280);
and UO_986 (O_986,N_28738,N_25721);
nor UO_987 (O_987,N_28676,N_27297);
and UO_988 (O_988,N_26710,N_26500);
or UO_989 (O_989,N_27749,N_25634);
nor UO_990 (O_990,N_29772,N_26589);
nor UO_991 (O_991,N_26259,N_28782);
or UO_992 (O_992,N_28799,N_29031);
nor UO_993 (O_993,N_27357,N_25122);
or UO_994 (O_994,N_27638,N_26859);
nand UO_995 (O_995,N_28256,N_28756);
or UO_996 (O_996,N_29036,N_29444);
nand UO_997 (O_997,N_27967,N_27102);
nand UO_998 (O_998,N_28802,N_26951);
or UO_999 (O_999,N_29099,N_29151);
or UO_1000 (O_1000,N_28407,N_29297);
and UO_1001 (O_1001,N_27778,N_27155);
and UO_1002 (O_1002,N_26429,N_29872);
nand UO_1003 (O_1003,N_27758,N_28837);
and UO_1004 (O_1004,N_25526,N_27746);
and UO_1005 (O_1005,N_29486,N_26181);
nand UO_1006 (O_1006,N_26669,N_28259);
or UO_1007 (O_1007,N_27415,N_25888);
or UO_1008 (O_1008,N_28675,N_25770);
and UO_1009 (O_1009,N_27035,N_27498);
nand UO_1010 (O_1010,N_29629,N_27474);
nor UO_1011 (O_1011,N_25514,N_29435);
xor UO_1012 (O_1012,N_29900,N_29931);
or UO_1013 (O_1013,N_25880,N_25330);
nand UO_1014 (O_1014,N_25266,N_27651);
nand UO_1015 (O_1015,N_25169,N_27881);
and UO_1016 (O_1016,N_26525,N_27786);
xnor UO_1017 (O_1017,N_28056,N_28313);
and UO_1018 (O_1018,N_26677,N_28210);
and UO_1019 (O_1019,N_28709,N_26048);
xor UO_1020 (O_1020,N_26858,N_28929);
and UO_1021 (O_1021,N_28931,N_28839);
or UO_1022 (O_1022,N_25006,N_27731);
and UO_1023 (O_1023,N_29656,N_25370);
nor UO_1024 (O_1024,N_26319,N_26205);
xnor UO_1025 (O_1025,N_28906,N_26449);
nor UO_1026 (O_1026,N_27825,N_27656);
and UO_1027 (O_1027,N_27071,N_28013);
or UO_1028 (O_1028,N_27181,N_28575);
nand UO_1029 (O_1029,N_25363,N_25234);
nand UO_1030 (O_1030,N_28952,N_28160);
nor UO_1031 (O_1031,N_25620,N_25669);
or UO_1032 (O_1032,N_26590,N_25127);
nand UO_1033 (O_1033,N_29927,N_27588);
or UO_1034 (O_1034,N_27009,N_27824);
nand UO_1035 (O_1035,N_27503,N_26343);
or UO_1036 (O_1036,N_28921,N_29454);
and UO_1037 (O_1037,N_27607,N_28856);
nor UO_1038 (O_1038,N_29418,N_26255);
nor UO_1039 (O_1039,N_26748,N_25528);
and UO_1040 (O_1040,N_26528,N_25191);
or UO_1041 (O_1041,N_28728,N_26814);
nand UO_1042 (O_1042,N_28050,N_27570);
nor UO_1043 (O_1043,N_28038,N_28740);
nor UO_1044 (O_1044,N_28490,N_26227);
and UO_1045 (O_1045,N_26779,N_25183);
nand UO_1046 (O_1046,N_27810,N_26711);
or UO_1047 (O_1047,N_27685,N_29702);
xor UO_1048 (O_1048,N_28686,N_28228);
nand UO_1049 (O_1049,N_28159,N_25805);
nand UO_1050 (O_1050,N_26272,N_29576);
or UO_1051 (O_1051,N_26661,N_26456);
nand UO_1052 (O_1052,N_28028,N_25840);
nor UO_1053 (O_1053,N_27884,N_26591);
and UO_1054 (O_1054,N_29892,N_26875);
or UO_1055 (O_1055,N_29137,N_27060);
and UO_1056 (O_1056,N_26251,N_25150);
and UO_1057 (O_1057,N_29326,N_28267);
xnor UO_1058 (O_1058,N_29528,N_25233);
or UO_1059 (O_1059,N_26526,N_29624);
nor UO_1060 (O_1060,N_26260,N_26322);
or UO_1061 (O_1061,N_25885,N_28900);
nor UO_1062 (O_1062,N_27972,N_26407);
and UO_1063 (O_1063,N_28526,N_26006);
and UO_1064 (O_1064,N_27410,N_25010);
and UO_1065 (O_1065,N_29831,N_26911);
xnor UO_1066 (O_1066,N_29337,N_25976);
nand UO_1067 (O_1067,N_29690,N_27916);
or UO_1068 (O_1068,N_26515,N_26357);
or UO_1069 (O_1069,N_28075,N_26986);
and UO_1070 (O_1070,N_26372,N_25649);
nor UO_1071 (O_1071,N_28492,N_26157);
nor UO_1072 (O_1072,N_25225,N_26963);
or UO_1073 (O_1073,N_28979,N_27447);
xnor UO_1074 (O_1074,N_27205,N_26556);
nand UO_1075 (O_1075,N_27200,N_28795);
xnor UO_1076 (O_1076,N_29440,N_27219);
nor UO_1077 (O_1077,N_25968,N_29366);
nor UO_1078 (O_1078,N_29597,N_26641);
or UO_1079 (O_1079,N_28102,N_28623);
or UO_1080 (O_1080,N_27046,N_27517);
xor UO_1081 (O_1081,N_26870,N_26265);
nand UO_1082 (O_1082,N_26949,N_27397);
xnor UO_1083 (O_1083,N_27551,N_29683);
nand UO_1084 (O_1084,N_27254,N_27481);
and UO_1085 (O_1085,N_29648,N_29751);
xor UO_1086 (O_1086,N_29864,N_28925);
xnor UO_1087 (O_1087,N_27256,N_27584);
nand UO_1088 (O_1088,N_26247,N_28609);
and UO_1089 (O_1089,N_25778,N_26373);
and UO_1090 (O_1090,N_25857,N_28514);
and UO_1091 (O_1091,N_27428,N_29497);
and UO_1092 (O_1092,N_26129,N_28173);
or UO_1093 (O_1093,N_29924,N_28123);
and UO_1094 (O_1094,N_26773,N_25105);
or UO_1095 (O_1095,N_27868,N_29355);
and UO_1096 (O_1096,N_28970,N_29573);
nor UO_1097 (O_1097,N_25951,N_26880);
or UO_1098 (O_1098,N_25747,N_28645);
and UO_1099 (O_1099,N_25854,N_29837);
and UO_1100 (O_1100,N_29053,N_28330);
nand UO_1101 (O_1101,N_27414,N_27882);
nand UO_1102 (O_1102,N_28548,N_27709);
nand UO_1103 (O_1103,N_27193,N_27827);
or UO_1104 (O_1104,N_25252,N_27689);
nor UO_1105 (O_1105,N_27019,N_28234);
or UO_1106 (O_1106,N_26562,N_25811);
nor UO_1107 (O_1107,N_29672,N_29073);
or UO_1108 (O_1108,N_29545,N_29707);
nand UO_1109 (O_1109,N_29537,N_28318);
or UO_1110 (O_1110,N_28880,N_27218);
or UO_1111 (O_1111,N_25451,N_29547);
nand UO_1112 (O_1112,N_26457,N_28666);
nand UO_1113 (O_1113,N_25074,N_25900);
and UO_1114 (O_1114,N_26170,N_28955);
or UO_1115 (O_1115,N_29799,N_26782);
or UO_1116 (O_1116,N_28133,N_28329);
nor UO_1117 (O_1117,N_27795,N_29804);
xnor UO_1118 (O_1118,N_26709,N_29918);
and UO_1119 (O_1119,N_29863,N_25501);
nand UO_1120 (O_1120,N_26017,N_27500);
nor UO_1121 (O_1121,N_25062,N_28083);
nor UO_1122 (O_1122,N_28242,N_29131);
nor UO_1123 (O_1123,N_27433,N_29246);
and UO_1124 (O_1124,N_28388,N_27594);
or UO_1125 (O_1125,N_29641,N_27389);
or UO_1126 (O_1126,N_26529,N_29650);
and UO_1127 (O_1127,N_28442,N_29483);
and UO_1128 (O_1128,N_26825,N_29750);
or UO_1129 (O_1129,N_27435,N_29166);
and UO_1130 (O_1130,N_26819,N_25839);
xnor UO_1131 (O_1131,N_26293,N_25215);
nand UO_1132 (O_1132,N_25779,N_29919);
or UO_1133 (O_1133,N_28464,N_28291);
nor UO_1134 (O_1134,N_25064,N_28983);
nand UO_1135 (O_1135,N_28417,N_29187);
or UO_1136 (O_1136,N_27031,N_25553);
and UO_1137 (O_1137,N_28382,N_26329);
or UO_1138 (O_1138,N_26514,N_28190);
nand UO_1139 (O_1139,N_29677,N_26002);
or UO_1140 (O_1140,N_27124,N_25760);
or UO_1141 (O_1141,N_26239,N_27937);
nand UO_1142 (O_1142,N_28439,N_28484);
or UO_1143 (O_1143,N_26200,N_28263);
nand UO_1144 (O_1144,N_26279,N_26854);
nand UO_1145 (O_1145,N_27122,N_26886);
and UO_1146 (O_1146,N_29851,N_29554);
nor UO_1147 (O_1147,N_27739,N_29958);
and UO_1148 (O_1148,N_29413,N_27488);
and UO_1149 (O_1149,N_28004,N_29623);
nand UO_1150 (O_1150,N_28522,N_26957);
and UO_1151 (O_1151,N_28022,N_25642);
nor UO_1152 (O_1152,N_26415,N_28842);
xnor UO_1153 (O_1153,N_29598,N_28746);
or UO_1154 (O_1154,N_27048,N_25543);
nand UO_1155 (O_1155,N_26685,N_28107);
and UO_1156 (O_1156,N_26984,N_27834);
xnor UO_1157 (O_1157,N_25181,N_27732);
nand UO_1158 (O_1158,N_28523,N_26433);
nand UO_1159 (O_1159,N_25607,N_25966);
xnor UO_1160 (O_1160,N_27159,N_29417);
nand UO_1161 (O_1161,N_26945,N_29966);
xnor UO_1162 (O_1162,N_28917,N_28914);
nor UO_1163 (O_1163,N_28701,N_29180);
nand UO_1164 (O_1164,N_25993,N_29354);
or UO_1165 (O_1165,N_27870,N_29567);
nor UO_1166 (O_1166,N_25979,N_27684);
nor UO_1167 (O_1167,N_26008,N_26257);
nand UO_1168 (O_1168,N_28169,N_27032);
nor UO_1169 (O_1169,N_27332,N_28017);
or UO_1170 (O_1170,N_26096,N_27178);
nor UO_1171 (O_1171,N_25865,N_28804);
and UO_1172 (O_1172,N_26031,N_28893);
nor UO_1173 (O_1173,N_29555,N_25518);
nor UO_1174 (O_1174,N_28118,N_29243);
and UO_1175 (O_1175,N_28157,N_26176);
or UO_1176 (O_1176,N_25263,N_25369);
nand UO_1177 (O_1177,N_25853,N_27100);
nand UO_1178 (O_1178,N_27540,N_26401);
and UO_1179 (O_1179,N_27472,N_25521);
nand UO_1180 (O_1180,N_26804,N_26055);
xor UO_1181 (O_1181,N_28520,N_28136);
nand UO_1182 (O_1182,N_25170,N_26057);
and UO_1183 (O_1183,N_27308,N_25734);
and UO_1184 (O_1184,N_26212,N_27647);
or UO_1185 (O_1185,N_26396,N_29847);
nand UO_1186 (O_1186,N_29770,N_27422);
or UO_1187 (O_1187,N_28971,N_27366);
xor UO_1188 (O_1188,N_25769,N_29043);
xor UO_1189 (O_1189,N_26760,N_25384);
and UO_1190 (O_1190,N_26917,N_27493);
nand UO_1191 (O_1191,N_29333,N_25153);
or UO_1192 (O_1192,N_28419,N_28565);
and UO_1193 (O_1193,N_25499,N_29562);
or UO_1194 (O_1194,N_27177,N_27672);
xor UO_1195 (O_1195,N_27578,N_29041);
or UO_1196 (O_1196,N_28219,N_25039);
nor UO_1197 (O_1197,N_29939,N_29352);
nor UO_1198 (O_1198,N_29387,N_27105);
and UO_1199 (O_1199,N_27295,N_29029);
or UO_1200 (O_1200,N_25701,N_25789);
or UO_1201 (O_1201,N_27167,N_25344);
nand UO_1202 (O_1202,N_28315,N_26667);
or UO_1203 (O_1203,N_25359,N_26842);
nor UO_1204 (O_1204,N_29325,N_28134);
nand UO_1205 (O_1205,N_26996,N_28199);
or UO_1206 (O_1206,N_27127,N_28233);
nand UO_1207 (O_1207,N_27176,N_29451);
nor UO_1208 (O_1208,N_29433,N_25488);
nand UO_1209 (O_1209,N_27086,N_28733);
or UO_1210 (O_1210,N_25922,N_28348);
xnor UO_1211 (O_1211,N_28344,N_27089);
or UO_1212 (O_1212,N_27374,N_27487);
nor UO_1213 (O_1213,N_27172,N_27555);
and UO_1214 (O_1214,N_25254,N_29475);
nor UO_1215 (O_1215,N_25165,N_28834);
nand UO_1216 (O_1216,N_29298,N_28156);
and UO_1217 (O_1217,N_25549,N_25874);
nand UO_1218 (O_1218,N_29679,N_28081);
nor UO_1219 (O_1219,N_27307,N_26249);
or UO_1220 (O_1220,N_27146,N_25519);
nand UO_1221 (O_1221,N_26631,N_26737);
and UO_1222 (O_1222,N_27010,N_27040);
or UO_1223 (O_1223,N_25580,N_29637);
or UO_1224 (O_1224,N_25551,N_29681);
nand UO_1225 (O_1225,N_28489,N_29840);
nand UO_1226 (O_1226,N_26674,N_29664);
nand UO_1227 (O_1227,N_26207,N_25091);
and UO_1228 (O_1228,N_27612,N_25592);
nor UO_1229 (O_1229,N_28427,N_28086);
nor UO_1230 (O_1230,N_28787,N_27783);
or UO_1231 (O_1231,N_27252,N_29161);
nor UO_1232 (O_1232,N_28104,N_29170);
and UO_1233 (O_1233,N_28843,N_26971);
xor UO_1234 (O_1234,N_26139,N_25321);
nand UO_1235 (O_1235,N_27430,N_27963);
nor UO_1236 (O_1236,N_26498,N_25929);
and UO_1237 (O_1237,N_26156,N_26439);
nand UO_1238 (O_1238,N_28206,N_29982);
nor UO_1239 (O_1239,N_27547,N_27735);
nor UO_1240 (O_1240,N_26081,N_28657);
and UO_1241 (O_1241,N_25332,N_29586);
nor UO_1242 (O_1242,N_28786,N_26505);
and UO_1243 (O_1243,N_28485,N_26112);
nand UO_1244 (O_1244,N_25877,N_25704);
or UO_1245 (O_1245,N_25496,N_29087);
and UO_1246 (O_1246,N_28803,N_28726);
nor UO_1247 (O_1247,N_27407,N_26934);
and UO_1248 (O_1248,N_29823,N_28079);
nor UO_1249 (O_1249,N_25378,N_27880);
or UO_1250 (O_1250,N_29696,N_25940);
nor UO_1251 (O_1251,N_26624,N_27016);
nand UO_1252 (O_1252,N_26419,N_28414);
nand UO_1253 (O_1253,N_27438,N_27274);
nor UO_1254 (O_1254,N_29129,N_28724);
xor UO_1255 (O_1255,N_29936,N_27244);
xnor UO_1256 (O_1256,N_26253,N_26411);
nor UO_1257 (O_1257,N_27210,N_29024);
or UO_1258 (O_1258,N_28729,N_26077);
nand UO_1259 (O_1259,N_26575,N_27793);
or UO_1260 (O_1260,N_25068,N_28261);
and UO_1261 (O_1261,N_27764,N_27277);
nor UO_1262 (O_1262,N_25997,N_29968);
nand UO_1263 (O_1263,N_29726,N_28470);
nor UO_1264 (O_1264,N_29756,N_27395);
and UO_1265 (O_1265,N_26233,N_26676);
nor UO_1266 (O_1266,N_25031,N_25697);
and UO_1267 (O_1267,N_28444,N_27335);
and UO_1268 (O_1268,N_29711,N_25147);
nor UO_1269 (O_1269,N_25199,N_29249);
nand UO_1270 (O_1270,N_26016,N_29231);
and UO_1271 (O_1271,N_28095,N_29269);
nand UO_1272 (O_1272,N_26131,N_26182);
and UO_1273 (O_1273,N_29950,N_29388);
nor UO_1274 (O_1274,N_27990,N_25078);
xnor UO_1275 (O_1275,N_29058,N_27759);
xor UO_1276 (O_1276,N_27267,N_28718);
and UO_1277 (O_1277,N_28783,N_27846);
nand UO_1278 (O_1278,N_25905,N_28998);
or UO_1279 (O_1279,N_28626,N_27344);
or UO_1280 (O_1280,N_25071,N_26503);
nand UO_1281 (O_1281,N_29773,N_29651);
nand UO_1282 (O_1282,N_27421,N_29882);
and UO_1283 (O_1283,N_27303,N_27352);
nor UO_1284 (O_1284,N_25602,N_28727);
and UO_1285 (O_1285,N_27372,N_25834);
or UO_1286 (O_1286,N_25046,N_28977);
and UO_1287 (O_1287,N_29270,N_26904);
nand UO_1288 (O_1288,N_29708,N_26108);
nor UO_1289 (O_1289,N_28827,N_28266);
nand UO_1290 (O_1290,N_27765,N_26068);
nand UO_1291 (O_1291,N_25567,N_26898);
and UO_1292 (O_1292,N_25599,N_26040);
or UO_1293 (O_1293,N_29828,N_28496);
nor UO_1294 (O_1294,N_25052,N_26406);
nor UO_1295 (O_1295,N_25351,N_29353);
nor UO_1296 (O_1296,N_29531,N_25633);
or UO_1297 (O_1297,N_26510,N_28933);
nand UO_1298 (O_1298,N_26268,N_26997);
or UO_1299 (O_1299,N_26046,N_25647);
nor UO_1300 (O_1300,N_29898,N_28494);
or UO_1301 (O_1301,N_25029,N_27593);
and UO_1302 (O_1302,N_26351,N_28231);
xnor UO_1303 (O_1303,N_25673,N_25610);
and UO_1304 (O_1304,N_29557,N_28680);
xnor UO_1305 (O_1305,N_25198,N_28708);
or UO_1306 (O_1306,N_25326,N_27736);
xnor UO_1307 (O_1307,N_29552,N_28863);
or UO_1308 (O_1308,N_26490,N_27229);
nand UO_1309 (O_1309,N_28905,N_26353);
nand UO_1310 (O_1310,N_25676,N_28528);
nor UO_1311 (O_1311,N_25023,N_29113);
or UO_1312 (O_1312,N_26387,N_25552);
and UO_1313 (O_1313,N_28006,N_25505);
and UO_1314 (O_1314,N_25085,N_29334);
nand UO_1315 (O_1315,N_26440,N_29263);
nor UO_1316 (O_1316,N_26820,N_27722);
nand UO_1317 (O_1317,N_26865,N_28861);
nor UO_1318 (O_1318,N_29928,N_28230);
and UO_1319 (O_1319,N_26733,N_29020);
or UO_1320 (O_1320,N_25816,N_25973);
nor UO_1321 (O_1321,N_29534,N_28188);
and UO_1322 (O_1322,N_28174,N_27260);
or UO_1323 (O_1323,N_29412,N_25079);
nor UO_1324 (O_1324,N_27320,N_28341);
nor UO_1325 (O_1325,N_25569,N_27492);
nor UO_1326 (O_1326,N_28148,N_27528);
xnor UO_1327 (O_1327,N_28816,N_28745);
nor UO_1328 (O_1328,N_29169,N_28166);
and UO_1329 (O_1329,N_29092,N_28904);
or UO_1330 (O_1330,N_27036,N_29915);
nor UO_1331 (O_1331,N_29916,N_28876);
nand UO_1332 (O_1332,N_29319,N_29172);
nor UO_1333 (O_1333,N_25856,N_29081);
nor UO_1334 (O_1334,N_26720,N_26305);
nor UO_1335 (O_1335,N_27569,N_28693);
or UO_1336 (O_1336,N_25405,N_29356);
or UO_1337 (O_1337,N_26116,N_25881);
and UO_1338 (O_1338,N_25665,N_26702);
and UO_1339 (O_1339,N_26093,N_27092);
and UO_1340 (O_1340,N_27711,N_28662);
nor UO_1341 (O_1341,N_28976,N_26645);
nand UO_1342 (O_1342,N_25832,N_26571);
or UO_1343 (O_1343,N_26700,N_27752);
or UO_1344 (O_1344,N_26325,N_26497);
nor UO_1345 (O_1345,N_27833,N_27767);
nand UO_1346 (O_1346,N_28918,N_29338);
or UO_1347 (O_1347,N_28519,N_27393);
or UO_1348 (O_1348,N_25325,N_25629);
or UO_1349 (O_1349,N_25406,N_25207);
xor UO_1350 (O_1350,N_26632,N_26561);
nand UO_1351 (O_1351,N_26294,N_26023);
or UO_1352 (O_1352,N_25764,N_26167);
or UO_1353 (O_1353,N_27148,N_28846);
nor UO_1354 (O_1354,N_26968,N_25981);
nor UO_1355 (O_1355,N_28320,N_28791);
xor UO_1356 (O_1356,N_26551,N_27929);
or UO_1357 (O_1357,N_27099,N_28652);
or UO_1358 (O_1358,N_25094,N_27708);
nor UO_1359 (O_1359,N_26502,N_25511);
nor UO_1360 (O_1360,N_28553,N_26158);
nand UO_1361 (O_1361,N_28094,N_29778);
or UO_1362 (O_1362,N_28332,N_29027);
nor UO_1363 (O_1363,N_25182,N_25600);
or UO_1364 (O_1364,N_27813,N_25641);
and UO_1365 (O_1365,N_25232,N_26203);
or UO_1366 (O_1366,N_26601,N_25368);
and UO_1367 (O_1367,N_29266,N_27991);
or UO_1368 (O_1368,N_28765,N_26462);
nor UO_1369 (O_1369,N_27710,N_25606);
or UO_1370 (O_1370,N_25655,N_25019);
and UO_1371 (O_1371,N_26656,N_29384);
nor UO_1372 (O_1372,N_28253,N_26536);
or UO_1373 (O_1373,N_28544,N_28562);
nor UO_1374 (O_1374,N_27780,N_29570);
or UO_1375 (O_1375,N_25783,N_28091);
or UO_1376 (O_1376,N_29709,N_25002);
nand UO_1377 (O_1377,N_26472,N_27038);
and UO_1378 (O_1378,N_25506,N_29981);
xor UO_1379 (O_1379,N_26290,N_28446);
and UO_1380 (O_1380,N_27989,N_26199);
or UO_1381 (O_1381,N_26019,N_27223);
nor UO_1382 (O_1382,N_26873,N_29487);
and UO_1383 (O_1383,N_25930,N_25598);
nor UO_1384 (O_1384,N_28702,N_29581);
nor UO_1385 (O_1385,N_25081,N_25849);
or UO_1386 (O_1386,N_28072,N_29731);
nand UO_1387 (O_1387,N_29277,N_29399);
or UO_1388 (O_1388,N_28950,N_25627);
nor UO_1389 (O_1389,N_26547,N_26906);
or UO_1390 (O_1390,N_27085,N_29165);
nand UO_1391 (O_1391,N_28269,N_28307);
and UO_1392 (O_1392,N_28154,N_27974);
or UO_1393 (O_1393,N_27098,N_26646);
and UO_1394 (O_1394,N_28385,N_26104);
xnor UO_1395 (O_1395,N_29588,N_26786);
or UO_1396 (O_1396,N_29862,N_28250);
nand UO_1397 (O_1397,N_28434,N_25423);
nand UO_1398 (O_1398,N_29200,N_28913);
or UO_1399 (O_1399,N_25621,N_27779);
or UO_1400 (O_1400,N_26989,N_26893);
and UO_1401 (O_1401,N_28466,N_29186);
nor UO_1402 (O_1402,N_27037,N_25276);
or UO_1403 (O_1403,N_27674,N_26833);
and UO_1404 (O_1404,N_26649,N_25028);
nor UO_1405 (O_1405,N_25358,N_29295);
or UO_1406 (O_1406,N_28506,N_26540);
and UO_1407 (O_1407,N_25267,N_28477);
and UO_1408 (O_1408,N_29901,N_25691);
nor UO_1409 (O_1409,N_25719,N_29402);
nor UO_1410 (O_1410,N_26028,N_27257);
nor UO_1411 (O_1411,N_26595,N_29071);
and UO_1412 (O_1412,N_25257,N_26839);
and UO_1413 (O_1413,N_29467,N_26881);
nand UO_1414 (O_1414,N_25664,N_29327);
xor UO_1415 (O_1415,N_25211,N_25443);
nand UO_1416 (O_1416,N_25593,N_29300);
or UO_1417 (O_1417,N_25860,N_27579);
or UO_1418 (O_1418,N_28498,N_26420);
nor UO_1419 (O_1419,N_25139,N_27132);
nor UO_1420 (O_1420,N_29710,N_26369);
and UO_1421 (O_1421,N_27396,N_25717);
nand UO_1422 (O_1422,N_29030,N_29101);
nand UO_1423 (O_1423,N_27693,N_25380);
or UO_1424 (O_1424,N_28633,N_26027);
or UO_1425 (O_1425,N_29155,N_28818);
nor UO_1426 (O_1426,N_28957,N_29111);
nor UO_1427 (O_1427,N_25293,N_26282);
nand UO_1428 (O_1428,N_25144,N_25696);
nand UO_1429 (O_1429,N_25509,N_27943);
and UO_1430 (O_1430,N_27486,N_28547);
nand UO_1431 (O_1431,N_27053,N_29427);
and UO_1432 (O_1432,N_25674,N_29644);
or UO_1433 (O_1433,N_29303,N_26136);
xnor UO_1434 (O_1434,N_25714,N_25975);
nand UO_1435 (O_1435,N_25092,N_26519);
nor UO_1436 (O_1436,N_29292,N_26036);
nand UO_1437 (O_1437,N_29742,N_27261);
or UO_1438 (O_1438,N_25912,N_29047);
nor UO_1439 (O_1439,N_29606,N_28966);
and UO_1440 (O_1440,N_27642,N_27631);
nor UO_1441 (O_1441,N_28678,N_25999);
nand UO_1442 (O_1442,N_27270,N_27062);
and UO_1443 (O_1443,N_29242,N_29767);
or UO_1444 (O_1444,N_26753,N_26939);
and UO_1445 (O_1445,N_29193,N_29472);
nand UO_1446 (O_1446,N_25485,N_27157);
or UO_1447 (O_1447,N_26975,N_27818);
nand UO_1448 (O_1448,N_27142,N_26564);
nor UO_1449 (O_1449,N_28114,N_29963);
and UO_1450 (O_1450,N_27278,N_25173);
and UO_1451 (O_1451,N_27897,N_27887);
or UO_1452 (O_1452,N_28262,N_26670);
or UO_1453 (O_1453,N_26297,N_27262);
nor UO_1454 (O_1454,N_26772,N_29985);
and UO_1455 (O_1455,N_28762,N_28425);
or UO_1456 (O_1456,N_29411,N_26442);
or UO_1457 (O_1457,N_26607,N_26430);
and UO_1458 (O_1458,N_25178,N_25360);
nand UO_1459 (O_1459,N_26012,N_25436);
nand UO_1460 (O_1460,N_27567,N_29496);
or UO_1461 (O_1461,N_26391,N_28438);
nand UO_1462 (O_1462,N_27442,N_25959);
nand UO_1463 (O_1463,N_29714,N_29234);
nor UO_1464 (O_1464,N_26074,N_28183);
and UO_1465 (O_1465,N_25845,N_27020);
nand UO_1466 (O_1466,N_26662,N_26594);
or UO_1467 (O_1467,N_26194,N_25013);
nand UO_1468 (O_1468,N_27912,N_28761);
and UO_1469 (O_1469,N_25463,N_25249);
nand UO_1470 (O_1470,N_28175,N_25863);
nor UO_1471 (O_1471,N_29687,N_26970);
and UO_1472 (O_1472,N_29022,N_25432);
xnor UO_1473 (O_1473,N_28031,N_29103);
xor UO_1474 (O_1474,N_29807,N_25892);
nand UO_1475 (O_1475,N_29146,N_27811);
nand UO_1476 (O_1476,N_25957,N_25540);
nand UO_1477 (O_1477,N_25980,N_27391);
and UO_1478 (O_1478,N_29878,N_27345);
xnor UO_1479 (O_1479,N_29199,N_25921);
nor UO_1480 (O_1480,N_29367,N_28486);
and UO_1481 (O_1481,N_28871,N_29846);
nor UO_1482 (O_1482,N_26085,N_26110);
and UO_1483 (O_1483,N_25901,N_27504);
xor UO_1484 (O_1484,N_26739,N_25914);
nor UO_1485 (O_1485,N_27054,N_26452);
and UO_1486 (O_1486,N_25571,N_27901);
and UO_1487 (O_1487,N_25268,N_28462);
nand UO_1488 (O_1488,N_28640,N_28358);
nand UO_1489 (O_1489,N_28170,N_26655);
nor UO_1490 (O_1490,N_25479,N_25372);
or UO_1491 (O_1491,N_25347,N_26221);
or UO_1492 (O_1492,N_27501,N_27363);
and UO_1493 (O_1493,N_29504,N_26360);
or UO_1494 (O_1494,N_28244,N_25045);
nand UO_1495 (O_1495,N_26777,N_26091);
nand UO_1496 (O_1496,N_27289,N_27401);
and UO_1497 (O_1497,N_26111,N_27556);
or UO_1498 (O_1498,N_25800,N_27973);
and UO_1499 (O_1499,N_26317,N_25188);
nor UO_1500 (O_1500,N_28637,N_28445);
nor UO_1501 (O_1501,N_26512,N_28699);
and UO_1502 (O_1502,N_29937,N_29673);
nand UO_1503 (O_1503,N_27522,N_28216);
xnor UO_1504 (O_1504,N_29806,N_28276);
nand UO_1505 (O_1505,N_28497,N_26835);
xnor UO_1506 (O_1506,N_28923,N_28710);
nand UO_1507 (O_1507,N_27392,N_28630);
and UO_1508 (O_1508,N_27950,N_25492);
and UO_1509 (O_1509,N_29021,N_28404);
or UO_1510 (O_1510,N_25809,N_26211);
or UO_1511 (O_1511,N_26926,N_26658);
xor UO_1512 (O_1512,N_26234,N_28058);
and UO_1513 (O_1513,N_29191,N_29238);
nand UO_1514 (O_1514,N_28636,N_26821);
nor UO_1515 (O_1515,N_29484,N_27911);
and UO_1516 (O_1516,N_25319,N_28026);
or UO_1517 (O_1517,N_29508,N_26013);
and UO_1518 (O_1518,N_26781,N_28771);
nand UO_1519 (O_1519,N_28472,N_29218);
nor UO_1520 (O_1520,N_29032,N_28302);
or UO_1521 (O_1521,N_26929,N_25725);
nand UO_1522 (O_1522,N_27806,N_27669);
and UO_1523 (O_1523,N_25135,N_25277);
nor UO_1524 (O_1524,N_26117,N_25898);
nand UO_1525 (O_1525,N_29996,N_25061);
nand UO_1526 (O_1526,N_28161,N_28127);
xor UO_1527 (O_1527,N_29790,N_28368);
or UO_1528 (O_1528,N_26458,N_28801);
nor UO_1529 (O_1529,N_26527,N_26948);
and UO_1530 (O_1530,N_29820,N_29390);
or UO_1531 (O_1531,N_28455,N_26907);
and UO_1532 (O_1532,N_29793,N_29142);
and UO_1533 (O_1533,N_28021,N_26788);
or UO_1534 (O_1534,N_28383,N_26228);
and UO_1535 (O_1535,N_25124,N_27683);
or UO_1536 (O_1536,N_28778,N_27217);
xor UO_1537 (O_1537,N_29825,N_27426);
and UO_1538 (O_1538,N_29594,N_25241);
xor UO_1539 (O_1539,N_27145,N_28852);
nand UO_1540 (O_1540,N_26920,N_28821);
nor UO_1541 (O_1541,N_28073,N_29728);
nand UO_1542 (O_1542,N_29610,N_29133);
or UO_1543 (O_1543,N_28482,N_27084);
or UO_1544 (O_1544,N_27757,N_26722);
and UO_1545 (O_1545,N_26778,N_29463);
nor UO_1546 (O_1546,N_28301,N_26585);
nor UO_1547 (O_1547,N_28085,N_28243);
nand UO_1548 (O_1548,N_27279,N_28113);
nor UO_1549 (O_1549,N_27039,N_26277);
nand UO_1550 (O_1550,N_28901,N_25906);
or UO_1551 (O_1551,N_29517,N_29007);
or UO_1552 (O_1552,N_26903,N_29328);
nor UO_1553 (O_1553,N_26344,N_28835);
and UO_1554 (O_1554,N_28779,N_26309);
and UO_1555 (O_1555,N_29194,N_29738);
nand UO_1556 (O_1556,N_28599,N_26470);
nand UO_1557 (O_1557,N_28014,N_27741);
xnor UO_1558 (O_1558,N_29420,N_27930);
or UO_1559 (O_1559,N_26130,N_27701);
and UO_1560 (O_1560,N_28606,N_26586);
nand UO_1561 (O_1561,N_27012,N_29320);
and UO_1562 (O_1562,N_25684,N_29258);
nand UO_1563 (O_1563,N_26427,N_27241);
nand UO_1564 (O_1564,N_25410,N_26405);
nand UO_1565 (O_1565,N_26800,N_28305);
xor UO_1566 (O_1566,N_26964,N_27726);
and UO_1567 (O_1567,N_25935,N_27871);
and UO_1568 (O_1568,N_26223,N_29676);
nand UO_1569 (O_1569,N_27064,N_26638);
xor UO_1570 (O_1570,N_25632,N_26463);
nor UO_1571 (O_1571,N_27878,N_26604);
and UO_1572 (O_1572,N_28926,N_27186);
and UO_1573 (O_1573,N_25777,N_27072);
nor UO_1574 (O_1574,N_29340,N_28264);
nor UO_1575 (O_1575,N_27686,N_27869);
and UO_1576 (O_1576,N_26569,N_29335);
and UO_1577 (O_1577,N_28560,N_28323);
nor UO_1578 (O_1578,N_26177,N_28289);
nor UO_1579 (O_1579,N_28480,N_28927);
nand UO_1580 (O_1580,N_28376,N_27707);
nand UO_1581 (O_1581,N_25175,N_25895);
or UO_1582 (O_1582,N_29196,N_28460);
nor UO_1583 (O_1583,N_28714,N_27542);
and UO_1584 (O_1584,N_27168,N_28974);
nand UO_1585 (O_1585,N_29114,N_28849);
or UO_1586 (O_1586,N_26813,N_25771);
and UO_1587 (O_1587,N_25659,N_25651);
or UO_1588 (O_1588,N_25403,N_28577);
and UO_1589 (O_1589,N_28690,N_26478);
and UO_1590 (O_1590,N_29291,N_28337);
and UO_1591 (O_1591,N_26192,N_26544);
or UO_1592 (O_1592,N_28649,N_28510);
nand UO_1593 (O_1593,N_27907,N_28359);
nor UO_1594 (O_1594,N_29992,N_29568);
nand UO_1595 (O_1595,N_27337,N_26332);
nor UO_1596 (O_1596,N_28430,N_28831);
and UO_1597 (O_1597,N_25909,N_27576);
and UO_1598 (O_1598,N_29822,N_26376);
nand UO_1599 (O_1599,N_26909,N_27836);
or UO_1600 (O_1600,N_27981,N_28665);
or UO_1601 (O_1601,N_27023,N_26454);
and UO_1602 (O_1602,N_28614,N_29577);
nor UO_1603 (O_1603,N_27423,N_29727);
nand UO_1604 (O_1604,N_29718,N_29000);
or UO_1605 (O_1605,N_29130,N_25123);
or UO_1606 (O_1606,N_28298,N_29720);
nand UO_1607 (O_1607,N_29744,N_29306);
and UO_1608 (O_1608,N_26365,N_25246);
or UO_1609 (O_1609,N_27520,N_26794);
nand UO_1610 (O_1610,N_28613,N_26692);
or UO_1611 (O_1611,N_25955,N_28008);
and UO_1612 (O_1612,N_28189,N_27889);
and UO_1613 (O_1613,N_28601,N_27713);
nand UO_1614 (O_1614,N_26118,N_27380);
nor UO_1615 (O_1615,N_26550,N_28691);
nand UO_1616 (O_1616,N_27774,N_27405);
nand UO_1617 (O_1617,N_26316,N_28595);
nand UO_1618 (O_1618,N_25177,N_26713);
nor UO_1619 (O_1619,N_28033,N_26746);
or UO_1620 (O_1620,N_29057,N_27033);
and UO_1621 (O_1621,N_26185,N_28668);
or UO_1622 (O_1622,N_26942,N_28643);
nor UO_1623 (O_1623,N_26400,N_26592);
or UO_1624 (O_1624,N_29313,N_25306);
nand UO_1625 (O_1625,N_27867,N_28592);
nor UO_1626 (O_1626,N_29946,N_27706);
xor UO_1627 (O_1627,N_28181,N_29120);
and UO_1628 (O_1628,N_25154,N_28236);
and UO_1629 (O_1629,N_28596,N_28529);
xor UO_1630 (O_1630,N_27959,N_28311);
nand UO_1631 (O_1631,N_29351,N_27017);
or UO_1632 (O_1632,N_26938,N_26847);
or UO_1633 (O_1633,N_27373,N_27886);
xnor UO_1634 (O_1634,N_26793,N_27185);
nand UO_1635 (O_1635,N_27518,N_28476);
nor UO_1636 (O_1636,N_27259,N_25759);
xnor UO_1637 (O_1637,N_27873,N_25352);
nor UO_1638 (O_1638,N_25862,N_25869);
xnor UO_1639 (O_1639,N_29375,N_27310);
or UO_1640 (O_1640,N_29771,N_29868);
nand UO_1641 (O_1641,N_26690,N_26054);
and UO_1642 (O_1642,N_26183,N_28624);
and UO_1643 (O_1643,N_27065,N_27738);
nand UO_1644 (O_1644,N_25698,N_25566);
xor UO_1645 (O_1645,N_26168,N_25424);
nor UO_1646 (O_1646,N_29932,N_27165);
nand UO_1647 (O_1647,N_26643,N_25538);
nand UO_1648 (O_1648,N_26468,N_26285);
and UO_1649 (O_1649,N_28800,N_26913);
nor UO_1650 (O_1650,N_26025,N_25947);
and UO_1651 (O_1651,N_25389,N_27558);
or UO_1652 (O_1652,N_25421,N_27008);
and UO_1653 (O_1653,N_26030,N_29509);
or UO_1654 (O_1654,N_27639,N_26026);
or UO_1655 (O_1655,N_29833,N_26523);
and UO_1656 (O_1656,N_25917,N_25381);
or UO_1657 (O_1657,N_29777,N_26555);
nand UO_1658 (O_1658,N_26072,N_28928);
or UO_1659 (O_1659,N_29814,N_27170);
nor UO_1660 (O_1660,N_26602,N_26483);
and UO_1661 (O_1661,N_28555,N_29818);
or UO_1662 (O_1662,N_27928,N_27496);
or UO_1663 (O_1663,N_26422,N_26273);
and UO_1664 (O_1664,N_29513,N_28057);
nor UO_1665 (O_1665,N_29859,N_28769);
nor UO_1666 (O_1666,N_29397,N_26301);
or UO_1667 (O_1667,N_25152,N_28764);
xnor UO_1668 (O_1668,N_29481,N_27860);
and UO_1669 (O_1669,N_27883,N_28187);
nor UO_1670 (O_1670,N_29748,N_29034);
nor UO_1671 (O_1671,N_28389,N_25155);
nor UO_1672 (O_1672,N_28671,N_27298);
nor UO_1673 (O_1673,N_27688,N_26303);
and UO_1674 (O_1674,N_25230,N_28279);
and UO_1675 (O_1675,N_25470,N_28479);
xor UO_1676 (O_1676,N_27378,N_29752);
nand UO_1677 (O_1677,N_28303,N_25586);
nor UO_1678 (O_1678,N_29437,N_27538);
and UO_1679 (O_1679,N_27953,N_29921);
nand UO_1680 (O_1680,N_27290,N_29345);
nor UO_1681 (O_1681,N_27814,N_27334);
and UO_1682 (O_1682,N_27747,N_29434);
nor UO_1683 (O_1683,N_27083,N_28903);
nor UO_1684 (O_1684,N_29665,N_28774);
nand UO_1685 (O_1685,N_26830,N_26380);
or UO_1686 (O_1686,N_25176,N_25099);
xnor UO_1687 (O_1687,N_25467,N_26993);
and UO_1688 (O_1688,N_29176,N_25196);
xor UO_1689 (O_1689,N_26487,N_29308);
and UO_1690 (O_1690,N_29124,N_26848);
nand UO_1691 (O_1691,N_25468,N_26245);
nor UO_1692 (O_1692,N_27108,N_27986);
nor UO_1693 (O_1693,N_29158,N_25590);
and UO_1694 (O_1694,N_29618,N_26368);
nand UO_1695 (O_1695,N_27411,N_29965);
nor UO_1696 (O_1696,N_26969,N_26007);
nor UO_1697 (O_1697,N_29289,N_25653);
and UO_1698 (O_1698,N_25035,N_25843);
nor UO_1699 (O_1699,N_29940,N_25603);
or UO_1700 (O_1700,N_25180,N_29736);
or UO_1701 (O_1701,N_27562,N_28938);
nor UO_1702 (O_1702,N_29501,N_26047);
nor UO_1703 (O_1703,N_29268,N_28574);
and UO_1704 (O_1704,N_25802,N_28222);
nand UO_1705 (O_1705,N_25715,N_29051);
nor UO_1706 (O_1706,N_26103,N_29876);
or UO_1707 (O_1707,N_29990,N_26437);
nor UO_1708 (O_1708,N_27982,N_25286);
and UO_1709 (O_1709,N_25965,N_25817);
nand UO_1710 (O_1710,N_25051,N_26267);
nor UO_1711 (O_1711,N_28682,N_27895);
and UO_1712 (O_1712,N_26890,N_28449);
nand UO_1713 (O_1713,N_25243,N_27460);
and UO_1714 (O_1714,N_27628,N_29093);
or UO_1715 (O_1715,N_29332,N_25273);
nor UO_1716 (O_1716,N_25650,N_29626);
nand UO_1717 (O_1717,N_29376,N_25310);
nand UO_1718 (O_1718,N_26435,N_28280);
nor UO_1719 (O_1719,N_27737,N_29693);
and UO_1720 (O_1720,N_28796,N_25285);
and UO_1721 (O_1721,N_27446,N_25116);
nand UO_1722 (O_1722,N_29348,N_29700);
or UO_1723 (O_1723,N_27018,N_27103);
and UO_1724 (O_1724,N_25502,N_26630);
nand UO_1725 (O_1725,N_25568,N_29239);
nand UO_1726 (O_1726,N_29970,N_27182);
or UO_1727 (O_1727,N_29934,N_26883);
xor UO_1728 (O_1728,N_29974,N_25420);
and UO_1729 (O_1729,N_27885,N_28912);
nor UO_1730 (O_1730,N_25808,N_28999);
nand UO_1731 (O_1731,N_26689,N_27842);
or UO_1732 (O_1732,N_27385,N_29865);
nand UO_1733 (O_1733,N_26480,N_29542);
nor UO_1734 (O_1734,N_29891,N_28907);
xor UO_1735 (O_1735,N_28504,N_25083);
and UO_1736 (O_1736,N_29459,N_29861);
nor UO_1737 (O_1737,N_29518,N_27835);
and UO_1738 (O_1738,N_28288,N_27531);
nor UO_1739 (O_1739,N_28176,N_29465);
or UO_1740 (O_1740,N_25560,N_29759);
and UO_1741 (O_1741,N_27090,N_26599);
nor UO_1742 (O_1742,N_25466,N_26568);
and UO_1743 (O_1743,N_29706,N_29370);
nand UO_1744 (O_1744,N_25654,N_26988);
xnor UO_1745 (O_1745,N_28249,N_26694);
nor UO_1746 (O_1746,N_25156,N_28284);
nor UO_1747 (O_1747,N_28268,N_29107);
or UO_1748 (O_1748,N_28525,N_27754);
or UO_1749 (O_1749,N_27920,N_29905);
nand UO_1750 (O_1750,N_27899,N_29490);
or UO_1751 (O_1751,N_26754,N_28712);
and UO_1752 (O_1752,N_27574,N_29079);
or UO_1753 (O_1753,N_26864,N_27888);
or UO_1754 (O_1754,N_27644,N_26750);
nand UO_1755 (O_1755,N_26021,N_29949);
xor UO_1756 (O_1756,N_27029,N_29406);
nor UO_1757 (O_1757,N_25012,N_26593);
and UO_1758 (O_1758,N_27679,N_28372);
nand UO_1759 (O_1759,N_27061,N_27586);
and UO_1760 (O_1760,N_28300,N_27440);
and UO_1761 (O_1761,N_25628,N_25385);
or UO_1762 (O_1762,N_27078,N_29926);
or UO_1763 (O_1763,N_26186,N_28798);
nor UO_1764 (O_1764,N_25658,N_29888);
nand UO_1765 (O_1765,N_28297,N_25836);
or UO_1766 (O_1766,N_27206,N_25168);
nand UO_1767 (O_1767,N_26154,N_25386);
nand UO_1768 (O_1768,N_27394,N_27156);
and UO_1769 (O_1769,N_27275,N_25097);
and UO_1770 (O_1770,N_26445,N_29539);
and UO_1771 (O_1771,N_27482,N_26197);
or UO_1772 (O_1772,N_25040,N_25383);
and UO_1773 (O_1773,N_25348,N_27605);
and UO_1774 (O_1774,N_28295,N_28347);
and UO_1775 (O_1775,N_29018,N_28829);
nor UO_1776 (O_1776,N_27690,N_26133);
nor UO_1777 (O_1777,N_26095,N_25577);
nand UO_1778 (O_1778,N_28369,N_28141);
nand UO_1779 (O_1779,N_28890,N_26235);
xnor UO_1780 (O_1780,N_29747,N_28517);
nor UO_1781 (O_1781,N_25594,N_26269);
or UO_1782 (O_1782,N_29153,N_25539);
nand UO_1783 (O_1783,N_29553,N_29042);
and UO_1784 (O_1784,N_26231,N_25998);
or UO_1785 (O_1785,N_25038,N_27368);
or UO_1786 (O_1786,N_27794,N_29894);
xnor UO_1787 (O_1787,N_26213,N_27450);
nor UO_1788 (O_1788,N_29209,N_27941);
xor UO_1789 (O_1789,N_27224,N_26163);
or UO_1790 (O_1790,N_26767,N_25848);
and UO_1791 (O_1791,N_29017,N_26654);
or UO_1792 (O_1792,N_29520,N_25242);
nor UO_1793 (O_1793,N_26202,N_26122);
nand UO_1794 (O_1794,N_28168,N_28569);
nand UO_1795 (O_1795,N_28836,N_27301);
nor UO_1796 (O_1796,N_29210,N_25737);
xnor UO_1797 (O_1797,N_27495,N_28793);
xor UO_1798 (O_1798,N_28792,N_27312);
or UO_1799 (O_1799,N_28556,N_26747);
nand UO_1800 (O_1800,N_29717,N_27681);
nand UO_1801 (O_1801,N_29359,N_27383);
xnor UO_1802 (O_1802,N_28981,N_28615);
and UO_1803 (O_1803,N_27789,N_28908);
and UO_1804 (O_1804,N_28223,N_25815);
nand UO_1805 (O_1805,N_26524,N_25708);
xnor UO_1806 (O_1806,N_29149,N_25248);
nand UO_1807 (O_1807,N_26665,N_25342);
or UO_1808 (O_1808,N_28047,N_29097);
nand UO_1809 (O_1809,N_27281,N_26933);
and UO_1810 (O_1810,N_29680,N_27606);
or UO_1811 (O_1811,N_27180,N_28597);
nand UO_1812 (O_1812,N_28003,N_26878);
or UO_1813 (O_1813,N_25404,N_28619);
nand UO_1814 (O_1814,N_28719,N_29118);
nand UO_1815 (O_1815,N_26414,N_29059);
and UO_1816 (O_1816,N_27221,N_25864);
nand UO_1817 (O_1817,N_25855,N_25962);
nand UO_1818 (O_1818,N_27233,N_29947);
and UO_1819 (O_1819,N_25272,N_26399);
and UO_1820 (O_1820,N_27287,N_26324);
nor UO_1821 (O_1821,N_27826,N_26291);
xnor UO_1822 (O_1822,N_27595,N_29850);
nand UO_1823 (O_1823,N_29911,N_26310);
nor UO_1824 (O_1824,N_27138,N_27467);
nor UO_1825 (O_1825,N_27875,N_29183);
and UO_1826 (O_1826,N_28377,N_29563);
nor UO_1827 (O_1827,N_25823,N_26625);
or UO_1828 (O_1828,N_26460,N_28993);
or UO_1829 (O_1829,N_27231,N_27114);
nor UO_1830 (O_1830,N_25336,N_28144);
nor UO_1831 (O_1831,N_26808,N_29975);
and UO_1832 (O_1832,N_26080,N_27166);
and UO_1833 (O_1833,N_28384,N_25197);
nand UO_1834 (O_1834,N_26732,N_26075);
nand UO_1835 (O_1835,N_27510,N_26326);
nand UO_1836 (O_1836,N_26384,N_25299);
nor UO_1837 (O_1837,N_25736,N_28469);
nand UO_1838 (O_1838,N_27388,N_25004);
nor UO_1839 (O_1839,N_28667,N_29446);
nor UO_1840 (O_1840,N_27264,N_29009);
or UO_1841 (O_1841,N_26620,N_26832);
or UO_1842 (O_1842,N_26553,N_28147);
or UO_1843 (O_1843,N_25794,N_25622);
xnor UO_1844 (O_1844,N_25780,N_28878);
and UO_1845 (O_1845,N_26307,N_27057);
nor UO_1846 (O_1846,N_28848,N_25090);
nand UO_1847 (O_1847,N_26761,N_25333);
nand UO_1848 (O_1848,N_25657,N_25195);
nor UO_1849 (O_1849,N_25281,N_25804);
and UO_1850 (O_1850,N_28650,N_29012);
xor UO_1851 (O_1851,N_26142,N_26298);
xor UO_1852 (O_1852,N_29855,N_28830);
and UO_1853 (O_1853,N_25866,N_28432);
nor UO_1854 (O_1854,N_26443,N_25739);
nand UO_1855 (O_1855,N_26570,N_29995);
xnor UO_1856 (O_1856,N_27109,N_29920);
or UO_1857 (O_1857,N_26682,N_25417);
or UO_1858 (O_1858,N_26741,N_26836);
and UO_1859 (O_1859,N_25416,N_29422);
and UO_1860 (O_1860,N_28576,N_25619);
nand UO_1861 (O_1861,N_28429,N_28240);
or UO_1862 (O_1862,N_29252,N_29439);
and UO_1863 (O_1863,N_28899,N_28967);
nor UO_1864 (O_1864,N_25584,N_25337);
and UO_1865 (O_1865,N_28789,N_26611);
or UO_1866 (O_1866,N_25812,N_26717);
and UO_1867 (O_1867,N_25744,N_26140);
nand UO_1868 (O_1868,N_28964,N_26274);
xor UO_1869 (O_1869,N_28213,N_27524);
nor UO_1870 (O_1870,N_26209,N_26596);
or UO_1871 (O_1871,N_29363,N_25430);
or UO_1872 (O_1872,N_25356,N_26153);
nand UO_1873 (O_1873,N_27798,N_26097);
or UO_1874 (O_1874,N_27976,N_26126);
xor UO_1875 (O_1875,N_27861,N_29424);
nor UO_1876 (O_1876,N_27675,N_27465);
nand UO_1877 (O_1877,N_25920,N_27742);
nand UO_1878 (O_1878,N_25205,N_28887);
and UO_1879 (O_1879,N_25875,N_25562);
or UO_1880 (O_1880,N_29616,N_26807);
xnor UO_1881 (O_1881,N_28963,N_25903);
nand UO_1882 (O_1882,N_27613,N_25946);
nor UO_1883 (O_1883,N_25001,N_28683);
nand UO_1884 (O_1884,N_28943,N_26627);
nor UO_1885 (O_1885,N_25838,N_25512);
nand UO_1886 (O_1886,N_25490,N_28994);
nand UO_1887 (O_1887,N_28068,N_25967);
nand UO_1888 (O_1888,N_29023,N_25411);
and UO_1889 (O_1889,N_26758,N_25515);
or UO_1890 (O_1890,N_28197,N_27247);
nand UO_1891 (O_1891,N_28387,N_28937);
or UO_1892 (O_1892,N_25387,N_27615);
nor UO_1893 (O_1893,N_27021,N_26979);
and UO_1894 (O_1894,N_25861,N_27243);
or UO_1895 (O_1895,N_28512,N_28605);
or UO_1896 (O_1896,N_26379,N_27413);
nand UO_1897 (O_1897,N_27284,N_25465);
and UO_1898 (O_1898,N_27666,N_28410);
nand UO_1899 (O_1899,N_25660,N_28278);
xor UO_1900 (O_1900,N_29845,N_27533);
or UO_1901 (O_1901,N_27149,N_29395);
nor UO_1902 (O_1902,N_26287,N_25775);
nor UO_1903 (O_1903,N_27698,N_25036);
nor UO_1904 (O_1904,N_28207,N_29584);
or UO_1905 (O_1905,N_29478,N_29469);
and UO_1906 (O_1906,N_26499,N_25773);
and UO_1907 (O_1907,N_25952,N_25943);
nor UO_1908 (O_1908,N_27505,N_29257);
nand UO_1909 (O_1909,N_28707,N_26954);
and UO_1910 (O_1910,N_28891,N_27582);
nand UO_1911 (O_1911,N_25145,N_28658);
nand UO_1912 (O_1912,N_25219,N_29470);
nand UO_1913 (O_1913,N_28324,N_27110);
nor UO_1914 (O_1914,N_29519,N_25617);
nor UO_1915 (O_1915,N_25542,N_29548);
or UO_1916 (O_1916,N_27232,N_26763);
and UO_1917 (O_1917,N_27341,N_26471);
nand UO_1918 (O_1918,N_27877,N_29766);
or UO_1919 (O_1919,N_26724,N_28378);
nor UO_1920 (O_1920,N_28019,N_26867);
and UO_1921 (O_1921,N_28350,N_26393);
nand UO_1922 (O_1922,N_27164,N_25556);
nor UO_1923 (O_1923,N_25870,N_27667);
nand UO_1924 (O_1924,N_28426,N_26271);
or UO_1925 (O_1925,N_28958,N_28229);
and UO_1926 (O_1926,N_29797,N_26609);
and UO_1927 (O_1927,N_29495,N_27215);
nor UO_1928 (O_1928,N_26695,N_29449);
or UO_1929 (O_1929,N_27478,N_28025);
nand UO_1930 (O_1930,N_26306,N_28461);
xnor UO_1931 (O_1931,N_29350,N_29589);
or UO_1932 (O_1932,N_25756,N_25315);
nand UO_1933 (O_1933,N_25648,N_29203);
and UO_1934 (O_1934,N_27074,N_28447);
nand UO_1935 (O_1935,N_27627,N_27113);
nand UO_1936 (O_1936,N_26436,N_29897);
and UO_1937 (O_1937,N_28227,N_25226);
and UO_1938 (O_1938,N_25361,N_28367);
xnor UO_1939 (O_1939,N_25695,N_29247);
and UO_1940 (O_1940,N_26390,N_26634);
nor UO_1941 (O_1941,N_28853,N_25948);
or UO_1942 (O_1942,N_28103,N_27425);
nand UO_1943 (O_1943,N_28984,N_28217);
and UO_1944 (O_1944,N_28186,N_25026);
or UO_1945 (O_1945,N_25126,N_25572);
and UO_1946 (O_1946,N_27591,N_28696);
nand UO_1947 (O_1947,N_25630,N_27782);
and UO_1948 (O_1948,N_29675,N_27321);
nor UO_1949 (O_1949,N_27597,N_28568);
nand UO_1950 (O_1950,N_29426,N_26577);
nand UO_1951 (O_1951,N_27997,N_28627);
or UO_1952 (O_1952,N_27313,N_25537);
nor UO_1953 (O_1953,N_26461,N_27760);
and UO_1954 (O_1954,N_29374,N_29784);
or UO_1955 (O_1955,N_27263,N_25726);
or UO_1956 (O_1956,N_25899,N_27336);
or UO_1957 (O_1957,N_29123,N_26106);
nor UO_1958 (O_1958,N_28314,N_25883);
nand UO_1959 (O_1959,N_29010,N_27718);
and UO_1960 (O_1960,N_26918,N_27362);
and UO_1961 (O_1961,N_29296,N_27566);
and UO_1962 (O_1962,N_29482,N_26908);
and UO_1963 (O_1963,N_27418,N_26238);
or UO_1964 (O_1964,N_25904,N_28043);
nor UO_1965 (O_1965,N_29603,N_25807);
or UO_1966 (O_1966,N_25558,N_26171);
xor UO_1967 (O_1967,N_25699,N_26359);
and UO_1968 (O_1968,N_29871,N_28810);
or UO_1969 (O_1969,N_27153,N_29582);
or UO_1970 (O_1970,N_27532,N_27641);
nor UO_1971 (O_1971,N_26612,N_29642);
and UO_1972 (O_1972,N_26849,N_29956);
xnor UO_1973 (O_1973,N_29403,N_29276);
and UO_1974 (O_1974,N_27379,N_28648);
and UO_1975 (O_1975,N_27022,N_29489);
nor UO_1976 (O_1976,N_29480,N_29115);
nor UO_1977 (O_1977,N_28589,N_25171);
nor UO_1978 (O_1978,N_25893,N_28135);
nand UO_1979 (O_1979,N_29054,N_29273);
nand UO_1980 (O_1980,N_25916,N_27966);
and UO_1981 (O_1981,N_29527,N_29096);
and UO_1982 (O_1982,N_29261,N_28062);
or UO_1983 (O_1983,N_27342,N_25437);
and UO_1984 (O_1984,N_29100,N_26622);
xnor UO_1985 (O_1985,N_28309,N_28401);
or UO_1986 (O_1986,N_26438,N_27491);
nand UO_1987 (O_1987,N_29400,N_27565);
and UO_1988 (O_1988,N_25331,N_27121);
or UO_1989 (O_1989,N_25339,N_28898);
nand UO_1990 (O_1990,N_26900,N_26990);
nor UO_1991 (O_1991,N_29324,N_26860);
or UO_1992 (O_1992,N_29450,N_27781);
or UO_1993 (O_1993,N_25350,N_27519);
or UO_1994 (O_1994,N_28146,N_28343);
or UO_1995 (O_1995,N_29617,N_29782);
and UO_1996 (O_1996,N_27052,N_27670);
or UO_1997 (O_1997,N_29964,N_26148);
xnor UO_1998 (O_1998,N_28573,N_26543);
xor UO_1999 (O_1999,N_25678,N_26366);
nand UO_2000 (O_2000,N_29740,N_26389);
and UO_2001 (O_2001,N_28617,N_27479);
nand UO_2002 (O_2002,N_28788,N_25640);
nor UO_2003 (O_2003,N_28679,N_28265);
and UO_2004 (O_2004,N_27266,N_28579);
nand UO_2005 (O_2005,N_26321,N_27601);
or UO_2006 (O_2006,N_29541,N_28294);
nand UO_2007 (O_2007,N_25536,N_27249);
and UO_2008 (O_2008,N_29080,N_28960);
nor UO_2009 (O_2009,N_28750,N_29160);
nor UO_2010 (O_2010,N_29048,N_26981);
nor UO_2011 (O_2011,N_28731,N_27464);
or UO_2012 (O_2012,N_26618,N_29003);
xnor UO_2013 (O_2013,N_29658,N_28360);
xor UO_2014 (O_2014,N_29801,N_29816);
and UO_2015 (O_2015,N_27841,N_25846);
or UO_2016 (O_2016,N_28612,N_27553);
nor UO_2017 (O_2017,N_28948,N_26520);
nor UO_2018 (O_2018,N_28936,N_29380);
or UO_2019 (O_2019,N_25103,N_29498);
nor UO_2020 (O_2020,N_26574,N_28546);
xnor UO_2021 (O_2021,N_25680,N_25050);
or UO_2022 (O_2022,N_27445,N_28339);
and UO_2023 (O_2023,N_28838,N_27288);
or UO_2024 (O_2024,N_26851,N_26715);
nor UO_2025 (O_2025,N_28537,N_26877);
nor UO_2026 (O_2026,N_29215,N_27451);
and UO_2027 (O_2027,N_27734,N_28670);
or UO_2028 (O_2028,N_25546,N_26208);
xor UO_2029 (O_2029,N_28695,N_29663);
nand UO_2030 (O_2030,N_27663,N_25231);
nand UO_2031 (O_2031,N_27636,N_28542);
nand UO_2032 (O_2032,N_27799,N_29647);
and UO_2033 (O_2033,N_27507,N_28832);
nor UO_2034 (O_2034,N_27471,N_28909);
nand UO_2035 (O_2035,N_26035,N_25643);
nand UO_2036 (O_2036,N_27323,N_25498);
nor UO_2037 (O_2037,N_25936,N_28143);
nor UO_2038 (O_2038,N_25963,N_26382);
or UO_2039 (O_2039,N_29571,N_27003);
nand UO_2040 (O_2040,N_25500,N_29314);
and UO_2041 (O_2041,N_27955,N_25375);
nand UO_2042 (O_2042,N_28403,N_28567);
or UO_2043 (O_2043,N_25440,N_26352);
and UO_2044 (O_2044,N_27001,N_29691);
nand UO_2045 (O_2045,N_25743,N_26776);
or UO_2046 (O_2046,N_27139,N_27444);
and UO_2047 (O_2047,N_29973,N_26518);
nand UO_2048 (O_2048,N_26375,N_26230);
and UO_2049 (O_2049,N_27030,N_27640);
nor UO_2050 (O_2050,N_28194,N_27964);
nor UO_2051 (O_2051,N_25290,N_25208);
and UO_2052 (O_2052,N_25786,N_27269);
nor UO_2053 (O_2053,N_28864,N_28082);
xor UO_2054 (O_2054,N_27454,N_27513);
nand UO_2055 (O_2055,N_27800,N_29109);
nor UO_2056 (O_2056,N_27891,N_28543);
or UO_2057 (O_2057,N_27080,N_29127);
and UO_2058 (O_2058,N_27691,N_29373);
nor UO_2059 (O_2059,N_28059,N_28833);
or UO_2060 (O_2060,N_29065,N_26121);
nand UO_2061 (O_2061,N_28956,N_27207);
nor UO_2062 (O_2062,N_29774,N_27135);
nand UO_2063 (O_2063,N_25279,N_28689);
or UO_2064 (O_2064,N_28503,N_28052);
nor UO_2065 (O_2065,N_26333,N_27516);
nand UO_2066 (O_2066,N_28646,N_29250);
and UO_2067 (O_2067,N_27740,N_28172);
nand UO_2068 (O_2068,N_27234,N_27617);
and UO_2069 (O_2069,N_27960,N_26491);
nor UO_2070 (O_2070,N_25037,N_28939);
nor UO_2071 (O_2071,N_28681,N_27349);
or UO_2072 (O_2072,N_28069,N_27620);
and UO_2073 (O_2073,N_29364,N_29565);
nor UO_2074 (O_2074,N_27076,N_29978);
or UO_2075 (O_2075,N_28335,N_28415);
xor UO_2076 (O_2076,N_27680,N_28638);
and UO_2077 (O_2077,N_29002,N_27854);
nand UO_2078 (O_2078,N_28386,N_27653);
and UO_2079 (O_2079,N_27213,N_28902);
and UO_2080 (O_2080,N_26600,N_27657);
or UO_2081 (O_2081,N_29674,N_29682);
and UO_2082 (O_2082,N_27333,N_25138);
nor UO_2083 (O_2083,N_29279,N_27541);
and UO_2084 (O_2084,N_26734,N_25200);
xor UO_2085 (O_2085,N_25435,N_29039);
nor UO_2086 (O_2086,N_26657,N_28894);
nand UO_2087 (O_2087,N_29037,N_29507);
nor UO_2088 (O_2088,N_26492,N_26339);
or UO_2089 (O_2089,N_29907,N_25557);
nand UO_2090 (O_2090,N_27603,N_29228);
and UO_2091 (O_2091,N_29473,N_28357);
or UO_2092 (O_2092,N_25785,N_25450);
and UO_2093 (O_2093,N_29503,N_28961);
nor UO_2094 (O_2094,N_26043,N_29944);
nand UO_2095 (O_2095,N_26897,N_29462);
nor UO_2096 (O_2096,N_27952,N_26509);
and UO_2097 (O_2097,N_27079,N_26178);
xor UO_2098 (O_2098,N_26206,N_25140);
xor UO_2099 (O_2099,N_27812,N_29620);
xnor UO_2100 (O_2100,N_27677,N_26284);
nor UO_2101 (O_2101,N_26288,N_29448);
and UO_2102 (O_2102,N_27797,N_27659);
nand UO_2103 (O_2103,N_26541,N_27821);
nor UO_2104 (O_2104,N_29293,N_27081);
nand UO_2105 (O_2105,N_26752,N_26371);
nor UO_2106 (O_2106,N_28200,N_29134);
nor UO_2107 (O_2107,N_26469,N_26823);
nand UO_2108 (O_2108,N_28046,N_29660);
and UO_2109 (O_2109,N_26798,N_28703);
nor UO_2110 (O_2110,N_26246,N_28272);
xnor UO_2111 (O_2111,N_28677,N_28884);
or UO_2112 (O_2112,N_27343,N_28772);
xnor UO_2113 (O_2113,N_26184,N_27984);
nand UO_2114 (O_2114,N_29253,N_25067);
nand UO_2115 (O_2115,N_26506,N_29237);
and UO_2116 (O_2116,N_29815,N_29207);
and UO_2117 (O_2117,N_27056,N_29538);
nor UO_2118 (O_2118,N_26522,N_28985);
or UO_2119 (O_2119,N_28749,N_29368);
or UO_2120 (O_2120,N_28060,N_29401);
nand UO_2121 (O_2121,N_26064,N_29961);
or UO_2122 (O_2122,N_27969,N_26635);
nor UO_2123 (O_2123,N_26331,N_28759);
or UO_2124 (O_2124,N_26950,N_25264);
nor UO_2125 (O_2125,N_28755,N_27309);
nand UO_2126 (O_2126,N_26342,N_25635);
xor UO_2127 (O_2127,N_28825,N_27719);
nor UO_2128 (O_2128,N_25681,N_26378);
and UO_2129 (O_2129,N_25136,N_26691);
nand UO_2130 (O_2130,N_26817,N_29734);
nand UO_2131 (O_2131,N_27848,N_26894);
or UO_2132 (O_2132,N_27455,N_27490);
and UO_2133 (O_2133,N_27857,N_27356);
and UO_2134 (O_2134,N_25237,N_28859);
or UO_2135 (O_2135,N_26977,N_26477);
nor UO_2136 (O_2136,N_25018,N_25327);
or UO_2137 (O_2137,N_27946,N_25939);
nand UO_2138 (O_2138,N_28775,N_27902);
nor UO_2139 (O_2139,N_28986,N_28475);
and UO_2140 (O_2140,N_25841,N_27998);
or UO_2141 (O_2141,N_28488,N_28039);
nand UO_2142 (O_2142,N_27850,N_29341);
and UO_2143 (O_2143,N_26314,N_27188);
nand UO_2144 (O_2144,N_25508,N_27441);
nor UO_2145 (O_2145,N_29028,N_25428);
nor UO_2146 (O_2146,N_28077,N_29383);
nand UO_2147 (O_2147,N_26358,N_26149);
nand UO_2148 (O_2148,N_28394,N_29812);
nand UO_2149 (O_2149,N_26787,N_29108);
and UO_2150 (O_2150,N_25596,N_29145);
nor UO_2151 (O_2151,N_25220,N_29188);
and UO_2152 (O_2152,N_29741,N_27258);
or UO_2153 (O_2153,N_29164,N_27822);
and UO_2154 (O_2154,N_25434,N_25803);
and UO_2155 (O_2155,N_28794,N_27043);
nand UO_2156 (O_2156,N_27494,N_29540);
and UO_2157 (O_2157,N_25668,N_26302);
xor UO_2158 (O_2158,N_28875,N_28706);
nand UO_2159 (O_2159,N_29391,N_27497);
nor UO_2160 (O_2160,N_29558,N_25842);
nor UO_2161 (O_2161,N_27987,N_28454);
nand UO_2162 (O_2162,N_26931,N_27633);
nand UO_2163 (O_2163,N_27900,N_25185);
nand UO_2164 (O_2164,N_29154,N_29045);
nor UO_2165 (O_2165,N_25374,N_27073);
nand UO_2166 (O_2166,N_28220,N_27047);
or UO_2167 (O_2167,N_25822,N_26127);
or UO_2168 (O_2168,N_27280,N_25427);
or UO_2169 (O_2169,N_27319,N_27803);
nand UO_2170 (O_2170,N_25218,N_26584);
xnor UO_2171 (O_2171,N_26745,N_28916);
and UO_2172 (O_2172,N_29511,N_27285);
and UO_2173 (O_2173,N_28593,N_28208);
or UO_2174 (O_2174,N_25151,N_29284);
and UO_2175 (O_2175,N_29765,N_26614);
and UO_2176 (O_2176,N_27255,N_27529);
nand UO_2177 (O_2177,N_27050,N_29220);
and UO_2178 (O_2178,N_27141,N_27240);
nand UO_2179 (O_2179,N_25460,N_27840);
and UO_2180 (O_2180,N_25288,N_25157);
or UO_2181 (O_2181,N_27005,N_25754);
nor UO_2182 (O_2182,N_26403,N_25991);
nor UO_2183 (O_2183,N_25510,N_25795);
nand UO_2184 (O_2184,N_29791,N_27851);
and UO_2185 (O_2185,N_25187,N_26680);
and UO_2186 (O_2186,N_28257,N_27346);
and UO_2187 (O_2187,N_27935,N_27554);
nor UO_2188 (O_2188,N_25748,N_25255);
and UO_2189 (O_2189,N_25772,N_25616);
nand UO_2190 (O_2190,N_27449,N_27173);
xor UO_2191 (O_2191,N_27619,N_26650);
nor UO_2192 (O_2192,N_28822,N_29838);
or UO_2193 (O_2193,N_27429,N_29800);
or UO_2194 (O_2194,N_25503,N_29404);
nand UO_2195 (O_2195,N_29713,N_28725);
nor UO_2196 (O_2196,N_29522,N_29179);
and UO_2197 (O_2197,N_28502,N_29178);
xor UO_2198 (O_2198,N_27377,N_29787);
and UO_2199 (O_2199,N_25685,N_29698);
or UO_2200 (O_2200,N_28812,N_27523);
nor UO_2201 (O_2201,N_29147,N_25114);
xor UO_2202 (O_2202,N_27931,N_25894);
and UO_2203 (O_2203,N_27563,N_29116);
xnor UO_2204 (O_2204,N_25300,N_28639);
and UO_2205 (O_2205,N_27331,N_27804);
xor UO_2206 (O_2206,N_29809,N_29811);
nor UO_2207 (O_2207,N_28282,N_28934);
nand UO_2208 (O_2208,N_26137,N_27406);
and UO_2209 (O_2209,N_29128,N_26774);
and UO_2210 (O_2210,N_27296,N_27097);
and UO_2211 (O_2211,N_25988,N_27853);
nor UO_2212 (O_2212,N_28754,N_29205);
nor UO_2213 (O_2213,N_29358,N_26079);
and UO_2214 (O_2214,N_29302,N_28982);
or UO_2215 (O_2215,N_27216,N_26613);
and UO_2216 (O_2216,N_28001,N_25251);
or UO_2217 (O_2217,N_26446,N_25132);
xnor UO_2218 (O_2218,N_26721,N_28202);
or UO_2219 (O_2219,N_29699,N_29612);
or UO_2220 (O_2220,N_29866,N_25189);
or UO_2221 (O_2221,N_27242,N_29895);
nand UO_2222 (O_2222,N_28873,N_26134);
or UO_2223 (O_2223,N_27208,N_25700);
nand UO_2224 (O_2224,N_29544,N_25245);
nor UO_2225 (O_2225,N_29516,N_28163);
xnor UO_2226 (O_2226,N_26089,N_25897);
nand UO_2227 (O_2227,N_28588,N_25455);
nor UO_2228 (O_2228,N_29725,N_26151);
xor UO_2229 (O_2229,N_28672,N_28090);
nor UO_2230 (O_2230,N_28416,N_29769);
and UO_2231 (O_2231,N_25626,N_28697);
nor UO_2232 (O_2232,N_26252,N_28700);
nor UO_2233 (O_2233,N_27580,N_27273);
xnor UO_2234 (O_2234,N_29287,N_29984);
and UO_2235 (O_2235,N_29206,N_29074);
nand UO_2236 (O_2236,N_28549,N_29933);
or UO_2237 (O_2237,N_26320,N_27934);
nand UO_2238 (O_2238,N_28521,N_29564);
nand UO_2239 (O_2239,N_28987,N_25787);
nand UO_2240 (O_2240,N_28018,N_29646);
nor UO_2241 (O_2241,N_27589,N_25160);
and UO_2242 (O_2242,N_29421,N_26818);
or UO_2243 (O_2243,N_29514,N_25774);
nor UO_2244 (O_2244,N_27748,N_27914);
xor UO_2245 (O_2245,N_29954,N_28962);
nand UO_2246 (O_2246,N_29014,N_25235);
xnor UO_2247 (O_2247,N_27756,N_25827);
nor UO_2248 (O_2248,N_25977,N_28723);
nor UO_2249 (O_2249,N_25392,N_28845);
nor UO_2250 (O_2250,N_27293,N_29184);
nor UO_2251 (O_2251,N_27925,N_28584);
nand UO_2252 (O_2252,N_29156,N_28465);
and UO_2253 (O_2253,N_28855,N_27055);
nand UO_2254 (O_2254,N_26822,N_25194);
nor UO_2255 (O_2255,N_28408,N_29066);
nand UO_2256 (O_2256,N_28969,N_27625);
nand UO_2257 (O_2257,N_26243,N_29227);
nand UO_2258 (O_2258,N_25713,N_28500);
or UO_2259 (O_2259,N_27348,N_25813);
or UO_2260 (O_2260,N_25318,N_25645);
and UO_2261 (O_2261,N_25671,N_26729);
or UO_2262 (O_2262,N_29604,N_26495);
or UO_2263 (O_2263,N_26606,N_25688);
nor UO_2264 (O_2264,N_29217,N_25723);
nor UO_2265 (O_2265,N_27117,N_29902);
and UO_2266 (O_2266,N_28349,N_26193);
or UO_2267 (O_2267,N_26179,N_27203);
and UO_2268 (O_2268,N_26862,N_28539);
nor UO_2269 (O_2269,N_26726,N_28111);
nand UO_2270 (O_2270,N_27137,N_28040);
nor UO_2271 (O_2271,N_26546,N_26697);
or UO_2272 (O_2272,N_28572,N_26059);
nand UO_2273 (O_2273,N_27637,N_28024);
nand UO_2274 (O_2274,N_26262,N_25166);
and UO_2275 (O_2275,N_25971,N_29025);
and UO_2276 (O_2276,N_25618,N_25742);
or UO_2277 (O_2277,N_27755,N_25158);
and UO_2278 (O_2278,N_28124,N_28930);
and UO_2279 (O_2279,N_29638,N_29852);
nor UO_2280 (O_2280,N_27004,N_27723);
and UO_2281 (O_2281,N_25354,N_28336);
or UO_2282 (O_2282,N_27743,N_26286);
xor UO_2283 (O_2283,N_26644,N_27094);
nor UO_2284 (O_2284,N_25193,N_29089);
or UO_2285 (O_2285,N_25143,N_26829);
and UO_2286 (O_2286,N_25735,N_29311);
nor UO_2287 (O_2287,N_26775,N_26743);
nand UO_2288 (O_2288,N_28807,N_25371);
and UO_2289 (O_2289,N_27648,N_27985);
nor UO_2290 (O_2290,N_29315,N_25345);
nand UO_2291 (O_2291,N_28641,N_26220);
or UO_2292 (O_2292,N_27226,N_25240);
or UO_2293 (O_2293,N_28002,N_27564);
and UO_2294 (O_2294,N_27107,N_25782);
or UO_2295 (O_2295,N_29917,N_25429);
nand UO_2296 (O_2296,N_27075,N_29788);
nor UO_2297 (O_2297,N_25301,N_26548);
and UO_2298 (O_2298,N_28121,N_26356);
and UO_2299 (O_2299,N_25024,N_25703);
and UO_2300 (O_2300,N_26708,N_28600);
nor UO_2301 (O_2301,N_29285,N_27330);
nor UO_2302 (O_2302,N_26927,N_25522);
nand UO_2303 (O_2303,N_27979,N_27678);
nand UO_2304 (O_2304,N_26809,N_25312);
nand UO_2305 (O_2305,N_27761,N_25274);
nor UO_2306 (O_2306,N_29342,N_29786);
nand UO_2307 (O_2307,N_26554,N_26684);
and UO_2308 (O_2308,N_26330,N_25088);
or UO_2309 (O_2309,N_29425,N_25014);
nand UO_2310 (O_2310,N_25459,N_27424);
and UO_2311 (O_2311,N_26334,N_27832);
or UO_2312 (O_2312,N_28468,N_29499);
and UO_2313 (O_2313,N_27059,N_25407);
or UO_2314 (O_2314,N_28167,N_26001);
or UO_2315 (O_2315,N_28872,N_28353);
xor UO_2316 (O_2316,N_27291,N_28586);
nor UO_2317 (O_2317,N_29068,N_26995);
nand UO_2318 (O_2318,N_25201,N_25217);
and UO_2319 (O_2319,N_25030,N_27947);
nor UO_2320 (O_2320,N_28823,N_26162);
and UO_2321 (O_2321,N_25408,N_28119);
nor UO_2322 (O_2322,N_29078,N_29213);
xnor UO_2323 (O_2323,N_25341,N_28988);
nand UO_2324 (O_2324,N_25513,N_29086);
and UO_2325 (O_2325,N_27322,N_25472);
nor UO_2326 (O_2326,N_29659,N_29860);
nand UO_2327 (O_2327,N_26441,N_29785);
and UO_2328 (O_2328,N_25314,N_25216);
and UO_2329 (O_2329,N_25722,N_29602);
nand UO_2330 (O_2330,N_29724,N_28010);
or UO_2331 (O_2331,N_28570,N_26222);
or UO_2332 (O_2332,N_28032,N_28897);
and UO_2333 (O_2333,N_28865,N_28215);
or UO_2334 (O_2334,N_27525,N_28911);
nand UO_2335 (O_2335,N_28581,N_28137);
nor UO_2336 (O_2336,N_26488,N_29989);
nand UO_2337 (O_2337,N_28571,N_28423);
and UO_2338 (O_2338,N_29235,N_28399);
or UO_2339 (O_2339,N_27509,N_29006);
xnor UO_2340 (O_2340,N_26404,N_27175);
and UO_2341 (O_2341,N_25475,N_25689);
nor UO_2342 (O_2342,N_27041,N_29776);
and UO_2343 (O_2343,N_28420,N_26318);
nor UO_2344 (O_2344,N_27209,N_27419);
xor UO_2345 (O_2345,N_26476,N_27305);
and UO_2346 (O_2346,N_25307,N_28844);
or UO_2347 (O_2347,N_25497,N_27169);
xnor UO_2348 (O_2348,N_26701,N_29240);
xor UO_2349 (O_2349,N_25456,N_29697);
and UO_2350 (O_2350,N_26086,N_26648);
or UO_2351 (O_2351,N_27999,N_29305);
or UO_2352 (O_2352,N_28431,N_29190);
nand UO_2353 (O_2353,N_29625,N_25670);
and UO_2354 (O_2354,N_28122,N_25989);
or UO_2355 (O_2355,N_25585,N_29389);
or UO_2356 (O_2356,N_26315,N_26241);
or UO_2357 (O_2357,N_28248,N_26637);
nor UO_2358 (O_2358,N_25625,N_28881);
nor UO_2359 (O_2359,N_27272,N_25835);
nand UO_2360 (O_2360,N_25229,N_27660);
and UO_2361 (O_2361,N_27412,N_28515);
nor UO_2362 (O_2362,N_27271,N_26759);
nor UO_2363 (O_2363,N_28051,N_26312);
or UO_2364 (O_2364,N_26616,N_28201);
or UO_2365 (O_2365,N_29281,N_28941);
nor UO_2366 (O_2366,N_29082,N_25624);
or UO_2367 (O_2367,N_28178,N_29585);
and UO_2368 (O_2368,N_26513,N_25559);
nand UO_2369 (O_2369,N_26496,N_25727);
and UO_2370 (O_2370,N_29307,N_27843);
or UO_2371 (O_2371,N_27292,N_26278);
or UO_2372 (O_2372,N_29282,N_25433);
nand UO_2373 (O_2373,N_25868,N_25548);
xor UO_2374 (O_2374,N_29729,N_29102);
or UO_2375 (O_2375,N_28895,N_26910);
nor UO_2376 (O_2376,N_29157,N_28390);
and UO_2377 (O_2377,N_25401,N_25797);
nor UO_2378 (O_2378,N_25104,N_26501);
and UO_2379 (O_2379,N_25982,N_27230);
nand UO_2380 (O_2380,N_27437,N_25956);
and UO_2381 (O_2381,N_27120,N_25978);
and UO_2382 (O_2382,N_25949,N_25533);
or UO_2383 (O_2383,N_29382,N_29943);
nand UO_2384 (O_2384,N_26738,N_25377);
and UO_2385 (O_2385,N_25121,N_29369);
or UO_2386 (O_2386,N_29262,N_27286);
nand UO_2387 (O_2387,N_25395,N_28951);
nor UO_2388 (O_2388,N_28088,N_25184);
nor UO_2389 (O_2389,N_25639,N_28131);
and UO_2390 (O_2390,N_26716,N_26863);
nand UO_2391 (O_2391,N_27961,N_26250);
or UO_2392 (O_2392,N_26610,N_29177);
or UO_2393 (O_2393,N_26065,N_29225);
and UO_2394 (O_2394,N_28042,N_29991);
nand UO_2395 (O_2395,N_26135,N_25265);
and UO_2396 (O_2396,N_27592,N_28140);
or UO_2397 (O_2397,N_26094,N_28992);
nor UO_2398 (O_2398,N_27864,N_29596);
or UO_2399 (O_2399,N_25247,N_29843);
nand UO_2400 (O_2400,N_26549,N_26099);
nor UO_2401 (O_2401,N_28989,N_28463);
nor UO_2402 (O_2402,N_25093,N_27470);
nand UO_2403 (O_2403,N_25373,N_25224);
and UO_2404 (O_2404,N_25214,N_26785);
nor UO_2405 (O_2405,N_26448,N_25110);
nor UO_2406 (O_2406,N_28635,N_28235);
or UO_2407 (O_2407,N_29090,N_26398);
or UO_2408 (O_2408,N_28182,N_29512);
or UO_2409 (O_2409,N_29221,N_27314);
or UO_2410 (O_2410,N_27091,N_29505);
nor UO_2411 (O_2411,N_25974,N_26652);
or UO_2412 (O_2412,N_28551,N_25793);
and UO_2413 (O_2413,N_25033,N_28858);
nor UO_2414 (O_2414,N_25524,N_28561);
and UO_2415 (O_2415,N_27512,N_25137);
and UO_2416 (O_2416,N_25595,N_29428);
and UO_2417 (O_2417,N_25493,N_26485);
and UO_2418 (O_2418,N_27499,N_26744);
or UO_2419 (O_2419,N_27816,N_29737);
or UO_2420 (O_2420,N_28752,N_27434);
and UO_2421 (O_2421,N_29630,N_28620);
or UO_2422 (O_2422,N_29019,N_28882);
and UO_2423 (O_2423,N_29761,N_28106);
nor UO_2424 (O_2424,N_29525,N_28093);
nor UO_2425 (O_2425,N_27376,N_29657);
or UO_2426 (O_2426,N_28450,N_29222);
and UO_2427 (O_2427,N_26812,N_28607);
nor UO_2428 (O_2428,N_25457,N_27340);
nand UO_2429 (O_2429,N_27728,N_28673);
and UO_2430 (O_2430,N_26484,N_25950);
and UO_2431 (O_2431,N_28583,N_29749);
or UO_2432 (O_2432,N_25049,N_25588);
and UO_2433 (O_2433,N_28773,N_28041);
xnor UO_2434 (O_2434,N_28000,N_26578);
nand UO_2435 (O_2435,N_28212,N_28758);
nand UO_2436 (O_2436,N_25740,N_29867);
nand UO_2437 (O_2437,N_26901,N_29272);
or UO_2438 (O_2438,N_26924,N_27927);
nand UO_2439 (O_2439,N_25113,N_29796);
or UO_2440 (O_2440,N_29471,N_27382);
nand UO_2441 (O_2441,N_26755,N_29529);
and UO_2442 (O_2442,N_27431,N_26120);
nor UO_2443 (O_2443,N_25048,N_26757);
nor UO_2444 (O_2444,N_29085,N_29694);
nand UO_2445 (O_2445,N_28422,N_28973);
nand UO_2446 (O_2446,N_29278,N_27996);
or UO_2447 (O_2447,N_25547,N_25826);
or UO_2448 (O_2448,N_26041,N_29466);
nand UO_2449 (O_2449,N_28456,N_25442);
nor UO_2450 (O_2450,N_29762,N_26535);
or UO_2451 (O_2451,N_26038,N_26603);
nor UO_2452 (O_2452,N_28634,N_27770);
nor UO_2453 (O_2453,N_27327,N_29722);
and UO_2454 (O_2454,N_25661,N_26473);
or UO_2455 (O_2455,N_28409,N_25323);
nand UO_2456 (O_2456,N_27975,N_25439);
and UO_2457 (O_2457,N_28715,N_29967);
nand UO_2458 (O_2458,N_27126,N_25986);
and UO_2459 (O_2459,N_25075,N_28924);
and UO_2460 (O_2460,N_29794,N_26853);
and UO_2461 (O_2461,N_25532,N_29299);
and UO_2462 (O_2462,N_29795,N_25449);
and UO_2463 (O_2463,N_29091,N_29666);
nor UO_2464 (O_2464,N_27151,N_25720);
nor UO_2465 (O_2465,N_25289,N_28959);
nand UO_2466 (O_2466,N_26128,N_27485);
or UO_2467 (O_2467,N_29117,N_28474);
nor UO_2468 (O_2468,N_27317,N_29515);
or UO_2469 (O_2469,N_26796,N_27614);
nand UO_2470 (O_2470,N_25844,N_26921);
or UO_2471 (O_2471,N_29241,N_27859);
and UO_2472 (O_2472,N_29844,N_28730);
nor UO_2473 (O_2473,N_26516,N_29829);
nor UO_2474 (O_2474,N_29813,N_29208);
and UO_2475 (O_2475,N_27702,N_26229);
nand UO_2476 (O_2476,N_25065,N_29942);
and UO_2477 (O_2477,N_28066,N_27136);
nor UO_2478 (O_2478,N_25119,N_28591);
nor UO_2479 (O_2479,N_26300,N_29836);
or UO_2480 (O_2480,N_25829,N_25425);
nor UO_2481 (O_2481,N_27304,N_28084);
nand UO_2482 (O_2482,N_26857,N_29805);
nand UO_2483 (O_2483,N_27489,N_26159);
or UO_2484 (O_2484,N_28067,N_27692);
or UO_2485 (O_2485,N_27661,N_25644);
nor UO_2486 (O_2486,N_26902,N_25928);
nand UO_2487 (O_2487,N_29393,N_29409);
and UO_2488 (O_2488,N_26994,N_28373);
and UO_2489 (O_2489,N_28664,N_28883);
or UO_2490 (O_2490,N_26791,N_29322);
nor UO_2491 (O_2491,N_28281,N_26687);
and UO_2492 (O_2492,N_28819,N_28642);
and UO_2493 (O_2493,N_27214,N_25069);
xor UO_2494 (O_2494,N_27919,N_29835);
nor UO_2495 (O_2495,N_27462,N_25204);
or UO_2496 (O_2496,N_26925,N_26386);
or UO_2497 (O_2497,N_29265,N_29408);
and UO_2498 (O_2498,N_29889,N_29899);
or UO_2499 (O_2499,N_25601,N_27034);
nor UO_2500 (O_2500,N_29290,N_27201);
or UO_2501 (O_2501,N_29293,N_27174);
nor UO_2502 (O_2502,N_29488,N_27815);
or UO_2503 (O_2503,N_27768,N_27035);
and UO_2504 (O_2504,N_25749,N_28524);
or UO_2505 (O_2505,N_27703,N_25254);
or UO_2506 (O_2506,N_29729,N_29842);
nand UO_2507 (O_2507,N_26795,N_26540);
nand UO_2508 (O_2508,N_26720,N_27259);
or UO_2509 (O_2509,N_25796,N_29590);
and UO_2510 (O_2510,N_26822,N_29282);
xor UO_2511 (O_2511,N_25820,N_27852);
and UO_2512 (O_2512,N_28143,N_27701);
nor UO_2513 (O_2513,N_25756,N_26554);
nor UO_2514 (O_2514,N_27669,N_25533);
nor UO_2515 (O_2515,N_26893,N_26494);
nand UO_2516 (O_2516,N_27456,N_25823);
or UO_2517 (O_2517,N_26835,N_25115);
or UO_2518 (O_2518,N_26854,N_29466);
nor UO_2519 (O_2519,N_28175,N_28228);
and UO_2520 (O_2520,N_27127,N_29695);
or UO_2521 (O_2521,N_26209,N_28635);
and UO_2522 (O_2522,N_26787,N_29914);
or UO_2523 (O_2523,N_29331,N_28224);
nand UO_2524 (O_2524,N_27134,N_28889);
and UO_2525 (O_2525,N_26664,N_29301);
nand UO_2526 (O_2526,N_28502,N_26819);
nand UO_2527 (O_2527,N_28208,N_28796);
nor UO_2528 (O_2528,N_27998,N_26594);
nand UO_2529 (O_2529,N_29898,N_25089);
and UO_2530 (O_2530,N_26948,N_27123);
nor UO_2531 (O_2531,N_27831,N_27156);
nor UO_2532 (O_2532,N_29488,N_26197);
nand UO_2533 (O_2533,N_29249,N_29806);
and UO_2534 (O_2534,N_28591,N_28252);
xor UO_2535 (O_2535,N_29632,N_25546);
nand UO_2536 (O_2536,N_26976,N_27680);
nor UO_2537 (O_2537,N_28804,N_25542);
nor UO_2538 (O_2538,N_28674,N_27203);
and UO_2539 (O_2539,N_27891,N_27374);
or UO_2540 (O_2540,N_28904,N_25082);
nand UO_2541 (O_2541,N_27040,N_28769);
nand UO_2542 (O_2542,N_27219,N_26185);
nor UO_2543 (O_2543,N_26224,N_26049);
and UO_2544 (O_2544,N_27616,N_28802);
or UO_2545 (O_2545,N_29746,N_27983);
nor UO_2546 (O_2546,N_29286,N_26748);
and UO_2547 (O_2547,N_27225,N_26746);
or UO_2548 (O_2548,N_25973,N_27001);
nand UO_2549 (O_2549,N_27868,N_25364);
and UO_2550 (O_2550,N_25109,N_29472);
nor UO_2551 (O_2551,N_25555,N_26801);
or UO_2552 (O_2552,N_28740,N_26281);
nor UO_2553 (O_2553,N_28242,N_27173);
or UO_2554 (O_2554,N_29484,N_29727);
or UO_2555 (O_2555,N_25219,N_28737);
or UO_2556 (O_2556,N_27566,N_25200);
xor UO_2557 (O_2557,N_29856,N_28106);
nand UO_2558 (O_2558,N_28148,N_29688);
or UO_2559 (O_2559,N_27978,N_27942);
and UO_2560 (O_2560,N_25751,N_25620);
nor UO_2561 (O_2561,N_28562,N_27908);
and UO_2562 (O_2562,N_27824,N_28480);
xnor UO_2563 (O_2563,N_28917,N_25895);
nor UO_2564 (O_2564,N_28536,N_26972);
nor UO_2565 (O_2565,N_25009,N_26258);
nand UO_2566 (O_2566,N_25383,N_25357);
or UO_2567 (O_2567,N_26716,N_28510);
or UO_2568 (O_2568,N_27983,N_25508);
nand UO_2569 (O_2569,N_27953,N_27636);
or UO_2570 (O_2570,N_25079,N_29090);
and UO_2571 (O_2571,N_29152,N_28433);
xor UO_2572 (O_2572,N_25600,N_27179);
and UO_2573 (O_2573,N_26725,N_28545);
nor UO_2574 (O_2574,N_29604,N_28655);
or UO_2575 (O_2575,N_28034,N_25530);
and UO_2576 (O_2576,N_29123,N_27973);
nor UO_2577 (O_2577,N_28426,N_29387);
nand UO_2578 (O_2578,N_28016,N_26108);
or UO_2579 (O_2579,N_29919,N_25114);
and UO_2580 (O_2580,N_26611,N_25884);
and UO_2581 (O_2581,N_29429,N_28049);
nor UO_2582 (O_2582,N_28454,N_27747);
and UO_2583 (O_2583,N_25255,N_25953);
nand UO_2584 (O_2584,N_29063,N_27784);
nor UO_2585 (O_2585,N_28639,N_27481);
nor UO_2586 (O_2586,N_28947,N_27592);
or UO_2587 (O_2587,N_26469,N_29430);
or UO_2588 (O_2588,N_26663,N_26852);
and UO_2589 (O_2589,N_28580,N_28156);
nand UO_2590 (O_2590,N_29374,N_29322);
nor UO_2591 (O_2591,N_26442,N_25153);
and UO_2592 (O_2592,N_27575,N_25626);
and UO_2593 (O_2593,N_28500,N_25391);
nand UO_2594 (O_2594,N_28453,N_27602);
nor UO_2595 (O_2595,N_28952,N_26046);
nor UO_2596 (O_2596,N_28665,N_25790);
and UO_2597 (O_2597,N_29682,N_28556);
xor UO_2598 (O_2598,N_28345,N_27165);
xnor UO_2599 (O_2599,N_29112,N_25603);
or UO_2600 (O_2600,N_29057,N_28171);
and UO_2601 (O_2601,N_29965,N_25787);
or UO_2602 (O_2602,N_25430,N_27649);
and UO_2603 (O_2603,N_25669,N_26037);
nor UO_2604 (O_2604,N_28071,N_28191);
nand UO_2605 (O_2605,N_28401,N_29261);
nor UO_2606 (O_2606,N_29282,N_27200);
xnor UO_2607 (O_2607,N_25979,N_25667);
or UO_2608 (O_2608,N_25847,N_27173);
nor UO_2609 (O_2609,N_27308,N_29990);
nor UO_2610 (O_2610,N_25467,N_25800);
nand UO_2611 (O_2611,N_28103,N_26363);
nor UO_2612 (O_2612,N_29255,N_25080);
nor UO_2613 (O_2613,N_28406,N_28099);
nand UO_2614 (O_2614,N_29688,N_29530);
or UO_2615 (O_2615,N_29980,N_28193);
and UO_2616 (O_2616,N_27491,N_28889);
xnor UO_2617 (O_2617,N_27191,N_25513);
nor UO_2618 (O_2618,N_27257,N_28451);
and UO_2619 (O_2619,N_27811,N_27972);
and UO_2620 (O_2620,N_25418,N_27036);
nand UO_2621 (O_2621,N_26974,N_25552);
and UO_2622 (O_2622,N_26906,N_26207);
nor UO_2623 (O_2623,N_28292,N_27048);
and UO_2624 (O_2624,N_28920,N_27978);
nor UO_2625 (O_2625,N_28165,N_26084);
or UO_2626 (O_2626,N_29853,N_26836);
nor UO_2627 (O_2627,N_27937,N_28524);
nor UO_2628 (O_2628,N_28313,N_29189);
nand UO_2629 (O_2629,N_27299,N_28599);
nor UO_2630 (O_2630,N_28276,N_28550);
and UO_2631 (O_2631,N_25165,N_27446);
nor UO_2632 (O_2632,N_29566,N_28736);
or UO_2633 (O_2633,N_28429,N_27392);
or UO_2634 (O_2634,N_28362,N_27783);
nand UO_2635 (O_2635,N_25120,N_25172);
nand UO_2636 (O_2636,N_27482,N_25285);
or UO_2637 (O_2637,N_26663,N_29083);
nor UO_2638 (O_2638,N_27216,N_27555);
and UO_2639 (O_2639,N_28265,N_25795);
and UO_2640 (O_2640,N_27312,N_29437);
nand UO_2641 (O_2641,N_25179,N_26177);
xor UO_2642 (O_2642,N_25437,N_26342);
and UO_2643 (O_2643,N_27016,N_26052);
or UO_2644 (O_2644,N_28638,N_26259);
and UO_2645 (O_2645,N_26331,N_28156);
and UO_2646 (O_2646,N_27553,N_29575);
nor UO_2647 (O_2647,N_28356,N_26602);
or UO_2648 (O_2648,N_29121,N_28462);
or UO_2649 (O_2649,N_26718,N_28495);
nand UO_2650 (O_2650,N_25481,N_27021);
or UO_2651 (O_2651,N_26549,N_25764);
nand UO_2652 (O_2652,N_28583,N_25581);
and UO_2653 (O_2653,N_28873,N_26444);
nand UO_2654 (O_2654,N_25865,N_25654);
or UO_2655 (O_2655,N_27555,N_28260);
or UO_2656 (O_2656,N_28451,N_27045);
nor UO_2657 (O_2657,N_28928,N_27772);
or UO_2658 (O_2658,N_29000,N_27936);
nand UO_2659 (O_2659,N_25286,N_28832);
and UO_2660 (O_2660,N_26742,N_25025);
nor UO_2661 (O_2661,N_28156,N_28672);
or UO_2662 (O_2662,N_26784,N_27825);
and UO_2663 (O_2663,N_28641,N_25453);
or UO_2664 (O_2664,N_25188,N_25560);
xnor UO_2665 (O_2665,N_26076,N_25759);
xnor UO_2666 (O_2666,N_25123,N_27946);
nand UO_2667 (O_2667,N_25979,N_29450);
nand UO_2668 (O_2668,N_28331,N_28439);
nor UO_2669 (O_2669,N_27212,N_29483);
nand UO_2670 (O_2670,N_28521,N_29107);
or UO_2671 (O_2671,N_26486,N_29026);
nand UO_2672 (O_2672,N_25299,N_27014);
and UO_2673 (O_2673,N_29654,N_29862);
nor UO_2674 (O_2674,N_25599,N_27462);
nor UO_2675 (O_2675,N_28939,N_25930);
and UO_2676 (O_2676,N_26259,N_27466);
and UO_2677 (O_2677,N_26754,N_28885);
nand UO_2678 (O_2678,N_28407,N_26943);
or UO_2679 (O_2679,N_29364,N_25015);
or UO_2680 (O_2680,N_27598,N_27858);
nand UO_2681 (O_2681,N_28971,N_25346);
xnor UO_2682 (O_2682,N_25546,N_26117);
and UO_2683 (O_2683,N_29308,N_26365);
and UO_2684 (O_2684,N_29208,N_27452);
or UO_2685 (O_2685,N_27187,N_26487);
and UO_2686 (O_2686,N_27085,N_29237);
or UO_2687 (O_2687,N_28513,N_25153);
nand UO_2688 (O_2688,N_27135,N_29930);
xor UO_2689 (O_2689,N_29017,N_26120);
or UO_2690 (O_2690,N_28199,N_25046);
nor UO_2691 (O_2691,N_25607,N_27233);
nand UO_2692 (O_2692,N_28825,N_28418);
nor UO_2693 (O_2693,N_27619,N_25132);
nor UO_2694 (O_2694,N_26895,N_25089);
nand UO_2695 (O_2695,N_25013,N_27047);
nor UO_2696 (O_2696,N_26312,N_29034);
nor UO_2697 (O_2697,N_27945,N_28738);
nand UO_2698 (O_2698,N_28731,N_29891);
or UO_2699 (O_2699,N_26938,N_26918);
nand UO_2700 (O_2700,N_26974,N_28862);
nand UO_2701 (O_2701,N_28101,N_28318);
nand UO_2702 (O_2702,N_26779,N_27079);
and UO_2703 (O_2703,N_26143,N_26522);
nor UO_2704 (O_2704,N_27248,N_29361);
nand UO_2705 (O_2705,N_27102,N_28855);
and UO_2706 (O_2706,N_29901,N_28203);
and UO_2707 (O_2707,N_27905,N_27226);
nand UO_2708 (O_2708,N_26634,N_26952);
xor UO_2709 (O_2709,N_28044,N_29233);
or UO_2710 (O_2710,N_26580,N_26394);
nand UO_2711 (O_2711,N_26098,N_28821);
nand UO_2712 (O_2712,N_29932,N_26706);
and UO_2713 (O_2713,N_25591,N_29769);
nor UO_2714 (O_2714,N_28598,N_26377);
nor UO_2715 (O_2715,N_25255,N_26103);
or UO_2716 (O_2716,N_25414,N_29052);
or UO_2717 (O_2717,N_26172,N_29909);
and UO_2718 (O_2718,N_29414,N_27334);
or UO_2719 (O_2719,N_26708,N_27880);
and UO_2720 (O_2720,N_27436,N_29693);
or UO_2721 (O_2721,N_29393,N_29286);
nand UO_2722 (O_2722,N_28175,N_27181);
nor UO_2723 (O_2723,N_29596,N_26488);
nand UO_2724 (O_2724,N_29368,N_27812);
xor UO_2725 (O_2725,N_28986,N_26138);
or UO_2726 (O_2726,N_29890,N_28718);
xor UO_2727 (O_2727,N_27148,N_29584);
nor UO_2728 (O_2728,N_27008,N_27847);
and UO_2729 (O_2729,N_28026,N_25430);
and UO_2730 (O_2730,N_29934,N_26805);
and UO_2731 (O_2731,N_26519,N_25549);
and UO_2732 (O_2732,N_29047,N_25386);
and UO_2733 (O_2733,N_25282,N_27433);
nor UO_2734 (O_2734,N_27052,N_25557);
or UO_2735 (O_2735,N_29562,N_27577);
or UO_2736 (O_2736,N_25735,N_27167);
nor UO_2737 (O_2737,N_25029,N_27089);
and UO_2738 (O_2738,N_25674,N_27580);
nor UO_2739 (O_2739,N_26744,N_28110);
nand UO_2740 (O_2740,N_27173,N_25875);
nor UO_2741 (O_2741,N_29566,N_28974);
xor UO_2742 (O_2742,N_29158,N_27661);
and UO_2743 (O_2743,N_25612,N_26063);
nor UO_2744 (O_2744,N_27158,N_28473);
or UO_2745 (O_2745,N_26443,N_28229);
and UO_2746 (O_2746,N_28975,N_28587);
nand UO_2747 (O_2747,N_25026,N_28999);
and UO_2748 (O_2748,N_26048,N_27398);
and UO_2749 (O_2749,N_25597,N_25184);
or UO_2750 (O_2750,N_26055,N_26527);
nor UO_2751 (O_2751,N_28558,N_27104);
or UO_2752 (O_2752,N_28167,N_28550);
xor UO_2753 (O_2753,N_25083,N_29163);
and UO_2754 (O_2754,N_26730,N_25021);
xnor UO_2755 (O_2755,N_25611,N_27116);
and UO_2756 (O_2756,N_26857,N_29781);
or UO_2757 (O_2757,N_25395,N_25853);
or UO_2758 (O_2758,N_25546,N_28785);
or UO_2759 (O_2759,N_28747,N_25263);
and UO_2760 (O_2760,N_28668,N_28794);
or UO_2761 (O_2761,N_26715,N_28637);
or UO_2762 (O_2762,N_28153,N_27233);
or UO_2763 (O_2763,N_28641,N_26872);
and UO_2764 (O_2764,N_29482,N_27147);
nand UO_2765 (O_2765,N_26532,N_29357);
and UO_2766 (O_2766,N_25785,N_26542);
nand UO_2767 (O_2767,N_27864,N_26850);
and UO_2768 (O_2768,N_26103,N_29045);
and UO_2769 (O_2769,N_29392,N_25101);
or UO_2770 (O_2770,N_25035,N_28404);
xnor UO_2771 (O_2771,N_27273,N_27008);
or UO_2772 (O_2772,N_26454,N_29020);
nor UO_2773 (O_2773,N_26158,N_28169);
nor UO_2774 (O_2774,N_28384,N_28064);
xnor UO_2775 (O_2775,N_29853,N_28680);
nand UO_2776 (O_2776,N_25049,N_25017);
nor UO_2777 (O_2777,N_28936,N_28771);
nand UO_2778 (O_2778,N_25569,N_27845);
or UO_2779 (O_2779,N_25882,N_26854);
nor UO_2780 (O_2780,N_25478,N_29693);
nor UO_2781 (O_2781,N_26964,N_28885);
nor UO_2782 (O_2782,N_26912,N_28923);
and UO_2783 (O_2783,N_26430,N_26808);
and UO_2784 (O_2784,N_26459,N_28816);
or UO_2785 (O_2785,N_27983,N_25546);
or UO_2786 (O_2786,N_29785,N_29289);
nor UO_2787 (O_2787,N_28206,N_27249);
nor UO_2788 (O_2788,N_25332,N_29324);
nor UO_2789 (O_2789,N_29488,N_26062);
xnor UO_2790 (O_2790,N_28303,N_28971);
and UO_2791 (O_2791,N_29201,N_26366);
or UO_2792 (O_2792,N_26722,N_28493);
nand UO_2793 (O_2793,N_28318,N_27329);
nand UO_2794 (O_2794,N_29135,N_27262);
or UO_2795 (O_2795,N_28418,N_25897);
or UO_2796 (O_2796,N_29563,N_28288);
xnor UO_2797 (O_2797,N_27339,N_25865);
or UO_2798 (O_2798,N_27356,N_28034);
or UO_2799 (O_2799,N_26832,N_27330);
nand UO_2800 (O_2800,N_29819,N_28784);
or UO_2801 (O_2801,N_29803,N_25857);
or UO_2802 (O_2802,N_29096,N_25786);
nand UO_2803 (O_2803,N_29631,N_25940);
or UO_2804 (O_2804,N_28124,N_28553);
and UO_2805 (O_2805,N_25775,N_26240);
nor UO_2806 (O_2806,N_28639,N_27358);
nand UO_2807 (O_2807,N_28536,N_26535);
and UO_2808 (O_2808,N_28118,N_27069);
nor UO_2809 (O_2809,N_27838,N_25819);
nor UO_2810 (O_2810,N_28554,N_28624);
and UO_2811 (O_2811,N_25364,N_26089);
xor UO_2812 (O_2812,N_29028,N_28976);
and UO_2813 (O_2813,N_28750,N_28641);
nor UO_2814 (O_2814,N_26275,N_26160);
nand UO_2815 (O_2815,N_28664,N_27134);
nor UO_2816 (O_2816,N_26548,N_29853);
nor UO_2817 (O_2817,N_26532,N_27163);
nand UO_2818 (O_2818,N_27559,N_27790);
nor UO_2819 (O_2819,N_26064,N_25834);
xor UO_2820 (O_2820,N_29883,N_26643);
nor UO_2821 (O_2821,N_28055,N_25483);
and UO_2822 (O_2822,N_27141,N_26698);
xnor UO_2823 (O_2823,N_28239,N_27795);
or UO_2824 (O_2824,N_25391,N_28251);
nor UO_2825 (O_2825,N_27264,N_25957);
or UO_2826 (O_2826,N_28351,N_26205);
nand UO_2827 (O_2827,N_29636,N_27991);
and UO_2828 (O_2828,N_25970,N_28390);
nor UO_2829 (O_2829,N_26033,N_26226);
nor UO_2830 (O_2830,N_25223,N_25594);
nor UO_2831 (O_2831,N_27778,N_27026);
nor UO_2832 (O_2832,N_29550,N_26599);
and UO_2833 (O_2833,N_28368,N_29893);
nand UO_2834 (O_2834,N_26927,N_29969);
nor UO_2835 (O_2835,N_27618,N_26095);
and UO_2836 (O_2836,N_26183,N_29903);
nor UO_2837 (O_2837,N_28843,N_29444);
nor UO_2838 (O_2838,N_26089,N_29304);
or UO_2839 (O_2839,N_25465,N_27764);
nor UO_2840 (O_2840,N_28381,N_29400);
nor UO_2841 (O_2841,N_25651,N_27669);
nor UO_2842 (O_2842,N_28083,N_29758);
xnor UO_2843 (O_2843,N_26165,N_28669);
nand UO_2844 (O_2844,N_28689,N_29631);
xnor UO_2845 (O_2845,N_28378,N_29391);
nor UO_2846 (O_2846,N_29826,N_25200);
and UO_2847 (O_2847,N_29559,N_29413);
nand UO_2848 (O_2848,N_27146,N_25201);
nor UO_2849 (O_2849,N_28490,N_29098);
nand UO_2850 (O_2850,N_25840,N_26413);
or UO_2851 (O_2851,N_27247,N_26369);
or UO_2852 (O_2852,N_29517,N_27286);
or UO_2853 (O_2853,N_26066,N_29797);
or UO_2854 (O_2854,N_27845,N_25360);
or UO_2855 (O_2855,N_26038,N_25393);
or UO_2856 (O_2856,N_28323,N_29769);
xnor UO_2857 (O_2857,N_26698,N_28498);
or UO_2858 (O_2858,N_26128,N_27546);
xnor UO_2859 (O_2859,N_27219,N_25708);
nor UO_2860 (O_2860,N_26513,N_25382);
or UO_2861 (O_2861,N_25978,N_26153);
and UO_2862 (O_2862,N_25716,N_26971);
or UO_2863 (O_2863,N_28635,N_25188);
xnor UO_2864 (O_2864,N_28894,N_25851);
and UO_2865 (O_2865,N_27581,N_25461);
nor UO_2866 (O_2866,N_27233,N_28744);
or UO_2867 (O_2867,N_27538,N_27523);
nor UO_2868 (O_2868,N_28930,N_28438);
and UO_2869 (O_2869,N_29238,N_28519);
nor UO_2870 (O_2870,N_26474,N_28365);
and UO_2871 (O_2871,N_25372,N_26307);
or UO_2872 (O_2872,N_29225,N_25658);
and UO_2873 (O_2873,N_25140,N_29886);
nand UO_2874 (O_2874,N_29988,N_27347);
or UO_2875 (O_2875,N_27826,N_25905);
nor UO_2876 (O_2876,N_28350,N_28189);
and UO_2877 (O_2877,N_27467,N_25218);
nor UO_2878 (O_2878,N_27549,N_28442);
xnor UO_2879 (O_2879,N_29821,N_29407);
nor UO_2880 (O_2880,N_25184,N_27463);
nand UO_2881 (O_2881,N_27142,N_25283);
and UO_2882 (O_2882,N_26549,N_29207);
and UO_2883 (O_2883,N_28761,N_28519);
xnor UO_2884 (O_2884,N_25444,N_25851);
xor UO_2885 (O_2885,N_25845,N_29159);
or UO_2886 (O_2886,N_26829,N_27380);
or UO_2887 (O_2887,N_26587,N_25755);
nand UO_2888 (O_2888,N_29415,N_25597);
nand UO_2889 (O_2889,N_25100,N_27239);
nor UO_2890 (O_2890,N_26571,N_26379);
nor UO_2891 (O_2891,N_29164,N_26034);
nor UO_2892 (O_2892,N_29651,N_26334);
or UO_2893 (O_2893,N_28700,N_27718);
and UO_2894 (O_2894,N_27573,N_25787);
or UO_2895 (O_2895,N_29366,N_26746);
nand UO_2896 (O_2896,N_27003,N_27110);
xor UO_2897 (O_2897,N_27177,N_28861);
xor UO_2898 (O_2898,N_26950,N_25927);
nand UO_2899 (O_2899,N_27655,N_28214);
or UO_2900 (O_2900,N_29168,N_26386);
nand UO_2901 (O_2901,N_29813,N_26490);
nand UO_2902 (O_2902,N_27900,N_28459);
nand UO_2903 (O_2903,N_27972,N_28870);
nor UO_2904 (O_2904,N_26849,N_27093);
and UO_2905 (O_2905,N_28142,N_27420);
and UO_2906 (O_2906,N_26359,N_26817);
and UO_2907 (O_2907,N_29135,N_28210);
and UO_2908 (O_2908,N_26684,N_27414);
nor UO_2909 (O_2909,N_28579,N_29175);
nand UO_2910 (O_2910,N_25022,N_29963);
nor UO_2911 (O_2911,N_26712,N_25926);
nand UO_2912 (O_2912,N_25522,N_26575);
or UO_2913 (O_2913,N_29676,N_29049);
or UO_2914 (O_2914,N_26630,N_27026);
nand UO_2915 (O_2915,N_26631,N_27486);
or UO_2916 (O_2916,N_27768,N_29797);
and UO_2917 (O_2917,N_26229,N_27743);
xor UO_2918 (O_2918,N_28402,N_25388);
xnor UO_2919 (O_2919,N_26740,N_27538);
and UO_2920 (O_2920,N_29792,N_26922);
and UO_2921 (O_2921,N_29764,N_27133);
and UO_2922 (O_2922,N_28185,N_26989);
nand UO_2923 (O_2923,N_26817,N_25006);
nor UO_2924 (O_2924,N_26904,N_29432);
or UO_2925 (O_2925,N_25287,N_29891);
or UO_2926 (O_2926,N_26111,N_25975);
nor UO_2927 (O_2927,N_25786,N_28776);
nor UO_2928 (O_2928,N_25323,N_25773);
nand UO_2929 (O_2929,N_28297,N_25005);
and UO_2930 (O_2930,N_27731,N_27942);
or UO_2931 (O_2931,N_25118,N_26166);
and UO_2932 (O_2932,N_29090,N_26357);
nand UO_2933 (O_2933,N_29330,N_26569);
nor UO_2934 (O_2934,N_28365,N_29162);
nand UO_2935 (O_2935,N_25984,N_29406);
nand UO_2936 (O_2936,N_25692,N_27061);
nand UO_2937 (O_2937,N_28770,N_26673);
or UO_2938 (O_2938,N_26594,N_26609);
or UO_2939 (O_2939,N_26174,N_28945);
nand UO_2940 (O_2940,N_28565,N_25417);
and UO_2941 (O_2941,N_28257,N_28867);
nand UO_2942 (O_2942,N_29946,N_29857);
nand UO_2943 (O_2943,N_25669,N_27845);
and UO_2944 (O_2944,N_26224,N_28181);
nor UO_2945 (O_2945,N_27091,N_28431);
and UO_2946 (O_2946,N_26466,N_29827);
and UO_2947 (O_2947,N_27054,N_29664);
or UO_2948 (O_2948,N_25486,N_28564);
nand UO_2949 (O_2949,N_29436,N_26334);
nand UO_2950 (O_2950,N_29303,N_27048);
nor UO_2951 (O_2951,N_27429,N_25257);
nor UO_2952 (O_2952,N_29524,N_27909);
nor UO_2953 (O_2953,N_26360,N_26878);
and UO_2954 (O_2954,N_25272,N_27803);
nor UO_2955 (O_2955,N_28715,N_27089);
nand UO_2956 (O_2956,N_29303,N_28977);
xnor UO_2957 (O_2957,N_27632,N_25191);
nand UO_2958 (O_2958,N_29807,N_26925);
xnor UO_2959 (O_2959,N_29361,N_27213);
xnor UO_2960 (O_2960,N_26262,N_28803);
or UO_2961 (O_2961,N_28013,N_27104);
nor UO_2962 (O_2962,N_29851,N_25751);
nor UO_2963 (O_2963,N_25294,N_28104);
nand UO_2964 (O_2964,N_26802,N_29098);
nand UO_2965 (O_2965,N_25379,N_28875);
and UO_2966 (O_2966,N_29882,N_29205);
nand UO_2967 (O_2967,N_27756,N_26260);
or UO_2968 (O_2968,N_27883,N_28060);
nor UO_2969 (O_2969,N_26399,N_29636);
nor UO_2970 (O_2970,N_25953,N_29842);
or UO_2971 (O_2971,N_29595,N_26876);
or UO_2972 (O_2972,N_27158,N_25897);
or UO_2973 (O_2973,N_28552,N_27467);
and UO_2974 (O_2974,N_29885,N_27804);
or UO_2975 (O_2975,N_27480,N_25866);
or UO_2976 (O_2976,N_27573,N_25587);
or UO_2977 (O_2977,N_29938,N_29896);
nor UO_2978 (O_2978,N_25489,N_25316);
nor UO_2979 (O_2979,N_29104,N_26639);
nand UO_2980 (O_2980,N_29961,N_25110);
nor UO_2981 (O_2981,N_28105,N_27625);
nand UO_2982 (O_2982,N_26769,N_25907);
or UO_2983 (O_2983,N_26529,N_29134);
nor UO_2984 (O_2984,N_27573,N_28122);
nand UO_2985 (O_2985,N_27399,N_27801);
and UO_2986 (O_2986,N_26706,N_28792);
and UO_2987 (O_2987,N_28539,N_29029);
or UO_2988 (O_2988,N_25574,N_28601);
or UO_2989 (O_2989,N_28511,N_27541);
xnor UO_2990 (O_2990,N_27136,N_26277);
nand UO_2991 (O_2991,N_28078,N_25738);
xor UO_2992 (O_2992,N_27818,N_27456);
or UO_2993 (O_2993,N_25543,N_27475);
and UO_2994 (O_2994,N_29897,N_26316);
nand UO_2995 (O_2995,N_27449,N_25134);
nand UO_2996 (O_2996,N_28500,N_27736);
or UO_2997 (O_2997,N_27038,N_28881);
xnor UO_2998 (O_2998,N_26871,N_26014);
and UO_2999 (O_2999,N_27601,N_27141);
nand UO_3000 (O_3000,N_27087,N_26848);
nand UO_3001 (O_3001,N_27437,N_28346);
nand UO_3002 (O_3002,N_25002,N_26983);
and UO_3003 (O_3003,N_25946,N_26521);
xnor UO_3004 (O_3004,N_27458,N_26185);
nand UO_3005 (O_3005,N_25855,N_26660);
nand UO_3006 (O_3006,N_28241,N_29374);
and UO_3007 (O_3007,N_26116,N_28077);
or UO_3008 (O_3008,N_29997,N_29786);
nor UO_3009 (O_3009,N_26204,N_26132);
nand UO_3010 (O_3010,N_28523,N_27964);
and UO_3011 (O_3011,N_27489,N_27333);
or UO_3012 (O_3012,N_25104,N_28864);
nor UO_3013 (O_3013,N_27486,N_26282);
xnor UO_3014 (O_3014,N_26528,N_28582);
and UO_3015 (O_3015,N_26127,N_25312);
or UO_3016 (O_3016,N_28119,N_25714);
nor UO_3017 (O_3017,N_25434,N_26943);
nand UO_3018 (O_3018,N_27148,N_29518);
nand UO_3019 (O_3019,N_26222,N_25631);
and UO_3020 (O_3020,N_26432,N_29267);
nor UO_3021 (O_3021,N_27844,N_26047);
nand UO_3022 (O_3022,N_29931,N_25574);
nor UO_3023 (O_3023,N_25216,N_27986);
or UO_3024 (O_3024,N_26209,N_26023);
and UO_3025 (O_3025,N_25367,N_29808);
or UO_3026 (O_3026,N_28512,N_29435);
nor UO_3027 (O_3027,N_29112,N_25908);
and UO_3028 (O_3028,N_29163,N_28658);
and UO_3029 (O_3029,N_27738,N_27257);
xnor UO_3030 (O_3030,N_27068,N_29410);
nor UO_3031 (O_3031,N_25812,N_27235);
nor UO_3032 (O_3032,N_25333,N_28825);
and UO_3033 (O_3033,N_29021,N_25161);
nand UO_3034 (O_3034,N_29676,N_27546);
xor UO_3035 (O_3035,N_29915,N_27392);
nand UO_3036 (O_3036,N_29818,N_26089);
nor UO_3037 (O_3037,N_27447,N_27257);
nor UO_3038 (O_3038,N_28520,N_27630);
nor UO_3039 (O_3039,N_26978,N_26723);
nor UO_3040 (O_3040,N_27533,N_27398);
xnor UO_3041 (O_3041,N_26659,N_26117);
and UO_3042 (O_3042,N_26636,N_26643);
and UO_3043 (O_3043,N_28105,N_25599);
or UO_3044 (O_3044,N_27231,N_25038);
nand UO_3045 (O_3045,N_28458,N_26821);
or UO_3046 (O_3046,N_29828,N_29050);
or UO_3047 (O_3047,N_29303,N_26371);
nand UO_3048 (O_3048,N_26048,N_26021);
or UO_3049 (O_3049,N_25957,N_26660);
or UO_3050 (O_3050,N_25463,N_25164);
nand UO_3051 (O_3051,N_27403,N_26520);
or UO_3052 (O_3052,N_27506,N_26387);
nand UO_3053 (O_3053,N_25517,N_29926);
nor UO_3054 (O_3054,N_25071,N_27227);
nand UO_3055 (O_3055,N_27464,N_28075);
nand UO_3056 (O_3056,N_29265,N_26105);
nand UO_3057 (O_3057,N_27865,N_26706);
nand UO_3058 (O_3058,N_26196,N_29751);
or UO_3059 (O_3059,N_26077,N_29193);
or UO_3060 (O_3060,N_26746,N_25644);
nand UO_3061 (O_3061,N_29439,N_27371);
nand UO_3062 (O_3062,N_29629,N_25527);
nand UO_3063 (O_3063,N_28130,N_26560);
xor UO_3064 (O_3064,N_29960,N_27301);
xnor UO_3065 (O_3065,N_29366,N_27091);
or UO_3066 (O_3066,N_26307,N_26020);
and UO_3067 (O_3067,N_25320,N_28799);
nand UO_3068 (O_3068,N_29068,N_29406);
and UO_3069 (O_3069,N_29759,N_27525);
nor UO_3070 (O_3070,N_27953,N_29556);
xnor UO_3071 (O_3071,N_28953,N_29907);
or UO_3072 (O_3072,N_26915,N_27464);
nand UO_3073 (O_3073,N_29150,N_29138);
or UO_3074 (O_3074,N_25776,N_29638);
or UO_3075 (O_3075,N_27529,N_27171);
or UO_3076 (O_3076,N_27497,N_29738);
and UO_3077 (O_3077,N_25670,N_28707);
nand UO_3078 (O_3078,N_29129,N_29057);
nor UO_3079 (O_3079,N_25913,N_25220);
xnor UO_3080 (O_3080,N_25542,N_27514);
nand UO_3081 (O_3081,N_25311,N_27561);
nand UO_3082 (O_3082,N_29573,N_25608);
nand UO_3083 (O_3083,N_28532,N_29336);
and UO_3084 (O_3084,N_26940,N_26595);
nand UO_3085 (O_3085,N_25897,N_25661);
nand UO_3086 (O_3086,N_25541,N_25125);
or UO_3087 (O_3087,N_26414,N_28207);
nor UO_3088 (O_3088,N_25485,N_29287);
nor UO_3089 (O_3089,N_26263,N_26433);
and UO_3090 (O_3090,N_28884,N_26664);
nor UO_3091 (O_3091,N_25730,N_28349);
nand UO_3092 (O_3092,N_28282,N_25854);
or UO_3093 (O_3093,N_27891,N_25706);
nand UO_3094 (O_3094,N_27721,N_27504);
and UO_3095 (O_3095,N_27438,N_26607);
and UO_3096 (O_3096,N_28772,N_26256);
nor UO_3097 (O_3097,N_26810,N_28352);
nor UO_3098 (O_3098,N_26044,N_26536);
nor UO_3099 (O_3099,N_29769,N_27767);
and UO_3100 (O_3100,N_28213,N_28968);
or UO_3101 (O_3101,N_26914,N_25047);
and UO_3102 (O_3102,N_29403,N_29802);
xor UO_3103 (O_3103,N_28899,N_29346);
and UO_3104 (O_3104,N_29706,N_25980);
and UO_3105 (O_3105,N_29917,N_28794);
or UO_3106 (O_3106,N_25969,N_26199);
or UO_3107 (O_3107,N_26518,N_25393);
and UO_3108 (O_3108,N_28030,N_29593);
nand UO_3109 (O_3109,N_26620,N_26276);
nor UO_3110 (O_3110,N_26437,N_27066);
nand UO_3111 (O_3111,N_27546,N_25251);
and UO_3112 (O_3112,N_28543,N_25100);
or UO_3113 (O_3113,N_28294,N_27096);
or UO_3114 (O_3114,N_28707,N_25301);
and UO_3115 (O_3115,N_29055,N_25679);
and UO_3116 (O_3116,N_28153,N_25425);
and UO_3117 (O_3117,N_29129,N_28591);
and UO_3118 (O_3118,N_27029,N_27057);
or UO_3119 (O_3119,N_27920,N_26419);
nand UO_3120 (O_3120,N_27041,N_27488);
nand UO_3121 (O_3121,N_28687,N_28585);
and UO_3122 (O_3122,N_28503,N_26354);
nor UO_3123 (O_3123,N_26986,N_27188);
nand UO_3124 (O_3124,N_26682,N_27130);
and UO_3125 (O_3125,N_26653,N_28759);
or UO_3126 (O_3126,N_25275,N_26885);
or UO_3127 (O_3127,N_29377,N_25262);
and UO_3128 (O_3128,N_29240,N_29390);
and UO_3129 (O_3129,N_27570,N_28819);
and UO_3130 (O_3130,N_25251,N_27467);
nor UO_3131 (O_3131,N_26013,N_27914);
or UO_3132 (O_3132,N_28251,N_25396);
or UO_3133 (O_3133,N_29898,N_29379);
and UO_3134 (O_3134,N_26215,N_29811);
nor UO_3135 (O_3135,N_29660,N_25224);
nor UO_3136 (O_3136,N_26087,N_26996);
or UO_3137 (O_3137,N_27952,N_28970);
xnor UO_3138 (O_3138,N_26336,N_29525);
nor UO_3139 (O_3139,N_25782,N_29020);
nand UO_3140 (O_3140,N_26297,N_28997);
and UO_3141 (O_3141,N_26250,N_29984);
and UO_3142 (O_3142,N_25867,N_28194);
or UO_3143 (O_3143,N_29148,N_25533);
and UO_3144 (O_3144,N_29690,N_29753);
or UO_3145 (O_3145,N_28375,N_29930);
and UO_3146 (O_3146,N_26198,N_27276);
and UO_3147 (O_3147,N_29635,N_28705);
and UO_3148 (O_3148,N_25727,N_26814);
or UO_3149 (O_3149,N_26127,N_26237);
nand UO_3150 (O_3150,N_29967,N_29364);
nand UO_3151 (O_3151,N_28621,N_28170);
and UO_3152 (O_3152,N_28612,N_25478);
nand UO_3153 (O_3153,N_29854,N_29437);
or UO_3154 (O_3154,N_28075,N_26907);
xnor UO_3155 (O_3155,N_27826,N_25184);
nor UO_3156 (O_3156,N_27967,N_27541);
nor UO_3157 (O_3157,N_28504,N_29798);
xor UO_3158 (O_3158,N_28885,N_27637);
nand UO_3159 (O_3159,N_27172,N_27341);
nand UO_3160 (O_3160,N_25308,N_25574);
nand UO_3161 (O_3161,N_26418,N_27644);
or UO_3162 (O_3162,N_29220,N_27887);
or UO_3163 (O_3163,N_25783,N_26475);
or UO_3164 (O_3164,N_29215,N_27332);
nor UO_3165 (O_3165,N_26745,N_26821);
and UO_3166 (O_3166,N_27923,N_29150);
nor UO_3167 (O_3167,N_27682,N_28554);
xor UO_3168 (O_3168,N_27064,N_28723);
nor UO_3169 (O_3169,N_25224,N_25391);
or UO_3170 (O_3170,N_26285,N_26934);
or UO_3171 (O_3171,N_29012,N_26727);
xnor UO_3172 (O_3172,N_28915,N_25079);
or UO_3173 (O_3173,N_29719,N_29896);
or UO_3174 (O_3174,N_26060,N_29273);
and UO_3175 (O_3175,N_29613,N_28318);
or UO_3176 (O_3176,N_26100,N_27767);
xnor UO_3177 (O_3177,N_27845,N_25816);
nor UO_3178 (O_3178,N_27610,N_27803);
xor UO_3179 (O_3179,N_28078,N_29890);
and UO_3180 (O_3180,N_28466,N_28567);
and UO_3181 (O_3181,N_29789,N_26422);
xnor UO_3182 (O_3182,N_27987,N_27914);
nand UO_3183 (O_3183,N_26878,N_25896);
or UO_3184 (O_3184,N_27367,N_25446);
nand UO_3185 (O_3185,N_27149,N_26410);
nand UO_3186 (O_3186,N_27238,N_29087);
nand UO_3187 (O_3187,N_27529,N_25366);
or UO_3188 (O_3188,N_27563,N_29919);
nor UO_3189 (O_3189,N_27091,N_29834);
or UO_3190 (O_3190,N_29317,N_29471);
nor UO_3191 (O_3191,N_26283,N_27461);
nand UO_3192 (O_3192,N_28335,N_25892);
nor UO_3193 (O_3193,N_27176,N_25596);
xnor UO_3194 (O_3194,N_29307,N_27009);
or UO_3195 (O_3195,N_25820,N_26815);
xor UO_3196 (O_3196,N_27276,N_28170);
nor UO_3197 (O_3197,N_29311,N_27676);
or UO_3198 (O_3198,N_29944,N_26276);
and UO_3199 (O_3199,N_28437,N_27296);
or UO_3200 (O_3200,N_26384,N_26819);
and UO_3201 (O_3201,N_26685,N_25238);
nand UO_3202 (O_3202,N_26622,N_29763);
or UO_3203 (O_3203,N_27056,N_25588);
or UO_3204 (O_3204,N_29651,N_28969);
nand UO_3205 (O_3205,N_26965,N_29039);
or UO_3206 (O_3206,N_27462,N_28425);
nor UO_3207 (O_3207,N_28994,N_26339);
and UO_3208 (O_3208,N_26651,N_28485);
nand UO_3209 (O_3209,N_29781,N_26698);
and UO_3210 (O_3210,N_29070,N_28511);
and UO_3211 (O_3211,N_27682,N_27689);
and UO_3212 (O_3212,N_25143,N_25327);
and UO_3213 (O_3213,N_26532,N_29045);
xnor UO_3214 (O_3214,N_28806,N_26028);
nand UO_3215 (O_3215,N_29697,N_28847);
nor UO_3216 (O_3216,N_27071,N_28070);
nor UO_3217 (O_3217,N_27634,N_26120);
or UO_3218 (O_3218,N_28689,N_25831);
or UO_3219 (O_3219,N_29403,N_26016);
nor UO_3220 (O_3220,N_29122,N_27876);
or UO_3221 (O_3221,N_25524,N_29103);
and UO_3222 (O_3222,N_29706,N_26096);
nor UO_3223 (O_3223,N_26972,N_29857);
or UO_3224 (O_3224,N_29292,N_26029);
and UO_3225 (O_3225,N_29121,N_29568);
and UO_3226 (O_3226,N_26371,N_29094);
nor UO_3227 (O_3227,N_28426,N_28311);
and UO_3228 (O_3228,N_25187,N_29323);
and UO_3229 (O_3229,N_29923,N_27789);
or UO_3230 (O_3230,N_28658,N_26842);
or UO_3231 (O_3231,N_29461,N_28970);
or UO_3232 (O_3232,N_25404,N_25850);
nand UO_3233 (O_3233,N_27733,N_27314);
or UO_3234 (O_3234,N_26927,N_29314);
xnor UO_3235 (O_3235,N_28128,N_27959);
nor UO_3236 (O_3236,N_29589,N_27742);
nand UO_3237 (O_3237,N_28766,N_29781);
nand UO_3238 (O_3238,N_28766,N_25157);
and UO_3239 (O_3239,N_26834,N_29156);
or UO_3240 (O_3240,N_29366,N_28402);
nand UO_3241 (O_3241,N_28678,N_27611);
and UO_3242 (O_3242,N_25312,N_26140);
and UO_3243 (O_3243,N_27178,N_26140);
xor UO_3244 (O_3244,N_28542,N_26361);
nand UO_3245 (O_3245,N_29624,N_28085);
or UO_3246 (O_3246,N_29320,N_26643);
nand UO_3247 (O_3247,N_25953,N_29106);
nor UO_3248 (O_3248,N_26203,N_28736);
and UO_3249 (O_3249,N_27298,N_29901);
and UO_3250 (O_3250,N_25540,N_26376);
nand UO_3251 (O_3251,N_29937,N_29867);
nor UO_3252 (O_3252,N_29235,N_28532);
nor UO_3253 (O_3253,N_29659,N_27737);
nor UO_3254 (O_3254,N_25542,N_26986);
nor UO_3255 (O_3255,N_29317,N_27336);
and UO_3256 (O_3256,N_28675,N_29581);
xor UO_3257 (O_3257,N_26593,N_29223);
nand UO_3258 (O_3258,N_26661,N_25850);
and UO_3259 (O_3259,N_26789,N_26272);
nor UO_3260 (O_3260,N_26910,N_29731);
or UO_3261 (O_3261,N_25992,N_27397);
nand UO_3262 (O_3262,N_29084,N_25476);
nor UO_3263 (O_3263,N_26325,N_25414);
nand UO_3264 (O_3264,N_29157,N_27550);
and UO_3265 (O_3265,N_25147,N_29230);
nand UO_3266 (O_3266,N_27472,N_27132);
nor UO_3267 (O_3267,N_26779,N_25776);
nand UO_3268 (O_3268,N_26485,N_26160);
nand UO_3269 (O_3269,N_25070,N_26988);
xnor UO_3270 (O_3270,N_29785,N_27666);
or UO_3271 (O_3271,N_26436,N_26580);
nand UO_3272 (O_3272,N_28134,N_28737);
nor UO_3273 (O_3273,N_29546,N_26417);
or UO_3274 (O_3274,N_29055,N_26903);
nand UO_3275 (O_3275,N_26180,N_27195);
and UO_3276 (O_3276,N_29137,N_26491);
and UO_3277 (O_3277,N_27643,N_27212);
nand UO_3278 (O_3278,N_26112,N_25727);
and UO_3279 (O_3279,N_29578,N_26604);
nor UO_3280 (O_3280,N_29180,N_26412);
and UO_3281 (O_3281,N_25304,N_27435);
nand UO_3282 (O_3282,N_26175,N_28574);
and UO_3283 (O_3283,N_25298,N_26543);
nor UO_3284 (O_3284,N_27168,N_27582);
nor UO_3285 (O_3285,N_25211,N_27158);
and UO_3286 (O_3286,N_26119,N_27425);
nand UO_3287 (O_3287,N_26396,N_28489);
or UO_3288 (O_3288,N_28263,N_27464);
nand UO_3289 (O_3289,N_29264,N_28024);
or UO_3290 (O_3290,N_27411,N_26492);
nor UO_3291 (O_3291,N_27638,N_29089);
or UO_3292 (O_3292,N_29255,N_29121);
or UO_3293 (O_3293,N_27523,N_28227);
nand UO_3294 (O_3294,N_29801,N_27703);
nor UO_3295 (O_3295,N_28402,N_26361);
and UO_3296 (O_3296,N_29536,N_27633);
and UO_3297 (O_3297,N_29656,N_28503);
or UO_3298 (O_3298,N_29921,N_25493);
nor UO_3299 (O_3299,N_29372,N_28821);
and UO_3300 (O_3300,N_27562,N_28360);
and UO_3301 (O_3301,N_29434,N_27258);
or UO_3302 (O_3302,N_27348,N_27339);
nor UO_3303 (O_3303,N_29760,N_29477);
or UO_3304 (O_3304,N_27978,N_27454);
nand UO_3305 (O_3305,N_28515,N_26193);
nand UO_3306 (O_3306,N_28553,N_26965);
nor UO_3307 (O_3307,N_27444,N_27736);
and UO_3308 (O_3308,N_29982,N_29897);
nand UO_3309 (O_3309,N_28081,N_27675);
nand UO_3310 (O_3310,N_29271,N_26763);
nand UO_3311 (O_3311,N_25419,N_27564);
or UO_3312 (O_3312,N_25110,N_25603);
and UO_3313 (O_3313,N_28673,N_27849);
and UO_3314 (O_3314,N_29035,N_26223);
or UO_3315 (O_3315,N_25787,N_26642);
or UO_3316 (O_3316,N_29842,N_29245);
nand UO_3317 (O_3317,N_25559,N_27964);
or UO_3318 (O_3318,N_29467,N_27737);
or UO_3319 (O_3319,N_25312,N_26482);
nor UO_3320 (O_3320,N_25951,N_29199);
nor UO_3321 (O_3321,N_25563,N_25826);
nand UO_3322 (O_3322,N_26381,N_29913);
nand UO_3323 (O_3323,N_26183,N_28961);
nor UO_3324 (O_3324,N_29464,N_27131);
and UO_3325 (O_3325,N_29466,N_29440);
xnor UO_3326 (O_3326,N_27536,N_26906);
or UO_3327 (O_3327,N_28270,N_26550);
and UO_3328 (O_3328,N_26223,N_28995);
or UO_3329 (O_3329,N_29611,N_27883);
or UO_3330 (O_3330,N_28417,N_27887);
or UO_3331 (O_3331,N_26909,N_28541);
nor UO_3332 (O_3332,N_28314,N_29208);
and UO_3333 (O_3333,N_25923,N_29474);
nor UO_3334 (O_3334,N_27177,N_29756);
nand UO_3335 (O_3335,N_29484,N_27502);
xor UO_3336 (O_3336,N_26387,N_25864);
nor UO_3337 (O_3337,N_27541,N_28359);
or UO_3338 (O_3338,N_28853,N_25084);
and UO_3339 (O_3339,N_29005,N_29487);
nand UO_3340 (O_3340,N_25824,N_26615);
and UO_3341 (O_3341,N_29997,N_27869);
and UO_3342 (O_3342,N_29578,N_25367);
nand UO_3343 (O_3343,N_25455,N_28404);
and UO_3344 (O_3344,N_26779,N_28908);
nor UO_3345 (O_3345,N_26920,N_26336);
nor UO_3346 (O_3346,N_25106,N_25449);
nor UO_3347 (O_3347,N_28975,N_28439);
and UO_3348 (O_3348,N_29232,N_25017);
nor UO_3349 (O_3349,N_25133,N_27826);
and UO_3350 (O_3350,N_25353,N_29741);
and UO_3351 (O_3351,N_27916,N_27453);
nor UO_3352 (O_3352,N_26636,N_26416);
or UO_3353 (O_3353,N_26196,N_27172);
or UO_3354 (O_3354,N_25788,N_26852);
nand UO_3355 (O_3355,N_27490,N_27032);
or UO_3356 (O_3356,N_29211,N_27174);
nand UO_3357 (O_3357,N_27298,N_28062);
nand UO_3358 (O_3358,N_29878,N_29256);
or UO_3359 (O_3359,N_25024,N_28509);
and UO_3360 (O_3360,N_29981,N_27104);
nand UO_3361 (O_3361,N_27856,N_27630);
nor UO_3362 (O_3362,N_28554,N_28413);
and UO_3363 (O_3363,N_26735,N_28618);
and UO_3364 (O_3364,N_25801,N_29181);
and UO_3365 (O_3365,N_26964,N_26588);
or UO_3366 (O_3366,N_25541,N_28209);
or UO_3367 (O_3367,N_27877,N_29255);
nand UO_3368 (O_3368,N_26137,N_28757);
and UO_3369 (O_3369,N_26126,N_27929);
and UO_3370 (O_3370,N_26989,N_26633);
nor UO_3371 (O_3371,N_25570,N_26425);
or UO_3372 (O_3372,N_28397,N_26241);
nand UO_3373 (O_3373,N_27796,N_28628);
and UO_3374 (O_3374,N_27171,N_28463);
xor UO_3375 (O_3375,N_26867,N_25317);
nor UO_3376 (O_3376,N_25189,N_26217);
nand UO_3377 (O_3377,N_26623,N_27569);
nor UO_3378 (O_3378,N_25561,N_29542);
or UO_3379 (O_3379,N_27147,N_29702);
or UO_3380 (O_3380,N_29857,N_28091);
nor UO_3381 (O_3381,N_29406,N_25959);
or UO_3382 (O_3382,N_26360,N_28450);
nand UO_3383 (O_3383,N_28981,N_27046);
xnor UO_3384 (O_3384,N_29829,N_27148);
nand UO_3385 (O_3385,N_29132,N_25794);
nand UO_3386 (O_3386,N_25573,N_29355);
and UO_3387 (O_3387,N_25721,N_28267);
nor UO_3388 (O_3388,N_26079,N_29819);
xor UO_3389 (O_3389,N_25011,N_25908);
nor UO_3390 (O_3390,N_26450,N_26488);
and UO_3391 (O_3391,N_27947,N_29893);
nand UO_3392 (O_3392,N_29203,N_26201);
or UO_3393 (O_3393,N_27639,N_29176);
nor UO_3394 (O_3394,N_28233,N_29914);
and UO_3395 (O_3395,N_29296,N_27951);
xnor UO_3396 (O_3396,N_29225,N_26621);
xnor UO_3397 (O_3397,N_27546,N_26288);
nor UO_3398 (O_3398,N_27801,N_26972);
or UO_3399 (O_3399,N_29337,N_28991);
nand UO_3400 (O_3400,N_27163,N_28001);
nand UO_3401 (O_3401,N_28155,N_27141);
or UO_3402 (O_3402,N_27784,N_26130);
or UO_3403 (O_3403,N_27764,N_25404);
nor UO_3404 (O_3404,N_29175,N_29455);
or UO_3405 (O_3405,N_27062,N_26824);
nor UO_3406 (O_3406,N_25180,N_27807);
nand UO_3407 (O_3407,N_27275,N_29893);
nand UO_3408 (O_3408,N_25613,N_29374);
nand UO_3409 (O_3409,N_27218,N_25540);
and UO_3410 (O_3410,N_28628,N_28107);
nand UO_3411 (O_3411,N_28719,N_25342);
nor UO_3412 (O_3412,N_28529,N_25744);
and UO_3413 (O_3413,N_25097,N_26882);
xor UO_3414 (O_3414,N_29436,N_29361);
nand UO_3415 (O_3415,N_26356,N_25748);
and UO_3416 (O_3416,N_25517,N_27203);
and UO_3417 (O_3417,N_29539,N_25565);
or UO_3418 (O_3418,N_26176,N_27487);
nor UO_3419 (O_3419,N_25246,N_27054);
and UO_3420 (O_3420,N_25176,N_26917);
xor UO_3421 (O_3421,N_29765,N_25671);
or UO_3422 (O_3422,N_29720,N_26194);
or UO_3423 (O_3423,N_26628,N_26096);
nor UO_3424 (O_3424,N_27742,N_25417);
xor UO_3425 (O_3425,N_25458,N_27498);
or UO_3426 (O_3426,N_25571,N_27138);
or UO_3427 (O_3427,N_25351,N_26090);
and UO_3428 (O_3428,N_26855,N_26944);
nand UO_3429 (O_3429,N_26114,N_25442);
xor UO_3430 (O_3430,N_29651,N_26744);
or UO_3431 (O_3431,N_28107,N_26730);
nand UO_3432 (O_3432,N_29522,N_28593);
or UO_3433 (O_3433,N_28409,N_29511);
or UO_3434 (O_3434,N_25341,N_25546);
nor UO_3435 (O_3435,N_26205,N_25518);
or UO_3436 (O_3436,N_25489,N_29793);
nor UO_3437 (O_3437,N_27619,N_27647);
nor UO_3438 (O_3438,N_26971,N_26377);
or UO_3439 (O_3439,N_27798,N_28710);
or UO_3440 (O_3440,N_26515,N_26080);
xnor UO_3441 (O_3441,N_28446,N_28912);
and UO_3442 (O_3442,N_28007,N_25928);
nand UO_3443 (O_3443,N_27627,N_25972);
and UO_3444 (O_3444,N_29345,N_27969);
nand UO_3445 (O_3445,N_29118,N_27123);
and UO_3446 (O_3446,N_28951,N_26762);
nand UO_3447 (O_3447,N_29755,N_29646);
and UO_3448 (O_3448,N_28266,N_25397);
nor UO_3449 (O_3449,N_25478,N_28659);
or UO_3450 (O_3450,N_27527,N_28090);
nor UO_3451 (O_3451,N_26781,N_27794);
nand UO_3452 (O_3452,N_29026,N_28218);
and UO_3453 (O_3453,N_27918,N_27206);
nand UO_3454 (O_3454,N_25211,N_25713);
and UO_3455 (O_3455,N_28168,N_25967);
nand UO_3456 (O_3456,N_26089,N_27320);
nor UO_3457 (O_3457,N_27560,N_26937);
or UO_3458 (O_3458,N_28335,N_29684);
xnor UO_3459 (O_3459,N_28364,N_26834);
nor UO_3460 (O_3460,N_25378,N_25531);
or UO_3461 (O_3461,N_25350,N_29368);
xnor UO_3462 (O_3462,N_27753,N_28142);
xnor UO_3463 (O_3463,N_26505,N_28896);
and UO_3464 (O_3464,N_25779,N_29550);
nand UO_3465 (O_3465,N_26430,N_29419);
xor UO_3466 (O_3466,N_29542,N_29072);
nand UO_3467 (O_3467,N_27916,N_26667);
or UO_3468 (O_3468,N_28213,N_27426);
or UO_3469 (O_3469,N_26634,N_29447);
or UO_3470 (O_3470,N_28639,N_28017);
xnor UO_3471 (O_3471,N_29008,N_25114);
nor UO_3472 (O_3472,N_27969,N_29841);
and UO_3473 (O_3473,N_29196,N_27679);
nand UO_3474 (O_3474,N_25140,N_28494);
nand UO_3475 (O_3475,N_25907,N_27394);
or UO_3476 (O_3476,N_29979,N_28754);
xor UO_3477 (O_3477,N_27238,N_25533);
nor UO_3478 (O_3478,N_26889,N_27117);
nor UO_3479 (O_3479,N_27994,N_25207);
nand UO_3480 (O_3480,N_27928,N_26463);
and UO_3481 (O_3481,N_28886,N_25152);
nor UO_3482 (O_3482,N_28394,N_25418);
nor UO_3483 (O_3483,N_29540,N_27736);
or UO_3484 (O_3484,N_28341,N_27436);
nand UO_3485 (O_3485,N_29004,N_28181);
and UO_3486 (O_3486,N_29429,N_25940);
or UO_3487 (O_3487,N_26689,N_28073);
nand UO_3488 (O_3488,N_25343,N_29704);
or UO_3489 (O_3489,N_28084,N_28109);
and UO_3490 (O_3490,N_25670,N_28612);
xor UO_3491 (O_3491,N_27129,N_25478);
nor UO_3492 (O_3492,N_28842,N_25838);
and UO_3493 (O_3493,N_27856,N_27005);
nor UO_3494 (O_3494,N_25959,N_25825);
nand UO_3495 (O_3495,N_26888,N_29083);
nand UO_3496 (O_3496,N_29067,N_25628);
nand UO_3497 (O_3497,N_28127,N_27422);
nor UO_3498 (O_3498,N_28002,N_28938);
nand UO_3499 (O_3499,N_26775,N_29312);
endmodule