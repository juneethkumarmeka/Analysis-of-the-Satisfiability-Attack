module basic_500_3000_500_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_262,In_382);
nand U1 (N_1,In_238,In_430);
xor U2 (N_2,In_326,In_21);
xnor U3 (N_3,In_154,In_41);
nand U4 (N_4,In_65,In_414);
nand U5 (N_5,In_95,In_441);
and U6 (N_6,In_73,In_255);
and U7 (N_7,In_376,In_274);
xor U8 (N_8,In_481,In_13);
or U9 (N_9,In_102,In_74);
nand U10 (N_10,In_82,In_462);
nand U11 (N_11,In_169,In_84);
or U12 (N_12,In_339,In_19);
and U13 (N_13,In_223,In_325);
nand U14 (N_14,In_439,In_234);
and U15 (N_15,In_69,In_164);
xor U16 (N_16,In_400,In_444);
xnor U17 (N_17,In_307,In_277);
nand U18 (N_18,In_393,In_20);
xnor U19 (N_19,In_147,In_458);
nand U20 (N_20,In_429,In_124);
or U21 (N_21,In_91,In_348);
or U22 (N_22,In_12,In_197);
nand U23 (N_23,In_57,In_293);
xor U24 (N_24,In_346,In_345);
and U25 (N_25,In_297,In_121);
or U26 (N_26,In_296,In_130);
nor U27 (N_27,In_104,In_129);
or U28 (N_28,In_391,In_126);
nor U29 (N_29,In_192,In_39);
nor U30 (N_30,In_202,In_290);
or U31 (N_31,In_99,In_195);
and U32 (N_32,In_407,In_120);
nand U33 (N_33,In_261,In_96);
nor U34 (N_34,In_399,In_493);
nand U35 (N_35,In_236,In_210);
or U36 (N_36,In_272,In_162);
nand U37 (N_37,In_263,In_123);
nand U38 (N_38,In_14,In_50);
nor U39 (N_39,In_118,In_303);
and U40 (N_40,In_253,In_284);
nor U41 (N_41,In_377,In_258);
nand U42 (N_42,In_168,In_231);
nor U43 (N_43,In_16,In_285);
nand U44 (N_44,In_472,In_252);
nand U45 (N_45,In_338,In_219);
and U46 (N_46,In_45,In_352);
nand U47 (N_47,In_54,In_106);
and U48 (N_48,In_358,In_413);
nor U49 (N_49,In_271,In_469);
xnor U50 (N_50,In_101,In_471);
nor U51 (N_51,In_251,In_374);
or U52 (N_52,In_183,In_235);
nand U53 (N_53,In_136,In_283);
nor U54 (N_54,In_454,In_38);
and U55 (N_55,In_435,In_35);
or U56 (N_56,In_5,In_1);
or U57 (N_57,In_330,In_311);
nand U58 (N_58,In_117,In_90);
or U59 (N_59,In_294,In_308);
or U60 (N_60,In_301,In_9);
nand U61 (N_61,In_207,In_83);
nand U62 (N_62,In_89,In_402);
nand U63 (N_63,In_312,In_237);
nand U64 (N_64,In_131,In_476);
and U65 (N_65,In_447,In_81);
nor U66 (N_66,In_289,In_370);
nor U67 (N_67,In_394,In_424);
nand U68 (N_68,In_498,In_63);
or U69 (N_69,In_486,In_221);
nand U70 (N_70,In_317,In_55);
and U71 (N_71,In_386,In_440);
nand U72 (N_72,In_380,In_64);
nor U73 (N_73,In_280,In_178);
or U74 (N_74,In_319,In_482);
nor U75 (N_75,In_436,In_201);
and U76 (N_76,In_176,In_244);
xnor U77 (N_77,In_18,In_52);
and U78 (N_78,In_300,In_229);
nor U79 (N_79,In_480,In_72);
nand U80 (N_80,In_465,In_70);
nor U81 (N_81,In_165,In_298);
and U82 (N_82,In_97,In_29);
nand U83 (N_83,In_492,In_455);
or U84 (N_84,In_372,In_309);
and U85 (N_85,In_58,In_417);
nor U86 (N_86,In_384,In_357);
xnor U87 (N_87,In_7,In_149);
nand U88 (N_88,In_4,In_109);
xnor U89 (N_89,In_321,In_431);
or U90 (N_90,In_204,In_215);
and U91 (N_91,In_107,In_116);
nor U92 (N_92,In_71,In_496);
nor U93 (N_93,In_248,In_420);
nor U94 (N_94,In_410,In_485);
xor U95 (N_95,In_103,In_3);
or U96 (N_96,In_397,In_259);
or U97 (N_97,In_383,In_172);
nor U98 (N_98,In_134,In_278);
nor U99 (N_99,In_239,In_137);
or U100 (N_100,In_310,In_0);
xor U101 (N_101,In_214,In_155);
nor U102 (N_102,In_111,In_190);
and U103 (N_103,In_51,In_22);
nor U104 (N_104,In_142,In_228);
or U105 (N_105,In_443,In_459);
and U106 (N_106,In_257,In_246);
nand U107 (N_107,In_247,In_79);
and U108 (N_108,In_139,In_483);
xor U109 (N_109,In_135,In_334);
or U110 (N_110,In_368,In_464);
or U111 (N_111,In_249,In_23);
nor U112 (N_112,In_203,In_287);
or U113 (N_113,In_187,In_276);
and U114 (N_114,In_404,In_422);
nor U115 (N_115,In_456,In_318);
nor U116 (N_116,In_367,In_32);
or U117 (N_117,In_24,In_359);
nand U118 (N_118,In_491,In_484);
nor U119 (N_119,In_173,In_198);
xnor U120 (N_120,In_418,In_477);
nand U121 (N_121,In_411,In_378);
nand U122 (N_122,In_273,In_451);
and U123 (N_123,In_161,In_389);
xnor U124 (N_124,In_37,In_46);
nor U125 (N_125,In_408,In_344);
xor U126 (N_126,In_396,In_266);
nand U127 (N_127,In_67,In_220);
xnor U128 (N_128,In_113,In_185);
and U129 (N_129,In_353,In_398);
or U130 (N_130,In_405,In_85);
nor U131 (N_131,In_421,In_419);
and U132 (N_132,In_473,In_369);
xnor U133 (N_133,In_66,In_227);
and U134 (N_134,In_256,In_158);
xor U135 (N_135,In_145,In_475);
or U136 (N_136,In_150,In_94);
and U137 (N_137,In_365,In_241);
xor U138 (N_138,In_2,In_180);
nor U139 (N_139,In_270,In_445);
xor U140 (N_140,In_392,In_213);
or U141 (N_141,In_25,In_387);
nor U142 (N_142,In_371,In_434);
nor U143 (N_143,In_49,In_499);
nand U144 (N_144,In_80,In_163);
or U145 (N_145,In_160,In_98);
xnor U146 (N_146,In_157,In_390);
and U147 (N_147,In_152,In_138);
xnor U148 (N_148,In_487,In_110);
and U149 (N_149,In_243,In_115);
and U150 (N_150,In_184,In_175);
xor U151 (N_151,In_291,In_31);
nand U152 (N_152,In_450,In_416);
xor U153 (N_153,In_363,In_260);
and U154 (N_154,In_304,In_196);
nand U155 (N_155,In_224,In_395);
or U156 (N_156,In_93,In_448);
or U157 (N_157,In_490,In_488);
nand U158 (N_158,In_206,In_179);
xor U159 (N_159,In_43,In_170);
or U160 (N_160,In_17,In_375);
and U161 (N_161,In_36,In_267);
nor U162 (N_162,In_132,In_406);
nand U163 (N_163,In_356,In_225);
xor U164 (N_164,In_62,In_119);
nand U165 (N_165,In_211,In_342);
xor U166 (N_166,In_30,In_432);
nand U167 (N_167,In_320,In_86);
xnor U168 (N_168,In_331,In_388);
nand U169 (N_169,In_34,In_381);
nor U170 (N_170,In_379,In_460);
xnor U171 (N_171,In_279,In_474);
or U172 (N_172,In_327,In_423);
xnor U173 (N_173,In_350,In_347);
nand U174 (N_174,In_230,In_100);
nand U175 (N_175,In_114,In_478);
nand U176 (N_176,In_306,In_299);
xor U177 (N_177,In_452,In_105);
nor U178 (N_178,In_415,In_362);
and U179 (N_179,In_28,In_281);
nand U180 (N_180,In_186,In_15);
nand U181 (N_181,In_193,In_87);
nor U182 (N_182,In_288,In_122);
and U183 (N_183,In_153,In_323);
or U184 (N_184,In_181,In_442);
or U185 (N_185,In_470,In_302);
xor U186 (N_186,In_446,In_437);
nor U187 (N_187,In_254,In_305);
or U188 (N_188,In_159,In_76);
and U189 (N_189,In_316,In_112);
xor U190 (N_190,In_133,In_328);
nor U191 (N_191,In_194,In_292);
xnor U192 (N_192,In_68,In_453);
nand U193 (N_193,In_75,In_412);
and U194 (N_194,In_205,In_269);
xor U195 (N_195,In_264,In_212);
or U196 (N_196,In_322,In_240);
nor U197 (N_197,In_265,In_143);
and U198 (N_198,In_33,In_92);
nor U199 (N_199,In_218,In_324);
and U200 (N_200,In_140,In_349);
nor U201 (N_201,In_141,In_275);
nand U202 (N_202,In_385,In_341);
nand U203 (N_203,In_315,In_189);
nor U204 (N_204,In_127,In_242);
xnor U205 (N_205,In_336,In_335);
nand U206 (N_206,In_401,In_332);
and U207 (N_207,In_286,In_360);
nor U208 (N_208,In_427,In_182);
nor U209 (N_209,In_355,In_495);
and U210 (N_210,In_282,In_199);
and U211 (N_211,In_354,In_361);
nor U212 (N_212,In_148,In_177);
or U213 (N_213,In_48,In_438);
and U214 (N_214,In_366,In_216);
nor U215 (N_215,In_295,In_425);
or U216 (N_216,In_60,In_494);
xnor U217 (N_217,In_208,In_171);
nand U218 (N_218,In_466,In_428);
nand U219 (N_219,In_167,In_222);
or U220 (N_220,In_226,In_497);
xnor U221 (N_221,In_151,In_373);
xnor U222 (N_222,In_40,In_56);
and U223 (N_223,In_10,In_461);
and U224 (N_224,In_245,In_191);
or U225 (N_225,In_433,In_166);
and U226 (N_226,In_268,In_314);
xor U227 (N_227,In_449,In_8);
xor U228 (N_228,In_146,In_463);
nor U229 (N_229,In_313,In_78);
or U230 (N_230,In_26,In_364);
and U231 (N_231,In_53,In_489);
nor U232 (N_232,In_467,In_340);
nand U233 (N_233,In_108,In_217);
nor U234 (N_234,In_6,In_351);
nor U235 (N_235,In_403,In_209);
nor U236 (N_236,In_11,In_232);
nor U237 (N_237,In_329,In_426);
and U238 (N_238,In_44,In_174);
or U239 (N_239,In_125,In_47);
or U240 (N_240,In_59,In_128);
and U241 (N_241,In_42,In_27);
nand U242 (N_242,In_343,In_457);
nor U243 (N_243,In_333,In_144);
nor U244 (N_244,In_250,In_156);
nand U245 (N_245,In_200,In_409);
xnor U246 (N_246,In_188,In_337);
nand U247 (N_247,In_88,In_61);
nand U248 (N_248,In_77,In_479);
nor U249 (N_249,In_233,In_468);
nand U250 (N_250,In_454,In_133);
or U251 (N_251,In_496,In_85);
and U252 (N_252,In_279,In_89);
or U253 (N_253,In_354,In_138);
nand U254 (N_254,In_435,In_492);
or U255 (N_255,In_2,In_344);
and U256 (N_256,In_275,In_133);
or U257 (N_257,In_404,In_247);
or U258 (N_258,In_183,In_131);
nor U259 (N_259,In_452,In_171);
and U260 (N_260,In_329,In_373);
nor U261 (N_261,In_348,In_287);
and U262 (N_262,In_477,In_127);
nor U263 (N_263,In_323,In_0);
xor U264 (N_264,In_227,In_455);
or U265 (N_265,In_120,In_194);
nor U266 (N_266,In_263,In_94);
xnor U267 (N_267,In_187,In_493);
xnor U268 (N_268,In_345,In_321);
xnor U269 (N_269,In_231,In_22);
xor U270 (N_270,In_37,In_135);
xor U271 (N_271,In_27,In_141);
xor U272 (N_272,In_327,In_495);
nor U273 (N_273,In_457,In_209);
nand U274 (N_274,In_91,In_440);
and U275 (N_275,In_146,In_379);
or U276 (N_276,In_107,In_355);
and U277 (N_277,In_134,In_256);
nor U278 (N_278,In_147,In_382);
xnor U279 (N_279,In_128,In_251);
nand U280 (N_280,In_223,In_33);
nor U281 (N_281,In_36,In_12);
or U282 (N_282,In_33,In_230);
xnor U283 (N_283,In_122,In_404);
and U284 (N_284,In_463,In_64);
xor U285 (N_285,In_207,In_359);
nand U286 (N_286,In_111,In_169);
and U287 (N_287,In_443,In_286);
nor U288 (N_288,In_203,In_304);
nand U289 (N_289,In_296,In_252);
xor U290 (N_290,In_148,In_133);
nand U291 (N_291,In_404,In_237);
nand U292 (N_292,In_326,In_122);
or U293 (N_293,In_301,In_32);
nor U294 (N_294,In_319,In_145);
nand U295 (N_295,In_443,In_293);
xnor U296 (N_296,In_392,In_467);
nor U297 (N_297,In_220,In_75);
nand U298 (N_298,In_181,In_367);
or U299 (N_299,In_491,In_239);
or U300 (N_300,In_289,In_66);
nor U301 (N_301,In_128,In_476);
and U302 (N_302,In_424,In_374);
nand U303 (N_303,In_388,In_136);
and U304 (N_304,In_255,In_35);
or U305 (N_305,In_290,In_101);
or U306 (N_306,In_76,In_352);
nor U307 (N_307,In_307,In_212);
xor U308 (N_308,In_316,In_484);
or U309 (N_309,In_161,In_369);
xor U310 (N_310,In_290,In_31);
nor U311 (N_311,In_330,In_17);
xor U312 (N_312,In_462,In_50);
nand U313 (N_313,In_195,In_328);
and U314 (N_314,In_98,In_181);
and U315 (N_315,In_493,In_247);
nor U316 (N_316,In_369,In_144);
nand U317 (N_317,In_134,In_96);
nor U318 (N_318,In_409,In_147);
xnor U319 (N_319,In_3,In_51);
nand U320 (N_320,In_122,In_287);
nand U321 (N_321,In_198,In_111);
nor U322 (N_322,In_316,In_349);
nor U323 (N_323,In_90,In_195);
or U324 (N_324,In_318,In_295);
nor U325 (N_325,In_288,In_371);
xor U326 (N_326,In_233,In_62);
and U327 (N_327,In_338,In_20);
and U328 (N_328,In_229,In_155);
or U329 (N_329,In_421,In_433);
and U330 (N_330,In_284,In_412);
nand U331 (N_331,In_74,In_442);
or U332 (N_332,In_249,In_448);
or U333 (N_333,In_92,In_306);
nor U334 (N_334,In_137,In_346);
nor U335 (N_335,In_290,In_105);
or U336 (N_336,In_440,In_453);
nor U337 (N_337,In_380,In_235);
nand U338 (N_338,In_283,In_134);
or U339 (N_339,In_345,In_435);
nand U340 (N_340,In_363,In_252);
and U341 (N_341,In_396,In_200);
nand U342 (N_342,In_146,In_96);
xnor U343 (N_343,In_25,In_49);
xnor U344 (N_344,In_50,In_174);
nor U345 (N_345,In_399,In_192);
and U346 (N_346,In_441,In_188);
and U347 (N_347,In_158,In_412);
nor U348 (N_348,In_232,In_99);
nor U349 (N_349,In_153,In_401);
or U350 (N_350,In_346,In_350);
or U351 (N_351,In_282,In_266);
and U352 (N_352,In_425,In_40);
and U353 (N_353,In_301,In_33);
nand U354 (N_354,In_372,In_180);
nand U355 (N_355,In_231,In_483);
xor U356 (N_356,In_473,In_459);
and U357 (N_357,In_423,In_476);
xor U358 (N_358,In_366,In_300);
nor U359 (N_359,In_169,In_487);
nor U360 (N_360,In_402,In_218);
xor U361 (N_361,In_194,In_73);
nor U362 (N_362,In_461,In_51);
nor U363 (N_363,In_49,In_346);
and U364 (N_364,In_360,In_425);
xnor U365 (N_365,In_20,In_385);
nor U366 (N_366,In_183,In_426);
nand U367 (N_367,In_213,In_464);
nand U368 (N_368,In_195,In_66);
nor U369 (N_369,In_51,In_377);
or U370 (N_370,In_463,In_488);
nor U371 (N_371,In_367,In_363);
nor U372 (N_372,In_429,In_40);
nand U373 (N_373,In_292,In_458);
xor U374 (N_374,In_475,In_304);
nand U375 (N_375,In_137,In_306);
xnor U376 (N_376,In_412,In_450);
and U377 (N_377,In_10,In_121);
nor U378 (N_378,In_43,In_142);
xnor U379 (N_379,In_161,In_383);
xor U380 (N_380,In_15,In_132);
or U381 (N_381,In_48,In_312);
nor U382 (N_382,In_5,In_441);
xnor U383 (N_383,In_162,In_114);
and U384 (N_384,In_247,In_68);
and U385 (N_385,In_166,In_109);
nand U386 (N_386,In_252,In_311);
or U387 (N_387,In_173,In_362);
nand U388 (N_388,In_234,In_56);
or U389 (N_389,In_294,In_95);
or U390 (N_390,In_401,In_248);
and U391 (N_391,In_273,In_377);
and U392 (N_392,In_321,In_148);
or U393 (N_393,In_0,In_340);
or U394 (N_394,In_21,In_175);
nand U395 (N_395,In_349,In_152);
nor U396 (N_396,In_307,In_358);
xor U397 (N_397,In_189,In_303);
xor U398 (N_398,In_461,In_30);
nand U399 (N_399,In_21,In_212);
xor U400 (N_400,In_256,In_82);
and U401 (N_401,In_73,In_132);
or U402 (N_402,In_215,In_69);
and U403 (N_403,In_369,In_314);
nor U404 (N_404,In_473,In_355);
nand U405 (N_405,In_294,In_448);
or U406 (N_406,In_120,In_393);
and U407 (N_407,In_146,In_209);
and U408 (N_408,In_481,In_462);
or U409 (N_409,In_424,In_485);
nor U410 (N_410,In_352,In_181);
and U411 (N_411,In_234,In_448);
and U412 (N_412,In_206,In_119);
xnor U413 (N_413,In_436,In_422);
and U414 (N_414,In_200,In_99);
and U415 (N_415,In_48,In_487);
xor U416 (N_416,In_91,In_243);
xor U417 (N_417,In_409,In_325);
or U418 (N_418,In_428,In_444);
nor U419 (N_419,In_320,In_422);
and U420 (N_420,In_381,In_296);
or U421 (N_421,In_413,In_349);
nand U422 (N_422,In_41,In_200);
or U423 (N_423,In_64,In_119);
and U424 (N_424,In_279,In_175);
nand U425 (N_425,In_332,In_243);
nor U426 (N_426,In_400,In_470);
nor U427 (N_427,In_16,In_228);
nor U428 (N_428,In_344,In_255);
or U429 (N_429,In_496,In_246);
and U430 (N_430,In_462,In_385);
or U431 (N_431,In_484,In_421);
nor U432 (N_432,In_378,In_288);
nand U433 (N_433,In_265,In_183);
and U434 (N_434,In_244,In_296);
and U435 (N_435,In_415,In_280);
xor U436 (N_436,In_209,In_241);
nor U437 (N_437,In_12,In_181);
nor U438 (N_438,In_420,In_484);
xnor U439 (N_439,In_189,In_174);
and U440 (N_440,In_270,In_198);
nand U441 (N_441,In_138,In_393);
xnor U442 (N_442,In_117,In_77);
nand U443 (N_443,In_10,In_169);
and U444 (N_444,In_176,In_202);
nor U445 (N_445,In_492,In_374);
and U446 (N_446,In_4,In_71);
xor U447 (N_447,In_281,In_309);
nor U448 (N_448,In_225,In_49);
nand U449 (N_449,In_219,In_122);
and U450 (N_450,In_329,In_139);
nand U451 (N_451,In_470,In_20);
xor U452 (N_452,In_255,In_193);
and U453 (N_453,In_492,In_368);
or U454 (N_454,In_325,In_436);
nand U455 (N_455,In_204,In_265);
or U456 (N_456,In_470,In_298);
and U457 (N_457,In_430,In_321);
and U458 (N_458,In_76,In_188);
and U459 (N_459,In_191,In_125);
nor U460 (N_460,In_16,In_382);
xnor U461 (N_461,In_9,In_113);
and U462 (N_462,In_10,In_42);
or U463 (N_463,In_79,In_350);
nor U464 (N_464,In_85,In_497);
nor U465 (N_465,In_366,In_38);
xnor U466 (N_466,In_261,In_209);
xnor U467 (N_467,In_23,In_7);
or U468 (N_468,In_367,In_88);
nand U469 (N_469,In_280,In_455);
nand U470 (N_470,In_490,In_271);
nor U471 (N_471,In_339,In_160);
xnor U472 (N_472,In_49,In_429);
nand U473 (N_473,In_133,In_77);
nor U474 (N_474,In_444,In_322);
nand U475 (N_475,In_477,In_190);
and U476 (N_476,In_245,In_246);
nor U477 (N_477,In_322,In_17);
or U478 (N_478,In_152,In_496);
or U479 (N_479,In_225,In_29);
and U480 (N_480,In_171,In_250);
nand U481 (N_481,In_389,In_378);
and U482 (N_482,In_387,In_227);
nor U483 (N_483,In_31,In_332);
or U484 (N_484,In_273,In_189);
or U485 (N_485,In_479,In_256);
or U486 (N_486,In_64,In_332);
xor U487 (N_487,In_347,In_132);
nand U488 (N_488,In_357,In_99);
and U489 (N_489,In_247,In_300);
xor U490 (N_490,In_169,In_35);
or U491 (N_491,In_327,In_421);
or U492 (N_492,In_140,In_434);
nand U493 (N_493,In_197,In_482);
and U494 (N_494,In_364,In_240);
or U495 (N_495,In_176,In_207);
and U496 (N_496,In_93,In_426);
xor U497 (N_497,In_363,In_459);
and U498 (N_498,In_374,In_253);
and U499 (N_499,In_134,In_392);
or U500 (N_500,In_431,In_101);
nor U501 (N_501,In_365,In_375);
and U502 (N_502,In_107,In_406);
or U503 (N_503,In_447,In_349);
nand U504 (N_504,In_34,In_162);
nand U505 (N_505,In_440,In_304);
and U506 (N_506,In_89,In_433);
xnor U507 (N_507,In_363,In_250);
or U508 (N_508,In_178,In_305);
nand U509 (N_509,In_220,In_360);
or U510 (N_510,In_317,In_190);
and U511 (N_511,In_297,In_211);
or U512 (N_512,In_364,In_214);
and U513 (N_513,In_10,In_391);
nor U514 (N_514,In_112,In_164);
or U515 (N_515,In_176,In_367);
or U516 (N_516,In_32,In_67);
xnor U517 (N_517,In_132,In_109);
or U518 (N_518,In_341,In_456);
xor U519 (N_519,In_156,In_149);
and U520 (N_520,In_81,In_367);
nand U521 (N_521,In_376,In_115);
nor U522 (N_522,In_485,In_368);
and U523 (N_523,In_7,In_312);
nor U524 (N_524,In_408,In_399);
xor U525 (N_525,In_383,In_140);
xor U526 (N_526,In_326,In_194);
nand U527 (N_527,In_410,In_374);
or U528 (N_528,In_494,In_134);
or U529 (N_529,In_395,In_32);
nor U530 (N_530,In_465,In_264);
xnor U531 (N_531,In_464,In_293);
xor U532 (N_532,In_364,In_145);
or U533 (N_533,In_369,In_139);
and U534 (N_534,In_46,In_108);
nor U535 (N_535,In_2,In_414);
or U536 (N_536,In_64,In_101);
xor U537 (N_537,In_269,In_116);
or U538 (N_538,In_359,In_495);
or U539 (N_539,In_96,In_353);
xor U540 (N_540,In_410,In_5);
xnor U541 (N_541,In_383,In_199);
nor U542 (N_542,In_336,In_427);
nor U543 (N_543,In_0,In_142);
xnor U544 (N_544,In_15,In_417);
or U545 (N_545,In_119,In_34);
nand U546 (N_546,In_136,In_183);
xnor U547 (N_547,In_436,In_91);
and U548 (N_548,In_321,In_106);
nand U549 (N_549,In_459,In_185);
nor U550 (N_550,In_267,In_328);
nor U551 (N_551,In_388,In_52);
xnor U552 (N_552,In_131,In_450);
xnor U553 (N_553,In_446,In_125);
xor U554 (N_554,In_354,In_263);
xnor U555 (N_555,In_54,In_7);
and U556 (N_556,In_241,In_92);
xnor U557 (N_557,In_79,In_421);
or U558 (N_558,In_489,In_360);
nand U559 (N_559,In_165,In_345);
nor U560 (N_560,In_197,In_268);
and U561 (N_561,In_276,In_196);
xor U562 (N_562,In_443,In_358);
and U563 (N_563,In_270,In_338);
or U564 (N_564,In_124,In_152);
nor U565 (N_565,In_5,In_172);
or U566 (N_566,In_422,In_21);
or U567 (N_567,In_439,In_491);
and U568 (N_568,In_464,In_267);
and U569 (N_569,In_308,In_54);
xnor U570 (N_570,In_66,In_439);
nand U571 (N_571,In_35,In_199);
xor U572 (N_572,In_331,In_238);
nand U573 (N_573,In_221,In_101);
or U574 (N_574,In_74,In_494);
or U575 (N_575,In_312,In_468);
or U576 (N_576,In_219,In_91);
or U577 (N_577,In_346,In_318);
xnor U578 (N_578,In_178,In_345);
xnor U579 (N_579,In_207,In_418);
nor U580 (N_580,In_238,In_42);
or U581 (N_581,In_144,In_466);
nand U582 (N_582,In_496,In_353);
nand U583 (N_583,In_120,In_214);
xor U584 (N_584,In_70,In_142);
nand U585 (N_585,In_219,In_479);
nor U586 (N_586,In_287,In_153);
and U587 (N_587,In_28,In_349);
or U588 (N_588,In_137,In_148);
nor U589 (N_589,In_315,In_21);
nand U590 (N_590,In_388,In_362);
xnor U591 (N_591,In_26,In_66);
nor U592 (N_592,In_169,In_158);
and U593 (N_593,In_37,In_483);
xnor U594 (N_594,In_313,In_256);
or U595 (N_595,In_492,In_196);
or U596 (N_596,In_492,In_456);
nor U597 (N_597,In_499,In_24);
or U598 (N_598,In_50,In_90);
xnor U599 (N_599,In_276,In_169);
xnor U600 (N_600,N_183,N_391);
nand U601 (N_601,N_203,N_499);
nor U602 (N_602,N_558,N_540);
nor U603 (N_603,N_393,N_582);
xor U604 (N_604,N_416,N_563);
or U605 (N_605,N_147,N_326);
or U606 (N_606,N_265,N_418);
nand U607 (N_607,N_139,N_2);
or U608 (N_608,N_21,N_160);
xnor U609 (N_609,N_246,N_569);
xor U610 (N_610,N_306,N_439);
xor U611 (N_611,N_89,N_532);
nor U612 (N_612,N_130,N_87);
and U613 (N_613,N_403,N_599);
or U614 (N_614,N_457,N_320);
nor U615 (N_615,N_465,N_145);
xor U616 (N_616,N_433,N_374);
nor U617 (N_617,N_544,N_519);
and U618 (N_618,N_311,N_9);
nand U619 (N_619,N_435,N_204);
xor U620 (N_620,N_524,N_193);
nor U621 (N_621,N_76,N_578);
xor U622 (N_622,N_413,N_95);
xor U623 (N_623,N_502,N_564);
and U624 (N_624,N_53,N_247);
nor U625 (N_625,N_297,N_395);
nand U626 (N_626,N_31,N_192);
nor U627 (N_627,N_547,N_188);
xor U628 (N_628,N_267,N_245);
nand U629 (N_629,N_79,N_74);
or U630 (N_630,N_186,N_383);
or U631 (N_631,N_535,N_179);
nor U632 (N_632,N_64,N_234);
or U633 (N_633,N_423,N_560);
and U634 (N_634,N_48,N_241);
nand U635 (N_635,N_440,N_555);
nor U636 (N_636,N_18,N_200);
xor U637 (N_637,N_460,N_355);
xnor U638 (N_638,N_27,N_47);
or U639 (N_639,N_119,N_574);
or U640 (N_640,N_51,N_286);
xor U641 (N_641,N_511,N_288);
and U642 (N_642,N_552,N_135);
xnor U643 (N_643,N_581,N_436);
xnor U644 (N_644,N_597,N_128);
xor U645 (N_645,N_349,N_154);
and U646 (N_646,N_410,N_152);
or U647 (N_647,N_93,N_454);
or U648 (N_648,N_105,N_464);
and U649 (N_649,N_75,N_127);
or U650 (N_650,N_103,N_68);
nor U651 (N_651,N_591,N_120);
or U652 (N_652,N_449,N_42);
xnor U653 (N_653,N_224,N_59);
xnor U654 (N_654,N_8,N_61);
or U655 (N_655,N_308,N_168);
nor U656 (N_656,N_447,N_55);
nor U657 (N_657,N_507,N_111);
and U658 (N_658,N_253,N_453);
or U659 (N_659,N_594,N_376);
and U660 (N_660,N_57,N_536);
xor U661 (N_661,N_323,N_144);
or U662 (N_662,N_142,N_116);
nand U663 (N_663,N_561,N_533);
nand U664 (N_664,N_437,N_390);
xor U665 (N_665,N_573,N_271);
nand U666 (N_666,N_104,N_136);
nor U667 (N_667,N_406,N_585);
and U668 (N_668,N_595,N_377);
or U669 (N_669,N_178,N_404);
and U670 (N_670,N_41,N_263);
nor U671 (N_671,N_505,N_518);
nor U672 (N_672,N_516,N_209);
xnor U673 (N_673,N_463,N_314);
or U674 (N_674,N_356,N_24);
or U675 (N_675,N_327,N_228);
nor U676 (N_676,N_493,N_161);
nor U677 (N_677,N_443,N_25);
nor U678 (N_678,N_69,N_83);
xor U679 (N_679,N_233,N_239);
and U680 (N_680,N_92,N_114);
nand U681 (N_681,N_261,N_7);
or U682 (N_682,N_23,N_113);
xor U683 (N_683,N_219,N_295);
and U684 (N_684,N_354,N_19);
nand U685 (N_685,N_227,N_254);
nand U686 (N_686,N_210,N_415);
nor U687 (N_687,N_137,N_132);
or U688 (N_688,N_14,N_251);
and U689 (N_689,N_347,N_473);
or U690 (N_690,N_419,N_361);
nor U691 (N_691,N_77,N_469);
nor U692 (N_692,N_283,N_36);
nor U693 (N_693,N_548,N_369);
xnor U694 (N_694,N_151,N_387);
xor U695 (N_695,N_316,N_1);
or U696 (N_696,N_198,N_50);
xnor U697 (N_697,N_225,N_273);
nand U698 (N_698,N_513,N_72);
nor U699 (N_699,N_22,N_334);
xor U700 (N_700,N_495,N_501);
or U701 (N_701,N_452,N_315);
nor U702 (N_702,N_371,N_335);
nor U703 (N_703,N_54,N_546);
xnor U704 (N_704,N_397,N_264);
or U705 (N_705,N_166,N_551);
nor U706 (N_706,N_545,N_444);
nand U707 (N_707,N_214,N_509);
nor U708 (N_708,N_515,N_385);
or U709 (N_709,N_71,N_353);
nor U710 (N_710,N_290,N_12);
or U711 (N_711,N_141,N_49);
nor U712 (N_712,N_90,N_205);
or U713 (N_713,N_80,N_63);
or U714 (N_714,N_39,N_541);
nor U715 (N_715,N_429,N_34);
nand U716 (N_716,N_478,N_133);
or U717 (N_717,N_182,N_592);
or U718 (N_718,N_207,N_458);
or U719 (N_719,N_217,N_73);
xnor U720 (N_720,N_222,N_466);
nand U721 (N_721,N_62,N_490);
and U722 (N_722,N_520,N_242);
and U723 (N_723,N_375,N_474);
or U724 (N_724,N_521,N_483);
xor U725 (N_725,N_481,N_522);
xor U726 (N_726,N_13,N_324);
or U727 (N_727,N_331,N_567);
nor U728 (N_728,N_456,N_26);
and U729 (N_729,N_579,N_257);
xnor U730 (N_730,N_322,N_468);
xor U731 (N_731,N_216,N_17);
nor U732 (N_732,N_475,N_528);
nor U733 (N_733,N_538,N_367);
xnor U734 (N_734,N_379,N_85);
or U735 (N_735,N_46,N_235);
or U736 (N_736,N_184,N_492);
xor U737 (N_737,N_388,N_40);
nand U738 (N_738,N_302,N_471);
xor U739 (N_739,N_148,N_339);
xnor U740 (N_740,N_243,N_30);
nor U741 (N_741,N_523,N_576);
nand U742 (N_742,N_352,N_303);
or U743 (N_743,N_291,N_319);
or U744 (N_744,N_206,N_176);
and U745 (N_745,N_292,N_459);
or U746 (N_746,N_174,N_332);
nand U747 (N_747,N_351,N_328);
or U748 (N_748,N_67,N_15);
nand U749 (N_749,N_96,N_70);
nand U750 (N_750,N_195,N_212);
and U751 (N_751,N_321,N_190);
nand U752 (N_752,N_58,N_534);
and U753 (N_753,N_577,N_425);
and U754 (N_754,N_220,N_525);
and U755 (N_755,N_398,N_175);
or U756 (N_756,N_537,N_318);
nand U757 (N_757,N_421,N_260);
or U758 (N_758,N_81,N_237);
xor U759 (N_759,N_262,N_287);
nor U760 (N_760,N_97,N_543);
nand U761 (N_761,N_236,N_572);
nor U762 (N_762,N_238,N_294);
nand U763 (N_763,N_301,N_268);
and U764 (N_764,N_299,N_78);
and U765 (N_765,N_112,N_550);
nand U766 (N_766,N_480,N_244);
nor U767 (N_767,N_401,N_252);
xor U768 (N_768,N_0,N_442);
and U769 (N_769,N_357,N_35);
or U770 (N_770,N_562,N_110);
and U771 (N_771,N_337,N_146);
and U772 (N_772,N_100,N_280);
xor U773 (N_773,N_211,N_554);
and U774 (N_774,N_125,N_424);
or U775 (N_775,N_530,N_317);
and U776 (N_776,N_169,N_358);
or U777 (N_777,N_503,N_88);
nor U778 (N_778,N_117,N_307);
and U779 (N_779,N_402,N_341);
nand U780 (N_780,N_66,N_52);
xnor U781 (N_781,N_10,N_431);
and U782 (N_782,N_414,N_191);
nand U783 (N_783,N_427,N_434);
nor U784 (N_784,N_197,N_381);
xnor U785 (N_785,N_86,N_298);
or U786 (N_786,N_472,N_106);
xnor U787 (N_787,N_4,N_304);
xor U788 (N_788,N_494,N_138);
xor U789 (N_789,N_187,N_417);
nor U790 (N_790,N_226,N_173);
xor U791 (N_791,N_181,N_514);
nand U792 (N_792,N_539,N_568);
nor U793 (N_793,N_420,N_428);
or U794 (N_794,N_156,N_270);
xor U795 (N_795,N_272,N_486);
nand U796 (N_796,N_149,N_201);
and U797 (N_797,N_158,N_409);
xor U798 (N_798,N_504,N_279);
nand U799 (N_799,N_134,N_218);
xor U800 (N_800,N_43,N_422);
or U801 (N_801,N_467,N_556);
nor U802 (N_802,N_249,N_170);
nand U803 (N_803,N_445,N_412);
and U804 (N_804,N_529,N_510);
nand U805 (N_805,N_296,N_360);
nand U806 (N_806,N_250,N_482);
xnor U807 (N_807,N_60,N_359);
and U808 (N_808,N_99,N_259);
xnor U809 (N_809,N_598,N_194);
xor U810 (N_810,N_373,N_5);
nor U811 (N_811,N_571,N_150);
and U812 (N_812,N_549,N_98);
nand U813 (N_813,N_284,N_345);
or U814 (N_814,N_258,N_312);
or U815 (N_815,N_348,N_94);
nor U816 (N_816,N_285,N_407);
nand U817 (N_817,N_343,N_329);
or U818 (N_818,N_386,N_56);
nor U819 (N_819,N_338,N_340);
or U820 (N_820,N_140,N_196);
and U821 (N_821,N_432,N_587);
and U822 (N_822,N_44,N_526);
and U823 (N_823,N_350,N_248);
nand U824 (N_824,N_570,N_430);
nand U825 (N_825,N_131,N_155);
xor U826 (N_826,N_165,N_282);
xnor U827 (N_827,N_461,N_124);
and U828 (N_828,N_115,N_487);
and U829 (N_829,N_313,N_221);
nor U830 (N_830,N_37,N_500);
nor U831 (N_831,N_336,N_129);
nand U832 (N_832,N_531,N_91);
xnor U833 (N_833,N_333,N_185);
or U834 (N_834,N_394,N_450);
nand U835 (N_835,N_484,N_365);
xnor U836 (N_836,N_559,N_202);
nand U837 (N_837,N_363,N_274);
and U838 (N_838,N_344,N_389);
nor U839 (N_839,N_16,N_256);
nor U840 (N_840,N_384,N_527);
xor U841 (N_841,N_584,N_84);
xor U842 (N_842,N_588,N_300);
nand U843 (N_843,N_590,N_305);
nor U844 (N_844,N_45,N_122);
or U845 (N_845,N_266,N_215);
nand U846 (N_846,N_28,N_230);
nand U847 (N_847,N_489,N_189);
nor U848 (N_848,N_309,N_38);
or U849 (N_849,N_82,N_479);
nor U850 (N_850,N_172,N_566);
or U851 (N_851,N_372,N_157);
and U852 (N_852,N_153,N_293);
or U853 (N_853,N_396,N_485);
nand U854 (N_854,N_380,N_405);
nor U855 (N_855,N_593,N_232);
nor U856 (N_856,N_400,N_278);
nor U857 (N_857,N_330,N_240);
nand U858 (N_858,N_506,N_364);
nor U859 (N_859,N_143,N_596);
and U860 (N_860,N_426,N_11);
nand U861 (N_861,N_476,N_368);
nor U862 (N_862,N_448,N_65);
nand U863 (N_863,N_496,N_277);
xnor U864 (N_864,N_177,N_446);
nand U865 (N_865,N_441,N_107);
and U866 (N_866,N_3,N_346);
and U867 (N_867,N_382,N_508);
nand U868 (N_868,N_163,N_101);
xnor U869 (N_869,N_512,N_275);
and U870 (N_870,N_164,N_118);
xnor U871 (N_871,N_477,N_281);
nand U872 (N_872,N_159,N_325);
nor U873 (N_873,N_229,N_517);
or U874 (N_874,N_451,N_370);
or U875 (N_875,N_378,N_123);
nand U876 (N_876,N_102,N_589);
nand U877 (N_877,N_32,N_408);
nor U878 (N_878,N_167,N_171);
and U879 (N_879,N_162,N_575);
nand U880 (N_880,N_180,N_470);
or U881 (N_881,N_557,N_491);
nand U882 (N_882,N_553,N_121);
or U883 (N_883,N_362,N_586);
xnor U884 (N_884,N_583,N_542);
nand U885 (N_885,N_269,N_109);
nand U886 (N_886,N_33,N_276);
xor U887 (N_887,N_20,N_438);
nand U888 (N_888,N_231,N_310);
and U889 (N_889,N_108,N_392);
nand U890 (N_890,N_411,N_498);
and U891 (N_891,N_497,N_366);
and U892 (N_892,N_488,N_255);
nand U893 (N_893,N_213,N_462);
nor U894 (N_894,N_29,N_565);
nor U895 (N_895,N_399,N_455);
and U896 (N_896,N_223,N_6);
and U897 (N_897,N_342,N_126);
and U898 (N_898,N_580,N_289);
nor U899 (N_899,N_199,N_208);
nand U900 (N_900,N_89,N_144);
or U901 (N_901,N_320,N_169);
and U902 (N_902,N_438,N_229);
nand U903 (N_903,N_268,N_9);
and U904 (N_904,N_332,N_171);
and U905 (N_905,N_334,N_576);
xnor U906 (N_906,N_169,N_77);
or U907 (N_907,N_256,N_258);
xnor U908 (N_908,N_24,N_577);
and U909 (N_909,N_110,N_238);
and U910 (N_910,N_4,N_464);
or U911 (N_911,N_479,N_201);
nand U912 (N_912,N_499,N_206);
xor U913 (N_913,N_527,N_312);
or U914 (N_914,N_44,N_580);
or U915 (N_915,N_337,N_427);
xor U916 (N_916,N_312,N_59);
nand U917 (N_917,N_16,N_81);
or U918 (N_918,N_68,N_353);
nand U919 (N_919,N_522,N_73);
and U920 (N_920,N_445,N_202);
xnor U921 (N_921,N_46,N_264);
or U922 (N_922,N_3,N_146);
nor U923 (N_923,N_462,N_495);
nor U924 (N_924,N_440,N_450);
nor U925 (N_925,N_290,N_338);
xor U926 (N_926,N_283,N_246);
and U927 (N_927,N_222,N_401);
nor U928 (N_928,N_221,N_121);
and U929 (N_929,N_196,N_205);
and U930 (N_930,N_161,N_49);
nand U931 (N_931,N_223,N_140);
or U932 (N_932,N_555,N_354);
and U933 (N_933,N_504,N_224);
xor U934 (N_934,N_45,N_315);
or U935 (N_935,N_102,N_417);
nand U936 (N_936,N_94,N_595);
nor U937 (N_937,N_498,N_406);
nand U938 (N_938,N_262,N_353);
nor U939 (N_939,N_389,N_235);
nand U940 (N_940,N_350,N_520);
xnor U941 (N_941,N_472,N_522);
and U942 (N_942,N_500,N_181);
nor U943 (N_943,N_268,N_308);
and U944 (N_944,N_378,N_66);
nand U945 (N_945,N_478,N_439);
or U946 (N_946,N_412,N_346);
and U947 (N_947,N_144,N_343);
and U948 (N_948,N_483,N_441);
nand U949 (N_949,N_517,N_386);
or U950 (N_950,N_35,N_289);
nand U951 (N_951,N_427,N_282);
or U952 (N_952,N_12,N_79);
or U953 (N_953,N_57,N_10);
or U954 (N_954,N_567,N_560);
nand U955 (N_955,N_459,N_227);
or U956 (N_956,N_569,N_253);
nand U957 (N_957,N_353,N_157);
nor U958 (N_958,N_32,N_430);
or U959 (N_959,N_251,N_486);
and U960 (N_960,N_575,N_476);
nand U961 (N_961,N_395,N_29);
and U962 (N_962,N_478,N_107);
nor U963 (N_963,N_155,N_576);
and U964 (N_964,N_35,N_498);
nor U965 (N_965,N_95,N_110);
xnor U966 (N_966,N_20,N_449);
and U967 (N_967,N_435,N_85);
nand U968 (N_968,N_112,N_480);
nor U969 (N_969,N_191,N_174);
nand U970 (N_970,N_581,N_199);
and U971 (N_971,N_174,N_38);
or U972 (N_972,N_48,N_568);
xor U973 (N_973,N_25,N_165);
nor U974 (N_974,N_299,N_1);
or U975 (N_975,N_431,N_194);
or U976 (N_976,N_227,N_498);
nand U977 (N_977,N_202,N_208);
or U978 (N_978,N_257,N_436);
xor U979 (N_979,N_419,N_223);
xor U980 (N_980,N_178,N_257);
or U981 (N_981,N_585,N_498);
nor U982 (N_982,N_50,N_306);
nand U983 (N_983,N_583,N_439);
and U984 (N_984,N_394,N_599);
and U985 (N_985,N_436,N_458);
nor U986 (N_986,N_155,N_319);
nor U987 (N_987,N_184,N_227);
xor U988 (N_988,N_521,N_503);
xor U989 (N_989,N_510,N_122);
or U990 (N_990,N_442,N_251);
and U991 (N_991,N_74,N_55);
and U992 (N_992,N_28,N_488);
or U993 (N_993,N_210,N_187);
and U994 (N_994,N_50,N_356);
nor U995 (N_995,N_467,N_356);
or U996 (N_996,N_289,N_87);
and U997 (N_997,N_478,N_554);
or U998 (N_998,N_394,N_376);
and U999 (N_999,N_312,N_40);
xor U1000 (N_1000,N_269,N_422);
or U1001 (N_1001,N_582,N_251);
and U1002 (N_1002,N_159,N_278);
and U1003 (N_1003,N_543,N_222);
nand U1004 (N_1004,N_503,N_526);
xor U1005 (N_1005,N_588,N_4);
nand U1006 (N_1006,N_360,N_429);
and U1007 (N_1007,N_44,N_256);
xor U1008 (N_1008,N_420,N_419);
xor U1009 (N_1009,N_338,N_367);
nand U1010 (N_1010,N_422,N_74);
xnor U1011 (N_1011,N_317,N_291);
xnor U1012 (N_1012,N_534,N_344);
nor U1013 (N_1013,N_564,N_11);
nand U1014 (N_1014,N_213,N_477);
nor U1015 (N_1015,N_216,N_455);
and U1016 (N_1016,N_429,N_29);
nand U1017 (N_1017,N_97,N_318);
nor U1018 (N_1018,N_71,N_572);
or U1019 (N_1019,N_54,N_502);
nor U1020 (N_1020,N_333,N_419);
or U1021 (N_1021,N_57,N_9);
and U1022 (N_1022,N_432,N_277);
xor U1023 (N_1023,N_532,N_466);
nand U1024 (N_1024,N_472,N_369);
nor U1025 (N_1025,N_496,N_488);
nor U1026 (N_1026,N_109,N_408);
or U1027 (N_1027,N_307,N_160);
nand U1028 (N_1028,N_430,N_407);
xnor U1029 (N_1029,N_353,N_576);
and U1030 (N_1030,N_404,N_183);
xnor U1031 (N_1031,N_146,N_206);
nor U1032 (N_1032,N_352,N_177);
and U1033 (N_1033,N_519,N_99);
xnor U1034 (N_1034,N_435,N_547);
or U1035 (N_1035,N_31,N_512);
xor U1036 (N_1036,N_503,N_580);
nand U1037 (N_1037,N_420,N_291);
and U1038 (N_1038,N_128,N_589);
nor U1039 (N_1039,N_493,N_332);
xnor U1040 (N_1040,N_221,N_54);
xnor U1041 (N_1041,N_240,N_304);
xnor U1042 (N_1042,N_566,N_570);
nor U1043 (N_1043,N_105,N_514);
nor U1044 (N_1044,N_156,N_261);
nand U1045 (N_1045,N_195,N_87);
or U1046 (N_1046,N_278,N_26);
and U1047 (N_1047,N_117,N_445);
and U1048 (N_1048,N_42,N_256);
or U1049 (N_1049,N_319,N_571);
nor U1050 (N_1050,N_64,N_12);
nor U1051 (N_1051,N_544,N_452);
nand U1052 (N_1052,N_132,N_349);
and U1053 (N_1053,N_63,N_186);
nand U1054 (N_1054,N_33,N_224);
nor U1055 (N_1055,N_535,N_458);
nor U1056 (N_1056,N_394,N_496);
xnor U1057 (N_1057,N_359,N_194);
and U1058 (N_1058,N_145,N_556);
nand U1059 (N_1059,N_471,N_253);
nor U1060 (N_1060,N_48,N_16);
xnor U1061 (N_1061,N_468,N_3);
xor U1062 (N_1062,N_113,N_278);
xnor U1063 (N_1063,N_74,N_204);
or U1064 (N_1064,N_536,N_194);
xor U1065 (N_1065,N_217,N_59);
or U1066 (N_1066,N_253,N_375);
and U1067 (N_1067,N_543,N_29);
nor U1068 (N_1068,N_174,N_459);
nor U1069 (N_1069,N_233,N_397);
xnor U1070 (N_1070,N_337,N_446);
nand U1071 (N_1071,N_578,N_270);
nand U1072 (N_1072,N_552,N_546);
nand U1073 (N_1073,N_418,N_12);
or U1074 (N_1074,N_99,N_79);
nor U1075 (N_1075,N_204,N_270);
nor U1076 (N_1076,N_582,N_415);
and U1077 (N_1077,N_384,N_237);
and U1078 (N_1078,N_465,N_491);
or U1079 (N_1079,N_261,N_441);
and U1080 (N_1080,N_393,N_9);
nand U1081 (N_1081,N_289,N_384);
nand U1082 (N_1082,N_276,N_406);
and U1083 (N_1083,N_335,N_184);
nor U1084 (N_1084,N_586,N_437);
or U1085 (N_1085,N_288,N_95);
or U1086 (N_1086,N_541,N_473);
or U1087 (N_1087,N_65,N_101);
nor U1088 (N_1088,N_446,N_336);
or U1089 (N_1089,N_13,N_460);
and U1090 (N_1090,N_411,N_406);
nor U1091 (N_1091,N_475,N_314);
nor U1092 (N_1092,N_193,N_399);
or U1093 (N_1093,N_315,N_494);
or U1094 (N_1094,N_354,N_108);
or U1095 (N_1095,N_509,N_315);
or U1096 (N_1096,N_343,N_376);
nand U1097 (N_1097,N_17,N_429);
nor U1098 (N_1098,N_269,N_325);
nor U1099 (N_1099,N_308,N_427);
or U1100 (N_1100,N_225,N_315);
or U1101 (N_1101,N_14,N_394);
nand U1102 (N_1102,N_187,N_77);
nand U1103 (N_1103,N_265,N_217);
xnor U1104 (N_1104,N_235,N_33);
nand U1105 (N_1105,N_176,N_153);
nor U1106 (N_1106,N_451,N_306);
nand U1107 (N_1107,N_593,N_424);
nor U1108 (N_1108,N_567,N_400);
and U1109 (N_1109,N_476,N_108);
and U1110 (N_1110,N_289,N_151);
nand U1111 (N_1111,N_96,N_80);
xnor U1112 (N_1112,N_268,N_507);
nor U1113 (N_1113,N_327,N_455);
xor U1114 (N_1114,N_398,N_292);
nand U1115 (N_1115,N_121,N_86);
xor U1116 (N_1116,N_463,N_525);
nand U1117 (N_1117,N_480,N_481);
nand U1118 (N_1118,N_244,N_3);
and U1119 (N_1119,N_154,N_35);
nor U1120 (N_1120,N_454,N_209);
xnor U1121 (N_1121,N_425,N_27);
and U1122 (N_1122,N_476,N_124);
nand U1123 (N_1123,N_316,N_379);
nor U1124 (N_1124,N_562,N_375);
xor U1125 (N_1125,N_408,N_241);
xor U1126 (N_1126,N_10,N_586);
nor U1127 (N_1127,N_486,N_557);
nor U1128 (N_1128,N_401,N_415);
xnor U1129 (N_1129,N_518,N_135);
and U1130 (N_1130,N_119,N_197);
nor U1131 (N_1131,N_551,N_376);
xor U1132 (N_1132,N_429,N_489);
or U1133 (N_1133,N_206,N_2);
or U1134 (N_1134,N_475,N_347);
nand U1135 (N_1135,N_97,N_478);
nor U1136 (N_1136,N_161,N_520);
or U1137 (N_1137,N_354,N_38);
xnor U1138 (N_1138,N_220,N_498);
or U1139 (N_1139,N_482,N_301);
or U1140 (N_1140,N_332,N_570);
nor U1141 (N_1141,N_264,N_357);
or U1142 (N_1142,N_358,N_242);
and U1143 (N_1143,N_547,N_327);
or U1144 (N_1144,N_72,N_442);
nand U1145 (N_1145,N_556,N_421);
and U1146 (N_1146,N_161,N_322);
nor U1147 (N_1147,N_71,N_126);
xnor U1148 (N_1148,N_511,N_59);
nor U1149 (N_1149,N_370,N_453);
xor U1150 (N_1150,N_313,N_383);
nor U1151 (N_1151,N_407,N_562);
or U1152 (N_1152,N_538,N_542);
nor U1153 (N_1153,N_544,N_528);
nor U1154 (N_1154,N_106,N_359);
nor U1155 (N_1155,N_99,N_249);
nor U1156 (N_1156,N_565,N_302);
xnor U1157 (N_1157,N_551,N_154);
and U1158 (N_1158,N_182,N_580);
and U1159 (N_1159,N_10,N_476);
or U1160 (N_1160,N_236,N_295);
xor U1161 (N_1161,N_338,N_311);
and U1162 (N_1162,N_312,N_458);
or U1163 (N_1163,N_387,N_386);
nand U1164 (N_1164,N_26,N_120);
xor U1165 (N_1165,N_570,N_497);
xnor U1166 (N_1166,N_223,N_17);
nand U1167 (N_1167,N_11,N_586);
nand U1168 (N_1168,N_551,N_225);
and U1169 (N_1169,N_129,N_518);
xor U1170 (N_1170,N_34,N_84);
xnor U1171 (N_1171,N_280,N_498);
xnor U1172 (N_1172,N_36,N_561);
nand U1173 (N_1173,N_88,N_0);
or U1174 (N_1174,N_514,N_180);
xor U1175 (N_1175,N_585,N_475);
and U1176 (N_1176,N_220,N_211);
xor U1177 (N_1177,N_427,N_529);
nand U1178 (N_1178,N_349,N_495);
nor U1179 (N_1179,N_209,N_346);
xnor U1180 (N_1180,N_279,N_438);
or U1181 (N_1181,N_184,N_449);
or U1182 (N_1182,N_245,N_337);
and U1183 (N_1183,N_362,N_363);
nand U1184 (N_1184,N_594,N_347);
nand U1185 (N_1185,N_560,N_68);
or U1186 (N_1186,N_46,N_373);
xor U1187 (N_1187,N_564,N_343);
xnor U1188 (N_1188,N_499,N_84);
xnor U1189 (N_1189,N_208,N_263);
or U1190 (N_1190,N_365,N_302);
or U1191 (N_1191,N_403,N_119);
and U1192 (N_1192,N_150,N_363);
or U1193 (N_1193,N_508,N_243);
nand U1194 (N_1194,N_288,N_158);
xnor U1195 (N_1195,N_450,N_184);
and U1196 (N_1196,N_100,N_179);
xnor U1197 (N_1197,N_394,N_193);
and U1198 (N_1198,N_305,N_448);
nor U1199 (N_1199,N_572,N_164);
nand U1200 (N_1200,N_819,N_1044);
nand U1201 (N_1201,N_953,N_1006);
or U1202 (N_1202,N_888,N_1188);
nor U1203 (N_1203,N_663,N_868);
and U1204 (N_1204,N_951,N_1049);
and U1205 (N_1205,N_812,N_661);
or U1206 (N_1206,N_1136,N_689);
nand U1207 (N_1207,N_835,N_1091);
xor U1208 (N_1208,N_647,N_802);
nand U1209 (N_1209,N_1171,N_1076);
or U1210 (N_1210,N_1056,N_952);
or U1211 (N_1211,N_783,N_1126);
xnor U1212 (N_1212,N_902,N_1169);
nand U1213 (N_1213,N_822,N_636);
or U1214 (N_1214,N_635,N_771);
nor U1215 (N_1215,N_977,N_1102);
nor U1216 (N_1216,N_1035,N_796);
or U1217 (N_1217,N_1081,N_624);
xor U1218 (N_1218,N_1124,N_801);
or U1219 (N_1219,N_1163,N_1167);
and U1220 (N_1220,N_821,N_1038);
and U1221 (N_1221,N_757,N_954);
or U1222 (N_1222,N_1096,N_874);
nor U1223 (N_1223,N_1170,N_705);
nor U1224 (N_1224,N_713,N_745);
or U1225 (N_1225,N_621,N_804);
nor U1226 (N_1226,N_1045,N_708);
nor U1227 (N_1227,N_881,N_1024);
nand U1228 (N_1228,N_865,N_973);
nand U1229 (N_1229,N_926,N_1140);
xnor U1230 (N_1230,N_749,N_845);
or U1231 (N_1231,N_1037,N_982);
and U1232 (N_1232,N_1000,N_1069);
xor U1233 (N_1233,N_862,N_1041);
and U1234 (N_1234,N_660,N_808);
or U1235 (N_1235,N_731,N_712);
nand U1236 (N_1236,N_722,N_844);
xnor U1237 (N_1237,N_827,N_652);
xor U1238 (N_1238,N_627,N_1100);
and U1239 (N_1239,N_920,N_693);
or U1240 (N_1240,N_1180,N_943);
or U1241 (N_1241,N_1112,N_940);
or U1242 (N_1242,N_999,N_1178);
and U1243 (N_1243,N_891,N_662);
nand U1244 (N_1244,N_1048,N_645);
and U1245 (N_1245,N_746,N_738);
nand U1246 (N_1246,N_809,N_747);
or U1247 (N_1247,N_915,N_942);
or U1248 (N_1248,N_702,N_1017);
and U1249 (N_1249,N_1158,N_1125);
and U1250 (N_1250,N_728,N_733);
nand U1251 (N_1251,N_1004,N_840);
nand U1252 (N_1252,N_696,N_719);
nand U1253 (N_1253,N_1055,N_1011);
nor U1254 (N_1254,N_743,N_969);
nand U1255 (N_1255,N_721,N_695);
nand U1256 (N_1256,N_1007,N_836);
nand U1257 (N_1257,N_889,N_676);
and U1258 (N_1258,N_994,N_707);
xor U1259 (N_1259,N_741,N_1071);
nor U1260 (N_1260,N_1190,N_601);
nor U1261 (N_1261,N_1014,N_607);
nor U1262 (N_1262,N_1067,N_777);
nand U1263 (N_1263,N_1159,N_1144);
nor U1264 (N_1264,N_1064,N_780);
nor U1265 (N_1265,N_772,N_1122);
nor U1266 (N_1266,N_1111,N_671);
xor U1267 (N_1267,N_1120,N_970);
nor U1268 (N_1268,N_978,N_755);
or U1269 (N_1269,N_814,N_1090);
xnor U1270 (N_1270,N_632,N_622);
or U1271 (N_1271,N_798,N_1198);
and U1272 (N_1272,N_892,N_643);
nand U1273 (N_1273,N_818,N_870);
or U1274 (N_1274,N_1103,N_717);
nand U1275 (N_1275,N_1181,N_824);
nor U1276 (N_1276,N_1052,N_976);
xnor U1277 (N_1277,N_933,N_995);
and U1278 (N_1278,N_911,N_838);
or U1279 (N_1279,N_1105,N_826);
nand U1280 (N_1280,N_1191,N_616);
xnor U1281 (N_1281,N_816,N_828);
or U1282 (N_1282,N_1080,N_887);
nor U1283 (N_1283,N_972,N_1086);
nand U1284 (N_1284,N_834,N_1187);
and U1285 (N_1285,N_955,N_1147);
xnor U1286 (N_1286,N_817,N_986);
nor U1287 (N_1287,N_753,N_803);
xnor U1288 (N_1288,N_609,N_1095);
xnor U1289 (N_1289,N_856,N_992);
nor U1290 (N_1290,N_684,N_852);
nand U1291 (N_1291,N_1013,N_1097);
nor U1292 (N_1292,N_1012,N_1094);
nand U1293 (N_1293,N_989,N_767);
nor U1294 (N_1294,N_1059,N_993);
xor U1295 (N_1295,N_752,N_1110);
or U1296 (N_1296,N_651,N_1028);
nor U1297 (N_1297,N_1009,N_1173);
and U1298 (N_1298,N_659,N_1057);
nor U1299 (N_1299,N_829,N_691);
or U1300 (N_1300,N_965,N_1070);
nor U1301 (N_1301,N_629,N_681);
or U1302 (N_1302,N_1177,N_967);
or U1303 (N_1303,N_930,N_700);
or U1304 (N_1304,N_1050,N_1075);
and U1305 (N_1305,N_1164,N_825);
xor U1306 (N_1306,N_857,N_739);
nand U1307 (N_1307,N_639,N_1082);
or U1308 (N_1308,N_793,N_778);
nand U1309 (N_1309,N_883,N_984);
xnor U1310 (N_1310,N_1139,N_987);
and U1311 (N_1311,N_974,N_669);
nand U1312 (N_1312,N_1117,N_1099);
xnor U1313 (N_1313,N_1036,N_961);
or U1314 (N_1314,N_690,N_1032);
nor U1315 (N_1315,N_718,N_960);
and U1316 (N_1316,N_633,N_879);
nand U1317 (N_1317,N_805,N_1145);
nor U1318 (N_1318,N_626,N_935);
nor U1319 (N_1319,N_1039,N_895);
or U1320 (N_1320,N_763,N_667);
xor U1321 (N_1321,N_1186,N_664);
or U1322 (N_1322,N_637,N_958);
or U1323 (N_1323,N_1020,N_619);
and U1324 (N_1324,N_1153,N_656);
nand U1325 (N_1325,N_1029,N_921);
nand U1326 (N_1326,N_1134,N_864);
nor U1327 (N_1327,N_1098,N_668);
and U1328 (N_1328,N_1152,N_615);
xnor U1329 (N_1329,N_797,N_727);
and U1330 (N_1330,N_848,N_1054);
and U1331 (N_1331,N_1043,N_991);
or U1332 (N_1332,N_1137,N_628);
nor U1333 (N_1333,N_1130,N_1051);
or U1334 (N_1334,N_714,N_985);
nor U1335 (N_1335,N_674,N_610);
nand U1336 (N_1336,N_710,N_1109);
nand U1337 (N_1337,N_799,N_1063);
nand U1338 (N_1338,N_766,N_792);
nor U1339 (N_1339,N_1066,N_754);
xor U1340 (N_1340,N_631,N_841);
xnor U1341 (N_1341,N_878,N_861);
or U1342 (N_1342,N_704,N_751);
nand U1343 (N_1343,N_1128,N_945);
and U1344 (N_1344,N_996,N_882);
nand U1345 (N_1345,N_1085,N_897);
nand U1346 (N_1346,N_709,N_867);
and U1347 (N_1347,N_981,N_744);
nor U1348 (N_1348,N_927,N_903);
xnor U1349 (N_1349,N_800,N_618);
or U1350 (N_1350,N_877,N_658);
and U1351 (N_1351,N_711,N_697);
nor U1352 (N_1352,N_941,N_916);
nor U1353 (N_1353,N_1079,N_815);
or U1354 (N_1354,N_929,N_790);
xor U1355 (N_1355,N_1087,N_602);
xnor U1356 (N_1356,N_1197,N_1005);
and U1357 (N_1357,N_1101,N_979);
xor U1358 (N_1358,N_625,N_657);
nand U1359 (N_1359,N_1168,N_1175);
nor U1360 (N_1360,N_1018,N_880);
or U1361 (N_1361,N_795,N_923);
and U1362 (N_1362,N_1061,N_666);
or U1363 (N_1363,N_860,N_1001);
nor U1364 (N_1364,N_905,N_904);
or U1365 (N_1365,N_644,N_604);
and U1366 (N_1366,N_1053,N_837);
nor U1367 (N_1367,N_910,N_928);
nor U1368 (N_1368,N_638,N_931);
xor U1369 (N_1369,N_1021,N_724);
or U1370 (N_1370,N_1143,N_830);
nor U1371 (N_1371,N_1060,N_1192);
and U1372 (N_1372,N_641,N_894);
and U1373 (N_1373,N_823,N_1189);
nand U1374 (N_1374,N_855,N_850);
and U1375 (N_1375,N_1183,N_1078);
and U1376 (N_1376,N_901,N_1156);
xor U1377 (N_1377,N_925,N_898);
nor U1378 (N_1378,N_1114,N_1157);
nand U1379 (N_1379,N_703,N_1031);
nor U1380 (N_1380,N_948,N_715);
or U1381 (N_1381,N_936,N_938);
and U1382 (N_1382,N_1142,N_776);
and U1383 (N_1383,N_726,N_983);
or U1384 (N_1384,N_839,N_701);
xnor U1385 (N_1385,N_1148,N_842);
nand U1386 (N_1386,N_886,N_832);
nor U1387 (N_1387,N_1106,N_1022);
nor U1388 (N_1388,N_642,N_851);
or U1389 (N_1389,N_646,N_813);
xnor U1390 (N_1390,N_617,N_909);
nor U1391 (N_1391,N_1062,N_1104);
nand U1392 (N_1392,N_680,N_1123);
xor U1393 (N_1393,N_1182,N_1116);
nor U1394 (N_1394,N_863,N_846);
xor U1395 (N_1395,N_1166,N_1027);
and U1396 (N_1396,N_1184,N_975);
nand U1397 (N_1397,N_1015,N_1113);
or U1398 (N_1398,N_773,N_786);
nand U1399 (N_1399,N_620,N_914);
and U1400 (N_1400,N_736,N_1141);
xor U1401 (N_1401,N_1072,N_650);
xor U1402 (N_1402,N_768,N_716);
xnor U1403 (N_1403,N_988,N_956);
xnor U1404 (N_1404,N_765,N_922);
nor U1405 (N_1405,N_779,N_1160);
and U1406 (N_1406,N_730,N_1115);
nor U1407 (N_1407,N_678,N_756);
xnor U1408 (N_1408,N_694,N_748);
and U1409 (N_1409,N_1065,N_630);
and U1410 (N_1410,N_605,N_924);
or U1411 (N_1411,N_939,N_764);
nand U1412 (N_1412,N_675,N_912);
nor U1413 (N_1413,N_859,N_687);
xnor U1414 (N_1414,N_688,N_1146);
nand U1415 (N_1415,N_723,N_740);
or U1416 (N_1416,N_872,N_854);
or U1417 (N_1417,N_820,N_734);
nand U1418 (N_1418,N_1088,N_1058);
and U1419 (N_1419,N_1121,N_1155);
and U1420 (N_1420,N_1034,N_774);
nand U1421 (N_1421,N_1074,N_654);
and U1422 (N_1422,N_1084,N_634);
and U1423 (N_1423,N_699,N_866);
or U1424 (N_1424,N_770,N_1161);
xor U1425 (N_1425,N_1131,N_1119);
nand U1426 (N_1426,N_1127,N_937);
or U1427 (N_1427,N_1129,N_1083);
nand U1428 (N_1428,N_1151,N_735);
and U1429 (N_1429,N_871,N_869);
or U1430 (N_1430,N_784,N_962);
nand U1431 (N_1431,N_653,N_1077);
and U1432 (N_1432,N_677,N_1008);
nor U1433 (N_1433,N_1108,N_858);
xor U1434 (N_1434,N_758,N_1199);
nand U1435 (N_1435,N_762,N_1193);
or U1436 (N_1436,N_614,N_1165);
or U1437 (N_1437,N_785,N_1089);
nor U1438 (N_1438,N_890,N_1195);
nand U1439 (N_1439,N_665,N_1073);
nand U1440 (N_1440,N_876,N_794);
and U1441 (N_1441,N_791,N_811);
or U1442 (N_1442,N_698,N_692);
nand U1443 (N_1443,N_649,N_682);
or U1444 (N_1444,N_725,N_600);
xnor U1445 (N_1445,N_908,N_672);
nand U1446 (N_1446,N_1194,N_1042);
nand U1447 (N_1447,N_1016,N_750);
or U1448 (N_1448,N_963,N_1154);
nand U1449 (N_1449,N_907,N_980);
xnor U1450 (N_1450,N_685,N_623);
xnor U1451 (N_1451,N_1196,N_742);
xor U1452 (N_1452,N_906,N_1176);
nand U1453 (N_1453,N_606,N_1026);
xnor U1454 (N_1454,N_833,N_612);
xor U1455 (N_1455,N_608,N_946);
and U1456 (N_1456,N_673,N_949);
nor U1457 (N_1457,N_1133,N_831);
xnor U1458 (N_1458,N_843,N_1093);
xnor U1459 (N_1459,N_807,N_959);
nor U1460 (N_1460,N_810,N_613);
xnor U1461 (N_1461,N_679,N_875);
or U1462 (N_1462,N_1162,N_670);
nand U1463 (N_1463,N_950,N_968);
or U1464 (N_1464,N_917,N_782);
nor U1465 (N_1465,N_900,N_706);
nor U1466 (N_1466,N_1138,N_1172);
nand U1467 (N_1467,N_849,N_640);
nor U1468 (N_1468,N_932,N_759);
nand U1469 (N_1469,N_603,N_1046);
or U1470 (N_1470,N_997,N_1003);
or U1471 (N_1471,N_1132,N_1033);
nor U1472 (N_1472,N_885,N_847);
nand U1473 (N_1473,N_1047,N_913);
and U1474 (N_1474,N_611,N_760);
nand U1475 (N_1475,N_893,N_853);
nor U1476 (N_1476,N_769,N_1023);
nand U1477 (N_1477,N_884,N_964);
nand U1478 (N_1478,N_737,N_990);
or U1479 (N_1479,N_873,N_787);
and U1480 (N_1480,N_966,N_1010);
or U1481 (N_1481,N_1174,N_1030);
nand U1482 (N_1482,N_655,N_944);
xnor U1483 (N_1483,N_788,N_781);
xnor U1484 (N_1484,N_683,N_1107);
and U1485 (N_1485,N_1019,N_775);
and U1486 (N_1486,N_686,N_789);
nand U1487 (N_1487,N_919,N_1068);
and U1488 (N_1488,N_971,N_1185);
nor U1489 (N_1489,N_896,N_998);
nor U1490 (N_1490,N_806,N_934);
or U1491 (N_1491,N_732,N_957);
or U1492 (N_1492,N_720,N_1092);
nand U1493 (N_1493,N_1150,N_1135);
nor U1494 (N_1494,N_947,N_1025);
nand U1495 (N_1495,N_918,N_1002);
xor U1496 (N_1496,N_648,N_729);
nand U1497 (N_1497,N_1149,N_899);
nor U1498 (N_1498,N_1118,N_1040);
or U1499 (N_1499,N_761,N_1179);
nand U1500 (N_1500,N_872,N_669);
nand U1501 (N_1501,N_1071,N_732);
or U1502 (N_1502,N_1018,N_795);
or U1503 (N_1503,N_680,N_876);
or U1504 (N_1504,N_1151,N_1117);
nor U1505 (N_1505,N_1144,N_1098);
or U1506 (N_1506,N_1126,N_1081);
or U1507 (N_1507,N_1035,N_699);
xnor U1508 (N_1508,N_884,N_692);
nand U1509 (N_1509,N_747,N_734);
nor U1510 (N_1510,N_1050,N_652);
xnor U1511 (N_1511,N_625,N_656);
xor U1512 (N_1512,N_734,N_761);
or U1513 (N_1513,N_874,N_965);
and U1514 (N_1514,N_1129,N_903);
nand U1515 (N_1515,N_875,N_1038);
xnor U1516 (N_1516,N_1005,N_856);
nor U1517 (N_1517,N_1061,N_751);
xor U1518 (N_1518,N_986,N_1154);
and U1519 (N_1519,N_1065,N_1019);
xor U1520 (N_1520,N_1055,N_869);
nor U1521 (N_1521,N_1119,N_767);
or U1522 (N_1522,N_1064,N_783);
and U1523 (N_1523,N_905,N_1117);
nor U1524 (N_1524,N_796,N_625);
or U1525 (N_1525,N_1050,N_855);
nand U1526 (N_1526,N_650,N_931);
or U1527 (N_1527,N_605,N_831);
nor U1528 (N_1528,N_695,N_774);
nand U1529 (N_1529,N_696,N_605);
or U1530 (N_1530,N_676,N_933);
and U1531 (N_1531,N_1053,N_1147);
nand U1532 (N_1532,N_989,N_679);
nor U1533 (N_1533,N_1107,N_1153);
and U1534 (N_1534,N_711,N_1015);
nand U1535 (N_1535,N_1089,N_670);
or U1536 (N_1536,N_1096,N_707);
nand U1537 (N_1537,N_856,N_739);
xor U1538 (N_1538,N_759,N_1150);
nand U1539 (N_1539,N_1188,N_1171);
or U1540 (N_1540,N_848,N_729);
or U1541 (N_1541,N_1168,N_777);
or U1542 (N_1542,N_758,N_787);
nand U1543 (N_1543,N_1109,N_751);
or U1544 (N_1544,N_625,N_703);
and U1545 (N_1545,N_807,N_786);
and U1546 (N_1546,N_765,N_955);
or U1547 (N_1547,N_936,N_965);
and U1548 (N_1548,N_799,N_1085);
nor U1549 (N_1549,N_1152,N_785);
nand U1550 (N_1550,N_886,N_782);
nand U1551 (N_1551,N_1025,N_903);
nand U1552 (N_1552,N_980,N_1125);
and U1553 (N_1553,N_808,N_667);
xor U1554 (N_1554,N_621,N_849);
nand U1555 (N_1555,N_882,N_1075);
xor U1556 (N_1556,N_659,N_631);
or U1557 (N_1557,N_608,N_1187);
or U1558 (N_1558,N_765,N_759);
nand U1559 (N_1559,N_646,N_1032);
nand U1560 (N_1560,N_781,N_706);
nand U1561 (N_1561,N_810,N_1000);
or U1562 (N_1562,N_838,N_1102);
and U1563 (N_1563,N_937,N_649);
or U1564 (N_1564,N_884,N_1039);
xor U1565 (N_1565,N_730,N_759);
nor U1566 (N_1566,N_760,N_1051);
or U1567 (N_1567,N_610,N_613);
nor U1568 (N_1568,N_1077,N_917);
xor U1569 (N_1569,N_734,N_909);
and U1570 (N_1570,N_1058,N_867);
or U1571 (N_1571,N_883,N_720);
or U1572 (N_1572,N_717,N_898);
nor U1573 (N_1573,N_1115,N_725);
or U1574 (N_1574,N_655,N_984);
xor U1575 (N_1575,N_732,N_1083);
xor U1576 (N_1576,N_970,N_1140);
nor U1577 (N_1577,N_619,N_769);
and U1578 (N_1578,N_814,N_1075);
xnor U1579 (N_1579,N_943,N_671);
and U1580 (N_1580,N_1063,N_1034);
or U1581 (N_1581,N_1176,N_627);
xnor U1582 (N_1582,N_935,N_685);
nor U1583 (N_1583,N_638,N_649);
nor U1584 (N_1584,N_1026,N_625);
nor U1585 (N_1585,N_1045,N_647);
and U1586 (N_1586,N_755,N_1059);
xnor U1587 (N_1587,N_829,N_972);
nor U1588 (N_1588,N_1040,N_937);
xnor U1589 (N_1589,N_982,N_1156);
nor U1590 (N_1590,N_1163,N_973);
or U1591 (N_1591,N_946,N_1144);
nor U1592 (N_1592,N_988,N_897);
nor U1593 (N_1593,N_991,N_895);
and U1594 (N_1594,N_1003,N_827);
nand U1595 (N_1595,N_917,N_612);
nand U1596 (N_1596,N_745,N_1109);
xor U1597 (N_1597,N_1139,N_636);
and U1598 (N_1598,N_1065,N_640);
or U1599 (N_1599,N_657,N_999);
nor U1600 (N_1600,N_823,N_840);
xor U1601 (N_1601,N_737,N_750);
nor U1602 (N_1602,N_892,N_688);
nand U1603 (N_1603,N_761,N_1164);
or U1604 (N_1604,N_737,N_1049);
nor U1605 (N_1605,N_1069,N_1171);
nor U1606 (N_1606,N_730,N_896);
and U1607 (N_1607,N_739,N_765);
xor U1608 (N_1608,N_1121,N_1020);
nor U1609 (N_1609,N_863,N_815);
xnor U1610 (N_1610,N_1182,N_1055);
and U1611 (N_1611,N_751,N_927);
nor U1612 (N_1612,N_711,N_880);
xnor U1613 (N_1613,N_1096,N_875);
nand U1614 (N_1614,N_1112,N_872);
nor U1615 (N_1615,N_643,N_869);
xor U1616 (N_1616,N_817,N_660);
xnor U1617 (N_1617,N_1019,N_1191);
or U1618 (N_1618,N_1190,N_675);
or U1619 (N_1619,N_887,N_697);
and U1620 (N_1620,N_955,N_1190);
nand U1621 (N_1621,N_604,N_725);
or U1622 (N_1622,N_790,N_906);
or U1623 (N_1623,N_1024,N_1196);
xnor U1624 (N_1624,N_900,N_916);
nor U1625 (N_1625,N_1185,N_945);
nand U1626 (N_1626,N_1068,N_1073);
nor U1627 (N_1627,N_788,N_1121);
xor U1628 (N_1628,N_1112,N_783);
or U1629 (N_1629,N_778,N_1168);
xor U1630 (N_1630,N_617,N_1072);
and U1631 (N_1631,N_1157,N_1051);
xor U1632 (N_1632,N_790,N_1081);
nor U1633 (N_1633,N_975,N_1060);
nand U1634 (N_1634,N_1110,N_902);
or U1635 (N_1635,N_787,N_1154);
nor U1636 (N_1636,N_639,N_638);
and U1637 (N_1637,N_709,N_1151);
nor U1638 (N_1638,N_965,N_961);
nand U1639 (N_1639,N_1060,N_716);
xor U1640 (N_1640,N_696,N_694);
or U1641 (N_1641,N_655,N_868);
and U1642 (N_1642,N_774,N_603);
xor U1643 (N_1643,N_1077,N_873);
and U1644 (N_1644,N_957,N_1064);
xor U1645 (N_1645,N_1176,N_900);
xnor U1646 (N_1646,N_616,N_751);
nor U1647 (N_1647,N_690,N_661);
or U1648 (N_1648,N_781,N_839);
nor U1649 (N_1649,N_1114,N_857);
or U1650 (N_1650,N_1037,N_612);
or U1651 (N_1651,N_1104,N_1074);
and U1652 (N_1652,N_830,N_942);
xnor U1653 (N_1653,N_996,N_1022);
and U1654 (N_1654,N_1183,N_1049);
xnor U1655 (N_1655,N_1033,N_613);
or U1656 (N_1656,N_660,N_895);
nand U1657 (N_1657,N_862,N_703);
and U1658 (N_1658,N_996,N_994);
nand U1659 (N_1659,N_926,N_845);
nor U1660 (N_1660,N_698,N_702);
xnor U1661 (N_1661,N_1144,N_1077);
or U1662 (N_1662,N_606,N_1159);
nand U1663 (N_1663,N_748,N_813);
xor U1664 (N_1664,N_822,N_804);
xnor U1665 (N_1665,N_751,N_611);
or U1666 (N_1666,N_631,N_1001);
and U1667 (N_1667,N_1115,N_1022);
nor U1668 (N_1668,N_666,N_852);
nor U1669 (N_1669,N_801,N_1141);
xnor U1670 (N_1670,N_864,N_643);
or U1671 (N_1671,N_693,N_1122);
nand U1672 (N_1672,N_1085,N_1121);
nand U1673 (N_1673,N_907,N_744);
xor U1674 (N_1674,N_810,N_1034);
xnor U1675 (N_1675,N_885,N_937);
and U1676 (N_1676,N_741,N_661);
xnor U1677 (N_1677,N_814,N_787);
xnor U1678 (N_1678,N_853,N_850);
and U1679 (N_1679,N_1117,N_1025);
and U1680 (N_1680,N_1168,N_1083);
xnor U1681 (N_1681,N_858,N_869);
nand U1682 (N_1682,N_1129,N_995);
and U1683 (N_1683,N_701,N_739);
and U1684 (N_1684,N_751,N_792);
and U1685 (N_1685,N_1167,N_1196);
nand U1686 (N_1686,N_636,N_743);
nand U1687 (N_1687,N_916,N_616);
nand U1688 (N_1688,N_643,N_680);
and U1689 (N_1689,N_1057,N_865);
nand U1690 (N_1690,N_720,N_1120);
nor U1691 (N_1691,N_949,N_624);
or U1692 (N_1692,N_1152,N_729);
nor U1693 (N_1693,N_601,N_812);
and U1694 (N_1694,N_692,N_783);
nor U1695 (N_1695,N_1102,N_1122);
or U1696 (N_1696,N_689,N_745);
xor U1697 (N_1697,N_1144,N_681);
nor U1698 (N_1698,N_858,N_900);
or U1699 (N_1699,N_1193,N_699);
nor U1700 (N_1700,N_851,N_808);
nand U1701 (N_1701,N_1023,N_1107);
xor U1702 (N_1702,N_895,N_687);
or U1703 (N_1703,N_684,N_812);
or U1704 (N_1704,N_848,N_738);
or U1705 (N_1705,N_1157,N_693);
xnor U1706 (N_1706,N_1151,N_1144);
or U1707 (N_1707,N_1003,N_604);
and U1708 (N_1708,N_907,N_663);
or U1709 (N_1709,N_701,N_742);
and U1710 (N_1710,N_929,N_818);
nand U1711 (N_1711,N_1195,N_671);
or U1712 (N_1712,N_684,N_864);
or U1713 (N_1713,N_1186,N_798);
nor U1714 (N_1714,N_1134,N_1173);
or U1715 (N_1715,N_816,N_867);
and U1716 (N_1716,N_649,N_1087);
nor U1717 (N_1717,N_611,N_918);
and U1718 (N_1718,N_755,N_1071);
nand U1719 (N_1719,N_696,N_829);
nand U1720 (N_1720,N_625,N_802);
nand U1721 (N_1721,N_799,N_910);
nor U1722 (N_1722,N_916,N_841);
and U1723 (N_1723,N_1079,N_819);
nand U1724 (N_1724,N_659,N_638);
or U1725 (N_1725,N_601,N_1015);
and U1726 (N_1726,N_918,N_1069);
xnor U1727 (N_1727,N_796,N_987);
or U1728 (N_1728,N_772,N_765);
or U1729 (N_1729,N_1084,N_727);
nor U1730 (N_1730,N_682,N_737);
and U1731 (N_1731,N_972,N_640);
xor U1732 (N_1732,N_1041,N_709);
nor U1733 (N_1733,N_1197,N_1031);
nor U1734 (N_1734,N_1009,N_904);
xor U1735 (N_1735,N_912,N_690);
nor U1736 (N_1736,N_812,N_676);
nor U1737 (N_1737,N_996,N_767);
nor U1738 (N_1738,N_1157,N_795);
or U1739 (N_1739,N_904,N_640);
or U1740 (N_1740,N_940,N_915);
nand U1741 (N_1741,N_905,N_1023);
nand U1742 (N_1742,N_1183,N_1057);
nor U1743 (N_1743,N_1056,N_805);
and U1744 (N_1744,N_829,N_1093);
xnor U1745 (N_1745,N_871,N_1190);
nor U1746 (N_1746,N_856,N_1053);
or U1747 (N_1747,N_676,N_1040);
nor U1748 (N_1748,N_794,N_676);
and U1749 (N_1749,N_973,N_909);
nand U1750 (N_1750,N_752,N_793);
nand U1751 (N_1751,N_1086,N_806);
nand U1752 (N_1752,N_742,N_859);
nand U1753 (N_1753,N_603,N_1159);
xnor U1754 (N_1754,N_1186,N_942);
and U1755 (N_1755,N_672,N_1080);
and U1756 (N_1756,N_635,N_779);
nor U1757 (N_1757,N_1023,N_706);
xor U1758 (N_1758,N_699,N_897);
nor U1759 (N_1759,N_734,N_783);
nand U1760 (N_1760,N_1165,N_1070);
or U1761 (N_1761,N_775,N_741);
and U1762 (N_1762,N_609,N_885);
and U1763 (N_1763,N_616,N_624);
nand U1764 (N_1764,N_902,N_914);
xnor U1765 (N_1765,N_673,N_1006);
nor U1766 (N_1766,N_989,N_1020);
nor U1767 (N_1767,N_683,N_1031);
nor U1768 (N_1768,N_1137,N_636);
nand U1769 (N_1769,N_753,N_663);
xor U1770 (N_1770,N_957,N_831);
or U1771 (N_1771,N_1123,N_1106);
and U1772 (N_1772,N_778,N_1111);
and U1773 (N_1773,N_1076,N_744);
xor U1774 (N_1774,N_1091,N_1197);
nand U1775 (N_1775,N_889,N_1034);
and U1776 (N_1776,N_623,N_968);
nor U1777 (N_1777,N_782,N_984);
nand U1778 (N_1778,N_696,N_842);
nor U1779 (N_1779,N_1128,N_957);
xnor U1780 (N_1780,N_898,N_1071);
nand U1781 (N_1781,N_1096,N_762);
nor U1782 (N_1782,N_734,N_1183);
xor U1783 (N_1783,N_1021,N_632);
nor U1784 (N_1784,N_621,N_1159);
xnor U1785 (N_1785,N_1103,N_614);
nor U1786 (N_1786,N_1078,N_1137);
nor U1787 (N_1787,N_830,N_850);
xnor U1788 (N_1788,N_685,N_1015);
or U1789 (N_1789,N_866,N_690);
or U1790 (N_1790,N_823,N_982);
nand U1791 (N_1791,N_641,N_650);
xnor U1792 (N_1792,N_1005,N_637);
and U1793 (N_1793,N_1100,N_676);
and U1794 (N_1794,N_950,N_750);
or U1795 (N_1795,N_1079,N_649);
or U1796 (N_1796,N_937,N_713);
and U1797 (N_1797,N_1053,N_1031);
nor U1798 (N_1798,N_1182,N_1127);
and U1799 (N_1799,N_960,N_836);
nand U1800 (N_1800,N_1353,N_1682);
and U1801 (N_1801,N_1606,N_1403);
nor U1802 (N_1802,N_1748,N_1709);
and U1803 (N_1803,N_1303,N_1674);
nor U1804 (N_1804,N_1678,N_1433);
nand U1805 (N_1805,N_1579,N_1321);
nand U1806 (N_1806,N_1635,N_1699);
xnor U1807 (N_1807,N_1411,N_1268);
or U1808 (N_1808,N_1778,N_1218);
nand U1809 (N_1809,N_1581,N_1336);
nand U1810 (N_1810,N_1421,N_1286);
and U1811 (N_1811,N_1607,N_1554);
xnor U1812 (N_1812,N_1762,N_1314);
or U1813 (N_1813,N_1477,N_1618);
nand U1814 (N_1814,N_1670,N_1383);
or U1815 (N_1815,N_1739,N_1728);
xnor U1816 (N_1816,N_1451,N_1436);
xnor U1817 (N_1817,N_1380,N_1253);
nand U1818 (N_1818,N_1462,N_1331);
and U1819 (N_1819,N_1333,N_1575);
nand U1820 (N_1820,N_1794,N_1453);
nor U1821 (N_1821,N_1495,N_1206);
xor U1822 (N_1822,N_1561,N_1463);
nor U1823 (N_1823,N_1422,N_1360);
nor U1824 (N_1824,N_1492,N_1370);
xor U1825 (N_1825,N_1744,N_1538);
and U1826 (N_1826,N_1666,N_1793);
nor U1827 (N_1827,N_1750,N_1279);
xor U1828 (N_1828,N_1284,N_1202);
and U1829 (N_1829,N_1473,N_1511);
nand U1830 (N_1830,N_1297,N_1797);
xor U1831 (N_1831,N_1387,N_1469);
nand U1832 (N_1832,N_1251,N_1273);
nor U1833 (N_1833,N_1700,N_1454);
and U1834 (N_1834,N_1371,N_1540);
and U1835 (N_1835,N_1656,N_1316);
nand U1836 (N_1836,N_1727,N_1757);
xnor U1837 (N_1837,N_1358,N_1576);
nor U1838 (N_1838,N_1388,N_1708);
or U1839 (N_1839,N_1236,N_1614);
xnor U1840 (N_1840,N_1252,N_1330);
nand U1841 (N_1841,N_1207,N_1694);
nor U1842 (N_1842,N_1776,N_1685);
or U1843 (N_1843,N_1315,N_1419);
or U1844 (N_1844,N_1256,N_1265);
or U1845 (N_1845,N_1213,N_1470);
or U1846 (N_1846,N_1342,N_1692);
or U1847 (N_1847,N_1429,N_1501);
xor U1848 (N_1848,N_1633,N_1450);
or U1849 (N_1849,N_1209,N_1483);
and U1850 (N_1850,N_1444,N_1246);
and U1851 (N_1851,N_1766,N_1737);
nor U1852 (N_1852,N_1667,N_1537);
nor U1853 (N_1853,N_1276,N_1407);
nor U1854 (N_1854,N_1617,N_1263);
nor U1855 (N_1855,N_1736,N_1296);
and U1856 (N_1856,N_1564,N_1516);
and U1857 (N_1857,N_1731,N_1711);
nor U1858 (N_1858,N_1362,N_1327);
xor U1859 (N_1859,N_1313,N_1690);
or U1860 (N_1860,N_1285,N_1597);
and U1861 (N_1861,N_1269,N_1572);
xor U1862 (N_1862,N_1544,N_1582);
xnor U1863 (N_1863,N_1496,N_1488);
or U1864 (N_1864,N_1241,N_1220);
nor U1865 (N_1865,N_1248,N_1704);
nand U1866 (N_1866,N_1229,N_1514);
xnor U1867 (N_1867,N_1590,N_1386);
or U1868 (N_1868,N_1465,N_1616);
and U1869 (N_1869,N_1416,N_1442);
xnor U1870 (N_1870,N_1567,N_1243);
nor U1871 (N_1871,N_1369,N_1782);
and U1872 (N_1872,N_1714,N_1536);
or U1873 (N_1873,N_1308,N_1623);
xor U1874 (N_1874,N_1584,N_1780);
or U1875 (N_1875,N_1266,N_1522);
xor U1876 (N_1876,N_1476,N_1726);
or U1877 (N_1877,N_1325,N_1508);
nand U1878 (N_1878,N_1233,N_1751);
nor U1879 (N_1879,N_1557,N_1529);
and U1880 (N_1880,N_1660,N_1424);
nor U1881 (N_1881,N_1441,N_1250);
nand U1882 (N_1882,N_1217,N_1293);
nor U1883 (N_1883,N_1264,N_1348);
nor U1884 (N_1884,N_1790,N_1351);
nor U1885 (N_1885,N_1368,N_1449);
nand U1886 (N_1886,N_1472,N_1578);
and U1887 (N_1887,N_1772,N_1795);
and U1888 (N_1888,N_1211,N_1281);
or U1889 (N_1889,N_1423,N_1773);
nor U1890 (N_1890,N_1254,N_1376);
and U1891 (N_1891,N_1410,N_1418);
xnor U1892 (N_1892,N_1231,N_1585);
and U1893 (N_1893,N_1555,N_1588);
or U1894 (N_1894,N_1735,N_1701);
xor U1895 (N_1895,N_1447,N_1659);
nand U1896 (N_1896,N_1372,N_1577);
nor U1897 (N_1897,N_1689,N_1509);
nand U1898 (N_1898,N_1783,N_1662);
or U1899 (N_1899,N_1551,N_1791);
nor U1900 (N_1900,N_1671,N_1713);
xor U1901 (N_1901,N_1324,N_1752);
xor U1902 (N_1902,N_1535,N_1755);
or U1903 (N_1903,N_1499,N_1389);
nor U1904 (N_1904,N_1352,N_1219);
nor U1905 (N_1905,N_1657,N_1636);
xor U1906 (N_1906,N_1628,N_1366);
and U1907 (N_1907,N_1474,N_1702);
nor U1908 (N_1908,N_1796,N_1640);
and U1909 (N_1909,N_1638,N_1603);
or U1910 (N_1910,N_1365,N_1367);
and U1911 (N_1911,N_1663,N_1210);
xnor U1912 (N_1912,N_1381,N_1393);
and U1913 (N_1913,N_1507,N_1271);
nand U1914 (N_1914,N_1409,N_1771);
nand U1915 (N_1915,N_1503,N_1758);
nand U1916 (N_1916,N_1347,N_1350);
nand U1917 (N_1917,N_1763,N_1767);
nor U1918 (N_1918,N_1677,N_1550);
nand U1919 (N_1919,N_1738,N_1642);
nand U1920 (N_1920,N_1486,N_1502);
nor U1921 (N_1921,N_1539,N_1326);
xor U1922 (N_1922,N_1759,N_1497);
nor U1923 (N_1923,N_1619,N_1641);
nor U1924 (N_1924,N_1718,N_1729);
nor U1925 (N_1925,N_1300,N_1375);
nor U1926 (N_1926,N_1634,N_1417);
nor U1927 (N_1927,N_1452,N_1290);
or U1928 (N_1928,N_1420,N_1295);
xnor U1929 (N_1929,N_1257,N_1777);
and U1930 (N_1930,N_1475,N_1494);
xnor U1931 (N_1931,N_1505,N_1430);
xnor U1932 (N_1932,N_1481,N_1683);
or U1933 (N_1933,N_1741,N_1428);
nand U1934 (N_1934,N_1563,N_1392);
and U1935 (N_1935,N_1456,N_1569);
or U1936 (N_1936,N_1272,N_1439);
xor U1937 (N_1937,N_1547,N_1570);
or U1938 (N_1938,N_1255,N_1598);
xnor U1939 (N_1939,N_1599,N_1604);
and U1940 (N_1940,N_1394,N_1792);
nor U1941 (N_1941,N_1756,N_1523);
xnor U1942 (N_1942,N_1247,N_1697);
nand U1943 (N_1943,N_1349,N_1785);
nor U1944 (N_1944,N_1361,N_1200);
nand U1945 (N_1945,N_1427,N_1515);
and U1946 (N_1946,N_1222,N_1500);
nand U1947 (N_1947,N_1455,N_1464);
nor U1948 (N_1948,N_1304,N_1629);
nor U1949 (N_1949,N_1631,N_1299);
nor U1950 (N_1950,N_1687,N_1594);
nand U1951 (N_1951,N_1707,N_1580);
or U1952 (N_1952,N_1489,N_1406);
xor U1953 (N_1953,N_1373,N_1328);
or U1954 (N_1954,N_1291,N_1412);
nand U1955 (N_1955,N_1356,N_1637);
xnor U1956 (N_1956,N_1695,N_1329);
nor U1957 (N_1957,N_1747,N_1437);
nand U1958 (N_1958,N_1467,N_1223);
xnor U1959 (N_1959,N_1586,N_1408);
xor U1960 (N_1960,N_1224,N_1644);
xor U1961 (N_1961,N_1379,N_1562);
xnor U1962 (N_1962,N_1274,N_1658);
nand U1963 (N_1963,N_1298,N_1743);
or U1964 (N_1964,N_1566,N_1346);
and U1965 (N_1965,N_1688,N_1775);
xnor U1966 (N_1966,N_1774,N_1239);
nand U1967 (N_1967,N_1676,N_1354);
or U1968 (N_1968,N_1705,N_1768);
and U1969 (N_1969,N_1201,N_1431);
and U1970 (N_1970,N_1595,N_1591);
and U1971 (N_1971,N_1405,N_1652);
nand U1972 (N_1972,N_1510,N_1238);
or U1973 (N_1973,N_1587,N_1232);
xnor U1974 (N_1974,N_1560,N_1395);
nand U1975 (N_1975,N_1542,N_1568);
nand U1976 (N_1976,N_1673,N_1675);
nor U1977 (N_1977,N_1753,N_1337);
and U1978 (N_1978,N_1205,N_1443);
nand U1979 (N_1979,N_1684,N_1769);
or U1980 (N_1980,N_1305,N_1459);
and U1981 (N_1981,N_1789,N_1363);
and U1982 (N_1982,N_1519,N_1301);
and U1983 (N_1983,N_1445,N_1779);
xnor U1984 (N_1984,N_1335,N_1306);
and U1985 (N_1985,N_1765,N_1620);
nor U1986 (N_1986,N_1400,N_1258);
and U1987 (N_1987,N_1528,N_1530);
nor U1988 (N_1988,N_1706,N_1309);
or U1989 (N_1989,N_1237,N_1602);
xnor U1990 (N_1990,N_1654,N_1307);
nor U1991 (N_1991,N_1203,N_1526);
nand U1992 (N_1992,N_1553,N_1781);
xor U1993 (N_1993,N_1533,N_1754);
nor U1994 (N_1994,N_1415,N_1357);
or U1995 (N_1995,N_1468,N_1230);
or U1996 (N_1996,N_1532,N_1214);
nor U1997 (N_1997,N_1506,N_1630);
or U1998 (N_1998,N_1745,N_1277);
nand U1999 (N_1999,N_1627,N_1319);
and U2000 (N_2000,N_1491,N_1204);
or U2001 (N_2001,N_1498,N_1490);
nand U2002 (N_2002,N_1399,N_1438);
or U2003 (N_2003,N_1693,N_1712);
and U2004 (N_2004,N_1615,N_1504);
nand U2005 (N_2005,N_1260,N_1359);
nor U2006 (N_2006,N_1249,N_1318);
xnor U2007 (N_2007,N_1402,N_1294);
nor U2008 (N_2008,N_1334,N_1716);
and U2009 (N_2009,N_1679,N_1471);
and U2010 (N_2010,N_1466,N_1364);
xnor U2011 (N_2011,N_1565,N_1653);
xnor U2012 (N_2012,N_1338,N_1404);
xor U2013 (N_2013,N_1548,N_1686);
nor U2014 (N_2014,N_1261,N_1655);
nor U2015 (N_2015,N_1228,N_1749);
nor U2016 (N_2016,N_1245,N_1788);
xnor U2017 (N_2017,N_1478,N_1262);
xor U2018 (N_2018,N_1596,N_1320);
or U2019 (N_2019,N_1698,N_1681);
or U2020 (N_2020,N_1721,N_1287);
nor U2021 (N_2021,N_1760,N_1518);
nor U2022 (N_2022,N_1649,N_1374);
and U2023 (N_2023,N_1643,N_1534);
nand U2024 (N_2024,N_1446,N_1341);
or U2025 (N_2025,N_1432,N_1696);
and U2026 (N_2026,N_1323,N_1742);
or U2027 (N_2027,N_1512,N_1278);
nand U2028 (N_2028,N_1527,N_1552);
and U2029 (N_2029,N_1270,N_1770);
nand U2030 (N_2030,N_1391,N_1216);
nand U2031 (N_2031,N_1622,N_1267);
xnor U2032 (N_2032,N_1339,N_1344);
or U2033 (N_2033,N_1669,N_1545);
and U2034 (N_2034,N_1398,N_1317);
and U2035 (N_2035,N_1244,N_1240);
and U2036 (N_2036,N_1613,N_1382);
and U2037 (N_2037,N_1384,N_1493);
nand U2038 (N_2038,N_1259,N_1460);
or U2039 (N_2039,N_1720,N_1608);
and U2040 (N_2040,N_1734,N_1396);
nand U2041 (N_2041,N_1647,N_1571);
and U2042 (N_2042,N_1457,N_1730);
xnor U2043 (N_2043,N_1715,N_1605);
nor U2044 (N_2044,N_1517,N_1280);
or U2045 (N_2045,N_1413,N_1672);
xor U2046 (N_2046,N_1343,N_1345);
nor U2047 (N_2047,N_1226,N_1541);
nor U2048 (N_2048,N_1225,N_1513);
nand U2049 (N_2049,N_1601,N_1625);
xnor U2050 (N_2050,N_1664,N_1480);
nand U2051 (N_2051,N_1626,N_1725);
xnor U2052 (N_2052,N_1546,N_1612);
and U2053 (N_2053,N_1556,N_1458);
nand U2054 (N_2054,N_1302,N_1549);
nor U2055 (N_2055,N_1288,N_1646);
nand U2056 (N_2056,N_1787,N_1680);
nand U2057 (N_2057,N_1275,N_1227);
nand U2058 (N_2058,N_1434,N_1668);
or U2059 (N_2059,N_1722,N_1559);
xor U2060 (N_2060,N_1558,N_1385);
nor U2061 (N_2061,N_1799,N_1650);
nand U2062 (N_2062,N_1624,N_1632);
and U2063 (N_2063,N_1401,N_1414);
nor U2064 (N_2064,N_1589,N_1740);
or U2065 (N_2065,N_1212,N_1234);
and U2066 (N_2066,N_1583,N_1524);
xnor U2067 (N_2067,N_1661,N_1651);
nor U2068 (N_2068,N_1377,N_1531);
nor U2069 (N_2069,N_1482,N_1435);
nor U2070 (N_2070,N_1221,N_1322);
nor U2071 (N_2071,N_1242,N_1798);
xnor U2072 (N_2072,N_1733,N_1425);
nand U2073 (N_2073,N_1610,N_1440);
or U2074 (N_2074,N_1312,N_1282);
xnor U2075 (N_2075,N_1390,N_1479);
or U2076 (N_2076,N_1761,N_1645);
and U2077 (N_2077,N_1543,N_1215);
xnor U2078 (N_2078,N_1355,N_1691);
nor U2079 (N_2079,N_1310,N_1525);
nor U2080 (N_2080,N_1719,N_1724);
xnor U2081 (N_2081,N_1723,N_1520);
nor U2082 (N_2082,N_1786,N_1311);
or U2083 (N_2083,N_1484,N_1665);
xor U2084 (N_2084,N_1784,N_1289);
nand U2085 (N_2085,N_1521,N_1340);
and U2086 (N_2086,N_1426,N_1600);
or U2087 (N_2087,N_1397,N_1378);
nand U2088 (N_2088,N_1593,N_1710);
or U2089 (N_2089,N_1703,N_1487);
nor U2090 (N_2090,N_1461,N_1621);
or U2091 (N_2091,N_1732,N_1717);
or U2092 (N_2092,N_1292,N_1283);
nor U2093 (N_2093,N_1485,N_1611);
or U2094 (N_2094,N_1208,N_1764);
or U2095 (N_2095,N_1609,N_1648);
nand U2096 (N_2096,N_1332,N_1235);
nand U2097 (N_2097,N_1592,N_1746);
and U2098 (N_2098,N_1448,N_1639);
nand U2099 (N_2099,N_1573,N_1574);
nor U2100 (N_2100,N_1698,N_1238);
nor U2101 (N_2101,N_1549,N_1655);
or U2102 (N_2102,N_1753,N_1376);
or U2103 (N_2103,N_1630,N_1613);
nand U2104 (N_2104,N_1565,N_1419);
or U2105 (N_2105,N_1757,N_1376);
and U2106 (N_2106,N_1579,N_1598);
and U2107 (N_2107,N_1505,N_1473);
nor U2108 (N_2108,N_1259,N_1609);
and U2109 (N_2109,N_1392,N_1716);
nor U2110 (N_2110,N_1229,N_1739);
and U2111 (N_2111,N_1331,N_1517);
xor U2112 (N_2112,N_1382,N_1252);
and U2113 (N_2113,N_1579,N_1739);
nand U2114 (N_2114,N_1277,N_1798);
nand U2115 (N_2115,N_1797,N_1623);
nand U2116 (N_2116,N_1644,N_1559);
and U2117 (N_2117,N_1598,N_1643);
xor U2118 (N_2118,N_1476,N_1750);
nand U2119 (N_2119,N_1400,N_1396);
nand U2120 (N_2120,N_1409,N_1336);
or U2121 (N_2121,N_1519,N_1371);
nor U2122 (N_2122,N_1492,N_1643);
nand U2123 (N_2123,N_1480,N_1344);
and U2124 (N_2124,N_1797,N_1443);
nand U2125 (N_2125,N_1266,N_1513);
nor U2126 (N_2126,N_1573,N_1540);
xnor U2127 (N_2127,N_1406,N_1214);
nor U2128 (N_2128,N_1746,N_1541);
and U2129 (N_2129,N_1676,N_1580);
xnor U2130 (N_2130,N_1383,N_1789);
xor U2131 (N_2131,N_1227,N_1262);
and U2132 (N_2132,N_1456,N_1691);
and U2133 (N_2133,N_1578,N_1649);
nor U2134 (N_2134,N_1620,N_1764);
and U2135 (N_2135,N_1436,N_1364);
nand U2136 (N_2136,N_1444,N_1521);
and U2137 (N_2137,N_1415,N_1529);
or U2138 (N_2138,N_1651,N_1392);
xor U2139 (N_2139,N_1708,N_1276);
xor U2140 (N_2140,N_1759,N_1575);
nand U2141 (N_2141,N_1555,N_1675);
and U2142 (N_2142,N_1266,N_1358);
and U2143 (N_2143,N_1265,N_1370);
and U2144 (N_2144,N_1439,N_1751);
xnor U2145 (N_2145,N_1398,N_1586);
nand U2146 (N_2146,N_1520,N_1302);
nor U2147 (N_2147,N_1331,N_1752);
and U2148 (N_2148,N_1407,N_1624);
nand U2149 (N_2149,N_1719,N_1797);
xnor U2150 (N_2150,N_1606,N_1421);
and U2151 (N_2151,N_1482,N_1317);
nor U2152 (N_2152,N_1373,N_1529);
nor U2153 (N_2153,N_1296,N_1509);
nand U2154 (N_2154,N_1474,N_1205);
or U2155 (N_2155,N_1338,N_1709);
xnor U2156 (N_2156,N_1753,N_1349);
nand U2157 (N_2157,N_1403,N_1255);
nand U2158 (N_2158,N_1464,N_1406);
nand U2159 (N_2159,N_1606,N_1438);
and U2160 (N_2160,N_1386,N_1456);
nand U2161 (N_2161,N_1328,N_1536);
nor U2162 (N_2162,N_1426,N_1705);
nand U2163 (N_2163,N_1450,N_1358);
nand U2164 (N_2164,N_1733,N_1603);
nand U2165 (N_2165,N_1533,N_1613);
nand U2166 (N_2166,N_1706,N_1453);
and U2167 (N_2167,N_1249,N_1486);
or U2168 (N_2168,N_1236,N_1458);
nor U2169 (N_2169,N_1483,N_1687);
or U2170 (N_2170,N_1507,N_1732);
xor U2171 (N_2171,N_1627,N_1469);
nand U2172 (N_2172,N_1381,N_1710);
or U2173 (N_2173,N_1257,N_1472);
xor U2174 (N_2174,N_1379,N_1690);
or U2175 (N_2175,N_1738,N_1525);
xor U2176 (N_2176,N_1781,N_1417);
and U2177 (N_2177,N_1777,N_1577);
xor U2178 (N_2178,N_1506,N_1473);
and U2179 (N_2179,N_1704,N_1387);
or U2180 (N_2180,N_1358,N_1457);
or U2181 (N_2181,N_1239,N_1482);
xor U2182 (N_2182,N_1246,N_1717);
xnor U2183 (N_2183,N_1752,N_1520);
xor U2184 (N_2184,N_1203,N_1502);
xor U2185 (N_2185,N_1271,N_1323);
nor U2186 (N_2186,N_1374,N_1723);
nand U2187 (N_2187,N_1685,N_1320);
and U2188 (N_2188,N_1559,N_1407);
xor U2189 (N_2189,N_1450,N_1399);
xor U2190 (N_2190,N_1629,N_1560);
and U2191 (N_2191,N_1312,N_1424);
and U2192 (N_2192,N_1650,N_1765);
and U2193 (N_2193,N_1551,N_1671);
nand U2194 (N_2194,N_1362,N_1395);
xor U2195 (N_2195,N_1736,N_1249);
or U2196 (N_2196,N_1390,N_1481);
and U2197 (N_2197,N_1527,N_1486);
xnor U2198 (N_2198,N_1308,N_1577);
or U2199 (N_2199,N_1659,N_1457);
nand U2200 (N_2200,N_1793,N_1571);
xnor U2201 (N_2201,N_1378,N_1774);
and U2202 (N_2202,N_1491,N_1600);
xnor U2203 (N_2203,N_1625,N_1795);
nand U2204 (N_2204,N_1446,N_1759);
or U2205 (N_2205,N_1463,N_1389);
nor U2206 (N_2206,N_1266,N_1317);
and U2207 (N_2207,N_1374,N_1552);
nor U2208 (N_2208,N_1245,N_1676);
nand U2209 (N_2209,N_1589,N_1741);
nor U2210 (N_2210,N_1322,N_1254);
nand U2211 (N_2211,N_1301,N_1204);
or U2212 (N_2212,N_1773,N_1505);
nor U2213 (N_2213,N_1325,N_1414);
xnor U2214 (N_2214,N_1758,N_1513);
nand U2215 (N_2215,N_1772,N_1433);
nand U2216 (N_2216,N_1473,N_1708);
and U2217 (N_2217,N_1380,N_1375);
nand U2218 (N_2218,N_1435,N_1745);
nor U2219 (N_2219,N_1277,N_1390);
nor U2220 (N_2220,N_1609,N_1649);
nor U2221 (N_2221,N_1760,N_1532);
and U2222 (N_2222,N_1546,N_1605);
nand U2223 (N_2223,N_1514,N_1752);
xor U2224 (N_2224,N_1733,N_1372);
and U2225 (N_2225,N_1282,N_1249);
xnor U2226 (N_2226,N_1230,N_1778);
xor U2227 (N_2227,N_1256,N_1612);
and U2228 (N_2228,N_1401,N_1208);
nand U2229 (N_2229,N_1754,N_1597);
and U2230 (N_2230,N_1294,N_1533);
or U2231 (N_2231,N_1668,N_1473);
and U2232 (N_2232,N_1609,N_1435);
xor U2233 (N_2233,N_1288,N_1561);
nand U2234 (N_2234,N_1691,N_1617);
nand U2235 (N_2235,N_1371,N_1346);
or U2236 (N_2236,N_1632,N_1753);
nand U2237 (N_2237,N_1538,N_1413);
or U2238 (N_2238,N_1353,N_1233);
or U2239 (N_2239,N_1509,N_1281);
and U2240 (N_2240,N_1630,N_1511);
or U2241 (N_2241,N_1265,N_1429);
or U2242 (N_2242,N_1418,N_1791);
xor U2243 (N_2243,N_1639,N_1464);
xnor U2244 (N_2244,N_1279,N_1382);
or U2245 (N_2245,N_1213,N_1505);
nor U2246 (N_2246,N_1752,N_1344);
and U2247 (N_2247,N_1438,N_1353);
nor U2248 (N_2248,N_1799,N_1340);
and U2249 (N_2249,N_1426,N_1606);
nor U2250 (N_2250,N_1742,N_1759);
nand U2251 (N_2251,N_1716,N_1599);
nand U2252 (N_2252,N_1349,N_1435);
or U2253 (N_2253,N_1331,N_1454);
and U2254 (N_2254,N_1313,N_1666);
xor U2255 (N_2255,N_1331,N_1516);
and U2256 (N_2256,N_1286,N_1524);
or U2257 (N_2257,N_1369,N_1358);
xnor U2258 (N_2258,N_1612,N_1657);
and U2259 (N_2259,N_1799,N_1282);
and U2260 (N_2260,N_1379,N_1584);
nand U2261 (N_2261,N_1303,N_1778);
or U2262 (N_2262,N_1259,N_1637);
or U2263 (N_2263,N_1683,N_1652);
nand U2264 (N_2264,N_1512,N_1717);
nand U2265 (N_2265,N_1362,N_1257);
or U2266 (N_2266,N_1689,N_1782);
and U2267 (N_2267,N_1775,N_1410);
or U2268 (N_2268,N_1674,N_1455);
and U2269 (N_2269,N_1603,N_1329);
or U2270 (N_2270,N_1375,N_1638);
nand U2271 (N_2271,N_1579,N_1559);
or U2272 (N_2272,N_1784,N_1365);
or U2273 (N_2273,N_1255,N_1751);
nor U2274 (N_2274,N_1377,N_1245);
nand U2275 (N_2275,N_1658,N_1647);
xor U2276 (N_2276,N_1669,N_1539);
xor U2277 (N_2277,N_1254,N_1670);
or U2278 (N_2278,N_1399,N_1684);
xnor U2279 (N_2279,N_1384,N_1636);
xnor U2280 (N_2280,N_1351,N_1373);
and U2281 (N_2281,N_1275,N_1595);
nand U2282 (N_2282,N_1280,N_1535);
and U2283 (N_2283,N_1544,N_1767);
xnor U2284 (N_2284,N_1633,N_1513);
xor U2285 (N_2285,N_1537,N_1209);
and U2286 (N_2286,N_1550,N_1420);
and U2287 (N_2287,N_1699,N_1247);
and U2288 (N_2288,N_1788,N_1538);
xnor U2289 (N_2289,N_1206,N_1546);
or U2290 (N_2290,N_1385,N_1219);
and U2291 (N_2291,N_1542,N_1797);
nor U2292 (N_2292,N_1506,N_1588);
nor U2293 (N_2293,N_1441,N_1357);
or U2294 (N_2294,N_1487,N_1452);
and U2295 (N_2295,N_1610,N_1200);
or U2296 (N_2296,N_1455,N_1615);
or U2297 (N_2297,N_1420,N_1661);
nand U2298 (N_2298,N_1683,N_1555);
and U2299 (N_2299,N_1478,N_1263);
nand U2300 (N_2300,N_1473,N_1302);
nand U2301 (N_2301,N_1556,N_1554);
xnor U2302 (N_2302,N_1792,N_1392);
or U2303 (N_2303,N_1691,N_1309);
xor U2304 (N_2304,N_1708,N_1284);
nor U2305 (N_2305,N_1602,N_1335);
nor U2306 (N_2306,N_1319,N_1783);
nor U2307 (N_2307,N_1788,N_1768);
xor U2308 (N_2308,N_1549,N_1440);
nor U2309 (N_2309,N_1333,N_1536);
or U2310 (N_2310,N_1722,N_1241);
nor U2311 (N_2311,N_1520,N_1765);
or U2312 (N_2312,N_1239,N_1652);
nor U2313 (N_2313,N_1460,N_1665);
or U2314 (N_2314,N_1633,N_1225);
nor U2315 (N_2315,N_1640,N_1710);
xor U2316 (N_2316,N_1640,N_1483);
nand U2317 (N_2317,N_1269,N_1702);
and U2318 (N_2318,N_1681,N_1320);
nor U2319 (N_2319,N_1240,N_1689);
xnor U2320 (N_2320,N_1656,N_1550);
nor U2321 (N_2321,N_1793,N_1748);
and U2322 (N_2322,N_1240,N_1382);
or U2323 (N_2323,N_1493,N_1369);
xor U2324 (N_2324,N_1746,N_1507);
or U2325 (N_2325,N_1538,N_1630);
and U2326 (N_2326,N_1427,N_1200);
or U2327 (N_2327,N_1259,N_1366);
nand U2328 (N_2328,N_1697,N_1420);
or U2329 (N_2329,N_1450,N_1507);
and U2330 (N_2330,N_1432,N_1740);
nor U2331 (N_2331,N_1724,N_1576);
xnor U2332 (N_2332,N_1695,N_1526);
or U2333 (N_2333,N_1704,N_1756);
xnor U2334 (N_2334,N_1580,N_1496);
and U2335 (N_2335,N_1242,N_1237);
nand U2336 (N_2336,N_1722,N_1793);
or U2337 (N_2337,N_1495,N_1645);
or U2338 (N_2338,N_1445,N_1295);
and U2339 (N_2339,N_1446,N_1469);
nand U2340 (N_2340,N_1274,N_1451);
and U2341 (N_2341,N_1595,N_1336);
and U2342 (N_2342,N_1549,N_1509);
nor U2343 (N_2343,N_1414,N_1341);
or U2344 (N_2344,N_1392,N_1734);
nand U2345 (N_2345,N_1645,N_1484);
nand U2346 (N_2346,N_1599,N_1481);
nand U2347 (N_2347,N_1604,N_1755);
or U2348 (N_2348,N_1346,N_1480);
or U2349 (N_2349,N_1293,N_1377);
and U2350 (N_2350,N_1433,N_1290);
and U2351 (N_2351,N_1265,N_1581);
or U2352 (N_2352,N_1759,N_1597);
nor U2353 (N_2353,N_1798,N_1404);
and U2354 (N_2354,N_1374,N_1322);
nor U2355 (N_2355,N_1311,N_1349);
nor U2356 (N_2356,N_1451,N_1421);
nand U2357 (N_2357,N_1673,N_1528);
xor U2358 (N_2358,N_1256,N_1312);
nand U2359 (N_2359,N_1660,N_1335);
and U2360 (N_2360,N_1412,N_1694);
and U2361 (N_2361,N_1741,N_1492);
and U2362 (N_2362,N_1285,N_1668);
and U2363 (N_2363,N_1740,N_1280);
nor U2364 (N_2364,N_1769,N_1730);
nor U2365 (N_2365,N_1582,N_1353);
nor U2366 (N_2366,N_1548,N_1489);
nand U2367 (N_2367,N_1682,N_1663);
nand U2368 (N_2368,N_1779,N_1471);
xor U2369 (N_2369,N_1604,N_1717);
nand U2370 (N_2370,N_1478,N_1430);
and U2371 (N_2371,N_1310,N_1462);
and U2372 (N_2372,N_1411,N_1216);
nor U2373 (N_2373,N_1557,N_1445);
and U2374 (N_2374,N_1742,N_1527);
nand U2375 (N_2375,N_1548,N_1520);
nor U2376 (N_2376,N_1717,N_1731);
or U2377 (N_2377,N_1691,N_1536);
xnor U2378 (N_2378,N_1363,N_1722);
and U2379 (N_2379,N_1673,N_1437);
xor U2380 (N_2380,N_1557,N_1278);
xor U2381 (N_2381,N_1286,N_1450);
xnor U2382 (N_2382,N_1537,N_1677);
nor U2383 (N_2383,N_1278,N_1248);
and U2384 (N_2384,N_1498,N_1263);
nand U2385 (N_2385,N_1645,N_1310);
and U2386 (N_2386,N_1738,N_1452);
or U2387 (N_2387,N_1494,N_1559);
or U2388 (N_2388,N_1284,N_1505);
xor U2389 (N_2389,N_1285,N_1774);
or U2390 (N_2390,N_1358,N_1515);
nor U2391 (N_2391,N_1317,N_1442);
nor U2392 (N_2392,N_1584,N_1251);
xnor U2393 (N_2393,N_1736,N_1602);
nand U2394 (N_2394,N_1693,N_1596);
xor U2395 (N_2395,N_1515,N_1281);
nor U2396 (N_2396,N_1489,N_1688);
nand U2397 (N_2397,N_1233,N_1786);
nand U2398 (N_2398,N_1404,N_1723);
or U2399 (N_2399,N_1561,N_1647);
xnor U2400 (N_2400,N_1822,N_2276);
and U2401 (N_2401,N_2168,N_2235);
nor U2402 (N_2402,N_2019,N_2368);
and U2403 (N_2403,N_2215,N_2154);
or U2404 (N_2404,N_2031,N_2283);
or U2405 (N_2405,N_2218,N_2327);
nor U2406 (N_2406,N_1915,N_1943);
nand U2407 (N_2407,N_2393,N_1936);
xor U2408 (N_2408,N_2317,N_2272);
nand U2409 (N_2409,N_1950,N_1859);
xnor U2410 (N_2410,N_1885,N_2208);
xor U2411 (N_2411,N_2281,N_2319);
and U2412 (N_2412,N_2043,N_1980);
and U2413 (N_2413,N_2112,N_1972);
and U2414 (N_2414,N_1820,N_2381);
nand U2415 (N_2415,N_2057,N_2324);
nor U2416 (N_2416,N_2159,N_2022);
nor U2417 (N_2417,N_2238,N_2289);
xor U2418 (N_2418,N_2050,N_2329);
nor U2419 (N_2419,N_2243,N_1862);
nand U2420 (N_2420,N_1854,N_2037);
or U2421 (N_2421,N_1933,N_1864);
or U2422 (N_2422,N_2011,N_2309);
and U2423 (N_2423,N_2378,N_2035);
and U2424 (N_2424,N_2107,N_1964);
or U2425 (N_2425,N_1957,N_2148);
nor U2426 (N_2426,N_1994,N_2040);
nor U2427 (N_2427,N_2030,N_2396);
or U2428 (N_2428,N_1969,N_2217);
xor U2429 (N_2429,N_1937,N_2113);
and U2430 (N_2430,N_2267,N_2178);
or U2431 (N_2431,N_2055,N_2326);
xnor U2432 (N_2432,N_1981,N_2245);
xor U2433 (N_2433,N_2012,N_2117);
and U2434 (N_2434,N_1817,N_2349);
or U2435 (N_2435,N_2280,N_1938);
nand U2436 (N_2436,N_1845,N_2269);
xnor U2437 (N_2437,N_1842,N_2375);
nor U2438 (N_2438,N_2071,N_1805);
xor U2439 (N_2439,N_2146,N_2253);
or U2440 (N_2440,N_2015,N_2351);
nor U2441 (N_2441,N_2268,N_1987);
xor U2442 (N_2442,N_1877,N_2194);
nand U2443 (N_2443,N_2129,N_2209);
nor U2444 (N_2444,N_2322,N_2158);
xnor U2445 (N_2445,N_1837,N_2186);
xnor U2446 (N_2446,N_1801,N_1907);
nor U2447 (N_2447,N_2231,N_2001);
xnor U2448 (N_2448,N_2330,N_2152);
and U2449 (N_2449,N_2101,N_1997);
nand U2450 (N_2450,N_1894,N_2360);
xor U2451 (N_2451,N_2213,N_1939);
xor U2452 (N_2452,N_2345,N_2108);
or U2453 (N_2453,N_2032,N_1878);
nor U2454 (N_2454,N_2303,N_1865);
or U2455 (N_2455,N_2034,N_2192);
or U2456 (N_2456,N_1901,N_1883);
or U2457 (N_2457,N_2080,N_2257);
and U2458 (N_2458,N_2271,N_1852);
nor U2459 (N_2459,N_2197,N_1839);
nand U2460 (N_2460,N_2102,N_2149);
or U2461 (N_2461,N_2394,N_2198);
and U2462 (N_2462,N_1869,N_1947);
and U2463 (N_2463,N_2275,N_2005);
or U2464 (N_2464,N_2266,N_2084);
and U2465 (N_2465,N_2041,N_1944);
nor U2466 (N_2466,N_1841,N_1985);
nand U2467 (N_2467,N_2020,N_2377);
xnor U2468 (N_2468,N_2311,N_2036);
or U2469 (N_2469,N_2286,N_2325);
and U2470 (N_2470,N_1871,N_2111);
and U2471 (N_2471,N_2347,N_1892);
nand U2472 (N_2472,N_1829,N_2344);
and U2473 (N_2473,N_1932,N_1834);
or U2474 (N_2474,N_1840,N_2078);
xnor U2475 (N_2475,N_2167,N_2210);
xor U2476 (N_2476,N_2230,N_1831);
nand U2477 (N_2477,N_1904,N_2128);
or U2478 (N_2478,N_2014,N_2250);
nor U2479 (N_2479,N_2323,N_2026);
or U2480 (N_2480,N_1847,N_2132);
and U2481 (N_2481,N_2064,N_1867);
xnor U2482 (N_2482,N_2023,N_1940);
nor U2483 (N_2483,N_1818,N_2008);
and U2484 (N_2484,N_2067,N_1860);
and U2485 (N_2485,N_1898,N_2140);
nor U2486 (N_2486,N_2348,N_2359);
nor U2487 (N_2487,N_2364,N_2139);
xnor U2488 (N_2488,N_1993,N_1962);
and U2489 (N_2489,N_2273,N_1927);
and U2490 (N_2490,N_2018,N_1814);
nor U2491 (N_2491,N_2204,N_2358);
xnor U2492 (N_2492,N_2085,N_2258);
or U2493 (N_2493,N_1870,N_2278);
xor U2494 (N_2494,N_1951,N_1881);
xor U2495 (N_2495,N_2246,N_2335);
and U2496 (N_2496,N_2308,N_1849);
or U2497 (N_2497,N_1931,N_2033);
or U2498 (N_2498,N_2207,N_2390);
nand U2499 (N_2499,N_2371,N_2002);
nor U2500 (N_2500,N_1922,N_1916);
nand U2501 (N_2501,N_1807,N_2196);
or U2502 (N_2502,N_2341,N_2389);
nor U2503 (N_2503,N_2174,N_1813);
nand U2504 (N_2504,N_1953,N_2123);
or U2505 (N_2505,N_2116,N_1911);
or U2506 (N_2506,N_1821,N_2316);
nor U2507 (N_2507,N_1810,N_2180);
and U2508 (N_2508,N_2165,N_2054);
nand U2509 (N_2509,N_2334,N_1857);
and U2510 (N_2510,N_2337,N_2095);
or U2511 (N_2511,N_2306,N_2096);
or U2512 (N_2512,N_2172,N_1971);
nand U2513 (N_2513,N_1966,N_2003);
or U2514 (N_2514,N_2224,N_1910);
and U2515 (N_2515,N_2321,N_2365);
nor U2516 (N_2516,N_2093,N_2259);
or U2517 (N_2517,N_2190,N_1887);
nand U2518 (N_2518,N_2133,N_1977);
and U2519 (N_2519,N_1844,N_1949);
xnor U2520 (N_2520,N_2274,N_2261);
or U2521 (N_2521,N_2297,N_2362);
or U2522 (N_2522,N_2070,N_2072);
xnor U2523 (N_2523,N_1815,N_1995);
xnor U2524 (N_2524,N_2075,N_2200);
nand U2525 (N_2525,N_2363,N_2162);
xor U2526 (N_2526,N_2328,N_2191);
and U2527 (N_2527,N_1986,N_2029);
nor U2528 (N_2528,N_1924,N_1923);
and U2529 (N_2529,N_1955,N_1876);
nand U2530 (N_2530,N_2109,N_2292);
xor U2531 (N_2531,N_2244,N_2024);
nor U2532 (N_2532,N_1999,N_1991);
nand U2533 (N_2533,N_2220,N_2179);
nor U2534 (N_2534,N_1976,N_2256);
xor U2535 (N_2535,N_2138,N_1975);
and U2536 (N_2536,N_1954,N_2212);
or U2537 (N_2537,N_2391,N_2193);
xnor U2538 (N_2538,N_2150,N_2287);
nand U2539 (N_2539,N_2352,N_2181);
xor U2540 (N_2540,N_2069,N_1811);
xnor U2541 (N_2541,N_1984,N_2232);
nor U2542 (N_2542,N_1982,N_2199);
nor U2543 (N_2543,N_1914,N_2300);
or U2544 (N_2544,N_1828,N_2115);
xor U2545 (N_2545,N_2277,N_1926);
nor U2546 (N_2546,N_2166,N_1921);
or U2547 (N_2547,N_2189,N_1956);
or U2548 (N_2548,N_2171,N_2373);
nand U2549 (N_2549,N_2065,N_2106);
or U2550 (N_2550,N_2385,N_2242);
nor U2551 (N_2551,N_2137,N_2114);
nand U2552 (N_2552,N_2060,N_2227);
or U2553 (N_2553,N_2157,N_2110);
xor U2554 (N_2554,N_2387,N_2290);
nand U2555 (N_2555,N_2270,N_1850);
or U2556 (N_2556,N_2251,N_2077);
nand U2557 (N_2557,N_2265,N_1800);
xor U2558 (N_2558,N_2136,N_2121);
nand U2559 (N_2559,N_2237,N_2384);
and U2560 (N_2560,N_1908,N_1802);
and U2561 (N_2561,N_1913,N_2051);
nor U2562 (N_2562,N_2331,N_2262);
xnor U2563 (N_2563,N_1965,N_1958);
xor U2564 (N_2564,N_2361,N_2376);
nand U2565 (N_2565,N_2062,N_2185);
and U2566 (N_2566,N_1882,N_1983);
nand U2567 (N_2567,N_2356,N_1930);
or U2568 (N_2568,N_1812,N_1906);
nor U2569 (N_2569,N_1928,N_2367);
or U2570 (N_2570,N_2169,N_1823);
nand U2571 (N_2571,N_2395,N_1884);
and U2572 (N_2572,N_1868,N_2017);
xor U2573 (N_2573,N_2059,N_2143);
nor U2574 (N_2574,N_1946,N_2013);
xnor U2575 (N_2575,N_2004,N_2058);
nor U2576 (N_2576,N_1886,N_1836);
xnor U2577 (N_2577,N_1934,N_1891);
xnor U2578 (N_2578,N_2155,N_2294);
nor U2579 (N_2579,N_2127,N_1959);
nor U2580 (N_2580,N_2130,N_1827);
xor U2581 (N_2581,N_2126,N_1967);
or U2582 (N_2582,N_2045,N_2228);
nand U2583 (N_2583,N_2254,N_1996);
and U2584 (N_2584,N_2214,N_1808);
and U2585 (N_2585,N_1905,N_1988);
and U2586 (N_2586,N_1896,N_1912);
and U2587 (N_2587,N_2061,N_2226);
nand U2588 (N_2588,N_2103,N_1968);
nand U2589 (N_2589,N_2343,N_2184);
nand U2590 (N_2590,N_1851,N_2006);
nor U2591 (N_2591,N_2177,N_2160);
and U2592 (N_2592,N_2225,N_2027);
nor U2593 (N_2593,N_2007,N_1816);
nor U2594 (N_2594,N_2163,N_2144);
nor U2595 (N_2595,N_2047,N_2142);
or U2596 (N_2596,N_2346,N_2288);
nand U2597 (N_2597,N_2120,N_2234);
xor U2598 (N_2598,N_2372,N_2170);
and U2599 (N_2599,N_1890,N_1832);
nand U2600 (N_2600,N_1889,N_2092);
and U2601 (N_2601,N_1853,N_2260);
xnor U2602 (N_2602,N_2336,N_1858);
or U2603 (N_2603,N_2241,N_1835);
or U2604 (N_2604,N_1929,N_2247);
xnor U2605 (N_2605,N_1843,N_2370);
nand U2606 (N_2606,N_1960,N_1963);
and U2607 (N_2607,N_2206,N_2151);
xnor U2608 (N_2608,N_1872,N_2314);
nor U2609 (N_2609,N_2091,N_2295);
nor U2610 (N_2610,N_1863,N_2074);
nand U2611 (N_2611,N_2118,N_1973);
nand U2612 (N_2612,N_2039,N_1948);
and U2613 (N_2613,N_2353,N_2105);
or U2614 (N_2614,N_2038,N_2307);
and U2615 (N_2615,N_1838,N_2125);
and U2616 (N_2616,N_2086,N_2182);
nand U2617 (N_2617,N_1879,N_2350);
nand U2618 (N_2618,N_2076,N_2399);
or U2619 (N_2619,N_2087,N_1806);
and U2620 (N_2620,N_1974,N_2122);
xor U2621 (N_2621,N_1846,N_2009);
xor U2622 (N_2622,N_2339,N_2318);
xnor U2623 (N_2623,N_1917,N_2049);
nand U2624 (N_2624,N_1918,N_1935);
nand U2625 (N_2625,N_2388,N_1925);
nand U2626 (N_2626,N_2223,N_2239);
nand U2627 (N_2627,N_2083,N_2383);
nand U2628 (N_2628,N_2028,N_1920);
or U2629 (N_2629,N_1990,N_1903);
nand U2630 (N_2630,N_2279,N_2380);
nor U2631 (N_2631,N_2342,N_2021);
nor U2632 (N_2632,N_2135,N_2134);
nand U2633 (N_2633,N_1866,N_2255);
nor U2634 (N_2634,N_2056,N_2221);
and U2635 (N_2635,N_2044,N_2183);
nor U2636 (N_2636,N_1826,N_2248);
nor U2637 (N_2637,N_2216,N_2355);
nor U2638 (N_2638,N_2285,N_2284);
xnor U2639 (N_2639,N_1970,N_2053);
xor U2640 (N_2640,N_2252,N_2392);
nor U2641 (N_2641,N_2298,N_2233);
xor U2642 (N_2642,N_2063,N_2161);
or U2643 (N_2643,N_1803,N_2097);
or U2644 (N_2644,N_2042,N_2124);
nand U2645 (N_2645,N_1919,N_1804);
nor U2646 (N_2646,N_2397,N_1833);
xnor U2647 (N_2647,N_1902,N_1961);
or U2648 (N_2648,N_1897,N_1873);
nor U2649 (N_2649,N_2340,N_2099);
or U2650 (N_2650,N_2305,N_1893);
nor U2651 (N_2651,N_2100,N_2203);
and U2652 (N_2652,N_2310,N_2240);
xnor U2653 (N_2653,N_2313,N_2131);
or U2654 (N_2654,N_2211,N_2293);
nand U2655 (N_2655,N_2374,N_2291);
nor U2656 (N_2656,N_1830,N_1945);
nor U2657 (N_2657,N_2052,N_2315);
nor U2658 (N_2658,N_2068,N_2164);
nand U2659 (N_2659,N_2141,N_2282);
and U2660 (N_2660,N_1861,N_1992);
xnor U2661 (N_2661,N_2089,N_2386);
nand U2662 (N_2662,N_2176,N_1855);
and U2663 (N_2663,N_1874,N_2299);
nor U2664 (N_2664,N_2382,N_1909);
nand U2665 (N_2665,N_2145,N_1952);
xnor U2666 (N_2666,N_1848,N_1900);
or U2667 (N_2667,N_2236,N_2369);
xor U2668 (N_2668,N_2104,N_2357);
and U2669 (N_2669,N_2025,N_2202);
or U2670 (N_2670,N_2333,N_2090);
xor U2671 (N_2671,N_2195,N_2147);
xor U2672 (N_2672,N_2229,N_2188);
nand U2673 (N_2673,N_1825,N_2010);
nor U2674 (N_2674,N_1942,N_1989);
and U2675 (N_2675,N_2301,N_2338);
or U2676 (N_2676,N_2354,N_1856);
or U2677 (N_2677,N_2156,N_1875);
xnor U2678 (N_2678,N_2296,N_2048);
xor U2679 (N_2679,N_2119,N_2332);
xnor U2680 (N_2680,N_1899,N_2082);
or U2681 (N_2681,N_2153,N_1880);
or U2682 (N_2682,N_2366,N_2249);
nor U2683 (N_2683,N_2219,N_1979);
and U2684 (N_2684,N_2088,N_2264);
nor U2685 (N_2685,N_2000,N_2046);
nor U2686 (N_2686,N_2175,N_2398);
nand U2687 (N_2687,N_2304,N_1809);
and U2688 (N_2688,N_1941,N_1824);
nand U2689 (N_2689,N_1895,N_2173);
or U2690 (N_2690,N_2079,N_1819);
nand U2691 (N_2691,N_2187,N_1978);
xor U2692 (N_2692,N_2201,N_2302);
or U2693 (N_2693,N_2016,N_1998);
and U2694 (N_2694,N_2222,N_2263);
and U2695 (N_2695,N_2073,N_2379);
nor U2696 (N_2696,N_1888,N_2081);
and U2697 (N_2697,N_2094,N_2098);
and U2698 (N_2698,N_2320,N_2205);
xor U2699 (N_2699,N_2066,N_2312);
nor U2700 (N_2700,N_2001,N_2337);
nor U2701 (N_2701,N_1995,N_2126);
xnor U2702 (N_2702,N_1854,N_2171);
nor U2703 (N_2703,N_2114,N_1918);
xor U2704 (N_2704,N_2220,N_2325);
or U2705 (N_2705,N_2284,N_2068);
or U2706 (N_2706,N_2322,N_2108);
and U2707 (N_2707,N_1952,N_1867);
or U2708 (N_2708,N_1833,N_1988);
nand U2709 (N_2709,N_1883,N_2289);
or U2710 (N_2710,N_2374,N_2087);
xor U2711 (N_2711,N_2200,N_1802);
or U2712 (N_2712,N_1975,N_1954);
or U2713 (N_2713,N_2237,N_1986);
and U2714 (N_2714,N_2364,N_2192);
or U2715 (N_2715,N_2211,N_1914);
nand U2716 (N_2716,N_2172,N_1852);
nand U2717 (N_2717,N_2091,N_1872);
nor U2718 (N_2718,N_2305,N_2194);
xor U2719 (N_2719,N_2081,N_2369);
and U2720 (N_2720,N_2205,N_2039);
or U2721 (N_2721,N_2315,N_2313);
nor U2722 (N_2722,N_2103,N_2354);
nand U2723 (N_2723,N_1994,N_1888);
nor U2724 (N_2724,N_2064,N_1977);
and U2725 (N_2725,N_2180,N_2314);
and U2726 (N_2726,N_2270,N_2205);
nor U2727 (N_2727,N_1960,N_2236);
or U2728 (N_2728,N_1936,N_2144);
nand U2729 (N_2729,N_2028,N_2370);
or U2730 (N_2730,N_2145,N_1866);
and U2731 (N_2731,N_2039,N_1898);
nor U2732 (N_2732,N_1948,N_2336);
or U2733 (N_2733,N_1856,N_2218);
nand U2734 (N_2734,N_2198,N_1965);
and U2735 (N_2735,N_2379,N_1882);
and U2736 (N_2736,N_2320,N_1995);
xor U2737 (N_2737,N_1826,N_2144);
xor U2738 (N_2738,N_1980,N_2054);
xor U2739 (N_2739,N_1815,N_2223);
or U2740 (N_2740,N_2110,N_1853);
nand U2741 (N_2741,N_1844,N_2009);
nand U2742 (N_2742,N_2226,N_2217);
xor U2743 (N_2743,N_1964,N_2369);
nor U2744 (N_2744,N_2022,N_1864);
or U2745 (N_2745,N_2217,N_1808);
nor U2746 (N_2746,N_2288,N_2175);
nor U2747 (N_2747,N_2063,N_2180);
nand U2748 (N_2748,N_2366,N_1897);
nor U2749 (N_2749,N_2338,N_2266);
nand U2750 (N_2750,N_2291,N_2164);
nor U2751 (N_2751,N_2253,N_1962);
nor U2752 (N_2752,N_1888,N_2382);
and U2753 (N_2753,N_1998,N_1902);
nor U2754 (N_2754,N_1962,N_1989);
or U2755 (N_2755,N_1897,N_2268);
nand U2756 (N_2756,N_1933,N_2124);
or U2757 (N_2757,N_1848,N_2312);
and U2758 (N_2758,N_1853,N_2271);
and U2759 (N_2759,N_2209,N_2176);
or U2760 (N_2760,N_1926,N_2178);
xnor U2761 (N_2761,N_2038,N_1830);
nand U2762 (N_2762,N_2331,N_2388);
or U2763 (N_2763,N_2051,N_1851);
or U2764 (N_2764,N_2282,N_1980);
and U2765 (N_2765,N_1929,N_2124);
or U2766 (N_2766,N_2244,N_2217);
and U2767 (N_2767,N_2398,N_2183);
or U2768 (N_2768,N_2365,N_2357);
and U2769 (N_2769,N_2220,N_2049);
and U2770 (N_2770,N_2109,N_1854);
nand U2771 (N_2771,N_1862,N_2368);
nand U2772 (N_2772,N_2230,N_2265);
xnor U2773 (N_2773,N_1840,N_2095);
and U2774 (N_2774,N_2321,N_2262);
xor U2775 (N_2775,N_2020,N_1816);
and U2776 (N_2776,N_1914,N_1927);
or U2777 (N_2777,N_2293,N_2020);
and U2778 (N_2778,N_2124,N_1939);
xnor U2779 (N_2779,N_2099,N_1860);
nor U2780 (N_2780,N_1991,N_1830);
xor U2781 (N_2781,N_2282,N_2396);
and U2782 (N_2782,N_2164,N_1832);
and U2783 (N_2783,N_2107,N_2307);
xor U2784 (N_2784,N_2343,N_2109);
and U2785 (N_2785,N_2056,N_2398);
xor U2786 (N_2786,N_2319,N_2101);
nor U2787 (N_2787,N_2174,N_1888);
xnor U2788 (N_2788,N_1966,N_2260);
or U2789 (N_2789,N_1938,N_2109);
xor U2790 (N_2790,N_2050,N_2251);
and U2791 (N_2791,N_1840,N_2258);
nand U2792 (N_2792,N_2135,N_2255);
and U2793 (N_2793,N_2277,N_1962);
or U2794 (N_2794,N_1807,N_1841);
and U2795 (N_2795,N_2012,N_2077);
xnor U2796 (N_2796,N_1925,N_2268);
and U2797 (N_2797,N_2038,N_1916);
xnor U2798 (N_2798,N_2234,N_1992);
and U2799 (N_2799,N_2101,N_1950);
or U2800 (N_2800,N_1852,N_2230);
nand U2801 (N_2801,N_1968,N_1861);
or U2802 (N_2802,N_1801,N_1966);
nor U2803 (N_2803,N_2219,N_1871);
and U2804 (N_2804,N_1871,N_2088);
and U2805 (N_2805,N_2222,N_2346);
xor U2806 (N_2806,N_1905,N_1840);
or U2807 (N_2807,N_2051,N_2084);
nand U2808 (N_2808,N_1981,N_2222);
nor U2809 (N_2809,N_1845,N_2302);
xor U2810 (N_2810,N_1884,N_2312);
nor U2811 (N_2811,N_1959,N_2072);
and U2812 (N_2812,N_1900,N_1876);
and U2813 (N_2813,N_2305,N_1810);
nand U2814 (N_2814,N_1840,N_2122);
nand U2815 (N_2815,N_1838,N_2189);
xnor U2816 (N_2816,N_2269,N_2190);
nand U2817 (N_2817,N_2248,N_2291);
xor U2818 (N_2818,N_2003,N_2215);
or U2819 (N_2819,N_2120,N_2176);
and U2820 (N_2820,N_2054,N_1849);
xor U2821 (N_2821,N_2185,N_1883);
or U2822 (N_2822,N_1873,N_2291);
xor U2823 (N_2823,N_2135,N_1839);
nor U2824 (N_2824,N_1882,N_2039);
nor U2825 (N_2825,N_2312,N_1995);
xnor U2826 (N_2826,N_1899,N_2045);
nor U2827 (N_2827,N_2139,N_2165);
and U2828 (N_2828,N_2238,N_1810);
and U2829 (N_2829,N_2277,N_2270);
nand U2830 (N_2830,N_2324,N_2235);
or U2831 (N_2831,N_2055,N_2284);
and U2832 (N_2832,N_1862,N_2050);
and U2833 (N_2833,N_2062,N_1807);
nand U2834 (N_2834,N_2387,N_2241);
or U2835 (N_2835,N_2285,N_2129);
and U2836 (N_2836,N_2323,N_1880);
and U2837 (N_2837,N_1949,N_1861);
xor U2838 (N_2838,N_2300,N_2040);
and U2839 (N_2839,N_2318,N_1853);
or U2840 (N_2840,N_2056,N_2089);
nor U2841 (N_2841,N_2245,N_2337);
or U2842 (N_2842,N_2080,N_2033);
xnor U2843 (N_2843,N_1849,N_2327);
or U2844 (N_2844,N_1996,N_2362);
and U2845 (N_2845,N_2196,N_2033);
nand U2846 (N_2846,N_2003,N_1944);
nor U2847 (N_2847,N_1911,N_2051);
and U2848 (N_2848,N_2278,N_1948);
nor U2849 (N_2849,N_2185,N_1936);
and U2850 (N_2850,N_2295,N_1890);
or U2851 (N_2851,N_2141,N_2087);
nor U2852 (N_2852,N_2155,N_2003);
nor U2853 (N_2853,N_2245,N_2335);
nor U2854 (N_2854,N_2223,N_1886);
nand U2855 (N_2855,N_1848,N_2212);
nor U2856 (N_2856,N_2321,N_2016);
xnor U2857 (N_2857,N_1899,N_2167);
nor U2858 (N_2858,N_2088,N_2174);
nand U2859 (N_2859,N_1851,N_2319);
nor U2860 (N_2860,N_1921,N_2285);
nand U2861 (N_2861,N_1978,N_1807);
nor U2862 (N_2862,N_2242,N_2065);
nand U2863 (N_2863,N_2164,N_2280);
and U2864 (N_2864,N_1823,N_2108);
nor U2865 (N_2865,N_1971,N_2147);
or U2866 (N_2866,N_1833,N_2239);
or U2867 (N_2867,N_2180,N_2047);
or U2868 (N_2868,N_1879,N_1867);
nor U2869 (N_2869,N_1809,N_2087);
or U2870 (N_2870,N_1917,N_1930);
or U2871 (N_2871,N_1965,N_2354);
nand U2872 (N_2872,N_2231,N_2365);
xor U2873 (N_2873,N_2299,N_2234);
nand U2874 (N_2874,N_2005,N_2196);
nor U2875 (N_2875,N_2049,N_2386);
nand U2876 (N_2876,N_2168,N_2068);
nand U2877 (N_2877,N_1998,N_2242);
or U2878 (N_2878,N_2195,N_2063);
and U2879 (N_2879,N_2140,N_1817);
nand U2880 (N_2880,N_2223,N_2209);
or U2881 (N_2881,N_2200,N_1976);
and U2882 (N_2882,N_2209,N_2226);
nand U2883 (N_2883,N_2252,N_2048);
nand U2884 (N_2884,N_1984,N_1844);
or U2885 (N_2885,N_2378,N_1847);
nor U2886 (N_2886,N_2367,N_2299);
or U2887 (N_2887,N_2313,N_1875);
xnor U2888 (N_2888,N_1884,N_2302);
nand U2889 (N_2889,N_1965,N_2318);
nor U2890 (N_2890,N_2357,N_2393);
xnor U2891 (N_2891,N_2115,N_1820);
or U2892 (N_2892,N_2275,N_2220);
and U2893 (N_2893,N_2383,N_2365);
xor U2894 (N_2894,N_2363,N_2225);
nor U2895 (N_2895,N_2271,N_2192);
nor U2896 (N_2896,N_2197,N_2002);
nor U2897 (N_2897,N_2340,N_2037);
xor U2898 (N_2898,N_2393,N_2027);
nand U2899 (N_2899,N_1890,N_2058);
and U2900 (N_2900,N_2228,N_1961);
and U2901 (N_2901,N_2086,N_2255);
xor U2902 (N_2902,N_2143,N_2169);
and U2903 (N_2903,N_1950,N_1968);
or U2904 (N_2904,N_1899,N_1994);
or U2905 (N_2905,N_2020,N_2086);
nand U2906 (N_2906,N_2354,N_2069);
or U2907 (N_2907,N_1906,N_2260);
nor U2908 (N_2908,N_2037,N_1900);
and U2909 (N_2909,N_1938,N_1916);
and U2910 (N_2910,N_1846,N_2105);
nand U2911 (N_2911,N_1904,N_2205);
xor U2912 (N_2912,N_2391,N_1874);
xor U2913 (N_2913,N_2325,N_2103);
or U2914 (N_2914,N_1902,N_2332);
nor U2915 (N_2915,N_1957,N_2257);
or U2916 (N_2916,N_2223,N_2285);
nand U2917 (N_2917,N_2258,N_1828);
nand U2918 (N_2918,N_2245,N_2287);
and U2919 (N_2919,N_1901,N_2073);
nor U2920 (N_2920,N_2015,N_2176);
and U2921 (N_2921,N_1991,N_1909);
or U2922 (N_2922,N_2231,N_2248);
or U2923 (N_2923,N_2011,N_1924);
and U2924 (N_2924,N_2118,N_1986);
xor U2925 (N_2925,N_2320,N_2111);
nand U2926 (N_2926,N_2379,N_1998);
xor U2927 (N_2927,N_2184,N_2163);
nor U2928 (N_2928,N_1824,N_2152);
and U2929 (N_2929,N_1840,N_2105);
or U2930 (N_2930,N_2289,N_2209);
nand U2931 (N_2931,N_2274,N_2139);
nand U2932 (N_2932,N_1921,N_1857);
xnor U2933 (N_2933,N_2007,N_1987);
nor U2934 (N_2934,N_1946,N_2381);
nand U2935 (N_2935,N_2107,N_2103);
xor U2936 (N_2936,N_2182,N_1805);
nand U2937 (N_2937,N_1923,N_1941);
nor U2938 (N_2938,N_2078,N_2250);
xnor U2939 (N_2939,N_2368,N_2263);
or U2940 (N_2940,N_1985,N_2252);
nor U2941 (N_2941,N_2019,N_1907);
and U2942 (N_2942,N_2163,N_2177);
or U2943 (N_2943,N_1803,N_2065);
xnor U2944 (N_2944,N_2336,N_2151);
and U2945 (N_2945,N_2397,N_1990);
xor U2946 (N_2946,N_1850,N_2112);
nand U2947 (N_2947,N_2305,N_1805);
and U2948 (N_2948,N_2056,N_2106);
or U2949 (N_2949,N_2050,N_2083);
xor U2950 (N_2950,N_2157,N_2239);
and U2951 (N_2951,N_2068,N_1930);
nor U2952 (N_2952,N_1962,N_2119);
nand U2953 (N_2953,N_2030,N_1839);
and U2954 (N_2954,N_1959,N_2066);
nand U2955 (N_2955,N_2066,N_2214);
nor U2956 (N_2956,N_2319,N_1918);
and U2957 (N_2957,N_1894,N_1822);
xnor U2958 (N_2958,N_2397,N_1845);
and U2959 (N_2959,N_1810,N_2121);
nor U2960 (N_2960,N_2344,N_2364);
nor U2961 (N_2961,N_2011,N_2355);
or U2962 (N_2962,N_1924,N_2092);
nand U2963 (N_2963,N_2021,N_2241);
and U2964 (N_2964,N_1840,N_1882);
and U2965 (N_2965,N_2088,N_1942);
xnor U2966 (N_2966,N_1964,N_2240);
and U2967 (N_2967,N_2174,N_2284);
and U2968 (N_2968,N_1827,N_2176);
and U2969 (N_2969,N_2367,N_2069);
xor U2970 (N_2970,N_2152,N_2392);
and U2971 (N_2971,N_2395,N_1835);
nand U2972 (N_2972,N_2371,N_2083);
nor U2973 (N_2973,N_1997,N_2331);
nand U2974 (N_2974,N_2083,N_1945);
nor U2975 (N_2975,N_1925,N_2021);
or U2976 (N_2976,N_1889,N_2049);
nor U2977 (N_2977,N_2382,N_2245);
nor U2978 (N_2978,N_2063,N_2184);
nor U2979 (N_2979,N_2195,N_2279);
and U2980 (N_2980,N_2297,N_1972);
nor U2981 (N_2981,N_1826,N_2281);
nand U2982 (N_2982,N_1808,N_2106);
nor U2983 (N_2983,N_2041,N_2033);
xnor U2984 (N_2984,N_2363,N_1924);
nor U2985 (N_2985,N_1835,N_1860);
nor U2986 (N_2986,N_1970,N_1972);
xor U2987 (N_2987,N_2325,N_1848);
xor U2988 (N_2988,N_2064,N_2130);
nand U2989 (N_2989,N_2276,N_1836);
nand U2990 (N_2990,N_1814,N_1849);
nor U2991 (N_2991,N_1952,N_2107);
or U2992 (N_2992,N_2133,N_1921);
xnor U2993 (N_2993,N_2102,N_2105);
or U2994 (N_2994,N_2304,N_2039);
nand U2995 (N_2995,N_2130,N_2095);
nand U2996 (N_2996,N_1814,N_2359);
and U2997 (N_2997,N_2359,N_2075);
or U2998 (N_2998,N_1895,N_1818);
or U2999 (N_2999,N_1827,N_1968);
nor UO_0 (O_0,N_2851,N_2854);
or UO_1 (O_1,N_2403,N_2775);
nand UO_2 (O_2,N_2913,N_2442);
nor UO_3 (O_3,N_2675,N_2724);
and UO_4 (O_4,N_2433,N_2762);
or UO_5 (O_5,N_2662,N_2964);
and UO_6 (O_6,N_2861,N_2549);
or UO_7 (O_7,N_2619,N_2535);
xor UO_8 (O_8,N_2435,N_2692);
or UO_9 (O_9,N_2527,N_2909);
nor UO_10 (O_10,N_2816,N_2559);
xnor UO_11 (O_11,N_2745,N_2994);
nor UO_12 (O_12,N_2834,N_2797);
or UO_13 (O_13,N_2479,N_2423);
xor UO_14 (O_14,N_2695,N_2783);
or UO_15 (O_15,N_2939,N_2575);
xor UO_16 (O_16,N_2464,N_2912);
or UO_17 (O_17,N_2924,N_2630);
and UO_18 (O_18,N_2734,N_2502);
nor UO_19 (O_19,N_2777,N_2709);
and UO_20 (O_20,N_2786,N_2910);
and UO_21 (O_21,N_2946,N_2426);
nand UO_22 (O_22,N_2576,N_2971);
or UO_23 (O_23,N_2699,N_2920);
and UO_24 (O_24,N_2658,N_2748);
or UO_25 (O_25,N_2635,N_2639);
and UO_26 (O_26,N_2523,N_2621);
xor UO_27 (O_27,N_2951,N_2989);
or UO_28 (O_28,N_2817,N_2430);
nor UO_29 (O_29,N_2967,N_2818);
and UO_30 (O_30,N_2450,N_2796);
or UO_31 (O_31,N_2992,N_2568);
xnor UO_32 (O_32,N_2809,N_2788);
or UO_33 (O_33,N_2585,N_2743);
xnor UO_34 (O_34,N_2518,N_2904);
nand UO_35 (O_35,N_2628,N_2470);
xnor UO_36 (O_36,N_2542,N_2750);
nor UO_37 (O_37,N_2729,N_2787);
nand UO_38 (O_38,N_2922,N_2570);
xor UO_39 (O_39,N_2666,N_2485);
nor UO_40 (O_40,N_2859,N_2804);
or UO_41 (O_41,N_2931,N_2451);
xor UO_42 (O_42,N_2521,N_2476);
or UO_43 (O_43,N_2401,N_2702);
and UO_44 (O_44,N_2896,N_2723);
or UO_45 (O_45,N_2656,N_2677);
nand UO_46 (O_46,N_2727,N_2615);
or UO_47 (O_47,N_2505,N_2599);
and UO_48 (O_48,N_2417,N_2751);
nor UO_49 (O_49,N_2540,N_2583);
nor UO_50 (O_50,N_2525,N_2932);
and UO_51 (O_51,N_2872,N_2508);
and UO_52 (O_52,N_2779,N_2892);
nor UO_53 (O_53,N_2721,N_2917);
xor UO_54 (O_54,N_2820,N_2986);
nand UO_55 (O_55,N_2482,N_2678);
nand UO_56 (O_56,N_2760,N_2554);
xnor UO_57 (O_57,N_2984,N_2857);
and UO_58 (O_58,N_2448,N_2815);
and UO_59 (O_59,N_2668,N_2853);
nor UO_60 (O_60,N_2586,N_2506);
nand UO_61 (O_61,N_2676,N_2694);
and UO_62 (O_62,N_2697,N_2819);
and UO_63 (O_63,N_2459,N_2772);
or UO_64 (O_64,N_2916,N_2925);
xor UO_65 (O_65,N_2940,N_2477);
and UO_66 (O_66,N_2611,N_2457);
or UO_67 (O_67,N_2564,N_2444);
nand UO_68 (O_68,N_2921,N_2773);
nand UO_69 (O_69,N_2483,N_2513);
or UO_70 (O_70,N_2858,N_2937);
and UO_71 (O_71,N_2891,N_2902);
nand UO_72 (O_72,N_2782,N_2973);
nand UO_73 (O_73,N_2999,N_2510);
xnor UO_74 (O_74,N_2860,N_2691);
xnor UO_75 (O_75,N_2453,N_2595);
xor UO_76 (O_76,N_2511,N_2597);
xnor UO_77 (O_77,N_2968,N_2446);
and UO_78 (O_78,N_2957,N_2997);
nand UO_79 (O_79,N_2841,N_2810);
or UO_80 (O_80,N_2991,N_2674);
or UO_81 (O_81,N_2722,N_2713);
nand UO_82 (O_82,N_2553,N_2660);
nand UO_83 (O_83,N_2731,N_2752);
nand UO_84 (O_84,N_2534,N_2962);
xnor UO_85 (O_85,N_2531,N_2929);
xnor UO_86 (O_86,N_2897,N_2785);
and UO_87 (O_87,N_2838,N_2411);
and UO_88 (O_88,N_2899,N_2715);
xnor UO_89 (O_89,N_2960,N_2689);
or UO_90 (O_90,N_2767,N_2687);
nand UO_91 (O_91,N_2831,N_2900);
nor UO_92 (O_92,N_2790,N_2494);
nand UO_93 (O_93,N_2690,N_2850);
or UO_94 (O_94,N_2529,N_2683);
nand UO_95 (O_95,N_2985,N_2768);
and UO_96 (O_96,N_2431,N_2871);
or UO_97 (O_97,N_2686,N_2799);
nand UO_98 (O_98,N_2737,N_2469);
nor UO_99 (O_99,N_2710,N_2617);
nand UO_100 (O_100,N_2906,N_2830);
and UO_101 (O_101,N_2606,N_2952);
xnor UO_102 (O_102,N_2927,N_2961);
nor UO_103 (O_103,N_2671,N_2682);
xnor UO_104 (O_104,N_2659,N_2440);
or UO_105 (O_105,N_2714,N_2524);
or UO_106 (O_106,N_2776,N_2551);
xnor UO_107 (O_107,N_2974,N_2942);
xnor UO_108 (O_108,N_2604,N_2918);
xnor UO_109 (O_109,N_2629,N_2579);
and UO_110 (O_110,N_2454,N_2837);
nor UO_111 (O_111,N_2996,N_2673);
nand UO_112 (O_112,N_2407,N_2811);
nand UO_113 (O_113,N_2725,N_2716);
and UO_114 (O_114,N_2624,N_2556);
or UO_115 (O_115,N_2712,N_2537);
nor UO_116 (O_116,N_2982,N_2574);
or UO_117 (O_117,N_2404,N_2565);
and UO_118 (O_118,N_2825,N_2626);
nor UO_119 (O_119,N_2744,N_2607);
nor UO_120 (O_120,N_2908,N_2756);
or UO_121 (O_121,N_2803,N_2732);
or UO_122 (O_122,N_2488,N_2949);
xor UO_123 (O_123,N_2515,N_2581);
nor UO_124 (O_124,N_2740,N_2526);
xnor UO_125 (O_125,N_2726,N_2418);
and UO_126 (O_126,N_2412,N_2907);
xor UO_127 (O_127,N_2684,N_2875);
or UO_128 (O_128,N_2465,N_2632);
and UO_129 (O_129,N_2852,N_2844);
xor UO_130 (O_130,N_2966,N_2594);
xnor UO_131 (O_131,N_2833,N_2636);
and UO_132 (O_132,N_2806,N_2481);
and UO_133 (O_133,N_2493,N_2763);
or UO_134 (O_134,N_2865,N_2990);
and UO_135 (O_135,N_2733,N_2774);
xnor UO_136 (O_136,N_2826,N_2500);
or UO_137 (O_137,N_2988,N_2823);
or UO_138 (O_138,N_2663,N_2958);
or UO_139 (O_139,N_2945,N_2846);
and UO_140 (O_140,N_2944,N_2573);
xnor UO_141 (O_141,N_2548,N_2580);
nand UO_142 (O_142,N_2864,N_2840);
nor UO_143 (O_143,N_2935,N_2601);
xnor UO_144 (O_144,N_2771,N_2679);
nor UO_145 (O_145,N_2784,N_2801);
nor UO_146 (O_146,N_2704,N_2643);
or UO_147 (O_147,N_2759,N_2592);
xnor UO_148 (O_148,N_2672,N_2600);
xor UO_149 (O_149,N_2693,N_2514);
and UO_150 (O_150,N_2648,N_2824);
nor UO_151 (O_151,N_2413,N_2923);
nand UO_152 (O_152,N_2654,N_2866);
nor UO_153 (O_153,N_2758,N_2447);
nor UO_154 (O_154,N_2764,N_2880);
or UO_155 (O_155,N_2463,N_2602);
nor UO_156 (O_156,N_2703,N_2953);
nor UO_157 (O_157,N_2855,N_2614);
xnor UO_158 (O_158,N_2425,N_2882);
and UO_159 (O_159,N_2998,N_2845);
nand UO_160 (O_160,N_2655,N_2577);
nand UO_161 (O_161,N_2983,N_2424);
and UO_162 (O_162,N_2888,N_2670);
nor UO_163 (O_163,N_2498,N_2653);
xnor UO_164 (O_164,N_2969,N_2761);
nand UO_165 (O_165,N_2749,N_2954);
nand UO_166 (O_166,N_2688,N_2955);
nand UO_167 (O_167,N_2685,N_2473);
or UO_168 (O_168,N_2598,N_2980);
xnor UO_169 (O_169,N_2795,N_2528);
and UO_170 (O_170,N_2416,N_2458);
or UO_171 (O_171,N_2665,N_2504);
nor UO_172 (O_172,N_2625,N_2769);
xnor UO_173 (O_173,N_2753,N_2428);
and UO_174 (O_174,N_2461,N_2455);
and UO_175 (O_175,N_2930,N_2868);
nor UO_176 (O_176,N_2589,N_2487);
and UO_177 (O_177,N_2647,N_2538);
and UO_178 (O_178,N_2836,N_2637);
nor UO_179 (O_179,N_2402,N_2813);
nor UO_180 (O_180,N_2432,N_2680);
nand UO_181 (O_181,N_2562,N_2541);
and UO_182 (O_182,N_2828,N_2445);
nor UO_183 (O_183,N_2472,N_2484);
and UO_184 (O_184,N_2452,N_2995);
nand UO_185 (O_185,N_2512,N_2429);
xnor UO_186 (O_186,N_2503,N_2972);
nand UO_187 (O_187,N_2478,N_2634);
and UO_188 (O_188,N_2754,N_2582);
xnor UO_189 (O_189,N_2856,N_2746);
nor UO_190 (O_190,N_2735,N_2893);
xnor UO_191 (O_191,N_2462,N_2843);
and UO_192 (O_192,N_2742,N_2947);
nand UO_193 (O_193,N_2561,N_2596);
nand UO_194 (O_194,N_2889,N_2890);
nor UO_195 (O_195,N_2622,N_2911);
nor UO_196 (O_196,N_2895,N_2842);
nand UO_197 (O_197,N_2547,N_2517);
or UO_198 (O_198,N_2495,N_2480);
nand UO_199 (O_199,N_2934,N_2489);
or UO_200 (O_200,N_2644,N_2884);
or UO_201 (O_201,N_2438,N_2827);
xnor UO_202 (O_202,N_2720,N_2701);
or UO_203 (O_203,N_2766,N_2590);
and UO_204 (O_204,N_2770,N_2791);
xor UO_205 (O_205,N_2566,N_2928);
nor UO_206 (O_206,N_2578,N_2550);
and UO_207 (O_207,N_2905,N_2543);
xor UO_208 (O_208,N_2456,N_2605);
nand UO_209 (O_209,N_2633,N_2886);
or UO_210 (O_210,N_2408,N_2400);
or UO_211 (O_211,N_2516,N_2497);
nand UO_212 (O_212,N_2981,N_2730);
and UO_213 (O_213,N_2747,N_2781);
nand UO_214 (O_214,N_2405,N_2977);
nand UO_215 (O_215,N_2419,N_2765);
nand UO_216 (O_216,N_2610,N_2422);
nor UO_217 (O_217,N_2616,N_2421);
nand UO_218 (O_218,N_2649,N_2593);
nand UO_219 (O_219,N_2708,N_2468);
or UO_220 (O_220,N_2466,N_2848);
or UO_221 (O_221,N_2420,N_2569);
nor UO_222 (O_222,N_2613,N_2976);
xor UO_223 (O_223,N_2664,N_2603);
xor UO_224 (O_224,N_2757,N_2807);
and UO_225 (O_225,N_2885,N_2443);
xor UO_226 (O_226,N_2645,N_2780);
nand UO_227 (O_227,N_2587,N_2975);
nand UO_228 (O_228,N_2965,N_2567);
and UO_229 (O_229,N_2427,N_2718);
and UO_230 (O_230,N_2956,N_2959);
xor UO_231 (O_231,N_2736,N_2698);
nor UO_232 (O_232,N_2835,N_2641);
nand UO_233 (O_233,N_2509,N_2609);
xnor UO_234 (O_234,N_2631,N_2406);
nor UO_235 (O_235,N_2873,N_2719);
nor UO_236 (O_236,N_2640,N_2874);
nor UO_237 (O_237,N_2862,N_2436);
and UO_238 (O_238,N_2546,N_2832);
or UO_239 (O_239,N_2938,N_2591);
and UO_240 (O_240,N_2970,N_2870);
and UO_241 (O_241,N_2642,N_2943);
nor UO_242 (O_242,N_2741,N_2987);
nor UO_243 (O_243,N_2558,N_2805);
or UO_244 (O_244,N_2474,N_2560);
or UO_245 (O_245,N_2486,N_2933);
xnor UO_246 (O_246,N_2792,N_2646);
nand UO_247 (O_247,N_2499,N_2681);
xor UO_248 (O_248,N_2867,N_2881);
and UO_249 (O_249,N_2555,N_2667);
and UO_250 (O_250,N_2434,N_2950);
xor UO_251 (O_251,N_2898,N_2963);
or UO_252 (O_252,N_2706,N_2941);
nor UO_253 (O_253,N_2492,N_2441);
nor UO_254 (O_254,N_2530,N_2661);
nand UO_255 (O_255,N_2869,N_2620);
nand UO_256 (O_256,N_2415,N_2496);
nand UO_257 (O_257,N_2449,N_2879);
or UO_258 (O_258,N_2812,N_2814);
xor UO_259 (O_259,N_2802,N_2738);
and UO_260 (O_260,N_2572,N_2728);
nor UO_261 (O_261,N_2901,N_2822);
nand UO_262 (O_262,N_2501,N_2849);
and UO_263 (O_263,N_2707,N_2490);
or UO_264 (O_264,N_2584,N_2739);
nor UO_265 (O_265,N_2808,N_2475);
xor UO_266 (O_266,N_2877,N_2519);
nor UO_267 (O_267,N_2948,N_2800);
nor UO_268 (O_268,N_2414,N_2700);
xor UO_269 (O_269,N_2979,N_2914);
nor UO_270 (O_270,N_2993,N_2711);
and UO_271 (O_271,N_2794,N_2847);
nor UO_272 (O_272,N_2544,N_2539);
nand UO_273 (O_273,N_2717,N_2552);
xor UO_274 (O_274,N_2520,N_2557);
or UO_275 (O_275,N_2878,N_2652);
nand UO_276 (O_276,N_2919,N_2793);
and UO_277 (O_277,N_2883,N_2650);
nor UO_278 (O_278,N_2533,N_2638);
and UO_279 (O_279,N_2978,N_2839);
xnor UO_280 (O_280,N_2627,N_2696);
nand UO_281 (O_281,N_2618,N_2439);
nand UO_282 (O_282,N_2588,N_2460);
nand UO_283 (O_283,N_2829,N_2612);
and UO_284 (O_284,N_2571,N_2936);
and UO_285 (O_285,N_2669,N_2522);
and UO_286 (O_286,N_2608,N_2410);
and UO_287 (O_287,N_2778,N_2887);
xnor UO_288 (O_288,N_2789,N_2471);
xor UO_289 (O_289,N_2755,N_2798);
nor UO_290 (O_290,N_2705,N_2623);
nor UO_291 (O_291,N_2903,N_2821);
nor UO_292 (O_292,N_2409,N_2657);
nand UO_293 (O_293,N_2536,N_2863);
or UO_294 (O_294,N_2491,N_2651);
xor UO_295 (O_295,N_2507,N_2532);
and UO_296 (O_296,N_2926,N_2545);
or UO_297 (O_297,N_2915,N_2437);
and UO_298 (O_298,N_2894,N_2876);
xor UO_299 (O_299,N_2467,N_2563);
or UO_300 (O_300,N_2961,N_2704);
or UO_301 (O_301,N_2557,N_2820);
nand UO_302 (O_302,N_2471,N_2418);
nand UO_303 (O_303,N_2421,N_2952);
xnor UO_304 (O_304,N_2758,N_2751);
and UO_305 (O_305,N_2623,N_2932);
and UO_306 (O_306,N_2796,N_2460);
and UO_307 (O_307,N_2415,N_2825);
or UO_308 (O_308,N_2610,N_2436);
nand UO_309 (O_309,N_2664,N_2709);
xor UO_310 (O_310,N_2991,N_2729);
nand UO_311 (O_311,N_2941,N_2608);
and UO_312 (O_312,N_2755,N_2530);
and UO_313 (O_313,N_2636,N_2475);
nor UO_314 (O_314,N_2694,N_2426);
and UO_315 (O_315,N_2889,N_2426);
and UO_316 (O_316,N_2569,N_2948);
and UO_317 (O_317,N_2583,N_2947);
xnor UO_318 (O_318,N_2539,N_2643);
nand UO_319 (O_319,N_2509,N_2691);
nor UO_320 (O_320,N_2996,N_2741);
and UO_321 (O_321,N_2496,N_2954);
and UO_322 (O_322,N_2660,N_2694);
xnor UO_323 (O_323,N_2514,N_2415);
xor UO_324 (O_324,N_2503,N_2506);
or UO_325 (O_325,N_2482,N_2754);
nand UO_326 (O_326,N_2931,N_2548);
and UO_327 (O_327,N_2573,N_2771);
or UO_328 (O_328,N_2432,N_2655);
or UO_329 (O_329,N_2943,N_2983);
xnor UO_330 (O_330,N_2618,N_2991);
nor UO_331 (O_331,N_2836,N_2897);
xnor UO_332 (O_332,N_2640,N_2993);
xnor UO_333 (O_333,N_2650,N_2426);
xnor UO_334 (O_334,N_2418,N_2682);
and UO_335 (O_335,N_2603,N_2898);
nand UO_336 (O_336,N_2705,N_2564);
nor UO_337 (O_337,N_2656,N_2923);
or UO_338 (O_338,N_2702,N_2917);
nand UO_339 (O_339,N_2952,N_2954);
or UO_340 (O_340,N_2618,N_2500);
nand UO_341 (O_341,N_2661,N_2629);
nand UO_342 (O_342,N_2646,N_2977);
and UO_343 (O_343,N_2498,N_2507);
and UO_344 (O_344,N_2836,N_2654);
xnor UO_345 (O_345,N_2433,N_2413);
or UO_346 (O_346,N_2750,N_2558);
nand UO_347 (O_347,N_2907,N_2519);
xnor UO_348 (O_348,N_2530,N_2662);
xnor UO_349 (O_349,N_2762,N_2728);
nor UO_350 (O_350,N_2438,N_2868);
xnor UO_351 (O_351,N_2454,N_2983);
nand UO_352 (O_352,N_2988,N_2903);
nor UO_353 (O_353,N_2823,N_2603);
nand UO_354 (O_354,N_2440,N_2612);
or UO_355 (O_355,N_2534,N_2661);
nand UO_356 (O_356,N_2553,N_2805);
and UO_357 (O_357,N_2681,N_2745);
nand UO_358 (O_358,N_2426,N_2898);
xnor UO_359 (O_359,N_2744,N_2833);
or UO_360 (O_360,N_2893,N_2655);
or UO_361 (O_361,N_2417,N_2721);
and UO_362 (O_362,N_2654,N_2917);
or UO_363 (O_363,N_2994,N_2404);
nand UO_364 (O_364,N_2610,N_2970);
xnor UO_365 (O_365,N_2889,N_2575);
and UO_366 (O_366,N_2918,N_2766);
nor UO_367 (O_367,N_2985,N_2988);
nor UO_368 (O_368,N_2673,N_2981);
or UO_369 (O_369,N_2896,N_2982);
nand UO_370 (O_370,N_2401,N_2820);
or UO_371 (O_371,N_2838,N_2918);
nand UO_372 (O_372,N_2617,N_2513);
nor UO_373 (O_373,N_2963,N_2427);
xnor UO_374 (O_374,N_2943,N_2661);
and UO_375 (O_375,N_2878,N_2561);
and UO_376 (O_376,N_2577,N_2766);
nand UO_377 (O_377,N_2616,N_2618);
and UO_378 (O_378,N_2645,N_2796);
nor UO_379 (O_379,N_2894,N_2521);
or UO_380 (O_380,N_2628,N_2835);
nand UO_381 (O_381,N_2791,N_2834);
or UO_382 (O_382,N_2619,N_2899);
nand UO_383 (O_383,N_2811,N_2615);
and UO_384 (O_384,N_2856,N_2456);
xnor UO_385 (O_385,N_2871,N_2544);
or UO_386 (O_386,N_2651,N_2824);
nand UO_387 (O_387,N_2405,N_2779);
and UO_388 (O_388,N_2417,N_2964);
or UO_389 (O_389,N_2469,N_2704);
nor UO_390 (O_390,N_2407,N_2587);
and UO_391 (O_391,N_2532,N_2458);
and UO_392 (O_392,N_2921,N_2816);
nor UO_393 (O_393,N_2506,N_2462);
xnor UO_394 (O_394,N_2631,N_2700);
and UO_395 (O_395,N_2836,N_2472);
nand UO_396 (O_396,N_2866,N_2474);
xnor UO_397 (O_397,N_2465,N_2562);
nand UO_398 (O_398,N_2802,N_2449);
xor UO_399 (O_399,N_2869,N_2408);
nand UO_400 (O_400,N_2876,N_2685);
and UO_401 (O_401,N_2488,N_2645);
or UO_402 (O_402,N_2612,N_2645);
nand UO_403 (O_403,N_2578,N_2488);
and UO_404 (O_404,N_2454,N_2953);
nand UO_405 (O_405,N_2677,N_2439);
or UO_406 (O_406,N_2561,N_2496);
nor UO_407 (O_407,N_2442,N_2952);
nand UO_408 (O_408,N_2443,N_2513);
and UO_409 (O_409,N_2590,N_2410);
nor UO_410 (O_410,N_2481,N_2478);
or UO_411 (O_411,N_2491,N_2947);
nor UO_412 (O_412,N_2565,N_2935);
and UO_413 (O_413,N_2869,N_2774);
and UO_414 (O_414,N_2999,N_2777);
nand UO_415 (O_415,N_2435,N_2531);
nand UO_416 (O_416,N_2572,N_2736);
xnor UO_417 (O_417,N_2835,N_2795);
nor UO_418 (O_418,N_2404,N_2487);
nor UO_419 (O_419,N_2750,N_2868);
and UO_420 (O_420,N_2406,N_2605);
xnor UO_421 (O_421,N_2758,N_2448);
nand UO_422 (O_422,N_2767,N_2492);
and UO_423 (O_423,N_2656,N_2817);
and UO_424 (O_424,N_2878,N_2569);
or UO_425 (O_425,N_2996,N_2820);
and UO_426 (O_426,N_2874,N_2500);
xnor UO_427 (O_427,N_2990,N_2762);
nand UO_428 (O_428,N_2646,N_2834);
and UO_429 (O_429,N_2630,N_2636);
or UO_430 (O_430,N_2724,N_2533);
and UO_431 (O_431,N_2876,N_2731);
xor UO_432 (O_432,N_2545,N_2788);
xnor UO_433 (O_433,N_2985,N_2598);
and UO_434 (O_434,N_2886,N_2751);
or UO_435 (O_435,N_2951,N_2875);
xnor UO_436 (O_436,N_2400,N_2512);
nor UO_437 (O_437,N_2755,N_2568);
and UO_438 (O_438,N_2570,N_2619);
xnor UO_439 (O_439,N_2802,N_2824);
xnor UO_440 (O_440,N_2822,N_2436);
nor UO_441 (O_441,N_2781,N_2676);
xor UO_442 (O_442,N_2483,N_2898);
xnor UO_443 (O_443,N_2762,N_2677);
or UO_444 (O_444,N_2425,N_2786);
xor UO_445 (O_445,N_2469,N_2544);
nor UO_446 (O_446,N_2721,N_2965);
nor UO_447 (O_447,N_2429,N_2477);
and UO_448 (O_448,N_2744,N_2609);
xor UO_449 (O_449,N_2857,N_2842);
or UO_450 (O_450,N_2825,N_2493);
nand UO_451 (O_451,N_2588,N_2511);
nand UO_452 (O_452,N_2805,N_2930);
and UO_453 (O_453,N_2973,N_2944);
nor UO_454 (O_454,N_2480,N_2820);
nand UO_455 (O_455,N_2445,N_2707);
nor UO_456 (O_456,N_2850,N_2733);
nor UO_457 (O_457,N_2969,N_2538);
or UO_458 (O_458,N_2666,N_2888);
and UO_459 (O_459,N_2933,N_2527);
and UO_460 (O_460,N_2748,N_2512);
xnor UO_461 (O_461,N_2461,N_2751);
nor UO_462 (O_462,N_2758,N_2620);
or UO_463 (O_463,N_2475,N_2942);
or UO_464 (O_464,N_2719,N_2747);
and UO_465 (O_465,N_2598,N_2401);
or UO_466 (O_466,N_2964,N_2788);
and UO_467 (O_467,N_2824,N_2480);
nor UO_468 (O_468,N_2526,N_2620);
and UO_469 (O_469,N_2596,N_2641);
xnor UO_470 (O_470,N_2872,N_2818);
nand UO_471 (O_471,N_2701,N_2862);
and UO_472 (O_472,N_2829,N_2479);
nor UO_473 (O_473,N_2651,N_2764);
nor UO_474 (O_474,N_2654,N_2508);
nand UO_475 (O_475,N_2638,N_2872);
and UO_476 (O_476,N_2878,N_2472);
nand UO_477 (O_477,N_2440,N_2734);
and UO_478 (O_478,N_2892,N_2472);
and UO_479 (O_479,N_2606,N_2742);
xnor UO_480 (O_480,N_2421,N_2639);
xnor UO_481 (O_481,N_2645,N_2867);
and UO_482 (O_482,N_2452,N_2779);
or UO_483 (O_483,N_2473,N_2840);
nand UO_484 (O_484,N_2605,N_2829);
or UO_485 (O_485,N_2765,N_2935);
or UO_486 (O_486,N_2946,N_2957);
nor UO_487 (O_487,N_2951,N_2708);
and UO_488 (O_488,N_2453,N_2613);
or UO_489 (O_489,N_2668,N_2778);
nand UO_490 (O_490,N_2839,N_2473);
nor UO_491 (O_491,N_2789,N_2707);
xor UO_492 (O_492,N_2970,N_2495);
or UO_493 (O_493,N_2600,N_2487);
and UO_494 (O_494,N_2926,N_2547);
xnor UO_495 (O_495,N_2990,N_2482);
nor UO_496 (O_496,N_2737,N_2837);
nand UO_497 (O_497,N_2707,N_2494);
nand UO_498 (O_498,N_2847,N_2523);
nor UO_499 (O_499,N_2401,N_2987);
endmodule