module basic_1500_15000_2000_75_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_650,In_1064);
and U1 (N_1,In_450,In_1456);
xnor U2 (N_2,In_169,In_1463);
nand U3 (N_3,In_1472,In_936);
nand U4 (N_4,In_572,In_863);
xor U5 (N_5,In_1460,In_856);
nor U6 (N_6,In_758,In_503);
nand U7 (N_7,In_1226,In_1451);
or U8 (N_8,In_873,In_747);
or U9 (N_9,In_1297,In_1464);
nor U10 (N_10,In_826,In_1115);
or U11 (N_11,In_619,In_432);
xnor U12 (N_12,In_256,In_116);
nand U13 (N_13,In_1305,In_1254);
xor U14 (N_14,In_664,In_1408);
nor U15 (N_15,In_858,In_1103);
nand U16 (N_16,In_1112,In_1342);
nor U17 (N_17,In_1190,In_679);
and U18 (N_18,In_104,In_206);
or U19 (N_19,In_1309,In_906);
and U20 (N_20,In_469,In_234);
nand U21 (N_21,In_887,In_1113);
nor U22 (N_22,In_594,In_221);
nor U23 (N_23,In_959,In_1400);
nand U24 (N_24,In_45,In_1248);
and U25 (N_25,In_705,In_796);
xor U26 (N_26,In_1052,In_1024);
or U27 (N_27,In_485,In_702);
and U28 (N_28,In_1166,In_93);
xor U29 (N_29,In_542,In_1159);
nand U30 (N_30,In_516,In_480);
nand U31 (N_31,In_1427,In_12);
xnor U32 (N_32,In_937,In_431);
and U33 (N_33,In_211,In_591);
nand U34 (N_34,In_1345,In_554);
and U35 (N_35,In_1347,In_547);
nor U36 (N_36,In_556,In_706);
nand U37 (N_37,In_955,In_451);
nor U38 (N_38,In_945,In_230);
and U39 (N_39,In_721,In_1186);
or U40 (N_40,In_1374,In_571);
xnor U41 (N_41,In_583,In_1475);
and U42 (N_42,In_279,In_1327);
nand U43 (N_43,In_1319,In_1257);
nand U44 (N_44,In_267,In_1314);
nor U45 (N_45,In_1390,In_555);
nand U46 (N_46,In_271,In_889);
or U47 (N_47,In_818,In_1388);
xnor U48 (N_48,In_445,In_1195);
nand U49 (N_49,In_967,In_546);
xor U50 (N_50,In_335,In_1059);
and U51 (N_51,In_395,In_691);
nand U52 (N_52,In_139,In_154);
or U53 (N_53,In_607,In_807);
nand U54 (N_54,In_96,In_6);
xnor U55 (N_55,In_91,In_1157);
or U56 (N_56,In_440,In_566);
xnor U57 (N_57,In_668,In_36);
and U58 (N_58,In_895,In_1287);
nand U59 (N_59,In_749,In_609);
nand U60 (N_60,In_95,In_797);
or U61 (N_61,In_220,In_760);
nor U62 (N_62,In_928,In_1030);
xnor U63 (N_63,In_1466,In_852);
or U64 (N_64,In_606,In_208);
xnor U65 (N_65,In_444,In_1152);
or U66 (N_66,In_295,In_1209);
xor U67 (N_67,In_1416,In_73);
nor U68 (N_68,In_1184,In_316);
nand U69 (N_69,In_202,In_1362);
nor U70 (N_70,In_223,In_57);
or U71 (N_71,In_832,In_833);
nand U72 (N_72,In_184,In_370);
or U73 (N_73,In_380,In_1123);
nand U74 (N_74,In_1426,In_851);
nand U75 (N_75,In_1470,In_1106);
nand U76 (N_76,In_1155,In_918);
or U77 (N_77,In_938,In_155);
nand U78 (N_78,In_412,In_734);
nor U79 (N_79,In_1352,In_1358);
nor U80 (N_80,In_1205,In_199);
nor U81 (N_81,In_977,In_795);
xor U82 (N_82,In_1100,In_142);
nor U83 (N_83,In_47,In_1192);
and U84 (N_84,In_437,In_1108);
and U85 (N_85,In_631,In_381);
nor U86 (N_86,In_136,In_909);
nand U87 (N_87,In_1215,In_284);
xnor U88 (N_88,In_932,In_44);
xor U89 (N_89,In_1445,In_775);
nand U90 (N_90,In_1057,In_1334);
nor U91 (N_91,In_1165,In_342);
nor U92 (N_92,In_0,In_1138);
nand U93 (N_93,In_1019,In_931);
nand U94 (N_94,In_912,In_964);
and U95 (N_95,In_1410,In_343);
nand U96 (N_96,In_35,In_701);
nor U97 (N_97,In_182,In_1009);
nor U98 (N_98,In_152,In_946);
and U99 (N_99,In_528,In_1259);
xor U100 (N_100,In_739,In_193);
and U101 (N_101,In_737,In_697);
and U102 (N_102,In_1424,In_1494);
and U103 (N_103,In_2,In_905);
xnor U104 (N_104,In_1432,In_1102);
xnor U105 (N_105,In_1012,In_1137);
xnor U106 (N_106,In_733,In_29);
or U107 (N_107,In_332,In_892);
or U108 (N_108,In_249,In_785);
nor U109 (N_109,In_559,In_644);
nor U110 (N_110,In_1022,In_318);
or U111 (N_111,In_400,In_232);
and U112 (N_112,In_423,In_1167);
xor U113 (N_113,In_1295,In_416);
nand U114 (N_114,In_1007,In_1201);
and U115 (N_115,In_855,In_1114);
nor U116 (N_116,In_458,In_159);
nand U117 (N_117,In_1056,In_1070);
nor U118 (N_118,In_1061,In_1355);
or U119 (N_119,In_317,In_1476);
and U120 (N_120,In_551,In_1111);
or U121 (N_121,In_1117,In_518);
xnor U122 (N_122,In_859,In_1055);
nor U123 (N_123,In_903,In_1407);
and U124 (N_124,In_286,In_258);
xor U125 (N_125,In_237,In_327);
and U126 (N_126,In_1350,In_1083);
and U127 (N_127,In_1200,In_179);
xor U128 (N_128,In_1177,In_1373);
and U129 (N_129,In_686,In_470);
xnor U130 (N_130,In_465,In_790);
nand U131 (N_131,In_1044,In_1396);
xnor U132 (N_132,In_200,In_21);
xnor U133 (N_133,In_1037,In_974);
nor U134 (N_134,In_351,In_735);
nand U135 (N_135,In_862,In_1153);
and U136 (N_136,In_1339,In_1176);
xor U137 (N_137,In_369,In_756);
xnor U138 (N_138,In_798,In_118);
xor U139 (N_139,In_1238,In_1497);
xnor U140 (N_140,In_923,In_1285);
nor U141 (N_141,In_1054,In_751);
xnor U142 (N_142,In_865,In_1169);
nor U143 (N_143,In_1191,In_212);
and U144 (N_144,In_672,In_1130);
or U145 (N_145,In_553,In_127);
or U146 (N_146,In_1371,In_1178);
or U147 (N_147,In_627,In_1078);
or U148 (N_148,In_446,In_1122);
xnor U149 (N_149,In_973,In_1378);
and U150 (N_150,In_949,In_951);
and U151 (N_151,In_427,In_505);
nor U152 (N_152,In_770,In_292);
nor U153 (N_153,In_934,In_1359);
or U154 (N_154,In_1299,In_539);
nor U155 (N_155,In_1003,In_779);
and U156 (N_156,In_744,In_532);
and U157 (N_157,In_134,In_1174);
nand U158 (N_158,In_430,In_759);
nor U159 (N_159,In_941,In_1376);
or U160 (N_160,In_80,In_828);
xor U161 (N_161,In_1428,In_117);
xor U162 (N_162,In_1193,In_55);
nor U163 (N_163,In_525,In_498);
and U164 (N_164,In_1409,In_1032);
nand U165 (N_165,In_394,In_996);
nor U166 (N_166,In_1288,In_1364);
nand U167 (N_167,In_1382,In_658);
or U168 (N_168,In_1025,In_41);
or U169 (N_169,In_1236,In_573);
nor U170 (N_170,In_490,In_1239);
xnor U171 (N_171,In_868,In_85);
or U172 (N_172,In_215,In_313);
xnor U173 (N_173,In_120,In_1270);
nor U174 (N_174,In_1049,In_893);
or U175 (N_175,In_961,In_389);
xnor U176 (N_176,In_277,In_675);
xnor U177 (N_177,In_1194,In_1233);
or U178 (N_178,In_950,In_628);
nand U179 (N_179,In_1218,In_1490);
xor U180 (N_180,In_1439,In_291);
nor U181 (N_181,In_1062,In_1333);
nor U182 (N_182,In_763,In_263);
xor U183 (N_183,In_989,In_500);
or U184 (N_184,In_1302,In_884);
xnor U185 (N_185,In_520,In_1413);
or U186 (N_186,In_306,In_1320);
and U187 (N_187,In_1141,In_259);
and U188 (N_188,In_602,In_1045);
or U189 (N_189,In_1247,In_605);
or U190 (N_190,In_1094,In_71);
and U191 (N_191,In_683,In_501);
or U192 (N_192,In_283,In_665);
nor U193 (N_193,In_1038,In_1394);
or U194 (N_194,In_1487,In_718);
nand U195 (N_195,In_471,In_1391);
or U196 (N_196,In_1154,In_364);
nor U197 (N_197,In_59,In_687);
nor U198 (N_198,In_131,In_1245);
or U199 (N_199,In_767,In_1453);
xor U200 (N_200,In_107,In_639);
nand U201 (N_201,In_1047,In_56);
xor U202 (N_202,In_1395,N_41);
and U203 (N_203,In_789,In_694);
nor U204 (N_204,In_1118,In_1099);
and U205 (N_205,In_971,N_96);
and U206 (N_206,In_980,In_1457);
nand U207 (N_207,In_882,N_80);
and U208 (N_208,In_344,In_920);
xnor U209 (N_209,N_109,In_1124);
and U210 (N_210,In_890,N_112);
nand U211 (N_211,In_487,In_1323);
and U212 (N_212,In_523,In_1);
xnor U213 (N_213,In_62,In_746);
xor U214 (N_214,In_1210,In_219);
nor U215 (N_215,In_519,In_561);
nand U216 (N_216,In_496,In_1207);
and U217 (N_217,In_810,In_413);
and U218 (N_218,N_24,In_769);
or U219 (N_219,In_294,In_1372);
nand U220 (N_220,In_170,In_1348);
nor U221 (N_221,In_682,In_830);
and U222 (N_222,In_926,N_149);
nand U223 (N_223,In_84,In_1286);
and U224 (N_224,In_1172,In_589);
nand U225 (N_225,In_58,In_517);
nand U226 (N_226,In_302,In_368);
and U227 (N_227,In_1104,In_545);
nor U228 (N_228,N_33,In_876);
xnor U229 (N_229,In_1081,In_990);
nand U230 (N_230,In_1317,In_1324);
nor U231 (N_231,In_738,In_1046);
and U232 (N_232,N_114,In_726);
nand U233 (N_233,In_409,In_816);
nand U234 (N_234,In_37,In_23);
xor U235 (N_235,In_712,In_399);
nand U236 (N_236,In_210,N_105);
nand U237 (N_237,N_134,In_160);
nor U238 (N_238,In_171,In_53);
and U239 (N_239,In_1255,In_424);
nor U240 (N_240,In_1143,In_264);
and U241 (N_241,In_26,In_997);
and U242 (N_242,In_929,In_173);
or U243 (N_243,N_12,In_1219);
nor U244 (N_244,In_1173,N_99);
or U245 (N_245,N_32,In_715);
xor U246 (N_246,In_698,In_640);
nand U247 (N_247,In_275,In_1351);
nand U248 (N_248,N_167,In_253);
or U249 (N_249,In_1363,In_457);
xor U250 (N_250,In_891,N_72);
or U251 (N_251,In_841,In_1232);
xor U252 (N_252,In_829,In_720);
xor U253 (N_253,In_293,In_764);
xor U254 (N_254,In_418,In_922);
nand U255 (N_255,N_146,N_39);
and U256 (N_256,In_1459,In_1423);
nor U257 (N_257,In_988,N_63);
nand U258 (N_258,In_878,In_753);
xor U259 (N_259,In_1203,In_8);
xor U260 (N_260,In_667,In_825);
xor U261 (N_261,N_44,In_97);
xnor U262 (N_262,N_76,N_43);
xnor U263 (N_263,N_61,In_422);
and U264 (N_264,In_18,N_158);
nor U265 (N_265,In_761,In_1448);
nor U266 (N_266,In_1150,N_126);
or U267 (N_267,In_508,In_146);
and U268 (N_268,In_269,In_1343);
and U269 (N_269,In_1392,In_809);
or U270 (N_270,In_315,In_1399);
nand U271 (N_271,In_48,In_417);
xor U272 (N_272,In_460,N_170);
nor U273 (N_273,N_68,In_579);
and U274 (N_274,In_1251,In_580);
or U275 (N_275,In_1202,N_162);
nor U276 (N_276,N_133,In_333);
and U277 (N_277,In_587,In_771);
or U278 (N_278,In_1188,N_123);
nor U279 (N_279,In_1134,In_7);
and U280 (N_280,In_630,In_1311);
and U281 (N_281,In_301,In_1105);
xnor U282 (N_282,In_535,In_1214);
xnor U283 (N_283,In_222,In_558);
nand U284 (N_284,In_406,In_1266);
nor U285 (N_285,N_42,N_66);
xor U286 (N_286,In_499,In_289);
nor U287 (N_287,In_30,N_48);
and U288 (N_288,In_736,In_953);
or U289 (N_289,In_947,In_382);
xor U290 (N_290,In_625,In_987);
or U291 (N_291,In_958,In_99);
nand U292 (N_292,In_1300,In_415);
nor U293 (N_293,In_162,In_727);
nand U294 (N_294,N_31,In_285);
and U295 (N_295,In_1405,In_1496);
nand U296 (N_296,In_1075,In_657);
xor U297 (N_297,In_994,N_94);
nand U298 (N_298,In_1278,In_1208);
and U299 (N_299,In_1268,In_1036);
nor U300 (N_300,In_1340,In_1312);
or U301 (N_301,In_113,In_729);
or U302 (N_302,In_1135,In_1216);
xnor U303 (N_303,In_728,In_75);
nor U304 (N_304,In_1223,In_149);
and U305 (N_305,In_647,In_960);
nor U306 (N_306,In_1000,In_633);
xnor U307 (N_307,In_1318,In_1147);
xor U308 (N_308,N_184,In_618);
or U309 (N_309,In_392,In_611);
and U310 (N_310,In_970,N_161);
and U311 (N_311,In_984,In_1144);
nor U312 (N_312,In_904,In_1020);
xor U313 (N_313,N_129,In_1386);
xnor U314 (N_314,In_385,In_896);
nor U315 (N_315,In_1263,N_67);
nor U316 (N_316,In_1240,In_731);
nor U317 (N_317,In_1262,In_72);
or U318 (N_318,In_1485,In_557);
xor U319 (N_319,In_600,N_69);
xnor U320 (N_320,In_158,In_309);
xnor U321 (N_321,In_130,In_1465);
nor U322 (N_322,In_1441,In_638);
xnor U323 (N_323,In_1258,In_1478);
xnor U324 (N_324,In_323,In_662);
or U325 (N_325,In_340,In_915);
and U326 (N_326,In_77,In_255);
or U327 (N_327,In_1074,N_21);
and U328 (N_328,In_786,In_540);
xor U329 (N_329,N_108,In_483);
or U330 (N_330,In_1269,N_92);
xor U331 (N_331,In_447,In_121);
and U332 (N_332,In_883,In_1087);
nand U333 (N_333,N_19,N_166);
or U334 (N_334,In_100,In_1005);
xnor U335 (N_335,In_653,In_353);
and U336 (N_336,In_801,In_1480);
xnor U337 (N_337,N_119,In_943);
nand U338 (N_338,In_711,In_1002);
nor U339 (N_339,In_198,In_637);
nand U340 (N_340,In_108,In_398);
nor U341 (N_341,In_684,In_1484);
nand U342 (N_342,In_710,In_805);
nand U343 (N_343,In_995,N_124);
xor U344 (N_344,In_879,In_745);
xnor U345 (N_345,In_1462,In_156);
and U346 (N_346,In_1298,In_1127);
or U347 (N_347,In_673,In_515);
xnor U348 (N_348,N_196,In_1101);
nor U349 (N_349,In_396,In_707);
and U350 (N_350,In_1016,In_565);
and U351 (N_351,In_1289,N_51);
nor U352 (N_352,In_814,In_1161);
nand U353 (N_353,N_83,In_473);
and U354 (N_354,In_656,In_1293);
xor U355 (N_355,N_11,In_260);
xnor U356 (N_356,In_504,In_109);
or U357 (N_357,In_524,In_529);
and U358 (N_358,In_300,In_132);
nor U359 (N_359,In_1282,In_429);
nand U360 (N_360,In_854,In_1095);
and U361 (N_361,In_695,In_593);
nand U362 (N_362,N_187,In_308);
xnor U363 (N_363,In_1415,In_11);
xnor U364 (N_364,In_383,In_740);
nor U365 (N_365,In_1160,In_438);
or U366 (N_366,In_1301,In_1069);
nand U367 (N_367,N_171,In_864);
xnor U368 (N_368,In_15,In_838);
and U369 (N_369,In_373,In_419);
xnor U370 (N_370,In_303,In_456);
or U371 (N_371,In_282,In_900);
nand U372 (N_372,N_137,N_38);
nor U373 (N_373,In_115,In_1316);
and U374 (N_374,In_195,In_972);
or U375 (N_375,In_231,In_346);
xnor U376 (N_376,In_550,In_240);
xnor U377 (N_377,In_236,In_1211);
nor U378 (N_378,In_22,In_511);
xnor U379 (N_379,In_1313,In_703);
nand U380 (N_380,In_992,In_671);
nand U381 (N_381,In_965,In_1136);
nand U382 (N_382,In_1043,In_408);
nand U383 (N_383,In_599,In_1084);
or U384 (N_384,N_174,In_948);
or U385 (N_385,In_213,In_966);
xnor U386 (N_386,In_261,In_513);
xor U387 (N_387,N_40,In_227);
xnor U388 (N_388,In_362,N_157);
and U389 (N_389,In_1291,In_455);
and U390 (N_390,In_708,In_881);
nand U391 (N_391,In_1421,In_1060);
xnor U392 (N_392,In_356,In_624);
or U393 (N_393,In_843,In_357);
and U394 (N_394,In_491,N_29);
and U395 (N_395,In_1442,In_842);
nand U396 (N_396,In_280,N_136);
or U397 (N_397,In_350,N_53);
or U398 (N_398,In_360,In_1495);
xnor U399 (N_399,In_942,N_60);
nor U400 (N_400,In_1429,In_526);
nand U401 (N_401,In_886,In_397);
nor U402 (N_402,In_632,N_323);
xnor U403 (N_403,N_389,N_73);
nor U404 (N_404,In_1474,In_441);
xor U405 (N_405,In_614,In_1418);
or U406 (N_406,In_867,N_177);
nand U407 (N_407,In_297,In_1072);
nor U408 (N_408,In_70,N_181);
and U409 (N_409,In_386,In_1158);
xor U410 (N_410,In_774,N_262);
xor U411 (N_411,In_781,In_1170);
nand U412 (N_412,In_1241,N_282);
xor U413 (N_413,N_128,N_365);
xor U414 (N_414,N_204,N_203);
nor U415 (N_415,In_244,N_13);
and U416 (N_416,In_612,In_128);
or U417 (N_417,N_106,In_1337);
xnor U418 (N_418,In_150,N_366);
nor U419 (N_419,N_292,In_521);
xor U420 (N_420,In_866,In_669);
or U421 (N_421,In_1116,In_390);
xnor U422 (N_422,In_899,In_713);
and U423 (N_423,N_224,In_1092);
xnor U424 (N_424,N_289,In_243);
nand U425 (N_425,In_1129,N_144);
nand U426 (N_426,N_229,In_19);
or U427 (N_427,In_914,N_261);
nand U428 (N_428,In_1227,In_1486);
nor U429 (N_429,In_1133,N_291);
and U430 (N_430,In_462,N_393);
and U431 (N_431,In_510,In_850);
or U432 (N_432,In_319,N_168);
nand U433 (N_433,N_14,N_26);
xor U434 (N_434,In_1326,N_185);
nand U435 (N_435,In_322,N_78);
nor U436 (N_436,In_461,In_1249);
or U437 (N_437,In_1354,In_1014);
nand U438 (N_438,N_192,In_336);
and U439 (N_439,In_811,In_1179);
nor U440 (N_440,N_260,In_1403);
or U441 (N_441,In_1066,N_209);
or U442 (N_442,N_254,N_5);
nand U443 (N_443,N_86,In_768);
xnor U444 (N_444,In_1204,In_32);
and U445 (N_445,In_1366,In_347);
xor U446 (N_446,In_813,In_1435);
nand U447 (N_447,In_636,N_71);
nor U448 (N_448,In_681,In_1353);
or U449 (N_449,In_777,N_182);
nand U450 (N_450,N_276,In_723);
and U451 (N_451,N_234,N_142);
and U452 (N_452,N_20,In_138);
or U453 (N_453,In_897,N_300);
xnor U454 (N_454,N_110,N_315);
xnor U455 (N_455,In_262,N_55);
or U456 (N_456,In_1234,In_1398);
and U457 (N_457,N_238,In_981);
nand U458 (N_458,In_564,In_1110);
nor U459 (N_459,N_207,In_148);
xnor U460 (N_460,In_328,N_214);
nand U461 (N_461,N_147,N_74);
nor U462 (N_462,In_87,N_259);
and U463 (N_463,N_369,N_28);
nor U464 (N_464,N_297,In_1296);
or U465 (N_465,In_819,In_144);
and U466 (N_466,In_326,N_225);
and U467 (N_467,N_165,N_372);
nor U468 (N_468,N_235,In_772);
xnor U469 (N_469,In_741,In_1213);
or U470 (N_470,In_475,N_285);
or U471 (N_471,N_352,N_397);
xor U472 (N_472,N_373,N_347);
or U473 (N_473,In_224,In_50);
nand U474 (N_474,N_304,In_324);
and U475 (N_475,N_183,In_110);
and U476 (N_476,N_223,In_288);
and U477 (N_477,N_339,In_1265);
nor U478 (N_478,In_1217,In_478);
or U479 (N_479,N_267,N_160);
or U480 (N_480,N_172,In_871);
and U481 (N_481,N_59,In_651);
xor U482 (N_482,In_575,N_163);
and U483 (N_483,In_925,In_1284);
or U484 (N_484,N_311,In_366);
nand U485 (N_485,In_844,In_1021);
xor U486 (N_486,N_202,In_860);
nor U487 (N_487,In_1369,In_861);
and U488 (N_488,In_420,In_355);
and U489 (N_489,N_322,In_1182);
xor U490 (N_490,In_352,In_1368);
or U491 (N_491,In_428,In_217);
xor U492 (N_492,In_1246,In_836);
xnor U493 (N_493,N_251,N_386);
nand U494 (N_494,N_272,In_81);
or U495 (N_495,In_752,In_1385);
nand U496 (N_496,In_82,N_97);
nor U497 (N_497,In_1449,N_194);
nand U498 (N_498,In_659,In_1029);
or U499 (N_499,In_304,N_127);
and U500 (N_500,N_221,In_434);
or U501 (N_501,N_394,In_1142);
or U502 (N_502,N_257,In_233);
or U503 (N_503,In_25,In_595);
xor U504 (N_504,In_1017,In_238);
nor U505 (N_505,N_310,N_248);
xnor U506 (N_506,In_617,In_824);
nand U507 (N_507,In_257,In_1162);
nor U508 (N_508,In_652,In_31);
xnor U509 (N_509,In_1187,In_1389);
nand U510 (N_510,N_327,In_278);
or U511 (N_511,In_34,N_1);
nand U512 (N_512,N_353,N_191);
xnor U513 (N_513,N_175,In_161);
nor U514 (N_514,N_93,In_13);
and U515 (N_515,N_379,In_1097);
xnor U516 (N_516,In_1349,N_263);
nor U517 (N_517,In_377,N_22);
or U518 (N_518,In_578,In_151);
nand U519 (N_519,N_271,N_299);
or U520 (N_520,In_716,N_9);
or U521 (N_521,In_167,In_645);
nor U522 (N_522,In_1053,In_1175);
or U523 (N_523,N_15,In_1065);
and U524 (N_524,N_312,In_472);
and U525 (N_525,N_46,In_562);
xor U526 (N_526,In_33,In_700);
nand U527 (N_527,In_163,N_141);
and U528 (N_528,In_192,In_803);
nand U529 (N_529,In_90,In_827);
and U530 (N_530,N_309,In_402);
xor U531 (N_531,In_812,N_87);
or U532 (N_532,In_86,In_126);
or U533 (N_533,In_822,In_207);
or U534 (N_534,In_512,N_16);
xor U535 (N_535,In_1151,In_661);
xor U536 (N_536,In_800,In_1098);
or U537 (N_537,In_1252,In_1163);
nor U538 (N_538,In_1183,In_766);
xnor U539 (N_539,N_91,In_178);
or U540 (N_540,In_1067,N_36);
or U541 (N_541,In_376,In_1425);
nand U542 (N_542,N_363,In_52);
xor U543 (N_543,In_930,N_336);
nor U544 (N_544,In_1015,N_189);
nor U545 (N_545,In_1126,In_1189);
nand U546 (N_546,In_305,N_2);
or U547 (N_547,N_375,N_398);
and U548 (N_548,In_643,In_985);
nand U549 (N_549,In_9,In_670);
nand U550 (N_550,In_405,In_1380);
xor U551 (N_551,In_106,In_1050);
and U552 (N_552,N_200,In_648);
nor U553 (N_553,N_302,N_199);
xnor U554 (N_554,In_135,In_911);
nand U555 (N_555,In_1011,In_509);
and U556 (N_556,In_788,In_363);
or U557 (N_557,In_674,N_385);
xor U558 (N_558,In_757,In_464);
nor U559 (N_559,N_269,N_340);
nor U560 (N_560,N_252,N_329);
or U561 (N_561,In_1477,In_1275);
or U562 (N_562,In_1264,In_534);
or U563 (N_563,In_1467,In_613);
nor U564 (N_564,In_42,In_1454);
or U565 (N_565,N_103,In_685);
nor U566 (N_566,In_365,In_835);
xor U567 (N_567,In_452,In_1406);
nand U568 (N_568,In_699,In_348);
or U569 (N_569,N_159,In_172);
xor U570 (N_570,In_1292,In_902);
nand U571 (N_571,In_299,In_1082);
and U572 (N_572,In_1080,In_1220);
and U573 (N_573,In_913,In_401);
xnor U574 (N_574,In_626,N_3);
xor U575 (N_575,In_1237,In_153);
xnor U576 (N_576,N_65,In_792);
and U577 (N_577,In_51,In_1109);
and U578 (N_578,N_213,In_489);
and U579 (N_579,In_907,N_102);
or U580 (N_580,In_649,In_433);
nor U581 (N_581,In_834,In_894);
xor U582 (N_582,N_132,In_494);
nand U583 (N_583,In_1308,In_1276);
or U584 (N_584,In_1341,N_290);
nor U585 (N_585,N_356,In_1498);
xor U586 (N_586,In_979,N_348);
and U587 (N_587,In_1492,N_151);
or U588 (N_588,N_391,N_239);
nor U589 (N_589,N_280,In_1093);
nor U590 (N_590,In_388,In_14);
nand U591 (N_591,In_63,In_1048);
nor U592 (N_592,In_103,In_888);
nor U593 (N_593,N_342,In_762);
or U594 (N_594,In_1212,In_680);
and U595 (N_595,In_1419,In_1004);
nand U596 (N_596,In_1452,N_81);
and U597 (N_597,N_115,In_901);
nand U598 (N_598,In_732,In_1279);
nand U599 (N_599,In_704,N_173);
nand U600 (N_600,In_853,N_409);
and U601 (N_601,N_429,N_337);
xnor U602 (N_602,In_849,N_432);
xnor U603 (N_603,N_537,N_79);
xnor U604 (N_604,N_104,In_831);
or U605 (N_605,In_1051,In_616);
xnor U606 (N_606,In_875,In_982);
xor U607 (N_607,N_428,In_1433);
and U608 (N_608,In_1307,N_510);
or U609 (N_609,In_541,In_773);
nor U610 (N_610,N_57,In_1401);
nor U611 (N_611,In_425,In_426);
and U612 (N_612,N_459,In_374);
or U613 (N_613,N_460,In_1383);
nand U614 (N_614,In_604,N_335);
and U615 (N_615,N_232,In_585);
or U616 (N_616,N_569,N_378);
xnor U617 (N_617,N_334,In_821);
nor U618 (N_618,In_1196,N_499);
or U619 (N_619,In_174,N_509);
nor U620 (N_620,N_574,N_488);
and U621 (N_621,In_1414,N_581);
and U622 (N_622,In_1277,In_17);
nand U623 (N_623,In_1444,In_321);
or U624 (N_624,In_124,In_569);
and U625 (N_625,N_454,In_1121);
nor U626 (N_626,In_1006,In_1273);
xnor U627 (N_627,In_765,In_307);
xor U628 (N_628,N_294,N_82);
and U629 (N_629,In_1253,In_1076);
and U630 (N_630,In_635,N_421);
and U631 (N_631,In_459,In_367);
and U632 (N_632,In_1330,In_1197);
or U633 (N_633,N_449,N_8);
nor U634 (N_634,N_402,N_361);
nand U635 (N_635,N_169,In_1171);
or U636 (N_636,N_359,In_448);
xor U637 (N_637,N_273,In_1280);
nor U638 (N_638,In_252,In_1039);
and U639 (N_639,N_417,N_475);
nand U640 (N_640,In_1281,N_591);
xnor U641 (N_641,N_461,In_272);
nor U642 (N_642,In_592,N_407);
or U643 (N_643,N_433,In_1086);
and U644 (N_644,In_338,In_102);
nor U645 (N_645,N_399,In_530);
and U646 (N_646,N_583,N_512);
nor U647 (N_647,N_388,In_177);
nor U648 (N_648,In_666,In_1322);
nor U649 (N_649,N_500,In_536);
nor U650 (N_650,In_1430,In_802);
nor U651 (N_651,N_278,In_436);
xnor U652 (N_652,In_474,N_561);
and U653 (N_653,In_4,N_331);
nand U654 (N_654,In_235,N_562);
nand U655 (N_655,N_592,In_64);
or U656 (N_656,N_457,In_778);
xor U657 (N_657,N_400,N_298);
xnor U658 (N_658,In_1089,In_486);
or U659 (N_659,In_754,In_354);
nand U660 (N_660,In_105,In_76);
xnor U661 (N_661,N_90,In_840);
xnor U662 (N_662,In_1393,In_1085);
or U663 (N_663,N_571,N_484);
nor U664 (N_664,In_20,In_78);
and U665 (N_665,In_114,N_117);
nand U666 (N_666,In_1328,In_1365);
nor U667 (N_667,In_372,N_406);
xor U668 (N_668,N_513,In_481);
xnor U669 (N_669,In_1242,In_654);
nor U670 (N_670,In_1443,In_1198);
or U671 (N_671,N_525,N_101);
nor U672 (N_672,In_189,In_567);
and U673 (N_673,In_581,In_1387);
or U674 (N_674,In_1091,In_755);
nand U675 (N_675,In_349,In_1356);
xor U676 (N_676,N_326,N_296);
xnor U677 (N_677,N_477,In_939);
xnor U678 (N_678,N_351,In_497);
and U679 (N_679,N_469,N_476);
xnor U680 (N_680,In_924,N_18);
xnor U681 (N_681,N_383,In_1440);
nand U682 (N_682,N_597,N_565);
nand U683 (N_683,N_424,In_1431);
nand U684 (N_684,N_303,N_266);
xnor U685 (N_685,N_503,In_247);
nor U686 (N_686,In_1360,In_1303);
nand U687 (N_687,In_1469,N_211);
xnor U688 (N_688,N_295,N_566);
nor U689 (N_689,In_1491,N_116);
and U690 (N_690,N_522,N_528);
xnor U691 (N_691,In_49,In_1120);
and U692 (N_692,In_476,In_1128);
nand U693 (N_693,In_92,N_230);
nor U694 (N_694,N_594,In_544);
and U695 (N_695,In_537,In_641);
and U696 (N_696,In_620,N_478);
and U697 (N_697,N_56,In_688);
and U698 (N_698,N_466,N_568);
or U699 (N_699,In_634,In_678);
and U700 (N_700,In_952,N_198);
or U701 (N_701,In_466,N_504);
nor U702 (N_702,In_180,In_83);
and U703 (N_703,In_1244,In_1206);
or U704 (N_704,N_416,N_575);
or U705 (N_705,In_310,In_1221);
xnor U706 (N_706,In_1058,N_468);
or U707 (N_707,N_554,In_145);
xor U708 (N_708,N_62,In_576);
xnor U709 (N_709,N_555,In_330);
or U710 (N_710,In_933,N_392);
nor U711 (N_711,In_1181,N_438);
xnor U712 (N_712,In_1436,N_544);
xnor U713 (N_713,In_998,N_593);
or U714 (N_714,In_341,In_248);
xor U715 (N_715,N_10,N_535);
or U716 (N_716,N_236,N_412);
or U717 (N_717,N_228,In_1294);
xor U718 (N_718,N_529,In_1132);
nor U719 (N_719,N_307,N_405);
or U720 (N_720,N_27,In_40);
nand U721 (N_721,In_748,In_414);
and U722 (N_722,In_325,In_848);
xor U723 (N_723,N_547,N_135);
and U724 (N_724,N_49,In_68);
or U725 (N_725,N_573,In_548);
and U726 (N_726,N_448,In_140);
nor U727 (N_727,In_1235,In_791);
and U728 (N_728,In_719,N_464);
or U729 (N_729,N_390,N_494);
nand U730 (N_730,In_239,In_725);
xor U731 (N_731,In_251,N_502);
nor U732 (N_732,In_1357,In_969);
nor U733 (N_733,N_107,In_586);
nor U734 (N_734,In_225,N_131);
or U735 (N_735,In_1335,In_181);
xnor U736 (N_736,In_968,In_815);
and U737 (N_737,N_180,In_101);
xnor U738 (N_738,N_47,In_1402);
xnor U739 (N_739,N_330,In_1473);
xor U740 (N_740,In_978,In_442);
nand U741 (N_741,In_1332,In_1139);
xnor U742 (N_742,N_495,N_576);
and U743 (N_743,N_368,In_568);
nor U744 (N_744,N_64,N_420);
nand U745 (N_745,N_441,N_121);
or U746 (N_746,In_880,In_783);
nor U747 (N_747,In_226,In_857);
xnor U748 (N_748,N_306,N_358);
or U749 (N_749,N_283,In_1437);
xor U750 (N_750,N_215,In_927);
or U751 (N_751,In_187,N_384);
nand U752 (N_752,In_250,N_270);
xnor U753 (N_753,In_677,In_10);
or U754 (N_754,In_1073,N_538);
and U755 (N_755,In_137,In_404);
nand U756 (N_756,In_1031,In_281);
nor U757 (N_757,In_845,In_125);
xnor U758 (N_758,In_1411,In_910);
and U759 (N_759,In_1438,N_563);
or U760 (N_760,In_24,In_393);
or U761 (N_761,N_524,In_1304);
xor U762 (N_762,In_603,N_195);
xnor U763 (N_763,In_492,In_621);
nand U764 (N_764,In_1145,N_589);
and U765 (N_765,N_564,In_1325);
or U766 (N_766,In_1471,In_722);
and U767 (N_767,In_164,N_212);
or U768 (N_768,In_582,N_100);
nor U769 (N_769,In_1140,In_379);
and U770 (N_770,In_1420,N_531);
xnor U771 (N_771,In_1260,In_359);
or U772 (N_772,N_250,N_410);
xor U773 (N_773,N_34,N_458);
xnor U774 (N_774,In_506,N_288);
and U775 (N_775,N_186,In_820);
and U776 (N_776,In_287,N_152);
and U777 (N_777,N_534,N_344);
nand U778 (N_778,In_67,In_54);
nor U779 (N_779,In_1283,N_244);
nor U780 (N_780,In_3,In_794);
xnor U781 (N_781,N_491,In_407);
and U782 (N_782,N_139,In_387);
or U783 (N_783,In_94,N_140);
or U784 (N_784,In_804,N_560);
nand U785 (N_785,N_552,In_1370);
or U786 (N_786,In_298,In_311);
xor U787 (N_787,In_1397,In_358);
nor U788 (N_788,N_243,In_1229);
xnor U789 (N_789,In_241,N_546);
and U790 (N_790,In_66,N_287);
and U791 (N_791,N_258,In_454);
xnor U792 (N_792,In_186,N_328);
xor U793 (N_793,N_401,N_367);
nor U794 (N_794,In_61,In_717);
nor U795 (N_795,In_290,N_413);
and U796 (N_796,N_508,In_482);
xnor U797 (N_797,N_493,N_305);
nor U798 (N_798,N_532,N_588);
or U799 (N_799,N_450,N_440);
or U800 (N_800,N_559,In_266);
nand U801 (N_801,In_320,N_764);
or U802 (N_802,N_617,N_422);
or U803 (N_803,N_427,N_320);
nor U804 (N_804,N_624,In_435);
nand U805 (N_805,N_598,N_542);
xnor U806 (N_806,N_426,N_242);
xnor U807 (N_807,N_775,In_629);
nand U808 (N_808,N_643,N_75);
xnor U809 (N_809,In_265,In_1310);
or U810 (N_810,In_1346,N_687);
nor U811 (N_811,In_676,In_218);
xnor U812 (N_812,In_839,In_276);
and U813 (N_813,N_719,N_463);
nor U814 (N_814,N_619,N_790);
or U815 (N_815,N_275,In_1243);
and U816 (N_816,In_1417,N_490);
or U817 (N_817,In_921,In_935);
and U818 (N_818,N_455,In_1344);
nor U819 (N_819,N_241,N_343);
and U820 (N_820,N_692,N_319);
or U821 (N_821,In_1035,N_553);
or U822 (N_822,N_150,N_467);
and U823 (N_823,In_274,N_54);
nor U824 (N_824,In_484,N_725);
xor U825 (N_825,In_538,In_514);
xor U826 (N_826,N_148,N_694);
or U827 (N_827,In_986,In_1228);
xnor U828 (N_828,N_474,In_1149);
or U829 (N_829,N_52,N_506);
nand U830 (N_830,N_370,N_138);
or U831 (N_831,In_689,N_541);
or U832 (N_832,N_498,N_627);
or U833 (N_833,In_43,In_27);
or U834 (N_834,N_596,N_540);
and U835 (N_835,N_473,In_714);
or U836 (N_836,N_155,N_762);
xnor U837 (N_837,N_345,In_190);
nor U838 (N_838,In_74,In_5);
or U839 (N_839,N_445,N_631);
nand U840 (N_840,In_1185,N_621);
nor U841 (N_841,In_378,In_122);
and U842 (N_842,N_277,N_655);
or U843 (N_843,In_1222,In_742);
or U844 (N_844,N_425,N_645);
and U845 (N_845,N_550,N_746);
nor U846 (N_846,N_84,N_620);
nor U847 (N_847,In_1028,N_113);
nor U848 (N_848,N_201,N_190);
or U849 (N_849,N_497,N_613);
or U850 (N_850,N_684,N_713);
and U851 (N_851,N_750,N_556);
nor U852 (N_852,In_1250,N_797);
nor U853 (N_853,In_957,N_768);
and U854 (N_854,N_614,N_111);
nor U855 (N_855,N_471,N_118);
nand U856 (N_856,N_122,N_453);
and U857 (N_857,N_639,In_1384);
or U858 (N_858,N_220,N_206);
nor U859 (N_859,N_233,N_663);
or U860 (N_860,N_362,In_375);
xnor U861 (N_861,N_761,In_1180);
xor U862 (N_862,In_693,In_1493);
xor U863 (N_863,In_623,N_634);
and U864 (N_864,N_660,In_1225);
nand U865 (N_865,N_264,N_25);
xnor U866 (N_866,In_1447,N_268);
nand U867 (N_867,In_1224,In_467);
and U868 (N_868,N_88,N_346);
and U869 (N_869,In_46,In_123);
nor U870 (N_870,N_794,In_1455);
nand U871 (N_871,N_696,N_654);
nand U872 (N_872,N_324,In_956);
or U873 (N_873,N_515,In_185);
nor U874 (N_874,In_391,N_465);
nor U875 (N_875,N_772,In_877);
xnor U876 (N_876,In_1131,N_325);
nand U877 (N_877,N_740,N_770);
and U878 (N_878,N_675,In_983);
or U879 (N_879,N_710,N_676);
and U880 (N_880,N_249,In_1034);
and U881 (N_881,N_293,N_403);
nand U882 (N_882,In_194,In_183);
xor U883 (N_883,N_247,In_622);
nor U884 (N_884,N_431,N_567);
and U885 (N_885,In_808,In_549);
or U886 (N_886,In_780,In_750);
nor U887 (N_887,In_119,In_16);
nor U888 (N_888,N_418,In_1090);
nor U889 (N_889,In_111,In_1168);
and U890 (N_890,N_349,In_1482);
nand U891 (N_891,N_193,In_176);
or U892 (N_892,In_1119,N_482);
nand U893 (N_893,In_784,In_1018);
nand U894 (N_894,N_30,N_527);
xnor U895 (N_895,N_89,In_502);
xnor U896 (N_896,N_179,In_166);
or U897 (N_897,N_154,N_360);
or U898 (N_898,N_788,N_557);
nor U899 (N_899,N_253,In_847);
nand U900 (N_900,N_626,N_789);
or U901 (N_901,N_314,In_312);
nand U902 (N_902,N_164,N_666);
and U903 (N_903,In_570,In_690);
xnor U904 (N_904,N_782,N_671);
nor U905 (N_905,N_237,In_1010);
nand U906 (N_906,N_579,N_197);
nor U907 (N_907,N_609,N_443);
nor U908 (N_908,N_649,N_6);
and U909 (N_909,N_670,N_724);
or U910 (N_910,N_387,In_228);
or U911 (N_911,N_721,In_823);
and U912 (N_912,N_667,N_691);
or U913 (N_913,N_767,In_1321);
or U914 (N_914,N_751,In_1077);
nor U915 (N_915,N_795,N_735);
or U916 (N_916,N_545,N_357);
or U917 (N_917,N_364,N_395);
xor U918 (N_918,In_1458,N_774);
xnor U919 (N_919,In_1461,N_702);
or U920 (N_920,N_599,In_940);
or U921 (N_921,N_616,In_493);
xor U922 (N_922,N_487,In_584);
nand U923 (N_923,In_1008,In_799);
xor U924 (N_924,In_782,In_724);
and U925 (N_925,In_1481,In_898);
nand U926 (N_926,N_58,In_1336);
and U927 (N_927,N_727,In_314);
nand U928 (N_928,N_377,N_771);
nand U929 (N_929,N_658,In_1361);
nand U930 (N_930,N_451,N_143);
and U931 (N_931,N_281,N_729);
xnor U932 (N_932,In_1231,N_622);
nor U933 (N_933,N_125,N_0);
or U934 (N_934,N_683,In_533);
nand U935 (N_935,N_798,In_188);
xor U936 (N_936,In_175,In_597);
and U937 (N_937,N_217,N_321);
nor U938 (N_938,N_50,In_147);
nand U939 (N_939,N_668,N_483);
xnor U940 (N_940,In_642,N_444);
xor U941 (N_941,In_1488,In_885);
and U942 (N_942,In_1148,N_793);
and U943 (N_943,N_739,N_640);
nor U944 (N_944,In_495,N_706);
xor U945 (N_945,N_700,N_578);
nor U946 (N_946,In_1164,In_655);
nor U947 (N_947,In_1041,N_437);
nand U948 (N_948,N_648,N_759);
and U949 (N_949,N_618,N_4);
nor U950 (N_950,N_633,In_196);
and U951 (N_951,N_404,N_712);
nand U952 (N_952,N_610,N_690);
or U953 (N_953,N_741,N_265);
and U954 (N_954,In_660,In_1063);
xnor U955 (N_955,In_1042,N_763);
and U956 (N_956,N_787,In_214);
nor U957 (N_957,N_430,N_396);
xor U958 (N_958,N_623,N_611);
nand U959 (N_959,In_1412,N_585);
or U960 (N_960,In_596,N_605);
or U961 (N_961,In_522,In_1199);
and U962 (N_962,N_717,In_1375);
nand U963 (N_963,In_112,In_1271);
and U964 (N_964,In_709,N_681);
xor U965 (N_965,In_787,N_786);
nor U966 (N_966,In_1381,In_361);
nand U967 (N_967,N_210,In_345);
xor U968 (N_968,N_776,N_374);
and U969 (N_969,In_837,In_1256);
and U970 (N_970,In_743,N_641);
and U971 (N_971,In_999,N_756);
xor U972 (N_972,N_35,In_598);
or U973 (N_973,N_586,In_488);
nor U974 (N_974,In_1156,In_439);
nor U975 (N_975,In_165,N_766);
or U976 (N_976,In_975,In_1422);
xnor U977 (N_977,In_38,N_682);
and U978 (N_978,In_477,N_85);
nor U979 (N_979,N_604,N_501);
nand U980 (N_980,In_1040,In_692);
nand U981 (N_981,N_246,N_673);
xnor U982 (N_982,N_37,In_962);
xnor U983 (N_983,N_745,N_720);
or U984 (N_984,N_587,N_695);
nand U985 (N_985,N_240,In_191);
and U986 (N_986,N_791,In_1315);
or U987 (N_987,N_301,N_549);
nor U988 (N_988,N_218,N_595);
xnor U989 (N_989,In_443,N_635);
or U990 (N_990,In_1027,N_350);
nor U991 (N_991,N_145,N_630);
and U992 (N_992,In_1125,N_354);
or U993 (N_993,In_1479,In_411);
nor U994 (N_994,In_229,In_610);
nor U995 (N_995,In_552,N_274);
and U996 (N_996,N_737,N_130);
nor U997 (N_997,In_870,In_157);
and U998 (N_998,In_65,N_615);
nor U999 (N_999,N_376,In_421);
nand U1000 (N_1000,N_156,N_874);
or U1001 (N_1001,N_582,N_742);
nand U1002 (N_1002,N_636,N_932);
nor U1003 (N_1003,N_452,N_840);
nor U1004 (N_1004,N_859,N_827);
nand U1005 (N_1005,N_881,N_644);
nand U1006 (N_1006,N_653,N_792);
and U1007 (N_1007,In_403,N_950);
and U1008 (N_1008,In_143,N_646);
nand U1009 (N_1009,N_434,N_678);
xnor U1010 (N_1010,N_955,N_948);
or U1011 (N_1011,In_869,N_908);
and U1012 (N_1012,N_849,N_867);
nand U1013 (N_1013,N_338,N_659);
and U1014 (N_1014,In_268,N_965);
xor U1015 (N_1015,N_558,In_254);
and U1016 (N_1016,In_1230,N_805);
xor U1017 (N_1017,N_205,N_414);
and U1018 (N_1018,N_98,N_960);
xnor U1019 (N_1019,In_1446,N_925);
xor U1020 (N_1020,N_927,In_1001);
nor U1021 (N_1021,N_308,N_732);
and U1022 (N_1022,In_588,In_133);
nand U1023 (N_1023,In_874,N_479);
xor U1024 (N_1024,N_255,N_958);
and U1025 (N_1025,N_333,N_901);
or U1026 (N_1026,In_1026,In_201);
and U1027 (N_1027,N_523,N_677);
xor U1028 (N_1028,In_663,N_912);
and U1029 (N_1029,N_880,In_1483);
nor U1030 (N_1030,N_590,N_456);
nand U1031 (N_1031,In_1071,N_834);
nand U1032 (N_1032,In_954,In_1023);
or U1033 (N_1033,In_69,N_817);
xor U1034 (N_1034,In_168,N_996);
nor U1035 (N_1035,N_521,N_208);
and U1036 (N_1036,N_778,N_853);
and U1037 (N_1037,N_946,In_197);
nand U1038 (N_1038,N_885,In_209);
or U1039 (N_1039,N_911,N_884);
and U1040 (N_1040,N_906,In_468);
or U1041 (N_1041,N_647,N_808);
xor U1042 (N_1042,N_577,In_963);
xnor U1043 (N_1043,N_758,N_813);
nand U1044 (N_1044,N_802,In_944);
xor U1045 (N_1045,N_227,N_652);
and U1046 (N_1046,N_882,N_699);
xor U1047 (N_1047,In_216,N_415);
xor U1048 (N_1048,N_889,N_752);
nand U1049 (N_1049,In_1267,N_847);
or U1050 (N_1050,N_707,N_178);
nor U1051 (N_1051,N_219,N_730);
or U1052 (N_1052,N_883,In_89);
and U1053 (N_1053,N_686,N_820);
xnor U1054 (N_1054,N_969,N_472);
and U1055 (N_1055,N_905,In_916);
xnor U1056 (N_1056,N_868,N_811);
nor U1057 (N_1057,N_704,N_600);
nor U1058 (N_1058,N_45,N_753);
or U1059 (N_1059,N_994,N_919);
and U1060 (N_1060,N_841,N_176);
xor U1061 (N_1061,In_334,N_381);
or U1062 (N_1062,N_843,In_371);
xnor U1063 (N_1063,In_590,N_899);
or U1064 (N_1064,N_470,N_679);
xor U1065 (N_1065,In_1272,N_818);
xor U1066 (N_1066,N_507,N_726);
xnor U1067 (N_1067,N_992,N_602);
nor U1068 (N_1068,N_738,In_242);
xnor U1069 (N_1069,In_1146,N_530);
xor U1070 (N_1070,In_507,In_1107);
nand U1071 (N_1071,In_245,N_715);
nor U1072 (N_1072,N_954,N_978);
nand U1073 (N_1073,N_341,N_519);
and U1074 (N_1074,N_777,In_204);
xnor U1075 (N_1075,In_1096,N_814);
and U1076 (N_1076,N_313,N_962);
nand U1077 (N_1077,N_548,N_672);
or U1078 (N_1078,N_650,In_776);
xor U1079 (N_1079,N_765,N_380);
or U1080 (N_1080,N_935,N_539);
nor U1081 (N_1081,N_976,N_988);
and U1082 (N_1082,N_966,In_1499);
xor U1083 (N_1083,N_701,In_543);
and U1084 (N_1084,N_865,In_646);
or U1085 (N_1085,N_816,In_1468);
and U1086 (N_1086,In_129,N_998);
nor U1087 (N_1087,N_999,In_1274);
nor U1088 (N_1088,N_973,N_982);
xnor U1089 (N_1089,N_823,N_986);
nand U1090 (N_1090,N_810,N_222);
nor U1091 (N_1091,N_806,N_734);
and U1092 (N_1092,N_606,N_708);
xnor U1093 (N_1093,N_875,N_711);
nand U1094 (N_1094,N_980,N_371);
nor U1095 (N_1095,N_832,N_895);
xnor U1096 (N_1096,N_943,N_780);
nand U1097 (N_1097,In_601,N_815);
nand U1098 (N_1098,N_743,N_625);
nor U1099 (N_1099,In_1306,N_917);
or U1100 (N_1100,N_855,N_858);
or U1101 (N_1101,N_669,N_940);
or U1102 (N_1102,N_942,N_436);
or U1103 (N_1103,N_796,N_245);
nand U1104 (N_1104,In_337,N_419);
xor U1105 (N_1105,N_723,N_951);
xnor U1106 (N_1106,In_296,In_246);
nor U1107 (N_1107,In_463,N_749);
nor U1108 (N_1108,In_203,N_733);
nand U1109 (N_1109,N_607,N_862);
nand U1110 (N_1110,N_878,N_904);
nand U1111 (N_1111,N_848,N_781);
or U1112 (N_1112,In_560,N_879);
nor U1113 (N_1113,N_584,N_638);
or U1114 (N_1114,N_511,N_572);
or U1115 (N_1115,In_79,N_907);
and U1116 (N_1116,N_941,N_842);
nor U1117 (N_1117,N_709,N_698);
nand U1118 (N_1118,N_231,N_863);
nor U1119 (N_1119,N_977,In_1033);
nand U1120 (N_1120,In_577,N_286);
nand U1121 (N_1121,In_453,N_915);
nor U1122 (N_1122,N_850,In_1079);
nor U1123 (N_1123,In_872,In_817);
nand U1124 (N_1124,In_1434,N_961);
and U1125 (N_1125,In_329,N_930);
nor U1126 (N_1126,In_479,In_1379);
and U1127 (N_1127,N_662,N_608);
and U1128 (N_1128,N_665,N_824);
and U1129 (N_1129,N_570,N_17);
nand U1130 (N_1130,N_846,In_908);
or U1131 (N_1131,N_543,N_989);
or U1132 (N_1132,N_979,N_924);
or U1133 (N_1133,N_945,N_731);
and U1134 (N_1134,N_95,N_918);
nor U1135 (N_1135,N_520,N_914);
or U1136 (N_1136,N_423,N_153);
xnor U1137 (N_1137,N_489,N_803);
or U1138 (N_1138,N_496,N_505);
xor U1139 (N_1139,N_316,N_804);
xnor U1140 (N_1140,N_800,N_872);
or U1141 (N_1141,N_382,N_983);
nand U1142 (N_1142,In_1013,N_809);
nand U1143 (N_1143,N_900,N_516);
xor U1144 (N_1144,N_896,N_829);
xnor U1145 (N_1145,N_744,In_563);
or U1146 (N_1146,N_931,N_718);
or U1147 (N_1147,N_871,In_273);
or U1148 (N_1148,N_486,N_831);
xnor U1149 (N_1149,N_819,N_963);
or U1150 (N_1150,N_705,N_922);
nor U1151 (N_1151,N_447,In_917);
and U1152 (N_1152,N_933,N_974);
xnor U1153 (N_1153,N_332,In_88);
nand U1154 (N_1154,N_722,N_799);
nor U1155 (N_1155,N_188,N_870);
or U1156 (N_1156,N_481,In_339);
nor U1157 (N_1157,In_1088,N_408);
and U1158 (N_1158,In_28,N_897);
or U1159 (N_1159,N_833,N_664);
nor U1160 (N_1160,N_852,N_807);
and U1161 (N_1161,N_887,N_517);
and U1162 (N_1162,N_838,N_975);
or U1163 (N_1163,In_730,In_527);
and U1164 (N_1164,N_877,N_844);
and U1165 (N_1165,N_836,In_1338);
nor U1166 (N_1166,N_861,In_410);
and U1167 (N_1167,N_629,In_60);
and U1168 (N_1168,N_514,N_317);
xor U1169 (N_1169,N_769,In_384);
and U1170 (N_1170,N_485,N_891);
nor U1171 (N_1171,N_462,N_714);
xor U1172 (N_1172,N_957,N_601);
and U1173 (N_1173,N_866,N_812);
and U1174 (N_1174,N_318,N_902);
or U1175 (N_1175,N_216,In_806);
and U1176 (N_1176,N_972,N_697);
or U1177 (N_1177,N_580,N_674);
nor U1178 (N_1178,N_355,N_773);
nor U1179 (N_1179,N_826,In_615);
nand U1180 (N_1180,N_953,N_728);
nand U1181 (N_1181,In_1404,N_839);
nor U1182 (N_1182,N_893,N_226);
nand U1183 (N_1183,In_531,N_637);
and U1184 (N_1184,N_929,In_141);
xnor U1185 (N_1185,N_910,In_574);
nand U1186 (N_1186,N_120,N_856);
nand U1187 (N_1187,N_435,N_754);
xor U1188 (N_1188,N_693,N_876);
or U1189 (N_1189,N_956,N_688);
xor U1190 (N_1190,N_703,N_801);
and U1191 (N_1191,N_411,N_492);
nor U1192 (N_1192,N_920,N_939);
nand U1193 (N_1193,In_449,In_1331);
nor U1194 (N_1194,N_936,N_987);
xor U1195 (N_1195,N_985,N_760);
nand U1196 (N_1196,In_98,N_959);
or U1197 (N_1197,N_680,N_890);
nand U1198 (N_1198,N_921,N_928);
xor U1199 (N_1199,N_916,N_903);
and U1200 (N_1200,N_1057,N_1132);
nor U1201 (N_1201,N_603,N_1130);
and U1202 (N_1202,N_1155,N_1027);
nand U1203 (N_1203,N_1018,N_1137);
xor U1204 (N_1204,N_1154,N_612);
and U1205 (N_1205,N_971,N_1047);
xnor U1206 (N_1206,N_23,N_1003);
nand U1207 (N_1207,N_1169,N_785);
xor U1208 (N_1208,N_1085,N_1103);
nor U1209 (N_1209,N_1091,N_1141);
or U1210 (N_1210,N_1134,N_1095);
xor U1211 (N_1211,N_1008,N_1032);
and U1212 (N_1212,N_1054,N_70);
xor U1213 (N_1213,N_783,N_1135);
nand U1214 (N_1214,N_1138,N_1055);
nor U1215 (N_1215,N_1009,N_1168);
xor U1216 (N_1216,N_892,N_1139);
nand U1217 (N_1217,N_1126,N_656);
and U1218 (N_1218,N_860,N_926);
or U1219 (N_1219,N_1053,N_651);
nor U1220 (N_1220,N_1063,N_1046);
xor U1221 (N_1221,N_1038,N_1026);
xnor U1222 (N_1222,N_1024,N_1186);
or U1223 (N_1223,N_1156,N_77);
nor U1224 (N_1224,N_1084,N_1035);
nor U1225 (N_1225,N_480,In_919);
nor U1226 (N_1226,N_964,N_1140);
xor U1227 (N_1227,N_1101,N_1187);
or U1228 (N_1228,N_1111,N_1174);
or U1229 (N_1229,N_1013,N_1121);
or U1230 (N_1230,In_1489,N_446);
and U1231 (N_1231,N_533,N_873);
xnor U1232 (N_1232,N_991,N_894);
xnor U1233 (N_1233,N_1124,N_1184);
xor U1234 (N_1234,In_1068,N_886);
nand U1235 (N_1235,N_1185,N_1039);
nand U1236 (N_1236,N_1192,N_1160);
xor U1237 (N_1237,N_1172,N_1064);
and U1238 (N_1238,N_997,In_1290);
xnor U1239 (N_1239,N_1110,N_1113);
xnor U1240 (N_1240,N_1128,N_536);
nor U1241 (N_1241,N_748,N_1157);
xnor U1242 (N_1242,N_1058,N_898);
and U1243 (N_1243,N_1081,N_716);
and U1244 (N_1244,N_1114,N_990);
or U1245 (N_1245,N_1076,N_1043);
and U1246 (N_1246,In_39,N_851);
nand U1247 (N_1247,N_1000,N_1015);
or U1248 (N_1248,N_1044,N_551);
nand U1249 (N_1249,N_970,In_993);
nor U1250 (N_1250,N_632,N_1096);
or U1251 (N_1251,N_822,N_1198);
nand U1252 (N_1252,N_1183,N_1164);
xnor U1253 (N_1253,N_1078,N_1014);
and U1254 (N_1254,N_1167,N_1123);
nor U1255 (N_1255,N_1161,N_1059);
nand U1256 (N_1256,N_1071,N_845);
nor U1257 (N_1257,In_696,N_1031);
xnor U1258 (N_1258,N_1056,N_1119);
or U1259 (N_1259,N_689,N_1116);
nor U1260 (N_1260,N_1005,N_1067);
and U1261 (N_1261,N_1173,N_1080);
nand U1262 (N_1262,N_736,N_1023);
and U1263 (N_1263,N_968,N_747);
or U1264 (N_1264,N_937,N_828);
nand U1265 (N_1265,N_1131,N_1049);
nand U1266 (N_1266,N_1040,N_830);
xor U1267 (N_1267,N_256,N_1175);
nor U1268 (N_1268,N_1033,N_938);
nand U1269 (N_1269,N_1176,N_1147);
xor U1270 (N_1270,N_1051,N_1118);
nand U1271 (N_1271,N_967,N_1041);
xnor U1272 (N_1272,In_205,N_1087);
or U1273 (N_1273,N_1106,N_1045);
nand U1274 (N_1274,N_1099,N_909);
and U1275 (N_1275,N_1143,N_1102);
nand U1276 (N_1276,N_857,N_1083);
and U1277 (N_1277,N_1117,N_1180);
and U1278 (N_1278,N_1142,N_864);
or U1279 (N_1279,In_846,N_1019);
nor U1280 (N_1280,N_1146,N_1065);
nor U1281 (N_1281,N_1197,In_1377);
nand U1282 (N_1282,N_1165,N_279);
nor U1283 (N_1283,N_1098,N_1199);
and U1284 (N_1284,N_1171,N_1034);
nor U1285 (N_1285,N_1127,N_923);
nand U1286 (N_1286,N_1089,N_1028);
xor U1287 (N_1287,N_1068,N_1148);
nand U1288 (N_1288,N_1152,N_642);
nand U1289 (N_1289,N_1159,N_952);
nor U1290 (N_1290,In_331,N_661);
nor U1291 (N_1291,N_1037,N_1149);
nor U1292 (N_1292,N_1088,N_7);
and U1293 (N_1293,N_1066,N_993);
nor U1294 (N_1294,N_1097,N_1109);
or U1295 (N_1295,N_1129,N_755);
nor U1296 (N_1296,N_1162,N_949);
and U1297 (N_1297,N_981,N_518);
nor U1298 (N_1298,In_793,N_1151);
and U1299 (N_1299,N_1100,N_1125);
or U1300 (N_1300,N_854,N_526);
xnor U1301 (N_1301,N_685,N_757);
nor U1302 (N_1302,N_1011,N_1190);
nor U1303 (N_1303,N_1029,N_1074);
nand U1304 (N_1304,N_1104,N_1191);
or U1305 (N_1305,N_1122,N_1030);
nand U1306 (N_1306,N_1107,N_1115);
or U1307 (N_1307,In_1329,N_1079);
xor U1308 (N_1308,N_1086,N_1050);
and U1309 (N_1309,N_934,N_1108);
or U1310 (N_1310,N_1092,N_821);
nand U1311 (N_1311,N_1052,N_657);
xnor U1312 (N_1312,N_779,N_1145);
xor U1313 (N_1313,N_995,In_608);
or U1314 (N_1314,N_1178,N_1189);
and U1315 (N_1315,N_784,N_1012);
or U1316 (N_1316,In_270,N_1112);
nor U1317 (N_1317,N_837,N_442);
xnor U1318 (N_1318,N_1188,N_1010);
and U1319 (N_1319,N_1001,N_913);
or U1320 (N_1320,N_1177,In_1450);
nor U1321 (N_1321,N_1007,N_1195);
and U1322 (N_1322,N_1006,N_1194);
nand U1323 (N_1323,N_1153,N_1158);
xor U1324 (N_1324,N_1166,N_1070);
or U1325 (N_1325,N_1090,N_1004);
nor U1326 (N_1326,In_976,N_1022);
and U1327 (N_1327,N_1073,N_1061);
or U1328 (N_1328,N_1133,N_835);
and U1329 (N_1329,N_1170,N_1082);
nand U1330 (N_1330,N_1105,N_1069);
or U1331 (N_1331,N_984,N_1163);
nor U1332 (N_1332,In_1367,N_1036);
nand U1333 (N_1333,N_628,N_1144);
nand U1334 (N_1334,N_1077,N_1060);
xnor U1335 (N_1335,N_1094,In_991);
nor U1336 (N_1336,N_284,N_439);
xor U1337 (N_1337,N_1136,N_1042);
xor U1338 (N_1338,In_1261,N_888);
and U1339 (N_1339,N_1017,N_1016);
and U1340 (N_1340,N_1021,N_944);
or U1341 (N_1341,N_1193,N_947);
nand U1342 (N_1342,N_1002,N_1025);
and U1343 (N_1343,N_825,N_1182);
nor U1344 (N_1344,N_1120,N_1181);
nor U1345 (N_1345,N_1196,N_1075);
nand U1346 (N_1346,N_869,N_1150);
nand U1347 (N_1347,N_1093,N_1072);
nor U1348 (N_1348,N_1020,N_1179);
and U1349 (N_1349,N_1048,N_1062);
or U1350 (N_1350,N_1021,N_949);
xor U1351 (N_1351,N_1183,N_1108);
and U1352 (N_1352,N_1182,N_1128);
nor U1353 (N_1353,N_1028,N_1019);
and U1354 (N_1354,N_1053,N_995);
xnor U1355 (N_1355,N_1095,N_1121);
or U1356 (N_1356,N_1013,N_526);
xor U1357 (N_1357,N_551,N_1116);
nor U1358 (N_1358,N_1186,N_1055);
nor U1359 (N_1359,N_1171,N_1003);
xor U1360 (N_1360,N_1044,N_1166);
and U1361 (N_1361,N_1076,N_1080);
nor U1362 (N_1362,N_1004,N_1124);
xor U1363 (N_1363,N_1166,N_830);
xor U1364 (N_1364,N_1093,N_1073);
nor U1365 (N_1365,In_270,N_944);
nand U1366 (N_1366,In_331,N_1139);
nor U1367 (N_1367,N_1007,N_1082);
xor U1368 (N_1368,N_1128,N_1033);
xnor U1369 (N_1369,N_1064,N_968);
nand U1370 (N_1370,N_518,N_1074);
nor U1371 (N_1371,In_1329,N_1070);
nand U1372 (N_1372,N_1051,N_439);
nand U1373 (N_1373,N_1132,In_1367);
xor U1374 (N_1374,N_1060,N_1051);
and U1375 (N_1375,N_854,N_1064);
and U1376 (N_1376,N_1132,N_1134);
and U1377 (N_1377,N_991,N_1164);
nor U1378 (N_1378,N_1014,N_1176);
xor U1379 (N_1379,N_1020,N_1122);
nor U1380 (N_1380,N_1182,N_1070);
xnor U1381 (N_1381,N_1027,N_1104);
nor U1382 (N_1382,N_1140,N_1060);
and U1383 (N_1383,N_1195,In_1489);
nor U1384 (N_1384,N_1198,N_1063);
or U1385 (N_1385,N_1016,In_1329);
nor U1386 (N_1386,N_736,N_284);
and U1387 (N_1387,N_1186,N_1031);
nor U1388 (N_1388,N_1099,N_757);
xor U1389 (N_1389,N_1172,N_1196);
xor U1390 (N_1390,N_1118,N_439);
or U1391 (N_1391,N_1094,N_1018);
and U1392 (N_1392,N_1074,N_892);
and U1393 (N_1393,N_1045,N_612);
or U1394 (N_1394,N_1008,N_1090);
nor U1395 (N_1395,N_1113,N_1183);
or U1396 (N_1396,N_1158,N_442);
xnor U1397 (N_1397,N_964,N_685);
nor U1398 (N_1398,N_1136,N_913);
and U1399 (N_1399,N_1159,N_1141);
xnor U1400 (N_1400,N_1302,N_1297);
nand U1401 (N_1401,N_1309,N_1397);
nor U1402 (N_1402,N_1257,N_1399);
nor U1403 (N_1403,N_1279,N_1294);
or U1404 (N_1404,N_1238,N_1317);
and U1405 (N_1405,N_1291,N_1272);
nor U1406 (N_1406,N_1336,N_1237);
or U1407 (N_1407,N_1305,N_1235);
nor U1408 (N_1408,N_1250,N_1395);
and U1409 (N_1409,N_1204,N_1220);
nand U1410 (N_1410,N_1206,N_1210);
nand U1411 (N_1411,N_1260,N_1222);
xnor U1412 (N_1412,N_1378,N_1278);
and U1413 (N_1413,N_1361,N_1383);
or U1414 (N_1414,N_1229,N_1375);
nor U1415 (N_1415,N_1218,N_1387);
nor U1416 (N_1416,N_1354,N_1345);
and U1417 (N_1417,N_1228,N_1219);
nor U1418 (N_1418,N_1363,N_1271);
and U1419 (N_1419,N_1332,N_1385);
nand U1420 (N_1420,N_1311,N_1256);
xor U1421 (N_1421,N_1348,N_1239);
and U1422 (N_1422,N_1299,N_1356);
xnor U1423 (N_1423,N_1288,N_1337);
xor U1424 (N_1424,N_1236,N_1381);
nand U1425 (N_1425,N_1212,N_1333);
nand U1426 (N_1426,N_1371,N_1328);
nor U1427 (N_1427,N_1200,N_1281);
nand U1428 (N_1428,N_1326,N_1284);
nor U1429 (N_1429,N_1319,N_1254);
nand U1430 (N_1430,N_1308,N_1380);
xnor U1431 (N_1431,N_1230,N_1316);
and U1432 (N_1432,N_1293,N_1350);
nor U1433 (N_1433,N_1394,N_1392);
or U1434 (N_1434,N_1231,N_1384);
nor U1435 (N_1435,N_1285,N_1241);
nand U1436 (N_1436,N_1211,N_1262);
and U1437 (N_1437,N_1259,N_1252);
nand U1438 (N_1438,N_1359,N_1217);
xor U1439 (N_1439,N_1227,N_1379);
and U1440 (N_1440,N_1346,N_1244);
nand U1441 (N_1441,N_1301,N_1360);
nor U1442 (N_1442,N_1327,N_1268);
nor U1443 (N_1443,N_1353,N_1357);
xnor U1444 (N_1444,N_1269,N_1355);
and U1445 (N_1445,N_1292,N_1338);
nand U1446 (N_1446,N_1276,N_1325);
nand U1447 (N_1447,N_1307,N_1286);
or U1448 (N_1448,N_1267,N_1282);
nand U1449 (N_1449,N_1213,N_1358);
nor U1450 (N_1450,N_1369,N_1232);
nor U1451 (N_1451,N_1266,N_1334);
xor U1452 (N_1452,N_1340,N_1234);
nor U1453 (N_1453,N_1270,N_1341);
or U1454 (N_1454,N_1201,N_1249);
xor U1455 (N_1455,N_1388,N_1223);
nor U1456 (N_1456,N_1310,N_1330);
or U1457 (N_1457,N_1209,N_1300);
nand U1458 (N_1458,N_1243,N_1221);
nor U1459 (N_1459,N_1331,N_1208);
and U1460 (N_1460,N_1290,N_1389);
nor U1461 (N_1461,N_1248,N_1374);
and U1462 (N_1462,N_1321,N_1245);
nor U1463 (N_1463,N_1215,N_1233);
nand U1464 (N_1464,N_1362,N_1329);
or U1465 (N_1465,N_1370,N_1277);
nor U1466 (N_1466,N_1261,N_1275);
and U1467 (N_1467,N_1365,N_1376);
nand U1468 (N_1468,N_1226,N_1349);
nor U1469 (N_1469,N_1298,N_1214);
nor U1470 (N_1470,N_1390,N_1313);
or U1471 (N_1471,N_1240,N_1382);
xor U1472 (N_1472,N_1306,N_1373);
xnor U1473 (N_1473,N_1289,N_1372);
nor U1474 (N_1474,N_1246,N_1322);
and U1475 (N_1475,N_1242,N_1205);
and U1476 (N_1476,N_1303,N_1347);
and U1477 (N_1477,N_1258,N_1255);
or U1478 (N_1478,N_1314,N_1202);
xor U1479 (N_1479,N_1203,N_1295);
nand U1480 (N_1480,N_1391,N_1274);
or U1481 (N_1481,N_1396,N_1335);
nor U1482 (N_1482,N_1318,N_1339);
and U1483 (N_1483,N_1366,N_1324);
nand U1484 (N_1484,N_1352,N_1377);
xor U1485 (N_1485,N_1263,N_1315);
or U1486 (N_1486,N_1367,N_1224);
nand U1487 (N_1487,N_1304,N_1323);
or U1488 (N_1488,N_1225,N_1264);
nor U1489 (N_1489,N_1253,N_1283);
nand U1490 (N_1490,N_1265,N_1251);
nand U1491 (N_1491,N_1273,N_1368);
nand U1492 (N_1492,N_1343,N_1247);
xor U1493 (N_1493,N_1312,N_1386);
nor U1494 (N_1494,N_1342,N_1351);
or U1495 (N_1495,N_1216,N_1287);
xor U1496 (N_1496,N_1320,N_1398);
nor U1497 (N_1497,N_1207,N_1296);
xnor U1498 (N_1498,N_1393,N_1280);
nor U1499 (N_1499,N_1344,N_1364);
and U1500 (N_1500,N_1269,N_1215);
or U1501 (N_1501,N_1273,N_1355);
or U1502 (N_1502,N_1375,N_1236);
and U1503 (N_1503,N_1330,N_1229);
nand U1504 (N_1504,N_1391,N_1281);
nor U1505 (N_1505,N_1310,N_1362);
or U1506 (N_1506,N_1386,N_1256);
nor U1507 (N_1507,N_1276,N_1240);
nor U1508 (N_1508,N_1384,N_1295);
xnor U1509 (N_1509,N_1231,N_1397);
xnor U1510 (N_1510,N_1246,N_1397);
and U1511 (N_1511,N_1297,N_1384);
xnor U1512 (N_1512,N_1245,N_1309);
or U1513 (N_1513,N_1300,N_1227);
or U1514 (N_1514,N_1201,N_1312);
nand U1515 (N_1515,N_1215,N_1258);
xnor U1516 (N_1516,N_1326,N_1240);
nand U1517 (N_1517,N_1254,N_1301);
nand U1518 (N_1518,N_1396,N_1389);
nor U1519 (N_1519,N_1205,N_1331);
nor U1520 (N_1520,N_1335,N_1224);
nand U1521 (N_1521,N_1376,N_1383);
xor U1522 (N_1522,N_1360,N_1248);
and U1523 (N_1523,N_1257,N_1232);
xnor U1524 (N_1524,N_1242,N_1355);
or U1525 (N_1525,N_1274,N_1338);
nand U1526 (N_1526,N_1349,N_1322);
xnor U1527 (N_1527,N_1298,N_1327);
xnor U1528 (N_1528,N_1354,N_1356);
nor U1529 (N_1529,N_1382,N_1280);
or U1530 (N_1530,N_1363,N_1356);
and U1531 (N_1531,N_1361,N_1363);
nand U1532 (N_1532,N_1218,N_1379);
or U1533 (N_1533,N_1209,N_1217);
and U1534 (N_1534,N_1331,N_1303);
or U1535 (N_1535,N_1277,N_1323);
nand U1536 (N_1536,N_1314,N_1219);
or U1537 (N_1537,N_1326,N_1224);
and U1538 (N_1538,N_1255,N_1281);
xnor U1539 (N_1539,N_1216,N_1379);
or U1540 (N_1540,N_1369,N_1391);
xnor U1541 (N_1541,N_1336,N_1278);
or U1542 (N_1542,N_1328,N_1257);
xnor U1543 (N_1543,N_1275,N_1257);
and U1544 (N_1544,N_1367,N_1225);
xor U1545 (N_1545,N_1249,N_1237);
nor U1546 (N_1546,N_1304,N_1204);
and U1547 (N_1547,N_1275,N_1367);
nor U1548 (N_1548,N_1399,N_1350);
nand U1549 (N_1549,N_1387,N_1263);
nor U1550 (N_1550,N_1301,N_1362);
and U1551 (N_1551,N_1398,N_1266);
nand U1552 (N_1552,N_1322,N_1255);
or U1553 (N_1553,N_1314,N_1359);
nand U1554 (N_1554,N_1331,N_1266);
nand U1555 (N_1555,N_1333,N_1379);
and U1556 (N_1556,N_1350,N_1336);
nand U1557 (N_1557,N_1264,N_1235);
nor U1558 (N_1558,N_1217,N_1354);
nor U1559 (N_1559,N_1393,N_1390);
and U1560 (N_1560,N_1304,N_1301);
or U1561 (N_1561,N_1298,N_1389);
and U1562 (N_1562,N_1276,N_1381);
xnor U1563 (N_1563,N_1339,N_1289);
nand U1564 (N_1564,N_1223,N_1231);
nor U1565 (N_1565,N_1200,N_1333);
nor U1566 (N_1566,N_1255,N_1344);
nor U1567 (N_1567,N_1335,N_1356);
nand U1568 (N_1568,N_1216,N_1339);
nor U1569 (N_1569,N_1323,N_1366);
or U1570 (N_1570,N_1291,N_1359);
nor U1571 (N_1571,N_1287,N_1219);
nor U1572 (N_1572,N_1363,N_1226);
nand U1573 (N_1573,N_1374,N_1381);
or U1574 (N_1574,N_1341,N_1350);
and U1575 (N_1575,N_1200,N_1388);
or U1576 (N_1576,N_1293,N_1224);
or U1577 (N_1577,N_1293,N_1203);
nand U1578 (N_1578,N_1242,N_1367);
nor U1579 (N_1579,N_1287,N_1382);
nor U1580 (N_1580,N_1298,N_1344);
or U1581 (N_1581,N_1242,N_1398);
xnor U1582 (N_1582,N_1384,N_1301);
and U1583 (N_1583,N_1203,N_1228);
xor U1584 (N_1584,N_1247,N_1384);
xnor U1585 (N_1585,N_1212,N_1315);
nand U1586 (N_1586,N_1231,N_1238);
and U1587 (N_1587,N_1263,N_1389);
nor U1588 (N_1588,N_1374,N_1235);
and U1589 (N_1589,N_1387,N_1315);
nor U1590 (N_1590,N_1290,N_1214);
nand U1591 (N_1591,N_1303,N_1329);
xor U1592 (N_1592,N_1328,N_1332);
and U1593 (N_1593,N_1367,N_1220);
nand U1594 (N_1594,N_1322,N_1376);
xnor U1595 (N_1595,N_1351,N_1298);
nand U1596 (N_1596,N_1205,N_1297);
and U1597 (N_1597,N_1335,N_1380);
or U1598 (N_1598,N_1208,N_1270);
nor U1599 (N_1599,N_1219,N_1245);
nand U1600 (N_1600,N_1471,N_1457);
nand U1601 (N_1601,N_1512,N_1483);
nand U1602 (N_1602,N_1420,N_1593);
nor U1603 (N_1603,N_1418,N_1433);
and U1604 (N_1604,N_1507,N_1545);
and U1605 (N_1605,N_1570,N_1562);
nor U1606 (N_1606,N_1495,N_1442);
nand U1607 (N_1607,N_1500,N_1521);
xnor U1608 (N_1608,N_1590,N_1536);
and U1609 (N_1609,N_1416,N_1489);
or U1610 (N_1610,N_1514,N_1564);
nor U1611 (N_1611,N_1499,N_1488);
or U1612 (N_1612,N_1427,N_1421);
nand U1613 (N_1613,N_1534,N_1410);
or U1614 (N_1614,N_1525,N_1535);
nor U1615 (N_1615,N_1451,N_1468);
nand U1616 (N_1616,N_1419,N_1559);
xnor U1617 (N_1617,N_1437,N_1494);
or U1618 (N_1618,N_1490,N_1448);
and U1619 (N_1619,N_1588,N_1439);
nand U1620 (N_1620,N_1557,N_1572);
xnor U1621 (N_1621,N_1578,N_1596);
and U1622 (N_1622,N_1482,N_1458);
and U1623 (N_1623,N_1585,N_1541);
nor U1624 (N_1624,N_1577,N_1543);
nor U1625 (N_1625,N_1462,N_1426);
xor U1626 (N_1626,N_1425,N_1402);
nand U1627 (N_1627,N_1527,N_1445);
and U1628 (N_1628,N_1444,N_1414);
or U1629 (N_1629,N_1574,N_1424);
nor U1630 (N_1630,N_1520,N_1484);
nand U1631 (N_1631,N_1502,N_1432);
nand U1632 (N_1632,N_1528,N_1563);
nand U1633 (N_1633,N_1455,N_1508);
nand U1634 (N_1634,N_1591,N_1544);
or U1635 (N_1635,N_1517,N_1523);
and U1636 (N_1636,N_1400,N_1430);
or U1637 (N_1637,N_1554,N_1459);
nand U1638 (N_1638,N_1558,N_1581);
or U1639 (N_1639,N_1532,N_1542);
xor U1640 (N_1640,N_1547,N_1479);
or U1641 (N_1641,N_1415,N_1453);
and U1642 (N_1642,N_1515,N_1481);
nand U1643 (N_1643,N_1452,N_1465);
or U1644 (N_1644,N_1549,N_1589);
and U1645 (N_1645,N_1524,N_1472);
nand U1646 (N_1646,N_1551,N_1565);
and U1647 (N_1647,N_1441,N_1503);
and U1648 (N_1648,N_1568,N_1412);
and U1649 (N_1649,N_1449,N_1566);
xnor U1650 (N_1650,N_1576,N_1560);
or U1651 (N_1651,N_1417,N_1539);
nand U1652 (N_1652,N_1413,N_1550);
nor U1653 (N_1653,N_1595,N_1586);
nand U1654 (N_1654,N_1582,N_1493);
nor U1655 (N_1655,N_1429,N_1450);
nor U1656 (N_1656,N_1580,N_1460);
nor U1657 (N_1657,N_1469,N_1599);
and U1658 (N_1658,N_1466,N_1475);
xnor U1659 (N_1659,N_1485,N_1511);
and U1660 (N_1660,N_1467,N_1516);
nand U1661 (N_1661,N_1510,N_1497);
nand U1662 (N_1662,N_1401,N_1478);
or U1663 (N_1663,N_1509,N_1403);
and U1664 (N_1664,N_1538,N_1487);
xor U1665 (N_1665,N_1587,N_1531);
xor U1666 (N_1666,N_1533,N_1409);
nor U1667 (N_1667,N_1546,N_1592);
and U1668 (N_1668,N_1513,N_1438);
nor U1669 (N_1669,N_1405,N_1519);
nand U1670 (N_1670,N_1548,N_1522);
nor U1671 (N_1671,N_1575,N_1431);
nor U1672 (N_1672,N_1561,N_1594);
and U1673 (N_1673,N_1434,N_1447);
xor U1674 (N_1674,N_1537,N_1474);
xnor U1675 (N_1675,N_1470,N_1598);
nand U1676 (N_1676,N_1553,N_1529);
nor U1677 (N_1677,N_1571,N_1404);
or U1678 (N_1678,N_1501,N_1486);
nand U1679 (N_1679,N_1428,N_1492);
xnor U1680 (N_1680,N_1408,N_1443);
nor U1681 (N_1681,N_1491,N_1518);
nor U1682 (N_1682,N_1526,N_1440);
nand U1683 (N_1683,N_1506,N_1556);
nor U1684 (N_1684,N_1436,N_1411);
xnor U1685 (N_1685,N_1579,N_1477);
or U1686 (N_1686,N_1406,N_1435);
nand U1687 (N_1687,N_1584,N_1461);
and U1688 (N_1688,N_1422,N_1463);
and U1689 (N_1689,N_1496,N_1446);
and U1690 (N_1690,N_1498,N_1530);
or U1691 (N_1691,N_1555,N_1569);
xnor U1692 (N_1692,N_1505,N_1464);
and U1693 (N_1693,N_1476,N_1583);
xor U1694 (N_1694,N_1454,N_1597);
or U1695 (N_1695,N_1504,N_1567);
xor U1696 (N_1696,N_1573,N_1540);
and U1697 (N_1697,N_1473,N_1423);
and U1698 (N_1698,N_1552,N_1456);
and U1699 (N_1699,N_1407,N_1480);
xnor U1700 (N_1700,N_1403,N_1499);
or U1701 (N_1701,N_1488,N_1555);
or U1702 (N_1702,N_1500,N_1414);
xnor U1703 (N_1703,N_1452,N_1569);
and U1704 (N_1704,N_1518,N_1481);
nor U1705 (N_1705,N_1480,N_1535);
xor U1706 (N_1706,N_1565,N_1504);
xor U1707 (N_1707,N_1589,N_1574);
nand U1708 (N_1708,N_1494,N_1432);
and U1709 (N_1709,N_1555,N_1473);
or U1710 (N_1710,N_1479,N_1553);
and U1711 (N_1711,N_1503,N_1459);
and U1712 (N_1712,N_1486,N_1447);
nor U1713 (N_1713,N_1448,N_1488);
and U1714 (N_1714,N_1444,N_1417);
nor U1715 (N_1715,N_1473,N_1519);
or U1716 (N_1716,N_1406,N_1487);
xor U1717 (N_1717,N_1417,N_1532);
xor U1718 (N_1718,N_1457,N_1583);
nor U1719 (N_1719,N_1578,N_1551);
xor U1720 (N_1720,N_1567,N_1563);
nor U1721 (N_1721,N_1415,N_1527);
and U1722 (N_1722,N_1424,N_1561);
xor U1723 (N_1723,N_1573,N_1463);
nand U1724 (N_1724,N_1568,N_1542);
xor U1725 (N_1725,N_1434,N_1430);
xnor U1726 (N_1726,N_1521,N_1473);
and U1727 (N_1727,N_1437,N_1442);
and U1728 (N_1728,N_1444,N_1412);
xnor U1729 (N_1729,N_1414,N_1441);
nand U1730 (N_1730,N_1475,N_1523);
and U1731 (N_1731,N_1540,N_1564);
and U1732 (N_1732,N_1410,N_1411);
xor U1733 (N_1733,N_1594,N_1491);
xor U1734 (N_1734,N_1586,N_1460);
nand U1735 (N_1735,N_1452,N_1473);
or U1736 (N_1736,N_1597,N_1414);
nand U1737 (N_1737,N_1554,N_1584);
nor U1738 (N_1738,N_1508,N_1511);
or U1739 (N_1739,N_1451,N_1440);
xnor U1740 (N_1740,N_1586,N_1559);
xnor U1741 (N_1741,N_1489,N_1412);
nand U1742 (N_1742,N_1507,N_1558);
or U1743 (N_1743,N_1598,N_1407);
nor U1744 (N_1744,N_1460,N_1502);
or U1745 (N_1745,N_1482,N_1422);
and U1746 (N_1746,N_1417,N_1475);
nor U1747 (N_1747,N_1484,N_1466);
and U1748 (N_1748,N_1502,N_1489);
nor U1749 (N_1749,N_1527,N_1438);
nand U1750 (N_1750,N_1549,N_1418);
xor U1751 (N_1751,N_1419,N_1587);
or U1752 (N_1752,N_1534,N_1519);
and U1753 (N_1753,N_1584,N_1510);
nor U1754 (N_1754,N_1484,N_1474);
nor U1755 (N_1755,N_1490,N_1546);
nand U1756 (N_1756,N_1498,N_1463);
nand U1757 (N_1757,N_1496,N_1594);
or U1758 (N_1758,N_1418,N_1499);
nand U1759 (N_1759,N_1578,N_1463);
and U1760 (N_1760,N_1585,N_1432);
and U1761 (N_1761,N_1484,N_1401);
and U1762 (N_1762,N_1538,N_1452);
nand U1763 (N_1763,N_1545,N_1516);
nand U1764 (N_1764,N_1581,N_1464);
and U1765 (N_1765,N_1589,N_1426);
or U1766 (N_1766,N_1433,N_1534);
and U1767 (N_1767,N_1499,N_1599);
nand U1768 (N_1768,N_1419,N_1414);
nor U1769 (N_1769,N_1548,N_1479);
nand U1770 (N_1770,N_1427,N_1594);
xnor U1771 (N_1771,N_1522,N_1486);
nand U1772 (N_1772,N_1401,N_1438);
nor U1773 (N_1773,N_1502,N_1465);
or U1774 (N_1774,N_1523,N_1593);
or U1775 (N_1775,N_1445,N_1504);
or U1776 (N_1776,N_1451,N_1429);
nand U1777 (N_1777,N_1428,N_1436);
and U1778 (N_1778,N_1536,N_1496);
nor U1779 (N_1779,N_1574,N_1453);
or U1780 (N_1780,N_1495,N_1537);
or U1781 (N_1781,N_1511,N_1443);
xnor U1782 (N_1782,N_1513,N_1573);
or U1783 (N_1783,N_1473,N_1404);
or U1784 (N_1784,N_1578,N_1589);
nor U1785 (N_1785,N_1508,N_1471);
or U1786 (N_1786,N_1401,N_1549);
or U1787 (N_1787,N_1531,N_1581);
nand U1788 (N_1788,N_1404,N_1570);
nand U1789 (N_1789,N_1477,N_1476);
or U1790 (N_1790,N_1590,N_1496);
nor U1791 (N_1791,N_1476,N_1483);
and U1792 (N_1792,N_1516,N_1451);
nand U1793 (N_1793,N_1538,N_1433);
nor U1794 (N_1794,N_1590,N_1414);
xnor U1795 (N_1795,N_1471,N_1527);
or U1796 (N_1796,N_1559,N_1538);
xnor U1797 (N_1797,N_1483,N_1436);
nor U1798 (N_1798,N_1570,N_1529);
xnor U1799 (N_1799,N_1483,N_1549);
xor U1800 (N_1800,N_1780,N_1686);
or U1801 (N_1801,N_1661,N_1609);
and U1802 (N_1802,N_1719,N_1631);
xnor U1803 (N_1803,N_1668,N_1738);
nand U1804 (N_1804,N_1603,N_1643);
or U1805 (N_1805,N_1684,N_1663);
nor U1806 (N_1806,N_1646,N_1783);
or U1807 (N_1807,N_1605,N_1698);
or U1808 (N_1808,N_1731,N_1674);
and U1809 (N_1809,N_1768,N_1673);
and U1810 (N_1810,N_1737,N_1718);
and U1811 (N_1811,N_1720,N_1650);
xor U1812 (N_1812,N_1680,N_1742);
nand U1813 (N_1813,N_1728,N_1745);
or U1814 (N_1814,N_1608,N_1774);
or U1815 (N_1815,N_1610,N_1788);
and U1816 (N_1816,N_1704,N_1653);
or U1817 (N_1817,N_1724,N_1725);
or U1818 (N_1818,N_1716,N_1658);
nor U1819 (N_1819,N_1775,N_1722);
nor U1820 (N_1820,N_1621,N_1613);
and U1821 (N_1821,N_1797,N_1776);
xor U1822 (N_1822,N_1607,N_1601);
nor U1823 (N_1823,N_1675,N_1623);
or U1824 (N_1824,N_1679,N_1652);
nor U1825 (N_1825,N_1729,N_1767);
or U1826 (N_1826,N_1714,N_1670);
xor U1827 (N_1827,N_1699,N_1666);
nor U1828 (N_1828,N_1696,N_1622);
and U1829 (N_1829,N_1772,N_1693);
xnor U1830 (N_1830,N_1787,N_1701);
xnor U1831 (N_1831,N_1739,N_1754);
xnor U1832 (N_1832,N_1659,N_1749);
nor U1833 (N_1833,N_1752,N_1638);
xor U1834 (N_1834,N_1784,N_1723);
and U1835 (N_1835,N_1604,N_1662);
xor U1836 (N_1836,N_1747,N_1636);
xnor U1837 (N_1837,N_1769,N_1602);
xor U1838 (N_1838,N_1763,N_1672);
xnor U1839 (N_1839,N_1649,N_1606);
and U1840 (N_1840,N_1789,N_1678);
xor U1841 (N_1841,N_1644,N_1667);
nand U1842 (N_1842,N_1713,N_1671);
nand U1843 (N_1843,N_1727,N_1624);
or U1844 (N_1844,N_1695,N_1700);
nand U1845 (N_1845,N_1798,N_1779);
and U1846 (N_1846,N_1721,N_1746);
nand U1847 (N_1847,N_1755,N_1757);
nand U1848 (N_1848,N_1681,N_1703);
or U1849 (N_1849,N_1732,N_1615);
nor U1850 (N_1850,N_1656,N_1785);
xnor U1851 (N_1851,N_1614,N_1765);
nor U1852 (N_1852,N_1733,N_1654);
xor U1853 (N_1853,N_1630,N_1707);
xor U1854 (N_1854,N_1759,N_1611);
or U1855 (N_1855,N_1682,N_1793);
nor U1856 (N_1856,N_1628,N_1710);
nand U1857 (N_1857,N_1619,N_1766);
nand U1858 (N_1858,N_1753,N_1690);
or U1859 (N_1859,N_1773,N_1726);
xnor U1860 (N_1860,N_1758,N_1688);
nand U1861 (N_1861,N_1647,N_1626);
nand U1862 (N_1862,N_1794,N_1734);
nor U1863 (N_1863,N_1655,N_1778);
nand U1864 (N_1864,N_1786,N_1634);
nand U1865 (N_1865,N_1730,N_1687);
and U1866 (N_1866,N_1744,N_1795);
xor U1867 (N_1867,N_1632,N_1669);
nor U1868 (N_1868,N_1705,N_1651);
nand U1869 (N_1869,N_1748,N_1777);
or U1870 (N_1870,N_1642,N_1637);
nor U1871 (N_1871,N_1665,N_1717);
nand U1872 (N_1872,N_1640,N_1639);
or U1873 (N_1873,N_1625,N_1618);
nand U1874 (N_1874,N_1782,N_1741);
xnor U1875 (N_1875,N_1633,N_1697);
nor U1876 (N_1876,N_1600,N_1616);
and U1877 (N_1877,N_1709,N_1711);
or U1878 (N_1878,N_1676,N_1712);
nor U1879 (N_1879,N_1617,N_1751);
xnor U1880 (N_1880,N_1683,N_1708);
xor U1881 (N_1881,N_1694,N_1796);
and U1882 (N_1882,N_1770,N_1677);
nor U1883 (N_1883,N_1781,N_1627);
or U1884 (N_1884,N_1706,N_1660);
and U1885 (N_1885,N_1762,N_1689);
and U1886 (N_1886,N_1629,N_1635);
and U1887 (N_1887,N_1692,N_1743);
nand U1888 (N_1888,N_1791,N_1736);
xor U1889 (N_1889,N_1685,N_1645);
and U1890 (N_1890,N_1691,N_1750);
nor U1891 (N_1891,N_1620,N_1792);
and U1892 (N_1892,N_1641,N_1799);
and U1893 (N_1893,N_1764,N_1761);
or U1894 (N_1894,N_1735,N_1612);
or U1895 (N_1895,N_1756,N_1771);
or U1896 (N_1896,N_1648,N_1702);
and U1897 (N_1897,N_1664,N_1715);
and U1898 (N_1898,N_1790,N_1657);
nor U1899 (N_1899,N_1760,N_1740);
nor U1900 (N_1900,N_1798,N_1614);
xnor U1901 (N_1901,N_1655,N_1638);
and U1902 (N_1902,N_1766,N_1697);
and U1903 (N_1903,N_1734,N_1634);
nand U1904 (N_1904,N_1760,N_1768);
nand U1905 (N_1905,N_1734,N_1688);
nand U1906 (N_1906,N_1719,N_1606);
or U1907 (N_1907,N_1711,N_1793);
or U1908 (N_1908,N_1770,N_1750);
xor U1909 (N_1909,N_1715,N_1619);
or U1910 (N_1910,N_1731,N_1687);
nor U1911 (N_1911,N_1682,N_1670);
xor U1912 (N_1912,N_1603,N_1758);
xnor U1913 (N_1913,N_1614,N_1760);
and U1914 (N_1914,N_1766,N_1779);
nand U1915 (N_1915,N_1634,N_1671);
and U1916 (N_1916,N_1780,N_1663);
and U1917 (N_1917,N_1615,N_1721);
or U1918 (N_1918,N_1667,N_1708);
or U1919 (N_1919,N_1799,N_1751);
xnor U1920 (N_1920,N_1631,N_1658);
nand U1921 (N_1921,N_1782,N_1612);
nor U1922 (N_1922,N_1621,N_1796);
xor U1923 (N_1923,N_1666,N_1694);
or U1924 (N_1924,N_1743,N_1724);
nor U1925 (N_1925,N_1615,N_1760);
nand U1926 (N_1926,N_1601,N_1638);
nand U1927 (N_1927,N_1675,N_1690);
and U1928 (N_1928,N_1744,N_1799);
xnor U1929 (N_1929,N_1677,N_1673);
xor U1930 (N_1930,N_1679,N_1764);
nand U1931 (N_1931,N_1710,N_1754);
xor U1932 (N_1932,N_1687,N_1640);
or U1933 (N_1933,N_1789,N_1745);
nand U1934 (N_1934,N_1754,N_1605);
nor U1935 (N_1935,N_1657,N_1678);
nor U1936 (N_1936,N_1602,N_1741);
nor U1937 (N_1937,N_1793,N_1696);
or U1938 (N_1938,N_1663,N_1616);
and U1939 (N_1939,N_1643,N_1765);
or U1940 (N_1940,N_1625,N_1728);
nor U1941 (N_1941,N_1678,N_1719);
xor U1942 (N_1942,N_1694,N_1690);
nand U1943 (N_1943,N_1689,N_1640);
nand U1944 (N_1944,N_1609,N_1796);
or U1945 (N_1945,N_1729,N_1760);
or U1946 (N_1946,N_1614,N_1618);
nand U1947 (N_1947,N_1727,N_1735);
nor U1948 (N_1948,N_1671,N_1759);
or U1949 (N_1949,N_1710,N_1709);
xnor U1950 (N_1950,N_1799,N_1637);
nor U1951 (N_1951,N_1760,N_1611);
nor U1952 (N_1952,N_1604,N_1771);
nand U1953 (N_1953,N_1789,N_1700);
nor U1954 (N_1954,N_1629,N_1601);
or U1955 (N_1955,N_1704,N_1750);
and U1956 (N_1956,N_1712,N_1779);
or U1957 (N_1957,N_1753,N_1666);
and U1958 (N_1958,N_1626,N_1740);
or U1959 (N_1959,N_1600,N_1745);
nand U1960 (N_1960,N_1603,N_1633);
and U1961 (N_1961,N_1628,N_1788);
xnor U1962 (N_1962,N_1783,N_1678);
nor U1963 (N_1963,N_1669,N_1664);
nor U1964 (N_1964,N_1754,N_1771);
and U1965 (N_1965,N_1628,N_1719);
or U1966 (N_1966,N_1614,N_1707);
xor U1967 (N_1967,N_1689,N_1710);
nor U1968 (N_1968,N_1781,N_1733);
or U1969 (N_1969,N_1682,N_1604);
nor U1970 (N_1970,N_1677,N_1768);
nand U1971 (N_1971,N_1628,N_1718);
or U1972 (N_1972,N_1649,N_1715);
or U1973 (N_1973,N_1647,N_1718);
and U1974 (N_1974,N_1687,N_1697);
or U1975 (N_1975,N_1757,N_1611);
and U1976 (N_1976,N_1754,N_1667);
nor U1977 (N_1977,N_1745,N_1671);
and U1978 (N_1978,N_1627,N_1639);
nand U1979 (N_1979,N_1758,N_1727);
nand U1980 (N_1980,N_1601,N_1753);
and U1981 (N_1981,N_1612,N_1747);
nand U1982 (N_1982,N_1669,N_1640);
nand U1983 (N_1983,N_1711,N_1744);
xnor U1984 (N_1984,N_1714,N_1643);
and U1985 (N_1985,N_1702,N_1767);
nand U1986 (N_1986,N_1643,N_1654);
nor U1987 (N_1987,N_1696,N_1736);
and U1988 (N_1988,N_1691,N_1605);
nand U1989 (N_1989,N_1600,N_1605);
nor U1990 (N_1990,N_1649,N_1711);
or U1991 (N_1991,N_1703,N_1716);
or U1992 (N_1992,N_1794,N_1788);
nand U1993 (N_1993,N_1750,N_1777);
xnor U1994 (N_1994,N_1741,N_1727);
nor U1995 (N_1995,N_1626,N_1608);
or U1996 (N_1996,N_1763,N_1639);
xor U1997 (N_1997,N_1638,N_1617);
xor U1998 (N_1998,N_1725,N_1782);
xor U1999 (N_1999,N_1789,N_1770);
or U2000 (N_2000,N_1850,N_1807);
xor U2001 (N_2001,N_1989,N_1917);
and U2002 (N_2002,N_1809,N_1911);
and U2003 (N_2003,N_1842,N_1889);
nand U2004 (N_2004,N_1866,N_1940);
xnor U2005 (N_2005,N_1855,N_1975);
and U2006 (N_2006,N_1851,N_1860);
nand U2007 (N_2007,N_1991,N_1966);
xor U2008 (N_2008,N_1884,N_1928);
or U2009 (N_2009,N_1969,N_1956);
and U2010 (N_2010,N_1978,N_1857);
nand U2011 (N_2011,N_1952,N_1909);
and U2012 (N_2012,N_1921,N_1823);
and U2013 (N_2013,N_1983,N_1895);
xor U2014 (N_2014,N_1915,N_1878);
or U2015 (N_2015,N_1804,N_1879);
xnor U2016 (N_2016,N_1979,N_1930);
xnor U2017 (N_2017,N_1932,N_1924);
nor U2018 (N_2018,N_1998,N_1808);
nor U2019 (N_2019,N_1962,N_1972);
nor U2020 (N_2020,N_1913,N_1916);
and U2021 (N_2021,N_1936,N_1933);
and U2022 (N_2022,N_1902,N_1992);
and U2023 (N_2023,N_1896,N_1904);
nand U2024 (N_2024,N_1965,N_1869);
nand U2025 (N_2025,N_1802,N_1854);
and U2026 (N_2026,N_1838,N_1931);
and U2027 (N_2027,N_1818,N_1987);
nand U2028 (N_2028,N_1832,N_1872);
and U2029 (N_2029,N_1970,N_1834);
nor U2030 (N_2030,N_1980,N_1927);
nor U2031 (N_2031,N_1893,N_1835);
or U2032 (N_2032,N_1946,N_1988);
and U2033 (N_2033,N_1883,N_1891);
and U2034 (N_2034,N_1925,N_1918);
nor U2035 (N_2035,N_1929,N_1887);
nand U2036 (N_2036,N_1863,N_1945);
nor U2037 (N_2037,N_1938,N_1859);
or U2038 (N_2038,N_1999,N_1821);
xnor U2039 (N_2039,N_1953,N_1833);
and U2040 (N_2040,N_1840,N_1901);
and U2041 (N_2041,N_1812,N_1955);
or U2042 (N_2042,N_1981,N_1995);
nor U2043 (N_2043,N_1881,N_1903);
xor U2044 (N_2044,N_1957,N_1964);
xor U2045 (N_2045,N_1888,N_1845);
xor U2046 (N_2046,N_1828,N_1967);
nor U2047 (N_2047,N_1826,N_1907);
and U2048 (N_2048,N_1856,N_1825);
nand U2049 (N_2049,N_1852,N_1947);
nand U2050 (N_2050,N_1865,N_1900);
nand U2051 (N_2051,N_1977,N_1942);
xnor U2052 (N_2052,N_1959,N_1926);
nor U2053 (N_2053,N_1906,N_1831);
nor U2054 (N_2054,N_1993,N_1912);
and U2055 (N_2055,N_1963,N_1814);
nor U2056 (N_2056,N_1968,N_1829);
and U2057 (N_2057,N_1886,N_1811);
or U2058 (N_2058,N_1876,N_1853);
nand U2059 (N_2059,N_1892,N_1919);
or U2060 (N_2060,N_1848,N_1815);
nand U2061 (N_2061,N_1836,N_1923);
nand U2062 (N_2062,N_1849,N_1867);
nand U2063 (N_2063,N_1871,N_1841);
nand U2064 (N_2064,N_1997,N_1875);
or U2065 (N_2065,N_1939,N_1824);
xnor U2066 (N_2066,N_1974,N_1973);
and U2067 (N_2067,N_1864,N_1934);
xnor U2068 (N_2068,N_1820,N_1844);
or U2069 (N_2069,N_1996,N_1873);
nand U2070 (N_2070,N_1994,N_1908);
and U2071 (N_2071,N_1874,N_1800);
xor U2072 (N_2072,N_1894,N_1958);
and U2073 (N_2073,N_1941,N_1954);
nand U2074 (N_2074,N_1862,N_1898);
or U2075 (N_2075,N_1803,N_1949);
and U2076 (N_2076,N_1897,N_1805);
and U2077 (N_2077,N_1961,N_1806);
nor U2078 (N_2078,N_1948,N_1935);
nand U2079 (N_2079,N_1861,N_1817);
nor U2080 (N_2080,N_1827,N_1971);
or U2081 (N_2081,N_1882,N_1985);
xor U2082 (N_2082,N_1951,N_1885);
and U2083 (N_2083,N_1984,N_1868);
xor U2084 (N_2084,N_1837,N_1846);
xnor U2085 (N_2085,N_1890,N_1870);
nand U2086 (N_2086,N_1990,N_1843);
and U2087 (N_2087,N_1950,N_1910);
nor U2088 (N_2088,N_1960,N_1816);
nor U2089 (N_2089,N_1914,N_1982);
nand U2090 (N_2090,N_1920,N_1822);
nand U2091 (N_2091,N_1986,N_1944);
xor U2092 (N_2092,N_1937,N_1877);
nand U2093 (N_2093,N_1880,N_1839);
or U2094 (N_2094,N_1819,N_1810);
nor U2095 (N_2095,N_1813,N_1830);
or U2096 (N_2096,N_1943,N_1976);
or U2097 (N_2097,N_1899,N_1801);
nor U2098 (N_2098,N_1858,N_1922);
or U2099 (N_2099,N_1905,N_1847);
xnor U2100 (N_2100,N_1930,N_1983);
nor U2101 (N_2101,N_1996,N_1971);
xor U2102 (N_2102,N_1877,N_1986);
xnor U2103 (N_2103,N_1803,N_1819);
nand U2104 (N_2104,N_1852,N_1833);
or U2105 (N_2105,N_1838,N_1996);
nor U2106 (N_2106,N_1803,N_1969);
nand U2107 (N_2107,N_1818,N_1843);
xor U2108 (N_2108,N_1964,N_1896);
xor U2109 (N_2109,N_1915,N_1812);
nor U2110 (N_2110,N_1860,N_1930);
nor U2111 (N_2111,N_1882,N_1837);
and U2112 (N_2112,N_1969,N_1821);
nand U2113 (N_2113,N_1919,N_1900);
nor U2114 (N_2114,N_1994,N_1848);
nor U2115 (N_2115,N_1846,N_1952);
or U2116 (N_2116,N_1974,N_1824);
and U2117 (N_2117,N_1802,N_1879);
or U2118 (N_2118,N_1828,N_1976);
nor U2119 (N_2119,N_1992,N_1935);
xnor U2120 (N_2120,N_1919,N_1995);
nand U2121 (N_2121,N_1953,N_1857);
and U2122 (N_2122,N_1978,N_1925);
nand U2123 (N_2123,N_1949,N_1878);
nor U2124 (N_2124,N_1897,N_1850);
and U2125 (N_2125,N_1895,N_1808);
nand U2126 (N_2126,N_1842,N_1849);
nand U2127 (N_2127,N_1817,N_1844);
nand U2128 (N_2128,N_1861,N_1828);
and U2129 (N_2129,N_1851,N_1906);
nand U2130 (N_2130,N_1824,N_1934);
and U2131 (N_2131,N_1862,N_1922);
nor U2132 (N_2132,N_1982,N_1907);
nor U2133 (N_2133,N_1818,N_1811);
or U2134 (N_2134,N_1888,N_1904);
nand U2135 (N_2135,N_1940,N_1935);
or U2136 (N_2136,N_1922,N_1933);
or U2137 (N_2137,N_1809,N_1806);
nor U2138 (N_2138,N_1843,N_1922);
nor U2139 (N_2139,N_1963,N_1826);
xnor U2140 (N_2140,N_1900,N_1975);
and U2141 (N_2141,N_1864,N_1825);
xor U2142 (N_2142,N_1849,N_1936);
xnor U2143 (N_2143,N_1929,N_1963);
or U2144 (N_2144,N_1828,N_1924);
nor U2145 (N_2145,N_1836,N_1835);
and U2146 (N_2146,N_1866,N_1925);
and U2147 (N_2147,N_1849,N_1831);
and U2148 (N_2148,N_1918,N_1880);
and U2149 (N_2149,N_1929,N_1897);
and U2150 (N_2150,N_1881,N_1937);
and U2151 (N_2151,N_1871,N_1816);
xor U2152 (N_2152,N_1926,N_1937);
nand U2153 (N_2153,N_1992,N_1852);
or U2154 (N_2154,N_1975,N_1836);
nor U2155 (N_2155,N_1838,N_1840);
nand U2156 (N_2156,N_1845,N_1997);
xor U2157 (N_2157,N_1910,N_1899);
xnor U2158 (N_2158,N_1805,N_1926);
xnor U2159 (N_2159,N_1924,N_1859);
and U2160 (N_2160,N_1950,N_1962);
and U2161 (N_2161,N_1934,N_1875);
or U2162 (N_2162,N_1933,N_1885);
xnor U2163 (N_2163,N_1839,N_1829);
xnor U2164 (N_2164,N_1874,N_1926);
xnor U2165 (N_2165,N_1972,N_1827);
and U2166 (N_2166,N_1836,N_1958);
xnor U2167 (N_2167,N_1830,N_1835);
and U2168 (N_2168,N_1941,N_1985);
nand U2169 (N_2169,N_1832,N_1825);
xor U2170 (N_2170,N_1932,N_1827);
and U2171 (N_2171,N_1895,N_1824);
or U2172 (N_2172,N_1899,N_1828);
and U2173 (N_2173,N_1900,N_1883);
and U2174 (N_2174,N_1922,N_1979);
nand U2175 (N_2175,N_1944,N_1915);
and U2176 (N_2176,N_1880,N_1824);
and U2177 (N_2177,N_1935,N_1962);
xor U2178 (N_2178,N_1873,N_1973);
nand U2179 (N_2179,N_1874,N_1967);
or U2180 (N_2180,N_1829,N_1926);
nor U2181 (N_2181,N_1925,N_1824);
and U2182 (N_2182,N_1910,N_1988);
nand U2183 (N_2183,N_1819,N_1961);
nor U2184 (N_2184,N_1846,N_1967);
nor U2185 (N_2185,N_1991,N_1861);
nor U2186 (N_2186,N_1898,N_1872);
or U2187 (N_2187,N_1927,N_1852);
xnor U2188 (N_2188,N_1967,N_1815);
nor U2189 (N_2189,N_1867,N_1971);
and U2190 (N_2190,N_1889,N_1986);
nor U2191 (N_2191,N_1809,N_1857);
and U2192 (N_2192,N_1986,N_1824);
nand U2193 (N_2193,N_1826,N_1945);
xnor U2194 (N_2194,N_1807,N_1968);
nand U2195 (N_2195,N_1937,N_1943);
or U2196 (N_2196,N_1906,N_1938);
xor U2197 (N_2197,N_1984,N_1889);
nor U2198 (N_2198,N_1890,N_1944);
xnor U2199 (N_2199,N_1975,N_1986);
nand U2200 (N_2200,N_2149,N_2074);
xor U2201 (N_2201,N_2128,N_2068);
or U2202 (N_2202,N_2197,N_2043);
and U2203 (N_2203,N_2104,N_2111);
or U2204 (N_2204,N_2057,N_2193);
nand U2205 (N_2205,N_2113,N_2140);
xnor U2206 (N_2206,N_2069,N_2064);
nand U2207 (N_2207,N_2053,N_2150);
and U2208 (N_2208,N_2060,N_2083);
and U2209 (N_2209,N_2198,N_2117);
nand U2210 (N_2210,N_2100,N_2004);
and U2211 (N_2211,N_2186,N_2147);
and U2212 (N_2212,N_2110,N_2070);
nand U2213 (N_2213,N_2001,N_2123);
xnor U2214 (N_2214,N_2167,N_2031);
and U2215 (N_2215,N_2177,N_2036);
nor U2216 (N_2216,N_2054,N_2007);
nand U2217 (N_2217,N_2194,N_2042);
nand U2218 (N_2218,N_2178,N_2181);
xnor U2219 (N_2219,N_2163,N_2089);
nor U2220 (N_2220,N_2059,N_2121);
xor U2221 (N_2221,N_2095,N_2009);
nor U2222 (N_2222,N_2021,N_2152);
nor U2223 (N_2223,N_2048,N_2000);
xnor U2224 (N_2224,N_2024,N_2073);
and U2225 (N_2225,N_2169,N_2046);
nand U2226 (N_2226,N_2188,N_2142);
or U2227 (N_2227,N_2184,N_2028);
xor U2228 (N_2228,N_2047,N_2067);
xor U2229 (N_2229,N_2094,N_2006);
or U2230 (N_2230,N_2081,N_2032);
nand U2231 (N_2231,N_2187,N_2016);
nand U2232 (N_2232,N_2190,N_2130);
nor U2233 (N_2233,N_2191,N_2002);
nand U2234 (N_2234,N_2141,N_2118);
nand U2235 (N_2235,N_2015,N_2099);
or U2236 (N_2236,N_2139,N_2168);
nand U2237 (N_2237,N_2058,N_2122);
nor U2238 (N_2238,N_2125,N_2120);
nor U2239 (N_2239,N_2146,N_2020);
or U2240 (N_2240,N_2077,N_2138);
nand U2241 (N_2241,N_2162,N_2106);
nand U2242 (N_2242,N_2018,N_2112);
or U2243 (N_2243,N_2011,N_2029);
xor U2244 (N_2244,N_2008,N_2101);
nand U2245 (N_2245,N_2185,N_2116);
nor U2246 (N_2246,N_2055,N_2156);
nor U2247 (N_2247,N_2012,N_2086);
or U2248 (N_2248,N_2171,N_2026);
xor U2249 (N_2249,N_2154,N_2153);
nand U2250 (N_2250,N_2033,N_2082);
or U2251 (N_2251,N_2037,N_2114);
nand U2252 (N_2252,N_2051,N_2005);
or U2253 (N_2253,N_2124,N_2131);
nand U2254 (N_2254,N_2078,N_2105);
nand U2255 (N_2255,N_2103,N_2133);
and U2256 (N_2256,N_2136,N_2061);
and U2257 (N_2257,N_2102,N_2161);
xnor U2258 (N_2258,N_2003,N_2041);
nand U2259 (N_2259,N_2052,N_2148);
or U2260 (N_2260,N_2062,N_2092);
nor U2261 (N_2261,N_2071,N_2172);
or U2262 (N_2262,N_2050,N_2196);
or U2263 (N_2263,N_2158,N_2044);
or U2264 (N_2264,N_2175,N_2035);
and U2265 (N_2265,N_2066,N_2049);
nor U2266 (N_2266,N_2065,N_2179);
nor U2267 (N_2267,N_2084,N_2090);
nor U2268 (N_2268,N_2091,N_2159);
nor U2269 (N_2269,N_2034,N_2025);
and U2270 (N_2270,N_2030,N_2098);
nand U2271 (N_2271,N_2109,N_2119);
or U2272 (N_2272,N_2108,N_2038);
xor U2273 (N_2273,N_2165,N_2027);
and U2274 (N_2274,N_2155,N_2063);
nand U2275 (N_2275,N_2097,N_2166);
nor U2276 (N_2276,N_2072,N_2039);
or U2277 (N_2277,N_2144,N_2022);
xor U2278 (N_2278,N_2173,N_2085);
or U2279 (N_2279,N_2157,N_2134);
or U2280 (N_2280,N_2013,N_2174);
nor U2281 (N_2281,N_2132,N_2096);
nor U2282 (N_2282,N_2087,N_2129);
xnor U2283 (N_2283,N_2080,N_2145);
and U2284 (N_2284,N_2010,N_2107);
nor U2285 (N_2285,N_2164,N_2183);
or U2286 (N_2286,N_2176,N_2199);
and U2287 (N_2287,N_2115,N_2045);
xor U2288 (N_2288,N_2180,N_2076);
xor U2289 (N_2289,N_2192,N_2127);
nand U2290 (N_2290,N_2079,N_2182);
nand U2291 (N_2291,N_2170,N_2137);
xor U2292 (N_2292,N_2056,N_2126);
nand U2293 (N_2293,N_2143,N_2040);
nand U2294 (N_2294,N_2088,N_2023);
or U2295 (N_2295,N_2135,N_2017);
nor U2296 (N_2296,N_2019,N_2160);
and U2297 (N_2297,N_2014,N_2189);
or U2298 (N_2298,N_2151,N_2093);
xnor U2299 (N_2299,N_2195,N_2075);
nor U2300 (N_2300,N_2015,N_2028);
nand U2301 (N_2301,N_2058,N_2031);
and U2302 (N_2302,N_2075,N_2048);
nand U2303 (N_2303,N_2138,N_2000);
and U2304 (N_2304,N_2042,N_2051);
or U2305 (N_2305,N_2184,N_2135);
xnor U2306 (N_2306,N_2033,N_2109);
nor U2307 (N_2307,N_2025,N_2127);
xnor U2308 (N_2308,N_2009,N_2082);
and U2309 (N_2309,N_2071,N_2194);
nor U2310 (N_2310,N_2020,N_2123);
and U2311 (N_2311,N_2048,N_2149);
and U2312 (N_2312,N_2111,N_2082);
and U2313 (N_2313,N_2093,N_2035);
or U2314 (N_2314,N_2194,N_2113);
nor U2315 (N_2315,N_2148,N_2030);
and U2316 (N_2316,N_2113,N_2164);
xor U2317 (N_2317,N_2105,N_2053);
or U2318 (N_2318,N_2003,N_2020);
xor U2319 (N_2319,N_2107,N_2158);
and U2320 (N_2320,N_2151,N_2068);
nand U2321 (N_2321,N_2020,N_2050);
and U2322 (N_2322,N_2127,N_2161);
and U2323 (N_2323,N_2183,N_2059);
xnor U2324 (N_2324,N_2173,N_2058);
or U2325 (N_2325,N_2198,N_2158);
nand U2326 (N_2326,N_2070,N_2105);
xor U2327 (N_2327,N_2116,N_2166);
xnor U2328 (N_2328,N_2056,N_2034);
nand U2329 (N_2329,N_2135,N_2155);
and U2330 (N_2330,N_2193,N_2150);
and U2331 (N_2331,N_2070,N_2168);
nand U2332 (N_2332,N_2195,N_2042);
or U2333 (N_2333,N_2192,N_2092);
xnor U2334 (N_2334,N_2043,N_2054);
xor U2335 (N_2335,N_2158,N_2173);
xnor U2336 (N_2336,N_2015,N_2145);
xor U2337 (N_2337,N_2103,N_2109);
and U2338 (N_2338,N_2177,N_2186);
nor U2339 (N_2339,N_2073,N_2138);
and U2340 (N_2340,N_2164,N_2199);
or U2341 (N_2341,N_2189,N_2060);
xor U2342 (N_2342,N_2070,N_2122);
xnor U2343 (N_2343,N_2166,N_2041);
nor U2344 (N_2344,N_2076,N_2022);
nand U2345 (N_2345,N_2020,N_2140);
or U2346 (N_2346,N_2141,N_2116);
xnor U2347 (N_2347,N_2141,N_2040);
nand U2348 (N_2348,N_2135,N_2029);
nand U2349 (N_2349,N_2163,N_2127);
nor U2350 (N_2350,N_2119,N_2103);
nor U2351 (N_2351,N_2042,N_2177);
nor U2352 (N_2352,N_2094,N_2189);
nand U2353 (N_2353,N_2014,N_2037);
nand U2354 (N_2354,N_2163,N_2181);
or U2355 (N_2355,N_2130,N_2003);
and U2356 (N_2356,N_2054,N_2077);
or U2357 (N_2357,N_2116,N_2031);
nand U2358 (N_2358,N_2046,N_2196);
or U2359 (N_2359,N_2108,N_2155);
xor U2360 (N_2360,N_2157,N_2012);
nor U2361 (N_2361,N_2059,N_2155);
nand U2362 (N_2362,N_2122,N_2130);
or U2363 (N_2363,N_2072,N_2032);
nor U2364 (N_2364,N_2045,N_2091);
or U2365 (N_2365,N_2135,N_2043);
or U2366 (N_2366,N_2110,N_2024);
or U2367 (N_2367,N_2114,N_2018);
nand U2368 (N_2368,N_2199,N_2099);
xnor U2369 (N_2369,N_2120,N_2080);
xnor U2370 (N_2370,N_2180,N_2017);
and U2371 (N_2371,N_2117,N_2078);
xnor U2372 (N_2372,N_2014,N_2155);
or U2373 (N_2373,N_2038,N_2071);
or U2374 (N_2374,N_2147,N_2090);
nor U2375 (N_2375,N_2078,N_2011);
or U2376 (N_2376,N_2154,N_2028);
nand U2377 (N_2377,N_2150,N_2198);
and U2378 (N_2378,N_2060,N_2179);
or U2379 (N_2379,N_2153,N_2043);
nand U2380 (N_2380,N_2019,N_2116);
nand U2381 (N_2381,N_2138,N_2045);
or U2382 (N_2382,N_2016,N_2129);
nand U2383 (N_2383,N_2157,N_2195);
xnor U2384 (N_2384,N_2048,N_2081);
xnor U2385 (N_2385,N_2096,N_2151);
or U2386 (N_2386,N_2031,N_2081);
nor U2387 (N_2387,N_2063,N_2152);
and U2388 (N_2388,N_2027,N_2129);
nor U2389 (N_2389,N_2188,N_2112);
xnor U2390 (N_2390,N_2080,N_2143);
xor U2391 (N_2391,N_2016,N_2095);
or U2392 (N_2392,N_2119,N_2165);
nor U2393 (N_2393,N_2064,N_2032);
xnor U2394 (N_2394,N_2109,N_2077);
xor U2395 (N_2395,N_2134,N_2012);
nor U2396 (N_2396,N_2034,N_2008);
nand U2397 (N_2397,N_2001,N_2194);
and U2398 (N_2398,N_2144,N_2113);
nor U2399 (N_2399,N_2119,N_2181);
xor U2400 (N_2400,N_2238,N_2283);
nand U2401 (N_2401,N_2287,N_2278);
nand U2402 (N_2402,N_2267,N_2268);
and U2403 (N_2403,N_2348,N_2277);
nand U2404 (N_2404,N_2366,N_2223);
xor U2405 (N_2405,N_2334,N_2376);
nand U2406 (N_2406,N_2386,N_2211);
nand U2407 (N_2407,N_2378,N_2212);
nor U2408 (N_2408,N_2328,N_2347);
and U2409 (N_2409,N_2266,N_2219);
or U2410 (N_2410,N_2203,N_2246);
or U2411 (N_2411,N_2375,N_2396);
nand U2412 (N_2412,N_2292,N_2352);
nand U2413 (N_2413,N_2325,N_2356);
or U2414 (N_2414,N_2202,N_2382);
nand U2415 (N_2415,N_2363,N_2354);
nor U2416 (N_2416,N_2216,N_2385);
or U2417 (N_2417,N_2384,N_2231);
xnor U2418 (N_2418,N_2389,N_2339);
nor U2419 (N_2419,N_2372,N_2313);
nand U2420 (N_2420,N_2380,N_2275);
and U2421 (N_2421,N_2254,N_2258);
xnor U2422 (N_2422,N_2239,N_2324);
xnor U2423 (N_2423,N_2321,N_2322);
and U2424 (N_2424,N_2251,N_2377);
xnor U2425 (N_2425,N_2227,N_2320);
or U2426 (N_2426,N_2312,N_2236);
and U2427 (N_2427,N_2242,N_2263);
and U2428 (N_2428,N_2333,N_2346);
xnor U2429 (N_2429,N_2337,N_2374);
and U2430 (N_2430,N_2270,N_2280);
xor U2431 (N_2431,N_2255,N_2341);
nand U2432 (N_2432,N_2397,N_2234);
xnor U2433 (N_2433,N_2391,N_2226);
nor U2434 (N_2434,N_2210,N_2332);
nand U2435 (N_2435,N_2379,N_2349);
nor U2436 (N_2436,N_2230,N_2300);
nand U2437 (N_2437,N_2273,N_2284);
nor U2438 (N_2438,N_2303,N_2271);
nor U2439 (N_2439,N_2276,N_2235);
nand U2440 (N_2440,N_2344,N_2297);
nor U2441 (N_2441,N_2381,N_2316);
nand U2442 (N_2442,N_2357,N_2318);
nor U2443 (N_2443,N_2317,N_2248);
nand U2444 (N_2444,N_2304,N_2253);
xnor U2445 (N_2445,N_2359,N_2388);
nor U2446 (N_2446,N_2244,N_2250);
nand U2447 (N_2447,N_2286,N_2272);
or U2448 (N_2448,N_2314,N_2308);
and U2449 (N_2449,N_2338,N_2310);
xor U2450 (N_2450,N_2257,N_2285);
xor U2451 (N_2451,N_2256,N_2241);
and U2452 (N_2452,N_2383,N_2201);
and U2453 (N_2453,N_2259,N_2370);
nor U2454 (N_2454,N_2291,N_2247);
or U2455 (N_2455,N_2398,N_2206);
and U2456 (N_2456,N_2262,N_2387);
or U2457 (N_2457,N_2243,N_2340);
nor U2458 (N_2458,N_2331,N_2290);
nor U2459 (N_2459,N_2245,N_2336);
nand U2460 (N_2460,N_2369,N_2345);
xnor U2461 (N_2461,N_2204,N_2302);
and U2462 (N_2462,N_2252,N_2289);
nor U2463 (N_2463,N_2295,N_2205);
nand U2464 (N_2464,N_2335,N_2364);
and U2465 (N_2465,N_2265,N_2360);
and U2466 (N_2466,N_2233,N_2309);
or U2467 (N_2467,N_2373,N_2330);
nand U2468 (N_2468,N_2208,N_2293);
xnor U2469 (N_2469,N_2240,N_2368);
or U2470 (N_2470,N_2367,N_2319);
and U2471 (N_2471,N_2260,N_2294);
xor U2472 (N_2472,N_2323,N_2281);
xnor U2473 (N_2473,N_2269,N_2249);
xor U2474 (N_2474,N_2355,N_2307);
nand U2475 (N_2475,N_2301,N_2299);
nor U2476 (N_2476,N_2288,N_2298);
nor U2477 (N_2477,N_2214,N_2264);
nand U2478 (N_2478,N_2315,N_2221);
xnor U2479 (N_2479,N_2343,N_2327);
or U2480 (N_2480,N_2358,N_2353);
nand U2481 (N_2481,N_2200,N_2225);
and U2482 (N_2482,N_2362,N_2279);
xor U2483 (N_2483,N_2213,N_2220);
or U2484 (N_2484,N_2274,N_2390);
nand U2485 (N_2485,N_2394,N_2305);
nor U2486 (N_2486,N_2296,N_2311);
or U2487 (N_2487,N_2399,N_2224);
or U2488 (N_2488,N_2361,N_2326);
nor U2489 (N_2489,N_2207,N_2342);
and U2490 (N_2490,N_2237,N_2393);
or U2491 (N_2491,N_2228,N_2395);
and U2492 (N_2492,N_2232,N_2218);
nor U2493 (N_2493,N_2351,N_2371);
nor U2494 (N_2494,N_2306,N_2365);
or U2495 (N_2495,N_2261,N_2217);
or U2496 (N_2496,N_2282,N_2215);
and U2497 (N_2497,N_2229,N_2392);
and U2498 (N_2498,N_2209,N_2350);
nor U2499 (N_2499,N_2222,N_2329);
nand U2500 (N_2500,N_2377,N_2253);
nand U2501 (N_2501,N_2213,N_2366);
nand U2502 (N_2502,N_2337,N_2286);
and U2503 (N_2503,N_2273,N_2398);
xor U2504 (N_2504,N_2380,N_2351);
nor U2505 (N_2505,N_2337,N_2200);
or U2506 (N_2506,N_2301,N_2226);
nor U2507 (N_2507,N_2224,N_2270);
nand U2508 (N_2508,N_2301,N_2319);
xnor U2509 (N_2509,N_2281,N_2352);
xor U2510 (N_2510,N_2277,N_2259);
nand U2511 (N_2511,N_2351,N_2363);
nor U2512 (N_2512,N_2231,N_2274);
nor U2513 (N_2513,N_2305,N_2278);
nand U2514 (N_2514,N_2324,N_2255);
xnor U2515 (N_2515,N_2232,N_2332);
nand U2516 (N_2516,N_2261,N_2255);
nand U2517 (N_2517,N_2320,N_2394);
nand U2518 (N_2518,N_2370,N_2397);
nand U2519 (N_2519,N_2268,N_2373);
nor U2520 (N_2520,N_2243,N_2322);
xnor U2521 (N_2521,N_2322,N_2287);
and U2522 (N_2522,N_2216,N_2243);
nor U2523 (N_2523,N_2318,N_2379);
or U2524 (N_2524,N_2369,N_2299);
nor U2525 (N_2525,N_2300,N_2253);
xnor U2526 (N_2526,N_2274,N_2215);
nor U2527 (N_2527,N_2300,N_2257);
xnor U2528 (N_2528,N_2371,N_2377);
and U2529 (N_2529,N_2215,N_2239);
and U2530 (N_2530,N_2395,N_2279);
or U2531 (N_2531,N_2240,N_2366);
xor U2532 (N_2532,N_2366,N_2395);
xnor U2533 (N_2533,N_2278,N_2362);
nand U2534 (N_2534,N_2271,N_2215);
and U2535 (N_2535,N_2257,N_2319);
and U2536 (N_2536,N_2337,N_2253);
or U2537 (N_2537,N_2242,N_2295);
nor U2538 (N_2538,N_2233,N_2386);
or U2539 (N_2539,N_2340,N_2328);
and U2540 (N_2540,N_2276,N_2229);
nor U2541 (N_2541,N_2300,N_2378);
and U2542 (N_2542,N_2386,N_2339);
xnor U2543 (N_2543,N_2354,N_2345);
or U2544 (N_2544,N_2298,N_2229);
nand U2545 (N_2545,N_2332,N_2353);
or U2546 (N_2546,N_2258,N_2304);
nand U2547 (N_2547,N_2356,N_2312);
and U2548 (N_2548,N_2272,N_2297);
xor U2549 (N_2549,N_2266,N_2284);
nand U2550 (N_2550,N_2349,N_2290);
nand U2551 (N_2551,N_2377,N_2365);
nand U2552 (N_2552,N_2366,N_2359);
nor U2553 (N_2553,N_2309,N_2354);
nor U2554 (N_2554,N_2389,N_2320);
nor U2555 (N_2555,N_2234,N_2386);
nand U2556 (N_2556,N_2338,N_2340);
nor U2557 (N_2557,N_2282,N_2309);
nand U2558 (N_2558,N_2231,N_2329);
nand U2559 (N_2559,N_2338,N_2231);
and U2560 (N_2560,N_2288,N_2203);
and U2561 (N_2561,N_2367,N_2270);
nand U2562 (N_2562,N_2278,N_2319);
nand U2563 (N_2563,N_2347,N_2217);
xnor U2564 (N_2564,N_2326,N_2370);
xor U2565 (N_2565,N_2308,N_2313);
nor U2566 (N_2566,N_2346,N_2203);
and U2567 (N_2567,N_2364,N_2242);
nand U2568 (N_2568,N_2272,N_2394);
and U2569 (N_2569,N_2380,N_2321);
nor U2570 (N_2570,N_2266,N_2375);
xnor U2571 (N_2571,N_2316,N_2240);
and U2572 (N_2572,N_2386,N_2370);
and U2573 (N_2573,N_2313,N_2327);
nor U2574 (N_2574,N_2262,N_2305);
and U2575 (N_2575,N_2316,N_2274);
and U2576 (N_2576,N_2340,N_2303);
xnor U2577 (N_2577,N_2265,N_2355);
nand U2578 (N_2578,N_2216,N_2335);
nor U2579 (N_2579,N_2231,N_2250);
xor U2580 (N_2580,N_2280,N_2372);
xnor U2581 (N_2581,N_2302,N_2395);
xnor U2582 (N_2582,N_2333,N_2377);
nor U2583 (N_2583,N_2315,N_2332);
and U2584 (N_2584,N_2254,N_2370);
nor U2585 (N_2585,N_2320,N_2310);
or U2586 (N_2586,N_2264,N_2387);
nand U2587 (N_2587,N_2285,N_2269);
nor U2588 (N_2588,N_2383,N_2213);
and U2589 (N_2589,N_2386,N_2267);
nor U2590 (N_2590,N_2305,N_2220);
nor U2591 (N_2591,N_2225,N_2395);
nand U2592 (N_2592,N_2385,N_2349);
xor U2593 (N_2593,N_2338,N_2237);
xnor U2594 (N_2594,N_2315,N_2326);
and U2595 (N_2595,N_2301,N_2391);
nand U2596 (N_2596,N_2321,N_2294);
and U2597 (N_2597,N_2291,N_2372);
or U2598 (N_2598,N_2330,N_2341);
and U2599 (N_2599,N_2360,N_2243);
xnor U2600 (N_2600,N_2578,N_2501);
and U2601 (N_2601,N_2446,N_2593);
nor U2602 (N_2602,N_2573,N_2544);
or U2603 (N_2603,N_2525,N_2478);
xnor U2604 (N_2604,N_2435,N_2418);
or U2605 (N_2605,N_2451,N_2471);
or U2606 (N_2606,N_2519,N_2511);
nand U2607 (N_2607,N_2590,N_2551);
xor U2608 (N_2608,N_2595,N_2427);
nor U2609 (N_2609,N_2434,N_2528);
nand U2610 (N_2610,N_2537,N_2543);
nor U2611 (N_2611,N_2524,N_2444);
and U2612 (N_2612,N_2574,N_2514);
xor U2613 (N_2613,N_2438,N_2422);
and U2614 (N_2614,N_2547,N_2483);
xnor U2615 (N_2615,N_2541,N_2405);
nand U2616 (N_2616,N_2414,N_2439);
nand U2617 (N_2617,N_2469,N_2576);
nor U2618 (N_2618,N_2538,N_2581);
and U2619 (N_2619,N_2443,N_2430);
and U2620 (N_2620,N_2489,N_2415);
and U2621 (N_2621,N_2557,N_2496);
nand U2622 (N_2622,N_2515,N_2424);
xor U2623 (N_2623,N_2485,N_2456);
or U2624 (N_2624,N_2417,N_2440);
and U2625 (N_2625,N_2453,N_2532);
nor U2626 (N_2626,N_2487,N_2416);
nor U2627 (N_2627,N_2502,N_2400);
or U2628 (N_2628,N_2539,N_2466);
nand U2629 (N_2629,N_2568,N_2580);
nand U2630 (N_2630,N_2570,N_2500);
or U2631 (N_2631,N_2591,N_2582);
nand U2632 (N_2632,N_2504,N_2512);
nand U2633 (N_2633,N_2429,N_2455);
nand U2634 (N_2634,N_2413,N_2472);
or U2635 (N_2635,N_2588,N_2594);
and U2636 (N_2636,N_2470,N_2592);
xnor U2637 (N_2637,N_2481,N_2490);
xnor U2638 (N_2638,N_2571,N_2423);
and U2639 (N_2639,N_2495,N_2565);
nor U2640 (N_2640,N_2403,N_2549);
nor U2641 (N_2641,N_2503,N_2412);
xor U2642 (N_2642,N_2420,N_2529);
or U2643 (N_2643,N_2499,N_2513);
and U2644 (N_2644,N_2535,N_2561);
or U2645 (N_2645,N_2461,N_2542);
xnor U2646 (N_2646,N_2583,N_2431);
or U2647 (N_2647,N_2520,N_2493);
and U2648 (N_2648,N_2567,N_2458);
or U2649 (N_2649,N_2559,N_2584);
or U2650 (N_2650,N_2505,N_2476);
xnor U2651 (N_2651,N_2442,N_2441);
and U2652 (N_2652,N_2425,N_2509);
nand U2653 (N_2653,N_2468,N_2596);
and U2654 (N_2654,N_2457,N_2460);
nand U2655 (N_2655,N_2421,N_2419);
or U2656 (N_2656,N_2477,N_2527);
and U2657 (N_2657,N_2564,N_2410);
or U2658 (N_2658,N_2552,N_2506);
nand U2659 (N_2659,N_2569,N_2406);
xnor U2660 (N_2660,N_2550,N_2518);
and U2661 (N_2661,N_2562,N_2560);
and U2662 (N_2662,N_2548,N_2599);
and U2663 (N_2663,N_2467,N_2597);
nor U2664 (N_2664,N_2407,N_2587);
or U2665 (N_2665,N_2436,N_2409);
nor U2666 (N_2666,N_2450,N_2426);
nand U2667 (N_2667,N_2445,N_2598);
nor U2668 (N_2668,N_2517,N_2411);
or U2669 (N_2669,N_2531,N_2523);
or U2670 (N_2670,N_2526,N_2579);
and U2671 (N_2671,N_2482,N_2408);
or U2672 (N_2672,N_2516,N_2558);
and U2673 (N_2673,N_2473,N_2463);
and U2674 (N_2674,N_2586,N_2454);
xnor U2675 (N_2675,N_2452,N_2572);
nor U2676 (N_2676,N_2554,N_2556);
nor U2677 (N_2677,N_2491,N_2459);
nor U2678 (N_2678,N_2494,N_2585);
nand U2679 (N_2679,N_2534,N_2464);
nand U2680 (N_2680,N_2589,N_2486);
xnor U2681 (N_2681,N_2566,N_2428);
and U2682 (N_2682,N_2546,N_2510);
or U2683 (N_2683,N_2449,N_2484);
or U2684 (N_2684,N_2507,N_2479);
xnor U2685 (N_2685,N_2480,N_2540);
and U2686 (N_2686,N_2488,N_2475);
nor U2687 (N_2687,N_2577,N_2437);
nor U2688 (N_2688,N_2497,N_2563);
nor U2689 (N_2689,N_2498,N_2521);
and U2690 (N_2690,N_2522,N_2508);
and U2691 (N_2691,N_2492,N_2402);
nand U2692 (N_2692,N_2575,N_2474);
xnor U2693 (N_2693,N_2404,N_2462);
xnor U2694 (N_2694,N_2530,N_2433);
and U2695 (N_2695,N_2401,N_2555);
and U2696 (N_2696,N_2536,N_2553);
or U2697 (N_2697,N_2545,N_2533);
xor U2698 (N_2698,N_2447,N_2448);
nor U2699 (N_2699,N_2465,N_2432);
xor U2700 (N_2700,N_2507,N_2481);
and U2701 (N_2701,N_2411,N_2514);
and U2702 (N_2702,N_2428,N_2538);
nor U2703 (N_2703,N_2409,N_2435);
and U2704 (N_2704,N_2509,N_2424);
or U2705 (N_2705,N_2539,N_2544);
and U2706 (N_2706,N_2507,N_2510);
nand U2707 (N_2707,N_2429,N_2524);
or U2708 (N_2708,N_2482,N_2590);
nor U2709 (N_2709,N_2595,N_2494);
xnor U2710 (N_2710,N_2520,N_2564);
or U2711 (N_2711,N_2541,N_2457);
xor U2712 (N_2712,N_2511,N_2597);
nand U2713 (N_2713,N_2491,N_2564);
or U2714 (N_2714,N_2517,N_2465);
and U2715 (N_2715,N_2519,N_2427);
and U2716 (N_2716,N_2410,N_2520);
nor U2717 (N_2717,N_2527,N_2521);
and U2718 (N_2718,N_2409,N_2575);
or U2719 (N_2719,N_2411,N_2585);
or U2720 (N_2720,N_2556,N_2405);
or U2721 (N_2721,N_2543,N_2584);
nor U2722 (N_2722,N_2408,N_2575);
nand U2723 (N_2723,N_2429,N_2431);
nand U2724 (N_2724,N_2417,N_2557);
and U2725 (N_2725,N_2486,N_2540);
nor U2726 (N_2726,N_2414,N_2470);
nor U2727 (N_2727,N_2556,N_2569);
nor U2728 (N_2728,N_2456,N_2565);
or U2729 (N_2729,N_2443,N_2416);
nor U2730 (N_2730,N_2587,N_2446);
or U2731 (N_2731,N_2529,N_2485);
and U2732 (N_2732,N_2596,N_2525);
xnor U2733 (N_2733,N_2582,N_2552);
xnor U2734 (N_2734,N_2501,N_2486);
xnor U2735 (N_2735,N_2486,N_2518);
nor U2736 (N_2736,N_2449,N_2415);
nor U2737 (N_2737,N_2556,N_2524);
xnor U2738 (N_2738,N_2420,N_2461);
nor U2739 (N_2739,N_2511,N_2513);
and U2740 (N_2740,N_2575,N_2573);
or U2741 (N_2741,N_2406,N_2519);
xor U2742 (N_2742,N_2427,N_2594);
xor U2743 (N_2743,N_2446,N_2490);
and U2744 (N_2744,N_2424,N_2560);
nor U2745 (N_2745,N_2507,N_2474);
xor U2746 (N_2746,N_2526,N_2521);
or U2747 (N_2747,N_2459,N_2596);
xor U2748 (N_2748,N_2597,N_2588);
and U2749 (N_2749,N_2434,N_2499);
and U2750 (N_2750,N_2534,N_2567);
and U2751 (N_2751,N_2596,N_2450);
and U2752 (N_2752,N_2465,N_2481);
nor U2753 (N_2753,N_2505,N_2448);
nor U2754 (N_2754,N_2573,N_2444);
nand U2755 (N_2755,N_2492,N_2543);
xor U2756 (N_2756,N_2480,N_2411);
and U2757 (N_2757,N_2450,N_2405);
xor U2758 (N_2758,N_2568,N_2436);
nor U2759 (N_2759,N_2453,N_2442);
and U2760 (N_2760,N_2585,N_2453);
and U2761 (N_2761,N_2512,N_2555);
or U2762 (N_2762,N_2490,N_2428);
xnor U2763 (N_2763,N_2488,N_2532);
xnor U2764 (N_2764,N_2533,N_2551);
xnor U2765 (N_2765,N_2444,N_2458);
xnor U2766 (N_2766,N_2447,N_2485);
xor U2767 (N_2767,N_2519,N_2436);
and U2768 (N_2768,N_2579,N_2477);
or U2769 (N_2769,N_2531,N_2535);
xnor U2770 (N_2770,N_2463,N_2461);
nor U2771 (N_2771,N_2573,N_2588);
nor U2772 (N_2772,N_2419,N_2457);
nor U2773 (N_2773,N_2567,N_2594);
or U2774 (N_2774,N_2426,N_2491);
xnor U2775 (N_2775,N_2401,N_2473);
or U2776 (N_2776,N_2583,N_2559);
xnor U2777 (N_2777,N_2416,N_2576);
xor U2778 (N_2778,N_2455,N_2511);
and U2779 (N_2779,N_2447,N_2425);
and U2780 (N_2780,N_2422,N_2501);
nand U2781 (N_2781,N_2440,N_2536);
nor U2782 (N_2782,N_2590,N_2465);
and U2783 (N_2783,N_2464,N_2508);
nand U2784 (N_2784,N_2565,N_2418);
nor U2785 (N_2785,N_2509,N_2572);
or U2786 (N_2786,N_2510,N_2569);
xor U2787 (N_2787,N_2492,N_2498);
nor U2788 (N_2788,N_2450,N_2406);
xor U2789 (N_2789,N_2428,N_2544);
nand U2790 (N_2790,N_2575,N_2547);
xor U2791 (N_2791,N_2441,N_2467);
and U2792 (N_2792,N_2462,N_2581);
and U2793 (N_2793,N_2590,N_2544);
xnor U2794 (N_2794,N_2407,N_2476);
xnor U2795 (N_2795,N_2414,N_2563);
xnor U2796 (N_2796,N_2434,N_2495);
xor U2797 (N_2797,N_2511,N_2591);
nor U2798 (N_2798,N_2533,N_2425);
nor U2799 (N_2799,N_2567,N_2577);
nor U2800 (N_2800,N_2654,N_2673);
nor U2801 (N_2801,N_2604,N_2773);
nor U2802 (N_2802,N_2707,N_2767);
nor U2803 (N_2803,N_2786,N_2632);
nand U2804 (N_2804,N_2778,N_2792);
xnor U2805 (N_2805,N_2657,N_2629);
nand U2806 (N_2806,N_2749,N_2603);
nor U2807 (N_2807,N_2753,N_2710);
xor U2808 (N_2808,N_2759,N_2745);
nand U2809 (N_2809,N_2634,N_2631);
xnor U2810 (N_2810,N_2601,N_2765);
nand U2811 (N_2811,N_2690,N_2635);
nand U2812 (N_2812,N_2656,N_2639);
nor U2813 (N_2813,N_2748,N_2770);
and U2814 (N_2814,N_2682,N_2734);
and U2815 (N_2815,N_2642,N_2691);
xor U2816 (N_2816,N_2703,N_2640);
nor U2817 (N_2817,N_2617,N_2645);
nor U2818 (N_2818,N_2660,N_2780);
nor U2819 (N_2819,N_2696,N_2731);
or U2820 (N_2820,N_2714,N_2769);
or U2821 (N_2821,N_2671,N_2764);
nor U2822 (N_2822,N_2685,N_2641);
nand U2823 (N_2823,N_2698,N_2791);
nor U2824 (N_2824,N_2697,N_2782);
and U2825 (N_2825,N_2742,N_2646);
and U2826 (N_2826,N_2775,N_2721);
nor U2827 (N_2827,N_2716,N_2612);
xnor U2828 (N_2828,N_2738,N_2677);
and U2829 (N_2829,N_2608,N_2679);
nor U2830 (N_2830,N_2616,N_2625);
or U2831 (N_2831,N_2665,N_2674);
nor U2832 (N_2832,N_2711,N_2638);
nor U2833 (N_2833,N_2757,N_2722);
and U2834 (N_2834,N_2649,N_2650);
or U2835 (N_2835,N_2672,N_2626);
or U2836 (N_2836,N_2662,N_2676);
nand U2837 (N_2837,N_2720,N_2723);
and U2838 (N_2838,N_2797,N_2655);
nor U2839 (N_2839,N_2648,N_2746);
and U2840 (N_2840,N_2725,N_2661);
and U2841 (N_2841,N_2663,N_2693);
nand U2842 (N_2842,N_2796,N_2686);
or U2843 (N_2843,N_2763,N_2614);
and U2844 (N_2844,N_2669,N_2605);
nand U2845 (N_2845,N_2618,N_2607);
nor U2846 (N_2846,N_2728,N_2613);
xor U2847 (N_2847,N_2666,N_2718);
xnor U2848 (N_2848,N_2730,N_2623);
or U2849 (N_2849,N_2627,N_2611);
or U2850 (N_2850,N_2799,N_2622);
nor U2851 (N_2851,N_2702,N_2606);
and U2852 (N_2852,N_2705,N_2790);
or U2853 (N_2853,N_2701,N_2699);
or U2854 (N_2854,N_2761,N_2647);
nand U2855 (N_2855,N_2681,N_2704);
nor U2856 (N_2856,N_2740,N_2772);
nor U2857 (N_2857,N_2758,N_2785);
xnor U2858 (N_2858,N_2793,N_2755);
nand U2859 (N_2859,N_2788,N_2624);
and U2860 (N_2860,N_2658,N_2692);
xor U2861 (N_2861,N_2715,N_2610);
and U2862 (N_2862,N_2687,N_2651);
xnor U2863 (N_2863,N_2644,N_2779);
or U2864 (N_2864,N_2736,N_2615);
or U2865 (N_2865,N_2621,N_2694);
xnor U2866 (N_2866,N_2771,N_2652);
and U2867 (N_2867,N_2795,N_2678);
nor U2868 (N_2868,N_2768,N_2751);
nand U2869 (N_2869,N_2739,N_2643);
xor U2870 (N_2870,N_2600,N_2668);
xor U2871 (N_2871,N_2619,N_2675);
nor U2872 (N_2872,N_2719,N_2709);
or U2873 (N_2873,N_2774,N_2752);
nand U2874 (N_2874,N_2787,N_2750);
and U2875 (N_2875,N_2637,N_2733);
xor U2876 (N_2876,N_2688,N_2747);
nor U2877 (N_2877,N_2781,N_2762);
nor U2878 (N_2878,N_2717,N_2680);
xor U2879 (N_2879,N_2737,N_2602);
nor U2880 (N_2880,N_2609,N_2784);
and U2881 (N_2881,N_2630,N_2798);
or U2882 (N_2882,N_2756,N_2713);
xor U2883 (N_2883,N_2744,N_2794);
nand U2884 (N_2884,N_2743,N_2729);
nor U2885 (N_2885,N_2776,N_2724);
xnor U2886 (N_2886,N_2783,N_2712);
nand U2887 (N_2887,N_2628,N_2735);
and U2888 (N_2888,N_2706,N_2741);
and U2889 (N_2889,N_2695,N_2653);
and U2890 (N_2890,N_2633,N_2777);
or U2891 (N_2891,N_2689,N_2659);
nand U2892 (N_2892,N_2766,N_2684);
nand U2893 (N_2893,N_2620,N_2727);
nor U2894 (N_2894,N_2664,N_2700);
nor U2895 (N_2895,N_2683,N_2760);
nor U2896 (N_2896,N_2636,N_2732);
and U2897 (N_2897,N_2726,N_2667);
nand U2898 (N_2898,N_2670,N_2789);
xnor U2899 (N_2899,N_2708,N_2754);
and U2900 (N_2900,N_2743,N_2774);
nor U2901 (N_2901,N_2761,N_2681);
or U2902 (N_2902,N_2798,N_2656);
nor U2903 (N_2903,N_2754,N_2793);
xnor U2904 (N_2904,N_2795,N_2661);
nor U2905 (N_2905,N_2761,N_2682);
nor U2906 (N_2906,N_2628,N_2741);
and U2907 (N_2907,N_2751,N_2709);
nand U2908 (N_2908,N_2781,N_2618);
and U2909 (N_2909,N_2757,N_2666);
nand U2910 (N_2910,N_2698,N_2735);
xnor U2911 (N_2911,N_2612,N_2722);
nand U2912 (N_2912,N_2749,N_2714);
nand U2913 (N_2913,N_2626,N_2682);
nand U2914 (N_2914,N_2786,N_2648);
nand U2915 (N_2915,N_2763,N_2736);
and U2916 (N_2916,N_2780,N_2772);
nor U2917 (N_2917,N_2639,N_2723);
xnor U2918 (N_2918,N_2617,N_2763);
or U2919 (N_2919,N_2714,N_2737);
nor U2920 (N_2920,N_2628,N_2607);
nand U2921 (N_2921,N_2637,N_2627);
nand U2922 (N_2922,N_2708,N_2737);
xor U2923 (N_2923,N_2664,N_2723);
or U2924 (N_2924,N_2621,N_2698);
and U2925 (N_2925,N_2799,N_2777);
nor U2926 (N_2926,N_2790,N_2627);
or U2927 (N_2927,N_2681,N_2780);
nand U2928 (N_2928,N_2644,N_2788);
or U2929 (N_2929,N_2692,N_2619);
xor U2930 (N_2930,N_2761,N_2694);
nor U2931 (N_2931,N_2636,N_2658);
xnor U2932 (N_2932,N_2625,N_2786);
and U2933 (N_2933,N_2680,N_2637);
or U2934 (N_2934,N_2787,N_2757);
nand U2935 (N_2935,N_2672,N_2652);
xor U2936 (N_2936,N_2675,N_2652);
xnor U2937 (N_2937,N_2732,N_2705);
nand U2938 (N_2938,N_2671,N_2649);
or U2939 (N_2939,N_2644,N_2730);
or U2940 (N_2940,N_2775,N_2785);
nor U2941 (N_2941,N_2742,N_2708);
xor U2942 (N_2942,N_2749,N_2716);
or U2943 (N_2943,N_2653,N_2680);
xnor U2944 (N_2944,N_2762,N_2706);
xor U2945 (N_2945,N_2654,N_2691);
nor U2946 (N_2946,N_2644,N_2637);
and U2947 (N_2947,N_2725,N_2677);
xnor U2948 (N_2948,N_2761,N_2612);
xor U2949 (N_2949,N_2625,N_2622);
or U2950 (N_2950,N_2660,N_2619);
nand U2951 (N_2951,N_2697,N_2671);
or U2952 (N_2952,N_2772,N_2613);
xor U2953 (N_2953,N_2787,N_2659);
and U2954 (N_2954,N_2729,N_2768);
xor U2955 (N_2955,N_2729,N_2660);
nor U2956 (N_2956,N_2742,N_2603);
nand U2957 (N_2957,N_2637,N_2736);
nor U2958 (N_2958,N_2746,N_2706);
or U2959 (N_2959,N_2754,N_2631);
nand U2960 (N_2960,N_2676,N_2661);
xnor U2961 (N_2961,N_2643,N_2676);
nor U2962 (N_2962,N_2778,N_2742);
or U2963 (N_2963,N_2760,N_2770);
nor U2964 (N_2964,N_2642,N_2700);
nor U2965 (N_2965,N_2731,N_2635);
nand U2966 (N_2966,N_2649,N_2652);
and U2967 (N_2967,N_2693,N_2653);
and U2968 (N_2968,N_2653,N_2752);
and U2969 (N_2969,N_2611,N_2790);
xor U2970 (N_2970,N_2722,N_2683);
nor U2971 (N_2971,N_2683,N_2689);
or U2972 (N_2972,N_2707,N_2755);
or U2973 (N_2973,N_2731,N_2721);
and U2974 (N_2974,N_2748,N_2669);
xor U2975 (N_2975,N_2769,N_2708);
nor U2976 (N_2976,N_2776,N_2632);
or U2977 (N_2977,N_2722,N_2666);
xor U2978 (N_2978,N_2747,N_2686);
xor U2979 (N_2979,N_2636,N_2708);
or U2980 (N_2980,N_2750,N_2636);
nand U2981 (N_2981,N_2701,N_2787);
or U2982 (N_2982,N_2732,N_2767);
and U2983 (N_2983,N_2700,N_2759);
and U2984 (N_2984,N_2636,N_2763);
and U2985 (N_2985,N_2639,N_2749);
xnor U2986 (N_2986,N_2605,N_2600);
nand U2987 (N_2987,N_2725,N_2706);
and U2988 (N_2988,N_2706,N_2635);
nor U2989 (N_2989,N_2743,N_2797);
nand U2990 (N_2990,N_2633,N_2797);
and U2991 (N_2991,N_2705,N_2653);
and U2992 (N_2992,N_2605,N_2702);
nand U2993 (N_2993,N_2683,N_2658);
nor U2994 (N_2994,N_2799,N_2612);
and U2995 (N_2995,N_2665,N_2688);
and U2996 (N_2996,N_2644,N_2700);
nor U2997 (N_2997,N_2638,N_2768);
xnor U2998 (N_2998,N_2692,N_2758);
nor U2999 (N_2999,N_2672,N_2685);
and U3000 (N_3000,N_2936,N_2963);
and U3001 (N_3001,N_2983,N_2915);
and U3002 (N_3002,N_2951,N_2985);
and U3003 (N_3003,N_2855,N_2834);
nor U3004 (N_3004,N_2836,N_2984);
nand U3005 (N_3005,N_2952,N_2959);
or U3006 (N_3006,N_2989,N_2816);
and U3007 (N_3007,N_2998,N_2870);
and U3008 (N_3008,N_2886,N_2958);
nor U3009 (N_3009,N_2923,N_2882);
nor U3010 (N_3010,N_2953,N_2843);
and U3011 (N_3011,N_2960,N_2949);
nor U3012 (N_3012,N_2817,N_2954);
nor U3013 (N_3013,N_2999,N_2971);
and U3014 (N_3014,N_2838,N_2916);
nor U3015 (N_3015,N_2890,N_2864);
nor U3016 (N_3016,N_2909,N_2903);
nand U3017 (N_3017,N_2850,N_2905);
xnor U3018 (N_3018,N_2866,N_2868);
or U3019 (N_3019,N_2941,N_2848);
and U3020 (N_3020,N_2815,N_2993);
or U3021 (N_3021,N_2986,N_2940);
xor U3022 (N_3022,N_2837,N_2825);
nor U3023 (N_3023,N_2947,N_2877);
nor U3024 (N_3024,N_2853,N_2884);
or U3025 (N_3025,N_2921,N_2812);
nor U3026 (N_3026,N_2946,N_2926);
xnor U3027 (N_3027,N_2930,N_2803);
xor U3028 (N_3028,N_2874,N_2879);
nand U3029 (N_3029,N_2867,N_2965);
xor U3030 (N_3030,N_2906,N_2974);
nand U3031 (N_3031,N_2865,N_2944);
nor U3032 (N_3032,N_2831,N_2811);
nor U3033 (N_3033,N_2939,N_2937);
and U3034 (N_3034,N_2943,N_2980);
xnor U3035 (N_3035,N_2829,N_2847);
xnor U3036 (N_3036,N_2804,N_2988);
and U3037 (N_3037,N_2822,N_2977);
or U3038 (N_3038,N_2917,N_2854);
xnor U3039 (N_3039,N_2970,N_2826);
or U3040 (N_3040,N_2919,N_2852);
xnor U3041 (N_3041,N_2885,N_2914);
xnor U3042 (N_3042,N_2860,N_2912);
nor U3043 (N_3043,N_2844,N_2895);
and U3044 (N_3044,N_2927,N_2821);
and U3045 (N_3045,N_2918,N_2904);
nor U3046 (N_3046,N_2840,N_2839);
and U3047 (N_3047,N_2898,N_2932);
or U3048 (N_3048,N_2934,N_2966);
and U3049 (N_3049,N_2888,N_2832);
nor U3050 (N_3050,N_2935,N_2880);
or U3051 (N_3051,N_2842,N_2819);
nand U3052 (N_3052,N_2964,N_2992);
and U3053 (N_3053,N_2911,N_2828);
xor U3054 (N_3054,N_2810,N_2979);
xnor U3055 (N_3055,N_2814,N_2857);
xnor U3056 (N_3056,N_2813,N_2929);
or U3057 (N_3057,N_2994,N_2807);
nor U3058 (N_3058,N_2861,N_2872);
xnor U3059 (N_3059,N_2887,N_2823);
xnor U3060 (N_3060,N_2871,N_2875);
and U3061 (N_3061,N_2801,N_2824);
and U3062 (N_3062,N_2925,N_2878);
nand U3063 (N_3063,N_2968,N_2869);
nand U3064 (N_3064,N_2893,N_2802);
xor U3065 (N_3065,N_2995,N_2990);
nand U3066 (N_3066,N_2891,N_2902);
and U3067 (N_3067,N_2800,N_2962);
xnor U3068 (N_3068,N_2883,N_2806);
and U3069 (N_3069,N_2851,N_2928);
nand U3070 (N_3070,N_2830,N_2862);
nor U3071 (N_3071,N_2938,N_2901);
and U3072 (N_3072,N_2910,N_2973);
and U3073 (N_3073,N_2845,N_2863);
or U3074 (N_3074,N_2924,N_2897);
nand U3075 (N_3075,N_2835,N_2913);
and U3076 (N_3076,N_2894,N_2987);
nand U3077 (N_3077,N_2881,N_2849);
nand U3078 (N_3078,N_2945,N_2975);
and U3079 (N_3079,N_2833,N_2859);
or U3080 (N_3080,N_2873,N_2955);
and U3081 (N_3081,N_2931,N_2972);
and U3082 (N_3082,N_2889,N_2996);
nor U3083 (N_3083,N_2808,N_2856);
nand U3084 (N_3084,N_2818,N_2991);
or U3085 (N_3085,N_2827,N_2933);
or U3086 (N_3086,N_2896,N_2997);
and U3087 (N_3087,N_2981,N_2908);
nor U3088 (N_3088,N_2978,N_2942);
xor U3089 (N_3089,N_2920,N_2892);
xor U3090 (N_3090,N_2820,N_2846);
xor U3091 (N_3091,N_2876,N_2841);
or U3092 (N_3092,N_2809,N_2956);
nand U3093 (N_3093,N_2969,N_2982);
and U3094 (N_3094,N_2805,N_2961);
xor U3095 (N_3095,N_2967,N_2922);
xnor U3096 (N_3096,N_2950,N_2858);
or U3097 (N_3097,N_2907,N_2948);
nor U3098 (N_3098,N_2957,N_2976);
nand U3099 (N_3099,N_2900,N_2899);
or U3100 (N_3100,N_2851,N_2802);
xor U3101 (N_3101,N_2920,N_2870);
nor U3102 (N_3102,N_2823,N_2811);
nand U3103 (N_3103,N_2935,N_2800);
or U3104 (N_3104,N_2819,N_2979);
and U3105 (N_3105,N_2887,N_2894);
nand U3106 (N_3106,N_2945,N_2863);
xor U3107 (N_3107,N_2917,N_2820);
and U3108 (N_3108,N_2825,N_2829);
xnor U3109 (N_3109,N_2957,N_2994);
or U3110 (N_3110,N_2886,N_2861);
or U3111 (N_3111,N_2908,N_2848);
and U3112 (N_3112,N_2913,N_2865);
xor U3113 (N_3113,N_2943,N_2903);
nand U3114 (N_3114,N_2880,N_2890);
xor U3115 (N_3115,N_2887,N_2969);
xnor U3116 (N_3116,N_2865,N_2863);
nand U3117 (N_3117,N_2816,N_2869);
nor U3118 (N_3118,N_2916,N_2917);
or U3119 (N_3119,N_2819,N_2912);
or U3120 (N_3120,N_2872,N_2838);
nand U3121 (N_3121,N_2808,N_2882);
or U3122 (N_3122,N_2956,N_2832);
xor U3123 (N_3123,N_2942,N_2946);
and U3124 (N_3124,N_2815,N_2891);
and U3125 (N_3125,N_2883,N_2936);
xnor U3126 (N_3126,N_2884,N_2815);
xnor U3127 (N_3127,N_2955,N_2856);
or U3128 (N_3128,N_2967,N_2833);
nor U3129 (N_3129,N_2815,N_2892);
or U3130 (N_3130,N_2905,N_2803);
nand U3131 (N_3131,N_2973,N_2945);
nand U3132 (N_3132,N_2999,N_2842);
or U3133 (N_3133,N_2850,N_2967);
and U3134 (N_3134,N_2998,N_2899);
or U3135 (N_3135,N_2992,N_2975);
or U3136 (N_3136,N_2971,N_2973);
and U3137 (N_3137,N_2923,N_2965);
and U3138 (N_3138,N_2935,N_2804);
nor U3139 (N_3139,N_2991,N_2808);
or U3140 (N_3140,N_2874,N_2886);
nor U3141 (N_3141,N_2978,N_2915);
xor U3142 (N_3142,N_2948,N_2810);
nor U3143 (N_3143,N_2842,N_2970);
and U3144 (N_3144,N_2865,N_2809);
and U3145 (N_3145,N_2918,N_2937);
nor U3146 (N_3146,N_2915,N_2883);
nor U3147 (N_3147,N_2844,N_2805);
or U3148 (N_3148,N_2975,N_2929);
nor U3149 (N_3149,N_2918,N_2897);
nand U3150 (N_3150,N_2968,N_2931);
xor U3151 (N_3151,N_2977,N_2864);
and U3152 (N_3152,N_2858,N_2983);
nor U3153 (N_3153,N_2913,N_2836);
or U3154 (N_3154,N_2938,N_2886);
nand U3155 (N_3155,N_2946,N_2801);
nand U3156 (N_3156,N_2990,N_2994);
nor U3157 (N_3157,N_2888,N_2993);
nor U3158 (N_3158,N_2966,N_2940);
nor U3159 (N_3159,N_2963,N_2812);
xor U3160 (N_3160,N_2951,N_2888);
nor U3161 (N_3161,N_2988,N_2866);
nand U3162 (N_3162,N_2816,N_2904);
nand U3163 (N_3163,N_2843,N_2865);
and U3164 (N_3164,N_2889,N_2937);
and U3165 (N_3165,N_2884,N_2914);
nand U3166 (N_3166,N_2894,N_2880);
xor U3167 (N_3167,N_2909,N_2885);
nor U3168 (N_3168,N_2840,N_2957);
xor U3169 (N_3169,N_2984,N_2866);
nand U3170 (N_3170,N_2957,N_2956);
nand U3171 (N_3171,N_2923,N_2822);
nand U3172 (N_3172,N_2847,N_2864);
nor U3173 (N_3173,N_2937,N_2829);
nand U3174 (N_3174,N_2811,N_2913);
nand U3175 (N_3175,N_2887,N_2824);
xor U3176 (N_3176,N_2977,N_2919);
xnor U3177 (N_3177,N_2976,N_2994);
or U3178 (N_3178,N_2956,N_2933);
xnor U3179 (N_3179,N_2872,N_2832);
or U3180 (N_3180,N_2880,N_2924);
nand U3181 (N_3181,N_2819,N_2938);
nor U3182 (N_3182,N_2981,N_2919);
and U3183 (N_3183,N_2941,N_2842);
nand U3184 (N_3184,N_2801,N_2947);
nor U3185 (N_3185,N_2895,N_2931);
nand U3186 (N_3186,N_2977,N_2955);
or U3187 (N_3187,N_2984,N_2845);
nand U3188 (N_3188,N_2899,N_2816);
xnor U3189 (N_3189,N_2859,N_2865);
nand U3190 (N_3190,N_2983,N_2998);
or U3191 (N_3191,N_2838,N_2905);
nand U3192 (N_3192,N_2950,N_2961);
xnor U3193 (N_3193,N_2805,N_2841);
nor U3194 (N_3194,N_2978,N_2906);
nand U3195 (N_3195,N_2975,N_2915);
or U3196 (N_3196,N_2969,N_2828);
and U3197 (N_3197,N_2947,N_2894);
xor U3198 (N_3198,N_2948,N_2956);
xor U3199 (N_3199,N_2898,N_2918);
and U3200 (N_3200,N_3155,N_3042);
xnor U3201 (N_3201,N_3021,N_3120);
or U3202 (N_3202,N_3002,N_3132);
and U3203 (N_3203,N_3057,N_3008);
nand U3204 (N_3204,N_3007,N_3195);
or U3205 (N_3205,N_3036,N_3037);
nand U3206 (N_3206,N_3016,N_3183);
or U3207 (N_3207,N_3006,N_3158);
xnor U3208 (N_3208,N_3129,N_3173);
and U3209 (N_3209,N_3093,N_3117);
xnor U3210 (N_3210,N_3064,N_3051);
nor U3211 (N_3211,N_3177,N_3055);
and U3212 (N_3212,N_3065,N_3060);
nor U3213 (N_3213,N_3154,N_3044);
and U3214 (N_3214,N_3098,N_3130);
and U3215 (N_3215,N_3199,N_3184);
xnor U3216 (N_3216,N_3135,N_3086);
nand U3217 (N_3217,N_3147,N_3152);
or U3218 (N_3218,N_3189,N_3041);
nand U3219 (N_3219,N_3115,N_3077);
nor U3220 (N_3220,N_3102,N_3197);
nor U3221 (N_3221,N_3112,N_3190);
xnor U3222 (N_3222,N_3046,N_3092);
xnor U3223 (N_3223,N_3123,N_3069);
xor U3224 (N_3224,N_3048,N_3164);
xnor U3225 (N_3225,N_3103,N_3150);
nor U3226 (N_3226,N_3104,N_3076);
xor U3227 (N_3227,N_3000,N_3003);
xor U3228 (N_3228,N_3078,N_3031);
xnor U3229 (N_3229,N_3089,N_3027);
nor U3230 (N_3230,N_3028,N_3185);
nand U3231 (N_3231,N_3105,N_3043);
and U3232 (N_3232,N_3163,N_3083);
or U3233 (N_3233,N_3179,N_3140);
and U3234 (N_3234,N_3080,N_3038);
xor U3235 (N_3235,N_3106,N_3128);
nor U3236 (N_3236,N_3013,N_3188);
xnor U3237 (N_3237,N_3171,N_3127);
nor U3238 (N_3238,N_3153,N_3099);
nor U3239 (N_3239,N_3066,N_3018);
or U3240 (N_3240,N_3012,N_3005);
nor U3241 (N_3241,N_3101,N_3170);
and U3242 (N_3242,N_3125,N_3111);
nor U3243 (N_3243,N_3119,N_3191);
and U3244 (N_3244,N_3095,N_3108);
nor U3245 (N_3245,N_3025,N_3161);
or U3246 (N_3246,N_3059,N_3074);
or U3247 (N_3247,N_3126,N_3040);
xnor U3248 (N_3248,N_3157,N_3050);
or U3249 (N_3249,N_3035,N_3091);
nor U3250 (N_3250,N_3151,N_3159);
and U3251 (N_3251,N_3133,N_3193);
and U3252 (N_3252,N_3107,N_3121);
and U3253 (N_3253,N_3049,N_3146);
nor U3254 (N_3254,N_3010,N_3024);
nand U3255 (N_3255,N_3052,N_3033);
xor U3256 (N_3256,N_3124,N_3196);
or U3257 (N_3257,N_3100,N_3187);
or U3258 (N_3258,N_3139,N_3058);
and U3259 (N_3259,N_3053,N_3081);
nand U3260 (N_3260,N_3014,N_3096);
nor U3261 (N_3261,N_3067,N_3165);
nor U3262 (N_3262,N_3145,N_3166);
and U3263 (N_3263,N_3039,N_3090);
xnor U3264 (N_3264,N_3180,N_3172);
or U3265 (N_3265,N_3182,N_3017);
xnor U3266 (N_3266,N_3148,N_3088);
and U3267 (N_3267,N_3068,N_3030);
and U3268 (N_3268,N_3032,N_3192);
xor U3269 (N_3269,N_3174,N_3168);
or U3270 (N_3270,N_3045,N_3142);
nor U3271 (N_3271,N_3019,N_3063);
or U3272 (N_3272,N_3056,N_3156);
xnor U3273 (N_3273,N_3079,N_3072);
and U3274 (N_3274,N_3162,N_3116);
or U3275 (N_3275,N_3073,N_3181);
nand U3276 (N_3276,N_3149,N_3061);
nand U3277 (N_3277,N_3023,N_3137);
or U3278 (N_3278,N_3175,N_3097);
nand U3279 (N_3279,N_3131,N_3198);
nand U3280 (N_3280,N_3122,N_3082);
xor U3281 (N_3281,N_3084,N_3009);
or U3282 (N_3282,N_3160,N_3071);
nor U3283 (N_3283,N_3194,N_3169);
nand U3284 (N_3284,N_3178,N_3136);
nand U3285 (N_3285,N_3029,N_3113);
and U3286 (N_3286,N_3026,N_3004);
and U3287 (N_3287,N_3094,N_3047);
nor U3288 (N_3288,N_3176,N_3186);
or U3289 (N_3289,N_3034,N_3022);
nor U3290 (N_3290,N_3110,N_3011);
or U3291 (N_3291,N_3015,N_3144);
or U3292 (N_3292,N_3001,N_3020);
xor U3293 (N_3293,N_3167,N_3075);
or U3294 (N_3294,N_3062,N_3109);
or U3295 (N_3295,N_3143,N_3054);
or U3296 (N_3296,N_3085,N_3138);
nand U3297 (N_3297,N_3070,N_3118);
or U3298 (N_3298,N_3087,N_3141);
nand U3299 (N_3299,N_3134,N_3114);
and U3300 (N_3300,N_3067,N_3179);
nor U3301 (N_3301,N_3031,N_3033);
and U3302 (N_3302,N_3141,N_3057);
xor U3303 (N_3303,N_3012,N_3170);
nor U3304 (N_3304,N_3134,N_3026);
or U3305 (N_3305,N_3140,N_3049);
xnor U3306 (N_3306,N_3094,N_3012);
or U3307 (N_3307,N_3016,N_3010);
nand U3308 (N_3308,N_3198,N_3123);
xnor U3309 (N_3309,N_3129,N_3098);
nand U3310 (N_3310,N_3194,N_3187);
and U3311 (N_3311,N_3076,N_3138);
nand U3312 (N_3312,N_3107,N_3034);
xnor U3313 (N_3313,N_3086,N_3039);
nand U3314 (N_3314,N_3005,N_3113);
xor U3315 (N_3315,N_3149,N_3160);
and U3316 (N_3316,N_3119,N_3175);
xor U3317 (N_3317,N_3170,N_3073);
nor U3318 (N_3318,N_3012,N_3172);
xor U3319 (N_3319,N_3049,N_3154);
xnor U3320 (N_3320,N_3191,N_3006);
xor U3321 (N_3321,N_3050,N_3021);
or U3322 (N_3322,N_3004,N_3146);
and U3323 (N_3323,N_3138,N_3181);
and U3324 (N_3324,N_3127,N_3151);
xor U3325 (N_3325,N_3054,N_3126);
nand U3326 (N_3326,N_3084,N_3057);
xor U3327 (N_3327,N_3082,N_3158);
xor U3328 (N_3328,N_3126,N_3175);
nand U3329 (N_3329,N_3121,N_3172);
xnor U3330 (N_3330,N_3011,N_3157);
nand U3331 (N_3331,N_3099,N_3136);
and U3332 (N_3332,N_3027,N_3185);
and U3333 (N_3333,N_3055,N_3188);
and U3334 (N_3334,N_3045,N_3069);
xor U3335 (N_3335,N_3065,N_3017);
nand U3336 (N_3336,N_3027,N_3031);
or U3337 (N_3337,N_3047,N_3087);
nor U3338 (N_3338,N_3081,N_3003);
xor U3339 (N_3339,N_3030,N_3042);
and U3340 (N_3340,N_3174,N_3089);
and U3341 (N_3341,N_3008,N_3175);
or U3342 (N_3342,N_3060,N_3073);
nand U3343 (N_3343,N_3077,N_3136);
nor U3344 (N_3344,N_3143,N_3059);
xnor U3345 (N_3345,N_3030,N_3166);
and U3346 (N_3346,N_3121,N_3108);
nand U3347 (N_3347,N_3070,N_3005);
xor U3348 (N_3348,N_3073,N_3103);
or U3349 (N_3349,N_3164,N_3037);
nand U3350 (N_3350,N_3058,N_3024);
xor U3351 (N_3351,N_3111,N_3192);
nor U3352 (N_3352,N_3016,N_3090);
xor U3353 (N_3353,N_3026,N_3096);
nand U3354 (N_3354,N_3046,N_3156);
nor U3355 (N_3355,N_3134,N_3083);
nand U3356 (N_3356,N_3110,N_3023);
nor U3357 (N_3357,N_3089,N_3044);
and U3358 (N_3358,N_3149,N_3113);
or U3359 (N_3359,N_3122,N_3003);
or U3360 (N_3360,N_3078,N_3056);
and U3361 (N_3361,N_3172,N_3199);
xnor U3362 (N_3362,N_3068,N_3152);
nand U3363 (N_3363,N_3150,N_3135);
xnor U3364 (N_3364,N_3080,N_3168);
and U3365 (N_3365,N_3128,N_3022);
and U3366 (N_3366,N_3095,N_3198);
nand U3367 (N_3367,N_3019,N_3107);
and U3368 (N_3368,N_3108,N_3072);
nor U3369 (N_3369,N_3090,N_3026);
and U3370 (N_3370,N_3070,N_3039);
xor U3371 (N_3371,N_3053,N_3185);
xor U3372 (N_3372,N_3181,N_3147);
nor U3373 (N_3373,N_3089,N_3179);
nand U3374 (N_3374,N_3050,N_3094);
or U3375 (N_3375,N_3138,N_3013);
xor U3376 (N_3376,N_3176,N_3141);
or U3377 (N_3377,N_3028,N_3177);
nor U3378 (N_3378,N_3027,N_3005);
xnor U3379 (N_3379,N_3165,N_3090);
or U3380 (N_3380,N_3195,N_3009);
and U3381 (N_3381,N_3174,N_3036);
or U3382 (N_3382,N_3039,N_3083);
or U3383 (N_3383,N_3068,N_3169);
and U3384 (N_3384,N_3172,N_3068);
nor U3385 (N_3385,N_3091,N_3164);
and U3386 (N_3386,N_3115,N_3007);
nand U3387 (N_3387,N_3133,N_3180);
xnor U3388 (N_3388,N_3061,N_3153);
nor U3389 (N_3389,N_3002,N_3090);
or U3390 (N_3390,N_3177,N_3052);
or U3391 (N_3391,N_3087,N_3110);
xor U3392 (N_3392,N_3160,N_3027);
nand U3393 (N_3393,N_3125,N_3042);
xor U3394 (N_3394,N_3043,N_3074);
or U3395 (N_3395,N_3041,N_3181);
and U3396 (N_3396,N_3058,N_3102);
xor U3397 (N_3397,N_3067,N_3114);
nor U3398 (N_3398,N_3077,N_3193);
nand U3399 (N_3399,N_3177,N_3063);
nand U3400 (N_3400,N_3368,N_3321);
nor U3401 (N_3401,N_3253,N_3353);
nor U3402 (N_3402,N_3394,N_3320);
nand U3403 (N_3403,N_3285,N_3331);
or U3404 (N_3404,N_3216,N_3206);
and U3405 (N_3405,N_3210,N_3395);
nand U3406 (N_3406,N_3278,N_3208);
nand U3407 (N_3407,N_3242,N_3222);
and U3408 (N_3408,N_3270,N_3301);
nor U3409 (N_3409,N_3305,N_3243);
and U3410 (N_3410,N_3289,N_3207);
or U3411 (N_3411,N_3311,N_3217);
and U3412 (N_3412,N_3239,N_3269);
or U3413 (N_3413,N_3310,N_3323);
nand U3414 (N_3414,N_3354,N_3360);
or U3415 (N_3415,N_3218,N_3226);
xor U3416 (N_3416,N_3380,N_3202);
nor U3417 (N_3417,N_3369,N_3225);
nand U3418 (N_3418,N_3357,N_3229);
and U3419 (N_3419,N_3374,N_3215);
xor U3420 (N_3420,N_3251,N_3336);
nor U3421 (N_3421,N_3297,N_3386);
or U3422 (N_3422,N_3306,N_3355);
nand U3423 (N_3423,N_3389,N_3340);
and U3424 (N_3424,N_3303,N_3378);
nand U3425 (N_3425,N_3308,N_3393);
nor U3426 (N_3426,N_3344,N_3284);
or U3427 (N_3427,N_3256,N_3347);
nor U3428 (N_3428,N_3282,N_3281);
nand U3429 (N_3429,N_3261,N_3268);
nor U3430 (N_3430,N_3304,N_3223);
or U3431 (N_3431,N_3376,N_3232);
xor U3432 (N_3432,N_3315,N_3264);
xor U3433 (N_3433,N_3392,N_3377);
nand U3434 (N_3434,N_3287,N_3341);
or U3435 (N_3435,N_3237,N_3205);
nand U3436 (N_3436,N_3338,N_3324);
and U3437 (N_3437,N_3348,N_3384);
or U3438 (N_3438,N_3335,N_3367);
xnor U3439 (N_3439,N_3312,N_3258);
and U3440 (N_3440,N_3337,N_3220);
and U3441 (N_3441,N_3313,N_3212);
or U3442 (N_3442,N_3352,N_3290);
nor U3443 (N_3443,N_3292,N_3314);
and U3444 (N_3444,N_3273,N_3288);
xnor U3445 (N_3445,N_3234,N_3398);
and U3446 (N_3446,N_3356,N_3241);
nand U3447 (N_3447,N_3366,N_3265);
or U3448 (N_3448,N_3370,N_3209);
and U3449 (N_3449,N_3309,N_3257);
xor U3450 (N_3450,N_3280,N_3249);
xnor U3451 (N_3451,N_3294,N_3224);
nor U3452 (N_3452,N_3327,N_3245);
nand U3453 (N_3453,N_3244,N_3221);
nor U3454 (N_3454,N_3351,N_3399);
and U3455 (N_3455,N_3339,N_3277);
nor U3456 (N_3456,N_3373,N_3259);
or U3457 (N_3457,N_3300,N_3298);
xnor U3458 (N_3458,N_3260,N_3214);
nand U3459 (N_3459,N_3295,N_3391);
or U3460 (N_3460,N_3385,N_3302);
nor U3461 (N_3461,N_3322,N_3211);
xnor U3462 (N_3462,N_3365,N_3274);
nor U3463 (N_3463,N_3203,N_3263);
nor U3464 (N_3464,N_3200,N_3272);
or U3465 (N_3465,N_3255,N_3387);
nor U3466 (N_3466,N_3227,N_3271);
nor U3467 (N_3467,N_3230,N_3228);
and U3468 (N_3468,N_3250,N_3262);
xnor U3469 (N_3469,N_3213,N_3329);
or U3470 (N_3470,N_3396,N_3361);
nand U3471 (N_3471,N_3316,N_3364);
nor U3472 (N_3472,N_3388,N_3350);
xor U3473 (N_3473,N_3359,N_3345);
or U3474 (N_3474,N_3296,N_3231);
nand U3475 (N_3475,N_3346,N_3201);
and U3476 (N_3476,N_3283,N_3236);
and U3477 (N_3477,N_3375,N_3238);
xnor U3478 (N_3478,N_3252,N_3343);
nand U3479 (N_3479,N_3247,N_3248);
xor U3480 (N_3480,N_3318,N_3240);
nand U3481 (N_3481,N_3319,N_3390);
or U3482 (N_3482,N_3235,N_3382);
or U3483 (N_3483,N_3293,N_3333);
nor U3484 (N_3484,N_3371,N_3381);
xnor U3485 (N_3485,N_3342,N_3307);
and U3486 (N_3486,N_3349,N_3363);
and U3487 (N_3487,N_3266,N_3267);
nand U3488 (N_3488,N_3254,N_3286);
xor U3489 (N_3489,N_3330,N_3279);
or U3490 (N_3490,N_3317,N_3358);
or U3491 (N_3491,N_3334,N_3275);
nand U3492 (N_3492,N_3332,N_3299);
or U3493 (N_3493,N_3276,N_3362);
xor U3494 (N_3494,N_3379,N_3372);
nand U3495 (N_3495,N_3383,N_3328);
xnor U3496 (N_3496,N_3246,N_3325);
or U3497 (N_3497,N_3219,N_3233);
or U3498 (N_3498,N_3397,N_3326);
nand U3499 (N_3499,N_3204,N_3291);
nand U3500 (N_3500,N_3355,N_3298);
xnor U3501 (N_3501,N_3296,N_3337);
nand U3502 (N_3502,N_3245,N_3207);
or U3503 (N_3503,N_3331,N_3207);
or U3504 (N_3504,N_3248,N_3218);
nand U3505 (N_3505,N_3261,N_3394);
nor U3506 (N_3506,N_3370,N_3285);
nor U3507 (N_3507,N_3390,N_3232);
or U3508 (N_3508,N_3288,N_3291);
xnor U3509 (N_3509,N_3290,N_3307);
xnor U3510 (N_3510,N_3295,N_3372);
nand U3511 (N_3511,N_3217,N_3270);
and U3512 (N_3512,N_3330,N_3393);
nand U3513 (N_3513,N_3205,N_3238);
and U3514 (N_3514,N_3361,N_3273);
xnor U3515 (N_3515,N_3317,N_3237);
nand U3516 (N_3516,N_3385,N_3205);
and U3517 (N_3517,N_3334,N_3279);
nand U3518 (N_3518,N_3299,N_3208);
nand U3519 (N_3519,N_3309,N_3393);
xor U3520 (N_3520,N_3332,N_3286);
nor U3521 (N_3521,N_3358,N_3204);
nor U3522 (N_3522,N_3363,N_3353);
nand U3523 (N_3523,N_3257,N_3345);
nor U3524 (N_3524,N_3386,N_3351);
nor U3525 (N_3525,N_3298,N_3390);
or U3526 (N_3526,N_3344,N_3236);
or U3527 (N_3527,N_3388,N_3206);
and U3528 (N_3528,N_3318,N_3267);
nand U3529 (N_3529,N_3349,N_3206);
and U3530 (N_3530,N_3291,N_3271);
xor U3531 (N_3531,N_3244,N_3235);
or U3532 (N_3532,N_3356,N_3248);
or U3533 (N_3533,N_3279,N_3392);
xor U3534 (N_3534,N_3251,N_3306);
xor U3535 (N_3535,N_3322,N_3342);
nor U3536 (N_3536,N_3274,N_3397);
nand U3537 (N_3537,N_3313,N_3347);
or U3538 (N_3538,N_3259,N_3273);
nand U3539 (N_3539,N_3344,N_3230);
nor U3540 (N_3540,N_3272,N_3380);
or U3541 (N_3541,N_3261,N_3337);
nor U3542 (N_3542,N_3256,N_3309);
xor U3543 (N_3543,N_3233,N_3346);
or U3544 (N_3544,N_3346,N_3322);
and U3545 (N_3545,N_3218,N_3208);
xnor U3546 (N_3546,N_3235,N_3323);
and U3547 (N_3547,N_3393,N_3368);
xnor U3548 (N_3548,N_3298,N_3240);
nand U3549 (N_3549,N_3317,N_3295);
and U3550 (N_3550,N_3276,N_3381);
or U3551 (N_3551,N_3254,N_3270);
nor U3552 (N_3552,N_3282,N_3384);
or U3553 (N_3553,N_3354,N_3356);
xor U3554 (N_3554,N_3234,N_3247);
or U3555 (N_3555,N_3248,N_3362);
nand U3556 (N_3556,N_3272,N_3284);
nor U3557 (N_3557,N_3258,N_3265);
or U3558 (N_3558,N_3267,N_3375);
xor U3559 (N_3559,N_3265,N_3317);
nor U3560 (N_3560,N_3382,N_3368);
nand U3561 (N_3561,N_3331,N_3381);
and U3562 (N_3562,N_3233,N_3258);
nor U3563 (N_3563,N_3230,N_3265);
nor U3564 (N_3564,N_3224,N_3259);
and U3565 (N_3565,N_3348,N_3361);
and U3566 (N_3566,N_3393,N_3224);
xnor U3567 (N_3567,N_3251,N_3327);
or U3568 (N_3568,N_3213,N_3223);
nand U3569 (N_3569,N_3285,N_3264);
nand U3570 (N_3570,N_3298,N_3286);
or U3571 (N_3571,N_3212,N_3257);
xnor U3572 (N_3572,N_3223,N_3284);
xnor U3573 (N_3573,N_3283,N_3241);
or U3574 (N_3574,N_3391,N_3280);
xnor U3575 (N_3575,N_3220,N_3354);
nand U3576 (N_3576,N_3282,N_3334);
nor U3577 (N_3577,N_3376,N_3333);
nand U3578 (N_3578,N_3248,N_3240);
xnor U3579 (N_3579,N_3390,N_3320);
nand U3580 (N_3580,N_3347,N_3281);
or U3581 (N_3581,N_3208,N_3372);
xnor U3582 (N_3582,N_3352,N_3236);
and U3583 (N_3583,N_3307,N_3215);
nor U3584 (N_3584,N_3207,N_3378);
xor U3585 (N_3585,N_3209,N_3268);
and U3586 (N_3586,N_3216,N_3396);
and U3587 (N_3587,N_3293,N_3273);
or U3588 (N_3588,N_3370,N_3264);
or U3589 (N_3589,N_3395,N_3240);
or U3590 (N_3590,N_3315,N_3236);
nand U3591 (N_3591,N_3273,N_3208);
and U3592 (N_3592,N_3384,N_3325);
nand U3593 (N_3593,N_3200,N_3271);
nor U3594 (N_3594,N_3275,N_3279);
xnor U3595 (N_3595,N_3308,N_3373);
nor U3596 (N_3596,N_3342,N_3233);
nor U3597 (N_3597,N_3223,N_3241);
and U3598 (N_3598,N_3251,N_3256);
xnor U3599 (N_3599,N_3303,N_3235);
xor U3600 (N_3600,N_3488,N_3493);
nor U3601 (N_3601,N_3547,N_3563);
nand U3602 (N_3602,N_3500,N_3437);
nor U3603 (N_3603,N_3432,N_3456);
and U3604 (N_3604,N_3404,N_3536);
and U3605 (N_3605,N_3453,N_3573);
or U3606 (N_3606,N_3520,N_3586);
and U3607 (N_3607,N_3485,N_3498);
or U3608 (N_3608,N_3525,N_3414);
and U3609 (N_3609,N_3440,N_3511);
or U3610 (N_3610,N_3489,N_3530);
or U3611 (N_3611,N_3544,N_3447);
or U3612 (N_3612,N_3473,N_3400);
nor U3613 (N_3613,N_3523,N_3477);
nand U3614 (N_3614,N_3581,N_3531);
and U3615 (N_3615,N_3425,N_3492);
and U3616 (N_3616,N_3592,N_3448);
and U3617 (N_3617,N_3574,N_3491);
xor U3618 (N_3618,N_3463,N_3513);
nand U3619 (N_3619,N_3571,N_3518);
nor U3620 (N_3620,N_3416,N_3468);
or U3621 (N_3621,N_3408,N_3593);
xor U3622 (N_3622,N_3564,N_3512);
nand U3623 (N_3623,N_3483,N_3539);
nand U3624 (N_3624,N_3508,N_3555);
nand U3625 (N_3625,N_3522,N_3538);
and U3626 (N_3626,N_3430,N_3553);
nand U3627 (N_3627,N_3598,N_3527);
and U3628 (N_3628,N_3433,N_3550);
xnor U3629 (N_3629,N_3501,N_3517);
nor U3630 (N_3630,N_3509,N_3418);
xnor U3631 (N_3631,N_3588,N_3549);
or U3632 (N_3632,N_3529,N_3545);
xor U3633 (N_3633,N_3476,N_3503);
and U3634 (N_3634,N_3454,N_3568);
or U3635 (N_3635,N_3505,N_3420);
and U3636 (N_3636,N_3466,N_3402);
nor U3637 (N_3637,N_3552,N_3541);
or U3638 (N_3638,N_3533,N_3490);
xnor U3639 (N_3639,N_3419,N_3566);
nor U3640 (N_3640,N_3532,N_3412);
or U3641 (N_3641,N_3471,N_3407);
or U3642 (N_3642,N_3583,N_3560);
xnor U3643 (N_3643,N_3507,N_3484);
and U3644 (N_3644,N_3478,N_3526);
or U3645 (N_3645,N_3562,N_3460);
xnor U3646 (N_3646,N_3482,N_3534);
nor U3647 (N_3647,N_3578,N_3472);
nor U3648 (N_3648,N_3557,N_3546);
xnor U3649 (N_3649,N_3423,N_3496);
or U3650 (N_3650,N_3446,N_3540);
xnor U3651 (N_3651,N_3594,N_3577);
nand U3652 (N_3652,N_3543,N_3428);
or U3653 (N_3653,N_3409,N_3474);
nand U3654 (N_3654,N_3426,N_3439);
nor U3655 (N_3655,N_3464,N_3470);
nor U3656 (N_3656,N_3579,N_3411);
or U3657 (N_3657,N_3410,N_3551);
nand U3658 (N_3658,N_3587,N_3591);
xor U3659 (N_3659,N_3450,N_3584);
xnor U3660 (N_3660,N_3444,N_3479);
nand U3661 (N_3661,N_3445,N_3401);
and U3662 (N_3662,N_3561,N_3558);
and U3663 (N_3663,N_3542,N_3495);
or U3664 (N_3664,N_3413,N_3504);
or U3665 (N_3665,N_3459,N_3417);
nand U3666 (N_3666,N_3441,N_3597);
and U3667 (N_3667,N_3434,N_3449);
or U3668 (N_3668,N_3569,N_3427);
or U3669 (N_3669,N_3462,N_3415);
nand U3670 (N_3670,N_3554,N_3590);
or U3671 (N_3671,N_3487,N_3519);
nand U3672 (N_3672,N_3502,N_3510);
nor U3673 (N_3673,N_3514,N_3580);
and U3674 (N_3674,N_3559,N_3486);
nor U3675 (N_3675,N_3521,N_3403);
and U3676 (N_3676,N_3455,N_3572);
xnor U3677 (N_3677,N_3452,N_3481);
or U3678 (N_3678,N_3436,N_3406);
or U3679 (N_3679,N_3435,N_3443);
and U3680 (N_3680,N_3405,N_3451);
xnor U3681 (N_3681,N_3424,N_3537);
xor U3682 (N_3682,N_3494,N_3457);
nor U3683 (N_3683,N_3429,N_3469);
and U3684 (N_3684,N_3515,N_3516);
xor U3685 (N_3685,N_3475,N_3465);
and U3686 (N_3686,N_3458,N_3589);
and U3687 (N_3687,N_3548,N_3524);
or U3688 (N_3688,N_3582,N_3595);
xor U3689 (N_3689,N_3570,N_3599);
nor U3690 (N_3690,N_3422,N_3556);
nand U3691 (N_3691,N_3576,N_3497);
nor U3692 (N_3692,N_3528,N_3480);
nand U3693 (N_3693,N_3596,N_3585);
nor U3694 (N_3694,N_3467,N_3575);
or U3695 (N_3695,N_3461,N_3431);
nor U3696 (N_3696,N_3499,N_3567);
nor U3697 (N_3697,N_3438,N_3565);
nand U3698 (N_3698,N_3442,N_3535);
nor U3699 (N_3699,N_3421,N_3506);
nand U3700 (N_3700,N_3570,N_3482);
and U3701 (N_3701,N_3589,N_3532);
nand U3702 (N_3702,N_3466,N_3536);
xnor U3703 (N_3703,N_3424,N_3582);
xor U3704 (N_3704,N_3521,N_3522);
nand U3705 (N_3705,N_3408,N_3515);
or U3706 (N_3706,N_3421,N_3468);
xor U3707 (N_3707,N_3563,N_3568);
nand U3708 (N_3708,N_3528,N_3463);
or U3709 (N_3709,N_3529,N_3565);
and U3710 (N_3710,N_3523,N_3423);
nor U3711 (N_3711,N_3411,N_3556);
or U3712 (N_3712,N_3512,N_3552);
nand U3713 (N_3713,N_3588,N_3536);
xnor U3714 (N_3714,N_3515,N_3577);
and U3715 (N_3715,N_3592,N_3578);
or U3716 (N_3716,N_3424,N_3461);
or U3717 (N_3717,N_3564,N_3563);
and U3718 (N_3718,N_3493,N_3469);
or U3719 (N_3719,N_3485,N_3479);
and U3720 (N_3720,N_3552,N_3557);
xor U3721 (N_3721,N_3473,N_3407);
nor U3722 (N_3722,N_3582,N_3454);
nand U3723 (N_3723,N_3419,N_3548);
xor U3724 (N_3724,N_3410,N_3563);
or U3725 (N_3725,N_3442,N_3528);
xor U3726 (N_3726,N_3515,N_3429);
xnor U3727 (N_3727,N_3418,N_3457);
or U3728 (N_3728,N_3573,N_3491);
nand U3729 (N_3729,N_3521,N_3566);
and U3730 (N_3730,N_3441,N_3409);
xor U3731 (N_3731,N_3509,N_3475);
and U3732 (N_3732,N_3411,N_3499);
nor U3733 (N_3733,N_3519,N_3404);
nor U3734 (N_3734,N_3512,N_3454);
or U3735 (N_3735,N_3504,N_3464);
xor U3736 (N_3736,N_3588,N_3555);
nor U3737 (N_3737,N_3588,N_3460);
and U3738 (N_3738,N_3590,N_3577);
nor U3739 (N_3739,N_3560,N_3445);
xnor U3740 (N_3740,N_3465,N_3598);
nor U3741 (N_3741,N_3431,N_3522);
xnor U3742 (N_3742,N_3432,N_3530);
xor U3743 (N_3743,N_3467,N_3440);
and U3744 (N_3744,N_3508,N_3542);
and U3745 (N_3745,N_3439,N_3463);
or U3746 (N_3746,N_3507,N_3542);
xnor U3747 (N_3747,N_3454,N_3496);
or U3748 (N_3748,N_3401,N_3511);
or U3749 (N_3749,N_3460,N_3402);
xor U3750 (N_3750,N_3462,N_3539);
or U3751 (N_3751,N_3541,N_3599);
xnor U3752 (N_3752,N_3573,N_3556);
nand U3753 (N_3753,N_3432,N_3476);
nor U3754 (N_3754,N_3586,N_3459);
or U3755 (N_3755,N_3480,N_3430);
nand U3756 (N_3756,N_3544,N_3471);
xor U3757 (N_3757,N_3564,N_3476);
xor U3758 (N_3758,N_3559,N_3470);
and U3759 (N_3759,N_3583,N_3490);
nand U3760 (N_3760,N_3459,N_3541);
and U3761 (N_3761,N_3595,N_3530);
nand U3762 (N_3762,N_3402,N_3500);
xor U3763 (N_3763,N_3419,N_3432);
nor U3764 (N_3764,N_3588,N_3424);
or U3765 (N_3765,N_3552,N_3504);
nand U3766 (N_3766,N_3436,N_3514);
or U3767 (N_3767,N_3575,N_3460);
and U3768 (N_3768,N_3405,N_3436);
or U3769 (N_3769,N_3540,N_3429);
or U3770 (N_3770,N_3529,N_3496);
nor U3771 (N_3771,N_3524,N_3568);
nor U3772 (N_3772,N_3449,N_3577);
and U3773 (N_3773,N_3563,N_3441);
nand U3774 (N_3774,N_3441,N_3493);
and U3775 (N_3775,N_3434,N_3562);
nor U3776 (N_3776,N_3419,N_3517);
xnor U3777 (N_3777,N_3509,N_3586);
nand U3778 (N_3778,N_3564,N_3420);
or U3779 (N_3779,N_3584,N_3588);
nand U3780 (N_3780,N_3446,N_3526);
xor U3781 (N_3781,N_3465,N_3593);
xnor U3782 (N_3782,N_3508,N_3571);
nand U3783 (N_3783,N_3562,N_3510);
xnor U3784 (N_3784,N_3567,N_3549);
nand U3785 (N_3785,N_3436,N_3467);
xnor U3786 (N_3786,N_3450,N_3543);
nand U3787 (N_3787,N_3558,N_3439);
or U3788 (N_3788,N_3571,N_3459);
nor U3789 (N_3789,N_3587,N_3427);
or U3790 (N_3790,N_3421,N_3540);
nand U3791 (N_3791,N_3576,N_3492);
nor U3792 (N_3792,N_3443,N_3472);
nand U3793 (N_3793,N_3403,N_3539);
xnor U3794 (N_3794,N_3402,N_3448);
nand U3795 (N_3795,N_3479,N_3527);
and U3796 (N_3796,N_3404,N_3558);
nor U3797 (N_3797,N_3524,N_3410);
nor U3798 (N_3798,N_3523,N_3507);
or U3799 (N_3799,N_3552,N_3580);
nand U3800 (N_3800,N_3778,N_3601);
nor U3801 (N_3801,N_3728,N_3693);
and U3802 (N_3802,N_3605,N_3672);
xnor U3803 (N_3803,N_3734,N_3647);
or U3804 (N_3804,N_3643,N_3727);
nor U3805 (N_3805,N_3718,N_3751);
or U3806 (N_3806,N_3660,N_3763);
xnor U3807 (N_3807,N_3754,N_3673);
nand U3808 (N_3808,N_3646,N_3619);
and U3809 (N_3809,N_3611,N_3769);
xor U3810 (N_3810,N_3635,N_3622);
nand U3811 (N_3811,N_3747,N_3710);
and U3812 (N_3812,N_3670,N_3793);
nor U3813 (N_3813,N_3698,N_3764);
or U3814 (N_3814,N_3796,N_3629);
xor U3815 (N_3815,N_3614,N_3640);
nand U3816 (N_3816,N_3636,N_3729);
or U3817 (N_3817,N_3697,N_3741);
xor U3818 (N_3818,N_3794,N_3624);
and U3819 (N_3819,N_3749,N_3694);
xor U3820 (N_3820,N_3687,N_3669);
nand U3821 (N_3821,N_3630,N_3633);
and U3822 (N_3822,N_3738,N_3665);
nor U3823 (N_3823,N_3655,N_3746);
nor U3824 (N_3824,N_3680,N_3617);
and U3825 (N_3825,N_3637,N_3705);
nand U3826 (N_3826,N_3773,N_3671);
and U3827 (N_3827,N_3604,N_3609);
and U3828 (N_3828,N_3788,N_3799);
xor U3829 (N_3829,N_3752,N_3780);
xor U3830 (N_3830,N_3714,N_3618);
xnor U3831 (N_3831,N_3739,N_3760);
or U3832 (N_3832,N_3613,N_3779);
and U3833 (N_3833,N_3674,N_3690);
nor U3834 (N_3834,N_3709,N_3707);
xor U3835 (N_3835,N_3677,N_3708);
nor U3836 (N_3836,N_3733,N_3731);
or U3837 (N_3837,N_3774,N_3716);
nand U3838 (N_3838,N_3756,N_3696);
nand U3839 (N_3839,N_3645,N_3666);
nor U3840 (N_3840,N_3688,N_3787);
or U3841 (N_3841,N_3686,N_3627);
or U3842 (N_3842,N_3663,N_3790);
or U3843 (N_3843,N_3600,N_3798);
and U3844 (N_3844,N_3650,N_3620);
nand U3845 (N_3845,N_3761,N_3681);
nand U3846 (N_3846,N_3654,N_3717);
xor U3847 (N_3847,N_3766,N_3712);
nor U3848 (N_3848,N_3723,N_3771);
nand U3849 (N_3849,N_3767,N_3626);
xor U3850 (N_3850,N_3699,N_3737);
nand U3851 (N_3851,N_3768,N_3695);
or U3852 (N_3852,N_3616,N_3782);
and U3853 (N_3853,N_3792,N_3607);
or U3854 (N_3854,N_3639,N_3719);
and U3855 (N_3855,N_3631,N_3772);
xor U3856 (N_3856,N_3797,N_3753);
or U3857 (N_3857,N_3726,N_3608);
nand U3858 (N_3858,N_3653,N_3750);
xnor U3859 (N_3859,N_3625,N_3634);
nand U3860 (N_3860,N_3675,N_3784);
xor U3861 (N_3861,N_3678,N_3721);
or U3862 (N_3862,N_3662,N_3612);
or U3863 (N_3863,N_3657,N_3668);
nor U3864 (N_3864,N_3623,N_3762);
nand U3865 (N_3865,N_3757,N_3759);
nand U3866 (N_3866,N_3786,N_3735);
nor U3867 (N_3867,N_3785,N_3685);
nand U3868 (N_3868,N_3664,N_3789);
and U3869 (N_3869,N_3791,N_3722);
and U3870 (N_3870,N_3676,N_3732);
or U3871 (N_3871,N_3667,N_3724);
nand U3872 (N_3872,N_3638,N_3725);
nand U3873 (N_3873,N_3706,N_3621);
or U3874 (N_3874,N_3736,N_3783);
nand U3875 (N_3875,N_3689,N_3682);
and U3876 (N_3876,N_3702,N_3720);
nand U3877 (N_3877,N_3603,N_3684);
nand U3878 (N_3878,N_3777,N_3651);
xnor U3879 (N_3879,N_3743,N_3776);
nand U3880 (N_3880,N_3704,N_3711);
nand U3881 (N_3881,N_3775,N_3656);
and U3882 (N_3882,N_3648,N_3703);
nand U3883 (N_3883,N_3644,N_3652);
or U3884 (N_3884,N_3713,N_3642);
nand U3885 (N_3885,N_3658,N_3755);
xnor U3886 (N_3886,N_3748,N_3795);
nand U3887 (N_3887,N_3606,N_3700);
and U3888 (N_3888,N_3730,N_3758);
and U3889 (N_3889,N_3615,N_3632);
and U3890 (N_3890,N_3661,N_3744);
nand U3891 (N_3891,N_3701,N_3745);
nand U3892 (N_3892,N_3740,N_3691);
and U3893 (N_3893,N_3715,N_3628);
nand U3894 (N_3894,N_3610,N_3770);
or U3895 (N_3895,N_3649,N_3742);
nand U3896 (N_3896,N_3683,N_3765);
nand U3897 (N_3897,N_3781,N_3692);
nand U3898 (N_3898,N_3602,N_3659);
nor U3899 (N_3899,N_3641,N_3679);
xor U3900 (N_3900,N_3668,N_3654);
and U3901 (N_3901,N_3647,N_3633);
or U3902 (N_3902,N_3675,N_3688);
nand U3903 (N_3903,N_3760,N_3642);
or U3904 (N_3904,N_3652,N_3725);
nor U3905 (N_3905,N_3630,N_3621);
nand U3906 (N_3906,N_3667,N_3725);
nor U3907 (N_3907,N_3685,N_3724);
or U3908 (N_3908,N_3773,N_3628);
xor U3909 (N_3909,N_3714,N_3649);
and U3910 (N_3910,N_3684,N_3726);
or U3911 (N_3911,N_3676,N_3646);
and U3912 (N_3912,N_3686,N_3723);
and U3913 (N_3913,N_3624,N_3782);
or U3914 (N_3914,N_3736,N_3643);
nand U3915 (N_3915,N_3701,N_3618);
nand U3916 (N_3916,N_3750,N_3640);
nand U3917 (N_3917,N_3715,N_3748);
and U3918 (N_3918,N_3652,N_3620);
and U3919 (N_3919,N_3670,N_3659);
or U3920 (N_3920,N_3622,N_3606);
nor U3921 (N_3921,N_3746,N_3722);
nor U3922 (N_3922,N_3691,N_3638);
xor U3923 (N_3923,N_3750,N_3686);
or U3924 (N_3924,N_3615,N_3734);
nand U3925 (N_3925,N_3734,N_3697);
and U3926 (N_3926,N_3658,N_3600);
xor U3927 (N_3927,N_3742,N_3734);
xnor U3928 (N_3928,N_3744,N_3713);
xor U3929 (N_3929,N_3670,N_3680);
nor U3930 (N_3930,N_3702,N_3790);
nor U3931 (N_3931,N_3715,N_3648);
nor U3932 (N_3932,N_3637,N_3616);
or U3933 (N_3933,N_3766,N_3659);
or U3934 (N_3934,N_3708,N_3797);
and U3935 (N_3935,N_3620,N_3689);
nand U3936 (N_3936,N_3763,N_3734);
and U3937 (N_3937,N_3789,N_3709);
nor U3938 (N_3938,N_3613,N_3740);
nor U3939 (N_3939,N_3760,N_3618);
or U3940 (N_3940,N_3705,N_3615);
and U3941 (N_3941,N_3624,N_3790);
nand U3942 (N_3942,N_3612,N_3736);
nor U3943 (N_3943,N_3744,N_3607);
and U3944 (N_3944,N_3657,N_3738);
nand U3945 (N_3945,N_3639,N_3709);
nor U3946 (N_3946,N_3748,N_3719);
or U3947 (N_3947,N_3731,N_3712);
or U3948 (N_3948,N_3785,N_3601);
nand U3949 (N_3949,N_3761,N_3710);
nand U3950 (N_3950,N_3775,N_3799);
or U3951 (N_3951,N_3685,N_3730);
and U3952 (N_3952,N_3767,N_3663);
xnor U3953 (N_3953,N_3653,N_3605);
and U3954 (N_3954,N_3668,N_3778);
or U3955 (N_3955,N_3792,N_3674);
and U3956 (N_3956,N_3693,N_3635);
nand U3957 (N_3957,N_3679,N_3689);
nor U3958 (N_3958,N_3722,N_3795);
xnor U3959 (N_3959,N_3620,N_3772);
and U3960 (N_3960,N_3643,N_3650);
and U3961 (N_3961,N_3736,N_3793);
xor U3962 (N_3962,N_3741,N_3628);
xor U3963 (N_3963,N_3620,N_3685);
or U3964 (N_3964,N_3720,N_3749);
xor U3965 (N_3965,N_3762,N_3768);
or U3966 (N_3966,N_3632,N_3618);
nand U3967 (N_3967,N_3602,N_3795);
nor U3968 (N_3968,N_3612,N_3761);
or U3969 (N_3969,N_3698,N_3789);
and U3970 (N_3970,N_3637,N_3727);
nor U3971 (N_3971,N_3720,N_3691);
xor U3972 (N_3972,N_3741,N_3714);
nor U3973 (N_3973,N_3612,N_3673);
nand U3974 (N_3974,N_3677,N_3657);
nand U3975 (N_3975,N_3607,N_3751);
nand U3976 (N_3976,N_3700,N_3699);
xnor U3977 (N_3977,N_3628,N_3799);
and U3978 (N_3978,N_3798,N_3763);
nand U3979 (N_3979,N_3624,N_3706);
nand U3980 (N_3980,N_3624,N_3676);
nor U3981 (N_3981,N_3773,N_3674);
or U3982 (N_3982,N_3711,N_3787);
xor U3983 (N_3983,N_3699,N_3746);
xor U3984 (N_3984,N_3695,N_3656);
and U3985 (N_3985,N_3674,N_3787);
or U3986 (N_3986,N_3651,N_3688);
xor U3987 (N_3987,N_3685,N_3757);
or U3988 (N_3988,N_3717,N_3631);
nor U3989 (N_3989,N_3678,N_3695);
nand U3990 (N_3990,N_3663,N_3711);
nand U3991 (N_3991,N_3758,N_3698);
nor U3992 (N_3992,N_3696,N_3747);
and U3993 (N_3993,N_3627,N_3613);
nor U3994 (N_3994,N_3721,N_3710);
nor U3995 (N_3995,N_3600,N_3797);
nor U3996 (N_3996,N_3643,N_3697);
and U3997 (N_3997,N_3655,N_3683);
nand U3998 (N_3998,N_3675,N_3742);
and U3999 (N_3999,N_3694,N_3767);
xnor U4000 (N_4000,N_3972,N_3929);
xnor U4001 (N_4001,N_3978,N_3871);
nand U4002 (N_4002,N_3825,N_3916);
nand U4003 (N_4003,N_3884,N_3936);
nor U4004 (N_4004,N_3974,N_3900);
and U4005 (N_4005,N_3836,N_3833);
and U4006 (N_4006,N_3939,N_3914);
and U4007 (N_4007,N_3860,N_3812);
nand U4008 (N_4008,N_3845,N_3906);
or U4009 (N_4009,N_3997,N_3928);
xnor U4010 (N_4010,N_3954,N_3941);
nor U4011 (N_4011,N_3927,N_3985);
nand U4012 (N_4012,N_3885,N_3951);
nor U4013 (N_4013,N_3804,N_3924);
and U4014 (N_4014,N_3926,N_3808);
nor U4015 (N_4015,N_3983,N_3887);
xor U4016 (N_4016,N_3908,N_3842);
xor U4017 (N_4017,N_3988,N_3953);
or U4018 (N_4018,N_3907,N_3990);
nand U4019 (N_4019,N_3805,N_3987);
or U4020 (N_4020,N_3854,N_3819);
xor U4021 (N_4021,N_3933,N_3981);
nand U4022 (N_4022,N_3940,N_3835);
xnor U4023 (N_4023,N_3991,N_3913);
xor U4024 (N_4024,N_3801,N_3866);
or U4025 (N_4025,N_3894,N_3868);
nor U4026 (N_4026,N_3862,N_3979);
nand U4027 (N_4027,N_3901,N_3920);
and U4028 (N_4028,N_3817,N_3899);
or U4029 (N_4029,N_3925,N_3896);
or U4030 (N_4030,N_3898,N_3861);
or U4031 (N_4031,N_3982,N_3856);
xnor U4032 (N_4032,N_3840,N_3917);
and U4033 (N_4033,N_3968,N_3932);
or U4034 (N_4034,N_3998,N_3930);
nor U4035 (N_4035,N_3943,N_3823);
and U4036 (N_4036,N_3904,N_3905);
or U4037 (N_4037,N_3975,N_3843);
and U4038 (N_4038,N_3877,N_3879);
nor U4039 (N_4039,N_3824,N_3820);
or U4040 (N_4040,N_3855,N_3977);
nor U4041 (N_4041,N_3865,N_3809);
nand U4042 (N_4042,N_3857,N_3910);
xnor U4043 (N_4043,N_3837,N_3955);
nand U4044 (N_4044,N_3918,N_3807);
and U4045 (N_4045,N_3969,N_3880);
nor U4046 (N_4046,N_3827,N_3959);
xor U4047 (N_4047,N_3851,N_3944);
xnor U4048 (N_4048,N_3986,N_3970);
nand U4049 (N_4049,N_3995,N_3922);
nand U4050 (N_4050,N_3889,N_3867);
nor U4051 (N_4051,N_3911,N_3859);
xnor U4052 (N_4052,N_3903,N_3996);
and U4053 (N_4053,N_3829,N_3844);
and U4054 (N_4054,N_3960,N_3912);
nand U4055 (N_4055,N_3878,N_3950);
nand U4056 (N_4056,N_3947,N_3846);
xnor U4057 (N_4057,N_3814,N_3942);
nand U4058 (N_4058,N_3923,N_3881);
nor U4059 (N_4059,N_3831,N_3803);
nand U4060 (N_4060,N_3957,N_3931);
or U4061 (N_4061,N_3921,N_3832);
nor U4062 (N_4062,N_3872,N_3875);
nor U4063 (N_4063,N_3863,N_3909);
xor U4064 (N_4064,N_3895,N_3853);
and U4065 (N_4065,N_3810,N_3902);
and U4066 (N_4066,N_3948,N_3848);
or U4067 (N_4067,N_3870,N_3811);
nand U4068 (N_4068,N_3993,N_3838);
or U4069 (N_4069,N_3828,N_3893);
or U4070 (N_4070,N_3873,N_3821);
and U4071 (N_4071,N_3883,N_3963);
nor U4072 (N_4072,N_3962,N_3800);
nand U4073 (N_4073,N_3984,N_3839);
xor U4074 (N_4074,N_3976,N_3806);
and U4075 (N_4075,N_3834,N_3864);
nor U4076 (N_4076,N_3965,N_3826);
or U4077 (N_4077,N_3992,N_3830);
nor U4078 (N_4078,N_3841,N_3888);
or U4079 (N_4079,N_3850,N_3946);
nand U4080 (N_4080,N_3937,N_3934);
nor U4081 (N_4081,N_3891,N_3869);
or U4082 (N_4082,N_3886,N_3994);
and U4083 (N_4083,N_3892,N_3938);
xnor U4084 (N_4084,N_3958,N_3999);
and U4085 (N_4085,N_3849,N_3816);
nand U4086 (N_4086,N_3973,N_3822);
xnor U4087 (N_4087,N_3874,N_3935);
or U4088 (N_4088,N_3945,N_3882);
nor U4089 (N_4089,N_3847,N_3964);
and U4090 (N_4090,N_3980,N_3802);
xnor U4091 (N_4091,N_3949,N_3952);
xnor U4092 (N_4092,N_3858,N_3915);
or U4093 (N_4093,N_3815,N_3971);
or U4094 (N_4094,N_3890,N_3989);
nand U4095 (N_4095,N_3897,N_3876);
and U4096 (N_4096,N_3818,N_3961);
xnor U4097 (N_4097,N_3967,N_3919);
nand U4098 (N_4098,N_3956,N_3852);
xor U4099 (N_4099,N_3966,N_3813);
or U4100 (N_4100,N_3853,N_3827);
nor U4101 (N_4101,N_3823,N_3941);
and U4102 (N_4102,N_3824,N_3815);
nor U4103 (N_4103,N_3893,N_3866);
or U4104 (N_4104,N_3846,N_3918);
nor U4105 (N_4105,N_3830,N_3859);
xor U4106 (N_4106,N_3862,N_3864);
nor U4107 (N_4107,N_3953,N_3995);
or U4108 (N_4108,N_3929,N_3870);
nor U4109 (N_4109,N_3918,N_3941);
nand U4110 (N_4110,N_3861,N_3948);
xor U4111 (N_4111,N_3872,N_3840);
nand U4112 (N_4112,N_3854,N_3974);
and U4113 (N_4113,N_3821,N_3858);
xnor U4114 (N_4114,N_3842,N_3910);
nand U4115 (N_4115,N_3857,N_3970);
or U4116 (N_4116,N_3810,N_3806);
and U4117 (N_4117,N_3826,N_3999);
nor U4118 (N_4118,N_3808,N_3806);
nand U4119 (N_4119,N_3810,N_3873);
and U4120 (N_4120,N_3983,N_3919);
xnor U4121 (N_4121,N_3833,N_3963);
nor U4122 (N_4122,N_3895,N_3801);
nor U4123 (N_4123,N_3875,N_3977);
and U4124 (N_4124,N_3880,N_3939);
xnor U4125 (N_4125,N_3904,N_3870);
nor U4126 (N_4126,N_3904,N_3932);
xnor U4127 (N_4127,N_3802,N_3977);
and U4128 (N_4128,N_3899,N_3896);
xnor U4129 (N_4129,N_3849,N_3883);
and U4130 (N_4130,N_3880,N_3887);
nand U4131 (N_4131,N_3873,N_3823);
or U4132 (N_4132,N_3903,N_3972);
xor U4133 (N_4133,N_3855,N_3967);
and U4134 (N_4134,N_3805,N_3925);
or U4135 (N_4135,N_3872,N_3958);
xor U4136 (N_4136,N_3949,N_3957);
or U4137 (N_4137,N_3975,N_3834);
xor U4138 (N_4138,N_3892,N_3919);
and U4139 (N_4139,N_3951,N_3869);
or U4140 (N_4140,N_3942,N_3949);
nor U4141 (N_4141,N_3979,N_3930);
nor U4142 (N_4142,N_3871,N_3866);
or U4143 (N_4143,N_3906,N_3985);
xor U4144 (N_4144,N_3917,N_3887);
or U4145 (N_4145,N_3861,N_3859);
xnor U4146 (N_4146,N_3900,N_3824);
and U4147 (N_4147,N_3897,N_3848);
and U4148 (N_4148,N_3994,N_3911);
and U4149 (N_4149,N_3822,N_3855);
nor U4150 (N_4150,N_3937,N_3905);
nor U4151 (N_4151,N_3945,N_3934);
nand U4152 (N_4152,N_3859,N_3996);
nor U4153 (N_4153,N_3844,N_3857);
and U4154 (N_4154,N_3835,N_3888);
and U4155 (N_4155,N_3922,N_3951);
nor U4156 (N_4156,N_3973,N_3899);
xnor U4157 (N_4157,N_3917,N_3825);
xnor U4158 (N_4158,N_3884,N_3862);
and U4159 (N_4159,N_3882,N_3849);
and U4160 (N_4160,N_3867,N_3866);
nor U4161 (N_4161,N_3959,N_3980);
and U4162 (N_4162,N_3958,N_3964);
and U4163 (N_4163,N_3864,N_3918);
xor U4164 (N_4164,N_3846,N_3911);
nor U4165 (N_4165,N_3893,N_3804);
xnor U4166 (N_4166,N_3813,N_3801);
nor U4167 (N_4167,N_3845,N_3836);
nor U4168 (N_4168,N_3874,N_3837);
and U4169 (N_4169,N_3827,N_3924);
or U4170 (N_4170,N_3967,N_3890);
xor U4171 (N_4171,N_3955,N_3951);
and U4172 (N_4172,N_3988,N_3898);
xnor U4173 (N_4173,N_3822,N_3804);
nor U4174 (N_4174,N_3951,N_3994);
xor U4175 (N_4175,N_3981,N_3915);
nor U4176 (N_4176,N_3829,N_3923);
xnor U4177 (N_4177,N_3991,N_3966);
and U4178 (N_4178,N_3875,N_3802);
or U4179 (N_4179,N_3941,N_3970);
and U4180 (N_4180,N_3878,N_3843);
or U4181 (N_4181,N_3876,N_3832);
xor U4182 (N_4182,N_3837,N_3818);
nand U4183 (N_4183,N_3868,N_3925);
nand U4184 (N_4184,N_3802,N_3940);
and U4185 (N_4185,N_3993,N_3816);
xor U4186 (N_4186,N_3879,N_3951);
and U4187 (N_4187,N_3922,N_3989);
xnor U4188 (N_4188,N_3814,N_3824);
xnor U4189 (N_4189,N_3800,N_3992);
nor U4190 (N_4190,N_3944,N_3932);
xor U4191 (N_4191,N_3883,N_3952);
nand U4192 (N_4192,N_3837,N_3946);
xnor U4193 (N_4193,N_3940,N_3804);
and U4194 (N_4194,N_3846,N_3977);
nand U4195 (N_4195,N_3893,N_3888);
or U4196 (N_4196,N_3948,N_3927);
nand U4197 (N_4197,N_3864,N_3856);
and U4198 (N_4198,N_3884,N_3801);
nand U4199 (N_4199,N_3924,N_3886);
nand U4200 (N_4200,N_4171,N_4005);
and U4201 (N_4201,N_4123,N_4010);
or U4202 (N_4202,N_4133,N_4075);
or U4203 (N_4203,N_4193,N_4114);
nor U4204 (N_4204,N_4197,N_4099);
and U4205 (N_4205,N_4032,N_4139);
xnor U4206 (N_4206,N_4122,N_4044);
xor U4207 (N_4207,N_4059,N_4194);
or U4208 (N_4208,N_4009,N_4104);
and U4209 (N_4209,N_4108,N_4036);
nand U4210 (N_4210,N_4024,N_4174);
xnor U4211 (N_4211,N_4021,N_4096);
nor U4212 (N_4212,N_4007,N_4144);
nor U4213 (N_4213,N_4074,N_4086);
xor U4214 (N_4214,N_4127,N_4110);
or U4215 (N_4215,N_4149,N_4196);
nor U4216 (N_4216,N_4152,N_4017);
nor U4217 (N_4217,N_4178,N_4120);
or U4218 (N_4218,N_4186,N_4091);
and U4219 (N_4219,N_4034,N_4172);
xor U4220 (N_4220,N_4160,N_4060);
or U4221 (N_4221,N_4042,N_4142);
nand U4222 (N_4222,N_4089,N_4100);
xor U4223 (N_4223,N_4015,N_4106);
and U4224 (N_4224,N_4198,N_4191);
or U4225 (N_4225,N_4169,N_4097);
and U4226 (N_4226,N_4061,N_4130);
nor U4227 (N_4227,N_4185,N_4033);
or U4228 (N_4228,N_4125,N_4037);
xnor U4229 (N_4229,N_4107,N_4181);
xnor U4230 (N_4230,N_4065,N_4039);
nor U4231 (N_4231,N_4078,N_4189);
nand U4232 (N_4232,N_4148,N_4051);
and U4233 (N_4233,N_4047,N_4093);
or U4234 (N_4234,N_4069,N_4068);
and U4235 (N_4235,N_4132,N_4111);
or U4236 (N_4236,N_4176,N_4105);
and U4237 (N_4237,N_4063,N_4043);
and U4238 (N_4238,N_4013,N_4118);
nand U4239 (N_4239,N_4066,N_4025);
nand U4240 (N_4240,N_4143,N_4035);
or U4241 (N_4241,N_4081,N_4006);
xnor U4242 (N_4242,N_4050,N_4150);
and U4243 (N_4243,N_4072,N_4048);
and U4244 (N_4244,N_4115,N_4195);
nor U4245 (N_4245,N_4022,N_4095);
nor U4246 (N_4246,N_4147,N_4012);
xnor U4247 (N_4247,N_4062,N_4164);
nand U4248 (N_4248,N_4016,N_4073);
nor U4249 (N_4249,N_4192,N_4056);
and U4250 (N_4250,N_4134,N_4151);
nor U4251 (N_4251,N_4136,N_4002);
or U4252 (N_4252,N_4071,N_4166);
nor U4253 (N_4253,N_4085,N_4019);
nor U4254 (N_4254,N_4087,N_4199);
nor U4255 (N_4255,N_4040,N_4029);
nand U4256 (N_4256,N_4156,N_4109);
or U4257 (N_4257,N_4161,N_4159);
or U4258 (N_4258,N_4020,N_4131);
nor U4259 (N_4259,N_4113,N_4102);
nor U4260 (N_4260,N_4090,N_4054);
nand U4261 (N_4261,N_4101,N_4018);
or U4262 (N_4262,N_4129,N_4182);
and U4263 (N_4263,N_4045,N_4146);
nor U4264 (N_4264,N_4011,N_4165);
xor U4265 (N_4265,N_4112,N_4121);
or U4266 (N_4266,N_4046,N_4076);
or U4267 (N_4267,N_4141,N_4162);
xnor U4268 (N_4268,N_4103,N_4094);
or U4269 (N_4269,N_4117,N_4180);
xnor U4270 (N_4270,N_4080,N_4053);
or U4271 (N_4271,N_4083,N_4135);
xnor U4272 (N_4272,N_4153,N_4052);
xnor U4273 (N_4273,N_4031,N_4023);
xnor U4274 (N_4274,N_4064,N_4155);
xnor U4275 (N_4275,N_4116,N_4077);
or U4276 (N_4276,N_4008,N_4167);
nor U4277 (N_4277,N_4168,N_4092);
xor U4278 (N_4278,N_4082,N_4026);
nand U4279 (N_4279,N_4014,N_4079);
and U4280 (N_4280,N_4030,N_4188);
nand U4281 (N_4281,N_4067,N_4070);
or U4282 (N_4282,N_4177,N_4098);
xor U4283 (N_4283,N_4184,N_4173);
nor U4284 (N_4284,N_4126,N_4058);
and U4285 (N_4285,N_4128,N_4004);
nor U4286 (N_4286,N_4183,N_4190);
nor U4287 (N_4287,N_4137,N_4154);
nor U4288 (N_4288,N_4084,N_4140);
xor U4289 (N_4289,N_4000,N_4049);
nor U4290 (N_4290,N_4163,N_4027);
nand U4291 (N_4291,N_4028,N_4001);
nor U4292 (N_4292,N_4145,N_4055);
and U4293 (N_4293,N_4124,N_4119);
or U4294 (N_4294,N_4138,N_4057);
xor U4295 (N_4295,N_4170,N_4003);
and U4296 (N_4296,N_4157,N_4158);
or U4297 (N_4297,N_4175,N_4041);
xnor U4298 (N_4298,N_4187,N_4088);
nand U4299 (N_4299,N_4038,N_4179);
nand U4300 (N_4300,N_4000,N_4135);
and U4301 (N_4301,N_4089,N_4015);
nor U4302 (N_4302,N_4171,N_4074);
nor U4303 (N_4303,N_4084,N_4148);
xnor U4304 (N_4304,N_4164,N_4007);
xor U4305 (N_4305,N_4125,N_4140);
and U4306 (N_4306,N_4031,N_4139);
nor U4307 (N_4307,N_4177,N_4159);
or U4308 (N_4308,N_4000,N_4148);
xor U4309 (N_4309,N_4110,N_4011);
nor U4310 (N_4310,N_4136,N_4080);
nand U4311 (N_4311,N_4187,N_4033);
nor U4312 (N_4312,N_4008,N_4080);
and U4313 (N_4313,N_4035,N_4005);
xor U4314 (N_4314,N_4032,N_4140);
and U4315 (N_4315,N_4149,N_4184);
nand U4316 (N_4316,N_4064,N_4143);
or U4317 (N_4317,N_4169,N_4035);
and U4318 (N_4318,N_4121,N_4186);
xor U4319 (N_4319,N_4192,N_4120);
nand U4320 (N_4320,N_4123,N_4072);
nand U4321 (N_4321,N_4042,N_4176);
xnor U4322 (N_4322,N_4046,N_4052);
xor U4323 (N_4323,N_4016,N_4176);
and U4324 (N_4324,N_4019,N_4162);
xnor U4325 (N_4325,N_4094,N_4039);
nand U4326 (N_4326,N_4041,N_4059);
nand U4327 (N_4327,N_4101,N_4093);
and U4328 (N_4328,N_4119,N_4189);
and U4329 (N_4329,N_4031,N_4035);
xor U4330 (N_4330,N_4029,N_4114);
nor U4331 (N_4331,N_4072,N_4148);
or U4332 (N_4332,N_4063,N_4141);
xor U4333 (N_4333,N_4007,N_4121);
nand U4334 (N_4334,N_4189,N_4179);
nand U4335 (N_4335,N_4011,N_4066);
or U4336 (N_4336,N_4198,N_4077);
nand U4337 (N_4337,N_4164,N_4017);
nand U4338 (N_4338,N_4182,N_4192);
nor U4339 (N_4339,N_4011,N_4139);
nor U4340 (N_4340,N_4180,N_4099);
or U4341 (N_4341,N_4126,N_4117);
nor U4342 (N_4342,N_4094,N_4182);
nand U4343 (N_4343,N_4195,N_4108);
nor U4344 (N_4344,N_4141,N_4175);
and U4345 (N_4345,N_4088,N_4143);
or U4346 (N_4346,N_4175,N_4066);
nor U4347 (N_4347,N_4122,N_4183);
or U4348 (N_4348,N_4040,N_4020);
xnor U4349 (N_4349,N_4194,N_4138);
nor U4350 (N_4350,N_4078,N_4012);
xor U4351 (N_4351,N_4004,N_4023);
nor U4352 (N_4352,N_4030,N_4016);
and U4353 (N_4353,N_4184,N_4176);
and U4354 (N_4354,N_4004,N_4131);
and U4355 (N_4355,N_4140,N_4110);
or U4356 (N_4356,N_4000,N_4017);
xor U4357 (N_4357,N_4043,N_4191);
nor U4358 (N_4358,N_4005,N_4084);
or U4359 (N_4359,N_4069,N_4102);
nand U4360 (N_4360,N_4129,N_4107);
xor U4361 (N_4361,N_4013,N_4055);
or U4362 (N_4362,N_4165,N_4002);
or U4363 (N_4363,N_4132,N_4054);
nor U4364 (N_4364,N_4082,N_4152);
xor U4365 (N_4365,N_4094,N_4012);
nand U4366 (N_4366,N_4110,N_4184);
nor U4367 (N_4367,N_4027,N_4167);
or U4368 (N_4368,N_4036,N_4123);
xor U4369 (N_4369,N_4147,N_4189);
nor U4370 (N_4370,N_4064,N_4022);
nor U4371 (N_4371,N_4056,N_4155);
nand U4372 (N_4372,N_4163,N_4138);
xor U4373 (N_4373,N_4093,N_4132);
nand U4374 (N_4374,N_4087,N_4017);
or U4375 (N_4375,N_4008,N_4067);
nand U4376 (N_4376,N_4088,N_4014);
nand U4377 (N_4377,N_4112,N_4172);
nor U4378 (N_4378,N_4182,N_4150);
nor U4379 (N_4379,N_4182,N_4081);
nand U4380 (N_4380,N_4193,N_4038);
or U4381 (N_4381,N_4167,N_4039);
or U4382 (N_4382,N_4114,N_4034);
nor U4383 (N_4383,N_4169,N_4055);
nor U4384 (N_4384,N_4116,N_4056);
and U4385 (N_4385,N_4046,N_4048);
or U4386 (N_4386,N_4190,N_4131);
or U4387 (N_4387,N_4017,N_4151);
nor U4388 (N_4388,N_4134,N_4033);
nand U4389 (N_4389,N_4113,N_4010);
or U4390 (N_4390,N_4161,N_4014);
and U4391 (N_4391,N_4094,N_4081);
nor U4392 (N_4392,N_4167,N_4062);
or U4393 (N_4393,N_4130,N_4175);
xnor U4394 (N_4394,N_4189,N_4145);
nand U4395 (N_4395,N_4077,N_4102);
or U4396 (N_4396,N_4078,N_4137);
nand U4397 (N_4397,N_4047,N_4065);
and U4398 (N_4398,N_4040,N_4197);
nand U4399 (N_4399,N_4011,N_4014);
and U4400 (N_4400,N_4270,N_4330);
or U4401 (N_4401,N_4357,N_4208);
or U4402 (N_4402,N_4314,N_4299);
and U4403 (N_4403,N_4252,N_4376);
nor U4404 (N_4404,N_4352,N_4259);
xor U4405 (N_4405,N_4277,N_4385);
nor U4406 (N_4406,N_4294,N_4204);
nand U4407 (N_4407,N_4214,N_4301);
nor U4408 (N_4408,N_4358,N_4390);
and U4409 (N_4409,N_4266,N_4386);
or U4410 (N_4410,N_4202,N_4219);
xor U4411 (N_4411,N_4273,N_4293);
xnor U4412 (N_4412,N_4364,N_4285);
nand U4413 (N_4413,N_4332,N_4227);
and U4414 (N_4414,N_4262,N_4324);
nor U4415 (N_4415,N_4297,N_4302);
or U4416 (N_4416,N_4278,N_4315);
xor U4417 (N_4417,N_4343,N_4247);
and U4418 (N_4418,N_4321,N_4329);
nand U4419 (N_4419,N_4393,N_4284);
or U4420 (N_4420,N_4215,N_4373);
nor U4421 (N_4421,N_4280,N_4379);
nor U4422 (N_4422,N_4375,N_4250);
and U4423 (N_4423,N_4355,N_4226);
or U4424 (N_4424,N_4229,N_4279);
nand U4425 (N_4425,N_4367,N_4241);
and U4426 (N_4426,N_4399,N_4256);
and U4427 (N_4427,N_4337,N_4394);
xnor U4428 (N_4428,N_4327,N_4395);
or U4429 (N_4429,N_4372,N_4397);
or U4430 (N_4430,N_4368,N_4272);
nor U4431 (N_4431,N_4307,N_4246);
nand U4432 (N_4432,N_4310,N_4360);
xor U4433 (N_4433,N_4371,N_4275);
nor U4434 (N_4434,N_4331,N_4291);
xor U4435 (N_4435,N_4362,N_4350);
or U4436 (N_4436,N_4220,N_4206);
xnor U4437 (N_4437,N_4378,N_4295);
or U4438 (N_4438,N_4290,N_4274);
nand U4439 (N_4439,N_4312,N_4354);
xnor U4440 (N_4440,N_4351,N_4213);
or U4441 (N_4441,N_4205,N_4269);
nand U4442 (N_4442,N_4369,N_4338);
xor U4443 (N_4443,N_4347,N_4305);
and U4444 (N_4444,N_4242,N_4257);
xor U4445 (N_4445,N_4359,N_4391);
nor U4446 (N_4446,N_4311,N_4382);
xnor U4447 (N_4447,N_4203,N_4230);
xnor U4448 (N_4448,N_4323,N_4335);
xor U4449 (N_4449,N_4344,N_4346);
or U4450 (N_4450,N_4328,N_4388);
xnor U4451 (N_4451,N_4210,N_4207);
nand U4452 (N_4452,N_4377,N_4313);
or U4453 (N_4453,N_4356,N_4211);
nand U4454 (N_4454,N_4339,N_4325);
nor U4455 (N_4455,N_4271,N_4392);
xor U4456 (N_4456,N_4248,N_4300);
xor U4457 (N_4457,N_4234,N_4387);
or U4458 (N_4458,N_4303,N_4308);
and U4459 (N_4459,N_4217,N_4288);
xor U4460 (N_4460,N_4260,N_4263);
xnor U4461 (N_4461,N_4232,N_4318);
and U4462 (N_4462,N_4365,N_4268);
and U4463 (N_4463,N_4363,N_4201);
xor U4464 (N_4464,N_4254,N_4340);
nor U4465 (N_4465,N_4243,N_4267);
and U4466 (N_4466,N_4304,N_4240);
or U4467 (N_4467,N_4228,N_4286);
and U4468 (N_4468,N_4233,N_4231);
and U4469 (N_4469,N_4341,N_4396);
and U4470 (N_4470,N_4381,N_4349);
nand U4471 (N_4471,N_4265,N_4366);
xor U4472 (N_4472,N_4353,N_4380);
and U4473 (N_4473,N_4389,N_4245);
xor U4474 (N_4474,N_4223,N_4336);
nand U4475 (N_4475,N_4342,N_4306);
xnor U4476 (N_4476,N_4289,N_4370);
xnor U4477 (N_4477,N_4225,N_4212);
nand U4478 (N_4478,N_4283,N_4296);
xor U4479 (N_4479,N_4345,N_4276);
and U4480 (N_4480,N_4218,N_4224);
and U4481 (N_4481,N_4281,N_4361);
or U4482 (N_4482,N_4322,N_4384);
xnor U4483 (N_4483,N_4239,N_4348);
nor U4484 (N_4484,N_4334,N_4316);
xor U4485 (N_4485,N_4255,N_4317);
xor U4486 (N_4486,N_4319,N_4216);
nand U4487 (N_4487,N_4249,N_4309);
xor U4488 (N_4488,N_4237,N_4258);
nor U4489 (N_4489,N_4238,N_4292);
and U4490 (N_4490,N_4236,N_4261);
and U4491 (N_4491,N_4298,N_4200);
and U4492 (N_4492,N_4221,N_4333);
and U4493 (N_4493,N_4383,N_4398);
or U4494 (N_4494,N_4244,N_4282);
nand U4495 (N_4495,N_4251,N_4222);
nand U4496 (N_4496,N_4253,N_4235);
and U4497 (N_4497,N_4209,N_4320);
nor U4498 (N_4498,N_4374,N_4264);
or U4499 (N_4499,N_4287,N_4326);
nand U4500 (N_4500,N_4279,N_4261);
nor U4501 (N_4501,N_4349,N_4243);
nor U4502 (N_4502,N_4362,N_4217);
or U4503 (N_4503,N_4290,N_4293);
and U4504 (N_4504,N_4224,N_4342);
and U4505 (N_4505,N_4361,N_4376);
nor U4506 (N_4506,N_4212,N_4268);
xnor U4507 (N_4507,N_4223,N_4284);
nand U4508 (N_4508,N_4298,N_4282);
or U4509 (N_4509,N_4312,N_4257);
or U4510 (N_4510,N_4342,N_4309);
and U4511 (N_4511,N_4233,N_4340);
xor U4512 (N_4512,N_4322,N_4352);
and U4513 (N_4513,N_4304,N_4217);
or U4514 (N_4514,N_4305,N_4314);
nor U4515 (N_4515,N_4397,N_4224);
or U4516 (N_4516,N_4220,N_4277);
nor U4517 (N_4517,N_4272,N_4396);
xnor U4518 (N_4518,N_4241,N_4307);
nor U4519 (N_4519,N_4369,N_4227);
and U4520 (N_4520,N_4225,N_4355);
nand U4521 (N_4521,N_4217,N_4222);
nor U4522 (N_4522,N_4395,N_4325);
nand U4523 (N_4523,N_4340,N_4317);
xor U4524 (N_4524,N_4300,N_4371);
and U4525 (N_4525,N_4379,N_4249);
or U4526 (N_4526,N_4248,N_4254);
xor U4527 (N_4527,N_4369,N_4239);
and U4528 (N_4528,N_4353,N_4213);
nand U4529 (N_4529,N_4217,N_4393);
nand U4530 (N_4530,N_4240,N_4384);
or U4531 (N_4531,N_4391,N_4242);
or U4532 (N_4532,N_4301,N_4293);
or U4533 (N_4533,N_4202,N_4203);
nor U4534 (N_4534,N_4250,N_4318);
nor U4535 (N_4535,N_4255,N_4280);
xor U4536 (N_4536,N_4343,N_4223);
nor U4537 (N_4537,N_4263,N_4353);
and U4538 (N_4538,N_4352,N_4389);
nand U4539 (N_4539,N_4275,N_4200);
nand U4540 (N_4540,N_4329,N_4322);
or U4541 (N_4541,N_4284,N_4266);
nand U4542 (N_4542,N_4217,N_4325);
nor U4543 (N_4543,N_4334,N_4366);
nor U4544 (N_4544,N_4329,N_4224);
or U4545 (N_4545,N_4228,N_4311);
xor U4546 (N_4546,N_4220,N_4236);
nor U4547 (N_4547,N_4275,N_4216);
or U4548 (N_4548,N_4380,N_4205);
nand U4549 (N_4549,N_4278,N_4375);
and U4550 (N_4550,N_4388,N_4398);
and U4551 (N_4551,N_4278,N_4210);
nor U4552 (N_4552,N_4303,N_4343);
nand U4553 (N_4553,N_4238,N_4356);
or U4554 (N_4554,N_4281,N_4265);
and U4555 (N_4555,N_4374,N_4364);
nor U4556 (N_4556,N_4340,N_4227);
and U4557 (N_4557,N_4380,N_4391);
nand U4558 (N_4558,N_4343,N_4300);
and U4559 (N_4559,N_4367,N_4382);
or U4560 (N_4560,N_4329,N_4259);
nor U4561 (N_4561,N_4201,N_4336);
nor U4562 (N_4562,N_4326,N_4344);
nor U4563 (N_4563,N_4275,N_4387);
nor U4564 (N_4564,N_4390,N_4279);
and U4565 (N_4565,N_4288,N_4239);
nor U4566 (N_4566,N_4327,N_4396);
or U4567 (N_4567,N_4221,N_4357);
or U4568 (N_4568,N_4210,N_4242);
nor U4569 (N_4569,N_4272,N_4338);
xor U4570 (N_4570,N_4376,N_4228);
xor U4571 (N_4571,N_4306,N_4360);
and U4572 (N_4572,N_4364,N_4336);
or U4573 (N_4573,N_4395,N_4233);
or U4574 (N_4574,N_4345,N_4205);
and U4575 (N_4575,N_4269,N_4325);
xor U4576 (N_4576,N_4324,N_4223);
nor U4577 (N_4577,N_4279,N_4373);
xnor U4578 (N_4578,N_4339,N_4274);
nor U4579 (N_4579,N_4356,N_4392);
nand U4580 (N_4580,N_4356,N_4397);
nand U4581 (N_4581,N_4262,N_4331);
nor U4582 (N_4582,N_4240,N_4362);
xor U4583 (N_4583,N_4246,N_4240);
xnor U4584 (N_4584,N_4305,N_4250);
nand U4585 (N_4585,N_4380,N_4208);
nor U4586 (N_4586,N_4316,N_4397);
nand U4587 (N_4587,N_4306,N_4344);
nand U4588 (N_4588,N_4245,N_4312);
nor U4589 (N_4589,N_4397,N_4312);
and U4590 (N_4590,N_4326,N_4217);
and U4591 (N_4591,N_4385,N_4380);
nand U4592 (N_4592,N_4335,N_4254);
nor U4593 (N_4593,N_4313,N_4251);
nand U4594 (N_4594,N_4311,N_4291);
and U4595 (N_4595,N_4380,N_4289);
and U4596 (N_4596,N_4217,N_4310);
nand U4597 (N_4597,N_4327,N_4224);
or U4598 (N_4598,N_4397,N_4215);
xnor U4599 (N_4599,N_4386,N_4233);
or U4600 (N_4600,N_4494,N_4542);
and U4601 (N_4601,N_4517,N_4401);
and U4602 (N_4602,N_4483,N_4468);
or U4603 (N_4603,N_4478,N_4546);
xor U4604 (N_4604,N_4568,N_4564);
nor U4605 (N_4605,N_4405,N_4411);
xnor U4606 (N_4606,N_4554,N_4524);
or U4607 (N_4607,N_4578,N_4558);
nor U4608 (N_4608,N_4476,N_4422);
or U4609 (N_4609,N_4572,N_4406);
xor U4610 (N_4610,N_4510,N_4444);
nor U4611 (N_4611,N_4427,N_4414);
nand U4612 (N_4612,N_4471,N_4532);
or U4613 (N_4613,N_4421,N_4435);
or U4614 (N_4614,N_4512,N_4434);
nor U4615 (N_4615,N_4561,N_4570);
nand U4616 (N_4616,N_4563,N_4553);
nand U4617 (N_4617,N_4590,N_4430);
xor U4618 (N_4618,N_4433,N_4449);
xnor U4619 (N_4619,N_4456,N_4577);
xnor U4620 (N_4620,N_4534,N_4574);
xnor U4621 (N_4621,N_4453,N_4519);
nand U4622 (N_4622,N_4598,N_4556);
xnor U4623 (N_4623,N_4535,N_4596);
nor U4624 (N_4624,N_4562,N_4423);
nor U4625 (N_4625,N_4439,N_4420);
nor U4626 (N_4626,N_4417,N_4486);
xnor U4627 (N_4627,N_4436,N_4429);
nand U4628 (N_4628,N_4593,N_4549);
and U4629 (N_4629,N_4543,N_4402);
xnor U4630 (N_4630,N_4432,N_4492);
xnor U4631 (N_4631,N_4477,N_4560);
or U4632 (N_4632,N_4567,N_4509);
or U4633 (N_4633,N_4413,N_4465);
and U4634 (N_4634,N_4499,N_4573);
or U4635 (N_4635,N_4475,N_4464);
xnor U4636 (N_4636,N_4498,N_4585);
or U4637 (N_4637,N_4511,N_4576);
nand U4638 (N_4638,N_4559,N_4502);
xnor U4639 (N_4639,N_4438,N_4548);
nand U4640 (N_4640,N_4536,N_4599);
xnor U4641 (N_4641,N_4595,N_4527);
xnor U4642 (N_4642,N_4550,N_4579);
nor U4643 (N_4643,N_4592,N_4445);
nor U4644 (N_4644,N_4426,N_4505);
nand U4645 (N_4645,N_4523,N_4407);
nand U4646 (N_4646,N_4516,N_4552);
and U4647 (N_4647,N_4479,N_4481);
and U4648 (N_4648,N_4533,N_4467);
nor U4649 (N_4649,N_4480,N_4518);
nand U4650 (N_4650,N_4591,N_4522);
nor U4651 (N_4651,N_4493,N_4501);
and U4652 (N_4652,N_4461,N_4412);
or U4653 (N_4653,N_4428,N_4525);
nor U4654 (N_4654,N_4544,N_4540);
and U4655 (N_4655,N_4587,N_4555);
nand U4656 (N_4656,N_4419,N_4557);
nor U4657 (N_4657,N_4504,N_4404);
xnor U4658 (N_4658,N_4490,N_4500);
nand U4659 (N_4659,N_4581,N_4495);
or U4660 (N_4660,N_4400,N_4448);
and U4661 (N_4661,N_4582,N_4425);
or U4662 (N_4662,N_4447,N_4459);
and U4663 (N_4663,N_4569,N_4586);
nand U4664 (N_4664,N_4487,N_4529);
nand U4665 (N_4665,N_4489,N_4450);
or U4666 (N_4666,N_4455,N_4463);
nand U4667 (N_4667,N_4474,N_4496);
and U4668 (N_4668,N_4528,N_4431);
xnor U4669 (N_4669,N_4485,N_4442);
or U4670 (N_4670,N_4488,N_4520);
nor U4671 (N_4671,N_4583,N_4537);
nor U4672 (N_4672,N_4441,N_4508);
nand U4673 (N_4673,N_4462,N_4515);
nor U4674 (N_4674,N_4513,N_4403);
nand U4675 (N_4675,N_4458,N_4589);
and U4676 (N_4676,N_4443,N_4457);
xor U4677 (N_4677,N_4526,N_4482);
nor U4678 (N_4678,N_4588,N_4521);
nor U4679 (N_4679,N_4424,N_4539);
or U4680 (N_4680,N_4418,N_4415);
nand U4681 (N_4681,N_4531,N_4454);
xnor U4682 (N_4682,N_4597,N_4446);
xnor U4683 (N_4683,N_4507,N_4547);
and U4684 (N_4684,N_4452,N_4408);
xor U4685 (N_4685,N_4571,N_4473);
nor U4686 (N_4686,N_4409,N_4551);
nand U4687 (N_4687,N_4484,N_4503);
xnor U4688 (N_4688,N_4594,N_4470);
or U4689 (N_4689,N_4541,N_4566);
nand U4690 (N_4690,N_4410,N_4565);
nand U4691 (N_4691,N_4437,N_4530);
nor U4692 (N_4692,N_4491,N_4497);
nor U4693 (N_4693,N_4440,N_4584);
xor U4694 (N_4694,N_4514,N_4580);
nand U4695 (N_4695,N_4460,N_4506);
and U4696 (N_4696,N_4545,N_4575);
nand U4697 (N_4697,N_4416,N_4472);
nand U4698 (N_4698,N_4466,N_4538);
or U4699 (N_4699,N_4451,N_4469);
xor U4700 (N_4700,N_4472,N_4468);
or U4701 (N_4701,N_4473,N_4407);
or U4702 (N_4702,N_4406,N_4455);
and U4703 (N_4703,N_4477,N_4468);
nand U4704 (N_4704,N_4584,N_4521);
and U4705 (N_4705,N_4430,N_4574);
or U4706 (N_4706,N_4576,N_4435);
nand U4707 (N_4707,N_4414,N_4445);
and U4708 (N_4708,N_4432,N_4405);
or U4709 (N_4709,N_4568,N_4550);
nor U4710 (N_4710,N_4558,N_4511);
nor U4711 (N_4711,N_4544,N_4480);
nand U4712 (N_4712,N_4565,N_4512);
nor U4713 (N_4713,N_4419,N_4578);
xnor U4714 (N_4714,N_4487,N_4485);
xor U4715 (N_4715,N_4524,N_4446);
or U4716 (N_4716,N_4564,N_4580);
xnor U4717 (N_4717,N_4436,N_4557);
nor U4718 (N_4718,N_4544,N_4534);
xor U4719 (N_4719,N_4551,N_4453);
nand U4720 (N_4720,N_4586,N_4595);
nand U4721 (N_4721,N_4518,N_4535);
nor U4722 (N_4722,N_4457,N_4432);
nand U4723 (N_4723,N_4446,N_4589);
and U4724 (N_4724,N_4596,N_4568);
xnor U4725 (N_4725,N_4490,N_4482);
nand U4726 (N_4726,N_4574,N_4441);
nor U4727 (N_4727,N_4512,N_4540);
and U4728 (N_4728,N_4533,N_4446);
or U4729 (N_4729,N_4431,N_4454);
nor U4730 (N_4730,N_4462,N_4416);
xor U4731 (N_4731,N_4420,N_4481);
nand U4732 (N_4732,N_4489,N_4468);
nor U4733 (N_4733,N_4433,N_4532);
and U4734 (N_4734,N_4405,N_4422);
xor U4735 (N_4735,N_4482,N_4541);
or U4736 (N_4736,N_4483,N_4456);
nand U4737 (N_4737,N_4411,N_4585);
nand U4738 (N_4738,N_4569,N_4441);
or U4739 (N_4739,N_4521,N_4556);
nor U4740 (N_4740,N_4512,N_4508);
nand U4741 (N_4741,N_4488,N_4503);
nand U4742 (N_4742,N_4538,N_4547);
nand U4743 (N_4743,N_4417,N_4491);
nor U4744 (N_4744,N_4563,N_4440);
nor U4745 (N_4745,N_4537,N_4403);
xnor U4746 (N_4746,N_4452,N_4413);
nor U4747 (N_4747,N_4595,N_4546);
xor U4748 (N_4748,N_4554,N_4430);
nand U4749 (N_4749,N_4496,N_4478);
nor U4750 (N_4750,N_4482,N_4500);
and U4751 (N_4751,N_4424,N_4541);
or U4752 (N_4752,N_4553,N_4485);
and U4753 (N_4753,N_4500,N_4532);
nand U4754 (N_4754,N_4563,N_4455);
nor U4755 (N_4755,N_4471,N_4445);
or U4756 (N_4756,N_4536,N_4479);
xor U4757 (N_4757,N_4556,N_4536);
or U4758 (N_4758,N_4418,N_4544);
nor U4759 (N_4759,N_4561,N_4500);
nor U4760 (N_4760,N_4565,N_4425);
or U4761 (N_4761,N_4476,N_4441);
nor U4762 (N_4762,N_4413,N_4444);
xor U4763 (N_4763,N_4590,N_4543);
nand U4764 (N_4764,N_4570,N_4548);
nor U4765 (N_4765,N_4565,N_4596);
nor U4766 (N_4766,N_4595,N_4569);
nor U4767 (N_4767,N_4567,N_4417);
or U4768 (N_4768,N_4491,N_4586);
and U4769 (N_4769,N_4468,N_4561);
xnor U4770 (N_4770,N_4514,N_4597);
nor U4771 (N_4771,N_4519,N_4469);
nand U4772 (N_4772,N_4449,N_4485);
nand U4773 (N_4773,N_4441,N_4430);
or U4774 (N_4774,N_4446,N_4430);
or U4775 (N_4775,N_4446,N_4458);
or U4776 (N_4776,N_4403,N_4400);
and U4777 (N_4777,N_4446,N_4448);
or U4778 (N_4778,N_4562,N_4406);
nand U4779 (N_4779,N_4479,N_4408);
xnor U4780 (N_4780,N_4567,N_4451);
nor U4781 (N_4781,N_4458,N_4513);
xor U4782 (N_4782,N_4569,N_4537);
or U4783 (N_4783,N_4553,N_4427);
nor U4784 (N_4784,N_4444,N_4598);
nand U4785 (N_4785,N_4588,N_4511);
xnor U4786 (N_4786,N_4497,N_4405);
nand U4787 (N_4787,N_4576,N_4468);
nor U4788 (N_4788,N_4462,N_4411);
nand U4789 (N_4789,N_4530,N_4568);
nor U4790 (N_4790,N_4590,N_4491);
xnor U4791 (N_4791,N_4545,N_4599);
xnor U4792 (N_4792,N_4591,N_4478);
or U4793 (N_4793,N_4546,N_4441);
nand U4794 (N_4794,N_4560,N_4481);
xor U4795 (N_4795,N_4564,N_4599);
nand U4796 (N_4796,N_4402,N_4435);
nor U4797 (N_4797,N_4548,N_4544);
and U4798 (N_4798,N_4474,N_4493);
or U4799 (N_4799,N_4415,N_4401);
or U4800 (N_4800,N_4674,N_4637);
nand U4801 (N_4801,N_4729,N_4740);
xor U4802 (N_4802,N_4624,N_4697);
nor U4803 (N_4803,N_4774,N_4645);
or U4804 (N_4804,N_4616,N_4696);
nand U4805 (N_4805,N_4601,N_4709);
nor U4806 (N_4806,N_4736,N_4606);
xnor U4807 (N_4807,N_4660,N_4786);
or U4808 (N_4808,N_4632,N_4742);
nor U4809 (N_4809,N_4627,N_4661);
nand U4810 (N_4810,N_4704,N_4698);
and U4811 (N_4811,N_4775,N_4779);
nand U4812 (N_4812,N_4600,N_4793);
xor U4813 (N_4813,N_4751,N_4630);
nand U4814 (N_4814,N_4728,N_4650);
or U4815 (N_4815,N_4790,N_4799);
and U4816 (N_4816,N_4602,N_4769);
nor U4817 (N_4817,N_4668,N_4703);
nor U4818 (N_4818,N_4721,N_4699);
nand U4819 (N_4819,N_4764,N_4797);
and U4820 (N_4820,N_4665,N_4663);
nor U4821 (N_4821,N_4615,N_4628);
xor U4822 (N_4822,N_4675,N_4792);
nand U4823 (N_4823,N_4622,N_4691);
or U4824 (N_4824,N_4684,N_4765);
nor U4825 (N_4825,N_4755,N_4784);
nand U4826 (N_4826,N_4763,N_4744);
or U4827 (N_4827,N_4638,N_4688);
nand U4828 (N_4828,N_4682,N_4727);
and U4829 (N_4829,N_4648,N_4679);
nand U4830 (N_4830,N_4635,N_4646);
nor U4831 (N_4831,N_4634,N_4772);
nor U4832 (N_4832,N_4641,N_4778);
nor U4833 (N_4833,N_4730,N_4748);
or U4834 (N_4834,N_4702,N_4692);
nand U4835 (N_4835,N_4644,N_4604);
or U4836 (N_4836,N_4788,N_4771);
nor U4837 (N_4837,N_4655,N_4656);
or U4838 (N_4838,N_4724,N_4794);
and U4839 (N_4839,N_4658,N_4700);
xor U4840 (N_4840,N_4780,N_4617);
nand U4841 (N_4841,N_4678,N_4666);
nand U4842 (N_4842,N_4783,N_4796);
xnor U4843 (N_4843,N_4732,N_4749);
nand U4844 (N_4844,N_4685,N_4639);
nand U4845 (N_4845,N_4714,N_4762);
nor U4846 (N_4846,N_4680,N_4777);
nand U4847 (N_4847,N_4670,N_4652);
nand U4848 (N_4848,N_4618,N_4647);
xor U4849 (N_4849,N_4686,N_4687);
nor U4850 (N_4850,N_4757,N_4766);
nand U4851 (N_4851,N_4695,N_4669);
nor U4852 (N_4852,N_4723,N_4657);
nand U4853 (N_4853,N_4613,N_4693);
nand U4854 (N_4854,N_4654,N_4708);
and U4855 (N_4855,N_4776,N_4725);
and U4856 (N_4856,N_4689,N_4629);
nand U4857 (N_4857,N_4718,N_4754);
and U4858 (N_4858,N_4798,N_4651);
nor U4859 (N_4859,N_4739,N_4672);
xnor U4860 (N_4860,N_4712,N_4734);
and U4861 (N_4861,N_4713,N_4760);
and U4862 (N_4862,N_4620,N_4640);
nand U4863 (N_4863,N_4789,N_4741);
xor U4864 (N_4864,N_4753,N_4717);
nand U4865 (N_4865,N_4770,N_4731);
and U4866 (N_4866,N_4773,N_4694);
and U4867 (N_4867,N_4608,N_4738);
nor U4868 (N_4868,N_4625,N_4611);
and U4869 (N_4869,N_4715,N_4759);
xnor U4870 (N_4870,N_4610,N_4683);
nand U4871 (N_4871,N_4720,N_4706);
nor U4872 (N_4872,N_4756,N_4782);
or U4873 (N_4873,N_4726,N_4653);
nand U4874 (N_4874,N_4667,N_4671);
and U4875 (N_4875,N_4609,N_4791);
and U4876 (N_4876,N_4623,N_4642);
and U4877 (N_4877,N_4636,N_4643);
or U4878 (N_4878,N_4735,N_4752);
nand U4879 (N_4879,N_4711,N_4612);
nor U4880 (N_4880,N_4722,N_4705);
nand U4881 (N_4881,N_4649,N_4710);
and U4882 (N_4882,N_4690,N_4745);
nand U4883 (N_4883,N_4716,N_4676);
xnor U4884 (N_4884,N_4781,N_4719);
or U4885 (N_4885,N_4787,N_4664);
and U4886 (N_4886,N_4733,N_4631);
and U4887 (N_4887,N_4677,N_4614);
and U4888 (N_4888,N_4750,N_4681);
nand U4889 (N_4889,N_4659,N_4737);
nor U4890 (N_4890,N_4747,N_4673);
and U4891 (N_4891,N_4746,N_4621);
xnor U4892 (N_4892,N_4603,N_4761);
nand U4893 (N_4893,N_4619,N_4785);
and U4894 (N_4894,N_4795,N_4607);
nand U4895 (N_4895,N_4768,N_4605);
or U4896 (N_4896,N_4743,N_4701);
xnor U4897 (N_4897,N_4626,N_4633);
nand U4898 (N_4898,N_4767,N_4707);
nand U4899 (N_4899,N_4758,N_4662);
nand U4900 (N_4900,N_4657,N_4719);
nor U4901 (N_4901,N_4715,N_4701);
nor U4902 (N_4902,N_4616,N_4722);
or U4903 (N_4903,N_4678,N_4630);
and U4904 (N_4904,N_4708,N_4670);
xnor U4905 (N_4905,N_4676,N_4786);
nor U4906 (N_4906,N_4652,N_4647);
nand U4907 (N_4907,N_4753,N_4798);
or U4908 (N_4908,N_4725,N_4710);
xor U4909 (N_4909,N_4654,N_4637);
or U4910 (N_4910,N_4651,N_4677);
nor U4911 (N_4911,N_4703,N_4652);
nor U4912 (N_4912,N_4772,N_4631);
nand U4913 (N_4913,N_4668,N_4600);
nand U4914 (N_4914,N_4759,N_4679);
nor U4915 (N_4915,N_4703,N_4741);
nand U4916 (N_4916,N_4655,N_4609);
and U4917 (N_4917,N_4618,N_4705);
or U4918 (N_4918,N_4662,N_4647);
xnor U4919 (N_4919,N_4796,N_4688);
or U4920 (N_4920,N_4712,N_4631);
or U4921 (N_4921,N_4667,N_4791);
nand U4922 (N_4922,N_4759,N_4766);
xor U4923 (N_4923,N_4744,N_4601);
nand U4924 (N_4924,N_4674,N_4780);
or U4925 (N_4925,N_4786,N_4726);
nor U4926 (N_4926,N_4611,N_4718);
nand U4927 (N_4927,N_4737,N_4660);
nand U4928 (N_4928,N_4659,N_4650);
and U4929 (N_4929,N_4654,N_4672);
nand U4930 (N_4930,N_4754,N_4750);
xnor U4931 (N_4931,N_4786,N_4637);
nor U4932 (N_4932,N_4640,N_4617);
xnor U4933 (N_4933,N_4699,N_4658);
nor U4934 (N_4934,N_4614,N_4635);
nand U4935 (N_4935,N_4792,N_4641);
or U4936 (N_4936,N_4652,N_4765);
or U4937 (N_4937,N_4760,N_4772);
xnor U4938 (N_4938,N_4710,N_4617);
or U4939 (N_4939,N_4736,N_4747);
and U4940 (N_4940,N_4753,N_4752);
nor U4941 (N_4941,N_4682,N_4738);
nor U4942 (N_4942,N_4741,N_4650);
xor U4943 (N_4943,N_4606,N_4742);
nor U4944 (N_4944,N_4748,N_4701);
nand U4945 (N_4945,N_4714,N_4766);
nor U4946 (N_4946,N_4739,N_4753);
or U4947 (N_4947,N_4773,N_4745);
nor U4948 (N_4948,N_4716,N_4678);
or U4949 (N_4949,N_4749,N_4784);
and U4950 (N_4950,N_4759,N_4633);
nand U4951 (N_4951,N_4638,N_4600);
nor U4952 (N_4952,N_4742,N_4601);
nor U4953 (N_4953,N_4689,N_4703);
nand U4954 (N_4954,N_4764,N_4682);
nor U4955 (N_4955,N_4776,N_4693);
and U4956 (N_4956,N_4709,N_4772);
or U4957 (N_4957,N_4651,N_4627);
nand U4958 (N_4958,N_4721,N_4617);
and U4959 (N_4959,N_4717,N_4792);
xnor U4960 (N_4960,N_4692,N_4760);
and U4961 (N_4961,N_4608,N_4785);
nand U4962 (N_4962,N_4754,N_4747);
xnor U4963 (N_4963,N_4794,N_4798);
xor U4964 (N_4964,N_4688,N_4774);
nand U4965 (N_4965,N_4772,N_4619);
xnor U4966 (N_4966,N_4647,N_4691);
nand U4967 (N_4967,N_4780,N_4728);
or U4968 (N_4968,N_4615,N_4623);
and U4969 (N_4969,N_4790,N_4787);
nor U4970 (N_4970,N_4685,N_4628);
nor U4971 (N_4971,N_4664,N_4649);
or U4972 (N_4972,N_4634,N_4666);
nor U4973 (N_4973,N_4668,N_4740);
nor U4974 (N_4974,N_4776,N_4782);
or U4975 (N_4975,N_4623,N_4718);
nand U4976 (N_4976,N_4644,N_4726);
xor U4977 (N_4977,N_4744,N_4623);
xor U4978 (N_4978,N_4700,N_4665);
xnor U4979 (N_4979,N_4739,N_4634);
nand U4980 (N_4980,N_4613,N_4783);
nand U4981 (N_4981,N_4759,N_4796);
and U4982 (N_4982,N_4661,N_4625);
or U4983 (N_4983,N_4797,N_4611);
nor U4984 (N_4984,N_4634,N_4707);
nand U4985 (N_4985,N_4694,N_4727);
and U4986 (N_4986,N_4748,N_4789);
or U4987 (N_4987,N_4793,N_4735);
xor U4988 (N_4988,N_4727,N_4684);
nand U4989 (N_4989,N_4788,N_4684);
and U4990 (N_4990,N_4625,N_4653);
nor U4991 (N_4991,N_4600,N_4690);
nand U4992 (N_4992,N_4726,N_4611);
xor U4993 (N_4993,N_4775,N_4663);
and U4994 (N_4994,N_4691,N_4786);
nand U4995 (N_4995,N_4735,N_4608);
xor U4996 (N_4996,N_4620,N_4664);
nor U4997 (N_4997,N_4766,N_4698);
nor U4998 (N_4998,N_4649,N_4754);
or U4999 (N_4999,N_4720,N_4721);
and U5000 (N_5000,N_4803,N_4854);
nor U5001 (N_5001,N_4892,N_4853);
nor U5002 (N_5002,N_4997,N_4889);
xnor U5003 (N_5003,N_4828,N_4888);
nor U5004 (N_5004,N_4863,N_4934);
or U5005 (N_5005,N_4847,N_4914);
nor U5006 (N_5006,N_4910,N_4984);
or U5007 (N_5007,N_4840,N_4965);
or U5008 (N_5008,N_4820,N_4981);
xor U5009 (N_5009,N_4931,N_4895);
xor U5010 (N_5010,N_4839,N_4806);
or U5011 (N_5011,N_4845,N_4979);
and U5012 (N_5012,N_4868,N_4901);
nand U5013 (N_5013,N_4831,N_4825);
xor U5014 (N_5014,N_4857,N_4954);
and U5015 (N_5015,N_4833,N_4841);
nand U5016 (N_5016,N_4826,N_4834);
xor U5017 (N_5017,N_4809,N_4813);
xor U5018 (N_5018,N_4844,N_4960);
nor U5019 (N_5019,N_4987,N_4913);
and U5020 (N_5020,N_4842,N_4969);
nor U5021 (N_5021,N_4909,N_4911);
nand U5022 (N_5022,N_4993,N_4881);
xor U5023 (N_5023,N_4967,N_4862);
and U5024 (N_5024,N_4922,N_4885);
or U5025 (N_5025,N_4898,N_4933);
or U5026 (N_5026,N_4947,N_4973);
or U5027 (N_5027,N_4968,N_4900);
xor U5028 (N_5028,N_4991,N_4985);
xnor U5029 (N_5029,N_4986,N_4812);
or U5030 (N_5030,N_4927,N_4938);
nand U5031 (N_5031,N_4821,N_4975);
nor U5032 (N_5032,N_4816,N_4846);
nand U5033 (N_5033,N_4920,N_4958);
nand U5034 (N_5034,N_4866,N_4830);
xnor U5035 (N_5035,N_4930,N_4849);
and U5036 (N_5036,N_4959,N_4990);
nor U5037 (N_5037,N_4891,N_4971);
and U5038 (N_5038,N_4872,N_4835);
nor U5039 (N_5039,N_4893,N_4869);
nand U5040 (N_5040,N_4867,N_4808);
xor U5041 (N_5041,N_4887,N_4980);
xnor U5042 (N_5042,N_4977,N_4929);
xnor U5043 (N_5043,N_4874,N_4878);
nand U5044 (N_5044,N_4858,N_4961);
xor U5045 (N_5045,N_4884,N_4957);
xnor U5046 (N_5046,N_4996,N_4917);
and U5047 (N_5047,N_4848,N_4902);
nor U5048 (N_5048,N_4836,N_4951);
nand U5049 (N_5049,N_4877,N_4906);
nor U5050 (N_5050,N_4948,N_4880);
nor U5051 (N_5051,N_4811,N_4800);
nor U5052 (N_5052,N_4974,N_4810);
or U5053 (N_5053,N_4864,N_4861);
nand U5054 (N_5054,N_4832,N_4890);
nor U5055 (N_5055,N_4804,N_4970);
and U5056 (N_5056,N_4817,N_4897);
xnor U5057 (N_5057,N_4851,N_4972);
or U5058 (N_5058,N_4903,N_4838);
nor U5059 (N_5059,N_4964,N_4807);
nand U5060 (N_5060,N_4956,N_4989);
and U5061 (N_5061,N_4915,N_4801);
nand U5062 (N_5062,N_4870,N_4945);
nand U5063 (N_5063,N_4827,N_4994);
and U5064 (N_5064,N_4805,N_4963);
xor U5065 (N_5065,N_4998,N_4924);
xnor U5066 (N_5066,N_4925,N_4935);
xnor U5067 (N_5067,N_4871,N_4982);
and U5068 (N_5068,N_4926,N_4999);
or U5069 (N_5069,N_4949,N_4823);
nand U5070 (N_5070,N_4941,N_4946);
nor U5071 (N_5071,N_4882,N_4995);
and U5072 (N_5072,N_4937,N_4876);
nand U5073 (N_5073,N_4904,N_4802);
nor U5074 (N_5074,N_4992,N_4978);
or U5075 (N_5075,N_4905,N_4837);
nor U5076 (N_5076,N_4916,N_4883);
nor U5077 (N_5077,N_4983,N_4875);
nor U5078 (N_5078,N_4952,N_4943);
nor U5079 (N_5079,N_4856,N_4886);
or U5080 (N_5080,N_4950,N_4944);
and U5081 (N_5081,N_4815,N_4908);
nand U5082 (N_5082,N_4936,N_4814);
or U5083 (N_5083,N_4918,N_4859);
nand U5084 (N_5084,N_4829,N_4919);
xnor U5085 (N_5085,N_4824,N_4899);
xnor U5086 (N_5086,N_4928,N_4940);
xnor U5087 (N_5087,N_4923,N_4819);
xor U5088 (N_5088,N_4879,N_4850);
nand U5089 (N_5089,N_4921,N_4896);
or U5090 (N_5090,N_4907,N_4843);
or U5091 (N_5091,N_4865,N_4912);
nor U5092 (N_5092,N_4988,N_4939);
nand U5093 (N_5093,N_4818,N_4953);
and U5094 (N_5094,N_4932,N_4966);
and U5095 (N_5095,N_4962,N_4894);
or U5096 (N_5096,N_4955,N_4942);
and U5097 (N_5097,N_4822,N_4873);
or U5098 (N_5098,N_4860,N_4855);
and U5099 (N_5099,N_4852,N_4976);
nor U5100 (N_5100,N_4855,N_4923);
and U5101 (N_5101,N_4971,N_4869);
xor U5102 (N_5102,N_4845,N_4869);
nand U5103 (N_5103,N_4884,N_4931);
xor U5104 (N_5104,N_4908,N_4988);
nor U5105 (N_5105,N_4915,N_4965);
nand U5106 (N_5106,N_4881,N_4914);
nor U5107 (N_5107,N_4883,N_4888);
nor U5108 (N_5108,N_4834,N_4863);
nand U5109 (N_5109,N_4868,N_4858);
xor U5110 (N_5110,N_4900,N_4800);
or U5111 (N_5111,N_4893,N_4828);
nand U5112 (N_5112,N_4811,N_4969);
nand U5113 (N_5113,N_4954,N_4903);
or U5114 (N_5114,N_4851,N_4886);
nand U5115 (N_5115,N_4826,N_4925);
and U5116 (N_5116,N_4895,N_4960);
nand U5117 (N_5117,N_4920,N_4815);
xnor U5118 (N_5118,N_4917,N_4929);
and U5119 (N_5119,N_4961,N_4812);
or U5120 (N_5120,N_4807,N_4847);
or U5121 (N_5121,N_4906,N_4802);
nor U5122 (N_5122,N_4918,N_4995);
xor U5123 (N_5123,N_4897,N_4805);
and U5124 (N_5124,N_4948,N_4938);
or U5125 (N_5125,N_4837,N_4801);
and U5126 (N_5126,N_4809,N_4832);
or U5127 (N_5127,N_4827,N_4902);
xnor U5128 (N_5128,N_4804,N_4822);
nand U5129 (N_5129,N_4988,N_4930);
nor U5130 (N_5130,N_4970,N_4921);
nand U5131 (N_5131,N_4998,N_4870);
or U5132 (N_5132,N_4942,N_4838);
and U5133 (N_5133,N_4962,N_4848);
nand U5134 (N_5134,N_4977,N_4895);
and U5135 (N_5135,N_4891,N_4825);
and U5136 (N_5136,N_4824,N_4982);
nand U5137 (N_5137,N_4912,N_4823);
or U5138 (N_5138,N_4967,N_4847);
xor U5139 (N_5139,N_4898,N_4868);
or U5140 (N_5140,N_4855,N_4862);
nor U5141 (N_5141,N_4961,N_4878);
nor U5142 (N_5142,N_4861,N_4974);
nor U5143 (N_5143,N_4895,N_4962);
and U5144 (N_5144,N_4932,N_4905);
or U5145 (N_5145,N_4810,N_4973);
nand U5146 (N_5146,N_4816,N_4890);
or U5147 (N_5147,N_4981,N_4951);
nor U5148 (N_5148,N_4901,N_4909);
nor U5149 (N_5149,N_4956,N_4801);
or U5150 (N_5150,N_4966,N_4956);
or U5151 (N_5151,N_4976,N_4953);
nor U5152 (N_5152,N_4896,N_4968);
nor U5153 (N_5153,N_4816,N_4822);
xor U5154 (N_5154,N_4951,N_4923);
xnor U5155 (N_5155,N_4824,N_4871);
nor U5156 (N_5156,N_4930,N_4874);
and U5157 (N_5157,N_4896,N_4853);
xor U5158 (N_5158,N_4939,N_4819);
xor U5159 (N_5159,N_4974,N_4892);
nor U5160 (N_5160,N_4919,N_4870);
nand U5161 (N_5161,N_4919,N_4964);
nor U5162 (N_5162,N_4879,N_4873);
nand U5163 (N_5163,N_4876,N_4963);
nand U5164 (N_5164,N_4892,N_4801);
nand U5165 (N_5165,N_4907,N_4973);
nand U5166 (N_5166,N_4873,N_4990);
nor U5167 (N_5167,N_4856,N_4843);
or U5168 (N_5168,N_4965,N_4851);
nor U5169 (N_5169,N_4818,N_4873);
xor U5170 (N_5170,N_4930,N_4941);
xor U5171 (N_5171,N_4995,N_4977);
xor U5172 (N_5172,N_4897,N_4927);
or U5173 (N_5173,N_4943,N_4807);
nand U5174 (N_5174,N_4946,N_4885);
xor U5175 (N_5175,N_4890,N_4838);
xor U5176 (N_5176,N_4886,N_4966);
xnor U5177 (N_5177,N_4944,N_4887);
nor U5178 (N_5178,N_4845,N_4935);
xor U5179 (N_5179,N_4982,N_4998);
or U5180 (N_5180,N_4866,N_4860);
and U5181 (N_5181,N_4808,N_4955);
xor U5182 (N_5182,N_4807,N_4882);
or U5183 (N_5183,N_4958,N_4971);
and U5184 (N_5184,N_4815,N_4917);
nor U5185 (N_5185,N_4945,N_4984);
nand U5186 (N_5186,N_4870,N_4990);
xnor U5187 (N_5187,N_4920,N_4938);
or U5188 (N_5188,N_4846,N_4977);
xor U5189 (N_5189,N_4843,N_4922);
xnor U5190 (N_5190,N_4821,N_4866);
xnor U5191 (N_5191,N_4864,N_4860);
and U5192 (N_5192,N_4878,N_4991);
nand U5193 (N_5193,N_4877,N_4807);
nand U5194 (N_5194,N_4977,N_4928);
or U5195 (N_5195,N_4807,N_4988);
nor U5196 (N_5196,N_4898,N_4956);
or U5197 (N_5197,N_4906,N_4814);
nand U5198 (N_5198,N_4868,N_4940);
nand U5199 (N_5199,N_4928,N_4911);
nand U5200 (N_5200,N_5136,N_5135);
nand U5201 (N_5201,N_5065,N_5055);
and U5202 (N_5202,N_5025,N_5153);
nor U5203 (N_5203,N_5035,N_5163);
or U5204 (N_5204,N_5124,N_5054);
or U5205 (N_5205,N_5062,N_5178);
xnor U5206 (N_5206,N_5121,N_5004);
or U5207 (N_5207,N_5097,N_5043);
nor U5208 (N_5208,N_5018,N_5078);
or U5209 (N_5209,N_5074,N_5028);
xnor U5210 (N_5210,N_5137,N_5128);
nor U5211 (N_5211,N_5016,N_5014);
or U5212 (N_5212,N_5113,N_5030);
or U5213 (N_5213,N_5131,N_5172);
xor U5214 (N_5214,N_5002,N_5126);
and U5215 (N_5215,N_5051,N_5185);
nand U5216 (N_5216,N_5129,N_5081);
xnor U5217 (N_5217,N_5053,N_5157);
and U5218 (N_5218,N_5063,N_5104);
xnor U5219 (N_5219,N_5156,N_5120);
nor U5220 (N_5220,N_5099,N_5125);
nor U5221 (N_5221,N_5013,N_5106);
or U5222 (N_5222,N_5031,N_5132);
xor U5223 (N_5223,N_5006,N_5039);
or U5224 (N_5224,N_5034,N_5161);
xor U5225 (N_5225,N_5147,N_5015);
and U5226 (N_5226,N_5189,N_5007);
or U5227 (N_5227,N_5042,N_5045);
and U5228 (N_5228,N_5192,N_5168);
nand U5229 (N_5229,N_5008,N_5079);
nand U5230 (N_5230,N_5038,N_5117);
or U5231 (N_5231,N_5020,N_5023);
and U5232 (N_5232,N_5155,N_5101);
xnor U5233 (N_5233,N_5159,N_5057);
or U5234 (N_5234,N_5198,N_5102);
nand U5235 (N_5235,N_5105,N_5027);
nand U5236 (N_5236,N_5067,N_5010);
xor U5237 (N_5237,N_5180,N_5096);
or U5238 (N_5238,N_5108,N_5177);
nor U5239 (N_5239,N_5071,N_5139);
xnor U5240 (N_5240,N_5036,N_5093);
xor U5241 (N_5241,N_5184,N_5083);
nor U5242 (N_5242,N_5060,N_5176);
and U5243 (N_5243,N_5114,N_5050);
or U5244 (N_5244,N_5085,N_5087);
or U5245 (N_5245,N_5151,N_5024);
nor U5246 (N_5246,N_5044,N_5009);
and U5247 (N_5247,N_5070,N_5100);
or U5248 (N_5248,N_5160,N_5032);
or U5249 (N_5249,N_5167,N_5092);
nand U5250 (N_5250,N_5191,N_5123);
nor U5251 (N_5251,N_5181,N_5149);
and U5252 (N_5252,N_5187,N_5186);
or U5253 (N_5253,N_5049,N_5047);
nand U5254 (N_5254,N_5143,N_5190);
nor U5255 (N_5255,N_5138,N_5154);
xor U5256 (N_5256,N_5072,N_5111);
nand U5257 (N_5257,N_5148,N_5182);
nand U5258 (N_5258,N_5029,N_5166);
xor U5259 (N_5259,N_5130,N_5040);
xor U5260 (N_5260,N_5011,N_5173);
or U5261 (N_5261,N_5001,N_5077);
or U5262 (N_5262,N_5012,N_5076);
and U5263 (N_5263,N_5056,N_5158);
nand U5264 (N_5264,N_5066,N_5165);
nor U5265 (N_5265,N_5005,N_5115);
nand U5266 (N_5266,N_5086,N_5058);
nor U5267 (N_5267,N_5194,N_5145);
or U5268 (N_5268,N_5048,N_5174);
xnor U5269 (N_5269,N_5195,N_5134);
and U5270 (N_5270,N_5094,N_5082);
xnor U5271 (N_5271,N_5109,N_5084);
xor U5272 (N_5272,N_5119,N_5152);
or U5273 (N_5273,N_5122,N_5019);
nor U5274 (N_5274,N_5142,N_5197);
or U5275 (N_5275,N_5141,N_5162);
or U5276 (N_5276,N_5112,N_5059);
xor U5277 (N_5277,N_5026,N_5091);
xnor U5278 (N_5278,N_5033,N_5171);
nor U5279 (N_5279,N_5017,N_5144);
or U5280 (N_5280,N_5116,N_5000);
xnor U5281 (N_5281,N_5041,N_5069);
nor U5282 (N_5282,N_5169,N_5064);
and U5283 (N_5283,N_5068,N_5150);
or U5284 (N_5284,N_5080,N_5003);
nand U5285 (N_5285,N_5089,N_5021);
or U5286 (N_5286,N_5022,N_5188);
and U5287 (N_5287,N_5199,N_5196);
nand U5288 (N_5288,N_5118,N_5140);
nor U5289 (N_5289,N_5133,N_5103);
nor U5290 (N_5290,N_5095,N_5107);
nor U5291 (N_5291,N_5037,N_5164);
xor U5292 (N_5292,N_5179,N_5127);
nand U5293 (N_5293,N_5052,N_5170);
xnor U5294 (N_5294,N_5110,N_5090);
nor U5295 (N_5295,N_5098,N_5075);
nor U5296 (N_5296,N_5061,N_5193);
or U5297 (N_5297,N_5073,N_5146);
nor U5298 (N_5298,N_5183,N_5046);
nor U5299 (N_5299,N_5088,N_5175);
xnor U5300 (N_5300,N_5133,N_5197);
nand U5301 (N_5301,N_5062,N_5167);
nand U5302 (N_5302,N_5176,N_5071);
nand U5303 (N_5303,N_5195,N_5084);
nor U5304 (N_5304,N_5134,N_5071);
nand U5305 (N_5305,N_5166,N_5106);
or U5306 (N_5306,N_5185,N_5040);
and U5307 (N_5307,N_5014,N_5032);
xnor U5308 (N_5308,N_5046,N_5124);
or U5309 (N_5309,N_5089,N_5195);
nor U5310 (N_5310,N_5123,N_5028);
xor U5311 (N_5311,N_5060,N_5001);
and U5312 (N_5312,N_5115,N_5069);
or U5313 (N_5313,N_5119,N_5063);
xor U5314 (N_5314,N_5118,N_5113);
or U5315 (N_5315,N_5133,N_5089);
and U5316 (N_5316,N_5176,N_5094);
and U5317 (N_5317,N_5061,N_5196);
or U5318 (N_5318,N_5154,N_5050);
xor U5319 (N_5319,N_5099,N_5178);
and U5320 (N_5320,N_5160,N_5012);
nand U5321 (N_5321,N_5051,N_5000);
and U5322 (N_5322,N_5130,N_5193);
and U5323 (N_5323,N_5199,N_5101);
and U5324 (N_5324,N_5017,N_5053);
nand U5325 (N_5325,N_5093,N_5007);
nor U5326 (N_5326,N_5128,N_5089);
nor U5327 (N_5327,N_5172,N_5004);
and U5328 (N_5328,N_5149,N_5021);
or U5329 (N_5329,N_5176,N_5198);
xnor U5330 (N_5330,N_5067,N_5146);
or U5331 (N_5331,N_5149,N_5183);
nand U5332 (N_5332,N_5178,N_5132);
and U5333 (N_5333,N_5023,N_5071);
xnor U5334 (N_5334,N_5165,N_5006);
xor U5335 (N_5335,N_5027,N_5185);
xor U5336 (N_5336,N_5168,N_5048);
nand U5337 (N_5337,N_5066,N_5182);
xnor U5338 (N_5338,N_5137,N_5133);
nor U5339 (N_5339,N_5002,N_5186);
and U5340 (N_5340,N_5099,N_5087);
xnor U5341 (N_5341,N_5056,N_5068);
or U5342 (N_5342,N_5180,N_5128);
and U5343 (N_5343,N_5095,N_5152);
and U5344 (N_5344,N_5114,N_5045);
xor U5345 (N_5345,N_5033,N_5191);
xnor U5346 (N_5346,N_5012,N_5011);
and U5347 (N_5347,N_5061,N_5000);
nor U5348 (N_5348,N_5143,N_5117);
nor U5349 (N_5349,N_5148,N_5101);
nor U5350 (N_5350,N_5015,N_5105);
nor U5351 (N_5351,N_5015,N_5027);
or U5352 (N_5352,N_5195,N_5090);
and U5353 (N_5353,N_5178,N_5174);
xnor U5354 (N_5354,N_5079,N_5006);
nand U5355 (N_5355,N_5103,N_5173);
or U5356 (N_5356,N_5075,N_5017);
nor U5357 (N_5357,N_5044,N_5173);
nor U5358 (N_5358,N_5042,N_5022);
or U5359 (N_5359,N_5089,N_5007);
or U5360 (N_5360,N_5197,N_5042);
nand U5361 (N_5361,N_5029,N_5193);
nor U5362 (N_5362,N_5071,N_5099);
nand U5363 (N_5363,N_5053,N_5104);
or U5364 (N_5364,N_5195,N_5098);
nand U5365 (N_5365,N_5080,N_5089);
or U5366 (N_5366,N_5135,N_5016);
nor U5367 (N_5367,N_5162,N_5017);
nor U5368 (N_5368,N_5196,N_5008);
and U5369 (N_5369,N_5177,N_5181);
nor U5370 (N_5370,N_5004,N_5047);
nand U5371 (N_5371,N_5057,N_5104);
nand U5372 (N_5372,N_5175,N_5023);
or U5373 (N_5373,N_5067,N_5104);
xor U5374 (N_5374,N_5107,N_5173);
nor U5375 (N_5375,N_5075,N_5055);
xor U5376 (N_5376,N_5192,N_5171);
nand U5377 (N_5377,N_5003,N_5144);
nand U5378 (N_5378,N_5053,N_5046);
xnor U5379 (N_5379,N_5011,N_5002);
nand U5380 (N_5380,N_5105,N_5061);
or U5381 (N_5381,N_5095,N_5050);
and U5382 (N_5382,N_5014,N_5106);
xnor U5383 (N_5383,N_5168,N_5027);
or U5384 (N_5384,N_5167,N_5113);
nand U5385 (N_5385,N_5192,N_5117);
nand U5386 (N_5386,N_5119,N_5032);
nor U5387 (N_5387,N_5182,N_5058);
nand U5388 (N_5388,N_5027,N_5022);
xor U5389 (N_5389,N_5103,N_5098);
nand U5390 (N_5390,N_5173,N_5122);
xnor U5391 (N_5391,N_5194,N_5170);
nand U5392 (N_5392,N_5010,N_5137);
nand U5393 (N_5393,N_5033,N_5132);
nand U5394 (N_5394,N_5046,N_5132);
and U5395 (N_5395,N_5076,N_5067);
nand U5396 (N_5396,N_5047,N_5131);
xor U5397 (N_5397,N_5006,N_5120);
or U5398 (N_5398,N_5007,N_5158);
and U5399 (N_5399,N_5142,N_5079);
nor U5400 (N_5400,N_5284,N_5309);
xor U5401 (N_5401,N_5343,N_5337);
xor U5402 (N_5402,N_5237,N_5346);
xnor U5403 (N_5403,N_5204,N_5318);
or U5404 (N_5404,N_5290,N_5390);
nor U5405 (N_5405,N_5260,N_5271);
nor U5406 (N_5406,N_5366,N_5244);
and U5407 (N_5407,N_5396,N_5247);
and U5408 (N_5408,N_5211,N_5317);
and U5409 (N_5409,N_5328,N_5349);
or U5410 (N_5410,N_5327,N_5221);
and U5411 (N_5411,N_5388,N_5348);
nand U5412 (N_5412,N_5391,N_5339);
nand U5413 (N_5413,N_5262,N_5238);
nand U5414 (N_5414,N_5331,N_5340);
and U5415 (N_5415,N_5356,N_5389);
or U5416 (N_5416,N_5245,N_5202);
xor U5417 (N_5417,N_5278,N_5376);
or U5418 (N_5418,N_5341,N_5275);
nand U5419 (N_5419,N_5207,N_5297);
or U5420 (N_5420,N_5323,N_5293);
or U5421 (N_5421,N_5344,N_5399);
nor U5422 (N_5422,N_5321,N_5325);
and U5423 (N_5423,N_5315,N_5274);
nand U5424 (N_5424,N_5350,N_5234);
xor U5425 (N_5425,N_5217,N_5383);
or U5426 (N_5426,N_5258,N_5353);
and U5427 (N_5427,N_5364,N_5215);
nor U5428 (N_5428,N_5397,N_5283);
xor U5429 (N_5429,N_5392,N_5395);
and U5430 (N_5430,N_5254,N_5307);
nor U5431 (N_5431,N_5324,N_5312);
and U5432 (N_5432,N_5305,N_5285);
or U5433 (N_5433,N_5322,N_5259);
nand U5434 (N_5434,N_5226,N_5239);
nand U5435 (N_5435,N_5298,N_5250);
and U5436 (N_5436,N_5203,N_5256);
nand U5437 (N_5437,N_5304,N_5360);
nand U5438 (N_5438,N_5306,N_5357);
nor U5439 (N_5439,N_5378,N_5362);
xnor U5440 (N_5440,N_5288,N_5382);
nor U5441 (N_5441,N_5335,N_5381);
nor U5442 (N_5442,N_5205,N_5265);
nor U5443 (N_5443,N_5365,N_5264);
and U5444 (N_5444,N_5246,N_5329);
nand U5445 (N_5445,N_5374,N_5216);
nand U5446 (N_5446,N_5229,N_5233);
or U5447 (N_5447,N_5308,N_5279);
or U5448 (N_5448,N_5241,N_5330);
or U5449 (N_5449,N_5261,N_5345);
xnor U5450 (N_5450,N_5296,N_5319);
xor U5451 (N_5451,N_5352,N_5268);
nand U5452 (N_5452,N_5359,N_5387);
and U5453 (N_5453,N_5347,N_5252);
or U5454 (N_5454,N_5231,N_5295);
nor U5455 (N_5455,N_5266,N_5313);
xor U5456 (N_5456,N_5301,N_5379);
or U5457 (N_5457,N_5334,N_5257);
nor U5458 (N_5458,N_5363,N_5236);
nor U5459 (N_5459,N_5302,N_5372);
nand U5460 (N_5460,N_5227,N_5263);
nor U5461 (N_5461,N_5281,N_5303);
xor U5462 (N_5462,N_5253,N_5316);
nand U5463 (N_5463,N_5218,N_5230);
nor U5464 (N_5464,N_5320,N_5311);
nor U5465 (N_5465,N_5371,N_5208);
nor U5466 (N_5466,N_5333,N_5338);
nor U5467 (N_5467,N_5251,N_5242);
xor U5468 (N_5468,N_5361,N_5326);
nand U5469 (N_5469,N_5277,N_5291);
or U5470 (N_5470,N_5269,N_5314);
or U5471 (N_5471,N_5342,N_5377);
and U5472 (N_5472,N_5380,N_5292);
xor U5473 (N_5473,N_5232,N_5255);
nand U5474 (N_5474,N_5210,N_5249);
and U5475 (N_5475,N_5394,N_5270);
nand U5476 (N_5476,N_5368,N_5370);
xor U5477 (N_5477,N_5355,N_5398);
nor U5478 (N_5478,N_5358,N_5332);
nor U5479 (N_5479,N_5225,N_5273);
or U5480 (N_5480,N_5209,N_5299);
nand U5481 (N_5481,N_5201,N_5369);
nand U5482 (N_5482,N_5289,N_5280);
and U5483 (N_5483,N_5336,N_5243);
and U5484 (N_5484,N_5219,N_5373);
xor U5485 (N_5485,N_5224,N_5300);
xor U5486 (N_5486,N_5294,N_5272);
and U5487 (N_5487,N_5276,N_5212);
nand U5488 (N_5488,N_5200,N_5228);
nand U5489 (N_5489,N_5240,N_5367);
nand U5490 (N_5490,N_5354,N_5310);
or U5491 (N_5491,N_5393,N_5375);
and U5492 (N_5492,N_5214,N_5223);
nor U5493 (N_5493,N_5213,N_5282);
and U5494 (N_5494,N_5386,N_5235);
or U5495 (N_5495,N_5267,N_5220);
xnor U5496 (N_5496,N_5351,N_5248);
or U5497 (N_5497,N_5206,N_5286);
or U5498 (N_5498,N_5384,N_5287);
nor U5499 (N_5499,N_5222,N_5385);
nand U5500 (N_5500,N_5294,N_5227);
nor U5501 (N_5501,N_5320,N_5314);
xnor U5502 (N_5502,N_5201,N_5222);
xnor U5503 (N_5503,N_5205,N_5258);
or U5504 (N_5504,N_5336,N_5235);
nand U5505 (N_5505,N_5265,N_5214);
or U5506 (N_5506,N_5332,N_5253);
nand U5507 (N_5507,N_5230,N_5236);
or U5508 (N_5508,N_5215,N_5201);
and U5509 (N_5509,N_5278,N_5263);
xor U5510 (N_5510,N_5340,N_5207);
xor U5511 (N_5511,N_5334,N_5288);
xnor U5512 (N_5512,N_5251,N_5322);
nor U5513 (N_5513,N_5238,N_5352);
and U5514 (N_5514,N_5216,N_5393);
and U5515 (N_5515,N_5362,N_5294);
nand U5516 (N_5516,N_5397,N_5215);
xor U5517 (N_5517,N_5387,N_5300);
xnor U5518 (N_5518,N_5201,N_5223);
nor U5519 (N_5519,N_5293,N_5229);
or U5520 (N_5520,N_5226,N_5344);
nand U5521 (N_5521,N_5228,N_5361);
or U5522 (N_5522,N_5216,N_5338);
xnor U5523 (N_5523,N_5237,N_5330);
and U5524 (N_5524,N_5278,N_5380);
nand U5525 (N_5525,N_5378,N_5351);
xnor U5526 (N_5526,N_5373,N_5339);
nand U5527 (N_5527,N_5357,N_5214);
nor U5528 (N_5528,N_5274,N_5260);
and U5529 (N_5529,N_5232,N_5324);
nand U5530 (N_5530,N_5336,N_5363);
nor U5531 (N_5531,N_5313,N_5234);
nor U5532 (N_5532,N_5294,N_5298);
xor U5533 (N_5533,N_5326,N_5260);
nor U5534 (N_5534,N_5212,N_5294);
nor U5535 (N_5535,N_5218,N_5277);
and U5536 (N_5536,N_5339,N_5337);
and U5537 (N_5537,N_5337,N_5285);
or U5538 (N_5538,N_5217,N_5397);
or U5539 (N_5539,N_5307,N_5362);
nand U5540 (N_5540,N_5358,N_5290);
and U5541 (N_5541,N_5217,N_5275);
xor U5542 (N_5542,N_5307,N_5354);
or U5543 (N_5543,N_5274,N_5391);
and U5544 (N_5544,N_5313,N_5364);
xor U5545 (N_5545,N_5284,N_5294);
and U5546 (N_5546,N_5396,N_5203);
nand U5547 (N_5547,N_5209,N_5292);
xnor U5548 (N_5548,N_5257,N_5325);
nand U5549 (N_5549,N_5263,N_5311);
or U5550 (N_5550,N_5266,N_5272);
nor U5551 (N_5551,N_5327,N_5264);
xnor U5552 (N_5552,N_5257,N_5357);
or U5553 (N_5553,N_5207,N_5345);
nand U5554 (N_5554,N_5390,N_5254);
nand U5555 (N_5555,N_5385,N_5252);
or U5556 (N_5556,N_5230,N_5387);
xnor U5557 (N_5557,N_5252,N_5383);
and U5558 (N_5558,N_5377,N_5285);
nand U5559 (N_5559,N_5218,N_5346);
and U5560 (N_5560,N_5381,N_5350);
nand U5561 (N_5561,N_5331,N_5213);
and U5562 (N_5562,N_5259,N_5372);
nand U5563 (N_5563,N_5230,N_5293);
xnor U5564 (N_5564,N_5214,N_5337);
nor U5565 (N_5565,N_5270,N_5278);
nand U5566 (N_5566,N_5382,N_5209);
nor U5567 (N_5567,N_5220,N_5384);
nor U5568 (N_5568,N_5302,N_5217);
and U5569 (N_5569,N_5313,N_5254);
nand U5570 (N_5570,N_5203,N_5243);
xor U5571 (N_5571,N_5303,N_5372);
and U5572 (N_5572,N_5317,N_5312);
nor U5573 (N_5573,N_5359,N_5342);
and U5574 (N_5574,N_5301,N_5203);
nand U5575 (N_5575,N_5333,N_5239);
or U5576 (N_5576,N_5367,N_5336);
and U5577 (N_5577,N_5381,N_5344);
and U5578 (N_5578,N_5323,N_5267);
xnor U5579 (N_5579,N_5323,N_5218);
nand U5580 (N_5580,N_5265,N_5374);
nand U5581 (N_5581,N_5248,N_5309);
nor U5582 (N_5582,N_5275,N_5324);
and U5583 (N_5583,N_5243,N_5216);
nor U5584 (N_5584,N_5235,N_5323);
and U5585 (N_5585,N_5253,N_5266);
nor U5586 (N_5586,N_5315,N_5391);
xor U5587 (N_5587,N_5317,N_5354);
xor U5588 (N_5588,N_5227,N_5373);
or U5589 (N_5589,N_5317,N_5212);
nand U5590 (N_5590,N_5223,N_5205);
and U5591 (N_5591,N_5232,N_5238);
nand U5592 (N_5592,N_5396,N_5305);
nor U5593 (N_5593,N_5286,N_5251);
nor U5594 (N_5594,N_5283,N_5389);
nor U5595 (N_5595,N_5399,N_5273);
and U5596 (N_5596,N_5325,N_5276);
or U5597 (N_5597,N_5229,N_5283);
nor U5598 (N_5598,N_5381,N_5288);
and U5599 (N_5599,N_5262,N_5316);
xor U5600 (N_5600,N_5474,N_5462);
nand U5601 (N_5601,N_5453,N_5521);
and U5602 (N_5602,N_5586,N_5419);
or U5603 (N_5603,N_5591,N_5593);
and U5604 (N_5604,N_5501,N_5523);
and U5605 (N_5605,N_5412,N_5438);
or U5606 (N_5606,N_5471,N_5448);
xnor U5607 (N_5607,N_5525,N_5481);
nand U5608 (N_5608,N_5426,N_5569);
nor U5609 (N_5609,N_5415,N_5581);
or U5610 (N_5610,N_5507,N_5416);
or U5611 (N_5611,N_5442,N_5440);
xnor U5612 (N_5612,N_5597,N_5499);
nor U5613 (N_5613,N_5497,N_5503);
nand U5614 (N_5614,N_5460,N_5445);
nor U5615 (N_5615,N_5577,N_5552);
xnor U5616 (N_5616,N_5439,N_5473);
and U5617 (N_5617,N_5541,N_5588);
nor U5618 (N_5618,N_5544,N_5598);
nand U5619 (N_5619,N_5432,N_5546);
and U5620 (N_5620,N_5464,N_5506);
nor U5621 (N_5621,N_5566,N_5530);
xnor U5622 (N_5622,N_5459,N_5553);
nor U5623 (N_5623,N_5492,N_5557);
nand U5624 (N_5624,N_5452,N_5511);
xnor U5625 (N_5625,N_5500,N_5517);
nor U5626 (N_5626,N_5455,N_5450);
xnor U5627 (N_5627,N_5595,N_5568);
nor U5628 (N_5628,N_5449,N_5466);
xnor U5629 (N_5629,N_5509,N_5512);
and U5630 (N_5630,N_5469,N_5428);
and U5631 (N_5631,N_5447,N_5522);
nand U5632 (N_5632,N_5413,N_5534);
and U5633 (N_5633,N_5502,N_5480);
xnor U5634 (N_5634,N_5582,N_5590);
nand U5635 (N_5635,N_5579,N_5527);
xnor U5636 (N_5636,N_5434,N_5536);
nand U5637 (N_5637,N_5491,N_5494);
nor U5638 (N_5638,N_5560,N_5468);
nand U5639 (N_5639,N_5547,N_5531);
and U5640 (N_5640,N_5488,N_5403);
and U5641 (N_5641,N_5524,N_5545);
and U5642 (N_5642,N_5558,N_5587);
or U5643 (N_5643,N_5549,N_5402);
and U5644 (N_5644,N_5574,N_5537);
or U5645 (N_5645,N_5562,N_5479);
or U5646 (N_5646,N_5457,N_5504);
and U5647 (N_5647,N_5478,N_5404);
nor U5648 (N_5648,N_5443,N_5554);
nand U5649 (N_5649,N_5423,N_5528);
xor U5650 (N_5650,N_5436,N_5421);
and U5651 (N_5651,N_5435,N_5508);
or U5652 (N_5652,N_5493,N_5465);
and U5653 (N_5653,N_5490,N_5446);
nor U5654 (N_5654,N_5540,N_5529);
nand U5655 (N_5655,N_5559,N_5429);
or U5656 (N_5656,N_5456,N_5437);
and U5657 (N_5657,N_5430,N_5475);
nand U5658 (N_5658,N_5418,N_5489);
and U5659 (N_5659,N_5519,N_5564);
xor U5660 (N_5660,N_5561,N_5496);
or U5661 (N_5661,N_5410,N_5476);
nor U5662 (N_5662,N_5411,N_5520);
or U5663 (N_5663,N_5461,N_5406);
nand U5664 (N_5664,N_5485,N_5414);
or U5665 (N_5665,N_5425,N_5484);
and U5666 (N_5666,N_5451,N_5583);
nor U5667 (N_5667,N_5589,N_5486);
nor U5668 (N_5668,N_5526,N_5567);
or U5669 (N_5669,N_5407,N_5599);
xor U5670 (N_5670,N_5482,N_5556);
nor U5671 (N_5671,N_5470,N_5515);
and U5672 (N_5672,N_5441,N_5575);
or U5673 (N_5673,N_5565,N_5563);
xor U5674 (N_5674,N_5498,N_5409);
and U5675 (N_5675,N_5467,N_5592);
and U5676 (N_5676,N_5408,N_5400);
nand U5677 (N_5677,N_5533,N_5514);
xor U5678 (N_5678,N_5477,N_5458);
xnor U5679 (N_5679,N_5510,N_5585);
nor U5680 (N_5680,N_5532,N_5516);
or U5681 (N_5681,N_5417,N_5594);
or U5682 (N_5682,N_5444,N_5551);
nor U5683 (N_5683,N_5405,N_5454);
and U5684 (N_5684,N_5570,N_5427);
nor U5685 (N_5685,N_5401,N_5422);
and U5686 (N_5686,N_5572,N_5518);
xnor U5687 (N_5687,N_5576,N_5538);
nand U5688 (N_5688,N_5431,N_5548);
and U5689 (N_5689,N_5584,N_5539);
nand U5690 (N_5690,N_5555,N_5573);
nor U5691 (N_5691,N_5571,N_5472);
and U5692 (N_5692,N_5424,N_5513);
nor U5693 (N_5693,N_5578,N_5550);
xor U5694 (N_5694,N_5483,N_5543);
or U5695 (N_5695,N_5433,N_5535);
nor U5696 (N_5696,N_5596,N_5463);
or U5697 (N_5697,N_5542,N_5580);
and U5698 (N_5698,N_5420,N_5495);
and U5699 (N_5699,N_5487,N_5505);
xor U5700 (N_5700,N_5543,N_5441);
or U5701 (N_5701,N_5420,N_5468);
and U5702 (N_5702,N_5570,N_5554);
or U5703 (N_5703,N_5550,N_5419);
nor U5704 (N_5704,N_5486,N_5406);
xnor U5705 (N_5705,N_5522,N_5437);
or U5706 (N_5706,N_5464,N_5531);
nor U5707 (N_5707,N_5532,N_5418);
or U5708 (N_5708,N_5489,N_5446);
nand U5709 (N_5709,N_5451,N_5461);
nand U5710 (N_5710,N_5445,N_5422);
nor U5711 (N_5711,N_5467,N_5513);
nor U5712 (N_5712,N_5556,N_5502);
nor U5713 (N_5713,N_5430,N_5485);
or U5714 (N_5714,N_5510,N_5548);
and U5715 (N_5715,N_5436,N_5519);
xnor U5716 (N_5716,N_5580,N_5460);
or U5717 (N_5717,N_5542,N_5470);
nand U5718 (N_5718,N_5433,N_5402);
nor U5719 (N_5719,N_5508,N_5473);
nor U5720 (N_5720,N_5527,N_5485);
or U5721 (N_5721,N_5440,N_5540);
or U5722 (N_5722,N_5563,N_5496);
or U5723 (N_5723,N_5490,N_5428);
nor U5724 (N_5724,N_5420,N_5545);
nand U5725 (N_5725,N_5431,N_5526);
nand U5726 (N_5726,N_5416,N_5444);
nand U5727 (N_5727,N_5546,N_5514);
nand U5728 (N_5728,N_5467,N_5459);
or U5729 (N_5729,N_5529,N_5511);
or U5730 (N_5730,N_5574,N_5518);
nor U5731 (N_5731,N_5455,N_5495);
nand U5732 (N_5732,N_5471,N_5571);
and U5733 (N_5733,N_5559,N_5481);
and U5734 (N_5734,N_5597,N_5490);
or U5735 (N_5735,N_5585,N_5500);
nand U5736 (N_5736,N_5497,N_5574);
nor U5737 (N_5737,N_5553,N_5451);
xor U5738 (N_5738,N_5508,N_5451);
and U5739 (N_5739,N_5448,N_5429);
nor U5740 (N_5740,N_5526,N_5460);
xnor U5741 (N_5741,N_5464,N_5530);
or U5742 (N_5742,N_5599,N_5420);
and U5743 (N_5743,N_5458,N_5538);
nor U5744 (N_5744,N_5578,N_5546);
nor U5745 (N_5745,N_5421,N_5534);
nand U5746 (N_5746,N_5530,N_5508);
nand U5747 (N_5747,N_5426,N_5543);
or U5748 (N_5748,N_5505,N_5450);
nor U5749 (N_5749,N_5464,N_5422);
and U5750 (N_5750,N_5589,N_5567);
and U5751 (N_5751,N_5564,N_5493);
xnor U5752 (N_5752,N_5426,N_5500);
nand U5753 (N_5753,N_5559,N_5462);
nor U5754 (N_5754,N_5558,N_5408);
xnor U5755 (N_5755,N_5410,N_5585);
and U5756 (N_5756,N_5550,N_5440);
nand U5757 (N_5757,N_5545,N_5573);
nor U5758 (N_5758,N_5582,N_5407);
xor U5759 (N_5759,N_5409,N_5530);
nand U5760 (N_5760,N_5494,N_5415);
and U5761 (N_5761,N_5576,N_5476);
nand U5762 (N_5762,N_5403,N_5414);
nand U5763 (N_5763,N_5510,N_5438);
nor U5764 (N_5764,N_5530,N_5476);
or U5765 (N_5765,N_5501,N_5560);
nor U5766 (N_5766,N_5525,N_5562);
and U5767 (N_5767,N_5515,N_5509);
and U5768 (N_5768,N_5476,N_5488);
and U5769 (N_5769,N_5506,N_5509);
or U5770 (N_5770,N_5408,N_5404);
and U5771 (N_5771,N_5478,N_5411);
or U5772 (N_5772,N_5483,N_5597);
and U5773 (N_5773,N_5472,N_5581);
nor U5774 (N_5774,N_5585,N_5419);
or U5775 (N_5775,N_5405,N_5450);
or U5776 (N_5776,N_5413,N_5561);
and U5777 (N_5777,N_5516,N_5411);
or U5778 (N_5778,N_5592,N_5500);
and U5779 (N_5779,N_5515,N_5514);
nor U5780 (N_5780,N_5545,N_5503);
nand U5781 (N_5781,N_5527,N_5418);
xnor U5782 (N_5782,N_5479,N_5489);
and U5783 (N_5783,N_5581,N_5453);
or U5784 (N_5784,N_5493,N_5592);
xnor U5785 (N_5785,N_5479,N_5442);
or U5786 (N_5786,N_5580,N_5502);
nor U5787 (N_5787,N_5426,N_5425);
xnor U5788 (N_5788,N_5430,N_5545);
nand U5789 (N_5789,N_5415,N_5501);
or U5790 (N_5790,N_5542,N_5436);
nand U5791 (N_5791,N_5569,N_5471);
nand U5792 (N_5792,N_5460,N_5555);
and U5793 (N_5793,N_5497,N_5516);
or U5794 (N_5794,N_5402,N_5566);
xor U5795 (N_5795,N_5470,N_5461);
nand U5796 (N_5796,N_5563,N_5486);
or U5797 (N_5797,N_5414,N_5506);
and U5798 (N_5798,N_5443,N_5404);
nor U5799 (N_5799,N_5548,N_5504);
xor U5800 (N_5800,N_5629,N_5710);
xnor U5801 (N_5801,N_5610,N_5720);
nand U5802 (N_5802,N_5664,N_5601);
or U5803 (N_5803,N_5766,N_5613);
xor U5804 (N_5804,N_5783,N_5646);
or U5805 (N_5805,N_5699,N_5623);
nand U5806 (N_5806,N_5672,N_5730);
and U5807 (N_5807,N_5787,N_5657);
or U5808 (N_5808,N_5729,N_5695);
nor U5809 (N_5809,N_5763,N_5683);
or U5810 (N_5810,N_5626,N_5640);
nor U5811 (N_5811,N_5693,N_5772);
nor U5812 (N_5812,N_5722,N_5671);
xnor U5813 (N_5813,N_5621,N_5706);
or U5814 (N_5814,N_5639,N_5619);
nand U5815 (N_5815,N_5785,N_5667);
nor U5816 (N_5816,N_5685,N_5603);
nand U5817 (N_5817,N_5617,N_5780);
xor U5818 (N_5818,N_5669,N_5745);
nand U5819 (N_5819,N_5694,N_5615);
and U5820 (N_5820,N_5677,N_5760);
and U5821 (N_5821,N_5734,N_5756);
or U5822 (N_5822,N_5779,N_5755);
and U5823 (N_5823,N_5781,N_5697);
xnor U5824 (N_5824,N_5684,N_5792);
nand U5825 (N_5825,N_5688,N_5707);
xnor U5826 (N_5826,N_5716,N_5743);
nand U5827 (N_5827,N_5658,N_5718);
nand U5828 (N_5828,N_5612,N_5659);
and U5829 (N_5829,N_5673,N_5773);
or U5830 (N_5830,N_5752,N_5618);
and U5831 (N_5831,N_5775,N_5696);
xnor U5832 (N_5832,N_5609,N_5634);
or U5833 (N_5833,N_5660,N_5776);
nand U5834 (N_5834,N_5627,N_5663);
and U5835 (N_5835,N_5633,N_5624);
and U5836 (N_5836,N_5717,N_5638);
and U5837 (N_5837,N_5794,N_5791);
and U5838 (N_5838,N_5749,N_5784);
nand U5839 (N_5839,N_5644,N_5630);
xnor U5840 (N_5840,N_5719,N_5681);
or U5841 (N_5841,N_5777,N_5698);
nand U5842 (N_5842,N_5747,N_5641);
nand U5843 (N_5843,N_5652,N_5762);
and U5844 (N_5844,N_5712,N_5628);
and U5845 (N_5845,N_5742,N_5705);
nand U5846 (N_5846,N_5757,N_5678);
or U5847 (N_5847,N_5625,N_5655);
and U5848 (N_5848,N_5758,N_5721);
or U5849 (N_5849,N_5748,N_5645);
nor U5850 (N_5850,N_5713,N_5797);
xor U5851 (N_5851,N_5774,N_5642);
nor U5852 (N_5852,N_5690,N_5701);
or U5853 (N_5853,N_5731,N_5631);
nand U5854 (N_5854,N_5620,N_5607);
xnor U5855 (N_5855,N_5753,N_5738);
nand U5856 (N_5856,N_5650,N_5796);
and U5857 (N_5857,N_5751,N_5715);
nand U5858 (N_5858,N_5602,N_5676);
or U5859 (N_5859,N_5704,N_5653);
xor U5860 (N_5860,N_5795,N_5793);
or U5861 (N_5861,N_5764,N_5636);
nor U5862 (N_5862,N_5703,N_5727);
nand U5863 (N_5863,N_5604,N_5771);
or U5864 (N_5864,N_5643,N_5674);
nand U5865 (N_5865,N_5782,N_5686);
and U5866 (N_5866,N_5790,N_5725);
nand U5867 (N_5867,N_5714,N_5679);
and U5868 (N_5868,N_5635,N_5737);
or U5869 (N_5869,N_5648,N_5765);
xnor U5870 (N_5870,N_5741,N_5744);
or U5871 (N_5871,N_5789,N_5759);
or U5872 (N_5872,N_5728,N_5735);
or U5873 (N_5873,N_5754,N_5649);
or U5874 (N_5874,N_5665,N_5799);
or U5875 (N_5875,N_5767,N_5739);
nor U5876 (N_5876,N_5798,N_5746);
or U5877 (N_5877,N_5632,N_5788);
and U5878 (N_5878,N_5668,N_5740);
and U5879 (N_5879,N_5723,N_5786);
nor U5880 (N_5880,N_5656,N_5770);
xnor U5881 (N_5881,N_5651,N_5661);
nor U5882 (N_5882,N_5733,N_5611);
and U5883 (N_5883,N_5605,N_5662);
and U5884 (N_5884,N_5666,N_5726);
and U5885 (N_5885,N_5675,N_5616);
nor U5886 (N_5886,N_5687,N_5608);
or U5887 (N_5887,N_5680,N_5700);
and U5888 (N_5888,N_5637,N_5606);
nor U5889 (N_5889,N_5670,N_5761);
nor U5890 (N_5890,N_5732,N_5708);
and U5891 (N_5891,N_5750,N_5600);
xnor U5892 (N_5892,N_5689,N_5702);
nand U5893 (N_5893,N_5614,N_5711);
nor U5894 (N_5894,N_5768,N_5736);
nand U5895 (N_5895,N_5778,N_5647);
and U5896 (N_5896,N_5769,N_5709);
or U5897 (N_5897,N_5692,N_5724);
or U5898 (N_5898,N_5654,N_5622);
nor U5899 (N_5899,N_5682,N_5691);
or U5900 (N_5900,N_5789,N_5755);
nand U5901 (N_5901,N_5724,N_5690);
xor U5902 (N_5902,N_5794,N_5714);
and U5903 (N_5903,N_5737,N_5604);
or U5904 (N_5904,N_5769,N_5786);
nand U5905 (N_5905,N_5697,N_5707);
xor U5906 (N_5906,N_5767,N_5727);
nand U5907 (N_5907,N_5719,N_5733);
or U5908 (N_5908,N_5771,N_5777);
nor U5909 (N_5909,N_5607,N_5788);
nor U5910 (N_5910,N_5710,N_5690);
and U5911 (N_5911,N_5707,N_5665);
xnor U5912 (N_5912,N_5700,N_5710);
xnor U5913 (N_5913,N_5749,N_5728);
xnor U5914 (N_5914,N_5602,N_5604);
or U5915 (N_5915,N_5725,N_5648);
xor U5916 (N_5916,N_5632,N_5693);
nor U5917 (N_5917,N_5678,N_5717);
or U5918 (N_5918,N_5691,N_5699);
nor U5919 (N_5919,N_5667,N_5660);
or U5920 (N_5920,N_5793,N_5605);
xor U5921 (N_5921,N_5734,N_5754);
xnor U5922 (N_5922,N_5704,N_5659);
and U5923 (N_5923,N_5756,N_5649);
nor U5924 (N_5924,N_5775,N_5677);
or U5925 (N_5925,N_5729,N_5720);
nand U5926 (N_5926,N_5638,N_5705);
nor U5927 (N_5927,N_5711,N_5766);
xor U5928 (N_5928,N_5780,N_5636);
xnor U5929 (N_5929,N_5606,N_5601);
nand U5930 (N_5930,N_5635,N_5763);
or U5931 (N_5931,N_5639,N_5601);
xor U5932 (N_5932,N_5704,N_5731);
nor U5933 (N_5933,N_5631,N_5646);
or U5934 (N_5934,N_5641,N_5742);
nor U5935 (N_5935,N_5757,N_5688);
nand U5936 (N_5936,N_5687,N_5626);
or U5937 (N_5937,N_5632,N_5620);
nor U5938 (N_5938,N_5705,N_5686);
and U5939 (N_5939,N_5769,N_5771);
nand U5940 (N_5940,N_5642,N_5779);
nand U5941 (N_5941,N_5687,N_5630);
nor U5942 (N_5942,N_5795,N_5760);
xnor U5943 (N_5943,N_5749,N_5611);
nor U5944 (N_5944,N_5711,N_5605);
nor U5945 (N_5945,N_5658,N_5791);
nand U5946 (N_5946,N_5751,N_5740);
nor U5947 (N_5947,N_5729,N_5734);
and U5948 (N_5948,N_5765,N_5695);
nand U5949 (N_5949,N_5673,N_5611);
xnor U5950 (N_5950,N_5606,N_5645);
xor U5951 (N_5951,N_5758,N_5625);
nand U5952 (N_5952,N_5615,N_5718);
xor U5953 (N_5953,N_5735,N_5747);
and U5954 (N_5954,N_5614,N_5603);
nand U5955 (N_5955,N_5682,N_5797);
nor U5956 (N_5956,N_5722,N_5600);
and U5957 (N_5957,N_5690,N_5647);
or U5958 (N_5958,N_5767,N_5694);
or U5959 (N_5959,N_5656,N_5615);
nand U5960 (N_5960,N_5675,N_5659);
nor U5961 (N_5961,N_5652,N_5682);
xnor U5962 (N_5962,N_5693,N_5760);
xnor U5963 (N_5963,N_5719,N_5716);
nor U5964 (N_5964,N_5672,N_5680);
nor U5965 (N_5965,N_5766,N_5656);
and U5966 (N_5966,N_5623,N_5745);
nor U5967 (N_5967,N_5658,N_5657);
xnor U5968 (N_5968,N_5694,N_5763);
and U5969 (N_5969,N_5677,N_5765);
and U5970 (N_5970,N_5646,N_5637);
xor U5971 (N_5971,N_5740,N_5783);
or U5972 (N_5972,N_5697,N_5746);
xor U5973 (N_5973,N_5742,N_5684);
xnor U5974 (N_5974,N_5603,N_5781);
and U5975 (N_5975,N_5740,N_5734);
nand U5976 (N_5976,N_5676,N_5641);
nand U5977 (N_5977,N_5788,N_5669);
nand U5978 (N_5978,N_5644,N_5791);
and U5979 (N_5979,N_5784,N_5739);
or U5980 (N_5980,N_5703,N_5794);
or U5981 (N_5981,N_5609,N_5786);
and U5982 (N_5982,N_5722,N_5646);
or U5983 (N_5983,N_5777,N_5657);
and U5984 (N_5984,N_5616,N_5722);
nor U5985 (N_5985,N_5692,N_5719);
nor U5986 (N_5986,N_5725,N_5645);
nand U5987 (N_5987,N_5629,N_5619);
and U5988 (N_5988,N_5643,N_5682);
nor U5989 (N_5989,N_5748,N_5731);
and U5990 (N_5990,N_5797,N_5703);
nand U5991 (N_5991,N_5605,N_5730);
and U5992 (N_5992,N_5715,N_5706);
or U5993 (N_5993,N_5639,N_5649);
xnor U5994 (N_5994,N_5602,N_5706);
and U5995 (N_5995,N_5790,N_5744);
xnor U5996 (N_5996,N_5783,N_5794);
nor U5997 (N_5997,N_5724,N_5624);
xnor U5998 (N_5998,N_5780,N_5753);
nand U5999 (N_5999,N_5704,N_5628);
xnor U6000 (N_6000,N_5925,N_5916);
nand U6001 (N_6001,N_5918,N_5803);
nor U6002 (N_6002,N_5818,N_5842);
nor U6003 (N_6003,N_5880,N_5962);
nand U6004 (N_6004,N_5977,N_5991);
nor U6005 (N_6005,N_5859,N_5834);
or U6006 (N_6006,N_5826,N_5914);
or U6007 (N_6007,N_5960,N_5922);
and U6008 (N_6008,N_5975,N_5974);
or U6009 (N_6009,N_5901,N_5985);
and U6010 (N_6010,N_5907,N_5822);
nand U6011 (N_6011,N_5838,N_5817);
and U6012 (N_6012,N_5820,N_5967);
nor U6013 (N_6013,N_5872,N_5980);
xor U6014 (N_6014,N_5845,N_5966);
xor U6015 (N_6015,N_5802,N_5807);
nand U6016 (N_6016,N_5969,N_5923);
and U6017 (N_6017,N_5879,N_5851);
nor U6018 (N_6018,N_5891,N_5868);
nor U6019 (N_6019,N_5979,N_5869);
and U6020 (N_6020,N_5849,N_5998);
xor U6021 (N_6021,N_5898,N_5941);
xnor U6022 (N_6022,N_5959,N_5877);
xnor U6023 (N_6023,N_5878,N_5992);
xor U6024 (N_6024,N_5801,N_5949);
nor U6025 (N_6025,N_5978,N_5847);
xnor U6026 (N_6026,N_5811,N_5899);
or U6027 (N_6027,N_5853,N_5964);
and U6028 (N_6028,N_5835,N_5823);
and U6029 (N_6029,N_5912,N_5804);
nor U6030 (N_6030,N_5881,N_5840);
xor U6031 (N_6031,N_5994,N_5893);
nor U6032 (N_6032,N_5933,N_5874);
and U6033 (N_6033,N_5816,N_5846);
nor U6034 (N_6034,N_5965,N_5837);
nand U6035 (N_6035,N_5865,N_5830);
xor U6036 (N_6036,N_5928,N_5982);
xnor U6037 (N_6037,N_5906,N_5932);
or U6038 (N_6038,N_5968,N_5937);
and U6039 (N_6039,N_5815,N_5809);
nand U6040 (N_6040,N_5839,N_5850);
and U6041 (N_6041,N_5813,N_5946);
and U6042 (N_6042,N_5973,N_5800);
and U6043 (N_6043,N_5950,N_5938);
or U6044 (N_6044,N_5940,N_5956);
nor U6045 (N_6045,N_5905,N_5911);
or U6046 (N_6046,N_5997,N_5870);
or U6047 (N_6047,N_5887,N_5805);
and U6048 (N_6048,N_5812,N_5951);
nor U6049 (N_6049,N_5958,N_5806);
xnor U6050 (N_6050,N_5934,N_5915);
and U6051 (N_6051,N_5957,N_5952);
nor U6052 (N_6052,N_5995,N_5990);
nand U6053 (N_6053,N_5873,N_5930);
or U6054 (N_6054,N_5882,N_5855);
xnor U6055 (N_6055,N_5909,N_5836);
and U6056 (N_6056,N_5866,N_5814);
nor U6057 (N_6057,N_5856,N_5854);
xnor U6058 (N_6058,N_5929,N_5983);
nor U6059 (N_6059,N_5919,N_5903);
and U6060 (N_6060,N_5875,N_5936);
or U6061 (N_6061,N_5889,N_5876);
and U6062 (N_6062,N_5970,N_5945);
and U6063 (N_6063,N_5961,N_5924);
nand U6064 (N_6064,N_5896,N_5831);
xor U6065 (N_6065,N_5939,N_5910);
nor U6066 (N_6066,N_5908,N_5848);
nor U6067 (N_6067,N_5864,N_5943);
and U6068 (N_6068,N_5935,N_5944);
xor U6069 (N_6069,N_5954,N_5871);
or U6070 (N_6070,N_5825,N_5858);
xor U6071 (N_6071,N_5986,N_5888);
or U6072 (N_6072,N_5884,N_5867);
xnor U6073 (N_6073,N_5988,N_5963);
and U6074 (N_6074,N_5843,N_5900);
and U6075 (N_6075,N_5942,N_5810);
or U6076 (N_6076,N_5993,N_5955);
and U6077 (N_6077,N_5987,N_5913);
xor U6078 (N_6078,N_5989,N_5844);
xnor U6079 (N_6079,N_5821,N_5833);
nand U6080 (N_6080,N_5921,N_5917);
xnor U6081 (N_6081,N_5852,N_5860);
and U6082 (N_6082,N_5948,N_5861);
xor U6083 (N_6083,N_5819,N_5895);
xor U6084 (N_6084,N_5824,N_5996);
or U6085 (N_6085,N_5894,N_5984);
and U6086 (N_6086,N_5890,N_5808);
or U6087 (N_6087,N_5862,N_5857);
and U6088 (N_6088,N_5972,N_5827);
nand U6089 (N_6089,N_5828,N_5902);
or U6090 (N_6090,N_5897,N_5886);
xnor U6091 (N_6091,N_5883,N_5981);
and U6092 (N_6092,N_5976,N_5904);
nor U6093 (N_6093,N_5926,N_5927);
xor U6094 (N_6094,N_5885,N_5832);
or U6095 (N_6095,N_5971,N_5931);
nand U6096 (N_6096,N_5829,N_5920);
nand U6097 (N_6097,N_5999,N_5892);
xor U6098 (N_6098,N_5841,N_5863);
xor U6099 (N_6099,N_5953,N_5947);
xor U6100 (N_6100,N_5983,N_5886);
xor U6101 (N_6101,N_5845,N_5836);
nand U6102 (N_6102,N_5915,N_5812);
or U6103 (N_6103,N_5808,N_5965);
and U6104 (N_6104,N_5895,N_5811);
nor U6105 (N_6105,N_5889,N_5853);
and U6106 (N_6106,N_5816,N_5924);
or U6107 (N_6107,N_5922,N_5877);
or U6108 (N_6108,N_5881,N_5937);
nor U6109 (N_6109,N_5842,N_5984);
or U6110 (N_6110,N_5902,N_5819);
or U6111 (N_6111,N_5927,N_5837);
and U6112 (N_6112,N_5975,N_5871);
or U6113 (N_6113,N_5909,N_5939);
nor U6114 (N_6114,N_5941,N_5890);
nor U6115 (N_6115,N_5915,N_5908);
or U6116 (N_6116,N_5889,N_5816);
nand U6117 (N_6117,N_5912,N_5879);
xor U6118 (N_6118,N_5817,N_5849);
or U6119 (N_6119,N_5912,N_5847);
or U6120 (N_6120,N_5965,N_5825);
nand U6121 (N_6121,N_5934,N_5902);
nand U6122 (N_6122,N_5971,N_5916);
nor U6123 (N_6123,N_5912,N_5837);
xor U6124 (N_6124,N_5969,N_5920);
and U6125 (N_6125,N_5804,N_5893);
nand U6126 (N_6126,N_5934,N_5920);
or U6127 (N_6127,N_5964,N_5925);
nand U6128 (N_6128,N_5829,N_5802);
nor U6129 (N_6129,N_5968,N_5931);
nor U6130 (N_6130,N_5832,N_5807);
or U6131 (N_6131,N_5829,N_5956);
and U6132 (N_6132,N_5907,N_5811);
and U6133 (N_6133,N_5970,N_5997);
nor U6134 (N_6134,N_5929,N_5885);
nand U6135 (N_6135,N_5939,N_5920);
xnor U6136 (N_6136,N_5921,N_5980);
nand U6137 (N_6137,N_5868,N_5864);
nor U6138 (N_6138,N_5820,N_5905);
nand U6139 (N_6139,N_5975,N_5810);
or U6140 (N_6140,N_5920,N_5925);
nor U6141 (N_6141,N_5858,N_5812);
nor U6142 (N_6142,N_5959,N_5888);
and U6143 (N_6143,N_5923,N_5825);
nand U6144 (N_6144,N_5862,N_5879);
nand U6145 (N_6145,N_5845,N_5832);
or U6146 (N_6146,N_5874,N_5828);
nand U6147 (N_6147,N_5916,N_5993);
or U6148 (N_6148,N_5816,N_5965);
and U6149 (N_6149,N_5927,N_5814);
nor U6150 (N_6150,N_5817,N_5860);
nand U6151 (N_6151,N_5878,N_5942);
or U6152 (N_6152,N_5988,N_5891);
nor U6153 (N_6153,N_5916,N_5951);
xnor U6154 (N_6154,N_5885,N_5870);
or U6155 (N_6155,N_5856,N_5853);
and U6156 (N_6156,N_5953,N_5968);
nor U6157 (N_6157,N_5884,N_5889);
nor U6158 (N_6158,N_5821,N_5968);
nor U6159 (N_6159,N_5956,N_5889);
xnor U6160 (N_6160,N_5920,N_5885);
and U6161 (N_6161,N_5975,N_5806);
and U6162 (N_6162,N_5959,N_5853);
or U6163 (N_6163,N_5831,N_5843);
nand U6164 (N_6164,N_5934,N_5879);
nand U6165 (N_6165,N_5838,N_5897);
nand U6166 (N_6166,N_5800,N_5890);
or U6167 (N_6167,N_5814,N_5947);
nor U6168 (N_6168,N_5845,N_5864);
and U6169 (N_6169,N_5848,N_5934);
nand U6170 (N_6170,N_5936,N_5980);
xor U6171 (N_6171,N_5905,N_5803);
nor U6172 (N_6172,N_5911,N_5970);
or U6173 (N_6173,N_5976,N_5986);
and U6174 (N_6174,N_5845,N_5894);
and U6175 (N_6175,N_5831,N_5878);
and U6176 (N_6176,N_5993,N_5964);
or U6177 (N_6177,N_5935,N_5987);
nor U6178 (N_6178,N_5966,N_5807);
or U6179 (N_6179,N_5887,N_5802);
and U6180 (N_6180,N_5855,N_5993);
nor U6181 (N_6181,N_5913,N_5945);
nand U6182 (N_6182,N_5861,N_5947);
or U6183 (N_6183,N_5988,N_5928);
nand U6184 (N_6184,N_5972,N_5804);
nor U6185 (N_6185,N_5862,N_5821);
xnor U6186 (N_6186,N_5921,N_5994);
and U6187 (N_6187,N_5922,N_5886);
nand U6188 (N_6188,N_5950,N_5987);
nand U6189 (N_6189,N_5889,N_5999);
or U6190 (N_6190,N_5899,N_5895);
nand U6191 (N_6191,N_5964,N_5937);
or U6192 (N_6192,N_5894,N_5919);
and U6193 (N_6193,N_5880,N_5915);
nand U6194 (N_6194,N_5802,N_5962);
and U6195 (N_6195,N_5977,N_5956);
and U6196 (N_6196,N_5932,N_5942);
and U6197 (N_6197,N_5931,N_5847);
nand U6198 (N_6198,N_5970,N_5963);
nor U6199 (N_6199,N_5982,N_5918);
and U6200 (N_6200,N_6015,N_6122);
nand U6201 (N_6201,N_6101,N_6126);
and U6202 (N_6202,N_6006,N_6099);
nand U6203 (N_6203,N_6117,N_6178);
nand U6204 (N_6204,N_6127,N_6153);
xor U6205 (N_6205,N_6156,N_6194);
xnor U6206 (N_6206,N_6092,N_6182);
and U6207 (N_6207,N_6150,N_6079);
xnor U6208 (N_6208,N_6164,N_6063);
xnor U6209 (N_6209,N_6142,N_6134);
nand U6210 (N_6210,N_6185,N_6031);
nor U6211 (N_6211,N_6149,N_6087);
nor U6212 (N_6212,N_6175,N_6109);
nor U6213 (N_6213,N_6165,N_6121);
nand U6214 (N_6214,N_6093,N_6035);
or U6215 (N_6215,N_6073,N_6118);
xor U6216 (N_6216,N_6089,N_6050);
nor U6217 (N_6217,N_6160,N_6029);
or U6218 (N_6218,N_6002,N_6147);
nand U6219 (N_6219,N_6046,N_6137);
or U6220 (N_6220,N_6159,N_6022);
nand U6221 (N_6221,N_6098,N_6025);
or U6222 (N_6222,N_6011,N_6168);
xnor U6223 (N_6223,N_6049,N_6053);
or U6224 (N_6224,N_6041,N_6067);
and U6225 (N_6225,N_6013,N_6197);
xor U6226 (N_6226,N_6177,N_6061);
nor U6227 (N_6227,N_6174,N_6019);
nor U6228 (N_6228,N_6032,N_6083);
nor U6229 (N_6229,N_6074,N_6173);
and U6230 (N_6230,N_6066,N_6044);
or U6231 (N_6231,N_6000,N_6082);
nor U6232 (N_6232,N_6119,N_6054);
nor U6233 (N_6233,N_6110,N_6155);
or U6234 (N_6234,N_6062,N_6162);
nor U6235 (N_6235,N_6161,N_6130);
nand U6236 (N_6236,N_6020,N_6014);
nand U6237 (N_6237,N_6116,N_6078);
or U6238 (N_6238,N_6143,N_6158);
nor U6239 (N_6239,N_6183,N_6199);
and U6240 (N_6240,N_6136,N_6179);
and U6241 (N_6241,N_6068,N_6094);
and U6242 (N_6242,N_6001,N_6154);
xnor U6243 (N_6243,N_6129,N_6166);
nand U6244 (N_6244,N_6071,N_6120);
nand U6245 (N_6245,N_6108,N_6133);
nand U6246 (N_6246,N_6193,N_6139);
xor U6247 (N_6247,N_6080,N_6023);
and U6248 (N_6248,N_6051,N_6091);
xor U6249 (N_6249,N_6111,N_6105);
and U6250 (N_6250,N_6005,N_6055);
nor U6251 (N_6251,N_6191,N_6172);
nand U6252 (N_6252,N_6010,N_6132);
or U6253 (N_6253,N_6180,N_6043);
nand U6254 (N_6254,N_6075,N_6057);
nor U6255 (N_6255,N_6077,N_6021);
and U6256 (N_6256,N_6038,N_6085);
nor U6257 (N_6257,N_6052,N_6123);
xor U6258 (N_6258,N_6072,N_6148);
or U6259 (N_6259,N_6036,N_6027);
or U6260 (N_6260,N_6151,N_6107);
nor U6261 (N_6261,N_6124,N_6115);
and U6262 (N_6262,N_6196,N_6138);
xnor U6263 (N_6263,N_6003,N_6028);
nor U6264 (N_6264,N_6114,N_6131);
xor U6265 (N_6265,N_6090,N_6039);
xnor U6266 (N_6266,N_6157,N_6084);
nand U6267 (N_6267,N_6152,N_6064);
nor U6268 (N_6268,N_6040,N_6033);
or U6269 (N_6269,N_6065,N_6135);
or U6270 (N_6270,N_6045,N_6144);
or U6271 (N_6271,N_6141,N_6018);
xnor U6272 (N_6272,N_6198,N_6070);
and U6273 (N_6273,N_6195,N_6181);
xnor U6274 (N_6274,N_6095,N_6081);
xnor U6275 (N_6275,N_6017,N_6034);
or U6276 (N_6276,N_6184,N_6190);
nand U6277 (N_6277,N_6112,N_6016);
or U6278 (N_6278,N_6103,N_6037);
and U6279 (N_6279,N_6096,N_6113);
or U6280 (N_6280,N_6146,N_6106);
and U6281 (N_6281,N_6102,N_6024);
xor U6282 (N_6282,N_6004,N_6088);
and U6283 (N_6283,N_6058,N_6030);
nand U6284 (N_6284,N_6128,N_6100);
nand U6285 (N_6285,N_6104,N_6176);
xor U6286 (N_6286,N_6076,N_6125);
and U6287 (N_6287,N_6012,N_6145);
xor U6288 (N_6288,N_6048,N_6026);
or U6289 (N_6289,N_6059,N_6167);
nand U6290 (N_6290,N_6086,N_6009);
nor U6291 (N_6291,N_6060,N_6140);
and U6292 (N_6292,N_6007,N_6047);
or U6293 (N_6293,N_6163,N_6187);
xor U6294 (N_6294,N_6069,N_6008);
nor U6295 (N_6295,N_6186,N_6189);
nand U6296 (N_6296,N_6097,N_6192);
xnor U6297 (N_6297,N_6188,N_6056);
xor U6298 (N_6298,N_6170,N_6042);
or U6299 (N_6299,N_6171,N_6169);
or U6300 (N_6300,N_6152,N_6021);
nor U6301 (N_6301,N_6107,N_6028);
and U6302 (N_6302,N_6137,N_6134);
or U6303 (N_6303,N_6100,N_6008);
and U6304 (N_6304,N_6074,N_6058);
xnor U6305 (N_6305,N_6165,N_6191);
nand U6306 (N_6306,N_6167,N_6182);
and U6307 (N_6307,N_6026,N_6001);
or U6308 (N_6308,N_6078,N_6119);
and U6309 (N_6309,N_6134,N_6185);
xnor U6310 (N_6310,N_6127,N_6050);
nand U6311 (N_6311,N_6197,N_6131);
nand U6312 (N_6312,N_6100,N_6007);
nand U6313 (N_6313,N_6004,N_6129);
nand U6314 (N_6314,N_6110,N_6166);
nor U6315 (N_6315,N_6118,N_6101);
xor U6316 (N_6316,N_6179,N_6008);
nand U6317 (N_6317,N_6134,N_6091);
nor U6318 (N_6318,N_6052,N_6165);
nand U6319 (N_6319,N_6074,N_6158);
nor U6320 (N_6320,N_6065,N_6120);
xnor U6321 (N_6321,N_6191,N_6041);
nand U6322 (N_6322,N_6075,N_6038);
xnor U6323 (N_6323,N_6007,N_6048);
nand U6324 (N_6324,N_6192,N_6183);
nor U6325 (N_6325,N_6113,N_6093);
and U6326 (N_6326,N_6146,N_6076);
or U6327 (N_6327,N_6114,N_6080);
nand U6328 (N_6328,N_6120,N_6031);
and U6329 (N_6329,N_6110,N_6124);
nand U6330 (N_6330,N_6168,N_6014);
xnor U6331 (N_6331,N_6141,N_6088);
xor U6332 (N_6332,N_6139,N_6000);
or U6333 (N_6333,N_6080,N_6186);
nand U6334 (N_6334,N_6062,N_6072);
nand U6335 (N_6335,N_6164,N_6047);
xor U6336 (N_6336,N_6004,N_6109);
and U6337 (N_6337,N_6151,N_6178);
or U6338 (N_6338,N_6051,N_6014);
xnor U6339 (N_6339,N_6126,N_6002);
nand U6340 (N_6340,N_6131,N_6122);
and U6341 (N_6341,N_6124,N_6044);
nand U6342 (N_6342,N_6124,N_6030);
xor U6343 (N_6343,N_6097,N_6193);
xor U6344 (N_6344,N_6130,N_6016);
or U6345 (N_6345,N_6084,N_6158);
and U6346 (N_6346,N_6063,N_6175);
nand U6347 (N_6347,N_6111,N_6187);
and U6348 (N_6348,N_6101,N_6141);
or U6349 (N_6349,N_6066,N_6072);
nand U6350 (N_6350,N_6086,N_6026);
nand U6351 (N_6351,N_6146,N_6050);
xnor U6352 (N_6352,N_6105,N_6070);
nand U6353 (N_6353,N_6178,N_6047);
or U6354 (N_6354,N_6111,N_6086);
nand U6355 (N_6355,N_6147,N_6178);
and U6356 (N_6356,N_6041,N_6159);
xnor U6357 (N_6357,N_6086,N_6143);
xnor U6358 (N_6358,N_6034,N_6114);
nor U6359 (N_6359,N_6107,N_6037);
and U6360 (N_6360,N_6109,N_6180);
nor U6361 (N_6361,N_6104,N_6007);
xor U6362 (N_6362,N_6082,N_6172);
or U6363 (N_6363,N_6154,N_6018);
and U6364 (N_6364,N_6110,N_6070);
nor U6365 (N_6365,N_6122,N_6085);
nor U6366 (N_6366,N_6032,N_6055);
nand U6367 (N_6367,N_6144,N_6163);
nor U6368 (N_6368,N_6194,N_6164);
or U6369 (N_6369,N_6188,N_6064);
nand U6370 (N_6370,N_6130,N_6047);
nand U6371 (N_6371,N_6022,N_6192);
or U6372 (N_6372,N_6189,N_6075);
nor U6373 (N_6373,N_6037,N_6013);
nor U6374 (N_6374,N_6020,N_6125);
and U6375 (N_6375,N_6069,N_6006);
and U6376 (N_6376,N_6011,N_6081);
xor U6377 (N_6377,N_6030,N_6028);
and U6378 (N_6378,N_6060,N_6188);
xnor U6379 (N_6379,N_6006,N_6147);
and U6380 (N_6380,N_6059,N_6080);
or U6381 (N_6381,N_6149,N_6031);
xnor U6382 (N_6382,N_6116,N_6085);
or U6383 (N_6383,N_6044,N_6091);
nand U6384 (N_6384,N_6037,N_6050);
nor U6385 (N_6385,N_6146,N_6126);
nand U6386 (N_6386,N_6042,N_6059);
and U6387 (N_6387,N_6119,N_6088);
or U6388 (N_6388,N_6086,N_6133);
or U6389 (N_6389,N_6176,N_6180);
xor U6390 (N_6390,N_6027,N_6037);
nand U6391 (N_6391,N_6153,N_6039);
nor U6392 (N_6392,N_6048,N_6190);
and U6393 (N_6393,N_6011,N_6023);
nand U6394 (N_6394,N_6112,N_6170);
xnor U6395 (N_6395,N_6064,N_6175);
or U6396 (N_6396,N_6139,N_6121);
or U6397 (N_6397,N_6064,N_6030);
xnor U6398 (N_6398,N_6197,N_6103);
nor U6399 (N_6399,N_6097,N_6146);
nor U6400 (N_6400,N_6287,N_6204);
xor U6401 (N_6401,N_6322,N_6267);
nand U6402 (N_6402,N_6378,N_6276);
and U6403 (N_6403,N_6302,N_6338);
and U6404 (N_6404,N_6230,N_6234);
nor U6405 (N_6405,N_6358,N_6272);
or U6406 (N_6406,N_6203,N_6206);
xnor U6407 (N_6407,N_6240,N_6334);
xor U6408 (N_6408,N_6355,N_6333);
nor U6409 (N_6409,N_6266,N_6235);
xor U6410 (N_6410,N_6379,N_6216);
and U6411 (N_6411,N_6306,N_6229);
nor U6412 (N_6412,N_6252,N_6382);
nor U6413 (N_6413,N_6324,N_6363);
or U6414 (N_6414,N_6353,N_6274);
nand U6415 (N_6415,N_6284,N_6359);
nor U6416 (N_6416,N_6291,N_6241);
nor U6417 (N_6417,N_6329,N_6370);
nor U6418 (N_6418,N_6288,N_6354);
nand U6419 (N_6419,N_6347,N_6351);
xor U6420 (N_6420,N_6392,N_6251);
nand U6421 (N_6421,N_6246,N_6280);
nor U6422 (N_6422,N_6228,N_6383);
nor U6423 (N_6423,N_6292,N_6256);
nor U6424 (N_6424,N_6231,N_6397);
or U6425 (N_6425,N_6242,N_6250);
nor U6426 (N_6426,N_6210,N_6224);
nor U6427 (N_6427,N_6296,N_6244);
xnor U6428 (N_6428,N_6258,N_6356);
and U6429 (N_6429,N_6261,N_6282);
and U6430 (N_6430,N_6336,N_6386);
nand U6431 (N_6431,N_6262,N_6344);
xnor U6432 (N_6432,N_6236,N_6398);
nor U6433 (N_6433,N_6289,N_6248);
xor U6434 (N_6434,N_6352,N_6384);
and U6435 (N_6435,N_6237,N_6254);
and U6436 (N_6436,N_6277,N_6215);
and U6437 (N_6437,N_6357,N_6260);
nor U6438 (N_6438,N_6326,N_6259);
and U6439 (N_6439,N_6270,N_6295);
or U6440 (N_6440,N_6394,N_6360);
nand U6441 (N_6441,N_6283,N_6209);
or U6442 (N_6442,N_6311,N_6279);
nor U6443 (N_6443,N_6389,N_6310);
and U6444 (N_6444,N_6393,N_6388);
nor U6445 (N_6445,N_6332,N_6369);
xnor U6446 (N_6446,N_6315,N_6249);
and U6447 (N_6447,N_6217,N_6211);
xor U6448 (N_6448,N_6313,N_6218);
nor U6449 (N_6449,N_6381,N_6387);
nand U6450 (N_6450,N_6297,N_6342);
and U6451 (N_6451,N_6376,N_6257);
or U6452 (N_6452,N_6390,N_6330);
and U6453 (N_6453,N_6349,N_6308);
or U6454 (N_6454,N_6346,N_6227);
nor U6455 (N_6455,N_6232,N_6331);
or U6456 (N_6456,N_6345,N_6214);
nor U6457 (N_6457,N_6278,N_6341);
xnor U6458 (N_6458,N_6255,N_6238);
nand U6459 (N_6459,N_6309,N_6264);
and U6460 (N_6460,N_6364,N_6371);
nand U6461 (N_6461,N_6375,N_6368);
or U6462 (N_6462,N_6233,N_6320);
or U6463 (N_6463,N_6286,N_6221);
nand U6464 (N_6464,N_6294,N_6367);
or U6465 (N_6465,N_6223,N_6208);
or U6466 (N_6466,N_6362,N_6391);
xnor U6467 (N_6467,N_6321,N_6380);
and U6468 (N_6468,N_6281,N_6339);
nor U6469 (N_6469,N_6207,N_6325);
nor U6470 (N_6470,N_6335,N_6318);
xnor U6471 (N_6471,N_6319,N_6374);
nor U6472 (N_6472,N_6300,N_6226);
nand U6473 (N_6473,N_6366,N_6202);
and U6474 (N_6474,N_6263,N_6213);
or U6475 (N_6475,N_6350,N_6312);
nand U6476 (N_6476,N_6299,N_6269);
xnor U6477 (N_6477,N_6201,N_6340);
and U6478 (N_6478,N_6307,N_6314);
xnor U6479 (N_6479,N_6385,N_6265);
xor U6480 (N_6480,N_6285,N_6301);
xnor U6481 (N_6481,N_6222,N_6220);
nor U6482 (N_6482,N_6348,N_6399);
nand U6483 (N_6483,N_6337,N_6243);
xnor U6484 (N_6484,N_6304,N_6273);
nand U6485 (N_6485,N_6247,N_6343);
or U6486 (N_6486,N_6239,N_6212);
or U6487 (N_6487,N_6268,N_6305);
or U6488 (N_6488,N_6219,N_6317);
xor U6489 (N_6489,N_6271,N_6365);
or U6490 (N_6490,N_6328,N_6245);
nand U6491 (N_6491,N_6395,N_6298);
and U6492 (N_6492,N_6377,N_6396);
and U6493 (N_6493,N_6293,N_6372);
and U6494 (N_6494,N_6373,N_6200);
xor U6495 (N_6495,N_6275,N_6290);
or U6496 (N_6496,N_6303,N_6361);
and U6497 (N_6497,N_6253,N_6323);
nand U6498 (N_6498,N_6205,N_6316);
and U6499 (N_6499,N_6327,N_6225);
xnor U6500 (N_6500,N_6214,N_6301);
or U6501 (N_6501,N_6390,N_6367);
nor U6502 (N_6502,N_6309,N_6370);
nor U6503 (N_6503,N_6277,N_6331);
xnor U6504 (N_6504,N_6237,N_6286);
xnor U6505 (N_6505,N_6259,N_6374);
or U6506 (N_6506,N_6339,N_6376);
xnor U6507 (N_6507,N_6398,N_6267);
nand U6508 (N_6508,N_6290,N_6292);
or U6509 (N_6509,N_6299,N_6233);
nand U6510 (N_6510,N_6349,N_6251);
nand U6511 (N_6511,N_6349,N_6219);
or U6512 (N_6512,N_6284,N_6247);
and U6513 (N_6513,N_6249,N_6259);
xor U6514 (N_6514,N_6345,N_6218);
xor U6515 (N_6515,N_6212,N_6206);
nor U6516 (N_6516,N_6220,N_6294);
xnor U6517 (N_6517,N_6217,N_6345);
xnor U6518 (N_6518,N_6379,N_6346);
or U6519 (N_6519,N_6361,N_6339);
or U6520 (N_6520,N_6383,N_6270);
and U6521 (N_6521,N_6223,N_6228);
xnor U6522 (N_6522,N_6274,N_6275);
and U6523 (N_6523,N_6301,N_6391);
xor U6524 (N_6524,N_6280,N_6316);
nor U6525 (N_6525,N_6386,N_6252);
xnor U6526 (N_6526,N_6314,N_6303);
or U6527 (N_6527,N_6383,N_6230);
xnor U6528 (N_6528,N_6370,N_6236);
and U6529 (N_6529,N_6210,N_6355);
xor U6530 (N_6530,N_6398,N_6294);
nor U6531 (N_6531,N_6256,N_6350);
xor U6532 (N_6532,N_6341,N_6202);
nand U6533 (N_6533,N_6304,N_6326);
xnor U6534 (N_6534,N_6379,N_6371);
xor U6535 (N_6535,N_6385,N_6326);
or U6536 (N_6536,N_6300,N_6307);
nor U6537 (N_6537,N_6346,N_6277);
xnor U6538 (N_6538,N_6394,N_6219);
xnor U6539 (N_6539,N_6209,N_6241);
nand U6540 (N_6540,N_6380,N_6269);
nand U6541 (N_6541,N_6281,N_6395);
xnor U6542 (N_6542,N_6203,N_6219);
nand U6543 (N_6543,N_6316,N_6289);
and U6544 (N_6544,N_6263,N_6317);
and U6545 (N_6545,N_6292,N_6248);
and U6546 (N_6546,N_6380,N_6349);
nor U6547 (N_6547,N_6325,N_6384);
or U6548 (N_6548,N_6307,N_6329);
and U6549 (N_6549,N_6202,N_6300);
xor U6550 (N_6550,N_6206,N_6358);
nand U6551 (N_6551,N_6219,N_6243);
and U6552 (N_6552,N_6317,N_6391);
or U6553 (N_6553,N_6347,N_6333);
or U6554 (N_6554,N_6219,N_6301);
nand U6555 (N_6555,N_6396,N_6367);
xnor U6556 (N_6556,N_6302,N_6326);
xor U6557 (N_6557,N_6290,N_6209);
nor U6558 (N_6558,N_6397,N_6358);
and U6559 (N_6559,N_6274,N_6277);
or U6560 (N_6560,N_6391,N_6371);
xor U6561 (N_6561,N_6282,N_6377);
and U6562 (N_6562,N_6271,N_6363);
nor U6563 (N_6563,N_6392,N_6273);
xnor U6564 (N_6564,N_6296,N_6275);
and U6565 (N_6565,N_6266,N_6242);
nand U6566 (N_6566,N_6271,N_6349);
and U6567 (N_6567,N_6307,N_6202);
xnor U6568 (N_6568,N_6302,N_6363);
or U6569 (N_6569,N_6210,N_6250);
nand U6570 (N_6570,N_6296,N_6276);
nor U6571 (N_6571,N_6290,N_6306);
xnor U6572 (N_6572,N_6379,N_6218);
nor U6573 (N_6573,N_6324,N_6281);
or U6574 (N_6574,N_6364,N_6272);
nand U6575 (N_6575,N_6362,N_6236);
and U6576 (N_6576,N_6376,N_6317);
and U6577 (N_6577,N_6376,N_6214);
or U6578 (N_6578,N_6313,N_6305);
nor U6579 (N_6579,N_6360,N_6395);
nor U6580 (N_6580,N_6295,N_6360);
nor U6581 (N_6581,N_6229,N_6378);
nand U6582 (N_6582,N_6356,N_6346);
xnor U6583 (N_6583,N_6232,N_6303);
nand U6584 (N_6584,N_6201,N_6282);
or U6585 (N_6585,N_6384,N_6218);
nand U6586 (N_6586,N_6318,N_6391);
and U6587 (N_6587,N_6222,N_6330);
xnor U6588 (N_6588,N_6231,N_6283);
nor U6589 (N_6589,N_6250,N_6338);
xnor U6590 (N_6590,N_6213,N_6226);
nor U6591 (N_6591,N_6355,N_6274);
or U6592 (N_6592,N_6367,N_6383);
or U6593 (N_6593,N_6308,N_6226);
or U6594 (N_6594,N_6385,N_6244);
nor U6595 (N_6595,N_6288,N_6213);
nand U6596 (N_6596,N_6260,N_6281);
nand U6597 (N_6597,N_6283,N_6370);
and U6598 (N_6598,N_6286,N_6321);
nand U6599 (N_6599,N_6397,N_6243);
nand U6600 (N_6600,N_6577,N_6482);
nor U6601 (N_6601,N_6425,N_6462);
nor U6602 (N_6602,N_6555,N_6562);
xor U6603 (N_6603,N_6568,N_6532);
xnor U6604 (N_6604,N_6585,N_6563);
and U6605 (N_6605,N_6435,N_6493);
xor U6606 (N_6606,N_6521,N_6561);
nor U6607 (N_6607,N_6444,N_6420);
or U6608 (N_6608,N_6508,N_6450);
nand U6609 (N_6609,N_6431,N_6480);
and U6610 (N_6610,N_6457,N_6557);
nor U6611 (N_6611,N_6570,N_6433);
nor U6612 (N_6612,N_6459,N_6447);
nand U6613 (N_6613,N_6412,N_6426);
nor U6614 (N_6614,N_6583,N_6468);
and U6615 (N_6615,N_6408,N_6522);
or U6616 (N_6616,N_6591,N_6416);
nor U6617 (N_6617,N_6476,N_6576);
or U6618 (N_6618,N_6534,N_6463);
xor U6619 (N_6619,N_6401,N_6481);
and U6620 (N_6620,N_6547,N_6573);
nand U6621 (N_6621,N_6513,N_6439);
nand U6622 (N_6622,N_6597,N_6550);
and U6623 (N_6623,N_6467,N_6470);
or U6624 (N_6624,N_6473,N_6543);
and U6625 (N_6625,N_6486,N_6437);
and U6626 (N_6626,N_6432,N_6469);
xor U6627 (N_6627,N_6428,N_6478);
nor U6628 (N_6628,N_6490,N_6403);
and U6629 (N_6629,N_6545,N_6495);
and U6630 (N_6630,N_6539,N_6590);
or U6631 (N_6631,N_6596,N_6441);
nand U6632 (N_6632,N_6501,N_6558);
or U6633 (N_6633,N_6588,N_6564);
xnor U6634 (N_6634,N_6488,N_6525);
or U6635 (N_6635,N_6537,N_6536);
and U6636 (N_6636,N_6593,N_6592);
nand U6637 (N_6637,N_6524,N_6415);
nor U6638 (N_6638,N_6571,N_6454);
or U6639 (N_6639,N_6465,N_6578);
xnor U6640 (N_6640,N_6413,N_6580);
nor U6641 (N_6641,N_6498,N_6472);
xnor U6642 (N_6642,N_6560,N_6511);
nand U6643 (N_6643,N_6485,N_6402);
or U6644 (N_6644,N_6479,N_6448);
nor U6645 (N_6645,N_6567,N_6405);
nand U6646 (N_6646,N_6523,N_6527);
nor U6647 (N_6647,N_6579,N_6458);
or U6648 (N_6648,N_6507,N_6406);
xor U6649 (N_6649,N_6410,N_6400);
xor U6650 (N_6650,N_6506,N_6464);
nand U6651 (N_6651,N_6492,N_6526);
xor U6652 (N_6652,N_6535,N_6471);
nand U6653 (N_6653,N_6436,N_6540);
nand U6654 (N_6654,N_6422,N_6512);
or U6655 (N_6655,N_6499,N_6598);
nor U6656 (N_6656,N_6531,N_6461);
or U6657 (N_6657,N_6409,N_6418);
nor U6658 (N_6658,N_6419,N_6502);
xnor U6659 (N_6659,N_6446,N_6440);
nand U6660 (N_6660,N_6569,N_6553);
nor U6661 (N_6661,N_6589,N_6411);
or U6662 (N_6662,N_6452,N_6556);
nor U6663 (N_6663,N_6496,N_6594);
xor U6664 (N_6664,N_6491,N_6430);
nand U6665 (N_6665,N_6423,N_6504);
nand U6666 (N_6666,N_6404,N_6538);
xor U6667 (N_6667,N_6434,N_6574);
nand U6668 (N_6668,N_6587,N_6421);
xnor U6669 (N_6669,N_6505,N_6575);
nor U6670 (N_6670,N_6566,N_6520);
nor U6671 (N_6671,N_6429,N_6581);
nand U6672 (N_6672,N_6474,N_6466);
nor U6673 (N_6673,N_6509,N_6424);
nor U6674 (N_6674,N_6542,N_6497);
xnor U6675 (N_6675,N_6494,N_6586);
nor U6676 (N_6676,N_6453,N_6417);
nand U6677 (N_6677,N_6427,N_6443);
xor U6678 (N_6678,N_6442,N_6451);
or U6679 (N_6679,N_6500,N_6548);
nor U6680 (N_6680,N_6559,N_6414);
or U6681 (N_6681,N_6514,N_6530);
or U6682 (N_6682,N_6572,N_6518);
and U6683 (N_6683,N_6503,N_6565);
and U6684 (N_6684,N_6554,N_6541);
nand U6685 (N_6685,N_6484,N_6533);
nand U6686 (N_6686,N_6582,N_6599);
nor U6687 (N_6687,N_6544,N_6528);
nand U6688 (N_6688,N_6460,N_6489);
xor U6689 (N_6689,N_6475,N_6477);
and U6690 (N_6690,N_6455,N_6407);
nand U6691 (N_6691,N_6517,N_6487);
nand U6692 (N_6692,N_6445,N_6549);
and U6693 (N_6693,N_6515,N_6449);
nand U6694 (N_6694,N_6552,N_6529);
and U6695 (N_6695,N_6551,N_6438);
or U6696 (N_6696,N_6595,N_6483);
nor U6697 (N_6697,N_6510,N_6456);
or U6698 (N_6698,N_6546,N_6516);
or U6699 (N_6699,N_6519,N_6584);
nand U6700 (N_6700,N_6583,N_6585);
xnor U6701 (N_6701,N_6425,N_6437);
nand U6702 (N_6702,N_6569,N_6572);
nor U6703 (N_6703,N_6529,N_6520);
or U6704 (N_6704,N_6507,N_6562);
or U6705 (N_6705,N_6575,N_6536);
nand U6706 (N_6706,N_6523,N_6486);
nand U6707 (N_6707,N_6578,N_6445);
or U6708 (N_6708,N_6411,N_6557);
or U6709 (N_6709,N_6515,N_6439);
and U6710 (N_6710,N_6550,N_6475);
or U6711 (N_6711,N_6429,N_6409);
or U6712 (N_6712,N_6597,N_6451);
or U6713 (N_6713,N_6508,N_6583);
xor U6714 (N_6714,N_6443,N_6414);
xor U6715 (N_6715,N_6469,N_6588);
and U6716 (N_6716,N_6584,N_6595);
nand U6717 (N_6717,N_6423,N_6445);
xor U6718 (N_6718,N_6458,N_6514);
xor U6719 (N_6719,N_6535,N_6411);
or U6720 (N_6720,N_6599,N_6508);
or U6721 (N_6721,N_6510,N_6440);
xnor U6722 (N_6722,N_6412,N_6435);
nand U6723 (N_6723,N_6545,N_6483);
nor U6724 (N_6724,N_6544,N_6553);
and U6725 (N_6725,N_6406,N_6431);
xor U6726 (N_6726,N_6466,N_6453);
or U6727 (N_6727,N_6554,N_6413);
nor U6728 (N_6728,N_6430,N_6513);
or U6729 (N_6729,N_6576,N_6555);
xnor U6730 (N_6730,N_6581,N_6522);
nor U6731 (N_6731,N_6449,N_6516);
or U6732 (N_6732,N_6598,N_6469);
nor U6733 (N_6733,N_6419,N_6427);
and U6734 (N_6734,N_6497,N_6587);
xor U6735 (N_6735,N_6542,N_6501);
nand U6736 (N_6736,N_6524,N_6590);
xor U6737 (N_6737,N_6464,N_6471);
or U6738 (N_6738,N_6466,N_6567);
nor U6739 (N_6739,N_6577,N_6466);
nand U6740 (N_6740,N_6486,N_6451);
and U6741 (N_6741,N_6580,N_6447);
xnor U6742 (N_6742,N_6440,N_6428);
nand U6743 (N_6743,N_6531,N_6424);
xnor U6744 (N_6744,N_6425,N_6586);
xnor U6745 (N_6745,N_6499,N_6526);
nor U6746 (N_6746,N_6536,N_6521);
nand U6747 (N_6747,N_6555,N_6541);
xnor U6748 (N_6748,N_6544,N_6488);
and U6749 (N_6749,N_6492,N_6438);
or U6750 (N_6750,N_6553,N_6483);
nand U6751 (N_6751,N_6410,N_6548);
and U6752 (N_6752,N_6531,N_6542);
or U6753 (N_6753,N_6561,N_6455);
or U6754 (N_6754,N_6570,N_6590);
xnor U6755 (N_6755,N_6572,N_6452);
nor U6756 (N_6756,N_6412,N_6526);
xnor U6757 (N_6757,N_6531,N_6587);
and U6758 (N_6758,N_6407,N_6587);
nand U6759 (N_6759,N_6516,N_6584);
or U6760 (N_6760,N_6545,N_6547);
nor U6761 (N_6761,N_6576,N_6418);
nor U6762 (N_6762,N_6525,N_6448);
and U6763 (N_6763,N_6513,N_6405);
nand U6764 (N_6764,N_6565,N_6415);
or U6765 (N_6765,N_6525,N_6561);
and U6766 (N_6766,N_6582,N_6517);
or U6767 (N_6767,N_6410,N_6408);
nand U6768 (N_6768,N_6563,N_6503);
or U6769 (N_6769,N_6572,N_6447);
or U6770 (N_6770,N_6445,N_6580);
and U6771 (N_6771,N_6510,N_6491);
nor U6772 (N_6772,N_6555,N_6590);
or U6773 (N_6773,N_6593,N_6428);
and U6774 (N_6774,N_6415,N_6505);
nor U6775 (N_6775,N_6577,N_6541);
nand U6776 (N_6776,N_6553,N_6429);
nand U6777 (N_6777,N_6585,N_6468);
nand U6778 (N_6778,N_6407,N_6428);
or U6779 (N_6779,N_6406,N_6559);
nand U6780 (N_6780,N_6447,N_6569);
nand U6781 (N_6781,N_6501,N_6401);
or U6782 (N_6782,N_6551,N_6411);
xnor U6783 (N_6783,N_6469,N_6451);
or U6784 (N_6784,N_6435,N_6564);
nor U6785 (N_6785,N_6597,N_6429);
or U6786 (N_6786,N_6438,N_6515);
and U6787 (N_6787,N_6498,N_6413);
or U6788 (N_6788,N_6459,N_6429);
nand U6789 (N_6789,N_6582,N_6433);
nor U6790 (N_6790,N_6521,N_6424);
xnor U6791 (N_6791,N_6435,N_6549);
xor U6792 (N_6792,N_6541,N_6504);
nor U6793 (N_6793,N_6570,N_6561);
nor U6794 (N_6794,N_6516,N_6433);
nand U6795 (N_6795,N_6514,N_6569);
nand U6796 (N_6796,N_6512,N_6547);
nor U6797 (N_6797,N_6513,N_6512);
and U6798 (N_6798,N_6480,N_6579);
xnor U6799 (N_6799,N_6448,N_6480);
and U6800 (N_6800,N_6798,N_6677);
nand U6801 (N_6801,N_6741,N_6728);
nor U6802 (N_6802,N_6754,N_6774);
or U6803 (N_6803,N_6799,N_6647);
and U6804 (N_6804,N_6657,N_6616);
xor U6805 (N_6805,N_6795,N_6797);
or U6806 (N_6806,N_6701,N_6634);
and U6807 (N_6807,N_6679,N_6653);
nor U6808 (N_6808,N_6787,N_6695);
and U6809 (N_6809,N_6637,N_6716);
nand U6810 (N_6810,N_6625,N_6609);
nor U6811 (N_6811,N_6707,N_6640);
or U6812 (N_6812,N_6614,N_6711);
xor U6813 (N_6813,N_6789,N_6786);
nor U6814 (N_6814,N_6780,N_6708);
and U6815 (N_6815,N_6683,N_6706);
xor U6816 (N_6816,N_6796,N_6749);
or U6817 (N_6817,N_6750,N_6615);
nand U6818 (N_6818,N_6758,N_6639);
xor U6819 (N_6819,N_6671,N_6755);
xnor U6820 (N_6820,N_6793,N_6746);
or U6821 (N_6821,N_6610,N_6691);
or U6822 (N_6822,N_6654,N_6611);
nand U6823 (N_6823,N_6763,N_6629);
or U6824 (N_6824,N_6698,N_6676);
nor U6825 (N_6825,N_6794,N_6636);
nand U6826 (N_6826,N_6735,N_6792);
and U6827 (N_6827,N_6772,N_6688);
or U6828 (N_6828,N_6649,N_6700);
or U6829 (N_6829,N_6689,N_6773);
or U6830 (N_6830,N_6760,N_6705);
or U6831 (N_6831,N_6680,N_6696);
nor U6832 (N_6832,N_6681,N_6646);
nor U6833 (N_6833,N_6608,N_6764);
and U6834 (N_6834,N_6778,N_6694);
nand U6835 (N_6835,N_6783,N_6687);
xnor U6836 (N_6836,N_6659,N_6630);
or U6837 (N_6837,N_6748,N_6651);
nand U6838 (N_6838,N_6620,N_6600);
nand U6839 (N_6839,N_6785,N_6712);
and U6840 (N_6840,N_6660,N_6720);
xnor U6841 (N_6841,N_6734,N_6624);
xnor U6842 (N_6842,N_6684,N_6726);
nand U6843 (N_6843,N_6658,N_6751);
or U6844 (N_6844,N_6784,N_6648);
or U6845 (N_6845,N_6669,N_6638);
or U6846 (N_6846,N_6767,N_6723);
nand U6847 (N_6847,N_6752,N_6673);
nor U6848 (N_6848,N_6775,N_6790);
xnor U6849 (N_6849,N_6744,N_6622);
and U6850 (N_6850,N_6612,N_6631);
and U6851 (N_6851,N_6766,N_6656);
nor U6852 (N_6852,N_6633,N_6663);
nor U6853 (N_6853,N_6777,N_6642);
xnor U6854 (N_6854,N_6718,N_6729);
nor U6855 (N_6855,N_6661,N_6645);
nor U6856 (N_6856,N_6621,N_6674);
nand U6857 (N_6857,N_6655,N_6740);
nand U6858 (N_6858,N_6601,N_6666);
and U6859 (N_6859,N_6628,N_6686);
or U6860 (N_6860,N_6664,N_6724);
and U6861 (N_6861,N_6690,N_6675);
or U6862 (N_6862,N_6733,N_6714);
nand U6863 (N_6863,N_6682,N_6619);
xnor U6864 (N_6864,N_6769,N_6779);
and U6865 (N_6865,N_6672,N_6721);
or U6866 (N_6866,N_6770,N_6670);
nand U6867 (N_6867,N_6730,N_6713);
and U6868 (N_6868,N_6737,N_6722);
nand U6869 (N_6869,N_6644,N_6791);
nor U6870 (N_6870,N_6715,N_6709);
and U6871 (N_6871,N_6776,N_6788);
xnor U6872 (N_6872,N_6736,N_6635);
nand U6873 (N_6873,N_6727,N_6604);
nor U6874 (N_6874,N_6692,N_6743);
nand U6875 (N_6875,N_6699,N_6665);
nor U6876 (N_6876,N_6765,N_6602);
nand U6877 (N_6877,N_6753,N_6782);
nor U6878 (N_6878,N_6747,N_6626);
nor U6879 (N_6879,N_6667,N_6739);
xnor U6880 (N_6880,N_6781,N_6759);
or U6881 (N_6881,N_6606,N_6756);
or U6882 (N_6882,N_6643,N_6702);
and U6883 (N_6883,N_6668,N_6607);
or U6884 (N_6884,N_6685,N_6704);
and U6885 (N_6885,N_6632,N_6771);
and U6886 (N_6886,N_6650,N_6617);
xnor U6887 (N_6887,N_6768,N_6662);
nor U6888 (N_6888,N_6717,N_6693);
nand U6889 (N_6889,N_6603,N_6762);
nor U6890 (N_6890,N_6703,N_6627);
nand U6891 (N_6891,N_6641,N_6761);
and U6892 (N_6892,N_6605,N_6710);
nor U6893 (N_6893,N_6745,N_6678);
nor U6894 (N_6894,N_6719,N_6652);
and U6895 (N_6895,N_6618,N_6725);
nand U6896 (N_6896,N_6732,N_6731);
and U6897 (N_6897,N_6742,N_6697);
xnor U6898 (N_6898,N_6757,N_6613);
and U6899 (N_6899,N_6623,N_6738);
nand U6900 (N_6900,N_6713,N_6683);
xnor U6901 (N_6901,N_6635,N_6697);
xnor U6902 (N_6902,N_6731,N_6650);
and U6903 (N_6903,N_6795,N_6651);
and U6904 (N_6904,N_6691,N_6659);
nor U6905 (N_6905,N_6708,N_6716);
and U6906 (N_6906,N_6637,N_6777);
or U6907 (N_6907,N_6607,N_6673);
nor U6908 (N_6908,N_6605,N_6602);
nand U6909 (N_6909,N_6747,N_6714);
xnor U6910 (N_6910,N_6680,N_6631);
nor U6911 (N_6911,N_6746,N_6684);
xnor U6912 (N_6912,N_6615,N_6673);
or U6913 (N_6913,N_6680,N_6727);
xor U6914 (N_6914,N_6679,N_6721);
or U6915 (N_6915,N_6753,N_6749);
nand U6916 (N_6916,N_6714,N_6795);
nand U6917 (N_6917,N_6642,N_6671);
nand U6918 (N_6918,N_6700,N_6621);
or U6919 (N_6919,N_6671,N_6686);
or U6920 (N_6920,N_6743,N_6751);
nand U6921 (N_6921,N_6756,N_6750);
and U6922 (N_6922,N_6685,N_6787);
xnor U6923 (N_6923,N_6729,N_6704);
nand U6924 (N_6924,N_6710,N_6614);
or U6925 (N_6925,N_6727,N_6754);
or U6926 (N_6926,N_6623,N_6726);
nor U6927 (N_6927,N_6766,N_6792);
nand U6928 (N_6928,N_6721,N_6749);
and U6929 (N_6929,N_6674,N_6643);
nand U6930 (N_6930,N_6690,N_6668);
or U6931 (N_6931,N_6766,N_6650);
and U6932 (N_6932,N_6677,N_6779);
xor U6933 (N_6933,N_6771,N_6758);
nand U6934 (N_6934,N_6678,N_6718);
nor U6935 (N_6935,N_6751,N_6752);
or U6936 (N_6936,N_6656,N_6769);
nor U6937 (N_6937,N_6632,N_6787);
xor U6938 (N_6938,N_6669,N_6694);
and U6939 (N_6939,N_6765,N_6613);
or U6940 (N_6940,N_6725,N_6710);
nand U6941 (N_6941,N_6780,N_6677);
or U6942 (N_6942,N_6792,N_6731);
nand U6943 (N_6943,N_6672,N_6788);
nor U6944 (N_6944,N_6743,N_6747);
nor U6945 (N_6945,N_6780,N_6646);
nor U6946 (N_6946,N_6708,N_6742);
xor U6947 (N_6947,N_6751,N_6795);
nor U6948 (N_6948,N_6675,N_6797);
and U6949 (N_6949,N_6796,N_6726);
nand U6950 (N_6950,N_6605,N_6649);
nand U6951 (N_6951,N_6611,N_6744);
nand U6952 (N_6952,N_6646,N_6761);
and U6953 (N_6953,N_6679,N_6745);
nand U6954 (N_6954,N_6792,N_6637);
and U6955 (N_6955,N_6708,N_6628);
and U6956 (N_6956,N_6745,N_6736);
xnor U6957 (N_6957,N_6694,N_6642);
nor U6958 (N_6958,N_6663,N_6643);
and U6959 (N_6959,N_6739,N_6636);
xor U6960 (N_6960,N_6714,N_6650);
and U6961 (N_6961,N_6696,N_6779);
or U6962 (N_6962,N_6778,N_6789);
and U6963 (N_6963,N_6680,N_6608);
or U6964 (N_6964,N_6723,N_6734);
or U6965 (N_6965,N_6697,N_6727);
or U6966 (N_6966,N_6679,N_6618);
xor U6967 (N_6967,N_6797,N_6759);
nor U6968 (N_6968,N_6715,N_6797);
nand U6969 (N_6969,N_6602,N_6624);
or U6970 (N_6970,N_6607,N_6757);
or U6971 (N_6971,N_6690,N_6770);
and U6972 (N_6972,N_6730,N_6681);
and U6973 (N_6973,N_6627,N_6717);
nor U6974 (N_6974,N_6676,N_6701);
xor U6975 (N_6975,N_6718,N_6685);
or U6976 (N_6976,N_6794,N_6624);
nor U6977 (N_6977,N_6679,N_6626);
nor U6978 (N_6978,N_6762,N_6675);
or U6979 (N_6979,N_6779,N_6782);
or U6980 (N_6980,N_6735,N_6760);
xnor U6981 (N_6981,N_6715,N_6748);
nor U6982 (N_6982,N_6765,N_6768);
nor U6983 (N_6983,N_6641,N_6617);
xor U6984 (N_6984,N_6733,N_6621);
nand U6985 (N_6985,N_6637,N_6672);
or U6986 (N_6986,N_6749,N_6653);
or U6987 (N_6987,N_6607,N_6653);
nor U6988 (N_6988,N_6697,N_6658);
and U6989 (N_6989,N_6647,N_6766);
nor U6990 (N_6990,N_6624,N_6629);
xnor U6991 (N_6991,N_6662,N_6623);
and U6992 (N_6992,N_6790,N_6686);
nand U6993 (N_6993,N_6702,N_6764);
and U6994 (N_6994,N_6649,N_6688);
nand U6995 (N_6995,N_6673,N_6743);
or U6996 (N_6996,N_6689,N_6603);
or U6997 (N_6997,N_6770,N_6730);
xnor U6998 (N_6998,N_6756,N_6700);
nand U6999 (N_6999,N_6607,N_6762);
nor U7000 (N_7000,N_6974,N_6937);
and U7001 (N_7001,N_6812,N_6986);
or U7002 (N_7002,N_6887,N_6818);
xnor U7003 (N_7003,N_6927,N_6824);
nand U7004 (N_7004,N_6869,N_6973);
nor U7005 (N_7005,N_6836,N_6923);
and U7006 (N_7006,N_6977,N_6805);
and U7007 (N_7007,N_6944,N_6890);
and U7008 (N_7008,N_6933,N_6826);
and U7009 (N_7009,N_6953,N_6823);
and U7010 (N_7010,N_6985,N_6817);
nor U7011 (N_7011,N_6811,N_6930);
or U7012 (N_7012,N_6881,N_6931);
or U7013 (N_7013,N_6911,N_6848);
xor U7014 (N_7014,N_6880,N_6834);
or U7015 (N_7015,N_6904,N_6903);
nor U7016 (N_7016,N_6987,N_6947);
nand U7017 (N_7017,N_6878,N_6963);
nand U7018 (N_7018,N_6981,N_6926);
xnor U7019 (N_7019,N_6957,N_6896);
nand U7020 (N_7020,N_6830,N_6821);
nor U7021 (N_7021,N_6858,N_6807);
nor U7022 (N_7022,N_6841,N_6813);
nor U7023 (N_7023,N_6932,N_6897);
or U7024 (N_7024,N_6856,N_6980);
and U7025 (N_7025,N_6968,N_6967);
and U7026 (N_7026,N_6855,N_6803);
and U7027 (N_7027,N_6820,N_6901);
xnor U7028 (N_7028,N_6994,N_6894);
xor U7029 (N_7029,N_6842,N_6915);
and U7030 (N_7030,N_6882,N_6935);
or U7031 (N_7031,N_6966,N_6867);
xor U7032 (N_7032,N_6802,N_6800);
xnor U7033 (N_7033,N_6877,N_6833);
and U7034 (N_7034,N_6857,N_6819);
or U7035 (N_7035,N_6845,N_6879);
nor U7036 (N_7036,N_6846,N_6864);
xor U7037 (N_7037,N_6874,N_6950);
xor U7038 (N_7038,N_6888,N_6847);
nor U7039 (N_7039,N_6893,N_6989);
nor U7040 (N_7040,N_6892,N_6899);
and U7041 (N_7041,N_6865,N_6815);
xor U7042 (N_7042,N_6850,N_6969);
nor U7043 (N_7043,N_6993,N_6891);
and U7044 (N_7044,N_6808,N_6999);
nand U7045 (N_7045,N_6851,N_6921);
nand U7046 (N_7046,N_6934,N_6996);
nand U7047 (N_7047,N_6884,N_6984);
or U7048 (N_7048,N_6804,N_6943);
or U7049 (N_7049,N_6849,N_6922);
nand U7050 (N_7050,N_6801,N_6941);
or U7051 (N_7051,N_6837,N_6936);
nand U7052 (N_7052,N_6997,N_6990);
nand U7053 (N_7053,N_6972,N_6832);
nand U7054 (N_7054,N_6952,N_6955);
and U7055 (N_7055,N_6853,N_6942);
or U7056 (N_7056,N_6983,N_6860);
or U7057 (N_7057,N_6866,N_6909);
and U7058 (N_7058,N_6905,N_6886);
and U7059 (N_7059,N_6924,N_6914);
xnor U7060 (N_7060,N_6954,N_6814);
nand U7061 (N_7061,N_6902,N_6960);
nand U7062 (N_7062,N_6844,N_6920);
or U7063 (N_7063,N_6859,N_6965);
nor U7064 (N_7064,N_6863,N_6883);
and U7065 (N_7065,N_6908,N_6948);
xor U7066 (N_7066,N_6828,N_6907);
nand U7067 (N_7067,N_6995,N_6939);
xor U7068 (N_7068,N_6962,N_6918);
nand U7069 (N_7069,N_6889,N_6991);
xnor U7070 (N_7070,N_6919,N_6916);
or U7071 (N_7071,N_6843,N_6979);
and U7072 (N_7072,N_6852,N_6970);
nand U7073 (N_7073,N_6825,N_6872);
xnor U7074 (N_7074,N_6861,N_6839);
and U7075 (N_7075,N_6925,N_6998);
nand U7076 (N_7076,N_6810,N_6978);
nand U7077 (N_7077,N_6871,N_6835);
xnor U7078 (N_7078,N_6917,N_6868);
xor U7079 (N_7079,N_6900,N_6898);
and U7080 (N_7080,N_6940,N_6971);
nand U7081 (N_7081,N_6876,N_6875);
nand U7082 (N_7082,N_6928,N_6929);
nor U7083 (N_7083,N_6951,N_6912);
and U7084 (N_7084,N_6809,N_6831);
or U7085 (N_7085,N_6827,N_6946);
or U7086 (N_7086,N_6829,N_6885);
or U7087 (N_7087,N_6906,N_6959);
or U7088 (N_7088,N_6958,N_6949);
nor U7089 (N_7089,N_6976,N_6982);
or U7090 (N_7090,N_6870,N_6964);
and U7091 (N_7091,N_6913,N_6910);
and U7092 (N_7092,N_6992,N_6988);
and U7093 (N_7093,N_6961,N_6956);
nor U7094 (N_7094,N_6838,N_6895);
or U7095 (N_7095,N_6822,N_6806);
nor U7096 (N_7096,N_6840,N_6862);
and U7097 (N_7097,N_6816,N_6854);
or U7098 (N_7098,N_6938,N_6873);
nand U7099 (N_7099,N_6975,N_6945);
nand U7100 (N_7100,N_6840,N_6879);
or U7101 (N_7101,N_6854,N_6908);
xnor U7102 (N_7102,N_6985,N_6907);
xnor U7103 (N_7103,N_6825,N_6988);
or U7104 (N_7104,N_6853,N_6875);
or U7105 (N_7105,N_6973,N_6944);
nor U7106 (N_7106,N_6938,N_6957);
xnor U7107 (N_7107,N_6848,N_6947);
or U7108 (N_7108,N_6876,N_6848);
nor U7109 (N_7109,N_6966,N_6854);
nor U7110 (N_7110,N_6900,N_6957);
nor U7111 (N_7111,N_6933,N_6847);
nor U7112 (N_7112,N_6840,N_6903);
xnor U7113 (N_7113,N_6966,N_6964);
and U7114 (N_7114,N_6994,N_6811);
nor U7115 (N_7115,N_6883,N_6989);
xor U7116 (N_7116,N_6963,N_6859);
nor U7117 (N_7117,N_6839,N_6989);
nor U7118 (N_7118,N_6806,N_6891);
nor U7119 (N_7119,N_6886,N_6806);
and U7120 (N_7120,N_6961,N_6806);
and U7121 (N_7121,N_6989,N_6801);
nand U7122 (N_7122,N_6965,N_6837);
nor U7123 (N_7123,N_6975,N_6839);
xor U7124 (N_7124,N_6899,N_6850);
and U7125 (N_7125,N_6964,N_6984);
and U7126 (N_7126,N_6919,N_6826);
xor U7127 (N_7127,N_6815,N_6876);
and U7128 (N_7128,N_6931,N_6867);
xnor U7129 (N_7129,N_6947,N_6808);
nor U7130 (N_7130,N_6986,N_6955);
xor U7131 (N_7131,N_6894,N_6851);
xnor U7132 (N_7132,N_6896,N_6815);
and U7133 (N_7133,N_6924,N_6995);
nor U7134 (N_7134,N_6849,N_6815);
and U7135 (N_7135,N_6844,N_6851);
nor U7136 (N_7136,N_6988,N_6959);
nand U7137 (N_7137,N_6809,N_6916);
or U7138 (N_7138,N_6859,N_6864);
xor U7139 (N_7139,N_6998,N_6909);
or U7140 (N_7140,N_6923,N_6936);
and U7141 (N_7141,N_6821,N_6902);
or U7142 (N_7142,N_6993,N_6839);
and U7143 (N_7143,N_6876,N_6860);
xor U7144 (N_7144,N_6905,N_6884);
nand U7145 (N_7145,N_6979,N_6901);
xnor U7146 (N_7146,N_6921,N_6878);
nand U7147 (N_7147,N_6805,N_6941);
nand U7148 (N_7148,N_6861,N_6942);
or U7149 (N_7149,N_6830,N_6935);
or U7150 (N_7150,N_6864,N_6832);
xor U7151 (N_7151,N_6855,N_6839);
nor U7152 (N_7152,N_6880,N_6897);
nand U7153 (N_7153,N_6993,N_6994);
xor U7154 (N_7154,N_6947,N_6906);
or U7155 (N_7155,N_6986,N_6881);
nand U7156 (N_7156,N_6812,N_6999);
xor U7157 (N_7157,N_6806,N_6916);
or U7158 (N_7158,N_6810,N_6963);
nor U7159 (N_7159,N_6816,N_6813);
xor U7160 (N_7160,N_6931,N_6846);
nand U7161 (N_7161,N_6861,N_6927);
nand U7162 (N_7162,N_6834,N_6995);
or U7163 (N_7163,N_6872,N_6939);
and U7164 (N_7164,N_6824,N_6919);
or U7165 (N_7165,N_6994,N_6956);
nor U7166 (N_7166,N_6838,N_6827);
or U7167 (N_7167,N_6977,N_6989);
or U7168 (N_7168,N_6893,N_6866);
xnor U7169 (N_7169,N_6835,N_6836);
nor U7170 (N_7170,N_6943,N_6873);
xor U7171 (N_7171,N_6970,N_6950);
nand U7172 (N_7172,N_6841,N_6878);
xor U7173 (N_7173,N_6879,N_6872);
nor U7174 (N_7174,N_6997,N_6861);
xnor U7175 (N_7175,N_6824,N_6810);
and U7176 (N_7176,N_6814,N_6870);
and U7177 (N_7177,N_6800,N_6820);
nor U7178 (N_7178,N_6953,N_6858);
nand U7179 (N_7179,N_6816,N_6843);
or U7180 (N_7180,N_6949,N_6847);
and U7181 (N_7181,N_6880,N_6971);
or U7182 (N_7182,N_6834,N_6811);
nand U7183 (N_7183,N_6817,N_6814);
or U7184 (N_7184,N_6920,N_6831);
nor U7185 (N_7185,N_6939,N_6862);
or U7186 (N_7186,N_6997,N_6945);
nand U7187 (N_7187,N_6972,N_6992);
nand U7188 (N_7188,N_6930,N_6869);
and U7189 (N_7189,N_6879,N_6949);
xor U7190 (N_7190,N_6990,N_6917);
xor U7191 (N_7191,N_6907,N_6834);
or U7192 (N_7192,N_6852,N_6836);
nor U7193 (N_7193,N_6938,N_6801);
or U7194 (N_7194,N_6869,N_6976);
and U7195 (N_7195,N_6842,N_6980);
nor U7196 (N_7196,N_6840,N_6898);
or U7197 (N_7197,N_6883,N_6841);
nor U7198 (N_7198,N_6843,N_6813);
nand U7199 (N_7199,N_6949,N_6887);
and U7200 (N_7200,N_7183,N_7100);
and U7201 (N_7201,N_7194,N_7175);
and U7202 (N_7202,N_7158,N_7148);
nand U7203 (N_7203,N_7163,N_7085);
or U7204 (N_7204,N_7076,N_7139);
xor U7205 (N_7205,N_7053,N_7147);
nor U7206 (N_7206,N_7131,N_7047);
and U7207 (N_7207,N_7149,N_7021);
xor U7208 (N_7208,N_7181,N_7126);
or U7209 (N_7209,N_7050,N_7162);
nand U7210 (N_7210,N_7055,N_7135);
and U7211 (N_7211,N_7015,N_7026);
or U7212 (N_7212,N_7129,N_7013);
nor U7213 (N_7213,N_7169,N_7111);
and U7214 (N_7214,N_7114,N_7193);
nor U7215 (N_7215,N_7065,N_7109);
or U7216 (N_7216,N_7187,N_7003);
xnor U7217 (N_7217,N_7098,N_7096);
and U7218 (N_7218,N_7144,N_7033);
nor U7219 (N_7219,N_7080,N_7006);
nor U7220 (N_7220,N_7072,N_7086);
or U7221 (N_7221,N_7171,N_7097);
nor U7222 (N_7222,N_7095,N_7176);
xor U7223 (N_7223,N_7174,N_7068);
and U7224 (N_7224,N_7010,N_7115);
nor U7225 (N_7225,N_7060,N_7164);
nand U7226 (N_7226,N_7107,N_7110);
or U7227 (N_7227,N_7178,N_7127);
nand U7228 (N_7228,N_7099,N_7198);
nor U7229 (N_7229,N_7014,N_7113);
nand U7230 (N_7230,N_7027,N_7190);
and U7231 (N_7231,N_7039,N_7069);
nand U7232 (N_7232,N_7035,N_7005);
nor U7233 (N_7233,N_7136,N_7017);
and U7234 (N_7234,N_7002,N_7157);
nand U7235 (N_7235,N_7121,N_7091);
xor U7236 (N_7236,N_7062,N_7106);
or U7237 (N_7237,N_7189,N_7167);
nand U7238 (N_7238,N_7061,N_7192);
nor U7239 (N_7239,N_7092,N_7152);
or U7240 (N_7240,N_7087,N_7078);
nor U7241 (N_7241,N_7140,N_7036);
nand U7242 (N_7242,N_7019,N_7191);
nand U7243 (N_7243,N_7022,N_7154);
and U7244 (N_7244,N_7004,N_7089);
nand U7245 (N_7245,N_7074,N_7030);
nor U7246 (N_7246,N_7180,N_7051);
nor U7247 (N_7247,N_7008,N_7123);
nand U7248 (N_7248,N_7186,N_7031);
xor U7249 (N_7249,N_7168,N_7138);
and U7250 (N_7250,N_7199,N_7116);
or U7251 (N_7251,N_7046,N_7119);
nor U7252 (N_7252,N_7182,N_7082);
nor U7253 (N_7253,N_7172,N_7128);
nand U7254 (N_7254,N_7118,N_7101);
nand U7255 (N_7255,N_7049,N_7064);
and U7256 (N_7256,N_7040,N_7038);
or U7257 (N_7257,N_7103,N_7052);
nand U7258 (N_7258,N_7108,N_7023);
nand U7259 (N_7259,N_7028,N_7009);
and U7260 (N_7260,N_7112,N_7122);
and U7261 (N_7261,N_7153,N_7161);
or U7262 (N_7262,N_7067,N_7124);
nand U7263 (N_7263,N_7073,N_7104);
nand U7264 (N_7264,N_7084,N_7025);
nand U7265 (N_7265,N_7081,N_7133);
nand U7266 (N_7266,N_7043,N_7054);
or U7267 (N_7267,N_7090,N_7141);
nand U7268 (N_7268,N_7057,N_7024);
or U7269 (N_7269,N_7155,N_7173);
xnor U7270 (N_7270,N_7029,N_7156);
xor U7271 (N_7271,N_7137,N_7120);
or U7272 (N_7272,N_7132,N_7071);
or U7273 (N_7273,N_7146,N_7196);
or U7274 (N_7274,N_7037,N_7032);
and U7275 (N_7275,N_7184,N_7170);
xnor U7276 (N_7276,N_7079,N_7011);
xor U7277 (N_7277,N_7125,N_7056);
xnor U7278 (N_7278,N_7177,N_7000);
or U7279 (N_7279,N_7020,N_7018);
xnor U7280 (N_7280,N_7083,N_7143);
nor U7281 (N_7281,N_7145,N_7166);
and U7282 (N_7282,N_7077,N_7188);
nor U7283 (N_7283,N_7041,N_7070);
and U7284 (N_7284,N_7093,N_7048);
xnor U7285 (N_7285,N_7130,N_7160);
nor U7286 (N_7286,N_7134,N_7105);
and U7287 (N_7287,N_7016,N_7102);
xor U7288 (N_7288,N_7165,N_7012);
nand U7289 (N_7289,N_7007,N_7034);
and U7290 (N_7290,N_7151,N_7075);
and U7291 (N_7291,N_7058,N_7045);
nand U7292 (N_7292,N_7066,N_7094);
nand U7293 (N_7293,N_7117,N_7150);
xnor U7294 (N_7294,N_7001,N_7195);
xnor U7295 (N_7295,N_7042,N_7159);
nor U7296 (N_7296,N_7088,N_7063);
or U7297 (N_7297,N_7142,N_7197);
and U7298 (N_7298,N_7185,N_7044);
and U7299 (N_7299,N_7059,N_7179);
nand U7300 (N_7300,N_7138,N_7072);
nor U7301 (N_7301,N_7167,N_7073);
nand U7302 (N_7302,N_7157,N_7149);
and U7303 (N_7303,N_7092,N_7055);
or U7304 (N_7304,N_7054,N_7052);
nand U7305 (N_7305,N_7001,N_7077);
xnor U7306 (N_7306,N_7152,N_7106);
or U7307 (N_7307,N_7170,N_7090);
or U7308 (N_7308,N_7189,N_7077);
nor U7309 (N_7309,N_7104,N_7087);
nand U7310 (N_7310,N_7126,N_7089);
xnor U7311 (N_7311,N_7113,N_7171);
nor U7312 (N_7312,N_7142,N_7075);
and U7313 (N_7313,N_7062,N_7098);
xor U7314 (N_7314,N_7084,N_7170);
nor U7315 (N_7315,N_7033,N_7114);
nand U7316 (N_7316,N_7106,N_7127);
and U7317 (N_7317,N_7174,N_7035);
nand U7318 (N_7318,N_7182,N_7131);
or U7319 (N_7319,N_7185,N_7096);
and U7320 (N_7320,N_7134,N_7067);
nor U7321 (N_7321,N_7199,N_7003);
and U7322 (N_7322,N_7131,N_7099);
nand U7323 (N_7323,N_7132,N_7171);
xnor U7324 (N_7324,N_7140,N_7097);
and U7325 (N_7325,N_7153,N_7174);
or U7326 (N_7326,N_7050,N_7033);
or U7327 (N_7327,N_7174,N_7181);
or U7328 (N_7328,N_7162,N_7048);
and U7329 (N_7329,N_7105,N_7002);
nor U7330 (N_7330,N_7045,N_7101);
and U7331 (N_7331,N_7080,N_7197);
xnor U7332 (N_7332,N_7130,N_7136);
and U7333 (N_7333,N_7067,N_7165);
or U7334 (N_7334,N_7015,N_7153);
nand U7335 (N_7335,N_7042,N_7069);
nand U7336 (N_7336,N_7192,N_7069);
nor U7337 (N_7337,N_7140,N_7069);
nor U7338 (N_7338,N_7166,N_7026);
or U7339 (N_7339,N_7007,N_7155);
and U7340 (N_7340,N_7002,N_7062);
nand U7341 (N_7341,N_7033,N_7020);
nor U7342 (N_7342,N_7027,N_7197);
nor U7343 (N_7343,N_7014,N_7184);
nand U7344 (N_7344,N_7192,N_7153);
xnor U7345 (N_7345,N_7110,N_7079);
xor U7346 (N_7346,N_7020,N_7195);
or U7347 (N_7347,N_7034,N_7053);
and U7348 (N_7348,N_7095,N_7043);
nand U7349 (N_7349,N_7033,N_7123);
xor U7350 (N_7350,N_7058,N_7091);
xor U7351 (N_7351,N_7131,N_7080);
or U7352 (N_7352,N_7104,N_7068);
or U7353 (N_7353,N_7023,N_7171);
nor U7354 (N_7354,N_7042,N_7182);
xnor U7355 (N_7355,N_7079,N_7119);
nor U7356 (N_7356,N_7181,N_7185);
nor U7357 (N_7357,N_7105,N_7057);
or U7358 (N_7358,N_7095,N_7188);
nor U7359 (N_7359,N_7078,N_7009);
or U7360 (N_7360,N_7120,N_7141);
or U7361 (N_7361,N_7082,N_7141);
nand U7362 (N_7362,N_7086,N_7132);
or U7363 (N_7363,N_7044,N_7102);
xnor U7364 (N_7364,N_7002,N_7055);
nor U7365 (N_7365,N_7045,N_7196);
nor U7366 (N_7366,N_7154,N_7004);
nor U7367 (N_7367,N_7104,N_7054);
xor U7368 (N_7368,N_7029,N_7190);
nand U7369 (N_7369,N_7094,N_7008);
nor U7370 (N_7370,N_7191,N_7055);
nand U7371 (N_7371,N_7174,N_7023);
or U7372 (N_7372,N_7147,N_7195);
nand U7373 (N_7373,N_7052,N_7135);
xor U7374 (N_7374,N_7135,N_7065);
or U7375 (N_7375,N_7045,N_7026);
xnor U7376 (N_7376,N_7004,N_7188);
nor U7377 (N_7377,N_7188,N_7087);
and U7378 (N_7378,N_7009,N_7019);
xor U7379 (N_7379,N_7154,N_7143);
or U7380 (N_7380,N_7143,N_7073);
and U7381 (N_7381,N_7184,N_7010);
nor U7382 (N_7382,N_7090,N_7133);
xnor U7383 (N_7383,N_7167,N_7120);
nand U7384 (N_7384,N_7048,N_7137);
or U7385 (N_7385,N_7124,N_7043);
or U7386 (N_7386,N_7170,N_7093);
xor U7387 (N_7387,N_7012,N_7198);
xor U7388 (N_7388,N_7199,N_7184);
and U7389 (N_7389,N_7163,N_7132);
nand U7390 (N_7390,N_7091,N_7086);
nor U7391 (N_7391,N_7140,N_7076);
and U7392 (N_7392,N_7123,N_7186);
or U7393 (N_7393,N_7158,N_7084);
nor U7394 (N_7394,N_7050,N_7090);
nor U7395 (N_7395,N_7055,N_7115);
xor U7396 (N_7396,N_7196,N_7127);
nand U7397 (N_7397,N_7109,N_7035);
nor U7398 (N_7398,N_7185,N_7182);
nand U7399 (N_7399,N_7057,N_7132);
xnor U7400 (N_7400,N_7208,N_7285);
nor U7401 (N_7401,N_7348,N_7366);
or U7402 (N_7402,N_7313,N_7314);
or U7403 (N_7403,N_7259,N_7280);
nand U7404 (N_7404,N_7257,N_7269);
or U7405 (N_7405,N_7340,N_7263);
nor U7406 (N_7406,N_7350,N_7364);
or U7407 (N_7407,N_7270,N_7338);
nand U7408 (N_7408,N_7223,N_7321);
nand U7409 (N_7409,N_7351,N_7382);
or U7410 (N_7410,N_7336,N_7297);
or U7411 (N_7411,N_7346,N_7354);
nand U7412 (N_7412,N_7323,N_7214);
nand U7413 (N_7413,N_7272,N_7247);
nor U7414 (N_7414,N_7282,N_7389);
nand U7415 (N_7415,N_7217,N_7376);
xnor U7416 (N_7416,N_7365,N_7300);
nor U7417 (N_7417,N_7238,N_7316);
nor U7418 (N_7418,N_7248,N_7250);
and U7419 (N_7419,N_7254,N_7356);
or U7420 (N_7420,N_7202,N_7230);
xor U7421 (N_7421,N_7375,N_7304);
and U7422 (N_7422,N_7265,N_7312);
nand U7423 (N_7423,N_7395,N_7324);
or U7424 (N_7424,N_7372,N_7262);
xnor U7425 (N_7425,N_7240,N_7251);
nand U7426 (N_7426,N_7319,N_7347);
nand U7427 (N_7427,N_7204,N_7311);
xnor U7428 (N_7428,N_7201,N_7349);
or U7429 (N_7429,N_7268,N_7390);
nand U7430 (N_7430,N_7246,N_7241);
or U7431 (N_7431,N_7235,N_7333);
and U7432 (N_7432,N_7374,N_7218);
nor U7433 (N_7433,N_7305,N_7275);
and U7434 (N_7434,N_7306,N_7233);
nor U7435 (N_7435,N_7224,N_7289);
nor U7436 (N_7436,N_7363,N_7332);
nor U7437 (N_7437,N_7274,N_7331);
or U7438 (N_7438,N_7264,N_7357);
or U7439 (N_7439,N_7337,N_7371);
nor U7440 (N_7440,N_7380,N_7244);
or U7441 (N_7441,N_7271,N_7373);
xor U7442 (N_7442,N_7277,N_7384);
xor U7443 (N_7443,N_7237,N_7386);
nand U7444 (N_7444,N_7385,N_7294);
or U7445 (N_7445,N_7261,N_7392);
xor U7446 (N_7446,N_7253,N_7362);
or U7447 (N_7447,N_7369,N_7358);
or U7448 (N_7448,N_7288,N_7236);
nand U7449 (N_7449,N_7360,N_7210);
or U7450 (N_7450,N_7342,N_7242);
or U7451 (N_7451,N_7334,N_7281);
nand U7452 (N_7452,N_7291,N_7229);
nor U7453 (N_7453,N_7231,N_7205);
or U7454 (N_7454,N_7326,N_7227);
and U7455 (N_7455,N_7345,N_7370);
xnor U7456 (N_7456,N_7381,N_7212);
nor U7457 (N_7457,N_7325,N_7317);
and U7458 (N_7458,N_7209,N_7252);
or U7459 (N_7459,N_7222,N_7255);
xor U7460 (N_7460,N_7328,N_7399);
and U7461 (N_7461,N_7391,N_7207);
nand U7462 (N_7462,N_7388,N_7387);
xnor U7463 (N_7463,N_7303,N_7213);
xnor U7464 (N_7464,N_7343,N_7279);
or U7465 (N_7465,N_7308,N_7302);
and U7466 (N_7466,N_7367,N_7393);
or U7467 (N_7467,N_7341,N_7301);
nand U7468 (N_7468,N_7234,N_7226);
and U7469 (N_7469,N_7245,N_7266);
xor U7470 (N_7470,N_7339,N_7377);
and U7471 (N_7471,N_7273,N_7203);
nor U7472 (N_7472,N_7287,N_7322);
or U7473 (N_7473,N_7307,N_7327);
xnor U7474 (N_7474,N_7200,N_7355);
and U7475 (N_7475,N_7215,N_7335);
or U7476 (N_7476,N_7396,N_7292);
and U7477 (N_7477,N_7318,N_7359);
or U7478 (N_7478,N_7276,N_7368);
nor U7479 (N_7479,N_7284,N_7397);
nor U7480 (N_7480,N_7353,N_7239);
and U7481 (N_7481,N_7258,N_7283);
nand U7482 (N_7482,N_7249,N_7286);
xor U7483 (N_7483,N_7228,N_7256);
xnor U7484 (N_7484,N_7225,N_7379);
xnor U7485 (N_7485,N_7394,N_7243);
nand U7486 (N_7486,N_7290,N_7221);
nand U7487 (N_7487,N_7267,N_7296);
nand U7488 (N_7488,N_7216,N_7398);
nor U7489 (N_7489,N_7329,N_7330);
or U7490 (N_7490,N_7211,N_7383);
nand U7491 (N_7491,N_7260,N_7299);
or U7492 (N_7492,N_7310,N_7278);
nor U7493 (N_7493,N_7293,N_7344);
and U7494 (N_7494,N_7219,N_7220);
xnor U7495 (N_7495,N_7295,N_7206);
nand U7496 (N_7496,N_7361,N_7378);
nor U7497 (N_7497,N_7315,N_7298);
and U7498 (N_7498,N_7352,N_7232);
xnor U7499 (N_7499,N_7309,N_7320);
nand U7500 (N_7500,N_7227,N_7270);
nand U7501 (N_7501,N_7216,N_7359);
nor U7502 (N_7502,N_7339,N_7232);
xor U7503 (N_7503,N_7311,N_7387);
nand U7504 (N_7504,N_7210,N_7233);
xor U7505 (N_7505,N_7311,N_7378);
or U7506 (N_7506,N_7366,N_7370);
nor U7507 (N_7507,N_7201,N_7335);
xnor U7508 (N_7508,N_7380,N_7324);
or U7509 (N_7509,N_7259,N_7350);
or U7510 (N_7510,N_7205,N_7365);
nor U7511 (N_7511,N_7382,N_7205);
nor U7512 (N_7512,N_7331,N_7365);
and U7513 (N_7513,N_7300,N_7233);
and U7514 (N_7514,N_7368,N_7260);
nor U7515 (N_7515,N_7238,N_7291);
xor U7516 (N_7516,N_7393,N_7239);
nand U7517 (N_7517,N_7341,N_7248);
xor U7518 (N_7518,N_7399,N_7392);
nand U7519 (N_7519,N_7244,N_7342);
or U7520 (N_7520,N_7223,N_7220);
nand U7521 (N_7521,N_7378,N_7247);
and U7522 (N_7522,N_7322,N_7388);
and U7523 (N_7523,N_7378,N_7302);
nor U7524 (N_7524,N_7328,N_7330);
and U7525 (N_7525,N_7373,N_7234);
xor U7526 (N_7526,N_7318,N_7326);
or U7527 (N_7527,N_7394,N_7396);
or U7528 (N_7528,N_7330,N_7259);
nor U7529 (N_7529,N_7358,N_7273);
nor U7530 (N_7530,N_7376,N_7320);
nand U7531 (N_7531,N_7301,N_7266);
xnor U7532 (N_7532,N_7324,N_7214);
or U7533 (N_7533,N_7329,N_7336);
or U7534 (N_7534,N_7387,N_7399);
nor U7535 (N_7535,N_7367,N_7341);
nor U7536 (N_7536,N_7202,N_7382);
nand U7537 (N_7537,N_7310,N_7266);
nor U7538 (N_7538,N_7201,N_7234);
xor U7539 (N_7539,N_7304,N_7373);
and U7540 (N_7540,N_7305,N_7315);
xnor U7541 (N_7541,N_7291,N_7391);
nor U7542 (N_7542,N_7332,N_7292);
nor U7543 (N_7543,N_7387,N_7230);
and U7544 (N_7544,N_7336,N_7348);
xor U7545 (N_7545,N_7206,N_7223);
xor U7546 (N_7546,N_7382,N_7295);
or U7547 (N_7547,N_7228,N_7274);
or U7548 (N_7548,N_7219,N_7241);
xnor U7549 (N_7549,N_7391,N_7260);
and U7550 (N_7550,N_7272,N_7209);
nand U7551 (N_7551,N_7213,N_7325);
xnor U7552 (N_7552,N_7372,N_7300);
xor U7553 (N_7553,N_7205,N_7257);
and U7554 (N_7554,N_7321,N_7268);
or U7555 (N_7555,N_7372,N_7267);
xnor U7556 (N_7556,N_7291,N_7237);
nor U7557 (N_7557,N_7324,N_7352);
nor U7558 (N_7558,N_7222,N_7359);
nor U7559 (N_7559,N_7214,N_7359);
nand U7560 (N_7560,N_7298,N_7374);
xnor U7561 (N_7561,N_7378,N_7307);
or U7562 (N_7562,N_7334,N_7220);
nor U7563 (N_7563,N_7303,N_7345);
nand U7564 (N_7564,N_7388,N_7264);
xor U7565 (N_7565,N_7330,N_7264);
nand U7566 (N_7566,N_7398,N_7289);
or U7567 (N_7567,N_7333,N_7348);
nor U7568 (N_7568,N_7369,N_7253);
nor U7569 (N_7569,N_7258,N_7264);
and U7570 (N_7570,N_7285,N_7331);
nand U7571 (N_7571,N_7361,N_7377);
nor U7572 (N_7572,N_7330,N_7380);
xor U7573 (N_7573,N_7345,N_7223);
nand U7574 (N_7574,N_7242,N_7320);
nand U7575 (N_7575,N_7305,N_7246);
or U7576 (N_7576,N_7312,N_7289);
and U7577 (N_7577,N_7245,N_7260);
nor U7578 (N_7578,N_7301,N_7271);
or U7579 (N_7579,N_7317,N_7309);
xor U7580 (N_7580,N_7213,N_7317);
or U7581 (N_7581,N_7339,N_7384);
nand U7582 (N_7582,N_7257,N_7360);
or U7583 (N_7583,N_7391,N_7236);
and U7584 (N_7584,N_7291,N_7257);
nand U7585 (N_7585,N_7294,N_7203);
and U7586 (N_7586,N_7225,N_7357);
nand U7587 (N_7587,N_7347,N_7266);
nor U7588 (N_7588,N_7232,N_7386);
nor U7589 (N_7589,N_7332,N_7230);
nand U7590 (N_7590,N_7371,N_7232);
or U7591 (N_7591,N_7280,N_7283);
nand U7592 (N_7592,N_7393,N_7229);
or U7593 (N_7593,N_7327,N_7320);
nor U7594 (N_7594,N_7316,N_7254);
xor U7595 (N_7595,N_7391,N_7304);
or U7596 (N_7596,N_7348,N_7397);
and U7597 (N_7597,N_7254,N_7342);
nand U7598 (N_7598,N_7310,N_7320);
nor U7599 (N_7599,N_7297,N_7395);
nand U7600 (N_7600,N_7596,N_7597);
xnor U7601 (N_7601,N_7449,N_7572);
and U7602 (N_7602,N_7456,N_7508);
nand U7603 (N_7603,N_7432,N_7419);
xnor U7604 (N_7604,N_7512,N_7423);
or U7605 (N_7605,N_7599,N_7586);
nand U7606 (N_7606,N_7438,N_7588);
or U7607 (N_7607,N_7479,N_7494);
nand U7608 (N_7608,N_7568,N_7540);
nand U7609 (N_7609,N_7519,N_7448);
nand U7610 (N_7610,N_7474,N_7516);
nor U7611 (N_7611,N_7504,N_7487);
nor U7612 (N_7612,N_7463,N_7400);
nor U7613 (N_7613,N_7493,N_7515);
or U7614 (N_7614,N_7427,N_7464);
nand U7615 (N_7615,N_7591,N_7480);
nand U7616 (N_7616,N_7574,N_7551);
nand U7617 (N_7617,N_7560,N_7499);
nor U7618 (N_7618,N_7453,N_7484);
xor U7619 (N_7619,N_7531,N_7433);
nor U7620 (N_7620,N_7429,N_7570);
and U7621 (N_7621,N_7500,N_7529);
nand U7622 (N_7622,N_7444,N_7584);
nor U7623 (N_7623,N_7497,N_7535);
nand U7624 (N_7624,N_7420,N_7502);
or U7625 (N_7625,N_7442,N_7407);
nand U7626 (N_7626,N_7485,N_7593);
xnor U7627 (N_7627,N_7475,N_7486);
or U7628 (N_7628,N_7507,N_7443);
or U7629 (N_7629,N_7537,N_7575);
and U7630 (N_7630,N_7476,N_7446);
nor U7631 (N_7631,N_7452,N_7521);
xnor U7632 (N_7632,N_7518,N_7532);
or U7633 (N_7633,N_7417,N_7431);
nand U7634 (N_7634,N_7583,N_7501);
and U7635 (N_7635,N_7526,N_7592);
nor U7636 (N_7636,N_7415,N_7585);
nand U7637 (N_7637,N_7582,N_7498);
and U7638 (N_7638,N_7425,N_7589);
and U7639 (N_7639,N_7577,N_7542);
nand U7640 (N_7640,N_7559,N_7470);
and U7641 (N_7641,N_7434,N_7513);
or U7642 (N_7642,N_7450,N_7418);
or U7643 (N_7643,N_7544,N_7550);
xnor U7644 (N_7644,N_7441,N_7509);
xor U7645 (N_7645,N_7598,N_7562);
xnor U7646 (N_7646,N_7469,N_7581);
or U7647 (N_7647,N_7492,N_7565);
and U7648 (N_7648,N_7538,N_7401);
xor U7649 (N_7649,N_7579,N_7528);
xor U7650 (N_7650,N_7483,N_7455);
nor U7651 (N_7651,N_7556,N_7408);
nand U7652 (N_7652,N_7541,N_7554);
nor U7653 (N_7653,N_7534,N_7522);
and U7654 (N_7654,N_7489,N_7536);
or U7655 (N_7655,N_7472,N_7404);
nor U7656 (N_7656,N_7488,N_7495);
nand U7657 (N_7657,N_7440,N_7520);
or U7658 (N_7658,N_7558,N_7414);
nor U7659 (N_7659,N_7523,N_7465);
nand U7660 (N_7660,N_7451,N_7481);
or U7661 (N_7661,N_7552,N_7445);
nand U7662 (N_7662,N_7496,N_7530);
xnor U7663 (N_7663,N_7426,N_7439);
nor U7664 (N_7664,N_7478,N_7563);
xor U7665 (N_7665,N_7460,N_7506);
and U7666 (N_7666,N_7457,N_7406);
xnor U7667 (N_7667,N_7473,N_7459);
or U7668 (N_7668,N_7503,N_7468);
nand U7669 (N_7669,N_7573,N_7514);
xnor U7670 (N_7670,N_7436,N_7539);
nand U7671 (N_7671,N_7482,N_7403);
xor U7672 (N_7672,N_7405,N_7549);
and U7673 (N_7673,N_7547,N_7548);
nor U7674 (N_7674,N_7458,N_7412);
or U7675 (N_7675,N_7477,N_7580);
xnor U7676 (N_7676,N_7511,N_7590);
or U7677 (N_7677,N_7578,N_7525);
or U7678 (N_7678,N_7428,N_7416);
nand U7679 (N_7679,N_7510,N_7527);
and U7680 (N_7680,N_7490,N_7545);
and U7681 (N_7681,N_7447,N_7435);
and U7682 (N_7682,N_7553,N_7421);
nand U7683 (N_7683,N_7461,N_7517);
nand U7684 (N_7684,N_7561,N_7524);
xnor U7685 (N_7685,N_7569,N_7411);
xnor U7686 (N_7686,N_7454,N_7413);
and U7687 (N_7687,N_7571,N_7587);
nand U7688 (N_7688,N_7555,N_7424);
nand U7689 (N_7689,N_7402,N_7594);
and U7690 (N_7690,N_7567,N_7437);
and U7691 (N_7691,N_7546,N_7422);
and U7692 (N_7692,N_7543,N_7566);
xor U7693 (N_7693,N_7410,N_7533);
xnor U7694 (N_7694,N_7576,N_7595);
or U7695 (N_7695,N_7409,N_7430);
or U7696 (N_7696,N_7466,N_7505);
xor U7697 (N_7697,N_7564,N_7467);
nand U7698 (N_7698,N_7557,N_7491);
nand U7699 (N_7699,N_7462,N_7471);
nor U7700 (N_7700,N_7459,N_7585);
and U7701 (N_7701,N_7560,N_7583);
nor U7702 (N_7702,N_7428,N_7525);
nand U7703 (N_7703,N_7517,N_7483);
xnor U7704 (N_7704,N_7518,N_7483);
nor U7705 (N_7705,N_7545,N_7572);
xnor U7706 (N_7706,N_7422,N_7483);
or U7707 (N_7707,N_7530,N_7565);
nor U7708 (N_7708,N_7597,N_7550);
and U7709 (N_7709,N_7438,N_7565);
nand U7710 (N_7710,N_7408,N_7512);
or U7711 (N_7711,N_7442,N_7564);
and U7712 (N_7712,N_7507,N_7418);
nor U7713 (N_7713,N_7503,N_7430);
and U7714 (N_7714,N_7532,N_7599);
or U7715 (N_7715,N_7526,N_7500);
or U7716 (N_7716,N_7555,N_7505);
or U7717 (N_7717,N_7409,N_7443);
or U7718 (N_7718,N_7573,N_7428);
xor U7719 (N_7719,N_7467,N_7429);
xor U7720 (N_7720,N_7509,N_7589);
xor U7721 (N_7721,N_7476,N_7520);
nand U7722 (N_7722,N_7497,N_7517);
xor U7723 (N_7723,N_7450,N_7403);
xor U7724 (N_7724,N_7536,N_7490);
and U7725 (N_7725,N_7474,N_7457);
nor U7726 (N_7726,N_7564,N_7514);
nor U7727 (N_7727,N_7553,N_7570);
xor U7728 (N_7728,N_7506,N_7573);
xnor U7729 (N_7729,N_7441,N_7445);
xnor U7730 (N_7730,N_7569,N_7414);
nand U7731 (N_7731,N_7469,N_7472);
or U7732 (N_7732,N_7445,N_7515);
xor U7733 (N_7733,N_7578,N_7455);
or U7734 (N_7734,N_7582,N_7530);
and U7735 (N_7735,N_7408,N_7519);
and U7736 (N_7736,N_7587,N_7582);
or U7737 (N_7737,N_7533,N_7405);
or U7738 (N_7738,N_7559,N_7403);
xnor U7739 (N_7739,N_7441,N_7491);
nor U7740 (N_7740,N_7544,N_7468);
and U7741 (N_7741,N_7567,N_7574);
xnor U7742 (N_7742,N_7439,N_7553);
or U7743 (N_7743,N_7495,N_7557);
and U7744 (N_7744,N_7488,N_7562);
and U7745 (N_7745,N_7571,N_7445);
nor U7746 (N_7746,N_7583,N_7418);
nor U7747 (N_7747,N_7414,N_7575);
nand U7748 (N_7748,N_7407,N_7566);
and U7749 (N_7749,N_7568,N_7555);
xnor U7750 (N_7750,N_7470,N_7406);
nand U7751 (N_7751,N_7583,N_7598);
nand U7752 (N_7752,N_7485,N_7410);
nor U7753 (N_7753,N_7464,N_7538);
nand U7754 (N_7754,N_7464,N_7476);
xnor U7755 (N_7755,N_7593,N_7447);
and U7756 (N_7756,N_7466,N_7424);
xnor U7757 (N_7757,N_7443,N_7481);
nor U7758 (N_7758,N_7541,N_7496);
nor U7759 (N_7759,N_7412,N_7447);
xor U7760 (N_7760,N_7467,N_7584);
nand U7761 (N_7761,N_7423,N_7433);
and U7762 (N_7762,N_7513,N_7521);
nor U7763 (N_7763,N_7431,N_7460);
xor U7764 (N_7764,N_7415,N_7521);
nand U7765 (N_7765,N_7504,N_7408);
or U7766 (N_7766,N_7562,N_7469);
nand U7767 (N_7767,N_7411,N_7547);
nand U7768 (N_7768,N_7432,N_7517);
or U7769 (N_7769,N_7528,N_7490);
xor U7770 (N_7770,N_7412,N_7513);
or U7771 (N_7771,N_7419,N_7559);
and U7772 (N_7772,N_7593,N_7543);
nand U7773 (N_7773,N_7434,N_7593);
or U7774 (N_7774,N_7544,N_7450);
nand U7775 (N_7775,N_7411,N_7510);
nor U7776 (N_7776,N_7446,N_7581);
xor U7777 (N_7777,N_7496,N_7403);
nor U7778 (N_7778,N_7515,N_7426);
xor U7779 (N_7779,N_7496,N_7584);
nand U7780 (N_7780,N_7481,N_7575);
nor U7781 (N_7781,N_7571,N_7559);
nor U7782 (N_7782,N_7516,N_7484);
xor U7783 (N_7783,N_7545,N_7426);
xnor U7784 (N_7784,N_7596,N_7442);
nand U7785 (N_7785,N_7462,N_7416);
nor U7786 (N_7786,N_7520,N_7453);
or U7787 (N_7787,N_7421,N_7578);
and U7788 (N_7788,N_7550,N_7446);
and U7789 (N_7789,N_7510,N_7531);
nor U7790 (N_7790,N_7588,N_7483);
nor U7791 (N_7791,N_7400,N_7571);
nand U7792 (N_7792,N_7477,N_7487);
nand U7793 (N_7793,N_7593,N_7500);
and U7794 (N_7794,N_7513,N_7517);
and U7795 (N_7795,N_7590,N_7473);
xor U7796 (N_7796,N_7521,N_7455);
nor U7797 (N_7797,N_7443,N_7579);
or U7798 (N_7798,N_7572,N_7590);
or U7799 (N_7799,N_7520,N_7553);
or U7800 (N_7800,N_7727,N_7665);
xnor U7801 (N_7801,N_7643,N_7710);
nand U7802 (N_7802,N_7766,N_7653);
xor U7803 (N_7803,N_7627,N_7636);
nor U7804 (N_7804,N_7763,N_7645);
nor U7805 (N_7805,N_7703,N_7729);
and U7806 (N_7806,N_7635,N_7774);
xnor U7807 (N_7807,N_7679,N_7600);
nand U7808 (N_7808,N_7637,N_7617);
nor U7809 (N_7809,N_7666,N_7744);
nor U7810 (N_7810,N_7644,N_7700);
or U7811 (N_7811,N_7614,N_7756);
nor U7812 (N_7812,N_7651,N_7610);
or U7813 (N_7813,N_7683,N_7717);
xor U7814 (N_7814,N_7702,N_7648);
or U7815 (N_7815,N_7798,N_7675);
nand U7816 (N_7816,N_7603,N_7799);
and U7817 (N_7817,N_7781,N_7623);
xnor U7818 (N_7818,N_7652,N_7661);
nor U7819 (N_7819,N_7792,N_7797);
and U7820 (N_7820,N_7716,N_7794);
or U7821 (N_7821,N_7668,N_7713);
and U7822 (N_7822,N_7787,N_7671);
nand U7823 (N_7823,N_7650,N_7676);
nor U7824 (N_7824,N_7712,N_7660);
or U7825 (N_7825,N_7632,N_7677);
and U7826 (N_7826,N_7620,N_7757);
xnor U7827 (N_7827,N_7642,N_7687);
nand U7828 (N_7828,N_7732,N_7725);
or U7829 (N_7829,N_7613,N_7695);
xor U7830 (N_7830,N_7696,N_7772);
or U7831 (N_7831,N_7754,N_7667);
nor U7832 (N_7832,N_7791,N_7601);
nor U7833 (N_7833,N_7747,N_7789);
nor U7834 (N_7834,N_7780,N_7674);
nor U7835 (N_7835,N_7638,N_7705);
and U7836 (N_7836,N_7689,N_7630);
xor U7837 (N_7837,N_7608,N_7646);
xnor U7838 (N_7838,N_7796,N_7621);
or U7839 (N_7839,N_7719,N_7670);
xnor U7840 (N_7840,N_7741,N_7698);
or U7841 (N_7841,N_7678,N_7618);
and U7842 (N_7842,N_7753,N_7742);
nand U7843 (N_7843,N_7720,N_7786);
nor U7844 (N_7844,N_7692,N_7771);
nand U7845 (N_7845,N_7748,N_7723);
xor U7846 (N_7846,N_7793,N_7659);
or U7847 (N_7847,N_7656,N_7782);
xor U7848 (N_7848,N_7609,N_7778);
xor U7849 (N_7849,N_7612,N_7697);
xor U7850 (N_7850,N_7728,N_7767);
nor U7851 (N_7851,N_7706,N_7699);
nor U7852 (N_7852,N_7770,N_7761);
nor U7853 (N_7853,N_7759,N_7730);
or U7854 (N_7854,N_7615,N_7714);
nor U7855 (N_7855,N_7611,N_7625);
and U7856 (N_7856,N_7624,N_7707);
nand U7857 (N_7857,N_7775,N_7731);
or U7858 (N_7858,N_7777,N_7790);
and U7859 (N_7859,N_7693,N_7783);
or U7860 (N_7860,N_7655,N_7746);
xnor U7861 (N_7861,N_7606,N_7721);
and U7862 (N_7862,N_7694,N_7633);
nor U7863 (N_7863,N_7752,N_7773);
and U7864 (N_7864,N_7631,N_7709);
or U7865 (N_7865,N_7724,N_7669);
and U7866 (N_7866,N_7640,N_7626);
xnor U7867 (N_7867,N_7736,N_7686);
xor U7868 (N_7868,N_7764,N_7647);
or U7869 (N_7869,N_7672,N_7641);
nand U7870 (N_7870,N_7784,N_7605);
nand U7871 (N_7871,N_7688,N_7739);
xor U7872 (N_7872,N_7788,N_7735);
and U7873 (N_7873,N_7649,N_7691);
or U7874 (N_7874,N_7682,N_7726);
nand U7875 (N_7875,N_7616,N_7629);
xnor U7876 (N_7876,N_7795,N_7762);
nand U7877 (N_7877,N_7628,N_7769);
xnor U7878 (N_7878,N_7684,N_7654);
or U7879 (N_7879,N_7768,N_7663);
nor U7880 (N_7880,N_7708,N_7738);
or U7881 (N_7881,N_7607,N_7737);
xor U7882 (N_7882,N_7785,N_7779);
nand U7883 (N_7883,N_7658,N_7634);
or U7884 (N_7884,N_7681,N_7680);
nand U7885 (N_7885,N_7733,N_7751);
or U7886 (N_7886,N_7602,N_7715);
nand U7887 (N_7887,N_7758,N_7673);
nor U7888 (N_7888,N_7743,N_7776);
and U7889 (N_7889,N_7619,N_7704);
xor U7890 (N_7890,N_7760,N_7755);
or U7891 (N_7891,N_7745,N_7740);
nand U7892 (N_7892,N_7664,N_7718);
nor U7893 (N_7893,N_7750,N_7711);
xor U7894 (N_7894,N_7639,N_7734);
nand U7895 (N_7895,N_7685,N_7604);
nand U7896 (N_7896,N_7662,N_7657);
nor U7897 (N_7897,N_7765,N_7722);
nor U7898 (N_7898,N_7749,N_7690);
nor U7899 (N_7899,N_7622,N_7701);
xor U7900 (N_7900,N_7748,N_7613);
nor U7901 (N_7901,N_7729,N_7600);
nand U7902 (N_7902,N_7757,N_7740);
and U7903 (N_7903,N_7705,N_7764);
or U7904 (N_7904,N_7695,N_7766);
xnor U7905 (N_7905,N_7738,N_7785);
or U7906 (N_7906,N_7799,N_7615);
xnor U7907 (N_7907,N_7653,N_7727);
xnor U7908 (N_7908,N_7631,N_7642);
nand U7909 (N_7909,N_7640,N_7658);
xnor U7910 (N_7910,N_7662,N_7743);
or U7911 (N_7911,N_7695,N_7674);
or U7912 (N_7912,N_7649,N_7664);
nor U7913 (N_7913,N_7757,N_7718);
and U7914 (N_7914,N_7614,N_7725);
or U7915 (N_7915,N_7705,N_7628);
xnor U7916 (N_7916,N_7625,N_7630);
xor U7917 (N_7917,N_7757,N_7614);
nor U7918 (N_7918,N_7617,N_7646);
and U7919 (N_7919,N_7712,N_7749);
nor U7920 (N_7920,N_7777,N_7626);
nor U7921 (N_7921,N_7760,N_7625);
nand U7922 (N_7922,N_7677,N_7727);
nand U7923 (N_7923,N_7789,N_7692);
nand U7924 (N_7924,N_7651,N_7685);
xnor U7925 (N_7925,N_7798,N_7767);
and U7926 (N_7926,N_7774,N_7667);
or U7927 (N_7927,N_7798,N_7751);
nand U7928 (N_7928,N_7708,N_7633);
or U7929 (N_7929,N_7714,N_7703);
xnor U7930 (N_7930,N_7718,N_7770);
xor U7931 (N_7931,N_7649,N_7749);
xor U7932 (N_7932,N_7758,N_7759);
nand U7933 (N_7933,N_7715,N_7791);
nand U7934 (N_7934,N_7661,N_7679);
or U7935 (N_7935,N_7754,N_7650);
nand U7936 (N_7936,N_7606,N_7735);
nand U7937 (N_7937,N_7661,N_7745);
or U7938 (N_7938,N_7678,N_7721);
and U7939 (N_7939,N_7763,N_7711);
or U7940 (N_7940,N_7672,N_7648);
nor U7941 (N_7941,N_7650,N_7640);
xnor U7942 (N_7942,N_7780,N_7668);
or U7943 (N_7943,N_7701,N_7663);
and U7944 (N_7944,N_7691,N_7642);
or U7945 (N_7945,N_7647,N_7641);
nand U7946 (N_7946,N_7611,N_7679);
nor U7947 (N_7947,N_7744,N_7664);
or U7948 (N_7948,N_7709,N_7719);
xor U7949 (N_7949,N_7733,N_7688);
and U7950 (N_7950,N_7724,N_7663);
nor U7951 (N_7951,N_7776,N_7648);
or U7952 (N_7952,N_7725,N_7796);
nor U7953 (N_7953,N_7649,N_7665);
nor U7954 (N_7954,N_7797,N_7714);
or U7955 (N_7955,N_7673,N_7651);
and U7956 (N_7956,N_7707,N_7726);
and U7957 (N_7957,N_7760,N_7646);
and U7958 (N_7958,N_7654,N_7664);
xnor U7959 (N_7959,N_7661,N_7626);
or U7960 (N_7960,N_7643,N_7759);
nand U7961 (N_7961,N_7726,N_7674);
nand U7962 (N_7962,N_7764,N_7635);
or U7963 (N_7963,N_7791,N_7793);
nor U7964 (N_7964,N_7685,N_7775);
or U7965 (N_7965,N_7604,N_7719);
nand U7966 (N_7966,N_7748,N_7773);
and U7967 (N_7967,N_7767,N_7740);
nor U7968 (N_7968,N_7722,N_7694);
nand U7969 (N_7969,N_7674,N_7753);
nand U7970 (N_7970,N_7789,N_7761);
nand U7971 (N_7971,N_7690,N_7773);
xnor U7972 (N_7972,N_7609,N_7704);
nor U7973 (N_7973,N_7724,N_7751);
xor U7974 (N_7974,N_7670,N_7674);
nor U7975 (N_7975,N_7637,N_7724);
nor U7976 (N_7976,N_7778,N_7733);
and U7977 (N_7977,N_7680,N_7676);
nor U7978 (N_7978,N_7674,N_7718);
nand U7979 (N_7979,N_7658,N_7626);
nand U7980 (N_7980,N_7719,N_7722);
nand U7981 (N_7981,N_7616,N_7601);
nor U7982 (N_7982,N_7720,N_7701);
and U7983 (N_7983,N_7607,N_7630);
and U7984 (N_7984,N_7792,N_7755);
nand U7985 (N_7985,N_7741,N_7648);
nor U7986 (N_7986,N_7629,N_7650);
nor U7987 (N_7987,N_7709,N_7661);
nand U7988 (N_7988,N_7785,N_7664);
xor U7989 (N_7989,N_7681,N_7778);
and U7990 (N_7990,N_7699,N_7700);
and U7991 (N_7991,N_7771,N_7610);
nor U7992 (N_7992,N_7751,N_7767);
or U7993 (N_7993,N_7709,N_7619);
or U7994 (N_7994,N_7698,N_7690);
nor U7995 (N_7995,N_7633,N_7641);
nand U7996 (N_7996,N_7756,N_7701);
and U7997 (N_7997,N_7754,N_7797);
nor U7998 (N_7998,N_7652,N_7646);
and U7999 (N_7999,N_7744,N_7730);
or U8000 (N_8000,N_7857,N_7963);
or U8001 (N_8001,N_7868,N_7951);
nand U8002 (N_8002,N_7960,N_7879);
nor U8003 (N_8003,N_7920,N_7804);
xnor U8004 (N_8004,N_7891,N_7840);
and U8005 (N_8005,N_7852,N_7832);
nor U8006 (N_8006,N_7926,N_7897);
nor U8007 (N_8007,N_7914,N_7904);
nor U8008 (N_8008,N_7883,N_7933);
xor U8009 (N_8009,N_7999,N_7885);
and U8010 (N_8010,N_7950,N_7820);
nor U8011 (N_8011,N_7859,N_7866);
nand U8012 (N_8012,N_7872,N_7818);
nand U8013 (N_8013,N_7887,N_7845);
and U8014 (N_8014,N_7819,N_7966);
nor U8015 (N_8015,N_7865,N_7830);
or U8016 (N_8016,N_7978,N_7844);
xor U8017 (N_8017,N_7921,N_7870);
nor U8018 (N_8018,N_7903,N_7803);
xor U8019 (N_8019,N_7871,N_7889);
nand U8020 (N_8020,N_7959,N_7900);
nand U8021 (N_8021,N_7888,N_7860);
xnor U8022 (N_8022,N_7997,N_7980);
and U8023 (N_8023,N_7800,N_7975);
nor U8024 (N_8024,N_7996,N_7829);
and U8025 (N_8025,N_7919,N_7934);
nor U8026 (N_8026,N_7922,N_7983);
nor U8027 (N_8027,N_7902,N_7946);
nor U8028 (N_8028,N_7935,N_7906);
or U8029 (N_8029,N_7989,N_7952);
nor U8030 (N_8030,N_7878,N_7849);
xnor U8031 (N_8031,N_7956,N_7968);
or U8032 (N_8032,N_7850,N_7886);
xor U8033 (N_8033,N_7974,N_7815);
nand U8034 (N_8034,N_7985,N_7958);
or U8035 (N_8035,N_7896,N_7979);
or U8036 (N_8036,N_7984,N_7831);
and U8037 (N_8037,N_7947,N_7907);
and U8038 (N_8038,N_7917,N_7801);
or U8039 (N_8039,N_7977,N_7987);
nor U8040 (N_8040,N_7937,N_7862);
nor U8041 (N_8041,N_7908,N_7940);
nand U8042 (N_8042,N_7967,N_7816);
nor U8043 (N_8043,N_7884,N_7838);
nand U8044 (N_8044,N_7976,N_7942);
xnor U8045 (N_8045,N_7825,N_7846);
and U8046 (N_8046,N_7964,N_7855);
nand U8047 (N_8047,N_7988,N_7808);
xnor U8048 (N_8048,N_7882,N_7923);
xnor U8049 (N_8049,N_7824,N_7913);
or U8050 (N_8050,N_7995,N_7848);
or U8051 (N_8051,N_7867,N_7991);
or U8052 (N_8052,N_7854,N_7938);
nor U8053 (N_8053,N_7861,N_7961);
or U8054 (N_8054,N_7955,N_7881);
xnor U8055 (N_8055,N_7924,N_7828);
nand U8056 (N_8056,N_7813,N_7895);
nand U8057 (N_8057,N_7842,N_7847);
nor U8058 (N_8058,N_7949,N_7863);
nand U8059 (N_8059,N_7982,N_7993);
xnor U8060 (N_8060,N_7998,N_7918);
xor U8061 (N_8061,N_7970,N_7823);
nand U8062 (N_8062,N_7817,N_7931);
or U8063 (N_8063,N_7927,N_7841);
and U8064 (N_8064,N_7853,N_7809);
xor U8065 (N_8065,N_7802,N_7930);
xnor U8066 (N_8066,N_7890,N_7836);
nor U8067 (N_8067,N_7972,N_7901);
or U8068 (N_8068,N_7894,N_7953);
nand U8069 (N_8069,N_7892,N_7945);
and U8070 (N_8070,N_7954,N_7874);
nor U8071 (N_8071,N_7909,N_7864);
nor U8072 (N_8072,N_7899,N_7827);
nor U8073 (N_8073,N_7925,N_7876);
xnor U8074 (N_8074,N_7806,N_7869);
and U8075 (N_8075,N_7835,N_7932);
nand U8076 (N_8076,N_7948,N_7973);
or U8077 (N_8077,N_7856,N_7994);
nand U8078 (N_8078,N_7969,N_7928);
nand U8079 (N_8079,N_7837,N_7851);
nor U8080 (N_8080,N_7877,N_7971);
nand U8081 (N_8081,N_7941,N_7939);
nor U8082 (N_8082,N_7986,N_7910);
nand U8083 (N_8083,N_7944,N_7929);
or U8084 (N_8084,N_7821,N_7834);
nand U8085 (N_8085,N_7905,N_7875);
nor U8086 (N_8086,N_7990,N_7880);
nor U8087 (N_8087,N_7981,N_7911);
nand U8088 (N_8088,N_7943,N_7957);
xnor U8089 (N_8089,N_7936,N_7812);
nand U8090 (N_8090,N_7805,N_7807);
nand U8091 (N_8091,N_7912,N_7858);
nand U8092 (N_8092,N_7814,N_7898);
and U8093 (N_8093,N_7962,N_7833);
and U8094 (N_8094,N_7811,N_7843);
nand U8095 (N_8095,N_7839,N_7965);
xor U8096 (N_8096,N_7873,N_7826);
and U8097 (N_8097,N_7810,N_7992);
nand U8098 (N_8098,N_7915,N_7822);
nand U8099 (N_8099,N_7893,N_7916);
or U8100 (N_8100,N_7843,N_7948);
xnor U8101 (N_8101,N_7973,N_7800);
and U8102 (N_8102,N_7833,N_7954);
xnor U8103 (N_8103,N_7913,N_7904);
nand U8104 (N_8104,N_7968,N_7834);
and U8105 (N_8105,N_7851,N_7939);
xnor U8106 (N_8106,N_7844,N_7879);
nand U8107 (N_8107,N_7850,N_7937);
nand U8108 (N_8108,N_7997,N_7855);
or U8109 (N_8109,N_7860,N_7806);
nor U8110 (N_8110,N_7932,N_7999);
xor U8111 (N_8111,N_7959,N_7906);
xnor U8112 (N_8112,N_7802,N_7952);
nor U8113 (N_8113,N_7996,N_7867);
nor U8114 (N_8114,N_7850,N_7992);
xnor U8115 (N_8115,N_7969,N_7949);
nand U8116 (N_8116,N_7880,N_7835);
and U8117 (N_8117,N_7848,N_7853);
nor U8118 (N_8118,N_7879,N_7855);
nor U8119 (N_8119,N_7923,N_7892);
or U8120 (N_8120,N_7971,N_7976);
nor U8121 (N_8121,N_7927,N_7944);
nand U8122 (N_8122,N_7837,N_7981);
nor U8123 (N_8123,N_7935,N_7808);
nand U8124 (N_8124,N_7936,N_7825);
or U8125 (N_8125,N_7903,N_7892);
and U8126 (N_8126,N_7931,N_7810);
xor U8127 (N_8127,N_7908,N_7802);
nand U8128 (N_8128,N_7831,N_7899);
and U8129 (N_8129,N_7920,N_7895);
and U8130 (N_8130,N_7830,N_7892);
nand U8131 (N_8131,N_7894,N_7914);
or U8132 (N_8132,N_7976,N_7983);
or U8133 (N_8133,N_7957,N_7876);
nand U8134 (N_8134,N_7986,N_7991);
and U8135 (N_8135,N_7817,N_7964);
and U8136 (N_8136,N_7903,N_7865);
nand U8137 (N_8137,N_7981,N_7810);
nand U8138 (N_8138,N_7993,N_7979);
and U8139 (N_8139,N_7868,N_7834);
and U8140 (N_8140,N_7927,N_7800);
or U8141 (N_8141,N_7922,N_7905);
or U8142 (N_8142,N_7980,N_7829);
and U8143 (N_8143,N_7972,N_7906);
and U8144 (N_8144,N_7831,N_7890);
xor U8145 (N_8145,N_7803,N_7812);
nor U8146 (N_8146,N_7893,N_7867);
nor U8147 (N_8147,N_7994,N_7997);
nand U8148 (N_8148,N_7855,N_7888);
xor U8149 (N_8149,N_7965,N_7843);
and U8150 (N_8150,N_7858,N_7964);
nor U8151 (N_8151,N_7916,N_7818);
or U8152 (N_8152,N_7878,N_7928);
nand U8153 (N_8153,N_7857,N_7914);
or U8154 (N_8154,N_7965,N_7804);
nor U8155 (N_8155,N_7974,N_7926);
nand U8156 (N_8156,N_7912,N_7837);
or U8157 (N_8157,N_7965,N_7847);
xnor U8158 (N_8158,N_7880,N_7967);
or U8159 (N_8159,N_7958,N_7828);
or U8160 (N_8160,N_7889,N_7917);
and U8161 (N_8161,N_7960,N_7891);
nor U8162 (N_8162,N_7990,N_7908);
or U8163 (N_8163,N_7931,N_7813);
nand U8164 (N_8164,N_7926,N_7887);
nor U8165 (N_8165,N_7839,N_7967);
nor U8166 (N_8166,N_7852,N_7870);
or U8167 (N_8167,N_7948,N_7815);
or U8168 (N_8168,N_7977,N_7877);
nand U8169 (N_8169,N_7939,N_7887);
and U8170 (N_8170,N_7989,N_7860);
or U8171 (N_8171,N_7833,N_7938);
and U8172 (N_8172,N_7807,N_7976);
and U8173 (N_8173,N_7906,N_7884);
and U8174 (N_8174,N_7871,N_7972);
nand U8175 (N_8175,N_7865,N_7985);
xor U8176 (N_8176,N_7828,N_7954);
or U8177 (N_8177,N_7977,N_7954);
nor U8178 (N_8178,N_7848,N_7824);
and U8179 (N_8179,N_7955,N_7860);
and U8180 (N_8180,N_7879,N_7942);
and U8181 (N_8181,N_7881,N_7976);
nor U8182 (N_8182,N_7841,N_7880);
nand U8183 (N_8183,N_7985,N_7878);
and U8184 (N_8184,N_7857,N_7844);
nand U8185 (N_8185,N_7988,N_7904);
nand U8186 (N_8186,N_7960,N_7874);
nand U8187 (N_8187,N_7919,N_7889);
and U8188 (N_8188,N_7885,N_7984);
nand U8189 (N_8189,N_7819,N_7967);
nor U8190 (N_8190,N_7883,N_7871);
xnor U8191 (N_8191,N_7867,N_7843);
or U8192 (N_8192,N_7882,N_7960);
nand U8193 (N_8193,N_7994,N_7989);
xor U8194 (N_8194,N_7907,N_7970);
xnor U8195 (N_8195,N_7828,N_7827);
nor U8196 (N_8196,N_7826,N_7893);
xor U8197 (N_8197,N_7911,N_7970);
xnor U8198 (N_8198,N_7873,N_7897);
nand U8199 (N_8199,N_7955,N_7832);
and U8200 (N_8200,N_8109,N_8065);
nor U8201 (N_8201,N_8030,N_8027);
or U8202 (N_8202,N_8114,N_8147);
xor U8203 (N_8203,N_8080,N_8063);
xnor U8204 (N_8204,N_8172,N_8037);
nor U8205 (N_8205,N_8005,N_8074);
or U8206 (N_8206,N_8150,N_8036);
nand U8207 (N_8207,N_8157,N_8155);
nor U8208 (N_8208,N_8044,N_8011);
xnor U8209 (N_8209,N_8035,N_8085);
nand U8210 (N_8210,N_8170,N_8015);
nand U8211 (N_8211,N_8033,N_8175);
xor U8212 (N_8212,N_8024,N_8107);
nand U8213 (N_8213,N_8019,N_8018);
xor U8214 (N_8214,N_8093,N_8095);
nor U8215 (N_8215,N_8016,N_8143);
or U8216 (N_8216,N_8053,N_8077);
or U8217 (N_8217,N_8195,N_8094);
and U8218 (N_8218,N_8086,N_8025);
xnor U8219 (N_8219,N_8180,N_8088);
nor U8220 (N_8220,N_8000,N_8101);
and U8221 (N_8221,N_8191,N_8042);
nor U8222 (N_8222,N_8091,N_8148);
nand U8223 (N_8223,N_8159,N_8022);
and U8224 (N_8224,N_8081,N_8198);
and U8225 (N_8225,N_8097,N_8104);
nor U8226 (N_8226,N_8039,N_8123);
xor U8227 (N_8227,N_8064,N_8145);
nand U8228 (N_8228,N_8013,N_8179);
nor U8229 (N_8229,N_8135,N_8003);
and U8230 (N_8230,N_8099,N_8133);
xnor U8231 (N_8231,N_8059,N_8112);
xor U8232 (N_8232,N_8158,N_8105);
xnor U8233 (N_8233,N_8152,N_8009);
nand U8234 (N_8234,N_8188,N_8066);
xnor U8235 (N_8235,N_8174,N_8178);
xor U8236 (N_8236,N_8144,N_8041);
and U8237 (N_8237,N_8128,N_8162);
xnor U8238 (N_8238,N_8167,N_8173);
nor U8239 (N_8239,N_8050,N_8168);
or U8240 (N_8240,N_8196,N_8048);
nor U8241 (N_8241,N_8113,N_8043);
nor U8242 (N_8242,N_8089,N_8138);
nor U8243 (N_8243,N_8082,N_8060);
or U8244 (N_8244,N_8054,N_8171);
or U8245 (N_8245,N_8186,N_8069);
or U8246 (N_8246,N_8079,N_8008);
or U8247 (N_8247,N_8068,N_8028);
nor U8248 (N_8248,N_8115,N_8141);
nand U8249 (N_8249,N_8119,N_8103);
or U8250 (N_8250,N_8197,N_8110);
and U8251 (N_8251,N_8100,N_8061);
nand U8252 (N_8252,N_8012,N_8132);
nor U8253 (N_8253,N_8125,N_8070);
nor U8254 (N_8254,N_8160,N_8038);
nand U8255 (N_8255,N_8182,N_8111);
nor U8256 (N_8256,N_8078,N_8031);
xnor U8257 (N_8257,N_8121,N_8154);
or U8258 (N_8258,N_8029,N_8140);
or U8259 (N_8259,N_8098,N_8149);
nor U8260 (N_8260,N_8151,N_8006);
xnor U8261 (N_8261,N_8153,N_8164);
nor U8262 (N_8262,N_8139,N_8076);
xor U8263 (N_8263,N_8004,N_8049);
xor U8264 (N_8264,N_8120,N_8166);
and U8265 (N_8265,N_8047,N_8106);
nor U8266 (N_8266,N_8165,N_8137);
or U8267 (N_8267,N_8046,N_8014);
nand U8268 (N_8268,N_8199,N_8102);
or U8269 (N_8269,N_8010,N_8072);
and U8270 (N_8270,N_8073,N_8183);
nor U8271 (N_8271,N_8087,N_8002);
and U8272 (N_8272,N_8116,N_8083);
and U8273 (N_8273,N_8055,N_8096);
or U8274 (N_8274,N_8026,N_8134);
and U8275 (N_8275,N_8130,N_8194);
or U8276 (N_8276,N_8127,N_8146);
and U8277 (N_8277,N_8161,N_8007);
nand U8278 (N_8278,N_8193,N_8021);
nor U8279 (N_8279,N_8040,N_8034);
xnor U8280 (N_8280,N_8001,N_8058);
nor U8281 (N_8281,N_8032,N_8187);
nand U8282 (N_8282,N_8108,N_8189);
nand U8283 (N_8283,N_8084,N_8090);
xor U8284 (N_8284,N_8136,N_8163);
nand U8285 (N_8285,N_8045,N_8156);
nor U8286 (N_8286,N_8071,N_8122);
xor U8287 (N_8287,N_8056,N_8131);
nand U8288 (N_8288,N_8169,N_8075);
nand U8289 (N_8289,N_8142,N_8184);
nand U8290 (N_8290,N_8017,N_8176);
nand U8291 (N_8291,N_8062,N_8057);
or U8292 (N_8292,N_8067,N_8192);
or U8293 (N_8293,N_8129,N_8020);
and U8294 (N_8294,N_8092,N_8052);
nor U8295 (N_8295,N_8126,N_8177);
nand U8296 (N_8296,N_8181,N_8118);
and U8297 (N_8297,N_8190,N_8124);
nor U8298 (N_8298,N_8185,N_8023);
xnor U8299 (N_8299,N_8051,N_8117);
nor U8300 (N_8300,N_8167,N_8146);
or U8301 (N_8301,N_8038,N_8018);
xor U8302 (N_8302,N_8017,N_8086);
and U8303 (N_8303,N_8001,N_8127);
xor U8304 (N_8304,N_8179,N_8169);
or U8305 (N_8305,N_8045,N_8019);
or U8306 (N_8306,N_8110,N_8033);
and U8307 (N_8307,N_8193,N_8067);
xnor U8308 (N_8308,N_8020,N_8004);
nor U8309 (N_8309,N_8078,N_8130);
nor U8310 (N_8310,N_8124,N_8127);
and U8311 (N_8311,N_8111,N_8046);
or U8312 (N_8312,N_8157,N_8105);
and U8313 (N_8313,N_8119,N_8172);
nor U8314 (N_8314,N_8104,N_8011);
xnor U8315 (N_8315,N_8059,N_8019);
nor U8316 (N_8316,N_8000,N_8085);
xnor U8317 (N_8317,N_8054,N_8155);
nor U8318 (N_8318,N_8072,N_8006);
nand U8319 (N_8319,N_8063,N_8091);
xor U8320 (N_8320,N_8021,N_8174);
nand U8321 (N_8321,N_8172,N_8020);
nand U8322 (N_8322,N_8003,N_8104);
nand U8323 (N_8323,N_8143,N_8129);
nor U8324 (N_8324,N_8006,N_8149);
nor U8325 (N_8325,N_8135,N_8060);
xor U8326 (N_8326,N_8179,N_8047);
or U8327 (N_8327,N_8015,N_8091);
xor U8328 (N_8328,N_8083,N_8149);
or U8329 (N_8329,N_8193,N_8042);
nor U8330 (N_8330,N_8182,N_8147);
and U8331 (N_8331,N_8049,N_8031);
and U8332 (N_8332,N_8012,N_8078);
nor U8333 (N_8333,N_8049,N_8150);
and U8334 (N_8334,N_8065,N_8070);
nor U8335 (N_8335,N_8106,N_8161);
or U8336 (N_8336,N_8114,N_8075);
xnor U8337 (N_8337,N_8050,N_8091);
or U8338 (N_8338,N_8072,N_8166);
nand U8339 (N_8339,N_8158,N_8052);
nor U8340 (N_8340,N_8088,N_8060);
xor U8341 (N_8341,N_8149,N_8089);
nand U8342 (N_8342,N_8080,N_8139);
or U8343 (N_8343,N_8185,N_8198);
or U8344 (N_8344,N_8134,N_8097);
or U8345 (N_8345,N_8036,N_8116);
and U8346 (N_8346,N_8137,N_8163);
and U8347 (N_8347,N_8081,N_8150);
nand U8348 (N_8348,N_8080,N_8126);
xor U8349 (N_8349,N_8094,N_8099);
nand U8350 (N_8350,N_8142,N_8038);
nor U8351 (N_8351,N_8180,N_8022);
nand U8352 (N_8352,N_8174,N_8049);
nor U8353 (N_8353,N_8078,N_8039);
and U8354 (N_8354,N_8141,N_8018);
and U8355 (N_8355,N_8064,N_8033);
nand U8356 (N_8356,N_8198,N_8103);
nand U8357 (N_8357,N_8079,N_8134);
or U8358 (N_8358,N_8137,N_8036);
nand U8359 (N_8359,N_8044,N_8145);
xnor U8360 (N_8360,N_8007,N_8082);
xor U8361 (N_8361,N_8159,N_8132);
xor U8362 (N_8362,N_8096,N_8060);
xnor U8363 (N_8363,N_8034,N_8168);
or U8364 (N_8364,N_8010,N_8060);
xnor U8365 (N_8365,N_8194,N_8054);
or U8366 (N_8366,N_8021,N_8046);
nand U8367 (N_8367,N_8122,N_8043);
xor U8368 (N_8368,N_8146,N_8138);
xor U8369 (N_8369,N_8170,N_8109);
and U8370 (N_8370,N_8142,N_8174);
nor U8371 (N_8371,N_8046,N_8117);
or U8372 (N_8372,N_8163,N_8046);
or U8373 (N_8373,N_8036,N_8109);
and U8374 (N_8374,N_8168,N_8171);
and U8375 (N_8375,N_8169,N_8160);
and U8376 (N_8376,N_8025,N_8035);
nor U8377 (N_8377,N_8196,N_8110);
nand U8378 (N_8378,N_8188,N_8115);
xnor U8379 (N_8379,N_8040,N_8068);
and U8380 (N_8380,N_8150,N_8008);
xor U8381 (N_8381,N_8070,N_8003);
or U8382 (N_8382,N_8016,N_8028);
xor U8383 (N_8383,N_8168,N_8162);
xnor U8384 (N_8384,N_8142,N_8154);
xnor U8385 (N_8385,N_8117,N_8006);
nand U8386 (N_8386,N_8065,N_8177);
or U8387 (N_8387,N_8142,N_8014);
nor U8388 (N_8388,N_8151,N_8057);
and U8389 (N_8389,N_8052,N_8023);
or U8390 (N_8390,N_8012,N_8085);
nor U8391 (N_8391,N_8086,N_8010);
xnor U8392 (N_8392,N_8093,N_8022);
or U8393 (N_8393,N_8104,N_8017);
xor U8394 (N_8394,N_8007,N_8020);
nor U8395 (N_8395,N_8095,N_8019);
or U8396 (N_8396,N_8102,N_8058);
and U8397 (N_8397,N_8088,N_8195);
nor U8398 (N_8398,N_8095,N_8111);
or U8399 (N_8399,N_8123,N_8067);
nand U8400 (N_8400,N_8292,N_8352);
xor U8401 (N_8401,N_8217,N_8357);
nand U8402 (N_8402,N_8371,N_8314);
and U8403 (N_8403,N_8315,N_8216);
nand U8404 (N_8404,N_8267,N_8387);
or U8405 (N_8405,N_8329,N_8251);
nand U8406 (N_8406,N_8369,N_8305);
nand U8407 (N_8407,N_8373,N_8259);
nor U8408 (N_8408,N_8330,N_8236);
or U8409 (N_8409,N_8263,N_8232);
nor U8410 (N_8410,N_8248,N_8244);
and U8411 (N_8411,N_8380,N_8331);
nand U8412 (N_8412,N_8328,N_8346);
nand U8413 (N_8413,N_8228,N_8250);
nand U8414 (N_8414,N_8212,N_8210);
and U8415 (N_8415,N_8301,N_8200);
nand U8416 (N_8416,N_8358,N_8270);
or U8417 (N_8417,N_8208,N_8264);
xor U8418 (N_8418,N_8275,N_8254);
and U8419 (N_8419,N_8283,N_8229);
nand U8420 (N_8420,N_8304,N_8245);
and U8421 (N_8421,N_8324,N_8391);
nor U8422 (N_8422,N_8388,N_8211);
nand U8423 (N_8423,N_8285,N_8295);
nand U8424 (N_8424,N_8379,N_8221);
nand U8425 (N_8425,N_8351,N_8306);
and U8426 (N_8426,N_8332,N_8239);
xor U8427 (N_8427,N_8226,N_8280);
nand U8428 (N_8428,N_8303,N_8320);
nand U8429 (N_8429,N_8213,N_8318);
and U8430 (N_8430,N_8282,N_8337);
or U8431 (N_8431,N_8365,N_8386);
and U8432 (N_8432,N_8345,N_8340);
nor U8433 (N_8433,N_8218,N_8268);
nor U8434 (N_8434,N_8246,N_8383);
nand U8435 (N_8435,N_8374,N_8396);
and U8436 (N_8436,N_8397,N_8399);
nand U8437 (N_8437,N_8209,N_8363);
xor U8438 (N_8438,N_8235,N_8203);
xor U8439 (N_8439,N_8290,N_8398);
nand U8440 (N_8440,N_8389,N_8243);
and U8441 (N_8441,N_8240,N_8261);
xor U8442 (N_8442,N_8287,N_8273);
nand U8443 (N_8443,N_8323,N_8327);
or U8444 (N_8444,N_8269,N_8255);
xnor U8445 (N_8445,N_8336,N_8207);
or U8446 (N_8446,N_8238,N_8308);
nor U8447 (N_8447,N_8321,N_8370);
and U8448 (N_8448,N_8341,N_8220);
nor U8449 (N_8449,N_8353,N_8249);
or U8450 (N_8450,N_8338,N_8241);
nor U8451 (N_8451,N_8281,N_8237);
or U8452 (N_8452,N_8349,N_8310);
nand U8453 (N_8453,N_8348,N_8205);
xor U8454 (N_8454,N_8376,N_8347);
and U8455 (N_8455,N_8364,N_8278);
xnor U8456 (N_8456,N_8289,N_8350);
nor U8457 (N_8457,N_8252,N_8272);
nor U8458 (N_8458,N_8260,N_8333);
and U8459 (N_8459,N_8395,N_8367);
nand U8460 (N_8460,N_8311,N_8277);
and U8461 (N_8461,N_8284,N_8247);
and U8462 (N_8462,N_8319,N_8293);
or U8463 (N_8463,N_8355,N_8392);
xor U8464 (N_8464,N_8325,N_8382);
xnor U8465 (N_8465,N_8368,N_8356);
or U8466 (N_8466,N_8343,N_8265);
xor U8467 (N_8467,N_8257,N_8242);
nand U8468 (N_8468,N_8344,N_8322);
and U8469 (N_8469,N_8309,N_8334);
xor U8470 (N_8470,N_8354,N_8366);
nand U8471 (N_8471,N_8223,N_8393);
or U8472 (N_8472,N_8359,N_8222);
xor U8473 (N_8473,N_8276,N_8316);
or U8474 (N_8474,N_8291,N_8230);
xor U8475 (N_8475,N_8384,N_8219);
and U8476 (N_8476,N_8271,N_8215);
nand U8477 (N_8477,N_8201,N_8375);
xnor U8478 (N_8478,N_8224,N_8326);
and U8479 (N_8479,N_8307,N_8253);
nor U8480 (N_8480,N_8225,N_8378);
nor U8481 (N_8481,N_8298,N_8342);
nor U8482 (N_8482,N_8361,N_8227);
and U8483 (N_8483,N_8296,N_8313);
xnor U8484 (N_8484,N_8234,N_8299);
xnor U8485 (N_8485,N_8274,N_8372);
nand U8486 (N_8486,N_8233,N_8231);
nor U8487 (N_8487,N_8288,N_8266);
nor U8488 (N_8488,N_8394,N_8377);
xor U8489 (N_8489,N_8302,N_8390);
nand U8490 (N_8490,N_8258,N_8312);
nand U8491 (N_8491,N_8214,N_8317);
xor U8492 (N_8492,N_8286,N_8206);
xor U8493 (N_8493,N_8294,N_8279);
nand U8494 (N_8494,N_8360,N_8297);
nor U8495 (N_8495,N_8202,N_8385);
and U8496 (N_8496,N_8335,N_8300);
nand U8497 (N_8497,N_8262,N_8339);
xor U8498 (N_8498,N_8362,N_8381);
and U8499 (N_8499,N_8256,N_8204);
nor U8500 (N_8500,N_8209,N_8257);
and U8501 (N_8501,N_8365,N_8326);
or U8502 (N_8502,N_8252,N_8338);
nor U8503 (N_8503,N_8221,N_8290);
xnor U8504 (N_8504,N_8350,N_8303);
or U8505 (N_8505,N_8288,N_8291);
xor U8506 (N_8506,N_8353,N_8271);
or U8507 (N_8507,N_8315,N_8217);
xnor U8508 (N_8508,N_8394,N_8261);
or U8509 (N_8509,N_8280,N_8284);
nand U8510 (N_8510,N_8291,N_8287);
nor U8511 (N_8511,N_8386,N_8247);
and U8512 (N_8512,N_8245,N_8223);
xor U8513 (N_8513,N_8257,N_8376);
nor U8514 (N_8514,N_8307,N_8353);
or U8515 (N_8515,N_8385,N_8296);
xor U8516 (N_8516,N_8354,N_8253);
and U8517 (N_8517,N_8254,N_8287);
or U8518 (N_8518,N_8369,N_8253);
or U8519 (N_8519,N_8337,N_8341);
nor U8520 (N_8520,N_8386,N_8244);
nand U8521 (N_8521,N_8206,N_8278);
nor U8522 (N_8522,N_8376,N_8259);
xnor U8523 (N_8523,N_8346,N_8248);
nor U8524 (N_8524,N_8394,N_8251);
and U8525 (N_8525,N_8284,N_8273);
xnor U8526 (N_8526,N_8245,N_8318);
nor U8527 (N_8527,N_8346,N_8339);
nor U8528 (N_8528,N_8208,N_8365);
nand U8529 (N_8529,N_8267,N_8203);
and U8530 (N_8530,N_8315,N_8229);
or U8531 (N_8531,N_8273,N_8279);
nand U8532 (N_8532,N_8386,N_8396);
nand U8533 (N_8533,N_8372,N_8342);
xor U8534 (N_8534,N_8303,N_8271);
nor U8535 (N_8535,N_8301,N_8220);
or U8536 (N_8536,N_8370,N_8378);
xnor U8537 (N_8537,N_8349,N_8290);
nor U8538 (N_8538,N_8367,N_8240);
and U8539 (N_8539,N_8223,N_8211);
nand U8540 (N_8540,N_8391,N_8328);
or U8541 (N_8541,N_8211,N_8382);
or U8542 (N_8542,N_8267,N_8269);
nand U8543 (N_8543,N_8254,N_8389);
nor U8544 (N_8544,N_8353,N_8344);
or U8545 (N_8545,N_8207,N_8287);
or U8546 (N_8546,N_8265,N_8311);
nor U8547 (N_8547,N_8324,N_8245);
or U8548 (N_8548,N_8340,N_8296);
nor U8549 (N_8549,N_8377,N_8239);
xor U8550 (N_8550,N_8238,N_8286);
nor U8551 (N_8551,N_8366,N_8275);
xor U8552 (N_8552,N_8306,N_8204);
nor U8553 (N_8553,N_8365,N_8237);
xor U8554 (N_8554,N_8355,N_8211);
and U8555 (N_8555,N_8207,N_8272);
or U8556 (N_8556,N_8215,N_8242);
nor U8557 (N_8557,N_8278,N_8318);
or U8558 (N_8558,N_8209,N_8272);
nor U8559 (N_8559,N_8309,N_8366);
nor U8560 (N_8560,N_8294,N_8323);
xor U8561 (N_8561,N_8203,N_8260);
or U8562 (N_8562,N_8237,N_8355);
nand U8563 (N_8563,N_8367,N_8220);
xor U8564 (N_8564,N_8342,N_8253);
nor U8565 (N_8565,N_8345,N_8311);
nand U8566 (N_8566,N_8257,N_8352);
nand U8567 (N_8567,N_8276,N_8397);
or U8568 (N_8568,N_8321,N_8384);
nand U8569 (N_8569,N_8285,N_8219);
nor U8570 (N_8570,N_8349,N_8329);
or U8571 (N_8571,N_8355,N_8315);
and U8572 (N_8572,N_8395,N_8296);
xor U8573 (N_8573,N_8293,N_8349);
nor U8574 (N_8574,N_8353,N_8228);
nor U8575 (N_8575,N_8354,N_8320);
and U8576 (N_8576,N_8323,N_8382);
and U8577 (N_8577,N_8208,N_8256);
and U8578 (N_8578,N_8375,N_8322);
and U8579 (N_8579,N_8388,N_8337);
nand U8580 (N_8580,N_8260,N_8234);
nand U8581 (N_8581,N_8273,N_8256);
nand U8582 (N_8582,N_8203,N_8353);
xor U8583 (N_8583,N_8372,N_8325);
and U8584 (N_8584,N_8229,N_8201);
xnor U8585 (N_8585,N_8327,N_8366);
nor U8586 (N_8586,N_8351,N_8336);
xor U8587 (N_8587,N_8320,N_8367);
xnor U8588 (N_8588,N_8391,N_8308);
xor U8589 (N_8589,N_8305,N_8300);
nor U8590 (N_8590,N_8344,N_8201);
and U8591 (N_8591,N_8381,N_8375);
nor U8592 (N_8592,N_8349,N_8227);
nand U8593 (N_8593,N_8280,N_8332);
xnor U8594 (N_8594,N_8346,N_8299);
or U8595 (N_8595,N_8283,N_8203);
or U8596 (N_8596,N_8333,N_8284);
or U8597 (N_8597,N_8322,N_8279);
nor U8598 (N_8598,N_8295,N_8231);
nor U8599 (N_8599,N_8211,N_8256);
xor U8600 (N_8600,N_8578,N_8498);
or U8601 (N_8601,N_8490,N_8564);
nand U8602 (N_8602,N_8444,N_8484);
or U8603 (N_8603,N_8571,N_8581);
xor U8604 (N_8604,N_8559,N_8537);
and U8605 (N_8605,N_8493,N_8523);
nand U8606 (N_8606,N_8451,N_8545);
nor U8607 (N_8607,N_8516,N_8476);
nor U8608 (N_8608,N_8457,N_8435);
or U8609 (N_8609,N_8464,N_8495);
xor U8610 (N_8610,N_8550,N_8400);
nor U8611 (N_8611,N_8416,N_8541);
nand U8612 (N_8612,N_8404,N_8549);
xor U8613 (N_8613,N_8483,N_8417);
and U8614 (N_8614,N_8494,N_8441);
and U8615 (N_8615,N_8401,N_8474);
nor U8616 (N_8616,N_8514,N_8518);
nor U8617 (N_8617,N_8566,N_8431);
nor U8618 (N_8618,N_8562,N_8467);
or U8619 (N_8619,N_8576,N_8411);
nor U8620 (N_8620,N_8515,N_8452);
and U8621 (N_8621,N_8413,N_8425);
xnor U8622 (N_8622,N_8499,N_8459);
and U8623 (N_8623,N_8478,N_8421);
xor U8624 (N_8624,N_8496,N_8487);
xnor U8625 (N_8625,N_8426,N_8430);
nand U8626 (N_8626,N_8589,N_8575);
nor U8627 (N_8627,N_8535,N_8528);
or U8628 (N_8628,N_8460,N_8597);
nor U8629 (N_8629,N_8412,N_8500);
or U8630 (N_8630,N_8472,N_8433);
or U8631 (N_8631,N_8480,N_8409);
xor U8632 (N_8632,N_8596,N_8463);
nand U8633 (N_8633,N_8469,N_8438);
and U8634 (N_8634,N_8415,N_8507);
nand U8635 (N_8635,N_8519,N_8486);
nand U8636 (N_8636,N_8403,N_8422);
nor U8637 (N_8637,N_8468,N_8572);
and U8638 (N_8638,N_8598,N_8553);
xor U8639 (N_8639,N_8447,N_8588);
nand U8640 (N_8640,N_8504,N_8585);
nand U8641 (N_8641,N_8561,N_8442);
nand U8642 (N_8642,N_8557,N_8456);
xnor U8643 (N_8643,N_8584,N_8551);
nor U8644 (N_8644,N_8592,N_8462);
or U8645 (N_8645,N_8445,N_8428);
and U8646 (N_8646,N_8558,N_8440);
nand U8647 (N_8647,N_8443,N_8534);
xnor U8648 (N_8648,N_8527,N_8524);
xor U8649 (N_8649,N_8570,N_8521);
xor U8650 (N_8650,N_8434,N_8473);
and U8651 (N_8651,N_8586,N_8525);
and U8652 (N_8652,N_8509,N_8548);
and U8653 (N_8653,N_8568,N_8567);
xor U8654 (N_8654,N_8419,N_8531);
nor U8655 (N_8655,N_8446,N_8579);
nor U8656 (N_8656,N_8492,N_8424);
and U8657 (N_8657,N_8520,N_8436);
or U8658 (N_8658,N_8530,N_8587);
nand U8659 (N_8659,N_8532,N_8569);
nand U8660 (N_8660,N_8407,N_8482);
and U8661 (N_8661,N_8503,N_8540);
nor U8662 (N_8662,N_8449,N_8529);
xnor U8663 (N_8663,N_8429,N_8533);
nand U8664 (N_8664,N_8573,N_8526);
and U8665 (N_8665,N_8497,N_8593);
or U8666 (N_8666,N_8554,N_8510);
nor U8667 (N_8667,N_8511,N_8544);
nor U8668 (N_8668,N_8506,N_8556);
xor U8669 (N_8669,N_8517,N_8546);
nand U8670 (N_8670,N_8439,N_8471);
nor U8671 (N_8671,N_8454,N_8577);
xor U8672 (N_8672,N_8475,N_8427);
xor U8673 (N_8673,N_8574,N_8539);
nand U8674 (N_8674,N_8555,N_8501);
nor U8675 (N_8675,N_8477,N_8420);
or U8676 (N_8676,N_8455,N_8453);
or U8677 (N_8677,N_8543,N_8485);
xor U8678 (N_8678,N_8470,N_8410);
and U8679 (N_8679,N_8538,N_8565);
and U8680 (N_8680,N_8488,N_8465);
or U8681 (N_8681,N_8432,N_8513);
nand U8682 (N_8682,N_8406,N_8580);
nor U8683 (N_8683,N_8512,N_8414);
nand U8684 (N_8684,N_8505,N_8491);
and U8685 (N_8685,N_8502,N_8536);
or U8686 (N_8686,N_8563,N_8594);
and U8687 (N_8687,N_8560,N_8591);
and U8688 (N_8688,N_8595,N_8481);
nor U8689 (N_8689,N_8542,N_8418);
or U8690 (N_8690,N_8423,N_8466);
xor U8691 (N_8691,N_8508,N_8450);
xnor U8692 (N_8692,N_8599,N_8583);
and U8693 (N_8693,N_8437,N_8582);
nor U8694 (N_8694,N_8590,N_8458);
nand U8695 (N_8695,N_8448,N_8489);
nand U8696 (N_8696,N_8547,N_8408);
and U8697 (N_8697,N_8522,N_8479);
xnor U8698 (N_8698,N_8552,N_8461);
and U8699 (N_8699,N_8402,N_8405);
xor U8700 (N_8700,N_8459,N_8556);
or U8701 (N_8701,N_8576,N_8548);
xor U8702 (N_8702,N_8418,N_8404);
nor U8703 (N_8703,N_8450,N_8563);
nand U8704 (N_8704,N_8491,N_8504);
nand U8705 (N_8705,N_8524,N_8403);
or U8706 (N_8706,N_8525,N_8537);
nor U8707 (N_8707,N_8471,N_8477);
nand U8708 (N_8708,N_8465,N_8577);
nor U8709 (N_8709,N_8509,N_8500);
and U8710 (N_8710,N_8436,N_8516);
nor U8711 (N_8711,N_8597,N_8535);
and U8712 (N_8712,N_8541,N_8510);
xor U8713 (N_8713,N_8547,N_8534);
or U8714 (N_8714,N_8450,N_8402);
nor U8715 (N_8715,N_8565,N_8530);
or U8716 (N_8716,N_8523,N_8457);
nand U8717 (N_8717,N_8542,N_8482);
nor U8718 (N_8718,N_8589,N_8420);
nand U8719 (N_8719,N_8564,N_8516);
and U8720 (N_8720,N_8472,N_8564);
and U8721 (N_8721,N_8475,N_8493);
xor U8722 (N_8722,N_8460,N_8529);
nor U8723 (N_8723,N_8446,N_8428);
nand U8724 (N_8724,N_8595,N_8556);
nor U8725 (N_8725,N_8576,N_8567);
or U8726 (N_8726,N_8462,N_8466);
and U8727 (N_8727,N_8417,N_8464);
xnor U8728 (N_8728,N_8549,N_8492);
nand U8729 (N_8729,N_8469,N_8530);
and U8730 (N_8730,N_8406,N_8442);
nand U8731 (N_8731,N_8483,N_8572);
xnor U8732 (N_8732,N_8402,N_8577);
xnor U8733 (N_8733,N_8512,N_8537);
nor U8734 (N_8734,N_8460,N_8459);
xor U8735 (N_8735,N_8400,N_8559);
or U8736 (N_8736,N_8496,N_8572);
nor U8737 (N_8737,N_8528,N_8488);
or U8738 (N_8738,N_8572,N_8597);
nor U8739 (N_8739,N_8568,N_8409);
xnor U8740 (N_8740,N_8455,N_8445);
or U8741 (N_8741,N_8540,N_8441);
nor U8742 (N_8742,N_8400,N_8567);
or U8743 (N_8743,N_8579,N_8523);
xnor U8744 (N_8744,N_8414,N_8426);
and U8745 (N_8745,N_8576,N_8503);
and U8746 (N_8746,N_8455,N_8505);
xor U8747 (N_8747,N_8504,N_8593);
and U8748 (N_8748,N_8472,N_8414);
and U8749 (N_8749,N_8451,N_8400);
nand U8750 (N_8750,N_8576,N_8401);
and U8751 (N_8751,N_8580,N_8506);
and U8752 (N_8752,N_8436,N_8424);
nand U8753 (N_8753,N_8472,N_8574);
or U8754 (N_8754,N_8447,N_8599);
or U8755 (N_8755,N_8425,N_8545);
or U8756 (N_8756,N_8563,N_8473);
xor U8757 (N_8757,N_8470,N_8529);
nand U8758 (N_8758,N_8596,N_8597);
nand U8759 (N_8759,N_8404,N_8541);
nor U8760 (N_8760,N_8435,N_8407);
nor U8761 (N_8761,N_8536,N_8486);
xor U8762 (N_8762,N_8532,N_8442);
nand U8763 (N_8763,N_8509,N_8409);
and U8764 (N_8764,N_8408,N_8496);
nand U8765 (N_8765,N_8593,N_8521);
nand U8766 (N_8766,N_8543,N_8437);
nor U8767 (N_8767,N_8512,N_8442);
xnor U8768 (N_8768,N_8531,N_8568);
nor U8769 (N_8769,N_8407,N_8442);
and U8770 (N_8770,N_8462,N_8570);
xnor U8771 (N_8771,N_8410,N_8451);
nand U8772 (N_8772,N_8428,N_8479);
or U8773 (N_8773,N_8491,N_8519);
xnor U8774 (N_8774,N_8491,N_8417);
or U8775 (N_8775,N_8563,N_8461);
nand U8776 (N_8776,N_8558,N_8568);
xor U8777 (N_8777,N_8433,N_8520);
or U8778 (N_8778,N_8598,N_8548);
nor U8779 (N_8779,N_8441,N_8543);
nand U8780 (N_8780,N_8447,N_8456);
nand U8781 (N_8781,N_8473,N_8409);
nand U8782 (N_8782,N_8488,N_8504);
or U8783 (N_8783,N_8527,N_8422);
and U8784 (N_8784,N_8467,N_8564);
nand U8785 (N_8785,N_8452,N_8491);
nand U8786 (N_8786,N_8568,N_8499);
xor U8787 (N_8787,N_8415,N_8521);
nand U8788 (N_8788,N_8412,N_8415);
and U8789 (N_8789,N_8488,N_8546);
xor U8790 (N_8790,N_8489,N_8593);
xnor U8791 (N_8791,N_8516,N_8507);
nor U8792 (N_8792,N_8587,N_8436);
or U8793 (N_8793,N_8450,N_8550);
nand U8794 (N_8794,N_8452,N_8419);
nand U8795 (N_8795,N_8547,N_8544);
or U8796 (N_8796,N_8403,N_8407);
and U8797 (N_8797,N_8438,N_8523);
or U8798 (N_8798,N_8566,N_8449);
nor U8799 (N_8799,N_8535,N_8520);
nand U8800 (N_8800,N_8790,N_8789);
nor U8801 (N_8801,N_8780,N_8623);
or U8802 (N_8802,N_8798,N_8708);
or U8803 (N_8803,N_8713,N_8601);
nor U8804 (N_8804,N_8638,N_8744);
nor U8805 (N_8805,N_8706,N_8689);
nor U8806 (N_8806,N_8752,N_8709);
and U8807 (N_8807,N_8625,N_8653);
nand U8808 (N_8808,N_8616,N_8721);
xnor U8809 (N_8809,N_8639,N_8640);
xor U8810 (N_8810,N_8655,N_8705);
or U8811 (N_8811,N_8676,N_8756);
nor U8812 (N_8812,N_8604,N_8611);
and U8813 (N_8813,N_8762,N_8624);
nand U8814 (N_8814,N_8675,N_8658);
nor U8815 (N_8815,N_8618,N_8696);
or U8816 (N_8816,N_8626,N_8636);
nand U8817 (N_8817,N_8677,N_8628);
nand U8818 (N_8818,N_8695,N_8702);
and U8819 (N_8819,N_8612,N_8667);
nand U8820 (N_8820,N_8759,N_8620);
xnor U8821 (N_8821,N_8645,N_8678);
and U8822 (N_8822,N_8686,N_8615);
xor U8823 (N_8823,N_8666,N_8783);
nor U8824 (N_8824,N_8730,N_8755);
and U8825 (N_8825,N_8734,N_8773);
xor U8826 (N_8826,N_8778,N_8766);
and U8827 (N_8827,N_8697,N_8673);
and U8828 (N_8828,N_8661,N_8793);
nor U8829 (N_8829,N_8745,N_8649);
nor U8830 (N_8830,N_8664,N_8605);
nor U8831 (N_8831,N_8725,N_8613);
and U8832 (N_8832,N_8719,N_8718);
nand U8833 (N_8833,N_8707,N_8796);
or U8834 (N_8834,N_8654,N_8632);
and U8835 (N_8835,N_8679,N_8672);
and U8836 (N_8836,N_8750,N_8600);
and U8837 (N_8837,N_8743,N_8629);
and U8838 (N_8838,N_8799,N_8746);
nor U8839 (N_8839,N_8668,N_8770);
and U8840 (N_8840,N_8619,N_8761);
and U8841 (N_8841,N_8650,N_8603);
or U8842 (N_8842,N_8665,N_8757);
and U8843 (N_8843,N_8610,N_8714);
xor U8844 (N_8844,N_8739,N_8726);
nor U8845 (N_8845,N_8776,N_8791);
nand U8846 (N_8846,N_8737,N_8728);
nand U8847 (N_8847,N_8662,N_8674);
nor U8848 (N_8848,N_8787,N_8720);
nor U8849 (N_8849,N_8749,N_8642);
nor U8850 (N_8850,N_8663,N_8742);
nor U8851 (N_8851,N_8758,N_8648);
or U8852 (N_8852,N_8711,N_8703);
xor U8853 (N_8853,N_8659,N_8701);
or U8854 (N_8854,N_8748,N_8797);
nor U8855 (N_8855,N_8607,N_8680);
nor U8856 (N_8856,N_8781,N_8777);
nor U8857 (N_8857,N_8753,N_8786);
and U8858 (N_8858,N_8691,N_8763);
or U8859 (N_8859,N_8670,N_8682);
and U8860 (N_8860,N_8699,N_8723);
or U8861 (N_8861,N_8602,N_8647);
nor U8862 (N_8862,N_8774,N_8657);
nor U8863 (N_8863,N_8710,N_8608);
nand U8864 (N_8864,N_8693,N_8754);
nand U8865 (N_8865,N_8617,N_8732);
nand U8866 (N_8866,N_8651,N_8733);
xor U8867 (N_8867,N_8768,N_8669);
and U8868 (N_8868,N_8769,N_8717);
and U8869 (N_8869,N_8627,N_8779);
xor U8870 (N_8870,N_8606,N_8643);
and U8871 (N_8871,N_8637,N_8614);
and U8872 (N_8872,N_8751,N_8767);
nand U8873 (N_8873,N_8631,N_8630);
or U8874 (N_8874,N_8688,N_8740);
xor U8875 (N_8875,N_8684,N_8634);
nand U8876 (N_8876,N_8722,N_8785);
xnor U8877 (N_8877,N_8681,N_8738);
and U8878 (N_8878,N_8788,N_8795);
xnor U8879 (N_8879,N_8741,N_8646);
nand U8880 (N_8880,N_8633,N_8644);
and U8881 (N_8881,N_8690,N_8635);
xnor U8882 (N_8882,N_8747,N_8764);
nor U8883 (N_8883,N_8671,N_8683);
and U8884 (N_8884,N_8724,N_8692);
or U8885 (N_8885,N_8784,N_8727);
and U8886 (N_8886,N_8735,N_8772);
or U8887 (N_8887,N_8609,N_8687);
nor U8888 (N_8888,N_8792,N_8729);
xnor U8889 (N_8889,N_8621,N_8694);
xor U8890 (N_8890,N_8656,N_8641);
and U8891 (N_8891,N_8760,N_8698);
xor U8892 (N_8892,N_8715,N_8771);
xor U8893 (N_8893,N_8736,N_8712);
nand U8894 (N_8894,N_8700,N_8652);
nand U8895 (N_8895,N_8716,N_8622);
nand U8896 (N_8896,N_8765,N_8731);
xor U8897 (N_8897,N_8685,N_8782);
nand U8898 (N_8898,N_8775,N_8704);
nor U8899 (N_8899,N_8794,N_8660);
nor U8900 (N_8900,N_8740,N_8733);
or U8901 (N_8901,N_8643,N_8657);
nor U8902 (N_8902,N_8736,N_8700);
and U8903 (N_8903,N_8609,N_8705);
or U8904 (N_8904,N_8660,N_8677);
and U8905 (N_8905,N_8787,N_8644);
and U8906 (N_8906,N_8615,N_8707);
nand U8907 (N_8907,N_8613,N_8600);
nor U8908 (N_8908,N_8614,N_8762);
xnor U8909 (N_8909,N_8620,N_8794);
and U8910 (N_8910,N_8747,N_8729);
nor U8911 (N_8911,N_8730,N_8712);
or U8912 (N_8912,N_8648,N_8792);
nor U8913 (N_8913,N_8780,N_8676);
nand U8914 (N_8914,N_8701,N_8727);
xnor U8915 (N_8915,N_8696,N_8660);
nor U8916 (N_8916,N_8627,N_8783);
or U8917 (N_8917,N_8615,N_8689);
xnor U8918 (N_8918,N_8681,N_8795);
and U8919 (N_8919,N_8665,N_8607);
nor U8920 (N_8920,N_8695,N_8602);
and U8921 (N_8921,N_8722,N_8742);
nand U8922 (N_8922,N_8616,N_8610);
nand U8923 (N_8923,N_8639,N_8737);
nor U8924 (N_8924,N_8638,N_8750);
xnor U8925 (N_8925,N_8687,N_8645);
nand U8926 (N_8926,N_8650,N_8623);
nor U8927 (N_8927,N_8772,N_8681);
and U8928 (N_8928,N_8614,N_8685);
nand U8929 (N_8929,N_8606,N_8717);
and U8930 (N_8930,N_8726,N_8799);
or U8931 (N_8931,N_8791,N_8680);
and U8932 (N_8932,N_8795,N_8777);
xnor U8933 (N_8933,N_8688,N_8664);
xnor U8934 (N_8934,N_8789,N_8776);
nand U8935 (N_8935,N_8642,N_8692);
xnor U8936 (N_8936,N_8685,N_8750);
xnor U8937 (N_8937,N_8682,N_8785);
xor U8938 (N_8938,N_8651,N_8619);
nor U8939 (N_8939,N_8729,N_8778);
xnor U8940 (N_8940,N_8714,N_8672);
and U8941 (N_8941,N_8610,N_8778);
xnor U8942 (N_8942,N_8650,N_8729);
or U8943 (N_8943,N_8761,N_8638);
xor U8944 (N_8944,N_8796,N_8714);
nor U8945 (N_8945,N_8661,N_8637);
nand U8946 (N_8946,N_8676,N_8771);
nor U8947 (N_8947,N_8783,N_8680);
xnor U8948 (N_8948,N_8641,N_8685);
or U8949 (N_8949,N_8655,N_8649);
xor U8950 (N_8950,N_8601,N_8633);
nand U8951 (N_8951,N_8670,N_8631);
or U8952 (N_8952,N_8672,N_8710);
and U8953 (N_8953,N_8640,N_8766);
xnor U8954 (N_8954,N_8662,N_8717);
or U8955 (N_8955,N_8642,N_8702);
or U8956 (N_8956,N_8783,N_8720);
and U8957 (N_8957,N_8743,N_8621);
or U8958 (N_8958,N_8602,N_8636);
or U8959 (N_8959,N_8767,N_8779);
and U8960 (N_8960,N_8694,N_8682);
or U8961 (N_8961,N_8760,N_8757);
nand U8962 (N_8962,N_8638,N_8664);
or U8963 (N_8963,N_8605,N_8614);
nor U8964 (N_8964,N_8744,N_8632);
or U8965 (N_8965,N_8703,N_8668);
nand U8966 (N_8966,N_8712,N_8624);
nand U8967 (N_8967,N_8690,N_8766);
nor U8968 (N_8968,N_8663,N_8764);
and U8969 (N_8969,N_8766,N_8765);
and U8970 (N_8970,N_8684,N_8734);
or U8971 (N_8971,N_8620,N_8601);
nor U8972 (N_8972,N_8717,N_8689);
xnor U8973 (N_8973,N_8735,N_8708);
nor U8974 (N_8974,N_8644,N_8677);
xor U8975 (N_8975,N_8732,N_8609);
xor U8976 (N_8976,N_8636,N_8794);
nor U8977 (N_8977,N_8701,N_8610);
or U8978 (N_8978,N_8789,N_8702);
nor U8979 (N_8979,N_8662,N_8759);
nor U8980 (N_8980,N_8651,N_8612);
nand U8981 (N_8981,N_8687,N_8748);
nor U8982 (N_8982,N_8606,N_8795);
nor U8983 (N_8983,N_8610,N_8666);
xnor U8984 (N_8984,N_8755,N_8622);
nor U8985 (N_8985,N_8784,N_8604);
and U8986 (N_8986,N_8758,N_8621);
and U8987 (N_8987,N_8718,N_8602);
or U8988 (N_8988,N_8761,N_8622);
nor U8989 (N_8989,N_8677,N_8688);
nor U8990 (N_8990,N_8675,N_8663);
xor U8991 (N_8991,N_8612,N_8639);
nor U8992 (N_8992,N_8660,N_8743);
xor U8993 (N_8993,N_8713,N_8618);
nand U8994 (N_8994,N_8757,N_8621);
or U8995 (N_8995,N_8764,N_8619);
nor U8996 (N_8996,N_8677,N_8734);
or U8997 (N_8997,N_8735,N_8762);
xnor U8998 (N_8998,N_8632,N_8771);
and U8999 (N_8999,N_8609,N_8601);
or U9000 (N_9000,N_8861,N_8800);
and U9001 (N_9001,N_8853,N_8995);
nor U9002 (N_9002,N_8848,N_8875);
and U9003 (N_9003,N_8865,N_8982);
nand U9004 (N_9004,N_8878,N_8887);
nor U9005 (N_9005,N_8916,N_8809);
nand U9006 (N_9006,N_8830,N_8872);
nor U9007 (N_9007,N_8844,N_8994);
and U9008 (N_9008,N_8979,N_8886);
nand U9009 (N_9009,N_8914,N_8836);
xnor U9010 (N_9010,N_8971,N_8907);
or U9011 (N_9011,N_8957,N_8975);
xnor U9012 (N_9012,N_8808,N_8877);
nor U9013 (N_9013,N_8821,N_8804);
nor U9014 (N_9014,N_8807,N_8850);
nor U9015 (N_9015,N_8978,N_8879);
or U9016 (N_9016,N_8984,N_8945);
nor U9017 (N_9017,N_8938,N_8827);
nand U9018 (N_9018,N_8963,N_8866);
or U9019 (N_9019,N_8841,N_8825);
nor U9020 (N_9020,N_8837,N_8968);
nand U9021 (N_9021,N_8838,N_8992);
or U9022 (N_9022,N_8986,N_8997);
or U9023 (N_9023,N_8983,N_8911);
or U9024 (N_9024,N_8927,N_8820);
nand U9025 (N_9025,N_8881,N_8976);
nor U9026 (N_9026,N_8828,N_8895);
xor U9027 (N_9027,N_8922,N_8989);
or U9028 (N_9028,N_8990,N_8977);
nand U9029 (N_9029,N_8954,N_8998);
nand U9030 (N_9030,N_8882,N_8965);
nor U9031 (N_9031,N_8919,N_8801);
nor U9032 (N_9032,N_8930,N_8867);
and U9033 (N_9033,N_8842,N_8924);
xor U9034 (N_9034,N_8833,N_8896);
nand U9035 (N_9035,N_8824,N_8869);
nor U9036 (N_9036,N_8901,N_8818);
nand U9037 (N_9037,N_8888,N_8910);
nand U9038 (N_9038,N_8811,N_8972);
nor U9039 (N_9039,N_8864,N_8857);
nor U9040 (N_9040,N_8943,N_8813);
nand U9041 (N_9041,N_8966,N_8880);
and U9042 (N_9042,N_8959,N_8862);
and U9043 (N_9043,N_8918,N_8906);
or U9044 (N_9044,N_8812,N_8900);
and U9045 (N_9045,N_8973,N_8981);
nand U9046 (N_9046,N_8958,N_8898);
nor U9047 (N_9047,N_8937,N_8969);
nor U9048 (N_9048,N_8894,N_8935);
or U9049 (N_9049,N_8939,N_8913);
nand U9050 (N_9050,N_8967,N_8846);
nand U9051 (N_9051,N_8993,N_8819);
xor U9052 (N_9052,N_8936,N_8917);
xor U9053 (N_9053,N_8823,N_8840);
and U9054 (N_9054,N_8929,N_8904);
nor U9055 (N_9055,N_8860,N_8934);
and U9056 (N_9056,N_8832,N_8970);
and U9057 (N_9057,N_8871,N_8834);
or U9058 (N_9058,N_8858,N_8814);
or U9059 (N_9059,N_8831,N_8933);
or U9060 (N_9060,N_8928,N_8946);
nand U9061 (N_9061,N_8817,N_8845);
xor U9062 (N_9062,N_8985,N_8892);
or U9063 (N_9063,N_8921,N_8893);
nor U9064 (N_9064,N_8868,N_8839);
nor U9065 (N_9065,N_8884,N_8950);
and U9066 (N_9066,N_8852,N_8903);
nand U9067 (N_9067,N_8932,N_8908);
nor U9068 (N_9068,N_8951,N_8961);
xor U9069 (N_9069,N_8905,N_8851);
xnor U9070 (N_9070,N_8854,N_8948);
or U9071 (N_9071,N_8835,N_8956);
and U9072 (N_9072,N_8806,N_8947);
and U9073 (N_9073,N_8964,N_8941);
and U9074 (N_9074,N_8876,N_8889);
or U9075 (N_9075,N_8909,N_8870);
nand U9076 (N_9076,N_8874,N_8859);
nor U9077 (N_9077,N_8829,N_8923);
nor U9078 (N_9078,N_8805,N_8897);
and U9079 (N_9079,N_8940,N_8952);
xor U9080 (N_9080,N_8942,N_8912);
nor U9081 (N_9081,N_8953,N_8926);
nand U9082 (N_9082,N_8944,N_8890);
nor U9083 (N_9083,N_8987,N_8999);
nor U9084 (N_9084,N_8980,N_8920);
and U9085 (N_9085,N_8974,N_8991);
nand U9086 (N_9086,N_8891,N_8988);
nand U9087 (N_9087,N_8962,N_8843);
xor U9088 (N_9088,N_8815,N_8931);
nor U9089 (N_9089,N_8810,N_8802);
nand U9090 (N_9090,N_8955,N_8960);
nor U9091 (N_9091,N_8863,N_8883);
or U9092 (N_9092,N_8816,N_8847);
xor U9093 (N_9093,N_8873,N_8826);
or U9094 (N_9094,N_8925,N_8803);
nor U9095 (N_9095,N_8856,N_8885);
nor U9096 (N_9096,N_8915,N_8855);
nand U9097 (N_9097,N_8902,N_8949);
nor U9098 (N_9098,N_8822,N_8899);
nor U9099 (N_9099,N_8849,N_8996);
and U9100 (N_9100,N_8812,N_8906);
and U9101 (N_9101,N_8820,N_8877);
nor U9102 (N_9102,N_8943,N_8965);
nor U9103 (N_9103,N_8842,N_8801);
nand U9104 (N_9104,N_8956,N_8963);
nor U9105 (N_9105,N_8893,N_8930);
nand U9106 (N_9106,N_8812,N_8854);
xnor U9107 (N_9107,N_8948,N_8890);
nor U9108 (N_9108,N_8825,N_8840);
nand U9109 (N_9109,N_8849,N_8941);
nor U9110 (N_9110,N_8873,N_8993);
nand U9111 (N_9111,N_8821,N_8834);
nor U9112 (N_9112,N_8877,N_8992);
and U9113 (N_9113,N_8871,N_8802);
nand U9114 (N_9114,N_8893,N_8957);
xnor U9115 (N_9115,N_8830,N_8957);
nor U9116 (N_9116,N_8895,N_8979);
xor U9117 (N_9117,N_8972,N_8948);
xor U9118 (N_9118,N_8801,N_8957);
nand U9119 (N_9119,N_8975,N_8823);
xnor U9120 (N_9120,N_8997,N_8830);
and U9121 (N_9121,N_8948,N_8899);
nand U9122 (N_9122,N_8832,N_8844);
and U9123 (N_9123,N_8973,N_8965);
nor U9124 (N_9124,N_8854,N_8983);
xor U9125 (N_9125,N_8890,N_8907);
and U9126 (N_9126,N_8848,N_8957);
and U9127 (N_9127,N_8817,N_8949);
xnor U9128 (N_9128,N_8891,N_8857);
xnor U9129 (N_9129,N_8836,N_8981);
or U9130 (N_9130,N_8951,N_8896);
and U9131 (N_9131,N_8928,N_8861);
or U9132 (N_9132,N_8962,N_8866);
xor U9133 (N_9133,N_8940,N_8931);
and U9134 (N_9134,N_8871,N_8982);
nand U9135 (N_9135,N_8808,N_8919);
xor U9136 (N_9136,N_8846,N_8833);
and U9137 (N_9137,N_8898,N_8933);
or U9138 (N_9138,N_8874,N_8961);
nor U9139 (N_9139,N_8937,N_8869);
or U9140 (N_9140,N_8977,N_8852);
nand U9141 (N_9141,N_8976,N_8902);
or U9142 (N_9142,N_8933,N_8814);
or U9143 (N_9143,N_8816,N_8806);
nor U9144 (N_9144,N_8904,N_8901);
nor U9145 (N_9145,N_8987,N_8815);
or U9146 (N_9146,N_8976,N_8985);
and U9147 (N_9147,N_8980,N_8889);
nand U9148 (N_9148,N_8979,N_8919);
nor U9149 (N_9149,N_8992,N_8821);
nor U9150 (N_9150,N_8967,N_8812);
or U9151 (N_9151,N_8975,N_8838);
or U9152 (N_9152,N_8950,N_8892);
nor U9153 (N_9153,N_8860,N_8872);
nand U9154 (N_9154,N_8935,N_8921);
xnor U9155 (N_9155,N_8950,N_8963);
xnor U9156 (N_9156,N_8832,N_8869);
nand U9157 (N_9157,N_8828,N_8906);
or U9158 (N_9158,N_8945,N_8866);
xor U9159 (N_9159,N_8803,N_8897);
nor U9160 (N_9160,N_8907,N_8910);
or U9161 (N_9161,N_8977,N_8943);
nor U9162 (N_9162,N_8891,N_8960);
xor U9163 (N_9163,N_8979,N_8855);
xor U9164 (N_9164,N_8936,N_8863);
or U9165 (N_9165,N_8956,N_8916);
or U9166 (N_9166,N_8937,N_8971);
nand U9167 (N_9167,N_8833,N_8881);
or U9168 (N_9168,N_8994,N_8949);
and U9169 (N_9169,N_8982,N_8826);
nor U9170 (N_9170,N_8840,N_8904);
nand U9171 (N_9171,N_8827,N_8849);
xor U9172 (N_9172,N_8934,N_8967);
nand U9173 (N_9173,N_8956,N_8803);
nand U9174 (N_9174,N_8847,N_8992);
nor U9175 (N_9175,N_8850,N_8927);
or U9176 (N_9176,N_8890,N_8993);
and U9177 (N_9177,N_8940,N_8848);
nor U9178 (N_9178,N_8902,N_8906);
nand U9179 (N_9179,N_8903,N_8810);
nor U9180 (N_9180,N_8938,N_8876);
and U9181 (N_9181,N_8833,N_8961);
xnor U9182 (N_9182,N_8940,N_8849);
xor U9183 (N_9183,N_8921,N_8950);
nor U9184 (N_9184,N_8933,N_8905);
nand U9185 (N_9185,N_8948,N_8827);
nor U9186 (N_9186,N_8925,N_8808);
or U9187 (N_9187,N_8916,N_8822);
nand U9188 (N_9188,N_8896,N_8979);
and U9189 (N_9189,N_8900,N_8845);
and U9190 (N_9190,N_8935,N_8975);
nor U9191 (N_9191,N_8913,N_8805);
nand U9192 (N_9192,N_8870,N_8849);
or U9193 (N_9193,N_8998,N_8875);
nand U9194 (N_9194,N_8998,N_8812);
and U9195 (N_9195,N_8926,N_8844);
nor U9196 (N_9196,N_8896,N_8830);
or U9197 (N_9197,N_8951,N_8994);
nand U9198 (N_9198,N_8892,N_8992);
nor U9199 (N_9199,N_8832,N_8939);
nor U9200 (N_9200,N_9071,N_9173);
and U9201 (N_9201,N_9106,N_9149);
or U9202 (N_9202,N_9096,N_9053);
and U9203 (N_9203,N_9188,N_9196);
xnor U9204 (N_9204,N_9075,N_9197);
nor U9205 (N_9205,N_9021,N_9044);
nor U9206 (N_9206,N_9034,N_9001);
nor U9207 (N_9207,N_9003,N_9008);
nor U9208 (N_9208,N_9059,N_9088);
or U9209 (N_9209,N_9028,N_9045);
nor U9210 (N_9210,N_9011,N_9054);
xor U9211 (N_9211,N_9010,N_9113);
nand U9212 (N_9212,N_9012,N_9142);
nand U9213 (N_9213,N_9024,N_9103);
and U9214 (N_9214,N_9018,N_9186);
nand U9215 (N_9215,N_9105,N_9157);
nand U9216 (N_9216,N_9079,N_9144);
nor U9217 (N_9217,N_9146,N_9027);
xnor U9218 (N_9218,N_9058,N_9162);
and U9219 (N_9219,N_9017,N_9181);
or U9220 (N_9220,N_9180,N_9099);
xor U9221 (N_9221,N_9118,N_9013);
nor U9222 (N_9222,N_9085,N_9155);
nand U9223 (N_9223,N_9168,N_9066);
or U9224 (N_9224,N_9092,N_9026);
nor U9225 (N_9225,N_9110,N_9035);
nand U9226 (N_9226,N_9137,N_9151);
nand U9227 (N_9227,N_9190,N_9081);
or U9228 (N_9228,N_9117,N_9154);
nand U9229 (N_9229,N_9130,N_9101);
nand U9230 (N_9230,N_9068,N_9089);
nand U9231 (N_9231,N_9177,N_9160);
xnor U9232 (N_9232,N_9098,N_9090);
nor U9233 (N_9233,N_9121,N_9172);
or U9234 (N_9234,N_9127,N_9174);
and U9235 (N_9235,N_9187,N_9124);
nand U9236 (N_9236,N_9108,N_9049);
and U9237 (N_9237,N_9133,N_9119);
xnor U9238 (N_9238,N_9025,N_9175);
or U9239 (N_9239,N_9120,N_9036);
nand U9240 (N_9240,N_9194,N_9063);
or U9241 (N_9241,N_9114,N_9007);
xnor U9242 (N_9242,N_9064,N_9166);
nor U9243 (N_9243,N_9082,N_9072);
xnor U9244 (N_9244,N_9163,N_9104);
and U9245 (N_9245,N_9009,N_9062);
xnor U9246 (N_9246,N_9037,N_9171);
or U9247 (N_9247,N_9057,N_9055);
xnor U9248 (N_9248,N_9023,N_9091);
nor U9249 (N_9249,N_9076,N_9086);
nor U9250 (N_9250,N_9165,N_9056);
or U9251 (N_9251,N_9147,N_9169);
or U9252 (N_9252,N_9067,N_9093);
xnor U9253 (N_9253,N_9183,N_9170);
nor U9254 (N_9254,N_9195,N_9191);
and U9255 (N_9255,N_9031,N_9061);
or U9256 (N_9256,N_9135,N_9116);
xnor U9257 (N_9257,N_9070,N_9129);
and U9258 (N_9258,N_9193,N_9131);
xor U9259 (N_9259,N_9159,N_9176);
xnor U9260 (N_9260,N_9128,N_9132);
nor U9261 (N_9261,N_9123,N_9178);
nor U9262 (N_9262,N_9014,N_9006);
and U9263 (N_9263,N_9094,N_9136);
nand U9264 (N_9264,N_9039,N_9115);
xnor U9265 (N_9265,N_9033,N_9029);
or U9266 (N_9266,N_9046,N_9185);
nor U9267 (N_9267,N_9153,N_9087);
nor U9268 (N_9268,N_9016,N_9140);
nand U9269 (N_9269,N_9002,N_9112);
xor U9270 (N_9270,N_9150,N_9005);
nand U9271 (N_9271,N_9161,N_9109);
nor U9272 (N_9272,N_9019,N_9138);
nand U9273 (N_9273,N_9041,N_9156);
and U9274 (N_9274,N_9148,N_9020);
nand U9275 (N_9275,N_9050,N_9189);
or U9276 (N_9276,N_9182,N_9032);
and U9277 (N_9277,N_9065,N_9083);
xnor U9278 (N_9278,N_9069,N_9000);
nand U9279 (N_9279,N_9122,N_9125);
or U9280 (N_9280,N_9184,N_9080);
and U9281 (N_9281,N_9152,N_9052);
nand U9282 (N_9282,N_9164,N_9084);
and U9283 (N_9283,N_9199,N_9145);
xnor U9284 (N_9284,N_9038,N_9179);
and U9285 (N_9285,N_9048,N_9167);
nor U9286 (N_9286,N_9047,N_9015);
and U9287 (N_9287,N_9107,N_9078);
nor U9288 (N_9288,N_9051,N_9192);
or U9289 (N_9289,N_9074,N_9043);
or U9290 (N_9290,N_9040,N_9060);
or U9291 (N_9291,N_9077,N_9022);
nor U9292 (N_9292,N_9134,N_9097);
and U9293 (N_9293,N_9095,N_9030);
or U9294 (N_9294,N_9042,N_9198);
nand U9295 (N_9295,N_9111,N_9126);
xnor U9296 (N_9296,N_9102,N_9141);
xnor U9297 (N_9297,N_9004,N_9139);
xor U9298 (N_9298,N_9073,N_9143);
nor U9299 (N_9299,N_9100,N_9158);
or U9300 (N_9300,N_9087,N_9048);
nor U9301 (N_9301,N_9035,N_9119);
or U9302 (N_9302,N_9056,N_9098);
nor U9303 (N_9303,N_9057,N_9064);
nor U9304 (N_9304,N_9139,N_9049);
and U9305 (N_9305,N_9138,N_9065);
and U9306 (N_9306,N_9129,N_9096);
or U9307 (N_9307,N_9107,N_9079);
xor U9308 (N_9308,N_9102,N_9068);
nor U9309 (N_9309,N_9138,N_9166);
nand U9310 (N_9310,N_9079,N_9080);
and U9311 (N_9311,N_9115,N_9008);
nor U9312 (N_9312,N_9185,N_9194);
nor U9313 (N_9313,N_9054,N_9166);
or U9314 (N_9314,N_9041,N_9036);
and U9315 (N_9315,N_9090,N_9023);
xnor U9316 (N_9316,N_9146,N_9137);
nand U9317 (N_9317,N_9147,N_9041);
nand U9318 (N_9318,N_9032,N_9037);
xnor U9319 (N_9319,N_9164,N_9089);
xnor U9320 (N_9320,N_9173,N_9191);
nand U9321 (N_9321,N_9001,N_9094);
nand U9322 (N_9322,N_9142,N_9179);
nor U9323 (N_9323,N_9159,N_9011);
or U9324 (N_9324,N_9087,N_9049);
or U9325 (N_9325,N_9045,N_9055);
and U9326 (N_9326,N_9042,N_9034);
nand U9327 (N_9327,N_9026,N_9022);
and U9328 (N_9328,N_9006,N_9089);
xnor U9329 (N_9329,N_9113,N_9018);
nand U9330 (N_9330,N_9057,N_9027);
and U9331 (N_9331,N_9101,N_9042);
xor U9332 (N_9332,N_9160,N_9182);
xor U9333 (N_9333,N_9012,N_9115);
or U9334 (N_9334,N_9012,N_9173);
and U9335 (N_9335,N_9055,N_9116);
nand U9336 (N_9336,N_9191,N_9084);
nand U9337 (N_9337,N_9065,N_9142);
nand U9338 (N_9338,N_9115,N_9015);
nand U9339 (N_9339,N_9196,N_9100);
xor U9340 (N_9340,N_9076,N_9071);
nand U9341 (N_9341,N_9005,N_9191);
nand U9342 (N_9342,N_9065,N_9042);
and U9343 (N_9343,N_9153,N_9079);
nand U9344 (N_9344,N_9102,N_9155);
xor U9345 (N_9345,N_9008,N_9004);
and U9346 (N_9346,N_9117,N_9188);
or U9347 (N_9347,N_9146,N_9111);
or U9348 (N_9348,N_9022,N_9120);
nand U9349 (N_9349,N_9120,N_9127);
nor U9350 (N_9350,N_9195,N_9078);
or U9351 (N_9351,N_9171,N_9022);
xor U9352 (N_9352,N_9045,N_9044);
or U9353 (N_9353,N_9092,N_9145);
or U9354 (N_9354,N_9139,N_9150);
nor U9355 (N_9355,N_9031,N_9149);
nor U9356 (N_9356,N_9111,N_9051);
and U9357 (N_9357,N_9159,N_9131);
or U9358 (N_9358,N_9171,N_9061);
and U9359 (N_9359,N_9181,N_9176);
xor U9360 (N_9360,N_9116,N_9016);
nor U9361 (N_9361,N_9016,N_9175);
xnor U9362 (N_9362,N_9160,N_9014);
nor U9363 (N_9363,N_9027,N_9148);
nand U9364 (N_9364,N_9161,N_9141);
nand U9365 (N_9365,N_9089,N_9025);
or U9366 (N_9366,N_9174,N_9005);
and U9367 (N_9367,N_9075,N_9021);
nor U9368 (N_9368,N_9018,N_9126);
nand U9369 (N_9369,N_9087,N_9017);
or U9370 (N_9370,N_9193,N_9006);
nand U9371 (N_9371,N_9167,N_9059);
nor U9372 (N_9372,N_9016,N_9022);
or U9373 (N_9373,N_9011,N_9039);
or U9374 (N_9374,N_9012,N_9180);
or U9375 (N_9375,N_9095,N_9055);
nand U9376 (N_9376,N_9143,N_9000);
and U9377 (N_9377,N_9019,N_9176);
nor U9378 (N_9378,N_9156,N_9010);
xnor U9379 (N_9379,N_9114,N_9130);
nor U9380 (N_9380,N_9196,N_9052);
or U9381 (N_9381,N_9065,N_9069);
nor U9382 (N_9382,N_9018,N_9044);
nor U9383 (N_9383,N_9134,N_9018);
and U9384 (N_9384,N_9146,N_9156);
and U9385 (N_9385,N_9015,N_9172);
nor U9386 (N_9386,N_9064,N_9030);
or U9387 (N_9387,N_9064,N_9077);
or U9388 (N_9388,N_9079,N_9176);
nor U9389 (N_9389,N_9102,N_9136);
and U9390 (N_9390,N_9032,N_9100);
and U9391 (N_9391,N_9092,N_9038);
and U9392 (N_9392,N_9009,N_9185);
and U9393 (N_9393,N_9124,N_9041);
xor U9394 (N_9394,N_9114,N_9140);
or U9395 (N_9395,N_9010,N_9030);
nand U9396 (N_9396,N_9170,N_9040);
nand U9397 (N_9397,N_9087,N_9064);
nand U9398 (N_9398,N_9107,N_9028);
xor U9399 (N_9399,N_9124,N_9132);
nand U9400 (N_9400,N_9242,N_9361);
nand U9401 (N_9401,N_9392,N_9397);
nor U9402 (N_9402,N_9266,N_9304);
nand U9403 (N_9403,N_9308,N_9319);
xor U9404 (N_9404,N_9366,N_9339);
nor U9405 (N_9405,N_9396,N_9325);
and U9406 (N_9406,N_9229,N_9281);
nor U9407 (N_9407,N_9323,N_9276);
and U9408 (N_9408,N_9215,N_9384);
or U9409 (N_9409,N_9399,N_9310);
nor U9410 (N_9410,N_9200,N_9327);
nand U9411 (N_9411,N_9303,N_9330);
xnor U9412 (N_9412,N_9243,N_9349);
xor U9413 (N_9413,N_9373,N_9360);
nor U9414 (N_9414,N_9237,N_9213);
nand U9415 (N_9415,N_9379,N_9205);
or U9416 (N_9416,N_9332,N_9282);
nand U9417 (N_9417,N_9317,N_9377);
nor U9418 (N_9418,N_9291,N_9220);
nor U9419 (N_9419,N_9395,N_9391);
nand U9420 (N_9420,N_9247,N_9259);
or U9421 (N_9421,N_9326,N_9324);
and U9422 (N_9422,N_9393,N_9212);
nor U9423 (N_9423,N_9275,N_9389);
nand U9424 (N_9424,N_9298,N_9255);
nor U9425 (N_9425,N_9257,N_9284);
nand U9426 (N_9426,N_9306,N_9348);
and U9427 (N_9427,N_9270,N_9353);
and U9428 (N_9428,N_9230,N_9253);
xnor U9429 (N_9429,N_9211,N_9309);
xnor U9430 (N_9430,N_9226,N_9394);
xor U9431 (N_9431,N_9370,N_9202);
xnor U9432 (N_9432,N_9254,N_9314);
and U9433 (N_9433,N_9374,N_9272);
xor U9434 (N_9434,N_9218,N_9346);
and U9435 (N_9435,N_9321,N_9358);
nor U9436 (N_9436,N_9355,N_9279);
nor U9437 (N_9437,N_9302,N_9273);
or U9438 (N_9438,N_9375,N_9288);
and U9439 (N_9439,N_9217,N_9268);
or U9440 (N_9440,N_9222,N_9381);
xor U9441 (N_9441,N_9250,N_9274);
and U9442 (N_9442,N_9277,N_9297);
and U9443 (N_9443,N_9296,N_9336);
nand U9444 (N_9444,N_9371,N_9283);
and U9445 (N_9445,N_9350,N_9345);
nand U9446 (N_9446,N_9278,N_9333);
xor U9447 (N_9447,N_9264,N_9285);
and U9448 (N_9448,N_9341,N_9347);
and U9449 (N_9449,N_9287,N_9357);
or U9450 (N_9450,N_9293,N_9311);
and U9451 (N_9451,N_9249,N_9224);
or U9452 (N_9452,N_9251,N_9385);
and U9453 (N_9453,N_9245,N_9322);
or U9454 (N_9454,N_9331,N_9235);
and U9455 (N_9455,N_9258,N_9263);
and U9456 (N_9456,N_9294,N_9378);
or U9457 (N_9457,N_9305,N_9221);
and U9458 (N_9458,N_9256,N_9313);
nand U9459 (N_9459,N_9398,N_9295);
xnor U9460 (N_9460,N_9340,N_9316);
nor U9461 (N_9461,N_9334,N_9388);
nand U9462 (N_9462,N_9338,N_9335);
xor U9463 (N_9463,N_9203,N_9301);
nand U9464 (N_9464,N_9239,N_9312);
xnor U9465 (N_9465,N_9367,N_9329);
xor U9466 (N_9466,N_9286,N_9364);
or U9467 (N_9467,N_9265,N_9351);
or U9468 (N_9468,N_9209,N_9269);
and U9469 (N_9469,N_9387,N_9290);
xor U9470 (N_9470,N_9260,N_9234);
nor U9471 (N_9471,N_9232,N_9289);
nor U9472 (N_9472,N_9204,N_9343);
or U9473 (N_9473,N_9280,N_9261);
and U9474 (N_9474,N_9362,N_9241);
nand U9475 (N_9475,N_9315,N_9354);
or U9476 (N_9476,N_9372,N_9225);
and U9477 (N_9477,N_9320,N_9252);
nand U9478 (N_9478,N_9267,N_9337);
nor U9479 (N_9479,N_9376,N_9201);
nor U9480 (N_9480,N_9363,N_9271);
xnor U9481 (N_9481,N_9365,N_9356);
and U9482 (N_9482,N_9299,N_9344);
nor U9483 (N_9483,N_9210,N_9207);
nand U9484 (N_9484,N_9383,N_9228);
nor U9485 (N_9485,N_9352,N_9206);
or U9486 (N_9486,N_9382,N_9246);
or U9487 (N_9487,N_9236,N_9342);
and U9488 (N_9488,N_9233,N_9240);
or U9489 (N_9489,N_9216,N_9238);
nand U9490 (N_9490,N_9219,N_9307);
or U9491 (N_9491,N_9328,N_9227);
xor U9492 (N_9492,N_9318,N_9231);
xnor U9493 (N_9493,N_9248,N_9214);
nor U9494 (N_9494,N_9262,N_9208);
nand U9495 (N_9495,N_9368,N_9380);
nor U9496 (N_9496,N_9292,N_9223);
and U9497 (N_9497,N_9359,N_9386);
nor U9498 (N_9498,N_9390,N_9244);
nor U9499 (N_9499,N_9369,N_9300);
or U9500 (N_9500,N_9239,N_9266);
nor U9501 (N_9501,N_9294,N_9326);
nor U9502 (N_9502,N_9215,N_9282);
or U9503 (N_9503,N_9230,N_9247);
xor U9504 (N_9504,N_9338,N_9257);
or U9505 (N_9505,N_9249,N_9227);
xnor U9506 (N_9506,N_9262,N_9225);
nor U9507 (N_9507,N_9294,N_9332);
nand U9508 (N_9508,N_9341,N_9363);
nand U9509 (N_9509,N_9312,N_9280);
xor U9510 (N_9510,N_9274,N_9366);
and U9511 (N_9511,N_9300,N_9296);
or U9512 (N_9512,N_9306,N_9386);
nor U9513 (N_9513,N_9331,N_9378);
or U9514 (N_9514,N_9288,N_9368);
or U9515 (N_9515,N_9310,N_9206);
nand U9516 (N_9516,N_9207,N_9322);
nand U9517 (N_9517,N_9387,N_9252);
or U9518 (N_9518,N_9261,N_9277);
nand U9519 (N_9519,N_9220,N_9232);
or U9520 (N_9520,N_9385,N_9299);
nand U9521 (N_9521,N_9201,N_9312);
nand U9522 (N_9522,N_9249,N_9337);
and U9523 (N_9523,N_9214,N_9342);
or U9524 (N_9524,N_9275,N_9331);
xor U9525 (N_9525,N_9363,N_9371);
and U9526 (N_9526,N_9218,N_9314);
and U9527 (N_9527,N_9201,N_9316);
or U9528 (N_9528,N_9369,N_9307);
nor U9529 (N_9529,N_9206,N_9356);
or U9530 (N_9530,N_9296,N_9225);
nand U9531 (N_9531,N_9223,N_9255);
nor U9532 (N_9532,N_9263,N_9278);
nand U9533 (N_9533,N_9251,N_9241);
nor U9534 (N_9534,N_9250,N_9243);
nand U9535 (N_9535,N_9308,N_9294);
or U9536 (N_9536,N_9349,N_9384);
or U9537 (N_9537,N_9235,N_9302);
nor U9538 (N_9538,N_9315,N_9394);
or U9539 (N_9539,N_9215,N_9251);
or U9540 (N_9540,N_9396,N_9310);
xor U9541 (N_9541,N_9344,N_9249);
nor U9542 (N_9542,N_9371,N_9206);
nor U9543 (N_9543,N_9341,N_9290);
xnor U9544 (N_9544,N_9367,N_9360);
nand U9545 (N_9545,N_9216,N_9208);
or U9546 (N_9546,N_9361,N_9393);
or U9547 (N_9547,N_9321,N_9275);
xnor U9548 (N_9548,N_9347,N_9320);
and U9549 (N_9549,N_9342,N_9232);
and U9550 (N_9550,N_9231,N_9345);
and U9551 (N_9551,N_9341,N_9307);
nand U9552 (N_9552,N_9219,N_9256);
nor U9553 (N_9553,N_9355,N_9311);
or U9554 (N_9554,N_9312,N_9366);
or U9555 (N_9555,N_9281,N_9227);
xnor U9556 (N_9556,N_9330,N_9212);
xnor U9557 (N_9557,N_9205,N_9288);
and U9558 (N_9558,N_9256,N_9382);
xor U9559 (N_9559,N_9370,N_9214);
nor U9560 (N_9560,N_9362,N_9204);
nand U9561 (N_9561,N_9213,N_9293);
nand U9562 (N_9562,N_9298,N_9272);
xor U9563 (N_9563,N_9370,N_9229);
or U9564 (N_9564,N_9356,N_9304);
or U9565 (N_9565,N_9289,N_9383);
or U9566 (N_9566,N_9350,N_9295);
and U9567 (N_9567,N_9340,N_9396);
xnor U9568 (N_9568,N_9329,N_9351);
nor U9569 (N_9569,N_9312,N_9325);
xnor U9570 (N_9570,N_9237,N_9324);
and U9571 (N_9571,N_9215,N_9264);
xnor U9572 (N_9572,N_9309,N_9213);
or U9573 (N_9573,N_9243,N_9343);
or U9574 (N_9574,N_9214,N_9383);
nand U9575 (N_9575,N_9337,N_9259);
nand U9576 (N_9576,N_9333,N_9359);
or U9577 (N_9577,N_9361,N_9301);
nor U9578 (N_9578,N_9380,N_9263);
xnor U9579 (N_9579,N_9335,N_9291);
nand U9580 (N_9580,N_9363,N_9359);
nand U9581 (N_9581,N_9317,N_9267);
nor U9582 (N_9582,N_9278,N_9253);
nor U9583 (N_9583,N_9353,N_9365);
and U9584 (N_9584,N_9369,N_9219);
or U9585 (N_9585,N_9276,N_9220);
xor U9586 (N_9586,N_9220,N_9237);
or U9587 (N_9587,N_9225,N_9351);
nor U9588 (N_9588,N_9243,N_9302);
xnor U9589 (N_9589,N_9314,N_9224);
and U9590 (N_9590,N_9347,N_9327);
or U9591 (N_9591,N_9316,N_9351);
nor U9592 (N_9592,N_9223,N_9215);
xor U9593 (N_9593,N_9257,N_9380);
and U9594 (N_9594,N_9241,N_9204);
and U9595 (N_9595,N_9237,N_9221);
nand U9596 (N_9596,N_9326,N_9315);
or U9597 (N_9597,N_9253,N_9334);
nand U9598 (N_9598,N_9337,N_9231);
nor U9599 (N_9599,N_9247,N_9265);
and U9600 (N_9600,N_9574,N_9496);
nor U9601 (N_9601,N_9507,N_9582);
or U9602 (N_9602,N_9588,N_9467);
xor U9603 (N_9603,N_9413,N_9476);
nor U9604 (N_9604,N_9552,N_9445);
and U9605 (N_9605,N_9428,N_9514);
nand U9606 (N_9606,N_9484,N_9433);
xor U9607 (N_9607,N_9500,N_9576);
or U9608 (N_9608,N_9418,N_9411);
or U9609 (N_9609,N_9403,N_9563);
nor U9610 (N_9610,N_9446,N_9452);
and U9611 (N_9611,N_9480,N_9422);
and U9612 (N_9612,N_9530,N_9572);
nor U9613 (N_9613,N_9498,N_9473);
xnor U9614 (N_9614,N_9585,N_9518);
xor U9615 (N_9615,N_9577,N_9405);
and U9616 (N_9616,N_9432,N_9584);
or U9617 (N_9617,N_9482,N_9559);
xnor U9618 (N_9618,N_9583,N_9575);
nor U9619 (N_9619,N_9503,N_9523);
or U9620 (N_9620,N_9497,N_9560);
nor U9621 (N_9621,N_9420,N_9404);
and U9622 (N_9622,N_9591,N_9434);
nand U9623 (N_9623,N_9407,N_9542);
nor U9624 (N_9624,N_9531,N_9548);
nand U9625 (N_9625,N_9544,N_9550);
nor U9626 (N_9626,N_9412,N_9541);
nand U9627 (N_9627,N_9400,N_9495);
nand U9628 (N_9628,N_9479,N_9491);
and U9629 (N_9629,N_9557,N_9421);
xnor U9630 (N_9630,N_9545,N_9468);
nor U9631 (N_9631,N_9546,N_9455);
nor U9632 (N_9632,N_9490,N_9424);
or U9633 (N_9633,N_9513,N_9538);
xor U9634 (N_9634,N_9558,N_9586);
or U9635 (N_9635,N_9595,N_9556);
nor U9636 (N_9636,N_9508,N_9458);
xor U9637 (N_9637,N_9554,N_9539);
and U9638 (N_9638,N_9505,N_9449);
and U9639 (N_9639,N_9415,N_9435);
nand U9640 (N_9640,N_9549,N_9506);
and U9641 (N_9641,N_9528,N_9442);
and U9642 (N_9642,N_9457,N_9517);
nand U9643 (N_9643,N_9440,N_9511);
and U9644 (N_9644,N_9562,N_9551);
xnor U9645 (N_9645,N_9499,N_9555);
or U9646 (N_9646,N_9561,N_9537);
nor U9647 (N_9647,N_9589,N_9571);
nor U9648 (N_9648,N_9597,N_9483);
nor U9649 (N_9649,N_9447,N_9454);
nand U9650 (N_9650,N_9520,N_9451);
xor U9651 (N_9651,N_9522,N_9533);
nor U9652 (N_9652,N_9580,N_9478);
or U9653 (N_9653,N_9450,N_9419);
or U9654 (N_9654,N_9475,N_9504);
or U9655 (N_9655,N_9417,N_9466);
nand U9656 (N_9656,N_9540,N_9423);
xor U9657 (N_9657,N_9462,N_9485);
and U9658 (N_9658,N_9566,N_9578);
nor U9659 (N_9659,N_9526,N_9427);
and U9660 (N_9660,N_9521,N_9524);
nand U9661 (N_9661,N_9567,N_9568);
and U9662 (N_9662,N_9470,N_9408);
nand U9663 (N_9663,N_9543,N_9444);
and U9664 (N_9664,N_9494,N_9509);
xor U9665 (N_9665,N_9515,N_9453);
and U9666 (N_9666,N_9430,N_9459);
and U9667 (N_9667,N_9471,N_9535);
nor U9668 (N_9668,N_9464,N_9488);
and U9669 (N_9669,N_9599,N_9465);
xor U9670 (N_9670,N_9426,N_9431);
nand U9671 (N_9671,N_9501,N_9410);
nor U9672 (N_9672,N_9487,N_9416);
or U9673 (N_9673,N_9493,N_9463);
xnor U9674 (N_9674,N_9414,N_9598);
nand U9675 (N_9675,N_9443,N_9469);
or U9676 (N_9676,N_9460,N_9581);
nand U9677 (N_9677,N_9579,N_9510);
or U9678 (N_9678,N_9402,N_9486);
nor U9679 (N_9679,N_9553,N_9570);
xor U9680 (N_9680,N_9564,N_9519);
xnor U9681 (N_9681,N_9472,N_9587);
or U9682 (N_9682,N_9448,N_9547);
or U9683 (N_9683,N_9401,N_9527);
and U9684 (N_9684,N_9437,N_9436);
xor U9685 (N_9685,N_9461,N_9439);
nand U9686 (N_9686,N_9532,N_9406);
nor U9687 (N_9687,N_9596,N_9456);
nor U9688 (N_9688,N_9536,N_9573);
xor U9689 (N_9689,N_9512,N_9429);
and U9690 (N_9690,N_9438,N_9425);
nand U9691 (N_9691,N_9502,N_9594);
xnor U9692 (N_9692,N_9409,N_9474);
nor U9693 (N_9693,N_9489,N_9492);
or U9694 (N_9694,N_9516,N_9593);
and U9695 (N_9695,N_9529,N_9534);
nor U9696 (N_9696,N_9592,N_9441);
and U9697 (N_9697,N_9525,N_9481);
nor U9698 (N_9698,N_9565,N_9590);
or U9699 (N_9699,N_9477,N_9569);
nand U9700 (N_9700,N_9587,N_9482);
or U9701 (N_9701,N_9435,N_9560);
nand U9702 (N_9702,N_9404,N_9406);
and U9703 (N_9703,N_9526,N_9575);
xnor U9704 (N_9704,N_9590,N_9429);
and U9705 (N_9705,N_9478,N_9432);
nand U9706 (N_9706,N_9559,N_9512);
nand U9707 (N_9707,N_9508,N_9449);
or U9708 (N_9708,N_9496,N_9434);
and U9709 (N_9709,N_9430,N_9576);
nor U9710 (N_9710,N_9497,N_9583);
nand U9711 (N_9711,N_9512,N_9552);
nand U9712 (N_9712,N_9511,N_9592);
nand U9713 (N_9713,N_9516,N_9552);
nand U9714 (N_9714,N_9489,N_9465);
nand U9715 (N_9715,N_9472,N_9526);
or U9716 (N_9716,N_9555,N_9447);
nor U9717 (N_9717,N_9407,N_9432);
nand U9718 (N_9718,N_9573,N_9493);
nor U9719 (N_9719,N_9400,N_9444);
xor U9720 (N_9720,N_9459,N_9478);
nor U9721 (N_9721,N_9452,N_9548);
xor U9722 (N_9722,N_9483,N_9431);
or U9723 (N_9723,N_9522,N_9549);
nor U9724 (N_9724,N_9420,N_9513);
and U9725 (N_9725,N_9419,N_9568);
and U9726 (N_9726,N_9407,N_9523);
nand U9727 (N_9727,N_9585,N_9457);
or U9728 (N_9728,N_9424,N_9445);
xnor U9729 (N_9729,N_9401,N_9498);
xor U9730 (N_9730,N_9533,N_9447);
and U9731 (N_9731,N_9475,N_9527);
nand U9732 (N_9732,N_9454,N_9450);
and U9733 (N_9733,N_9432,N_9518);
and U9734 (N_9734,N_9516,N_9527);
or U9735 (N_9735,N_9536,N_9497);
xnor U9736 (N_9736,N_9473,N_9507);
and U9737 (N_9737,N_9555,N_9524);
nand U9738 (N_9738,N_9594,N_9486);
xor U9739 (N_9739,N_9547,N_9437);
and U9740 (N_9740,N_9481,N_9498);
or U9741 (N_9741,N_9424,N_9517);
or U9742 (N_9742,N_9443,N_9446);
nor U9743 (N_9743,N_9576,N_9543);
nor U9744 (N_9744,N_9471,N_9534);
and U9745 (N_9745,N_9489,N_9441);
or U9746 (N_9746,N_9567,N_9500);
nand U9747 (N_9747,N_9500,N_9583);
nor U9748 (N_9748,N_9588,N_9530);
or U9749 (N_9749,N_9430,N_9547);
nand U9750 (N_9750,N_9421,N_9563);
xnor U9751 (N_9751,N_9525,N_9479);
and U9752 (N_9752,N_9454,N_9501);
and U9753 (N_9753,N_9494,N_9529);
nor U9754 (N_9754,N_9445,N_9461);
nand U9755 (N_9755,N_9479,N_9401);
or U9756 (N_9756,N_9576,N_9518);
or U9757 (N_9757,N_9516,N_9483);
xnor U9758 (N_9758,N_9479,N_9538);
and U9759 (N_9759,N_9412,N_9573);
or U9760 (N_9760,N_9449,N_9458);
and U9761 (N_9761,N_9455,N_9516);
nor U9762 (N_9762,N_9509,N_9577);
or U9763 (N_9763,N_9488,N_9521);
nor U9764 (N_9764,N_9563,N_9497);
and U9765 (N_9765,N_9466,N_9438);
nand U9766 (N_9766,N_9476,N_9472);
nand U9767 (N_9767,N_9552,N_9547);
or U9768 (N_9768,N_9417,N_9416);
or U9769 (N_9769,N_9571,N_9446);
nand U9770 (N_9770,N_9556,N_9515);
xnor U9771 (N_9771,N_9508,N_9445);
xor U9772 (N_9772,N_9442,N_9431);
or U9773 (N_9773,N_9503,N_9418);
or U9774 (N_9774,N_9423,N_9422);
and U9775 (N_9775,N_9532,N_9405);
and U9776 (N_9776,N_9568,N_9528);
nor U9777 (N_9777,N_9420,N_9563);
xnor U9778 (N_9778,N_9583,N_9421);
xor U9779 (N_9779,N_9581,N_9526);
or U9780 (N_9780,N_9570,N_9407);
xor U9781 (N_9781,N_9564,N_9586);
nor U9782 (N_9782,N_9551,N_9430);
nand U9783 (N_9783,N_9400,N_9587);
nor U9784 (N_9784,N_9568,N_9509);
and U9785 (N_9785,N_9572,N_9435);
or U9786 (N_9786,N_9568,N_9478);
and U9787 (N_9787,N_9477,N_9408);
xor U9788 (N_9788,N_9461,N_9591);
nand U9789 (N_9789,N_9455,N_9522);
nor U9790 (N_9790,N_9439,N_9483);
or U9791 (N_9791,N_9426,N_9596);
or U9792 (N_9792,N_9522,N_9504);
xor U9793 (N_9793,N_9595,N_9590);
nand U9794 (N_9794,N_9441,N_9572);
and U9795 (N_9795,N_9442,N_9510);
and U9796 (N_9796,N_9489,N_9554);
or U9797 (N_9797,N_9563,N_9502);
xnor U9798 (N_9798,N_9573,N_9571);
xnor U9799 (N_9799,N_9560,N_9566);
nand U9800 (N_9800,N_9618,N_9656);
xor U9801 (N_9801,N_9641,N_9620);
nand U9802 (N_9802,N_9676,N_9781);
or U9803 (N_9803,N_9717,N_9737);
and U9804 (N_9804,N_9790,N_9750);
and U9805 (N_9805,N_9740,N_9606);
xor U9806 (N_9806,N_9665,N_9742);
nand U9807 (N_9807,N_9622,N_9602);
xor U9808 (N_9808,N_9664,N_9733);
or U9809 (N_9809,N_9673,N_9772);
nor U9810 (N_9810,N_9741,N_9659);
or U9811 (N_9811,N_9612,N_9732);
or U9812 (N_9812,N_9768,N_9736);
or U9813 (N_9813,N_9642,N_9639);
or U9814 (N_9814,N_9766,N_9777);
or U9815 (N_9815,N_9713,N_9670);
nor U9816 (N_9816,N_9690,N_9650);
nor U9817 (N_9817,N_9702,N_9675);
or U9818 (N_9818,N_9603,N_9645);
xnor U9819 (N_9819,N_9720,N_9681);
or U9820 (N_9820,N_9700,N_9655);
and U9821 (N_9821,N_9685,N_9696);
or U9822 (N_9822,N_9704,N_9738);
xnor U9823 (N_9823,N_9794,N_9661);
xor U9824 (N_9824,N_9625,N_9747);
xnor U9825 (N_9825,N_9752,N_9744);
nand U9826 (N_9826,N_9629,N_9626);
xnor U9827 (N_9827,N_9708,N_9695);
or U9828 (N_9828,N_9701,N_9743);
or U9829 (N_9829,N_9709,N_9692);
or U9830 (N_9830,N_9764,N_9698);
nand U9831 (N_9831,N_9771,N_9746);
xor U9832 (N_9832,N_9632,N_9760);
nor U9833 (N_9833,N_9705,N_9666);
nor U9834 (N_9834,N_9761,N_9795);
and U9835 (N_9835,N_9782,N_9725);
or U9836 (N_9836,N_9763,N_9784);
xnor U9837 (N_9837,N_9694,N_9667);
and U9838 (N_9838,N_9652,N_9686);
and U9839 (N_9839,N_9614,N_9778);
nor U9840 (N_9840,N_9636,N_9793);
nand U9841 (N_9841,N_9789,N_9633);
or U9842 (N_9842,N_9723,N_9726);
and U9843 (N_9843,N_9788,N_9785);
xor U9844 (N_9844,N_9730,N_9697);
xor U9845 (N_9845,N_9658,N_9683);
and U9846 (N_9846,N_9631,N_9699);
or U9847 (N_9847,N_9647,N_9796);
nand U9848 (N_9848,N_9677,N_9649);
xnor U9849 (N_9849,N_9621,N_9765);
nand U9850 (N_9850,N_9753,N_9689);
nand U9851 (N_9851,N_9775,N_9751);
nor U9852 (N_9852,N_9748,N_9729);
or U9853 (N_9853,N_9734,N_9791);
or U9854 (N_9854,N_9786,N_9706);
nand U9855 (N_9855,N_9654,N_9638);
and U9856 (N_9856,N_9616,N_9783);
nor U9857 (N_9857,N_9711,N_9703);
and U9858 (N_9858,N_9773,N_9787);
or U9859 (N_9859,N_9610,N_9608);
and U9860 (N_9860,N_9719,N_9617);
nand U9861 (N_9861,N_9756,N_9600);
and U9862 (N_9862,N_9635,N_9798);
nand U9863 (N_9863,N_9669,N_9774);
and U9864 (N_9864,N_9758,N_9628);
and U9865 (N_9865,N_9714,N_9668);
nor U9866 (N_9866,N_9780,N_9797);
or U9867 (N_9867,N_9731,N_9754);
nand U9868 (N_9868,N_9678,N_9615);
and U9869 (N_9869,N_9671,N_9682);
and U9870 (N_9870,N_9646,N_9674);
nand U9871 (N_9871,N_9757,N_9634);
nor U9872 (N_9872,N_9770,N_9607);
and U9873 (N_9873,N_9707,N_9718);
nand U9874 (N_9874,N_9779,N_9662);
or U9875 (N_9875,N_9637,N_9688);
or U9876 (N_9876,N_9749,N_9693);
or U9877 (N_9877,N_9759,N_9648);
nand U9878 (N_9878,N_9716,N_9609);
or U9879 (N_9879,N_9611,N_9660);
or U9880 (N_9880,N_9684,N_9644);
and U9881 (N_9881,N_9767,N_9613);
and U9882 (N_9882,N_9679,N_9722);
nand U9883 (N_9883,N_9601,N_9630);
nand U9884 (N_9884,N_9710,N_9672);
nor U9885 (N_9885,N_9712,N_9640);
nor U9886 (N_9886,N_9745,N_9755);
or U9887 (N_9887,N_9627,N_9799);
nand U9888 (N_9888,N_9653,N_9715);
nor U9889 (N_9889,N_9739,N_9651);
nor U9890 (N_9890,N_9643,N_9605);
or U9891 (N_9891,N_9680,N_9735);
nor U9892 (N_9892,N_9691,N_9619);
nor U9893 (N_9893,N_9663,N_9721);
nor U9894 (N_9894,N_9604,N_9769);
xnor U9895 (N_9895,N_9657,N_9724);
nand U9896 (N_9896,N_9762,N_9623);
xor U9897 (N_9897,N_9728,N_9792);
xnor U9898 (N_9898,N_9624,N_9687);
or U9899 (N_9899,N_9776,N_9727);
nand U9900 (N_9900,N_9605,N_9655);
nand U9901 (N_9901,N_9696,N_9720);
or U9902 (N_9902,N_9709,N_9644);
or U9903 (N_9903,N_9605,N_9624);
xnor U9904 (N_9904,N_9661,N_9705);
nand U9905 (N_9905,N_9793,N_9732);
nand U9906 (N_9906,N_9652,N_9743);
nor U9907 (N_9907,N_9702,N_9776);
nor U9908 (N_9908,N_9735,N_9702);
nand U9909 (N_9909,N_9708,N_9794);
or U9910 (N_9910,N_9656,N_9722);
or U9911 (N_9911,N_9772,N_9625);
or U9912 (N_9912,N_9651,N_9639);
nand U9913 (N_9913,N_9712,N_9618);
and U9914 (N_9914,N_9663,N_9770);
nor U9915 (N_9915,N_9735,N_9714);
xnor U9916 (N_9916,N_9736,N_9778);
xnor U9917 (N_9917,N_9696,N_9688);
and U9918 (N_9918,N_9715,N_9667);
and U9919 (N_9919,N_9631,N_9700);
nor U9920 (N_9920,N_9763,N_9671);
or U9921 (N_9921,N_9649,N_9627);
nor U9922 (N_9922,N_9704,N_9646);
nand U9923 (N_9923,N_9642,N_9635);
and U9924 (N_9924,N_9658,N_9609);
and U9925 (N_9925,N_9625,N_9780);
xor U9926 (N_9926,N_9697,N_9631);
nor U9927 (N_9927,N_9673,N_9791);
nand U9928 (N_9928,N_9792,N_9738);
or U9929 (N_9929,N_9678,N_9776);
nor U9930 (N_9930,N_9645,N_9705);
nand U9931 (N_9931,N_9636,N_9785);
or U9932 (N_9932,N_9690,N_9662);
xor U9933 (N_9933,N_9781,N_9777);
xnor U9934 (N_9934,N_9767,N_9751);
nor U9935 (N_9935,N_9611,N_9792);
nand U9936 (N_9936,N_9663,N_9753);
xnor U9937 (N_9937,N_9778,N_9715);
or U9938 (N_9938,N_9714,N_9780);
and U9939 (N_9939,N_9642,N_9786);
and U9940 (N_9940,N_9788,N_9735);
nand U9941 (N_9941,N_9699,N_9673);
or U9942 (N_9942,N_9777,N_9618);
and U9943 (N_9943,N_9713,N_9789);
or U9944 (N_9944,N_9758,N_9715);
or U9945 (N_9945,N_9713,N_9734);
or U9946 (N_9946,N_9707,N_9688);
nand U9947 (N_9947,N_9786,N_9773);
and U9948 (N_9948,N_9782,N_9690);
or U9949 (N_9949,N_9628,N_9616);
nand U9950 (N_9950,N_9674,N_9767);
nor U9951 (N_9951,N_9694,N_9662);
or U9952 (N_9952,N_9739,N_9787);
nor U9953 (N_9953,N_9759,N_9674);
xnor U9954 (N_9954,N_9670,N_9655);
xor U9955 (N_9955,N_9732,N_9644);
xnor U9956 (N_9956,N_9783,N_9730);
nand U9957 (N_9957,N_9682,N_9779);
nor U9958 (N_9958,N_9764,N_9635);
and U9959 (N_9959,N_9603,N_9630);
or U9960 (N_9960,N_9622,N_9623);
nand U9961 (N_9961,N_9776,N_9650);
nor U9962 (N_9962,N_9776,N_9604);
nand U9963 (N_9963,N_9655,N_9759);
and U9964 (N_9964,N_9612,N_9747);
and U9965 (N_9965,N_9769,N_9787);
nor U9966 (N_9966,N_9749,N_9627);
nand U9967 (N_9967,N_9634,N_9637);
and U9968 (N_9968,N_9652,N_9723);
nor U9969 (N_9969,N_9771,N_9737);
and U9970 (N_9970,N_9738,N_9700);
xnor U9971 (N_9971,N_9639,N_9762);
and U9972 (N_9972,N_9775,N_9764);
nand U9973 (N_9973,N_9633,N_9702);
nor U9974 (N_9974,N_9610,N_9725);
or U9975 (N_9975,N_9760,N_9620);
nand U9976 (N_9976,N_9716,N_9734);
or U9977 (N_9977,N_9653,N_9670);
nand U9978 (N_9978,N_9763,N_9755);
nand U9979 (N_9979,N_9719,N_9671);
or U9980 (N_9980,N_9778,N_9683);
xor U9981 (N_9981,N_9698,N_9743);
xor U9982 (N_9982,N_9776,N_9744);
nor U9983 (N_9983,N_9719,N_9612);
and U9984 (N_9984,N_9642,N_9648);
or U9985 (N_9985,N_9660,N_9750);
xor U9986 (N_9986,N_9763,N_9722);
nor U9987 (N_9987,N_9793,N_9638);
nand U9988 (N_9988,N_9682,N_9792);
nor U9989 (N_9989,N_9666,N_9702);
or U9990 (N_9990,N_9620,N_9627);
or U9991 (N_9991,N_9645,N_9789);
and U9992 (N_9992,N_9653,N_9786);
or U9993 (N_9993,N_9748,N_9666);
or U9994 (N_9994,N_9601,N_9767);
or U9995 (N_9995,N_9731,N_9709);
nand U9996 (N_9996,N_9789,N_9625);
nor U9997 (N_9997,N_9628,N_9605);
xor U9998 (N_9998,N_9691,N_9659);
and U9999 (N_9999,N_9711,N_9715);
nand U10000 (N_10000,N_9939,N_9902);
nand U10001 (N_10001,N_9967,N_9908);
nand U10002 (N_10002,N_9837,N_9951);
xnor U10003 (N_10003,N_9913,N_9845);
xnor U10004 (N_10004,N_9835,N_9952);
nand U10005 (N_10005,N_9928,N_9893);
xor U10006 (N_10006,N_9876,N_9839);
or U10007 (N_10007,N_9915,N_9982);
xor U10008 (N_10008,N_9812,N_9936);
nor U10009 (N_10009,N_9820,N_9852);
and U10010 (N_10010,N_9833,N_9881);
or U10011 (N_10011,N_9977,N_9957);
or U10012 (N_10012,N_9942,N_9965);
nor U10013 (N_10013,N_9922,N_9879);
nand U10014 (N_10014,N_9849,N_9905);
and U10015 (N_10015,N_9918,N_9943);
xnor U10016 (N_10016,N_9920,N_9818);
and U10017 (N_10017,N_9948,N_9838);
xnor U10018 (N_10018,N_9828,N_9972);
or U10019 (N_10019,N_9978,N_9896);
and U10020 (N_10020,N_9937,N_9958);
and U10021 (N_10021,N_9945,N_9926);
xor U10022 (N_10022,N_9996,N_9816);
and U10023 (N_10023,N_9925,N_9955);
nor U10024 (N_10024,N_9840,N_9865);
nor U10025 (N_10025,N_9904,N_9993);
xnor U10026 (N_10026,N_9981,N_9882);
and U10027 (N_10027,N_9826,N_9931);
and U10028 (N_10028,N_9997,N_9813);
and U10029 (N_10029,N_9850,N_9827);
or U10030 (N_10030,N_9853,N_9964);
xor U10031 (N_10031,N_9807,N_9864);
xnor U10032 (N_10032,N_9974,N_9877);
and U10033 (N_10033,N_9801,N_9821);
nand U10034 (N_10034,N_9927,N_9988);
or U10035 (N_10035,N_9987,N_9971);
or U10036 (N_10036,N_9829,N_9874);
xor U10037 (N_10037,N_9998,N_9909);
and U10038 (N_10038,N_9891,N_9995);
nor U10039 (N_10039,N_9805,N_9851);
and U10040 (N_10040,N_9985,N_9941);
nor U10041 (N_10041,N_9836,N_9970);
nand U10042 (N_10042,N_9935,N_9871);
and U10043 (N_10043,N_9857,N_9932);
or U10044 (N_10044,N_9856,N_9832);
nor U10045 (N_10045,N_9815,N_9802);
nand U10046 (N_10046,N_9878,N_9953);
xnor U10047 (N_10047,N_9898,N_9809);
nor U10048 (N_10048,N_9870,N_9804);
or U10049 (N_10049,N_9841,N_9983);
nand U10050 (N_10050,N_9961,N_9884);
or U10051 (N_10051,N_9938,N_9875);
and U10052 (N_10052,N_9914,N_9994);
xnor U10053 (N_10053,N_9800,N_9854);
nor U10054 (N_10054,N_9962,N_9886);
xnor U10055 (N_10055,N_9861,N_9947);
and U10056 (N_10056,N_9989,N_9923);
nand U10057 (N_10057,N_9901,N_9842);
nand U10058 (N_10058,N_9917,N_9859);
xnor U10059 (N_10059,N_9959,N_9895);
nor U10060 (N_10060,N_9810,N_9900);
nor U10061 (N_10061,N_9944,N_9903);
or U10062 (N_10062,N_9949,N_9868);
and U10063 (N_10063,N_9986,N_9890);
or U10064 (N_10064,N_9894,N_9883);
nand U10065 (N_10065,N_9855,N_9831);
nor U10066 (N_10066,N_9808,N_9806);
xnor U10067 (N_10067,N_9858,N_9966);
or U10068 (N_10068,N_9814,N_9824);
or U10069 (N_10069,N_9906,N_9968);
xor U10070 (N_10070,N_9863,N_9822);
or U10071 (N_10071,N_9990,N_9975);
or U10072 (N_10072,N_9888,N_9892);
nand U10073 (N_10073,N_9817,N_9979);
and U10074 (N_10074,N_9811,N_9873);
or U10075 (N_10075,N_9991,N_9934);
and U10076 (N_10076,N_9999,N_9897);
nand U10077 (N_10077,N_9956,N_9919);
xor U10078 (N_10078,N_9963,N_9969);
or U10079 (N_10079,N_9946,N_9819);
nand U10080 (N_10080,N_9930,N_9848);
xor U10081 (N_10081,N_9933,N_9803);
nand U10082 (N_10082,N_9844,N_9867);
nor U10083 (N_10083,N_9976,N_9834);
nand U10084 (N_10084,N_9887,N_9924);
nand U10085 (N_10085,N_9911,N_9973);
and U10086 (N_10086,N_9899,N_9992);
or U10087 (N_10087,N_9912,N_9960);
or U10088 (N_10088,N_9869,N_9872);
nand U10089 (N_10089,N_9823,N_9954);
or U10090 (N_10090,N_9916,N_9889);
xnor U10091 (N_10091,N_9940,N_9846);
nand U10092 (N_10092,N_9866,N_9910);
nand U10093 (N_10093,N_9980,N_9862);
xor U10094 (N_10094,N_9843,N_9907);
nor U10095 (N_10095,N_9880,N_9830);
or U10096 (N_10096,N_9929,N_9847);
nand U10097 (N_10097,N_9984,N_9921);
nor U10098 (N_10098,N_9825,N_9885);
nand U10099 (N_10099,N_9950,N_9860);
xor U10100 (N_10100,N_9828,N_9832);
xor U10101 (N_10101,N_9856,N_9819);
or U10102 (N_10102,N_9846,N_9931);
nor U10103 (N_10103,N_9910,N_9953);
nand U10104 (N_10104,N_9829,N_9803);
xor U10105 (N_10105,N_9960,N_9972);
and U10106 (N_10106,N_9923,N_9835);
and U10107 (N_10107,N_9943,N_9868);
or U10108 (N_10108,N_9812,N_9895);
nand U10109 (N_10109,N_9907,N_9852);
xor U10110 (N_10110,N_9801,N_9958);
and U10111 (N_10111,N_9897,N_9914);
nand U10112 (N_10112,N_9853,N_9967);
nand U10113 (N_10113,N_9951,N_9890);
nand U10114 (N_10114,N_9998,N_9858);
or U10115 (N_10115,N_9887,N_9922);
nor U10116 (N_10116,N_9939,N_9940);
xor U10117 (N_10117,N_9895,N_9983);
xnor U10118 (N_10118,N_9801,N_9974);
xor U10119 (N_10119,N_9824,N_9810);
nand U10120 (N_10120,N_9974,N_9800);
nand U10121 (N_10121,N_9894,N_9971);
nand U10122 (N_10122,N_9886,N_9848);
and U10123 (N_10123,N_9947,N_9820);
and U10124 (N_10124,N_9990,N_9903);
nor U10125 (N_10125,N_9868,N_9984);
nand U10126 (N_10126,N_9834,N_9926);
and U10127 (N_10127,N_9883,N_9979);
or U10128 (N_10128,N_9830,N_9919);
or U10129 (N_10129,N_9893,N_9926);
nand U10130 (N_10130,N_9857,N_9846);
xnor U10131 (N_10131,N_9945,N_9943);
and U10132 (N_10132,N_9822,N_9803);
and U10133 (N_10133,N_9872,N_9913);
nor U10134 (N_10134,N_9868,N_9824);
and U10135 (N_10135,N_9800,N_9941);
nand U10136 (N_10136,N_9937,N_9922);
and U10137 (N_10137,N_9969,N_9936);
nand U10138 (N_10138,N_9954,N_9991);
or U10139 (N_10139,N_9946,N_9873);
nor U10140 (N_10140,N_9816,N_9850);
nand U10141 (N_10141,N_9906,N_9931);
and U10142 (N_10142,N_9826,N_9880);
nand U10143 (N_10143,N_9929,N_9972);
nand U10144 (N_10144,N_9881,N_9951);
nor U10145 (N_10145,N_9921,N_9987);
nor U10146 (N_10146,N_9844,N_9818);
and U10147 (N_10147,N_9967,N_9930);
nor U10148 (N_10148,N_9935,N_9868);
and U10149 (N_10149,N_9904,N_9879);
or U10150 (N_10150,N_9949,N_9834);
or U10151 (N_10151,N_9845,N_9998);
xnor U10152 (N_10152,N_9810,N_9953);
nand U10153 (N_10153,N_9931,N_9988);
or U10154 (N_10154,N_9958,N_9894);
nand U10155 (N_10155,N_9937,N_9858);
and U10156 (N_10156,N_9815,N_9935);
nand U10157 (N_10157,N_9909,N_9967);
nand U10158 (N_10158,N_9986,N_9835);
and U10159 (N_10159,N_9871,N_9843);
nor U10160 (N_10160,N_9962,N_9884);
xnor U10161 (N_10161,N_9841,N_9812);
xor U10162 (N_10162,N_9985,N_9846);
or U10163 (N_10163,N_9945,N_9800);
and U10164 (N_10164,N_9900,N_9814);
and U10165 (N_10165,N_9935,N_9840);
xor U10166 (N_10166,N_9986,N_9855);
nand U10167 (N_10167,N_9929,N_9927);
nor U10168 (N_10168,N_9973,N_9938);
or U10169 (N_10169,N_9964,N_9849);
or U10170 (N_10170,N_9960,N_9892);
xor U10171 (N_10171,N_9912,N_9829);
and U10172 (N_10172,N_9944,N_9868);
nor U10173 (N_10173,N_9866,N_9944);
and U10174 (N_10174,N_9859,N_9977);
nand U10175 (N_10175,N_9858,N_9923);
xnor U10176 (N_10176,N_9945,N_9989);
and U10177 (N_10177,N_9831,N_9973);
nand U10178 (N_10178,N_9868,N_9862);
xnor U10179 (N_10179,N_9873,N_9876);
nor U10180 (N_10180,N_9917,N_9922);
xor U10181 (N_10181,N_9821,N_9892);
or U10182 (N_10182,N_9807,N_9979);
nand U10183 (N_10183,N_9851,N_9923);
and U10184 (N_10184,N_9814,N_9802);
or U10185 (N_10185,N_9932,N_9978);
or U10186 (N_10186,N_9968,N_9816);
and U10187 (N_10187,N_9999,N_9802);
nand U10188 (N_10188,N_9917,N_9836);
or U10189 (N_10189,N_9940,N_9810);
xor U10190 (N_10190,N_9859,N_9918);
nand U10191 (N_10191,N_9894,N_9809);
xnor U10192 (N_10192,N_9823,N_9926);
or U10193 (N_10193,N_9963,N_9939);
nand U10194 (N_10194,N_9845,N_9951);
and U10195 (N_10195,N_9914,N_9917);
xnor U10196 (N_10196,N_9930,N_9886);
nand U10197 (N_10197,N_9807,N_9906);
or U10198 (N_10198,N_9982,N_9803);
nand U10199 (N_10199,N_9837,N_9859);
nor U10200 (N_10200,N_10010,N_10198);
and U10201 (N_10201,N_10091,N_10098);
xnor U10202 (N_10202,N_10104,N_10025);
nor U10203 (N_10203,N_10061,N_10177);
and U10204 (N_10204,N_10112,N_10037);
xnor U10205 (N_10205,N_10004,N_10014);
or U10206 (N_10206,N_10188,N_10175);
or U10207 (N_10207,N_10153,N_10065);
nor U10208 (N_10208,N_10088,N_10080);
or U10209 (N_10209,N_10149,N_10003);
nor U10210 (N_10210,N_10100,N_10064);
nand U10211 (N_10211,N_10157,N_10000);
and U10212 (N_10212,N_10108,N_10007);
or U10213 (N_10213,N_10047,N_10075);
nor U10214 (N_10214,N_10169,N_10039);
or U10215 (N_10215,N_10161,N_10148);
nor U10216 (N_10216,N_10070,N_10178);
or U10217 (N_10217,N_10027,N_10071);
and U10218 (N_10218,N_10019,N_10144);
and U10219 (N_10219,N_10170,N_10151);
or U10220 (N_10220,N_10183,N_10042);
and U10221 (N_10221,N_10165,N_10094);
or U10222 (N_10222,N_10097,N_10182);
nor U10223 (N_10223,N_10068,N_10032);
or U10224 (N_10224,N_10063,N_10073);
and U10225 (N_10225,N_10074,N_10180);
xnor U10226 (N_10226,N_10193,N_10185);
xor U10227 (N_10227,N_10168,N_10141);
and U10228 (N_10228,N_10124,N_10172);
nand U10229 (N_10229,N_10099,N_10067);
and U10230 (N_10230,N_10101,N_10048);
nor U10231 (N_10231,N_10125,N_10142);
and U10232 (N_10232,N_10166,N_10043);
nor U10233 (N_10233,N_10095,N_10044);
nand U10234 (N_10234,N_10111,N_10022);
and U10235 (N_10235,N_10085,N_10009);
xor U10236 (N_10236,N_10190,N_10053);
nand U10237 (N_10237,N_10143,N_10041);
nand U10238 (N_10238,N_10119,N_10107);
nand U10239 (N_10239,N_10150,N_10050);
nor U10240 (N_10240,N_10001,N_10158);
xor U10241 (N_10241,N_10139,N_10077);
and U10242 (N_10242,N_10028,N_10076);
nor U10243 (N_10243,N_10132,N_10059);
nor U10244 (N_10244,N_10136,N_10110);
and U10245 (N_10245,N_10083,N_10156);
xnor U10246 (N_10246,N_10194,N_10147);
xnor U10247 (N_10247,N_10018,N_10086);
and U10248 (N_10248,N_10121,N_10002);
and U10249 (N_10249,N_10049,N_10052);
or U10250 (N_10250,N_10105,N_10122);
xor U10251 (N_10251,N_10160,N_10033);
or U10252 (N_10252,N_10116,N_10102);
nand U10253 (N_10253,N_10024,N_10113);
or U10254 (N_10254,N_10045,N_10154);
nor U10255 (N_10255,N_10066,N_10195);
xor U10256 (N_10256,N_10056,N_10179);
nor U10257 (N_10257,N_10164,N_10159);
xnor U10258 (N_10258,N_10131,N_10118);
nand U10259 (N_10259,N_10181,N_10171);
xnor U10260 (N_10260,N_10079,N_10058);
nand U10261 (N_10261,N_10057,N_10031);
nor U10262 (N_10262,N_10012,N_10145);
nor U10263 (N_10263,N_10176,N_10084);
or U10264 (N_10264,N_10029,N_10146);
nor U10265 (N_10265,N_10026,N_10134);
xnor U10266 (N_10266,N_10103,N_10087);
nor U10267 (N_10267,N_10021,N_10138);
xor U10268 (N_10268,N_10152,N_10155);
and U10269 (N_10269,N_10006,N_10096);
nor U10270 (N_10270,N_10174,N_10192);
nand U10271 (N_10271,N_10186,N_10054);
nor U10272 (N_10272,N_10082,N_10081);
or U10273 (N_10273,N_10092,N_10008);
nor U10274 (N_10274,N_10187,N_10016);
nor U10275 (N_10275,N_10191,N_10051);
or U10276 (N_10276,N_10140,N_10015);
or U10277 (N_10277,N_10114,N_10013);
or U10278 (N_10278,N_10128,N_10196);
nor U10279 (N_10279,N_10120,N_10078);
or U10280 (N_10280,N_10035,N_10017);
nor U10281 (N_10281,N_10167,N_10127);
nand U10282 (N_10282,N_10005,N_10184);
nand U10283 (N_10283,N_10106,N_10023);
or U10284 (N_10284,N_10020,N_10197);
or U10285 (N_10285,N_10189,N_10046);
xnor U10286 (N_10286,N_10040,N_10126);
nor U10287 (N_10287,N_10090,N_10069);
and U10288 (N_10288,N_10133,N_10163);
nand U10289 (N_10289,N_10089,N_10199);
and U10290 (N_10290,N_10036,N_10135);
and U10291 (N_10291,N_10030,N_10137);
and U10292 (N_10292,N_10115,N_10060);
and U10293 (N_10293,N_10093,N_10055);
nand U10294 (N_10294,N_10129,N_10130);
nor U10295 (N_10295,N_10109,N_10123);
and U10296 (N_10296,N_10117,N_10072);
nand U10297 (N_10297,N_10162,N_10173);
or U10298 (N_10298,N_10011,N_10034);
or U10299 (N_10299,N_10038,N_10062);
nor U10300 (N_10300,N_10194,N_10000);
and U10301 (N_10301,N_10102,N_10115);
and U10302 (N_10302,N_10052,N_10061);
and U10303 (N_10303,N_10082,N_10175);
xor U10304 (N_10304,N_10173,N_10168);
xor U10305 (N_10305,N_10098,N_10042);
or U10306 (N_10306,N_10149,N_10189);
or U10307 (N_10307,N_10187,N_10035);
and U10308 (N_10308,N_10139,N_10174);
and U10309 (N_10309,N_10186,N_10014);
or U10310 (N_10310,N_10052,N_10019);
nor U10311 (N_10311,N_10134,N_10179);
and U10312 (N_10312,N_10128,N_10104);
nor U10313 (N_10313,N_10157,N_10067);
nand U10314 (N_10314,N_10189,N_10095);
xnor U10315 (N_10315,N_10126,N_10148);
or U10316 (N_10316,N_10002,N_10181);
and U10317 (N_10317,N_10145,N_10178);
nor U10318 (N_10318,N_10104,N_10091);
nor U10319 (N_10319,N_10136,N_10027);
or U10320 (N_10320,N_10053,N_10024);
xnor U10321 (N_10321,N_10067,N_10152);
xor U10322 (N_10322,N_10162,N_10092);
xnor U10323 (N_10323,N_10016,N_10008);
and U10324 (N_10324,N_10018,N_10017);
and U10325 (N_10325,N_10135,N_10083);
xnor U10326 (N_10326,N_10012,N_10065);
nand U10327 (N_10327,N_10040,N_10100);
or U10328 (N_10328,N_10047,N_10009);
nand U10329 (N_10329,N_10116,N_10172);
and U10330 (N_10330,N_10165,N_10031);
and U10331 (N_10331,N_10002,N_10075);
nand U10332 (N_10332,N_10188,N_10047);
and U10333 (N_10333,N_10100,N_10088);
xnor U10334 (N_10334,N_10015,N_10142);
or U10335 (N_10335,N_10038,N_10068);
and U10336 (N_10336,N_10184,N_10196);
and U10337 (N_10337,N_10145,N_10069);
and U10338 (N_10338,N_10098,N_10060);
or U10339 (N_10339,N_10081,N_10185);
and U10340 (N_10340,N_10139,N_10023);
nand U10341 (N_10341,N_10104,N_10144);
nand U10342 (N_10342,N_10188,N_10173);
nor U10343 (N_10343,N_10019,N_10091);
and U10344 (N_10344,N_10027,N_10177);
or U10345 (N_10345,N_10040,N_10096);
nand U10346 (N_10346,N_10172,N_10183);
and U10347 (N_10347,N_10103,N_10143);
nand U10348 (N_10348,N_10078,N_10106);
and U10349 (N_10349,N_10119,N_10168);
xor U10350 (N_10350,N_10109,N_10122);
nand U10351 (N_10351,N_10184,N_10180);
nand U10352 (N_10352,N_10104,N_10080);
xnor U10353 (N_10353,N_10051,N_10174);
or U10354 (N_10354,N_10114,N_10136);
nor U10355 (N_10355,N_10141,N_10104);
and U10356 (N_10356,N_10002,N_10131);
and U10357 (N_10357,N_10191,N_10145);
nand U10358 (N_10358,N_10194,N_10089);
nand U10359 (N_10359,N_10179,N_10147);
xor U10360 (N_10360,N_10163,N_10167);
or U10361 (N_10361,N_10163,N_10152);
nand U10362 (N_10362,N_10053,N_10131);
xnor U10363 (N_10363,N_10185,N_10052);
xnor U10364 (N_10364,N_10113,N_10109);
nand U10365 (N_10365,N_10037,N_10080);
and U10366 (N_10366,N_10005,N_10167);
and U10367 (N_10367,N_10157,N_10195);
or U10368 (N_10368,N_10178,N_10099);
xnor U10369 (N_10369,N_10102,N_10096);
nor U10370 (N_10370,N_10170,N_10179);
and U10371 (N_10371,N_10166,N_10072);
nand U10372 (N_10372,N_10180,N_10185);
and U10373 (N_10373,N_10184,N_10051);
and U10374 (N_10374,N_10061,N_10078);
nor U10375 (N_10375,N_10001,N_10064);
nor U10376 (N_10376,N_10124,N_10095);
nand U10377 (N_10377,N_10182,N_10159);
xnor U10378 (N_10378,N_10099,N_10045);
xor U10379 (N_10379,N_10168,N_10050);
nand U10380 (N_10380,N_10175,N_10183);
nand U10381 (N_10381,N_10001,N_10182);
or U10382 (N_10382,N_10094,N_10034);
xnor U10383 (N_10383,N_10045,N_10022);
or U10384 (N_10384,N_10158,N_10089);
nand U10385 (N_10385,N_10182,N_10046);
or U10386 (N_10386,N_10126,N_10170);
xnor U10387 (N_10387,N_10046,N_10031);
or U10388 (N_10388,N_10174,N_10132);
nand U10389 (N_10389,N_10058,N_10092);
and U10390 (N_10390,N_10132,N_10108);
or U10391 (N_10391,N_10131,N_10019);
nor U10392 (N_10392,N_10107,N_10124);
xor U10393 (N_10393,N_10114,N_10151);
nand U10394 (N_10394,N_10141,N_10090);
nor U10395 (N_10395,N_10123,N_10082);
nor U10396 (N_10396,N_10120,N_10007);
nand U10397 (N_10397,N_10009,N_10168);
xnor U10398 (N_10398,N_10132,N_10020);
xor U10399 (N_10399,N_10059,N_10047);
or U10400 (N_10400,N_10227,N_10279);
nand U10401 (N_10401,N_10204,N_10357);
nand U10402 (N_10402,N_10265,N_10262);
nand U10403 (N_10403,N_10318,N_10217);
nor U10404 (N_10404,N_10236,N_10307);
nand U10405 (N_10405,N_10292,N_10393);
and U10406 (N_10406,N_10297,N_10330);
nor U10407 (N_10407,N_10324,N_10243);
xor U10408 (N_10408,N_10367,N_10224);
nor U10409 (N_10409,N_10268,N_10310);
nor U10410 (N_10410,N_10364,N_10351);
and U10411 (N_10411,N_10216,N_10240);
and U10412 (N_10412,N_10349,N_10246);
nor U10413 (N_10413,N_10301,N_10396);
nor U10414 (N_10414,N_10370,N_10256);
nand U10415 (N_10415,N_10218,N_10321);
or U10416 (N_10416,N_10281,N_10341);
nand U10417 (N_10417,N_10336,N_10397);
or U10418 (N_10418,N_10372,N_10258);
xor U10419 (N_10419,N_10353,N_10275);
or U10420 (N_10420,N_10373,N_10305);
nand U10421 (N_10421,N_10222,N_10237);
and U10422 (N_10422,N_10298,N_10233);
or U10423 (N_10423,N_10394,N_10328);
nand U10424 (N_10424,N_10220,N_10302);
nor U10425 (N_10425,N_10366,N_10249);
nand U10426 (N_10426,N_10389,N_10391);
or U10427 (N_10427,N_10291,N_10337);
or U10428 (N_10428,N_10299,N_10230);
and U10429 (N_10429,N_10323,N_10280);
xor U10430 (N_10430,N_10311,N_10355);
xor U10431 (N_10431,N_10211,N_10270);
or U10432 (N_10432,N_10334,N_10374);
xor U10433 (N_10433,N_10360,N_10386);
xnor U10434 (N_10434,N_10207,N_10239);
xnor U10435 (N_10435,N_10362,N_10242);
nand U10436 (N_10436,N_10247,N_10329);
and U10437 (N_10437,N_10285,N_10284);
nor U10438 (N_10438,N_10325,N_10384);
xnor U10439 (N_10439,N_10331,N_10308);
nand U10440 (N_10440,N_10271,N_10276);
nor U10441 (N_10441,N_10335,N_10241);
nand U10442 (N_10442,N_10332,N_10273);
nor U10443 (N_10443,N_10382,N_10395);
or U10444 (N_10444,N_10206,N_10359);
and U10445 (N_10445,N_10277,N_10361);
or U10446 (N_10446,N_10322,N_10293);
xor U10447 (N_10447,N_10381,N_10288);
and U10448 (N_10448,N_10212,N_10201);
and U10449 (N_10449,N_10342,N_10315);
and U10450 (N_10450,N_10254,N_10223);
nor U10451 (N_10451,N_10289,N_10345);
or U10452 (N_10452,N_10225,N_10377);
nand U10453 (N_10453,N_10263,N_10229);
xor U10454 (N_10454,N_10253,N_10387);
and U10455 (N_10455,N_10304,N_10346);
xor U10456 (N_10456,N_10213,N_10363);
xnor U10457 (N_10457,N_10343,N_10278);
nor U10458 (N_10458,N_10252,N_10228);
or U10459 (N_10459,N_10221,N_10226);
and U10460 (N_10460,N_10269,N_10251);
nand U10461 (N_10461,N_10347,N_10309);
xor U10462 (N_10462,N_10290,N_10209);
or U10463 (N_10463,N_10295,N_10354);
and U10464 (N_10464,N_10303,N_10390);
nand U10465 (N_10465,N_10260,N_10385);
nor U10466 (N_10466,N_10344,N_10383);
nand U10467 (N_10467,N_10317,N_10375);
xnor U10468 (N_10468,N_10368,N_10286);
and U10469 (N_10469,N_10371,N_10264);
nor U10470 (N_10470,N_10338,N_10358);
or U10471 (N_10471,N_10378,N_10234);
xor U10472 (N_10472,N_10283,N_10215);
or U10473 (N_10473,N_10300,N_10294);
nand U10474 (N_10474,N_10365,N_10296);
nor U10475 (N_10475,N_10245,N_10244);
and U10476 (N_10476,N_10282,N_10261);
xnor U10477 (N_10477,N_10232,N_10339);
xor U10478 (N_10478,N_10219,N_10313);
nor U10479 (N_10479,N_10266,N_10314);
nor U10480 (N_10480,N_10312,N_10238);
nand U10481 (N_10481,N_10231,N_10274);
and U10482 (N_10482,N_10248,N_10235);
nand U10483 (N_10483,N_10200,N_10380);
nor U10484 (N_10484,N_10202,N_10327);
nand U10485 (N_10485,N_10306,N_10326);
and U10486 (N_10486,N_10255,N_10348);
nand U10487 (N_10487,N_10352,N_10203);
nand U10488 (N_10488,N_10267,N_10214);
nand U10489 (N_10489,N_10399,N_10259);
and U10490 (N_10490,N_10257,N_10208);
or U10491 (N_10491,N_10333,N_10205);
nand U10492 (N_10492,N_10210,N_10316);
nor U10493 (N_10493,N_10272,N_10379);
or U10494 (N_10494,N_10369,N_10250);
and U10495 (N_10495,N_10356,N_10376);
or U10496 (N_10496,N_10319,N_10340);
and U10497 (N_10497,N_10398,N_10392);
nor U10498 (N_10498,N_10320,N_10388);
nor U10499 (N_10499,N_10350,N_10287);
or U10500 (N_10500,N_10342,N_10369);
nor U10501 (N_10501,N_10284,N_10368);
nor U10502 (N_10502,N_10238,N_10325);
nor U10503 (N_10503,N_10319,N_10361);
and U10504 (N_10504,N_10297,N_10288);
nor U10505 (N_10505,N_10228,N_10340);
xor U10506 (N_10506,N_10324,N_10331);
and U10507 (N_10507,N_10288,N_10306);
and U10508 (N_10508,N_10223,N_10282);
nor U10509 (N_10509,N_10327,N_10254);
and U10510 (N_10510,N_10240,N_10325);
and U10511 (N_10511,N_10341,N_10295);
nand U10512 (N_10512,N_10368,N_10283);
nand U10513 (N_10513,N_10353,N_10225);
or U10514 (N_10514,N_10237,N_10335);
xnor U10515 (N_10515,N_10223,N_10219);
nor U10516 (N_10516,N_10223,N_10367);
nor U10517 (N_10517,N_10377,N_10301);
and U10518 (N_10518,N_10212,N_10231);
and U10519 (N_10519,N_10206,N_10224);
nor U10520 (N_10520,N_10232,N_10289);
or U10521 (N_10521,N_10288,N_10264);
and U10522 (N_10522,N_10273,N_10317);
xor U10523 (N_10523,N_10398,N_10259);
xor U10524 (N_10524,N_10341,N_10338);
xor U10525 (N_10525,N_10378,N_10289);
or U10526 (N_10526,N_10329,N_10378);
nand U10527 (N_10527,N_10353,N_10380);
xor U10528 (N_10528,N_10325,N_10256);
and U10529 (N_10529,N_10312,N_10382);
and U10530 (N_10530,N_10279,N_10253);
and U10531 (N_10531,N_10297,N_10253);
and U10532 (N_10532,N_10210,N_10204);
and U10533 (N_10533,N_10314,N_10345);
nand U10534 (N_10534,N_10239,N_10344);
nor U10535 (N_10535,N_10388,N_10368);
nand U10536 (N_10536,N_10223,N_10304);
and U10537 (N_10537,N_10373,N_10348);
nor U10538 (N_10538,N_10387,N_10206);
and U10539 (N_10539,N_10205,N_10397);
nand U10540 (N_10540,N_10273,N_10211);
xnor U10541 (N_10541,N_10265,N_10266);
xnor U10542 (N_10542,N_10301,N_10268);
and U10543 (N_10543,N_10381,N_10213);
or U10544 (N_10544,N_10260,N_10356);
nand U10545 (N_10545,N_10240,N_10362);
nand U10546 (N_10546,N_10303,N_10378);
nor U10547 (N_10547,N_10336,N_10284);
or U10548 (N_10548,N_10235,N_10220);
or U10549 (N_10549,N_10282,N_10390);
and U10550 (N_10550,N_10241,N_10248);
nand U10551 (N_10551,N_10280,N_10352);
and U10552 (N_10552,N_10282,N_10293);
or U10553 (N_10553,N_10201,N_10310);
or U10554 (N_10554,N_10265,N_10311);
and U10555 (N_10555,N_10207,N_10272);
and U10556 (N_10556,N_10364,N_10227);
xnor U10557 (N_10557,N_10351,N_10234);
xnor U10558 (N_10558,N_10234,N_10361);
xor U10559 (N_10559,N_10284,N_10378);
xor U10560 (N_10560,N_10298,N_10270);
and U10561 (N_10561,N_10255,N_10201);
nand U10562 (N_10562,N_10379,N_10273);
nor U10563 (N_10563,N_10310,N_10205);
and U10564 (N_10564,N_10396,N_10291);
nor U10565 (N_10565,N_10367,N_10270);
nand U10566 (N_10566,N_10393,N_10381);
xor U10567 (N_10567,N_10226,N_10207);
and U10568 (N_10568,N_10244,N_10320);
and U10569 (N_10569,N_10387,N_10261);
and U10570 (N_10570,N_10261,N_10219);
nor U10571 (N_10571,N_10308,N_10399);
or U10572 (N_10572,N_10310,N_10392);
xor U10573 (N_10573,N_10390,N_10269);
nand U10574 (N_10574,N_10380,N_10291);
or U10575 (N_10575,N_10353,N_10343);
nand U10576 (N_10576,N_10326,N_10320);
xnor U10577 (N_10577,N_10242,N_10383);
nor U10578 (N_10578,N_10219,N_10396);
nor U10579 (N_10579,N_10333,N_10229);
and U10580 (N_10580,N_10356,N_10223);
or U10581 (N_10581,N_10302,N_10261);
nand U10582 (N_10582,N_10222,N_10261);
and U10583 (N_10583,N_10355,N_10315);
and U10584 (N_10584,N_10212,N_10370);
nand U10585 (N_10585,N_10290,N_10363);
or U10586 (N_10586,N_10351,N_10229);
or U10587 (N_10587,N_10347,N_10244);
or U10588 (N_10588,N_10382,N_10342);
or U10589 (N_10589,N_10342,N_10329);
nand U10590 (N_10590,N_10356,N_10216);
nand U10591 (N_10591,N_10215,N_10393);
or U10592 (N_10592,N_10230,N_10207);
or U10593 (N_10593,N_10226,N_10255);
xor U10594 (N_10594,N_10204,N_10284);
nand U10595 (N_10595,N_10383,N_10318);
nor U10596 (N_10596,N_10270,N_10226);
or U10597 (N_10597,N_10238,N_10344);
or U10598 (N_10598,N_10311,N_10294);
and U10599 (N_10599,N_10361,N_10369);
xor U10600 (N_10600,N_10462,N_10408);
nand U10601 (N_10601,N_10458,N_10549);
and U10602 (N_10602,N_10596,N_10431);
nand U10603 (N_10603,N_10537,N_10435);
and U10604 (N_10604,N_10534,N_10580);
and U10605 (N_10605,N_10533,N_10539);
nand U10606 (N_10606,N_10532,N_10477);
nor U10607 (N_10607,N_10509,N_10540);
nor U10608 (N_10608,N_10516,N_10583);
and U10609 (N_10609,N_10470,N_10488);
nand U10610 (N_10610,N_10482,N_10418);
nor U10611 (N_10611,N_10444,N_10442);
nand U10612 (N_10612,N_10440,N_10581);
nor U10613 (N_10613,N_10510,N_10452);
nor U10614 (N_10614,N_10459,N_10475);
and U10615 (N_10615,N_10522,N_10529);
xnor U10616 (N_10616,N_10469,N_10541);
and U10617 (N_10617,N_10518,N_10437);
nand U10618 (N_10618,N_10557,N_10514);
or U10619 (N_10619,N_10584,N_10595);
nor U10620 (N_10620,N_10438,N_10515);
xnor U10621 (N_10621,N_10421,N_10519);
and U10622 (N_10622,N_10483,N_10547);
xor U10623 (N_10623,N_10496,N_10404);
nor U10624 (N_10624,N_10536,N_10552);
nand U10625 (N_10625,N_10570,N_10575);
nor U10626 (N_10626,N_10456,N_10490);
or U10627 (N_10627,N_10545,N_10463);
and U10628 (N_10628,N_10512,N_10531);
nand U10629 (N_10629,N_10402,N_10493);
nand U10630 (N_10630,N_10450,N_10585);
or U10631 (N_10631,N_10423,N_10484);
nor U10632 (N_10632,N_10426,N_10434);
or U10633 (N_10633,N_10525,N_10594);
nand U10634 (N_10634,N_10405,N_10568);
and U10635 (N_10635,N_10521,N_10553);
nor U10636 (N_10636,N_10400,N_10599);
and U10637 (N_10637,N_10411,N_10491);
xnor U10638 (N_10638,N_10507,N_10448);
and U10639 (N_10639,N_10429,N_10502);
nor U10640 (N_10640,N_10578,N_10406);
nor U10641 (N_10641,N_10466,N_10517);
and U10642 (N_10642,N_10453,N_10417);
or U10643 (N_10643,N_10454,N_10574);
nor U10644 (N_10644,N_10425,N_10576);
nor U10645 (N_10645,N_10443,N_10439);
or U10646 (N_10646,N_10546,N_10543);
and U10647 (N_10647,N_10455,N_10591);
or U10648 (N_10648,N_10449,N_10588);
or U10649 (N_10649,N_10415,N_10573);
and U10650 (N_10650,N_10587,N_10564);
nor U10651 (N_10651,N_10474,N_10447);
xor U10652 (N_10652,N_10446,N_10489);
xnor U10653 (N_10653,N_10562,N_10479);
and U10654 (N_10654,N_10542,N_10427);
nand U10655 (N_10655,N_10565,N_10577);
xnor U10656 (N_10656,N_10590,N_10555);
and U10657 (N_10657,N_10424,N_10481);
or U10658 (N_10658,N_10460,N_10551);
and U10659 (N_10659,N_10556,N_10480);
nand U10660 (N_10660,N_10433,N_10495);
nand U10661 (N_10661,N_10467,N_10486);
or U10662 (N_10662,N_10403,N_10410);
nor U10663 (N_10663,N_10511,N_10520);
nand U10664 (N_10664,N_10505,N_10451);
nand U10665 (N_10665,N_10506,N_10538);
or U10666 (N_10666,N_10544,N_10430);
and U10667 (N_10667,N_10476,N_10487);
xnor U10668 (N_10668,N_10571,N_10413);
or U10669 (N_10669,N_10428,N_10420);
or U10670 (N_10670,N_10558,N_10441);
xor U10671 (N_10671,N_10432,N_10500);
and U10672 (N_10672,N_10497,N_10414);
and U10673 (N_10673,N_10582,N_10485);
nand U10674 (N_10674,N_10407,N_10504);
nor U10675 (N_10675,N_10527,N_10567);
nor U10676 (N_10676,N_10503,N_10560);
nand U10677 (N_10677,N_10494,N_10561);
and U10678 (N_10678,N_10468,N_10501);
or U10679 (N_10679,N_10563,N_10461);
nor U10680 (N_10680,N_10589,N_10528);
xnor U10681 (N_10681,N_10492,N_10471);
and U10682 (N_10682,N_10566,N_10586);
or U10683 (N_10683,N_10550,N_10548);
xor U10684 (N_10684,N_10457,N_10593);
nand U10685 (N_10685,N_10523,N_10416);
xnor U10686 (N_10686,N_10530,N_10598);
nand U10687 (N_10687,N_10445,N_10535);
xnor U10688 (N_10688,N_10478,N_10401);
nor U10689 (N_10689,N_10409,N_10569);
or U10690 (N_10690,N_10508,N_10464);
nand U10691 (N_10691,N_10498,N_10499);
and U10692 (N_10692,N_10572,N_10513);
xor U10693 (N_10693,N_10526,N_10436);
xor U10694 (N_10694,N_10554,N_10419);
and U10695 (N_10695,N_10579,N_10592);
or U10696 (N_10696,N_10472,N_10422);
nand U10697 (N_10697,N_10597,N_10559);
or U10698 (N_10698,N_10412,N_10524);
or U10699 (N_10699,N_10465,N_10473);
xor U10700 (N_10700,N_10442,N_10534);
nor U10701 (N_10701,N_10489,N_10466);
nand U10702 (N_10702,N_10477,N_10499);
and U10703 (N_10703,N_10443,N_10515);
or U10704 (N_10704,N_10414,N_10560);
or U10705 (N_10705,N_10458,N_10578);
nor U10706 (N_10706,N_10477,N_10571);
nand U10707 (N_10707,N_10517,N_10461);
nand U10708 (N_10708,N_10479,N_10491);
and U10709 (N_10709,N_10479,N_10554);
or U10710 (N_10710,N_10412,N_10589);
nand U10711 (N_10711,N_10500,N_10441);
or U10712 (N_10712,N_10427,N_10502);
xor U10713 (N_10713,N_10592,N_10580);
nand U10714 (N_10714,N_10516,N_10401);
and U10715 (N_10715,N_10548,N_10498);
or U10716 (N_10716,N_10481,N_10572);
nand U10717 (N_10717,N_10498,N_10550);
xnor U10718 (N_10718,N_10442,N_10518);
or U10719 (N_10719,N_10513,N_10438);
nand U10720 (N_10720,N_10461,N_10579);
xor U10721 (N_10721,N_10419,N_10446);
and U10722 (N_10722,N_10458,N_10471);
and U10723 (N_10723,N_10419,N_10504);
or U10724 (N_10724,N_10564,N_10436);
xor U10725 (N_10725,N_10535,N_10577);
nor U10726 (N_10726,N_10479,N_10481);
nand U10727 (N_10727,N_10531,N_10488);
or U10728 (N_10728,N_10433,N_10514);
nand U10729 (N_10729,N_10599,N_10458);
nor U10730 (N_10730,N_10423,N_10451);
and U10731 (N_10731,N_10433,N_10448);
nand U10732 (N_10732,N_10476,N_10585);
nor U10733 (N_10733,N_10420,N_10563);
nand U10734 (N_10734,N_10530,N_10571);
nand U10735 (N_10735,N_10413,N_10514);
nand U10736 (N_10736,N_10434,N_10573);
nor U10737 (N_10737,N_10494,N_10436);
or U10738 (N_10738,N_10488,N_10450);
xnor U10739 (N_10739,N_10519,N_10432);
or U10740 (N_10740,N_10486,N_10490);
nor U10741 (N_10741,N_10596,N_10426);
xor U10742 (N_10742,N_10432,N_10431);
and U10743 (N_10743,N_10512,N_10598);
xnor U10744 (N_10744,N_10559,N_10551);
nand U10745 (N_10745,N_10554,N_10411);
and U10746 (N_10746,N_10491,N_10487);
nor U10747 (N_10747,N_10465,N_10447);
or U10748 (N_10748,N_10523,N_10560);
xnor U10749 (N_10749,N_10490,N_10408);
and U10750 (N_10750,N_10571,N_10551);
or U10751 (N_10751,N_10514,N_10446);
nor U10752 (N_10752,N_10566,N_10400);
nand U10753 (N_10753,N_10528,N_10499);
or U10754 (N_10754,N_10408,N_10410);
or U10755 (N_10755,N_10424,N_10495);
xnor U10756 (N_10756,N_10491,N_10594);
or U10757 (N_10757,N_10410,N_10532);
xnor U10758 (N_10758,N_10592,N_10515);
xor U10759 (N_10759,N_10571,N_10474);
nand U10760 (N_10760,N_10441,N_10449);
or U10761 (N_10761,N_10402,N_10589);
or U10762 (N_10762,N_10564,N_10478);
nor U10763 (N_10763,N_10589,N_10599);
xor U10764 (N_10764,N_10495,N_10595);
and U10765 (N_10765,N_10572,N_10412);
nand U10766 (N_10766,N_10502,N_10593);
xnor U10767 (N_10767,N_10488,N_10431);
nor U10768 (N_10768,N_10587,N_10543);
xnor U10769 (N_10769,N_10590,N_10430);
nand U10770 (N_10770,N_10544,N_10480);
xnor U10771 (N_10771,N_10591,N_10431);
and U10772 (N_10772,N_10509,N_10414);
xor U10773 (N_10773,N_10565,N_10483);
xor U10774 (N_10774,N_10476,N_10412);
and U10775 (N_10775,N_10402,N_10497);
xor U10776 (N_10776,N_10559,N_10547);
or U10777 (N_10777,N_10409,N_10465);
or U10778 (N_10778,N_10470,N_10478);
or U10779 (N_10779,N_10448,N_10509);
or U10780 (N_10780,N_10592,N_10582);
nor U10781 (N_10781,N_10479,N_10536);
xor U10782 (N_10782,N_10561,N_10599);
nor U10783 (N_10783,N_10532,N_10408);
nand U10784 (N_10784,N_10473,N_10530);
and U10785 (N_10785,N_10402,N_10561);
xor U10786 (N_10786,N_10419,N_10451);
or U10787 (N_10787,N_10464,N_10591);
nand U10788 (N_10788,N_10521,N_10427);
xor U10789 (N_10789,N_10586,N_10439);
nand U10790 (N_10790,N_10477,N_10412);
xor U10791 (N_10791,N_10529,N_10518);
nor U10792 (N_10792,N_10507,N_10466);
nor U10793 (N_10793,N_10521,N_10479);
xor U10794 (N_10794,N_10520,N_10563);
nor U10795 (N_10795,N_10436,N_10428);
and U10796 (N_10796,N_10564,N_10416);
and U10797 (N_10797,N_10401,N_10407);
nand U10798 (N_10798,N_10441,N_10406);
and U10799 (N_10799,N_10443,N_10502);
nand U10800 (N_10800,N_10774,N_10748);
and U10801 (N_10801,N_10775,N_10608);
nand U10802 (N_10802,N_10730,N_10684);
nor U10803 (N_10803,N_10744,N_10705);
xnor U10804 (N_10804,N_10767,N_10791);
nor U10805 (N_10805,N_10607,N_10788);
xnor U10806 (N_10806,N_10781,N_10639);
and U10807 (N_10807,N_10752,N_10689);
xor U10808 (N_10808,N_10606,N_10661);
nand U10809 (N_10809,N_10720,N_10642);
xnor U10810 (N_10810,N_10600,N_10611);
and U10811 (N_10811,N_10717,N_10778);
or U10812 (N_10812,N_10624,N_10612);
nor U10813 (N_10813,N_10754,N_10671);
or U10814 (N_10814,N_10602,N_10652);
or U10815 (N_10815,N_10763,N_10727);
nor U10816 (N_10816,N_10615,N_10732);
xor U10817 (N_10817,N_10660,N_10659);
and U10818 (N_10818,N_10790,N_10758);
and U10819 (N_10819,N_10726,N_10666);
and U10820 (N_10820,N_10632,N_10749);
and U10821 (N_10821,N_10703,N_10773);
nand U10822 (N_10822,N_10628,N_10690);
and U10823 (N_10823,N_10731,N_10698);
nand U10824 (N_10824,N_10765,N_10750);
nor U10825 (N_10825,N_10709,N_10658);
nand U10826 (N_10826,N_10616,N_10685);
or U10827 (N_10827,N_10793,N_10776);
nor U10828 (N_10828,N_10687,N_10777);
or U10829 (N_10829,N_10707,N_10795);
xnor U10830 (N_10830,N_10604,N_10619);
nor U10831 (N_10831,N_10649,N_10760);
nor U10832 (N_10832,N_10620,N_10710);
nor U10833 (N_10833,N_10735,N_10622);
xnor U10834 (N_10834,N_10654,N_10626);
nor U10835 (N_10835,N_10746,N_10677);
or U10836 (N_10836,N_10711,N_10673);
and U10837 (N_10837,N_10753,N_10734);
and U10838 (N_10838,N_10655,N_10609);
xnor U10839 (N_10839,N_10629,N_10702);
and U10840 (N_10840,N_10647,N_10798);
nand U10841 (N_10841,N_10761,N_10669);
or U10842 (N_10842,N_10693,N_10706);
or U10843 (N_10843,N_10739,N_10714);
or U10844 (N_10844,N_10621,N_10725);
nand U10845 (N_10845,N_10701,N_10796);
or U10846 (N_10846,N_10782,N_10623);
xor U10847 (N_10847,N_10724,N_10766);
nand U10848 (N_10848,N_10719,N_10665);
xor U10849 (N_10849,N_10715,N_10678);
xnor U10850 (N_10850,N_10713,N_10613);
nor U10851 (N_10851,N_10605,N_10721);
nand U10852 (N_10852,N_10716,N_10737);
and U10853 (N_10853,N_10764,N_10785);
and U10854 (N_10854,N_10745,N_10648);
xor U10855 (N_10855,N_10718,N_10797);
nor U10856 (N_10856,N_10601,N_10728);
nor U10857 (N_10857,N_10770,N_10771);
and U10858 (N_10858,N_10638,N_10683);
nand U10859 (N_10859,N_10614,N_10680);
nor U10860 (N_10860,N_10759,N_10769);
and U10861 (N_10861,N_10625,N_10653);
or U10862 (N_10862,N_10692,N_10668);
and U10863 (N_10863,N_10699,N_10787);
nor U10864 (N_10864,N_10603,N_10634);
or U10865 (N_10865,N_10741,N_10742);
nand U10866 (N_10866,N_10627,N_10700);
xnor U10867 (N_10867,N_10751,N_10743);
nand U10868 (N_10868,N_10786,N_10762);
nand U10869 (N_10869,N_10672,N_10682);
nand U10870 (N_10870,N_10662,N_10755);
nor U10871 (N_10871,N_10631,N_10756);
xnor U10872 (N_10872,N_10681,N_10617);
nor U10873 (N_10873,N_10779,N_10736);
xor U10874 (N_10874,N_10712,N_10768);
xnor U10875 (N_10875,N_10784,N_10723);
xor U10876 (N_10876,N_10694,N_10646);
xor U10877 (N_10877,N_10729,N_10792);
and U10878 (N_10878,N_10708,N_10722);
and U10879 (N_10879,N_10747,N_10618);
nand U10880 (N_10880,N_10686,N_10651);
nand U10881 (N_10881,N_10691,N_10645);
and U10882 (N_10882,N_10789,N_10664);
nor U10883 (N_10883,N_10667,N_10675);
nand U10884 (N_10884,N_10657,N_10610);
nand U10885 (N_10885,N_10641,N_10740);
nor U10886 (N_10886,N_10636,N_10780);
and U10887 (N_10887,N_10733,N_10696);
and U10888 (N_10888,N_10640,N_10674);
xnor U10889 (N_10889,N_10695,N_10783);
and U10890 (N_10890,N_10799,N_10644);
and U10891 (N_10891,N_10635,N_10688);
nand U10892 (N_10892,N_10704,N_10757);
or U10893 (N_10893,N_10794,N_10633);
xor U10894 (N_10894,N_10676,N_10650);
and U10895 (N_10895,N_10643,N_10772);
xnor U10896 (N_10896,N_10738,N_10630);
or U10897 (N_10897,N_10679,N_10637);
xnor U10898 (N_10898,N_10656,N_10670);
xnor U10899 (N_10899,N_10697,N_10663);
xor U10900 (N_10900,N_10691,N_10658);
nand U10901 (N_10901,N_10773,N_10720);
and U10902 (N_10902,N_10747,N_10764);
nand U10903 (N_10903,N_10655,N_10672);
xor U10904 (N_10904,N_10727,N_10784);
or U10905 (N_10905,N_10664,N_10726);
nor U10906 (N_10906,N_10625,N_10697);
nand U10907 (N_10907,N_10717,N_10654);
nor U10908 (N_10908,N_10695,N_10661);
nor U10909 (N_10909,N_10768,N_10680);
nor U10910 (N_10910,N_10727,N_10638);
nand U10911 (N_10911,N_10648,N_10604);
nand U10912 (N_10912,N_10747,N_10629);
or U10913 (N_10913,N_10675,N_10755);
or U10914 (N_10914,N_10791,N_10751);
and U10915 (N_10915,N_10635,N_10735);
nor U10916 (N_10916,N_10703,N_10664);
nor U10917 (N_10917,N_10738,N_10680);
nor U10918 (N_10918,N_10792,N_10688);
or U10919 (N_10919,N_10788,N_10731);
nand U10920 (N_10920,N_10636,N_10791);
or U10921 (N_10921,N_10681,N_10662);
or U10922 (N_10922,N_10603,N_10705);
and U10923 (N_10923,N_10673,N_10683);
and U10924 (N_10924,N_10611,N_10738);
nand U10925 (N_10925,N_10747,N_10750);
and U10926 (N_10926,N_10641,N_10745);
or U10927 (N_10927,N_10740,N_10609);
xnor U10928 (N_10928,N_10616,N_10602);
and U10929 (N_10929,N_10740,N_10621);
and U10930 (N_10930,N_10673,N_10763);
and U10931 (N_10931,N_10771,N_10672);
nor U10932 (N_10932,N_10627,N_10644);
nand U10933 (N_10933,N_10621,N_10615);
nand U10934 (N_10934,N_10631,N_10607);
nor U10935 (N_10935,N_10649,N_10671);
or U10936 (N_10936,N_10707,N_10659);
xor U10937 (N_10937,N_10780,N_10670);
or U10938 (N_10938,N_10683,N_10684);
nand U10939 (N_10939,N_10628,N_10644);
or U10940 (N_10940,N_10639,N_10690);
nand U10941 (N_10941,N_10667,N_10704);
and U10942 (N_10942,N_10688,N_10721);
or U10943 (N_10943,N_10785,N_10628);
nor U10944 (N_10944,N_10612,N_10756);
nand U10945 (N_10945,N_10786,N_10642);
xnor U10946 (N_10946,N_10626,N_10757);
xnor U10947 (N_10947,N_10792,N_10682);
xor U10948 (N_10948,N_10779,N_10754);
and U10949 (N_10949,N_10617,N_10763);
nand U10950 (N_10950,N_10675,N_10622);
xnor U10951 (N_10951,N_10642,N_10616);
xnor U10952 (N_10952,N_10604,N_10796);
nor U10953 (N_10953,N_10757,N_10709);
or U10954 (N_10954,N_10766,N_10660);
or U10955 (N_10955,N_10617,N_10737);
nor U10956 (N_10956,N_10669,N_10715);
nand U10957 (N_10957,N_10744,N_10766);
nand U10958 (N_10958,N_10632,N_10781);
nand U10959 (N_10959,N_10767,N_10625);
nor U10960 (N_10960,N_10679,N_10772);
nor U10961 (N_10961,N_10761,N_10659);
nor U10962 (N_10962,N_10780,N_10683);
nand U10963 (N_10963,N_10694,N_10748);
or U10964 (N_10964,N_10683,N_10737);
or U10965 (N_10965,N_10783,N_10660);
nor U10966 (N_10966,N_10770,N_10753);
xor U10967 (N_10967,N_10674,N_10649);
nor U10968 (N_10968,N_10780,N_10790);
nor U10969 (N_10969,N_10671,N_10641);
and U10970 (N_10970,N_10629,N_10662);
nand U10971 (N_10971,N_10729,N_10757);
or U10972 (N_10972,N_10683,N_10786);
nand U10973 (N_10973,N_10711,N_10766);
nor U10974 (N_10974,N_10687,N_10663);
or U10975 (N_10975,N_10781,N_10743);
xor U10976 (N_10976,N_10653,N_10701);
xor U10977 (N_10977,N_10701,N_10709);
or U10978 (N_10978,N_10787,N_10698);
nand U10979 (N_10979,N_10696,N_10734);
and U10980 (N_10980,N_10636,N_10760);
or U10981 (N_10981,N_10642,N_10740);
or U10982 (N_10982,N_10775,N_10730);
or U10983 (N_10983,N_10744,N_10669);
and U10984 (N_10984,N_10702,N_10675);
and U10985 (N_10985,N_10701,N_10670);
nor U10986 (N_10986,N_10716,N_10678);
or U10987 (N_10987,N_10786,N_10633);
nor U10988 (N_10988,N_10786,N_10655);
nor U10989 (N_10989,N_10640,N_10643);
and U10990 (N_10990,N_10708,N_10613);
xnor U10991 (N_10991,N_10751,N_10748);
nand U10992 (N_10992,N_10701,N_10703);
or U10993 (N_10993,N_10750,N_10650);
and U10994 (N_10994,N_10664,N_10612);
and U10995 (N_10995,N_10758,N_10632);
nand U10996 (N_10996,N_10624,N_10601);
xor U10997 (N_10997,N_10736,N_10671);
nand U10998 (N_10998,N_10798,N_10637);
nor U10999 (N_10999,N_10688,N_10665);
and U11000 (N_11000,N_10936,N_10942);
nor U11001 (N_11001,N_10969,N_10850);
and U11002 (N_11002,N_10987,N_10892);
or U11003 (N_11003,N_10950,N_10912);
and U11004 (N_11004,N_10851,N_10813);
nand U11005 (N_11005,N_10970,N_10983);
and U11006 (N_11006,N_10804,N_10800);
or U11007 (N_11007,N_10839,N_10894);
or U11008 (N_11008,N_10827,N_10842);
xnor U11009 (N_11009,N_10848,N_10844);
nand U11010 (N_11010,N_10869,N_10996);
nor U11011 (N_11011,N_10974,N_10958);
and U11012 (N_11012,N_10823,N_10986);
nand U11013 (N_11013,N_10917,N_10882);
or U11014 (N_11014,N_10954,N_10862);
or U11015 (N_11015,N_10973,N_10898);
nand U11016 (N_11016,N_10870,N_10856);
xnor U11017 (N_11017,N_10975,N_10901);
nand U11018 (N_11018,N_10841,N_10812);
xor U11019 (N_11019,N_10989,N_10854);
nor U11020 (N_11020,N_10884,N_10890);
nor U11021 (N_11021,N_10923,N_10941);
xnor U11022 (N_11022,N_10947,N_10944);
or U11023 (N_11023,N_10891,N_10935);
nand U11024 (N_11024,N_10913,N_10997);
and U11025 (N_11025,N_10979,N_10809);
and U11026 (N_11026,N_10904,N_10802);
nand U11027 (N_11027,N_10834,N_10853);
or U11028 (N_11028,N_10908,N_10963);
xnor U11029 (N_11029,N_10999,N_10879);
nor U11030 (N_11030,N_10876,N_10925);
and U11031 (N_11031,N_10980,N_10831);
and U11032 (N_11032,N_10982,N_10959);
and U11033 (N_11033,N_10865,N_10934);
xnor U11034 (N_11034,N_10808,N_10911);
nor U11035 (N_11035,N_10825,N_10992);
nand U11036 (N_11036,N_10822,N_10968);
or U11037 (N_11037,N_10920,N_10885);
or U11038 (N_11038,N_10860,N_10932);
nand U11039 (N_11039,N_10994,N_10810);
or U11040 (N_11040,N_10849,N_10918);
xnor U11041 (N_11041,N_10818,N_10868);
nand U11042 (N_11042,N_10875,N_10805);
and U11043 (N_11043,N_10962,N_10937);
or U11044 (N_11044,N_10919,N_10988);
and U11045 (N_11045,N_10815,N_10931);
and U11046 (N_11046,N_10867,N_10806);
nor U11047 (N_11047,N_10828,N_10964);
nand U11048 (N_11048,N_10859,N_10829);
nor U11049 (N_11049,N_10816,N_10840);
nand U11050 (N_11050,N_10993,N_10945);
xor U11051 (N_11051,N_10955,N_10826);
nor U11052 (N_11052,N_10921,N_10960);
nor U11053 (N_11053,N_10977,N_10837);
xnor U11054 (N_11054,N_10895,N_10863);
nand U11055 (N_11055,N_10916,N_10838);
and U11056 (N_11056,N_10928,N_10924);
xnor U11057 (N_11057,N_10910,N_10902);
xnor U11058 (N_11058,N_10817,N_10907);
or U11059 (N_11059,N_10887,N_10909);
nand U11060 (N_11060,N_10881,N_10933);
nand U11061 (N_11061,N_10940,N_10893);
nor U11062 (N_11062,N_10835,N_10801);
or U11063 (N_11063,N_10858,N_10845);
nor U11064 (N_11064,N_10833,N_10990);
or U11065 (N_11065,N_10998,N_10930);
nor U11066 (N_11066,N_10871,N_10900);
or U11067 (N_11067,N_10946,N_10939);
and U11068 (N_11068,N_10880,N_10814);
or U11069 (N_11069,N_10836,N_10803);
xor U11070 (N_11070,N_10807,N_10883);
nor U11071 (N_11071,N_10929,N_10972);
or U11072 (N_11072,N_10965,N_10906);
and U11073 (N_11073,N_10981,N_10866);
or U11074 (N_11074,N_10926,N_10889);
nand U11075 (N_11075,N_10857,N_10832);
xnor U11076 (N_11076,N_10984,N_10846);
xor U11077 (N_11077,N_10985,N_10943);
nor U11078 (N_11078,N_10886,N_10905);
and U11079 (N_11079,N_10878,N_10949);
xnor U11080 (N_11080,N_10967,N_10952);
xnor U11081 (N_11081,N_10976,N_10995);
nor U11082 (N_11082,N_10948,N_10873);
nor U11083 (N_11083,N_10847,N_10927);
and U11084 (N_11084,N_10899,N_10855);
and U11085 (N_11085,N_10861,N_10897);
or U11086 (N_11086,N_10821,N_10956);
and U11087 (N_11087,N_10978,N_10914);
xor U11088 (N_11088,N_10877,N_10991);
xnor U11089 (N_11089,N_10951,N_10896);
and U11090 (N_11090,N_10843,N_10819);
or U11091 (N_11091,N_10971,N_10961);
nand U11092 (N_11092,N_10874,N_10820);
or U11093 (N_11093,N_10811,N_10953);
nor U11094 (N_11094,N_10957,N_10888);
or U11095 (N_11095,N_10922,N_10864);
and U11096 (N_11096,N_10915,N_10830);
nor U11097 (N_11097,N_10903,N_10966);
or U11098 (N_11098,N_10938,N_10872);
nor U11099 (N_11099,N_10852,N_10824);
and U11100 (N_11100,N_10834,N_10920);
and U11101 (N_11101,N_10991,N_10812);
nand U11102 (N_11102,N_10999,N_10845);
or U11103 (N_11103,N_10961,N_10873);
nor U11104 (N_11104,N_10843,N_10972);
nand U11105 (N_11105,N_10927,N_10974);
xnor U11106 (N_11106,N_10803,N_10826);
or U11107 (N_11107,N_10970,N_10932);
xor U11108 (N_11108,N_10893,N_10887);
or U11109 (N_11109,N_10994,N_10988);
xnor U11110 (N_11110,N_10812,N_10854);
or U11111 (N_11111,N_10845,N_10961);
or U11112 (N_11112,N_10897,N_10960);
or U11113 (N_11113,N_10901,N_10966);
and U11114 (N_11114,N_10905,N_10802);
xor U11115 (N_11115,N_10997,N_10845);
xnor U11116 (N_11116,N_10998,N_10860);
nor U11117 (N_11117,N_10992,N_10969);
and U11118 (N_11118,N_10856,N_10875);
or U11119 (N_11119,N_10836,N_10915);
and U11120 (N_11120,N_10906,N_10905);
xnor U11121 (N_11121,N_10819,N_10968);
xnor U11122 (N_11122,N_10932,N_10905);
xnor U11123 (N_11123,N_10828,N_10982);
nor U11124 (N_11124,N_10902,N_10869);
nand U11125 (N_11125,N_10933,N_10948);
nand U11126 (N_11126,N_10934,N_10886);
nor U11127 (N_11127,N_10999,N_10870);
or U11128 (N_11128,N_10904,N_10998);
nand U11129 (N_11129,N_10867,N_10868);
xnor U11130 (N_11130,N_10888,N_10833);
xor U11131 (N_11131,N_10955,N_10847);
nor U11132 (N_11132,N_10989,N_10845);
or U11133 (N_11133,N_10908,N_10803);
and U11134 (N_11134,N_10972,N_10995);
nand U11135 (N_11135,N_10802,N_10820);
or U11136 (N_11136,N_10813,N_10880);
nand U11137 (N_11137,N_10819,N_10806);
nor U11138 (N_11138,N_10983,N_10944);
xnor U11139 (N_11139,N_10965,N_10832);
and U11140 (N_11140,N_10964,N_10891);
or U11141 (N_11141,N_10804,N_10838);
and U11142 (N_11142,N_10961,N_10813);
or U11143 (N_11143,N_10901,N_10900);
nor U11144 (N_11144,N_10967,N_10966);
nand U11145 (N_11145,N_10821,N_10911);
nor U11146 (N_11146,N_10993,N_10979);
nor U11147 (N_11147,N_10875,N_10903);
and U11148 (N_11148,N_10987,N_10937);
xor U11149 (N_11149,N_10833,N_10989);
nor U11150 (N_11150,N_10930,N_10882);
nand U11151 (N_11151,N_10879,N_10903);
and U11152 (N_11152,N_10889,N_10900);
and U11153 (N_11153,N_10941,N_10818);
nor U11154 (N_11154,N_10995,N_10954);
and U11155 (N_11155,N_10981,N_10884);
nand U11156 (N_11156,N_10803,N_10983);
xnor U11157 (N_11157,N_10909,N_10886);
xor U11158 (N_11158,N_10893,N_10903);
and U11159 (N_11159,N_10908,N_10983);
or U11160 (N_11160,N_10928,N_10923);
nor U11161 (N_11161,N_10815,N_10883);
nand U11162 (N_11162,N_10957,N_10809);
xor U11163 (N_11163,N_10913,N_10944);
nor U11164 (N_11164,N_10887,N_10852);
or U11165 (N_11165,N_10872,N_10805);
and U11166 (N_11166,N_10911,N_10895);
or U11167 (N_11167,N_10988,N_10959);
nor U11168 (N_11168,N_10864,N_10986);
and U11169 (N_11169,N_10891,N_10966);
or U11170 (N_11170,N_10920,N_10847);
or U11171 (N_11171,N_10857,N_10975);
and U11172 (N_11172,N_10923,N_10905);
nor U11173 (N_11173,N_10885,N_10811);
xor U11174 (N_11174,N_10952,N_10870);
nand U11175 (N_11175,N_10991,N_10996);
and U11176 (N_11176,N_10964,N_10934);
or U11177 (N_11177,N_10937,N_10809);
xor U11178 (N_11178,N_10834,N_10847);
xor U11179 (N_11179,N_10840,N_10939);
and U11180 (N_11180,N_10954,N_10833);
nand U11181 (N_11181,N_10878,N_10918);
nand U11182 (N_11182,N_10846,N_10857);
or U11183 (N_11183,N_10954,N_10919);
nor U11184 (N_11184,N_10990,N_10915);
and U11185 (N_11185,N_10917,N_10918);
and U11186 (N_11186,N_10997,N_10943);
nor U11187 (N_11187,N_10933,N_10930);
nor U11188 (N_11188,N_10903,N_10870);
and U11189 (N_11189,N_10926,N_10832);
nor U11190 (N_11190,N_10888,N_10800);
xor U11191 (N_11191,N_10867,N_10950);
xnor U11192 (N_11192,N_10956,N_10904);
nand U11193 (N_11193,N_10863,N_10837);
or U11194 (N_11194,N_10829,N_10803);
and U11195 (N_11195,N_10855,N_10924);
nand U11196 (N_11196,N_10910,N_10989);
nor U11197 (N_11197,N_10834,N_10825);
xor U11198 (N_11198,N_10947,N_10940);
nand U11199 (N_11199,N_10809,N_10892);
xor U11200 (N_11200,N_11039,N_11025);
or U11201 (N_11201,N_11097,N_11046);
and U11202 (N_11202,N_11145,N_11019);
nor U11203 (N_11203,N_11027,N_11095);
or U11204 (N_11204,N_11134,N_11100);
nor U11205 (N_11205,N_11191,N_11018);
nor U11206 (N_11206,N_11136,N_11031);
or U11207 (N_11207,N_11158,N_11092);
xnor U11208 (N_11208,N_11075,N_11020);
nor U11209 (N_11209,N_11198,N_11035);
xor U11210 (N_11210,N_11183,N_11115);
or U11211 (N_11211,N_11108,N_11012);
and U11212 (N_11212,N_11118,N_11194);
xnor U11213 (N_11213,N_11176,N_11143);
nand U11214 (N_11214,N_11036,N_11080);
or U11215 (N_11215,N_11008,N_11053);
and U11216 (N_11216,N_11014,N_11088);
xnor U11217 (N_11217,N_11180,N_11022);
nor U11218 (N_11218,N_11187,N_11041);
or U11219 (N_11219,N_11178,N_11166);
nand U11220 (N_11220,N_11101,N_11132);
nand U11221 (N_11221,N_11029,N_11123);
or U11222 (N_11222,N_11000,N_11077);
and U11223 (N_11223,N_11079,N_11148);
nor U11224 (N_11224,N_11156,N_11107);
nand U11225 (N_11225,N_11061,N_11151);
xnor U11226 (N_11226,N_11109,N_11131);
or U11227 (N_11227,N_11174,N_11150);
and U11228 (N_11228,N_11056,N_11162);
or U11229 (N_11229,N_11179,N_11116);
or U11230 (N_11230,N_11114,N_11023);
or U11231 (N_11231,N_11121,N_11138);
xnor U11232 (N_11232,N_11050,N_11047);
or U11233 (N_11233,N_11074,N_11129);
or U11234 (N_11234,N_11028,N_11152);
and U11235 (N_11235,N_11110,N_11146);
nand U11236 (N_11236,N_11163,N_11173);
or U11237 (N_11237,N_11044,N_11051);
nor U11238 (N_11238,N_11072,N_11172);
and U11239 (N_11239,N_11111,N_11052);
nor U11240 (N_11240,N_11124,N_11021);
nand U11241 (N_11241,N_11093,N_11113);
xor U11242 (N_11242,N_11057,N_11190);
and U11243 (N_11243,N_11155,N_11011);
nand U11244 (N_11244,N_11161,N_11032);
nand U11245 (N_11245,N_11071,N_11167);
or U11246 (N_11246,N_11004,N_11017);
nand U11247 (N_11247,N_11096,N_11182);
and U11248 (N_11248,N_11060,N_11013);
and U11249 (N_11249,N_11153,N_11104);
xor U11250 (N_11250,N_11103,N_11034);
and U11251 (N_11251,N_11122,N_11165);
nor U11252 (N_11252,N_11157,N_11144);
or U11253 (N_11253,N_11159,N_11049);
nor U11254 (N_11254,N_11065,N_11186);
xnor U11255 (N_11255,N_11007,N_11001);
nand U11256 (N_11256,N_11141,N_11058);
and U11257 (N_11257,N_11195,N_11086);
and U11258 (N_11258,N_11083,N_11030);
xnor U11259 (N_11259,N_11084,N_11085);
and U11260 (N_11260,N_11140,N_11081);
nand U11261 (N_11261,N_11016,N_11147);
xnor U11262 (N_11262,N_11139,N_11154);
and U11263 (N_11263,N_11015,N_11037);
or U11264 (N_11264,N_11119,N_11185);
nand U11265 (N_11265,N_11181,N_11076);
and U11266 (N_11266,N_11054,N_11135);
nor U11267 (N_11267,N_11199,N_11087);
nor U11268 (N_11268,N_11098,N_11005);
and U11269 (N_11269,N_11043,N_11171);
or U11270 (N_11270,N_11009,N_11073);
or U11271 (N_11271,N_11040,N_11137);
and U11272 (N_11272,N_11026,N_11188);
nand U11273 (N_11273,N_11130,N_11090);
nor U11274 (N_11274,N_11102,N_11067);
xor U11275 (N_11275,N_11045,N_11125);
xor U11276 (N_11276,N_11126,N_11059);
nand U11277 (N_11277,N_11033,N_11105);
and U11278 (N_11278,N_11070,N_11089);
nor U11279 (N_11279,N_11082,N_11133);
or U11280 (N_11280,N_11160,N_11069);
nor U11281 (N_11281,N_11038,N_11063);
or U11282 (N_11282,N_11055,N_11184);
nand U11283 (N_11283,N_11078,N_11024);
nand U11284 (N_11284,N_11042,N_11003);
or U11285 (N_11285,N_11197,N_11010);
nor U11286 (N_11286,N_11168,N_11106);
or U11287 (N_11287,N_11068,N_11164);
xor U11288 (N_11288,N_11002,N_11192);
or U11289 (N_11289,N_11048,N_11112);
nand U11290 (N_11290,N_11064,N_11062);
xnor U11291 (N_11291,N_11169,N_11177);
and U11292 (N_11292,N_11170,N_11127);
nand U11293 (N_11293,N_11066,N_11120);
nand U11294 (N_11294,N_11006,N_11149);
nand U11295 (N_11295,N_11128,N_11094);
xnor U11296 (N_11296,N_11175,N_11196);
xor U11297 (N_11297,N_11099,N_11142);
and U11298 (N_11298,N_11091,N_11189);
and U11299 (N_11299,N_11193,N_11117);
nor U11300 (N_11300,N_11159,N_11012);
nand U11301 (N_11301,N_11129,N_11035);
xnor U11302 (N_11302,N_11013,N_11086);
or U11303 (N_11303,N_11065,N_11063);
and U11304 (N_11304,N_11159,N_11077);
and U11305 (N_11305,N_11162,N_11067);
or U11306 (N_11306,N_11139,N_11137);
nand U11307 (N_11307,N_11136,N_11199);
nor U11308 (N_11308,N_11131,N_11107);
xnor U11309 (N_11309,N_11010,N_11132);
nand U11310 (N_11310,N_11029,N_11180);
nor U11311 (N_11311,N_11103,N_11076);
nand U11312 (N_11312,N_11072,N_11137);
nor U11313 (N_11313,N_11086,N_11148);
and U11314 (N_11314,N_11049,N_11153);
or U11315 (N_11315,N_11177,N_11030);
nand U11316 (N_11316,N_11134,N_11094);
and U11317 (N_11317,N_11139,N_11165);
and U11318 (N_11318,N_11150,N_11038);
xnor U11319 (N_11319,N_11024,N_11113);
nor U11320 (N_11320,N_11047,N_11141);
xnor U11321 (N_11321,N_11189,N_11041);
or U11322 (N_11322,N_11022,N_11124);
or U11323 (N_11323,N_11127,N_11006);
or U11324 (N_11324,N_11123,N_11131);
nor U11325 (N_11325,N_11142,N_11010);
and U11326 (N_11326,N_11040,N_11085);
or U11327 (N_11327,N_11016,N_11130);
or U11328 (N_11328,N_11093,N_11002);
and U11329 (N_11329,N_11061,N_11059);
or U11330 (N_11330,N_11130,N_11098);
and U11331 (N_11331,N_11111,N_11121);
and U11332 (N_11332,N_11048,N_11028);
xor U11333 (N_11333,N_11006,N_11028);
or U11334 (N_11334,N_11032,N_11141);
and U11335 (N_11335,N_11079,N_11155);
or U11336 (N_11336,N_11027,N_11150);
and U11337 (N_11337,N_11167,N_11194);
xnor U11338 (N_11338,N_11166,N_11181);
nand U11339 (N_11339,N_11076,N_11063);
and U11340 (N_11340,N_11152,N_11050);
and U11341 (N_11341,N_11176,N_11090);
or U11342 (N_11342,N_11010,N_11198);
or U11343 (N_11343,N_11078,N_11144);
and U11344 (N_11344,N_11139,N_11093);
xor U11345 (N_11345,N_11139,N_11133);
nor U11346 (N_11346,N_11059,N_11096);
nand U11347 (N_11347,N_11076,N_11101);
nor U11348 (N_11348,N_11097,N_11066);
and U11349 (N_11349,N_11187,N_11029);
nor U11350 (N_11350,N_11036,N_11089);
nor U11351 (N_11351,N_11161,N_11126);
and U11352 (N_11352,N_11100,N_11017);
xnor U11353 (N_11353,N_11174,N_11063);
or U11354 (N_11354,N_11171,N_11050);
nand U11355 (N_11355,N_11138,N_11092);
or U11356 (N_11356,N_11108,N_11177);
and U11357 (N_11357,N_11033,N_11100);
nor U11358 (N_11358,N_11154,N_11098);
or U11359 (N_11359,N_11134,N_11187);
or U11360 (N_11360,N_11136,N_11108);
nor U11361 (N_11361,N_11111,N_11110);
xor U11362 (N_11362,N_11094,N_11080);
and U11363 (N_11363,N_11070,N_11057);
and U11364 (N_11364,N_11131,N_11066);
and U11365 (N_11365,N_11101,N_11025);
or U11366 (N_11366,N_11136,N_11068);
nor U11367 (N_11367,N_11019,N_11040);
nor U11368 (N_11368,N_11000,N_11145);
and U11369 (N_11369,N_11168,N_11124);
xnor U11370 (N_11370,N_11136,N_11010);
xor U11371 (N_11371,N_11149,N_11100);
xnor U11372 (N_11372,N_11082,N_11121);
nor U11373 (N_11373,N_11003,N_11136);
nand U11374 (N_11374,N_11138,N_11170);
nor U11375 (N_11375,N_11172,N_11100);
or U11376 (N_11376,N_11160,N_11066);
xnor U11377 (N_11377,N_11078,N_11075);
nor U11378 (N_11378,N_11137,N_11157);
or U11379 (N_11379,N_11057,N_11053);
xnor U11380 (N_11380,N_11170,N_11115);
or U11381 (N_11381,N_11165,N_11029);
nor U11382 (N_11382,N_11145,N_11067);
and U11383 (N_11383,N_11046,N_11015);
xor U11384 (N_11384,N_11168,N_11096);
nor U11385 (N_11385,N_11027,N_11156);
nand U11386 (N_11386,N_11016,N_11173);
xor U11387 (N_11387,N_11041,N_11151);
nand U11388 (N_11388,N_11196,N_11172);
and U11389 (N_11389,N_11007,N_11066);
xnor U11390 (N_11390,N_11171,N_11133);
nand U11391 (N_11391,N_11197,N_11050);
or U11392 (N_11392,N_11156,N_11075);
and U11393 (N_11393,N_11085,N_11098);
nor U11394 (N_11394,N_11051,N_11037);
nor U11395 (N_11395,N_11130,N_11064);
xor U11396 (N_11396,N_11044,N_11161);
xor U11397 (N_11397,N_11004,N_11089);
xnor U11398 (N_11398,N_11142,N_11188);
or U11399 (N_11399,N_11001,N_11004);
nor U11400 (N_11400,N_11261,N_11316);
or U11401 (N_11401,N_11205,N_11323);
and U11402 (N_11402,N_11397,N_11273);
or U11403 (N_11403,N_11292,N_11245);
and U11404 (N_11404,N_11340,N_11398);
xnor U11405 (N_11405,N_11339,N_11239);
xor U11406 (N_11406,N_11229,N_11327);
or U11407 (N_11407,N_11221,N_11280);
or U11408 (N_11408,N_11289,N_11210);
or U11409 (N_11409,N_11347,N_11381);
nand U11410 (N_11410,N_11379,N_11212);
nor U11411 (N_11411,N_11356,N_11317);
and U11412 (N_11412,N_11399,N_11326);
and U11413 (N_11413,N_11308,N_11369);
xnor U11414 (N_11414,N_11258,N_11377);
nand U11415 (N_11415,N_11333,N_11311);
xnor U11416 (N_11416,N_11330,N_11386);
or U11417 (N_11417,N_11249,N_11274);
or U11418 (N_11418,N_11387,N_11259);
nand U11419 (N_11419,N_11354,N_11366);
and U11420 (N_11420,N_11237,N_11324);
xnor U11421 (N_11421,N_11305,N_11213);
xnor U11422 (N_11422,N_11337,N_11208);
xnor U11423 (N_11423,N_11359,N_11335);
nor U11424 (N_11424,N_11276,N_11263);
xnor U11425 (N_11425,N_11203,N_11296);
and U11426 (N_11426,N_11298,N_11270);
nand U11427 (N_11427,N_11376,N_11283);
xor U11428 (N_11428,N_11307,N_11243);
nand U11429 (N_11429,N_11312,N_11385);
or U11430 (N_11430,N_11220,N_11201);
or U11431 (N_11431,N_11288,N_11392);
and U11432 (N_11432,N_11267,N_11204);
nor U11433 (N_11433,N_11202,N_11368);
or U11434 (N_11434,N_11394,N_11351);
nand U11435 (N_11435,N_11375,N_11338);
or U11436 (N_11436,N_11269,N_11222);
nand U11437 (N_11437,N_11294,N_11299);
and U11438 (N_11438,N_11253,N_11309);
nor U11439 (N_11439,N_11236,N_11362);
nand U11440 (N_11440,N_11343,N_11371);
and U11441 (N_11441,N_11357,N_11272);
nor U11442 (N_11442,N_11279,N_11234);
xor U11443 (N_11443,N_11374,N_11364);
nor U11444 (N_11444,N_11380,N_11290);
nor U11445 (N_11445,N_11223,N_11257);
nand U11446 (N_11446,N_11382,N_11248);
and U11447 (N_11447,N_11389,N_11352);
nand U11448 (N_11448,N_11341,N_11282);
xor U11449 (N_11449,N_11293,N_11211);
nand U11450 (N_11450,N_11303,N_11235);
nor U11451 (N_11451,N_11278,N_11358);
xor U11452 (N_11452,N_11363,N_11281);
xor U11453 (N_11453,N_11232,N_11256);
or U11454 (N_11454,N_11391,N_11260);
xnor U11455 (N_11455,N_11342,N_11215);
xnor U11456 (N_11456,N_11393,N_11265);
xor U11457 (N_11457,N_11214,N_11285);
xnor U11458 (N_11458,N_11310,N_11329);
or U11459 (N_11459,N_11344,N_11346);
nand U11460 (N_11460,N_11350,N_11226);
nand U11461 (N_11461,N_11332,N_11328);
nand U11462 (N_11462,N_11384,N_11209);
nand U11463 (N_11463,N_11318,N_11297);
or U11464 (N_11464,N_11251,N_11304);
nand U11465 (N_11465,N_11200,N_11349);
nor U11466 (N_11466,N_11325,N_11216);
nand U11467 (N_11467,N_11336,N_11306);
xnor U11468 (N_11468,N_11334,N_11225);
and U11469 (N_11469,N_11314,N_11313);
or U11470 (N_11470,N_11390,N_11271);
xor U11471 (N_11471,N_11275,N_11320);
nor U11472 (N_11472,N_11250,N_11395);
or U11473 (N_11473,N_11233,N_11353);
or U11474 (N_11474,N_11230,N_11383);
and U11475 (N_11475,N_11302,N_11244);
and U11476 (N_11476,N_11217,N_11254);
nand U11477 (N_11477,N_11365,N_11242);
nor U11478 (N_11478,N_11378,N_11266);
and U11479 (N_11479,N_11207,N_11241);
and U11480 (N_11480,N_11300,N_11228);
and U11481 (N_11481,N_11262,N_11206);
nor U11482 (N_11482,N_11264,N_11321);
nor U11483 (N_11483,N_11367,N_11373);
nor U11484 (N_11484,N_11218,N_11291);
and U11485 (N_11485,N_11240,N_11331);
nand U11486 (N_11486,N_11219,N_11322);
or U11487 (N_11487,N_11370,N_11255);
and U11488 (N_11488,N_11247,N_11388);
xnor U11489 (N_11489,N_11295,N_11252);
nor U11490 (N_11490,N_11277,N_11345);
xor U11491 (N_11491,N_11348,N_11315);
nand U11492 (N_11492,N_11231,N_11287);
and U11493 (N_11493,N_11301,N_11372);
or U11494 (N_11494,N_11361,N_11396);
or U11495 (N_11495,N_11284,N_11286);
or U11496 (N_11496,N_11360,N_11268);
or U11497 (N_11497,N_11319,N_11227);
or U11498 (N_11498,N_11224,N_11246);
and U11499 (N_11499,N_11355,N_11238);
nor U11500 (N_11500,N_11327,N_11277);
nand U11501 (N_11501,N_11269,N_11209);
xor U11502 (N_11502,N_11380,N_11360);
nor U11503 (N_11503,N_11254,N_11298);
xor U11504 (N_11504,N_11386,N_11361);
xnor U11505 (N_11505,N_11322,N_11303);
or U11506 (N_11506,N_11308,N_11393);
nand U11507 (N_11507,N_11312,N_11258);
or U11508 (N_11508,N_11284,N_11298);
nand U11509 (N_11509,N_11368,N_11214);
xnor U11510 (N_11510,N_11319,N_11352);
nand U11511 (N_11511,N_11301,N_11341);
nand U11512 (N_11512,N_11295,N_11229);
or U11513 (N_11513,N_11268,N_11278);
xor U11514 (N_11514,N_11393,N_11287);
and U11515 (N_11515,N_11304,N_11298);
and U11516 (N_11516,N_11363,N_11243);
xor U11517 (N_11517,N_11388,N_11382);
and U11518 (N_11518,N_11343,N_11392);
nand U11519 (N_11519,N_11259,N_11294);
and U11520 (N_11520,N_11237,N_11369);
nand U11521 (N_11521,N_11339,N_11271);
nor U11522 (N_11522,N_11355,N_11316);
xor U11523 (N_11523,N_11224,N_11268);
or U11524 (N_11524,N_11342,N_11391);
xor U11525 (N_11525,N_11371,N_11378);
xnor U11526 (N_11526,N_11326,N_11343);
nand U11527 (N_11527,N_11312,N_11370);
nor U11528 (N_11528,N_11331,N_11314);
and U11529 (N_11529,N_11354,N_11293);
nor U11530 (N_11530,N_11352,N_11295);
nand U11531 (N_11531,N_11240,N_11317);
nor U11532 (N_11532,N_11271,N_11222);
nor U11533 (N_11533,N_11250,N_11326);
or U11534 (N_11534,N_11365,N_11328);
nor U11535 (N_11535,N_11265,N_11306);
nor U11536 (N_11536,N_11312,N_11271);
and U11537 (N_11537,N_11285,N_11274);
or U11538 (N_11538,N_11372,N_11370);
nand U11539 (N_11539,N_11355,N_11274);
xor U11540 (N_11540,N_11239,N_11286);
and U11541 (N_11541,N_11298,N_11378);
or U11542 (N_11542,N_11214,N_11258);
nor U11543 (N_11543,N_11335,N_11304);
or U11544 (N_11544,N_11302,N_11205);
xor U11545 (N_11545,N_11261,N_11343);
nand U11546 (N_11546,N_11327,N_11388);
or U11547 (N_11547,N_11338,N_11296);
nand U11548 (N_11548,N_11354,N_11246);
or U11549 (N_11549,N_11391,N_11210);
xnor U11550 (N_11550,N_11392,N_11251);
and U11551 (N_11551,N_11249,N_11251);
xor U11552 (N_11552,N_11253,N_11230);
and U11553 (N_11553,N_11276,N_11387);
nor U11554 (N_11554,N_11378,N_11207);
and U11555 (N_11555,N_11326,N_11202);
xnor U11556 (N_11556,N_11395,N_11294);
nor U11557 (N_11557,N_11239,N_11347);
nor U11558 (N_11558,N_11303,N_11336);
xor U11559 (N_11559,N_11291,N_11338);
and U11560 (N_11560,N_11362,N_11203);
and U11561 (N_11561,N_11325,N_11353);
and U11562 (N_11562,N_11367,N_11254);
xnor U11563 (N_11563,N_11376,N_11251);
nor U11564 (N_11564,N_11257,N_11378);
nor U11565 (N_11565,N_11382,N_11317);
and U11566 (N_11566,N_11307,N_11304);
and U11567 (N_11567,N_11277,N_11318);
and U11568 (N_11568,N_11277,N_11343);
nand U11569 (N_11569,N_11264,N_11208);
nand U11570 (N_11570,N_11227,N_11224);
or U11571 (N_11571,N_11352,N_11262);
xnor U11572 (N_11572,N_11284,N_11205);
or U11573 (N_11573,N_11269,N_11398);
or U11574 (N_11574,N_11301,N_11225);
and U11575 (N_11575,N_11353,N_11338);
xor U11576 (N_11576,N_11253,N_11218);
nor U11577 (N_11577,N_11370,N_11237);
nand U11578 (N_11578,N_11255,N_11312);
xnor U11579 (N_11579,N_11371,N_11235);
xnor U11580 (N_11580,N_11303,N_11382);
xnor U11581 (N_11581,N_11245,N_11340);
or U11582 (N_11582,N_11317,N_11337);
nor U11583 (N_11583,N_11382,N_11355);
and U11584 (N_11584,N_11241,N_11374);
nor U11585 (N_11585,N_11282,N_11365);
nand U11586 (N_11586,N_11217,N_11210);
nor U11587 (N_11587,N_11219,N_11252);
and U11588 (N_11588,N_11268,N_11242);
or U11589 (N_11589,N_11389,N_11319);
nor U11590 (N_11590,N_11349,N_11395);
nand U11591 (N_11591,N_11295,N_11245);
nor U11592 (N_11592,N_11229,N_11320);
and U11593 (N_11593,N_11359,N_11311);
nand U11594 (N_11594,N_11252,N_11277);
or U11595 (N_11595,N_11244,N_11386);
or U11596 (N_11596,N_11242,N_11234);
or U11597 (N_11597,N_11231,N_11326);
or U11598 (N_11598,N_11288,N_11287);
and U11599 (N_11599,N_11269,N_11394);
nand U11600 (N_11600,N_11505,N_11422);
or U11601 (N_11601,N_11461,N_11522);
nor U11602 (N_11602,N_11579,N_11587);
nor U11603 (N_11603,N_11431,N_11511);
nand U11604 (N_11604,N_11594,N_11451);
or U11605 (N_11605,N_11433,N_11529);
nand U11606 (N_11606,N_11557,N_11531);
nor U11607 (N_11607,N_11437,N_11490);
nand U11608 (N_11608,N_11464,N_11504);
or U11609 (N_11609,N_11542,N_11507);
and U11610 (N_11610,N_11537,N_11426);
or U11611 (N_11611,N_11552,N_11521);
nand U11612 (N_11612,N_11476,N_11446);
and U11613 (N_11613,N_11439,N_11584);
nor U11614 (N_11614,N_11427,N_11536);
and U11615 (N_11615,N_11517,N_11452);
nor U11616 (N_11616,N_11478,N_11496);
or U11617 (N_11617,N_11564,N_11487);
nor U11618 (N_11618,N_11534,N_11599);
and U11619 (N_11619,N_11486,N_11488);
and U11620 (N_11620,N_11567,N_11450);
and U11621 (N_11621,N_11449,N_11492);
or U11622 (N_11622,N_11489,N_11480);
nand U11623 (N_11623,N_11571,N_11458);
nor U11624 (N_11624,N_11498,N_11519);
nor U11625 (N_11625,N_11482,N_11565);
xnor U11626 (N_11626,N_11513,N_11506);
nand U11627 (N_11627,N_11589,N_11491);
xor U11628 (N_11628,N_11444,N_11595);
xor U11629 (N_11629,N_11548,N_11423);
and U11630 (N_11630,N_11479,N_11553);
nor U11631 (N_11631,N_11541,N_11575);
or U11632 (N_11632,N_11515,N_11429);
or U11633 (N_11633,N_11400,N_11471);
and U11634 (N_11634,N_11560,N_11483);
xor U11635 (N_11635,N_11583,N_11591);
and U11636 (N_11636,N_11481,N_11412);
nor U11637 (N_11637,N_11523,N_11550);
and U11638 (N_11638,N_11588,N_11445);
xnor U11639 (N_11639,N_11499,N_11405);
xor U11640 (N_11640,N_11554,N_11598);
or U11641 (N_11641,N_11475,N_11559);
and U11642 (N_11642,N_11474,N_11454);
xor U11643 (N_11643,N_11508,N_11545);
xor U11644 (N_11644,N_11572,N_11453);
nand U11645 (N_11645,N_11586,N_11593);
nor U11646 (N_11646,N_11447,N_11527);
and U11647 (N_11647,N_11404,N_11428);
nor U11648 (N_11648,N_11581,N_11477);
and U11649 (N_11649,N_11485,N_11555);
nand U11650 (N_11650,N_11528,N_11530);
or U11651 (N_11651,N_11424,N_11570);
nand U11652 (N_11652,N_11493,N_11409);
nor U11653 (N_11653,N_11585,N_11416);
and U11654 (N_11654,N_11503,N_11568);
and U11655 (N_11655,N_11561,N_11502);
and U11656 (N_11656,N_11500,N_11455);
nor U11657 (N_11657,N_11402,N_11540);
or U11658 (N_11658,N_11469,N_11543);
or U11659 (N_11659,N_11494,N_11401);
nand U11660 (N_11660,N_11547,N_11406);
nor U11661 (N_11661,N_11467,N_11563);
nand U11662 (N_11662,N_11518,N_11525);
xnor U11663 (N_11663,N_11435,N_11510);
or U11664 (N_11664,N_11425,N_11434);
nor U11665 (N_11665,N_11430,N_11463);
nor U11666 (N_11666,N_11442,N_11497);
or U11667 (N_11667,N_11440,N_11582);
or U11668 (N_11668,N_11438,N_11495);
nor U11669 (N_11669,N_11577,N_11443);
nor U11670 (N_11670,N_11512,N_11411);
or U11671 (N_11671,N_11516,N_11413);
and U11672 (N_11672,N_11408,N_11597);
nand U11673 (N_11673,N_11551,N_11470);
or U11674 (N_11674,N_11462,N_11417);
and U11675 (N_11675,N_11558,N_11466);
and U11676 (N_11676,N_11457,N_11468);
or U11677 (N_11677,N_11465,N_11472);
nand U11678 (N_11678,N_11420,N_11414);
nand U11679 (N_11679,N_11526,N_11460);
nand U11680 (N_11680,N_11592,N_11549);
and U11681 (N_11681,N_11448,N_11596);
nor U11682 (N_11682,N_11538,N_11441);
nor U11683 (N_11683,N_11418,N_11539);
and U11684 (N_11684,N_11459,N_11456);
nor U11685 (N_11685,N_11407,N_11514);
nand U11686 (N_11686,N_11436,N_11535);
nand U11687 (N_11687,N_11574,N_11576);
nand U11688 (N_11688,N_11524,N_11501);
xor U11689 (N_11689,N_11532,N_11421);
nor U11690 (N_11690,N_11410,N_11546);
nor U11691 (N_11691,N_11432,N_11473);
nor U11692 (N_11692,N_11509,N_11403);
and U11693 (N_11693,N_11533,N_11580);
xor U11694 (N_11694,N_11415,N_11556);
nand U11695 (N_11695,N_11544,N_11590);
nand U11696 (N_11696,N_11562,N_11573);
nand U11697 (N_11697,N_11578,N_11566);
nand U11698 (N_11698,N_11520,N_11419);
xnor U11699 (N_11699,N_11484,N_11569);
nor U11700 (N_11700,N_11495,N_11563);
and U11701 (N_11701,N_11588,N_11472);
and U11702 (N_11702,N_11567,N_11562);
nand U11703 (N_11703,N_11543,N_11537);
xor U11704 (N_11704,N_11413,N_11534);
or U11705 (N_11705,N_11505,N_11467);
xnor U11706 (N_11706,N_11512,N_11438);
or U11707 (N_11707,N_11439,N_11415);
or U11708 (N_11708,N_11576,N_11429);
or U11709 (N_11709,N_11543,N_11459);
or U11710 (N_11710,N_11445,N_11424);
and U11711 (N_11711,N_11484,N_11464);
xnor U11712 (N_11712,N_11451,N_11422);
xnor U11713 (N_11713,N_11493,N_11427);
or U11714 (N_11714,N_11503,N_11509);
nand U11715 (N_11715,N_11464,N_11525);
and U11716 (N_11716,N_11479,N_11402);
nand U11717 (N_11717,N_11503,N_11485);
and U11718 (N_11718,N_11486,N_11438);
nand U11719 (N_11719,N_11431,N_11512);
nand U11720 (N_11720,N_11512,N_11433);
and U11721 (N_11721,N_11492,N_11480);
xnor U11722 (N_11722,N_11537,N_11484);
or U11723 (N_11723,N_11557,N_11507);
xnor U11724 (N_11724,N_11457,N_11565);
nor U11725 (N_11725,N_11450,N_11570);
xor U11726 (N_11726,N_11497,N_11429);
nand U11727 (N_11727,N_11586,N_11493);
xor U11728 (N_11728,N_11451,N_11417);
nor U11729 (N_11729,N_11412,N_11523);
or U11730 (N_11730,N_11510,N_11500);
nand U11731 (N_11731,N_11587,N_11564);
nand U11732 (N_11732,N_11529,N_11476);
xor U11733 (N_11733,N_11446,N_11455);
nor U11734 (N_11734,N_11456,N_11465);
or U11735 (N_11735,N_11441,N_11505);
xor U11736 (N_11736,N_11530,N_11407);
nand U11737 (N_11737,N_11493,N_11452);
nand U11738 (N_11738,N_11427,N_11483);
xor U11739 (N_11739,N_11467,N_11405);
and U11740 (N_11740,N_11492,N_11587);
and U11741 (N_11741,N_11557,N_11425);
and U11742 (N_11742,N_11519,N_11492);
xnor U11743 (N_11743,N_11466,N_11475);
xnor U11744 (N_11744,N_11484,N_11405);
or U11745 (N_11745,N_11423,N_11441);
or U11746 (N_11746,N_11441,N_11439);
nand U11747 (N_11747,N_11402,N_11537);
nor U11748 (N_11748,N_11519,N_11460);
nor U11749 (N_11749,N_11422,N_11585);
nand U11750 (N_11750,N_11525,N_11524);
nor U11751 (N_11751,N_11499,N_11540);
xor U11752 (N_11752,N_11518,N_11413);
or U11753 (N_11753,N_11534,N_11467);
or U11754 (N_11754,N_11451,N_11449);
nor U11755 (N_11755,N_11556,N_11448);
and U11756 (N_11756,N_11573,N_11537);
nand U11757 (N_11757,N_11561,N_11508);
and U11758 (N_11758,N_11452,N_11526);
xnor U11759 (N_11759,N_11523,N_11572);
or U11760 (N_11760,N_11582,N_11434);
and U11761 (N_11761,N_11450,N_11485);
or U11762 (N_11762,N_11535,N_11474);
nand U11763 (N_11763,N_11455,N_11512);
nor U11764 (N_11764,N_11513,N_11510);
nand U11765 (N_11765,N_11435,N_11483);
xnor U11766 (N_11766,N_11569,N_11521);
nand U11767 (N_11767,N_11560,N_11574);
xor U11768 (N_11768,N_11570,N_11428);
and U11769 (N_11769,N_11511,N_11442);
nor U11770 (N_11770,N_11411,N_11480);
xnor U11771 (N_11771,N_11575,N_11501);
and U11772 (N_11772,N_11584,N_11461);
or U11773 (N_11773,N_11402,N_11410);
nor U11774 (N_11774,N_11561,N_11568);
nor U11775 (N_11775,N_11539,N_11477);
nor U11776 (N_11776,N_11577,N_11424);
or U11777 (N_11777,N_11557,N_11565);
xnor U11778 (N_11778,N_11421,N_11505);
or U11779 (N_11779,N_11421,N_11563);
nor U11780 (N_11780,N_11537,N_11526);
xnor U11781 (N_11781,N_11510,N_11533);
and U11782 (N_11782,N_11515,N_11475);
or U11783 (N_11783,N_11464,N_11416);
and U11784 (N_11784,N_11571,N_11438);
and U11785 (N_11785,N_11473,N_11533);
nand U11786 (N_11786,N_11573,N_11435);
or U11787 (N_11787,N_11515,N_11435);
nand U11788 (N_11788,N_11520,N_11437);
nor U11789 (N_11789,N_11425,N_11477);
xnor U11790 (N_11790,N_11425,N_11551);
nand U11791 (N_11791,N_11561,N_11494);
nand U11792 (N_11792,N_11562,N_11543);
nor U11793 (N_11793,N_11425,N_11432);
or U11794 (N_11794,N_11514,N_11456);
xnor U11795 (N_11795,N_11588,N_11431);
xnor U11796 (N_11796,N_11579,N_11542);
or U11797 (N_11797,N_11470,N_11596);
nand U11798 (N_11798,N_11566,N_11401);
xor U11799 (N_11799,N_11411,N_11518);
nor U11800 (N_11800,N_11701,N_11688);
or U11801 (N_11801,N_11696,N_11682);
or U11802 (N_11802,N_11675,N_11708);
xnor U11803 (N_11803,N_11799,N_11641);
nor U11804 (N_11804,N_11664,N_11668);
nand U11805 (N_11805,N_11703,N_11710);
or U11806 (N_11806,N_11709,N_11705);
nand U11807 (N_11807,N_11784,N_11736);
or U11808 (N_11808,N_11609,N_11734);
and U11809 (N_11809,N_11750,N_11731);
nand U11810 (N_11810,N_11671,N_11769);
nor U11811 (N_11811,N_11630,N_11713);
nor U11812 (N_11812,N_11667,N_11771);
and U11813 (N_11813,N_11794,N_11637);
and U11814 (N_11814,N_11715,N_11690);
xnor U11815 (N_11815,N_11720,N_11770);
nand U11816 (N_11816,N_11610,N_11792);
nand U11817 (N_11817,N_11748,N_11790);
nand U11818 (N_11818,N_11725,N_11718);
xor U11819 (N_11819,N_11670,N_11774);
nor U11820 (N_11820,N_11658,N_11782);
xor U11821 (N_11821,N_11741,N_11798);
xnor U11822 (N_11822,N_11661,N_11699);
xor U11823 (N_11823,N_11758,N_11729);
nor U11824 (N_11824,N_11751,N_11623);
or U11825 (N_11825,N_11716,N_11754);
nand U11826 (N_11826,N_11689,N_11753);
nand U11827 (N_11827,N_11732,N_11659);
nor U11828 (N_11828,N_11706,N_11644);
and U11829 (N_11829,N_11677,N_11698);
or U11830 (N_11830,N_11702,N_11605);
or U11831 (N_11831,N_11793,N_11607);
nand U11832 (N_11832,N_11622,N_11612);
nand U11833 (N_11833,N_11787,N_11645);
nand U11834 (N_11834,N_11763,N_11617);
nor U11835 (N_11835,N_11719,N_11765);
nor U11836 (N_11836,N_11752,N_11743);
nand U11837 (N_11837,N_11723,N_11797);
nor U11838 (N_11838,N_11744,N_11600);
and U11839 (N_11839,N_11683,N_11693);
and U11840 (N_11840,N_11783,N_11779);
nor U11841 (N_11841,N_11738,N_11767);
or U11842 (N_11842,N_11788,N_11614);
or U11843 (N_11843,N_11652,N_11733);
and U11844 (N_11844,N_11691,N_11674);
xnor U11845 (N_11845,N_11714,N_11633);
or U11846 (N_11846,N_11632,N_11745);
nand U11847 (N_11847,N_11649,N_11755);
or U11848 (N_11848,N_11781,N_11672);
xnor U11849 (N_11849,N_11640,N_11796);
and U11850 (N_11850,N_11786,N_11795);
xor U11851 (N_11851,N_11616,N_11618);
xor U11852 (N_11852,N_11648,N_11681);
and U11853 (N_11853,N_11651,N_11727);
nor U11854 (N_11854,N_11761,N_11739);
xnor U11855 (N_11855,N_11634,N_11757);
and U11856 (N_11856,N_11620,N_11773);
or U11857 (N_11857,N_11728,N_11747);
nor U11858 (N_11858,N_11695,N_11613);
and U11859 (N_11859,N_11759,N_11687);
or U11860 (N_11860,N_11791,N_11766);
nor U11861 (N_11861,N_11602,N_11657);
xnor U11862 (N_11862,N_11700,N_11722);
or U11863 (N_11863,N_11680,N_11603);
nor U11864 (N_11864,N_11746,N_11646);
nor U11865 (N_11865,N_11772,N_11717);
xnor U11866 (N_11866,N_11712,N_11704);
xnor U11867 (N_11867,N_11666,N_11673);
nand U11868 (N_11868,N_11656,N_11762);
and U11869 (N_11869,N_11789,N_11627);
nor U11870 (N_11870,N_11721,N_11685);
nand U11871 (N_11871,N_11760,N_11621);
and U11872 (N_11872,N_11697,N_11631);
and U11873 (N_11873,N_11647,N_11684);
or U11874 (N_11874,N_11749,N_11628);
nand U11875 (N_11875,N_11692,N_11676);
xor U11876 (N_11876,N_11669,N_11653);
xor U11877 (N_11877,N_11624,N_11778);
xor U11878 (N_11878,N_11665,N_11780);
nand U11879 (N_11879,N_11730,N_11678);
xor U11880 (N_11880,N_11663,N_11615);
nand U11881 (N_11881,N_11635,N_11606);
nor U11882 (N_11882,N_11650,N_11662);
nand U11883 (N_11883,N_11654,N_11601);
nor U11884 (N_11884,N_11777,N_11636);
or U11885 (N_11885,N_11686,N_11619);
or U11886 (N_11886,N_11742,N_11629);
xnor U11887 (N_11887,N_11604,N_11611);
or U11888 (N_11888,N_11639,N_11694);
and U11889 (N_11889,N_11764,N_11785);
nand U11890 (N_11890,N_11642,N_11626);
and U11891 (N_11891,N_11643,N_11776);
nor U11892 (N_11892,N_11740,N_11737);
nor U11893 (N_11893,N_11724,N_11768);
and U11894 (N_11894,N_11625,N_11707);
nor U11895 (N_11895,N_11655,N_11775);
nor U11896 (N_11896,N_11735,N_11726);
xnor U11897 (N_11897,N_11679,N_11638);
nand U11898 (N_11898,N_11711,N_11660);
xor U11899 (N_11899,N_11608,N_11756);
nor U11900 (N_11900,N_11631,N_11603);
nor U11901 (N_11901,N_11745,N_11621);
nor U11902 (N_11902,N_11664,N_11717);
nand U11903 (N_11903,N_11673,N_11675);
nand U11904 (N_11904,N_11627,N_11770);
xnor U11905 (N_11905,N_11602,N_11766);
or U11906 (N_11906,N_11799,N_11600);
nor U11907 (N_11907,N_11730,N_11622);
and U11908 (N_11908,N_11656,N_11713);
nor U11909 (N_11909,N_11614,N_11667);
nand U11910 (N_11910,N_11612,N_11688);
xor U11911 (N_11911,N_11704,N_11691);
and U11912 (N_11912,N_11773,N_11749);
or U11913 (N_11913,N_11781,N_11684);
nor U11914 (N_11914,N_11650,N_11762);
and U11915 (N_11915,N_11613,N_11703);
xnor U11916 (N_11916,N_11738,N_11671);
and U11917 (N_11917,N_11740,N_11720);
nand U11918 (N_11918,N_11676,N_11661);
xnor U11919 (N_11919,N_11725,N_11765);
xor U11920 (N_11920,N_11631,N_11777);
nand U11921 (N_11921,N_11729,N_11771);
and U11922 (N_11922,N_11617,N_11696);
nor U11923 (N_11923,N_11730,N_11725);
nand U11924 (N_11924,N_11652,N_11743);
nand U11925 (N_11925,N_11689,N_11621);
or U11926 (N_11926,N_11627,N_11636);
xnor U11927 (N_11927,N_11789,N_11613);
xor U11928 (N_11928,N_11615,N_11631);
nand U11929 (N_11929,N_11730,N_11663);
nand U11930 (N_11930,N_11636,N_11683);
nor U11931 (N_11931,N_11653,N_11685);
and U11932 (N_11932,N_11709,N_11608);
or U11933 (N_11933,N_11655,N_11770);
or U11934 (N_11934,N_11788,N_11791);
and U11935 (N_11935,N_11703,N_11757);
xor U11936 (N_11936,N_11667,N_11627);
nor U11937 (N_11937,N_11712,N_11648);
nand U11938 (N_11938,N_11740,N_11634);
nor U11939 (N_11939,N_11790,N_11782);
and U11940 (N_11940,N_11613,N_11746);
nor U11941 (N_11941,N_11707,N_11691);
nor U11942 (N_11942,N_11661,N_11741);
nand U11943 (N_11943,N_11650,N_11782);
xnor U11944 (N_11944,N_11693,N_11665);
nand U11945 (N_11945,N_11656,N_11698);
nor U11946 (N_11946,N_11774,N_11657);
nor U11947 (N_11947,N_11652,N_11689);
nor U11948 (N_11948,N_11768,N_11710);
or U11949 (N_11949,N_11752,N_11652);
xor U11950 (N_11950,N_11625,N_11797);
and U11951 (N_11951,N_11648,N_11628);
nor U11952 (N_11952,N_11608,N_11780);
nor U11953 (N_11953,N_11719,N_11720);
xor U11954 (N_11954,N_11697,N_11618);
xnor U11955 (N_11955,N_11618,N_11796);
xor U11956 (N_11956,N_11701,N_11686);
xor U11957 (N_11957,N_11782,N_11742);
or U11958 (N_11958,N_11797,N_11757);
or U11959 (N_11959,N_11634,N_11763);
nand U11960 (N_11960,N_11653,N_11754);
xor U11961 (N_11961,N_11667,N_11741);
or U11962 (N_11962,N_11635,N_11691);
and U11963 (N_11963,N_11747,N_11738);
and U11964 (N_11964,N_11725,N_11780);
or U11965 (N_11965,N_11778,N_11788);
and U11966 (N_11966,N_11742,N_11646);
nor U11967 (N_11967,N_11632,N_11623);
or U11968 (N_11968,N_11670,N_11643);
nor U11969 (N_11969,N_11691,N_11609);
nand U11970 (N_11970,N_11783,N_11603);
nor U11971 (N_11971,N_11700,N_11738);
and U11972 (N_11972,N_11728,N_11758);
nor U11973 (N_11973,N_11751,N_11790);
nor U11974 (N_11974,N_11635,N_11772);
xnor U11975 (N_11975,N_11718,N_11736);
and U11976 (N_11976,N_11629,N_11703);
nor U11977 (N_11977,N_11635,N_11674);
or U11978 (N_11978,N_11669,N_11757);
nand U11979 (N_11979,N_11627,N_11766);
nor U11980 (N_11980,N_11796,N_11632);
and U11981 (N_11981,N_11663,N_11611);
nor U11982 (N_11982,N_11643,N_11615);
nand U11983 (N_11983,N_11703,N_11667);
or U11984 (N_11984,N_11672,N_11779);
xor U11985 (N_11985,N_11607,N_11704);
nand U11986 (N_11986,N_11735,N_11661);
nor U11987 (N_11987,N_11759,N_11792);
and U11988 (N_11988,N_11727,N_11653);
nand U11989 (N_11989,N_11632,N_11708);
nor U11990 (N_11990,N_11653,N_11777);
and U11991 (N_11991,N_11731,N_11619);
nor U11992 (N_11992,N_11795,N_11645);
nor U11993 (N_11993,N_11787,N_11735);
xor U11994 (N_11994,N_11726,N_11756);
nand U11995 (N_11995,N_11606,N_11657);
and U11996 (N_11996,N_11736,N_11620);
nand U11997 (N_11997,N_11641,N_11774);
nand U11998 (N_11998,N_11797,N_11754);
xor U11999 (N_11999,N_11781,N_11783);
or U12000 (N_12000,N_11940,N_11904);
and U12001 (N_12001,N_11988,N_11960);
xor U12002 (N_12002,N_11920,N_11897);
nor U12003 (N_12003,N_11812,N_11827);
and U12004 (N_12004,N_11882,N_11978);
nand U12005 (N_12005,N_11905,N_11888);
and U12006 (N_12006,N_11866,N_11835);
or U12007 (N_12007,N_11895,N_11820);
and U12008 (N_12008,N_11911,N_11913);
nand U12009 (N_12009,N_11964,N_11823);
xor U12010 (N_12010,N_11957,N_11998);
and U12011 (N_12011,N_11894,N_11965);
xnor U12012 (N_12012,N_11868,N_11941);
or U12013 (N_12013,N_11831,N_11826);
nor U12014 (N_12014,N_11893,N_11805);
or U12015 (N_12015,N_11839,N_11983);
and U12016 (N_12016,N_11803,N_11930);
nor U12017 (N_12017,N_11929,N_11945);
nand U12018 (N_12018,N_11942,N_11900);
nor U12019 (N_12019,N_11944,N_11834);
nor U12020 (N_12020,N_11990,N_11809);
nor U12021 (N_12021,N_11921,N_11956);
xnor U12022 (N_12022,N_11914,N_11800);
xor U12023 (N_12023,N_11981,N_11973);
nand U12024 (N_12024,N_11959,N_11976);
nand U12025 (N_12025,N_11885,N_11898);
or U12026 (N_12026,N_11907,N_11933);
and U12027 (N_12027,N_11931,N_11849);
and U12028 (N_12028,N_11838,N_11875);
nor U12029 (N_12029,N_11985,N_11934);
nand U12030 (N_12030,N_11910,N_11979);
nand U12031 (N_12031,N_11887,N_11891);
nand U12032 (N_12032,N_11828,N_11922);
nor U12033 (N_12033,N_11917,N_11879);
nand U12034 (N_12034,N_11819,N_11952);
or U12035 (N_12035,N_11851,N_11840);
xnor U12036 (N_12036,N_11880,N_11858);
nand U12037 (N_12037,N_11939,N_11918);
nor U12038 (N_12038,N_11912,N_11899);
or U12039 (N_12039,N_11810,N_11909);
xnor U12040 (N_12040,N_11971,N_11916);
and U12041 (N_12041,N_11870,N_11968);
nand U12042 (N_12042,N_11989,N_11995);
xnor U12043 (N_12043,N_11861,N_11865);
nand U12044 (N_12044,N_11987,N_11873);
nor U12045 (N_12045,N_11984,N_11813);
nand U12046 (N_12046,N_11825,N_11932);
xnor U12047 (N_12047,N_11975,N_11871);
nor U12048 (N_12048,N_11997,N_11816);
xnor U12049 (N_12049,N_11853,N_11951);
nor U12050 (N_12050,N_11841,N_11806);
or U12051 (N_12051,N_11935,N_11993);
and U12052 (N_12052,N_11923,N_11906);
or U12053 (N_12053,N_11992,N_11850);
and U12054 (N_12054,N_11902,N_11947);
nor U12055 (N_12055,N_11948,N_11830);
and U12056 (N_12056,N_11829,N_11908);
nor U12057 (N_12057,N_11963,N_11889);
and U12058 (N_12058,N_11986,N_11878);
and U12059 (N_12059,N_11901,N_11802);
and U12060 (N_12060,N_11845,N_11807);
or U12061 (N_12061,N_11846,N_11822);
or U12062 (N_12062,N_11996,N_11982);
xor U12063 (N_12063,N_11974,N_11936);
xor U12064 (N_12064,N_11950,N_11869);
xnor U12065 (N_12065,N_11867,N_11970);
xor U12066 (N_12066,N_11877,N_11832);
nor U12067 (N_12067,N_11833,N_11969);
nand U12068 (N_12068,N_11967,N_11915);
xnor U12069 (N_12069,N_11972,N_11854);
xnor U12070 (N_12070,N_11883,N_11876);
nor U12071 (N_12071,N_11977,N_11818);
or U12072 (N_12072,N_11804,N_11954);
nor U12073 (N_12073,N_11860,N_11926);
nand U12074 (N_12074,N_11814,N_11863);
or U12075 (N_12075,N_11815,N_11928);
nand U12076 (N_12076,N_11844,N_11919);
or U12077 (N_12077,N_11943,N_11847);
or U12078 (N_12078,N_11842,N_11859);
nor U12079 (N_12079,N_11938,N_11925);
nor U12080 (N_12080,N_11949,N_11801);
xnor U12081 (N_12081,N_11836,N_11896);
or U12082 (N_12082,N_11994,N_11980);
nor U12083 (N_12083,N_11862,N_11937);
xnor U12084 (N_12084,N_11961,N_11817);
and U12085 (N_12085,N_11892,N_11955);
or U12086 (N_12086,N_11874,N_11962);
and U12087 (N_12087,N_11890,N_11884);
xnor U12088 (N_12088,N_11864,N_11966);
nor U12089 (N_12089,N_11855,N_11886);
nor U12090 (N_12090,N_11872,N_11811);
xnor U12091 (N_12091,N_11857,N_11848);
xor U12092 (N_12092,N_11953,N_11821);
nand U12093 (N_12093,N_11852,N_11903);
nand U12094 (N_12094,N_11856,N_11881);
nor U12095 (N_12095,N_11837,N_11958);
nand U12096 (N_12096,N_11843,N_11927);
xor U12097 (N_12097,N_11824,N_11808);
nand U12098 (N_12098,N_11946,N_11999);
xnor U12099 (N_12099,N_11991,N_11924);
nand U12100 (N_12100,N_11823,N_11839);
nor U12101 (N_12101,N_11997,N_11805);
nand U12102 (N_12102,N_11968,N_11906);
xor U12103 (N_12103,N_11810,N_11962);
nor U12104 (N_12104,N_11969,N_11981);
xnor U12105 (N_12105,N_11803,N_11929);
and U12106 (N_12106,N_11975,N_11886);
or U12107 (N_12107,N_11831,N_11988);
and U12108 (N_12108,N_11913,N_11814);
and U12109 (N_12109,N_11994,N_11951);
nor U12110 (N_12110,N_11880,N_11994);
or U12111 (N_12111,N_11983,N_11868);
nor U12112 (N_12112,N_11907,N_11838);
nand U12113 (N_12113,N_11883,N_11961);
and U12114 (N_12114,N_11909,N_11831);
or U12115 (N_12115,N_11802,N_11884);
and U12116 (N_12116,N_11960,N_11842);
nand U12117 (N_12117,N_11901,N_11827);
nand U12118 (N_12118,N_11873,N_11899);
and U12119 (N_12119,N_11868,N_11874);
xor U12120 (N_12120,N_11893,N_11834);
or U12121 (N_12121,N_11923,N_11891);
and U12122 (N_12122,N_11955,N_11950);
or U12123 (N_12123,N_11878,N_11936);
and U12124 (N_12124,N_11879,N_11800);
and U12125 (N_12125,N_11869,N_11986);
nor U12126 (N_12126,N_11850,N_11885);
xnor U12127 (N_12127,N_11875,N_11967);
or U12128 (N_12128,N_11972,N_11970);
and U12129 (N_12129,N_11887,N_11944);
nor U12130 (N_12130,N_11828,N_11995);
or U12131 (N_12131,N_11989,N_11899);
or U12132 (N_12132,N_11852,N_11851);
nand U12133 (N_12133,N_11929,N_11988);
nand U12134 (N_12134,N_11801,N_11942);
nand U12135 (N_12135,N_11838,N_11846);
nor U12136 (N_12136,N_11909,N_11806);
nand U12137 (N_12137,N_11989,N_11858);
and U12138 (N_12138,N_11951,N_11845);
nand U12139 (N_12139,N_11999,N_11958);
xnor U12140 (N_12140,N_11854,N_11955);
xnor U12141 (N_12141,N_11976,N_11885);
xnor U12142 (N_12142,N_11850,N_11995);
and U12143 (N_12143,N_11843,N_11847);
xnor U12144 (N_12144,N_11965,N_11877);
nand U12145 (N_12145,N_11926,N_11890);
xor U12146 (N_12146,N_11937,N_11838);
nor U12147 (N_12147,N_11822,N_11900);
nor U12148 (N_12148,N_11882,N_11915);
xnor U12149 (N_12149,N_11847,N_11842);
or U12150 (N_12150,N_11880,N_11850);
and U12151 (N_12151,N_11803,N_11925);
and U12152 (N_12152,N_11836,N_11958);
xnor U12153 (N_12153,N_11993,N_11969);
nor U12154 (N_12154,N_11830,N_11951);
nand U12155 (N_12155,N_11882,N_11813);
xnor U12156 (N_12156,N_11828,N_11809);
or U12157 (N_12157,N_11946,N_11821);
and U12158 (N_12158,N_11889,N_11973);
nor U12159 (N_12159,N_11841,N_11816);
nor U12160 (N_12160,N_11991,N_11805);
nand U12161 (N_12161,N_11824,N_11905);
and U12162 (N_12162,N_11901,N_11869);
xor U12163 (N_12163,N_11869,N_11902);
nor U12164 (N_12164,N_11878,N_11844);
or U12165 (N_12165,N_11881,N_11826);
nor U12166 (N_12166,N_11993,N_11800);
or U12167 (N_12167,N_11998,N_11991);
xnor U12168 (N_12168,N_11921,N_11959);
or U12169 (N_12169,N_11809,N_11998);
nor U12170 (N_12170,N_11929,N_11987);
nand U12171 (N_12171,N_11943,N_11842);
nand U12172 (N_12172,N_11978,N_11922);
or U12173 (N_12173,N_11921,N_11929);
and U12174 (N_12174,N_11806,N_11997);
or U12175 (N_12175,N_11922,N_11826);
or U12176 (N_12176,N_11958,N_11969);
and U12177 (N_12177,N_11995,N_11999);
nor U12178 (N_12178,N_11867,N_11933);
nor U12179 (N_12179,N_11897,N_11819);
and U12180 (N_12180,N_11913,N_11847);
xnor U12181 (N_12181,N_11963,N_11920);
nor U12182 (N_12182,N_11879,N_11988);
xor U12183 (N_12183,N_11967,N_11903);
nor U12184 (N_12184,N_11967,N_11832);
or U12185 (N_12185,N_11913,N_11920);
or U12186 (N_12186,N_11936,N_11922);
nor U12187 (N_12187,N_11952,N_11982);
nor U12188 (N_12188,N_11933,N_11955);
and U12189 (N_12189,N_11984,N_11879);
nand U12190 (N_12190,N_11840,N_11905);
nor U12191 (N_12191,N_11838,N_11969);
and U12192 (N_12192,N_11816,N_11873);
and U12193 (N_12193,N_11964,N_11976);
xnor U12194 (N_12194,N_11812,N_11879);
xor U12195 (N_12195,N_11916,N_11847);
and U12196 (N_12196,N_11829,N_11960);
or U12197 (N_12197,N_11802,N_11942);
and U12198 (N_12198,N_11805,N_11885);
nor U12199 (N_12199,N_11994,N_11984);
or U12200 (N_12200,N_12198,N_12183);
xnor U12201 (N_12201,N_12018,N_12151);
nand U12202 (N_12202,N_12037,N_12009);
nor U12203 (N_12203,N_12008,N_12094);
nand U12204 (N_12204,N_12015,N_12146);
or U12205 (N_12205,N_12049,N_12058);
or U12206 (N_12206,N_12010,N_12084);
or U12207 (N_12207,N_12180,N_12141);
xor U12208 (N_12208,N_12033,N_12078);
or U12209 (N_12209,N_12133,N_12056);
xor U12210 (N_12210,N_12095,N_12112);
nand U12211 (N_12211,N_12072,N_12155);
xor U12212 (N_12212,N_12177,N_12070);
and U12213 (N_12213,N_12006,N_12165);
nor U12214 (N_12214,N_12027,N_12069);
nor U12215 (N_12215,N_12127,N_12130);
or U12216 (N_12216,N_12044,N_12132);
and U12217 (N_12217,N_12040,N_12060);
xnor U12218 (N_12218,N_12175,N_12052);
or U12219 (N_12219,N_12091,N_12189);
or U12220 (N_12220,N_12039,N_12184);
xnor U12221 (N_12221,N_12107,N_12114);
xor U12222 (N_12222,N_12089,N_12170);
nor U12223 (N_12223,N_12081,N_12195);
nor U12224 (N_12224,N_12187,N_12048);
and U12225 (N_12225,N_12000,N_12092);
nand U12226 (N_12226,N_12131,N_12123);
nor U12227 (N_12227,N_12079,N_12128);
nor U12228 (N_12228,N_12088,N_12190);
nor U12229 (N_12229,N_12042,N_12164);
and U12230 (N_12230,N_12014,N_12090);
or U12231 (N_12231,N_12087,N_12113);
and U12232 (N_12232,N_12075,N_12016);
nand U12233 (N_12233,N_12102,N_12191);
xnor U12234 (N_12234,N_12098,N_12086);
or U12235 (N_12235,N_12196,N_12082);
and U12236 (N_12236,N_12176,N_12122);
xor U12237 (N_12237,N_12111,N_12197);
and U12238 (N_12238,N_12154,N_12173);
nand U12239 (N_12239,N_12101,N_12105);
or U12240 (N_12240,N_12030,N_12029);
nor U12241 (N_12241,N_12172,N_12021);
nor U12242 (N_12242,N_12194,N_12137);
nand U12243 (N_12243,N_12003,N_12062);
or U12244 (N_12244,N_12013,N_12077);
and U12245 (N_12245,N_12163,N_12119);
nand U12246 (N_12246,N_12053,N_12011);
nand U12247 (N_12247,N_12007,N_12036);
nand U12248 (N_12248,N_12032,N_12004);
or U12249 (N_12249,N_12152,N_12142);
nand U12250 (N_12250,N_12117,N_12147);
or U12251 (N_12251,N_12038,N_12020);
or U12252 (N_12252,N_12073,N_12076);
nand U12253 (N_12253,N_12185,N_12025);
xnor U12254 (N_12254,N_12182,N_12093);
and U12255 (N_12255,N_12178,N_12193);
or U12256 (N_12256,N_12167,N_12066);
nor U12257 (N_12257,N_12047,N_12083);
nor U12258 (N_12258,N_12012,N_12024);
and U12259 (N_12259,N_12041,N_12067);
and U12260 (N_12260,N_12174,N_12157);
nand U12261 (N_12261,N_12005,N_12134);
xnor U12262 (N_12262,N_12055,N_12192);
xnor U12263 (N_12263,N_12168,N_12103);
and U12264 (N_12264,N_12166,N_12068);
nand U12265 (N_12265,N_12023,N_12153);
xnor U12266 (N_12266,N_12045,N_12054);
nand U12267 (N_12267,N_12071,N_12138);
and U12268 (N_12268,N_12121,N_12001);
xor U12269 (N_12269,N_12050,N_12063);
and U12270 (N_12270,N_12085,N_12097);
and U12271 (N_12271,N_12125,N_12135);
nand U12272 (N_12272,N_12149,N_12145);
nand U12273 (N_12273,N_12118,N_12179);
or U12274 (N_12274,N_12096,N_12099);
nor U12275 (N_12275,N_12126,N_12028);
xor U12276 (N_12276,N_12169,N_12136);
and U12277 (N_12277,N_12162,N_12019);
xnor U12278 (N_12278,N_12057,N_12116);
and U12279 (N_12279,N_12104,N_12017);
or U12280 (N_12280,N_12031,N_12108);
and U12281 (N_12281,N_12158,N_12188);
nor U12282 (N_12282,N_12161,N_12043);
xnor U12283 (N_12283,N_12159,N_12144);
and U12284 (N_12284,N_12100,N_12065);
nand U12285 (N_12285,N_12059,N_12022);
and U12286 (N_12286,N_12034,N_12140);
nand U12287 (N_12287,N_12120,N_12106);
nand U12288 (N_12288,N_12199,N_12110);
xor U12289 (N_12289,N_12171,N_12026);
nor U12290 (N_12290,N_12002,N_12160);
nand U12291 (N_12291,N_12074,N_12051);
nand U12292 (N_12292,N_12186,N_12064);
or U12293 (N_12293,N_12148,N_12143);
or U12294 (N_12294,N_12115,N_12109);
xnor U12295 (N_12295,N_12124,N_12181);
xor U12296 (N_12296,N_12046,N_12156);
xor U12297 (N_12297,N_12080,N_12150);
xnor U12298 (N_12298,N_12129,N_12139);
xor U12299 (N_12299,N_12035,N_12061);
or U12300 (N_12300,N_12117,N_12193);
nor U12301 (N_12301,N_12190,N_12082);
xor U12302 (N_12302,N_12080,N_12192);
nor U12303 (N_12303,N_12170,N_12182);
nand U12304 (N_12304,N_12195,N_12042);
xor U12305 (N_12305,N_12034,N_12165);
nand U12306 (N_12306,N_12086,N_12070);
and U12307 (N_12307,N_12179,N_12106);
or U12308 (N_12308,N_12171,N_12021);
or U12309 (N_12309,N_12172,N_12114);
and U12310 (N_12310,N_12088,N_12034);
or U12311 (N_12311,N_12101,N_12129);
or U12312 (N_12312,N_12121,N_12058);
or U12313 (N_12313,N_12181,N_12135);
or U12314 (N_12314,N_12107,N_12137);
nor U12315 (N_12315,N_12091,N_12043);
and U12316 (N_12316,N_12121,N_12112);
or U12317 (N_12317,N_12165,N_12040);
nor U12318 (N_12318,N_12064,N_12097);
xnor U12319 (N_12319,N_12080,N_12165);
xnor U12320 (N_12320,N_12140,N_12192);
xnor U12321 (N_12321,N_12166,N_12030);
and U12322 (N_12322,N_12136,N_12078);
and U12323 (N_12323,N_12081,N_12065);
and U12324 (N_12324,N_12046,N_12037);
and U12325 (N_12325,N_12002,N_12053);
nor U12326 (N_12326,N_12125,N_12104);
xnor U12327 (N_12327,N_12012,N_12174);
and U12328 (N_12328,N_12033,N_12064);
nor U12329 (N_12329,N_12124,N_12074);
nand U12330 (N_12330,N_12077,N_12137);
and U12331 (N_12331,N_12155,N_12106);
or U12332 (N_12332,N_12101,N_12026);
or U12333 (N_12333,N_12136,N_12139);
nand U12334 (N_12334,N_12002,N_12025);
xor U12335 (N_12335,N_12025,N_12014);
or U12336 (N_12336,N_12181,N_12161);
xor U12337 (N_12337,N_12049,N_12180);
or U12338 (N_12338,N_12000,N_12066);
nor U12339 (N_12339,N_12023,N_12078);
and U12340 (N_12340,N_12113,N_12016);
and U12341 (N_12341,N_12159,N_12193);
nand U12342 (N_12342,N_12174,N_12016);
xor U12343 (N_12343,N_12051,N_12108);
nand U12344 (N_12344,N_12068,N_12165);
nand U12345 (N_12345,N_12005,N_12033);
nor U12346 (N_12346,N_12107,N_12038);
nand U12347 (N_12347,N_12011,N_12131);
xnor U12348 (N_12348,N_12049,N_12102);
or U12349 (N_12349,N_12014,N_12127);
or U12350 (N_12350,N_12045,N_12197);
or U12351 (N_12351,N_12193,N_12114);
xnor U12352 (N_12352,N_12103,N_12108);
nand U12353 (N_12353,N_12152,N_12005);
xor U12354 (N_12354,N_12008,N_12146);
nand U12355 (N_12355,N_12072,N_12056);
nor U12356 (N_12356,N_12049,N_12037);
and U12357 (N_12357,N_12127,N_12000);
nand U12358 (N_12358,N_12193,N_12066);
xor U12359 (N_12359,N_12185,N_12076);
or U12360 (N_12360,N_12159,N_12154);
and U12361 (N_12361,N_12006,N_12051);
nand U12362 (N_12362,N_12016,N_12100);
nor U12363 (N_12363,N_12082,N_12113);
and U12364 (N_12364,N_12075,N_12116);
xor U12365 (N_12365,N_12068,N_12168);
xnor U12366 (N_12366,N_12137,N_12080);
or U12367 (N_12367,N_12032,N_12050);
nand U12368 (N_12368,N_12088,N_12110);
or U12369 (N_12369,N_12162,N_12088);
nand U12370 (N_12370,N_12173,N_12106);
nor U12371 (N_12371,N_12113,N_12146);
nand U12372 (N_12372,N_12055,N_12086);
nor U12373 (N_12373,N_12068,N_12145);
and U12374 (N_12374,N_12197,N_12038);
nand U12375 (N_12375,N_12011,N_12193);
nor U12376 (N_12376,N_12078,N_12099);
nor U12377 (N_12377,N_12152,N_12067);
or U12378 (N_12378,N_12020,N_12074);
nor U12379 (N_12379,N_12086,N_12174);
nor U12380 (N_12380,N_12018,N_12122);
or U12381 (N_12381,N_12133,N_12053);
nor U12382 (N_12382,N_12065,N_12046);
nor U12383 (N_12383,N_12032,N_12141);
nor U12384 (N_12384,N_12149,N_12119);
and U12385 (N_12385,N_12163,N_12044);
or U12386 (N_12386,N_12015,N_12024);
and U12387 (N_12387,N_12144,N_12162);
nand U12388 (N_12388,N_12079,N_12152);
nand U12389 (N_12389,N_12113,N_12003);
nand U12390 (N_12390,N_12178,N_12195);
nand U12391 (N_12391,N_12162,N_12149);
or U12392 (N_12392,N_12037,N_12180);
and U12393 (N_12393,N_12007,N_12000);
xnor U12394 (N_12394,N_12162,N_12117);
nand U12395 (N_12395,N_12177,N_12106);
nand U12396 (N_12396,N_12198,N_12121);
xor U12397 (N_12397,N_12071,N_12160);
or U12398 (N_12398,N_12069,N_12090);
nor U12399 (N_12399,N_12034,N_12138);
nor U12400 (N_12400,N_12366,N_12342);
or U12401 (N_12401,N_12292,N_12223);
and U12402 (N_12402,N_12267,N_12382);
nor U12403 (N_12403,N_12391,N_12312);
nand U12404 (N_12404,N_12399,N_12254);
and U12405 (N_12405,N_12266,N_12316);
nor U12406 (N_12406,N_12373,N_12248);
or U12407 (N_12407,N_12355,N_12271);
nand U12408 (N_12408,N_12349,N_12361);
xor U12409 (N_12409,N_12304,N_12206);
or U12410 (N_12410,N_12379,N_12335);
or U12411 (N_12411,N_12241,N_12222);
and U12412 (N_12412,N_12238,N_12330);
nor U12413 (N_12413,N_12287,N_12270);
xnor U12414 (N_12414,N_12237,N_12381);
nor U12415 (N_12415,N_12376,N_12224);
nand U12416 (N_12416,N_12336,N_12377);
or U12417 (N_12417,N_12329,N_12268);
and U12418 (N_12418,N_12392,N_12305);
xnor U12419 (N_12419,N_12228,N_12244);
nand U12420 (N_12420,N_12341,N_12339);
and U12421 (N_12421,N_12256,N_12394);
nor U12422 (N_12422,N_12294,N_12365);
and U12423 (N_12423,N_12326,N_12286);
or U12424 (N_12424,N_12340,N_12347);
nor U12425 (N_12425,N_12378,N_12221);
and U12426 (N_12426,N_12273,N_12219);
nand U12427 (N_12427,N_12321,N_12334);
nor U12428 (N_12428,N_12317,N_12320);
xor U12429 (N_12429,N_12277,N_12310);
nor U12430 (N_12430,N_12315,N_12331);
and U12431 (N_12431,N_12390,N_12300);
nor U12432 (N_12432,N_12220,N_12232);
nand U12433 (N_12433,N_12370,N_12204);
and U12434 (N_12434,N_12261,N_12225);
xor U12435 (N_12435,N_12291,N_12397);
or U12436 (N_12436,N_12386,N_12203);
nor U12437 (N_12437,N_12293,N_12367);
nor U12438 (N_12438,N_12202,N_12313);
and U12439 (N_12439,N_12395,N_12250);
and U12440 (N_12440,N_12284,N_12360);
nand U12441 (N_12441,N_12280,N_12281);
and U12442 (N_12442,N_12388,N_12332);
or U12443 (N_12443,N_12299,N_12308);
nand U12444 (N_12444,N_12307,N_12283);
or U12445 (N_12445,N_12375,N_12201);
or U12446 (N_12446,N_12230,N_12252);
or U12447 (N_12447,N_12306,N_12318);
or U12448 (N_12448,N_12240,N_12311);
or U12449 (N_12449,N_12362,N_12322);
xor U12450 (N_12450,N_12364,N_12231);
or U12451 (N_12451,N_12380,N_12385);
or U12452 (N_12452,N_12288,N_12324);
nand U12453 (N_12453,N_12338,N_12212);
nor U12454 (N_12454,N_12272,N_12215);
nor U12455 (N_12455,N_12258,N_12337);
xnor U12456 (N_12456,N_12285,N_12290);
nand U12457 (N_12457,N_12298,N_12278);
xnor U12458 (N_12458,N_12343,N_12319);
or U12459 (N_12459,N_12207,N_12372);
xor U12460 (N_12460,N_12297,N_12302);
nand U12461 (N_12461,N_12333,N_12249);
xor U12462 (N_12462,N_12259,N_12327);
nand U12463 (N_12463,N_12214,N_12369);
and U12464 (N_12464,N_12236,N_12354);
and U12465 (N_12465,N_12371,N_12282);
nor U12466 (N_12466,N_12289,N_12279);
nor U12467 (N_12467,N_12227,N_12374);
xnor U12468 (N_12468,N_12384,N_12247);
or U12469 (N_12469,N_12368,N_12350);
nand U12470 (N_12470,N_12396,N_12216);
nor U12471 (N_12471,N_12210,N_12323);
or U12472 (N_12472,N_12262,N_12260);
nand U12473 (N_12473,N_12218,N_12296);
or U12474 (N_12474,N_12314,N_12276);
or U12475 (N_12475,N_12351,N_12245);
xor U12476 (N_12476,N_12295,N_12363);
or U12477 (N_12477,N_12255,N_12348);
nand U12478 (N_12478,N_12274,N_12200);
or U12479 (N_12479,N_12251,N_12263);
or U12480 (N_12480,N_12253,N_12234);
and U12481 (N_12481,N_12243,N_12275);
nor U12482 (N_12482,N_12358,N_12325);
or U12483 (N_12483,N_12301,N_12357);
or U12484 (N_12484,N_12269,N_12309);
nand U12485 (N_12485,N_12213,N_12352);
nand U12486 (N_12486,N_12235,N_12398);
or U12487 (N_12487,N_12328,N_12229);
nor U12488 (N_12488,N_12383,N_12389);
or U12489 (N_12489,N_12211,N_12226);
and U12490 (N_12490,N_12303,N_12239);
nand U12491 (N_12491,N_12345,N_12393);
xnor U12492 (N_12492,N_12344,N_12205);
xor U12493 (N_12493,N_12233,N_12353);
or U12494 (N_12494,N_12387,N_12217);
or U12495 (N_12495,N_12346,N_12264);
nor U12496 (N_12496,N_12242,N_12265);
nor U12497 (N_12497,N_12257,N_12246);
nand U12498 (N_12498,N_12208,N_12359);
and U12499 (N_12499,N_12209,N_12356);
xnor U12500 (N_12500,N_12210,N_12303);
nor U12501 (N_12501,N_12248,N_12200);
or U12502 (N_12502,N_12244,N_12347);
xor U12503 (N_12503,N_12258,N_12210);
nand U12504 (N_12504,N_12364,N_12229);
or U12505 (N_12505,N_12372,N_12378);
and U12506 (N_12506,N_12374,N_12365);
and U12507 (N_12507,N_12314,N_12223);
nand U12508 (N_12508,N_12371,N_12291);
and U12509 (N_12509,N_12379,N_12220);
nand U12510 (N_12510,N_12354,N_12208);
or U12511 (N_12511,N_12221,N_12275);
and U12512 (N_12512,N_12359,N_12251);
xor U12513 (N_12513,N_12346,N_12252);
and U12514 (N_12514,N_12376,N_12290);
nor U12515 (N_12515,N_12361,N_12330);
and U12516 (N_12516,N_12377,N_12249);
nand U12517 (N_12517,N_12271,N_12231);
or U12518 (N_12518,N_12232,N_12236);
nor U12519 (N_12519,N_12270,N_12201);
xor U12520 (N_12520,N_12378,N_12211);
xnor U12521 (N_12521,N_12348,N_12217);
xnor U12522 (N_12522,N_12289,N_12354);
and U12523 (N_12523,N_12353,N_12287);
or U12524 (N_12524,N_12356,N_12344);
nand U12525 (N_12525,N_12337,N_12278);
nor U12526 (N_12526,N_12256,N_12340);
nor U12527 (N_12527,N_12231,N_12273);
and U12528 (N_12528,N_12219,N_12302);
or U12529 (N_12529,N_12209,N_12256);
nand U12530 (N_12530,N_12370,N_12223);
xnor U12531 (N_12531,N_12355,N_12292);
nand U12532 (N_12532,N_12273,N_12335);
or U12533 (N_12533,N_12330,N_12220);
or U12534 (N_12534,N_12226,N_12295);
nor U12535 (N_12535,N_12366,N_12214);
nand U12536 (N_12536,N_12211,N_12295);
and U12537 (N_12537,N_12375,N_12398);
and U12538 (N_12538,N_12297,N_12357);
or U12539 (N_12539,N_12323,N_12309);
nand U12540 (N_12540,N_12271,N_12272);
nor U12541 (N_12541,N_12377,N_12247);
or U12542 (N_12542,N_12257,N_12397);
nand U12543 (N_12543,N_12280,N_12256);
xor U12544 (N_12544,N_12385,N_12223);
xor U12545 (N_12545,N_12310,N_12398);
and U12546 (N_12546,N_12207,N_12234);
nor U12547 (N_12547,N_12327,N_12217);
xnor U12548 (N_12548,N_12338,N_12245);
xnor U12549 (N_12549,N_12306,N_12234);
nand U12550 (N_12550,N_12358,N_12396);
and U12551 (N_12551,N_12278,N_12242);
xnor U12552 (N_12552,N_12307,N_12337);
nand U12553 (N_12553,N_12397,N_12284);
xor U12554 (N_12554,N_12352,N_12306);
nor U12555 (N_12555,N_12257,N_12322);
and U12556 (N_12556,N_12231,N_12370);
nand U12557 (N_12557,N_12327,N_12365);
and U12558 (N_12558,N_12365,N_12212);
nand U12559 (N_12559,N_12201,N_12358);
nor U12560 (N_12560,N_12360,N_12287);
nand U12561 (N_12561,N_12298,N_12383);
xor U12562 (N_12562,N_12257,N_12310);
nand U12563 (N_12563,N_12363,N_12342);
xnor U12564 (N_12564,N_12364,N_12383);
nor U12565 (N_12565,N_12292,N_12392);
nor U12566 (N_12566,N_12355,N_12269);
and U12567 (N_12567,N_12232,N_12313);
nand U12568 (N_12568,N_12271,N_12216);
or U12569 (N_12569,N_12295,N_12385);
xnor U12570 (N_12570,N_12215,N_12294);
or U12571 (N_12571,N_12213,N_12220);
nand U12572 (N_12572,N_12294,N_12290);
and U12573 (N_12573,N_12315,N_12317);
or U12574 (N_12574,N_12221,N_12257);
nand U12575 (N_12575,N_12329,N_12222);
xor U12576 (N_12576,N_12379,N_12206);
nor U12577 (N_12577,N_12289,N_12361);
xnor U12578 (N_12578,N_12391,N_12200);
and U12579 (N_12579,N_12233,N_12254);
and U12580 (N_12580,N_12281,N_12303);
nand U12581 (N_12581,N_12372,N_12277);
nor U12582 (N_12582,N_12327,N_12347);
nand U12583 (N_12583,N_12238,N_12209);
xor U12584 (N_12584,N_12207,N_12369);
nand U12585 (N_12585,N_12232,N_12207);
or U12586 (N_12586,N_12237,N_12244);
nor U12587 (N_12587,N_12353,N_12350);
nor U12588 (N_12588,N_12359,N_12297);
nor U12589 (N_12589,N_12213,N_12337);
xnor U12590 (N_12590,N_12362,N_12301);
xnor U12591 (N_12591,N_12310,N_12207);
xnor U12592 (N_12592,N_12270,N_12330);
xor U12593 (N_12593,N_12262,N_12283);
nor U12594 (N_12594,N_12260,N_12228);
or U12595 (N_12595,N_12376,N_12234);
or U12596 (N_12596,N_12308,N_12358);
or U12597 (N_12597,N_12281,N_12298);
and U12598 (N_12598,N_12226,N_12220);
and U12599 (N_12599,N_12364,N_12355);
and U12600 (N_12600,N_12582,N_12436);
or U12601 (N_12601,N_12427,N_12482);
nor U12602 (N_12602,N_12517,N_12463);
xnor U12603 (N_12603,N_12501,N_12485);
nand U12604 (N_12604,N_12464,N_12483);
nor U12605 (N_12605,N_12520,N_12444);
nor U12606 (N_12606,N_12434,N_12418);
or U12607 (N_12607,N_12553,N_12521);
nand U12608 (N_12608,N_12571,N_12402);
or U12609 (N_12609,N_12411,N_12596);
xnor U12610 (N_12610,N_12577,N_12471);
nor U12611 (N_12611,N_12557,N_12440);
or U12612 (N_12612,N_12462,N_12410);
or U12613 (N_12613,N_12495,N_12515);
and U12614 (N_12614,N_12468,N_12435);
xor U12615 (N_12615,N_12539,N_12429);
nand U12616 (N_12616,N_12524,N_12446);
or U12617 (N_12617,N_12533,N_12522);
and U12618 (N_12618,N_12589,N_12570);
nor U12619 (N_12619,N_12567,N_12592);
nand U12620 (N_12620,N_12544,N_12449);
xnor U12621 (N_12621,N_12555,N_12494);
nor U12622 (N_12622,N_12467,N_12564);
xor U12623 (N_12623,N_12525,N_12474);
nand U12624 (N_12624,N_12426,N_12447);
xnor U12625 (N_12625,N_12560,N_12587);
xnor U12626 (N_12626,N_12597,N_12537);
xor U12627 (N_12627,N_12512,N_12432);
and U12628 (N_12628,N_12419,N_12425);
nor U12629 (N_12629,N_12579,N_12409);
or U12630 (N_12630,N_12565,N_12451);
xnor U12631 (N_12631,N_12442,N_12413);
and U12632 (N_12632,N_12486,N_12572);
or U12633 (N_12633,N_12558,N_12545);
xnor U12634 (N_12634,N_12518,N_12478);
xor U12635 (N_12635,N_12508,N_12591);
xor U12636 (N_12636,N_12532,N_12450);
nor U12637 (N_12637,N_12531,N_12480);
nor U12638 (N_12638,N_12417,N_12458);
nand U12639 (N_12639,N_12552,N_12403);
xnor U12640 (N_12640,N_12408,N_12400);
and U12641 (N_12641,N_12519,N_12405);
nor U12642 (N_12642,N_12493,N_12433);
xnor U12643 (N_12643,N_12487,N_12543);
or U12644 (N_12644,N_12504,N_12470);
nand U12645 (N_12645,N_12430,N_12509);
and U12646 (N_12646,N_12412,N_12424);
nand U12647 (N_12647,N_12420,N_12594);
xor U12648 (N_12648,N_12489,N_12505);
or U12649 (N_12649,N_12473,N_12448);
nand U12650 (N_12650,N_12526,N_12406);
xor U12651 (N_12651,N_12583,N_12438);
or U12652 (N_12652,N_12529,N_12514);
xor U12653 (N_12653,N_12569,N_12441);
and U12654 (N_12654,N_12456,N_12439);
nor U12655 (N_12655,N_12499,N_12461);
nor U12656 (N_12656,N_12479,N_12598);
xor U12657 (N_12657,N_12538,N_12503);
xnor U12658 (N_12658,N_12414,N_12530);
or U12659 (N_12659,N_12575,N_12465);
nor U12660 (N_12660,N_12584,N_12466);
and U12661 (N_12661,N_12588,N_12542);
and U12662 (N_12662,N_12590,N_12585);
xor U12663 (N_12663,N_12556,N_12459);
xor U12664 (N_12664,N_12527,N_12428);
xor U12665 (N_12665,N_12554,N_12416);
or U12666 (N_12666,N_12511,N_12422);
xor U12667 (N_12667,N_12490,N_12415);
or U12668 (N_12668,N_12492,N_12578);
nand U12669 (N_12669,N_12563,N_12566);
nor U12670 (N_12670,N_12475,N_12401);
xnor U12671 (N_12671,N_12506,N_12502);
xnor U12672 (N_12672,N_12573,N_12443);
nor U12673 (N_12673,N_12550,N_12407);
and U12674 (N_12674,N_12536,N_12528);
and U12675 (N_12675,N_12455,N_12500);
xnor U12676 (N_12676,N_12574,N_12593);
or U12677 (N_12677,N_12580,N_12549);
nor U12678 (N_12678,N_12491,N_12454);
nand U12679 (N_12679,N_12516,N_12576);
and U12680 (N_12680,N_12421,N_12513);
or U12681 (N_12681,N_12534,N_12546);
nand U12682 (N_12682,N_12477,N_12453);
or U12683 (N_12683,N_12586,N_12562);
or U12684 (N_12684,N_12540,N_12484);
nor U12685 (N_12685,N_12452,N_12510);
nand U12686 (N_12686,N_12595,N_12581);
or U12687 (N_12687,N_12568,N_12535);
nor U12688 (N_12688,N_12437,N_12523);
nand U12689 (N_12689,N_12469,N_12498);
and U12690 (N_12690,N_12423,N_12488);
nand U12691 (N_12691,N_12481,N_12445);
nand U12692 (N_12692,N_12551,N_12599);
xor U12693 (N_12693,N_12561,N_12404);
nor U12694 (N_12694,N_12472,N_12476);
or U12695 (N_12695,N_12547,N_12496);
nor U12696 (N_12696,N_12460,N_12457);
and U12697 (N_12697,N_12541,N_12548);
and U12698 (N_12698,N_12497,N_12559);
nand U12699 (N_12699,N_12431,N_12507);
nor U12700 (N_12700,N_12519,N_12415);
nand U12701 (N_12701,N_12580,N_12449);
and U12702 (N_12702,N_12522,N_12403);
nor U12703 (N_12703,N_12523,N_12469);
or U12704 (N_12704,N_12463,N_12470);
xor U12705 (N_12705,N_12438,N_12452);
and U12706 (N_12706,N_12514,N_12484);
or U12707 (N_12707,N_12561,N_12443);
nor U12708 (N_12708,N_12501,N_12532);
xnor U12709 (N_12709,N_12501,N_12551);
nor U12710 (N_12710,N_12527,N_12489);
xor U12711 (N_12711,N_12427,N_12534);
nor U12712 (N_12712,N_12430,N_12565);
and U12713 (N_12713,N_12573,N_12467);
or U12714 (N_12714,N_12525,N_12466);
and U12715 (N_12715,N_12446,N_12556);
xor U12716 (N_12716,N_12485,N_12554);
and U12717 (N_12717,N_12426,N_12575);
nand U12718 (N_12718,N_12446,N_12578);
xnor U12719 (N_12719,N_12502,N_12597);
nand U12720 (N_12720,N_12528,N_12491);
or U12721 (N_12721,N_12430,N_12410);
nor U12722 (N_12722,N_12489,N_12541);
nor U12723 (N_12723,N_12520,N_12429);
nand U12724 (N_12724,N_12430,N_12452);
nand U12725 (N_12725,N_12443,N_12589);
nand U12726 (N_12726,N_12510,N_12425);
and U12727 (N_12727,N_12460,N_12401);
nand U12728 (N_12728,N_12528,N_12496);
nor U12729 (N_12729,N_12510,N_12563);
and U12730 (N_12730,N_12506,N_12431);
nor U12731 (N_12731,N_12459,N_12418);
nor U12732 (N_12732,N_12557,N_12588);
xnor U12733 (N_12733,N_12516,N_12402);
nor U12734 (N_12734,N_12484,N_12594);
nand U12735 (N_12735,N_12593,N_12492);
nor U12736 (N_12736,N_12543,N_12438);
nor U12737 (N_12737,N_12537,N_12522);
xnor U12738 (N_12738,N_12430,N_12527);
and U12739 (N_12739,N_12497,N_12491);
nand U12740 (N_12740,N_12463,N_12450);
xnor U12741 (N_12741,N_12530,N_12454);
and U12742 (N_12742,N_12549,N_12585);
and U12743 (N_12743,N_12508,N_12490);
xnor U12744 (N_12744,N_12591,N_12483);
nand U12745 (N_12745,N_12448,N_12456);
nor U12746 (N_12746,N_12424,N_12427);
and U12747 (N_12747,N_12456,N_12583);
xnor U12748 (N_12748,N_12497,N_12442);
or U12749 (N_12749,N_12453,N_12447);
nor U12750 (N_12750,N_12561,N_12448);
xnor U12751 (N_12751,N_12414,N_12535);
and U12752 (N_12752,N_12533,N_12465);
and U12753 (N_12753,N_12465,N_12543);
nor U12754 (N_12754,N_12463,N_12545);
nor U12755 (N_12755,N_12596,N_12544);
and U12756 (N_12756,N_12540,N_12404);
xnor U12757 (N_12757,N_12473,N_12528);
nor U12758 (N_12758,N_12517,N_12505);
nor U12759 (N_12759,N_12519,N_12498);
nand U12760 (N_12760,N_12598,N_12444);
or U12761 (N_12761,N_12583,N_12488);
nand U12762 (N_12762,N_12540,N_12423);
nand U12763 (N_12763,N_12591,N_12465);
nor U12764 (N_12764,N_12451,N_12423);
nand U12765 (N_12765,N_12470,N_12421);
or U12766 (N_12766,N_12408,N_12436);
and U12767 (N_12767,N_12446,N_12523);
nor U12768 (N_12768,N_12418,N_12496);
and U12769 (N_12769,N_12483,N_12590);
nor U12770 (N_12770,N_12492,N_12584);
nor U12771 (N_12771,N_12492,N_12452);
and U12772 (N_12772,N_12435,N_12593);
nor U12773 (N_12773,N_12527,N_12405);
or U12774 (N_12774,N_12533,N_12413);
or U12775 (N_12775,N_12581,N_12576);
or U12776 (N_12776,N_12525,N_12448);
and U12777 (N_12777,N_12522,N_12553);
and U12778 (N_12778,N_12549,N_12470);
and U12779 (N_12779,N_12593,N_12556);
nand U12780 (N_12780,N_12551,N_12583);
nand U12781 (N_12781,N_12555,N_12452);
and U12782 (N_12782,N_12530,N_12571);
and U12783 (N_12783,N_12558,N_12570);
nor U12784 (N_12784,N_12495,N_12412);
and U12785 (N_12785,N_12447,N_12400);
xor U12786 (N_12786,N_12424,N_12557);
and U12787 (N_12787,N_12574,N_12421);
xor U12788 (N_12788,N_12411,N_12428);
or U12789 (N_12789,N_12590,N_12443);
xnor U12790 (N_12790,N_12401,N_12543);
nand U12791 (N_12791,N_12460,N_12412);
or U12792 (N_12792,N_12587,N_12540);
nor U12793 (N_12793,N_12448,N_12498);
or U12794 (N_12794,N_12455,N_12479);
xnor U12795 (N_12795,N_12461,N_12540);
and U12796 (N_12796,N_12480,N_12570);
or U12797 (N_12797,N_12424,N_12567);
nand U12798 (N_12798,N_12529,N_12486);
nand U12799 (N_12799,N_12518,N_12414);
nand U12800 (N_12800,N_12639,N_12720);
or U12801 (N_12801,N_12625,N_12652);
or U12802 (N_12802,N_12605,N_12678);
nor U12803 (N_12803,N_12701,N_12765);
nand U12804 (N_12804,N_12798,N_12776);
xnor U12805 (N_12805,N_12729,N_12671);
and U12806 (N_12806,N_12621,N_12766);
and U12807 (N_12807,N_12731,N_12742);
nor U12808 (N_12808,N_12643,N_12761);
nor U12809 (N_12809,N_12688,N_12704);
nor U12810 (N_12810,N_12660,N_12709);
nand U12811 (N_12811,N_12767,N_12614);
or U12812 (N_12812,N_12751,N_12746);
or U12813 (N_12813,N_12724,N_12663);
xnor U12814 (N_12814,N_12747,N_12775);
nand U12815 (N_12815,N_12758,N_12735);
nand U12816 (N_12816,N_12732,N_12697);
nand U12817 (N_12817,N_12753,N_12672);
nor U12818 (N_12818,N_12604,N_12656);
and U12819 (N_12819,N_12730,N_12721);
nand U12820 (N_12820,N_12629,N_12777);
nand U12821 (N_12821,N_12785,N_12637);
nand U12822 (N_12822,N_12771,N_12794);
or U12823 (N_12823,N_12658,N_12715);
nand U12824 (N_12824,N_12670,N_12769);
nor U12825 (N_12825,N_12630,N_12608);
nor U12826 (N_12826,N_12644,N_12788);
and U12827 (N_12827,N_12628,N_12622);
and U12828 (N_12828,N_12783,N_12682);
xnor U12829 (N_12829,N_12712,N_12738);
xnor U12830 (N_12830,N_12737,N_12781);
or U12831 (N_12831,N_12687,N_12651);
nand U12832 (N_12832,N_12726,N_12619);
nand U12833 (N_12833,N_12645,N_12733);
nand U12834 (N_12834,N_12779,N_12631);
nor U12835 (N_12835,N_12603,N_12602);
and U12836 (N_12836,N_12680,N_12627);
nor U12837 (N_12837,N_12741,N_12790);
xnor U12838 (N_12838,N_12750,N_12649);
xnor U12839 (N_12839,N_12772,N_12612);
and U12840 (N_12840,N_12725,N_12617);
nand U12841 (N_12841,N_12700,N_12673);
nor U12842 (N_12842,N_12686,N_12734);
nor U12843 (N_12843,N_12748,N_12676);
or U12844 (N_12844,N_12694,N_12754);
xnor U12845 (N_12845,N_12623,N_12667);
and U12846 (N_12846,N_12762,N_12799);
or U12847 (N_12847,N_12787,N_12710);
or U12848 (N_12848,N_12632,N_12662);
xor U12849 (N_12849,N_12634,N_12760);
nand U12850 (N_12850,N_12665,N_12780);
and U12851 (N_12851,N_12666,N_12706);
xnor U12852 (N_12852,N_12718,N_12739);
or U12853 (N_12853,N_12606,N_12740);
or U12854 (N_12854,N_12770,N_12763);
nand U12855 (N_12855,N_12797,N_12698);
or U12856 (N_12856,N_12723,N_12640);
xor U12857 (N_12857,N_12655,N_12600);
nand U12858 (N_12858,N_12692,N_12638);
nor U12859 (N_12859,N_12719,N_12684);
xnor U12860 (N_12860,N_12752,N_12650);
or U12861 (N_12861,N_12657,N_12626);
and U12862 (N_12862,N_12743,N_12793);
nor U12863 (N_12863,N_12653,N_12659);
nand U12864 (N_12864,N_12620,N_12635);
nand U12865 (N_12865,N_12683,N_12641);
xor U12866 (N_12866,N_12642,N_12764);
nor U12867 (N_12867,N_12610,N_12696);
or U12868 (N_12868,N_12782,N_12690);
nor U12869 (N_12869,N_12654,N_12669);
xor U12870 (N_12870,N_12749,N_12786);
nor U12871 (N_12871,N_12722,N_12611);
nand U12872 (N_12872,N_12711,N_12736);
nand U12873 (N_12873,N_12609,N_12744);
or U12874 (N_12874,N_12661,N_12689);
and U12875 (N_12875,N_12681,N_12796);
xor U12876 (N_12876,N_12699,N_12615);
or U12877 (N_12877,N_12668,N_12607);
xnor U12878 (N_12878,N_12708,N_12784);
or U12879 (N_12879,N_12714,N_12792);
xor U12880 (N_12880,N_12618,N_12677);
nand U12881 (N_12881,N_12624,N_12646);
and U12882 (N_12882,N_12778,N_12727);
and U12883 (N_12883,N_12773,N_12675);
or U12884 (N_12884,N_12757,N_12728);
or U12885 (N_12885,N_12685,N_12648);
and U12886 (N_12886,N_12647,N_12613);
or U12887 (N_12887,N_12601,N_12707);
xnor U12888 (N_12888,N_12745,N_12755);
nor U12889 (N_12889,N_12664,N_12702);
xor U12890 (N_12890,N_12768,N_12703);
nor U12891 (N_12891,N_12674,N_12795);
or U12892 (N_12892,N_12679,N_12713);
or U12893 (N_12893,N_12691,N_12774);
nor U12894 (N_12894,N_12717,N_12756);
nor U12895 (N_12895,N_12789,N_12705);
nor U12896 (N_12896,N_12616,N_12791);
and U12897 (N_12897,N_12633,N_12695);
nor U12898 (N_12898,N_12716,N_12759);
xor U12899 (N_12899,N_12693,N_12636);
or U12900 (N_12900,N_12644,N_12704);
xor U12901 (N_12901,N_12635,N_12601);
nand U12902 (N_12902,N_12751,N_12791);
and U12903 (N_12903,N_12701,N_12737);
and U12904 (N_12904,N_12665,N_12790);
xnor U12905 (N_12905,N_12782,N_12629);
and U12906 (N_12906,N_12793,N_12796);
xor U12907 (N_12907,N_12742,N_12793);
or U12908 (N_12908,N_12617,N_12774);
or U12909 (N_12909,N_12703,N_12720);
xnor U12910 (N_12910,N_12623,N_12603);
nand U12911 (N_12911,N_12747,N_12784);
nor U12912 (N_12912,N_12641,N_12764);
and U12913 (N_12913,N_12626,N_12770);
xnor U12914 (N_12914,N_12719,N_12628);
nand U12915 (N_12915,N_12786,N_12603);
xnor U12916 (N_12916,N_12717,N_12797);
or U12917 (N_12917,N_12616,N_12782);
xnor U12918 (N_12918,N_12768,N_12724);
or U12919 (N_12919,N_12649,N_12653);
xor U12920 (N_12920,N_12638,N_12765);
or U12921 (N_12921,N_12684,N_12679);
or U12922 (N_12922,N_12789,N_12674);
nand U12923 (N_12923,N_12686,N_12685);
xnor U12924 (N_12924,N_12767,N_12671);
xor U12925 (N_12925,N_12690,N_12643);
nand U12926 (N_12926,N_12788,N_12737);
xnor U12927 (N_12927,N_12651,N_12731);
xor U12928 (N_12928,N_12747,N_12726);
or U12929 (N_12929,N_12758,N_12675);
and U12930 (N_12930,N_12702,N_12643);
nor U12931 (N_12931,N_12783,N_12665);
nand U12932 (N_12932,N_12764,N_12780);
xor U12933 (N_12933,N_12606,N_12780);
nand U12934 (N_12934,N_12728,N_12624);
nand U12935 (N_12935,N_12666,N_12624);
nand U12936 (N_12936,N_12729,N_12612);
or U12937 (N_12937,N_12707,N_12607);
and U12938 (N_12938,N_12736,N_12661);
and U12939 (N_12939,N_12794,N_12737);
or U12940 (N_12940,N_12665,N_12606);
and U12941 (N_12941,N_12673,N_12774);
nand U12942 (N_12942,N_12660,N_12736);
and U12943 (N_12943,N_12685,N_12689);
or U12944 (N_12944,N_12662,N_12700);
or U12945 (N_12945,N_12732,N_12679);
nor U12946 (N_12946,N_12692,N_12715);
nand U12947 (N_12947,N_12627,N_12734);
and U12948 (N_12948,N_12735,N_12786);
xnor U12949 (N_12949,N_12754,N_12690);
or U12950 (N_12950,N_12611,N_12629);
and U12951 (N_12951,N_12672,N_12738);
nor U12952 (N_12952,N_12692,N_12649);
xor U12953 (N_12953,N_12707,N_12631);
nor U12954 (N_12954,N_12772,N_12636);
xor U12955 (N_12955,N_12661,N_12658);
xnor U12956 (N_12956,N_12707,N_12672);
or U12957 (N_12957,N_12775,N_12760);
xnor U12958 (N_12958,N_12634,N_12718);
or U12959 (N_12959,N_12694,N_12756);
xor U12960 (N_12960,N_12639,N_12764);
nand U12961 (N_12961,N_12609,N_12615);
or U12962 (N_12962,N_12648,N_12642);
xnor U12963 (N_12963,N_12645,N_12646);
and U12964 (N_12964,N_12737,N_12634);
or U12965 (N_12965,N_12713,N_12739);
or U12966 (N_12966,N_12735,N_12621);
or U12967 (N_12967,N_12609,N_12724);
xor U12968 (N_12968,N_12789,N_12686);
nand U12969 (N_12969,N_12607,N_12676);
or U12970 (N_12970,N_12774,N_12747);
or U12971 (N_12971,N_12674,N_12764);
or U12972 (N_12972,N_12743,N_12699);
or U12973 (N_12973,N_12658,N_12754);
nor U12974 (N_12974,N_12776,N_12648);
nor U12975 (N_12975,N_12764,N_12640);
nand U12976 (N_12976,N_12649,N_12617);
and U12977 (N_12977,N_12722,N_12652);
nor U12978 (N_12978,N_12658,N_12674);
and U12979 (N_12979,N_12689,N_12746);
and U12980 (N_12980,N_12750,N_12701);
or U12981 (N_12981,N_12607,N_12646);
and U12982 (N_12982,N_12739,N_12641);
nor U12983 (N_12983,N_12725,N_12688);
xnor U12984 (N_12984,N_12672,N_12780);
xor U12985 (N_12985,N_12720,N_12603);
or U12986 (N_12986,N_12764,N_12792);
and U12987 (N_12987,N_12680,N_12724);
and U12988 (N_12988,N_12705,N_12606);
nor U12989 (N_12989,N_12640,N_12620);
nor U12990 (N_12990,N_12622,N_12778);
nand U12991 (N_12991,N_12791,N_12729);
nand U12992 (N_12992,N_12705,N_12769);
and U12993 (N_12993,N_12680,N_12620);
and U12994 (N_12994,N_12612,N_12697);
nor U12995 (N_12995,N_12706,N_12792);
xnor U12996 (N_12996,N_12675,N_12653);
or U12997 (N_12997,N_12690,N_12619);
or U12998 (N_12998,N_12783,N_12628);
xnor U12999 (N_12999,N_12634,N_12772);
or U13000 (N_13000,N_12898,N_12969);
xor U13001 (N_13001,N_12879,N_12802);
nor U13002 (N_13002,N_12952,N_12829);
and U13003 (N_13003,N_12864,N_12940);
and U13004 (N_13004,N_12984,N_12887);
nand U13005 (N_13005,N_12995,N_12822);
or U13006 (N_13006,N_12891,N_12811);
and U13007 (N_13007,N_12884,N_12907);
nand U13008 (N_13008,N_12973,N_12923);
and U13009 (N_13009,N_12855,N_12926);
or U13010 (N_13010,N_12806,N_12915);
and U13011 (N_13011,N_12854,N_12970);
nor U13012 (N_13012,N_12976,N_12983);
nor U13013 (N_13013,N_12828,N_12847);
nor U13014 (N_13014,N_12933,N_12904);
nand U13015 (N_13015,N_12908,N_12857);
xor U13016 (N_13016,N_12853,N_12895);
and U13017 (N_13017,N_12818,N_12964);
nor U13018 (N_13018,N_12963,N_12883);
nand U13019 (N_13019,N_12954,N_12922);
or U13020 (N_13020,N_12878,N_12856);
or U13021 (N_13021,N_12832,N_12929);
nand U13022 (N_13022,N_12928,N_12815);
nand U13023 (N_13023,N_12881,N_12956);
xnor U13024 (N_13024,N_12919,N_12998);
nand U13025 (N_13025,N_12987,N_12972);
nor U13026 (N_13026,N_12824,N_12851);
xnor U13027 (N_13027,N_12981,N_12812);
nand U13028 (N_13028,N_12863,N_12823);
xor U13029 (N_13029,N_12842,N_12994);
nand U13030 (N_13030,N_12844,N_12902);
nand U13031 (N_13031,N_12942,N_12916);
nand U13032 (N_13032,N_12809,N_12861);
or U13033 (N_13033,N_12803,N_12989);
nor U13034 (N_13034,N_12900,N_12839);
nand U13035 (N_13035,N_12938,N_12996);
and U13036 (N_13036,N_12949,N_12936);
xor U13037 (N_13037,N_12885,N_12991);
and U13038 (N_13038,N_12944,N_12937);
and U13039 (N_13039,N_12850,N_12912);
nand U13040 (N_13040,N_12924,N_12993);
nand U13041 (N_13041,N_12875,N_12961);
or U13042 (N_13042,N_12968,N_12921);
xnor U13043 (N_13043,N_12999,N_12886);
nand U13044 (N_13044,N_12841,N_12880);
xor U13045 (N_13045,N_12992,N_12914);
nor U13046 (N_13046,N_12862,N_12931);
and U13047 (N_13047,N_12830,N_12892);
nor U13048 (N_13048,N_12906,N_12953);
or U13049 (N_13049,N_12897,N_12939);
nand U13050 (N_13050,N_12934,N_12889);
xnor U13051 (N_13051,N_12913,N_12810);
and U13052 (N_13052,N_12985,N_12846);
nand U13053 (N_13053,N_12941,N_12888);
or U13054 (N_13054,N_12868,N_12866);
nor U13055 (N_13055,N_12882,N_12852);
xnor U13056 (N_13056,N_12894,N_12927);
xor U13057 (N_13057,N_12849,N_12971);
nand U13058 (N_13058,N_12979,N_12917);
nand U13059 (N_13059,N_12826,N_12825);
nand U13060 (N_13060,N_12905,N_12958);
xor U13061 (N_13061,N_12858,N_12813);
xor U13062 (N_13062,N_12876,N_12836);
xnor U13063 (N_13063,N_12808,N_12955);
and U13064 (N_13064,N_12834,N_12903);
nand U13065 (N_13065,N_12877,N_12965);
xnor U13066 (N_13066,N_12920,N_12957);
and U13067 (N_13067,N_12977,N_12932);
and U13068 (N_13068,N_12959,N_12980);
nand U13069 (N_13069,N_12950,N_12974);
nand U13070 (N_13070,N_12918,N_12873);
and U13071 (N_13071,N_12820,N_12837);
or U13072 (N_13072,N_12827,N_12833);
nor U13073 (N_13073,N_12948,N_12848);
xnor U13074 (N_13074,N_12860,N_12859);
xor U13075 (N_13075,N_12960,N_12967);
nand U13076 (N_13076,N_12978,N_12990);
xor U13077 (N_13077,N_12890,N_12816);
nand U13078 (N_13078,N_12870,N_12869);
and U13079 (N_13079,N_12843,N_12817);
nand U13080 (N_13080,N_12867,N_12865);
nand U13081 (N_13081,N_12831,N_12801);
xnor U13082 (N_13082,N_12871,N_12982);
xnor U13083 (N_13083,N_12930,N_12947);
or U13084 (N_13084,N_12997,N_12935);
nand U13085 (N_13085,N_12840,N_12951);
xnor U13086 (N_13086,N_12845,N_12814);
and U13087 (N_13087,N_12986,N_12874);
nand U13088 (N_13088,N_12821,N_12962);
nand U13089 (N_13089,N_12911,N_12872);
nand U13090 (N_13090,N_12909,N_12925);
nand U13091 (N_13091,N_12819,N_12966);
nand U13092 (N_13092,N_12805,N_12800);
nand U13093 (N_13093,N_12835,N_12943);
nor U13094 (N_13094,N_12901,N_12807);
nand U13095 (N_13095,N_12893,N_12899);
nand U13096 (N_13096,N_12910,N_12804);
and U13097 (N_13097,N_12988,N_12975);
nand U13098 (N_13098,N_12838,N_12946);
or U13099 (N_13099,N_12945,N_12896);
nor U13100 (N_13100,N_12816,N_12883);
and U13101 (N_13101,N_12967,N_12927);
and U13102 (N_13102,N_12834,N_12883);
and U13103 (N_13103,N_12902,N_12994);
and U13104 (N_13104,N_12931,N_12990);
and U13105 (N_13105,N_12972,N_12876);
nand U13106 (N_13106,N_12944,N_12821);
nor U13107 (N_13107,N_12816,N_12805);
xor U13108 (N_13108,N_12879,N_12815);
or U13109 (N_13109,N_12881,N_12948);
xor U13110 (N_13110,N_12834,N_12839);
nor U13111 (N_13111,N_12903,N_12970);
nand U13112 (N_13112,N_12941,N_12943);
and U13113 (N_13113,N_12834,N_12964);
nor U13114 (N_13114,N_12979,N_12856);
nor U13115 (N_13115,N_12879,N_12948);
xnor U13116 (N_13116,N_12954,N_12944);
nor U13117 (N_13117,N_12873,N_12854);
nor U13118 (N_13118,N_12957,N_12945);
and U13119 (N_13119,N_12829,N_12885);
and U13120 (N_13120,N_12909,N_12849);
and U13121 (N_13121,N_12913,N_12978);
nor U13122 (N_13122,N_12928,N_12922);
xor U13123 (N_13123,N_12893,N_12800);
xnor U13124 (N_13124,N_12966,N_12876);
or U13125 (N_13125,N_12894,N_12877);
and U13126 (N_13126,N_12939,N_12914);
and U13127 (N_13127,N_12818,N_12969);
or U13128 (N_13128,N_12831,N_12904);
or U13129 (N_13129,N_12862,N_12892);
and U13130 (N_13130,N_12857,N_12881);
xnor U13131 (N_13131,N_12975,N_12803);
nor U13132 (N_13132,N_12975,N_12820);
and U13133 (N_13133,N_12981,N_12886);
nor U13134 (N_13134,N_12927,N_12859);
nand U13135 (N_13135,N_12852,N_12843);
and U13136 (N_13136,N_12862,N_12814);
xnor U13137 (N_13137,N_12957,N_12948);
xor U13138 (N_13138,N_12807,N_12849);
xor U13139 (N_13139,N_12841,N_12852);
nand U13140 (N_13140,N_12840,N_12835);
or U13141 (N_13141,N_12917,N_12962);
and U13142 (N_13142,N_12915,N_12832);
and U13143 (N_13143,N_12833,N_12938);
or U13144 (N_13144,N_12982,N_12821);
and U13145 (N_13145,N_12834,N_12915);
and U13146 (N_13146,N_12854,N_12839);
nor U13147 (N_13147,N_12990,N_12815);
nor U13148 (N_13148,N_12842,N_12858);
and U13149 (N_13149,N_12909,N_12994);
nor U13150 (N_13150,N_12993,N_12856);
nor U13151 (N_13151,N_12966,N_12806);
and U13152 (N_13152,N_12904,N_12802);
xor U13153 (N_13153,N_12808,N_12809);
and U13154 (N_13154,N_12981,N_12964);
or U13155 (N_13155,N_12823,N_12860);
nand U13156 (N_13156,N_12907,N_12857);
xor U13157 (N_13157,N_12855,N_12961);
xor U13158 (N_13158,N_12808,N_12964);
xnor U13159 (N_13159,N_12820,N_12807);
and U13160 (N_13160,N_12983,N_12887);
nor U13161 (N_13161,N_12831,N_12918);
nand U13162 (N_13162,N_12950,N_12921);
and U13163 (N_13163,N_12971,N_12972);
and U13164 (N_13164,N_12851,N_12955);
or U13165 (N_13165,N_12821,N_12890);
or U13166 (N_13166,N_12912,N_12969);
or U13167 (N_13167,N_12942,N_12850);
nor U13168 (N_13168,N_12916,N_12948);
xnor U13169 (N_13169,N_12898,N_12881);
xor U13170 (N_13170,N_12939,N_12930);
or U13171 (N_13171,N_12848,N_12860);
nor U13172 (N_13172,N_12897,N_12962);
nor U13173 (N_13173,N_12872,N_12978);
nor U13174 (N_13174,N_12940,N_12821);
nand U13175 (N_13175,N_12822,N_12801);
nor U13176 (N_13176,N_12925,N_12977);
xor U13177 (N_13177,N_12844,N_12960);
or U13178 (N_13178,N_12849,N_12891);
and U13179 (N_13179,N_12927,N_12999);
or U13180 (N_13180,N_12893,N_12951);
or U13181 (N_13181,N_12883,N_12821);
and U13182 (N_13182,N_12874,N_12881);
nand U13183 (N_13183,N_12936,N_12867);
and U13184 (N_13184,N_12916,N_12906);
nand U13185 (N_13185,N_12927,N_12919);
xor U13186 (N_13186,N_12984,N_12987);
or U13187 (N_13187,N_12832,N_12997);
or U13188 (N_13188,N_12929,N_12934);
nor U13189 (N_13189,N_12939,N_12907);
xor U13190 (N_13190,N_12842,N_12996);
nand U13191 (N_13191,N_12845,N_12886);
nor U13192 (N_13192,N_12957,N_12839);
nand U13193 (N_13193,N_12817,N_12829);
xor U13194 (N_13194,N_12808,N_12918);
nor U13195 (N_13195,N_12922,N_12873);
and U13196 (N_13196,N_12919,N_12986);
or U13197 (N_13197,N_12823,N_12944);
or U13198 (N_13198,N_12898,N_12865);
and U13199 (N_13199,N_12845,N_12958);
nor U13200 (N_13200,N_13120,N_13046);
xor U13201 (N_13201,N_13169,N_13186);
xnor U13202 (N_13202,N_13172,N_13071);
or U13203 (N_13203,N_13072,N_13077);
and U13204 (N_13204,N_13003,N_13113);
and U13205 (N_13205,N_13069,N_13190);
xnor U13206 (N_13206,N_13165,N_13138);
or U13207 (N_13207,N_13006,N_13085);
nand U13208 (N_13208,N_13183,N_13056);
xor U13209 (N_13209,N_13157,N_13009);
nand U13210 (N_13210,N_13121,N_13164);
nor U13211 (N_13211,N_13055,N_13038);
nand U13212 (N_13212,N_13149,N_13089);
and U13213 (N_13213,N_13115,N_13131);
nand U13214 (N_13214,N_13080,N_13163);
xnor U13215 (N_13215,N_13041,N_13062);
and U13216 (N_13216,N_13057,N_13052);
nand U13217 (N_13217,N_13134,N_13037);
or U13218 (N_13218,N_13002,N_13122);
xnor U13219 (N_13219,N_13017,N_13195);
or U13220 (N_13220,N_13197,N_13192);
nand U13221 (N_13221,N_13029,N_13187);
or U13222 (N_13222,N_13030,N_13175);
nand U13223 (N_13223,N_13160,N_13083);
xnor U13224 (N_13224,N_13094,N_13012);
or U13225 (N_13225,N_13061,N_13132);
or U13226 (N_13226,N_13063,N_13060);
xnor U13227 (N_13227,N_13161,N_13128);
or U13228 (N_13228,N_13199,N_13173);
xnor U13229 (N_13229,N_13107,N_13098);
xnor U13230 (N_13230,N_13171,N_13068);
or U13231 (N_13231,N_13150,N_13036);
nor U13232 (N_13232,N_13188,N_13184);
nor U13233 (N_13233,N_13126,N_13176);
nand U13234 (N_13234,N_13043,N_13004);
xor U13235 (N_13235,N_13090,N_13170);
or U13236 (N_13236,N_13116,N_13148);
nor U13237 (N_13237,N_13130,N_13021);
or U13238 (N_13238,N_13162,N_13189);
and U13239 (N_13239,N_13099,N_13155);
nand U13240 (N_13240,N_13000,N_13102);
or U13241 (N_13241,N_13185,N_13025);
nor U13242 (N_13242,N_13023,N_13124);
xor U13243 (N_13243,N_13081,N_13118);
xor U13244 (N_13244,N_13014,N_13059);
nand U13245 (N_13245,N_13180,N_13167);
and U13246 (N_13246,N_13127,N_13112);
and U13247 (N_13247,N_13086,N_13074);
and U13248 (N_13248,N_13073,N_13026);
or U13249 (N_13249,N_13159,N_13140);
xnor U13250 (N_13250,N_13129,N_13178);
xnor U13251 (N_13251,N_13151,N_13136);
and U13252 (N_13252,N_13109,N_13103);
and U13253 (N_13253,N_13028,N_13123);
xor U13254 (N_13254,N_13154,N_13117);
nor U13255 (N_13255,N_13067,N_13007);
nand U13256 (N_13256,N_13047,N_13179);
nor U13257 (N_13257,N_13108,N_13042);
or U13258 (N_13258,N_13093,N_13181);
xor U13259 (N_13259,N_13044,N_13051);
xnor U13260 (N_13260,N_13079,N_13153);
and U13261 (N_13261,N_13152,N_13168);
nor U13262 (N_13262,N_13145,N_13104);
nand U13263 (N_13263,N_13084,N_13182);
or U13264 (N_13264,N_13193,N_13065);
nand U13265 (N_13265,N_13091,N_13125);
nand U13266 (N_13266,N_13054,N_13142);
nand U13267 (N_13267,N_13008,N_13137);
xnor U13268 (N_13268,N_13040,N_13027);
nand U13269 (N_13269,N_13194,N_13015);
nor U13270 (N_13270,N_13147,N_13166);
nor U13271 (N_13271,N_13031,N_13177);
nor U13272 (N_13272,N_13045,N_13053);
nand U13273 (N_13273,N_13144,N_13033);
nand U13274 (N_13274,N_13114,N_13066);
nand U13275 (N_13275,N_13101,N_13135);
xor U13276 (N_13276,N_13034,N_13049);
nor U13277 (N_13277,N_13097,N_13005);
or U13278 (N_13278,N_13133,N_13024);
nand U13279 (N_13279,N_13013,N_13050);
xor U13280 (N_13280,N_13143,N_13087);
xnor U13281 (N_13281,N_13032,N_13010);
nand U13282 (N_13282,N_13019,N_13088);
nand U13283 (N_13283,N_13070,N_13001);
or U13284 (N_13284,N_13110,N_13156);
nand U13285 (N_13285,N_13105,N_13039);
and U13286 (N_13286,N_13064,N_13022);
xor U13287 (N_13287,N_13020,N_13139);
or U13288 (N_13288,N_13082,N_13095);
and U13289 (N_13289,N_13106,N_13100);
and U13290 (N_13290,N_13111,N_13035);
and U13291 (N_13291,N_13048,N_13141);
nor U13292 (N_13292,N_13196,N_13075);
and U13293 (N_13293,N_13016,N_13076);
and U13294 (N_13294,N_13119,N_13018);
nor U13295 (N_13295,N_13092,N_13078);
or U13296 (N_13296,N_13096,N_13191);
xor U13297 (N_13297,N_13058,N_13146);
and U13298 (N_13298,N_13011,N_13158);
nand U13299 (N_13299,N_13174,N_13198);
and U13300 (N_13300,N_13071,N_13195);
nor U13301 (N_13301,N_13193,N_13109);
or U13302 (N_13302,N_13190,N_13060);
and U13303 (N_13303,N_13150,N_13193);
nand U13304 (N_13304,N_13032,N_13185);
and U13305 (N_13305,N_13118,N_13067);
nand U13306 (N_13306,N_13113,N_13105);
or U13307 (N_13307,N_13103,N_13198);
xor U13308 (N_13308,N_13102,N_13090);
nor U13309 (N_13309,N_13025,N_13150);
xnor U13310 (N_13310,N_13020,N_13098);
or U13311 (N_13311,N_13038,N_13017);
or U13312 (N_13312,N_13135,N_13076);
nor U13313 (N_13313,N_13058,N_13159);
xnor U13314 (N_13314,N_13148,N_13156);
and U13315 (N_13315,N_13089,N_13103);
xor U13316 (N_13316,N_13011,N_13147);
or U13317 (N_13317,N_13113,N_13190);
nor U13318 (N_13318,N_13165,N_13074);
xnor U13319 (N_13319,N_13030,N_13158);
or U13320 (N_13320,N_13083,N_13064);
xor U13321 (N_13321,N_13096,N_13189);
and U13322 (N_13322,N_13174,N_13005);
nand U13323 (N_13323,N_13133,N_13109);
and U13324 (N_13324,N_13048,N_13194);
nand U13325 (N_13325,N_13005,N_13073);
and U13326 (N_13326,N_13010,N_13117);
xor U13327 (N_13327,N_13044,N_13126);
nor U13328 (N_13328,N_13173,N_13165);
nor U13329 (N_13329,N_13126,N_13101);
or U13330 (N_13330,N_13032,N_13004);
and U13331 (N_13331,N_13111,N_13055);
and U13332 (N_13332,N_13085,N_13182);
nor U13333 (N_13333,N_13147,N_13022);
xnor U13334 (N_13334,N_13129,N_13099);
nor U13335 (N_13335,N_13053,N_13064);
nand U13336 (N_13336,N_13124,N_13187);
xor U13337 (N_13337,N_13042,N_13189);
and U13338 (N_13338,N_13133,N_13119);
nand U13339 (N_13339,N_13025,N_13191);
nor U13340 (N_13340,N_13139,N_13001);
nand U13341 (N_13341,N_13183,N_13057);
nor U13342 (N_13342,N_13115,N_13121);
xnor U13343 (N_13343,N_13158,N_13129);
or U13344 (N_13344,N_13084,N_13156);
nor U13345 (N_13345,N_13122,N_13077);
nand U13346 (N_13346,N_13129,N_13000);
nor U13347 (N_13347,N_13129,N_13093);
or U13348 (N_13348,N_13166,N_13036);
nor U13349 (N_13349,N_13156,N_13072);
xnor U13350 (N_13350,N_13008,N_13195);
nor U13351 (N_13351,N_13110,N_13179);
and U13352 (N_13352,N_13014,N_13155);
xnor U13353 (N_13353,N_13066,N_13031);
xor U13354 (N_13354,N_13063,N_13012);
nor U13355 (N_13355,N_13096,N_13057);
nor U13356 (N_13356,N_13163,N_13044);
nand U13357 (N_13357,N_13111,N_13110);
or U13358 (N_13358,N_13026,N_13121);
nor U13359 (N_13359,N_13013,N_13135);
or U13360 (N_13360,N_13151,N_13190);
nand U13361 (N_13361,N_13130,N_13088);
or U13362 (N_13362,N_13176,N_13140);
nand U13363 (N_13363,N_13090,N_13180);
or U13364 (N_13364,N_13160,N_13190);
and U13365 (N_13365,N_13166,N_13063);
nand U13366 (N_13366,N_13038,N_13023);
nor U13367 (N_13367,N_13091,N_13004);
nand U13368 (N_13368,N_13073,N_13185);
nand U13369 (N_13369,N_13134,N_13076);
xnor U13370 (N_13370,N_13092,N_13104);
nor U13371 (N_13371,N_13123,N_13134);
or U13372 (N_13372,N_13003,N_13078);
xnor U13373 (N_13373,N_13182,N_13130);
or U13374 (N_13374,N_13182,N_13016);
or U13375 (N_13375,N_13178,N_13122);
xnor U13376 (N_13376,N_13028,N_13175);
and U13377 (N_13377,N_13143,N_13028);
nor U13378 (N_13378,N_13002,N_13178);
or U13379 (N_13379,N_13170,N_13190);
xnor U13380 (N_13380,N_13169,N_13108);
xnor U13381 (N_13381,N_13182,N_13026);
nand U13382 (N_13382,N_13143,N_13111);
nand U13383 (N_13383,N_13004,N_13185);
and U13384 (N_13384,N_13101,N_13068);
and U13385 (N_13385,N_13172,N_13079);
xor U13386 (N_13386,N_13054,N_13083);
nand U13387 (N_13387,N_13143,N_13188);
and U13388 (N_13388,N_13138,N_13116);
xnor U13389 (N_13389,N_13152,N_13060);
nor U13390 (N_13390,N_13093,N_13065);
and U13391 (N_13391,N_13156,N_13026);
nand U13392 (N_13392,N_13112,N_13130);
and U13393 (N_13393,N_13040,N_13179);
or U13394 (N_13394,N_13082,N_13041);
nand U13395 (N_13395,N_13082,N_13148);
nor U13396 (N_13396,N_13169,N_13004);
xnor U13397 (N_13397,N_13042,N_13175);
nand U13398 (N_13398,N_13019,N_13106);
and U13399 (N_13399,N_13072,N_13073);
xor U13400 (N_13400,N_13321,N_13396);
nand U13401 (N_13401,N_13209,N_13300);
and U13402 (N_13402,N_13324,N_13373);
nor U13403 (N_13403,N_13335,N_13305);
or U13404 (N_13404,N_13260,N_13370);
nor U13405 (N_13405,N_13262,N_13268);
and U13406 (N_13406,N_13333,N_13377);
xnor U13407 (N_13407,N_13252,N_13243);
nor U13408 (N_13408,N_13390,N_13232);
xnor U13409 (N_13409,N_13277,N_13384);
or U13410 (N_13410,N_13225,N_13206);
and U13411 (N_13411,N_13281,N_13343);
nand U13412 (N_13412,N_13267,N_13381);
and U13413 (N_13413,N_13273,N_13353);
nand U13414 (N_13414,N_13347,N_13357);
nor U13415 (N_13415,N_13298,N_13207);
xor U13416 (N_13416,N_13272,N_13361);
nand U13417 (N_13417,N_13286,N_13253);
xor U13418 (N_13418,N_13226,N_13284);
and U13419 (N_13419,N_13244,N_13372);
or U13420 (N_13420,N_13307,N_13246);
nand U13421 (N_13421,N_13364,N_13247);
or U13422 (N_13422,N_13388,N_13329);
xor U13423 (N_13423,N_13261,N_13397);
nand U13424 (N_13424,N_13367,N_13234);
and U13425 (N_13425,N_13395,N_13229);
or U13426 (N_13426,N_13204,N_13205);
and U13427 (N_13427,N_13250,N_13269);
xnor U13428 (N_13428,N_13316,N_13241);
xor U13429 (N_13429,N_13289,N_13236);
xnor U13430 (N_13430,N_13215,N_13276);
xor U13431 (N_13431,N_13210,N_13263);
nand U13432 (N_13432,N_13201,N_13233);
and U13433 (N_13433,N_13203,N_13290);
nor U13434 (N_13434,N_13295,N_13320);
nand U13435 (N_13435,N_13327,N_13266);
xnor U13436 (N_13436,N_13214,N_13336);
nor U13437 (N_13437,N_13212,N_13238);
nor U13438 (N_13438,N_13223,N_13382);
xnor U13439 (N_13439,N_13369,N_13334);
and U13440 (N_13440,N_13285,N_13365);
or U13441 (N_13441,N_13271,N_13355);
xor U13442 (N_13442,N_13371,N_13317);
and U13443 (N_13443,N_13342,N_13322);
or U13444 (N_13444,N_13213,N_13311);
xnor U13445 (N_13445,N_13323,N_13339);
or U13446 (N_13446,N_13265,N_13315);
nand U13447 (N_13447,N_13296,N_13366);
nor U13448 (N_13448,N_13235,N_13376);
or U13449 (N_13449,N_13221,N_13287);
and U13450 (N_13450,N_13310,N_13356);
nor U13451 (N_13451,N_13256,N_13344);
and U13452 (N_13452,N_13304,N_13280);
or U13453 (N_13453,N_13332,N_13274);
nor U13454 (N_13454,N_13362,N_13378);
nand U13455 (N_13455,N_13351,N_13216);
and U13456 (N_13456,N_13313,N_13319);
nor U13457 (N_13457,N_13259,N_13391);
nor U13458 (N_13458,N_13314,N_13374);
nor U13459 (N_13459,N_13202,N_13218);
and U13460 (N_13460,N_13275,N_13392);
nand U13461 (N_13461,N_13340,N_13325);
and U13462 (N_13462,N_13346,N_13270);
or U13463 (N_13463,N_13352,N_13379);
or U13464 (N_13464,N_13345,N_13258);
nor U13465 (N_13465,N_13200,N_13331);
and U13466 (N_13466,N_13227,N_13228);
nor U13467 (N_13467,N_13308,N_13237);
nand U13468 (N_13468,N_13254,N_13398);
xor U13469 (N_13469,N_13348,N_13341);
and U13470 (N_13470,N_13282,N_13350);
xnor U13471 (N_13471,N_13299,N_13338);
or U13472 (N_13472,N_13309,N_13288);
and U13473 (N_13473,N_13255,N_13393);
or U13474 (N_13474,N_13303,N_13245);
nor U13475 (N_13475,N_13231,N_13302);
and U13476 (N_13476,N_13359,N_13358);
nand U13477 (N_13477,N_13363,N_13240);
nor U13478 (N_13478,N_13279,N_13297);
xnor U13479 (N_13479,N_13360,N_13354);
nand U13480 (N_13480,N_13399,N_13368);
and U13481 (N_13481,N_13318,N_13375);
and U13482 (N_13482,N_13385,N_13389);
nor U13483 (N_13483,N_13330,N_13383);
or U13484 (N_13484,N_13301,N_13283);
xnor U13485 (N_13485,N_13211,N_13312);
xnor U13486 (N_13486,N_13292,N_13217);
and U13487 (N_13487,N_13220,N_13224);
and U13488 (N_13488,N_13294,N_13222);
and U13489 (N_13489,N_13394,N_13337);
or U13490 (N_13490,N_13326,N_13257);
nor U13491 (N_13491,N_13291,N_13230);
or U13492 (N_13492,N_13278,N_13208);
and U13493 (N_13493,N_13249,N_13293);
nor U13494 (N_13494,N_13380,N_13264);
xnor U13495 (N_13495,N_13328,N_13349);
xnor U13496 (N_13496,N_13386,N_13251);
and U13497 (N_13497,N_13248,N_13239);
and U13498 (N_13498,N_13306,N_13242);
nand U13499 (N_13499,N_13219,N_13387);
xnor U13500 (N_13500,N_13274,N_13286);
xor U13501 (N_13501,N_13280,N_13265);
or U13502 (N_13502,N_13227,N_13259);
or U13503 (N_13503,N_13286,N_13314);
or U13504 (N_13504,N_13382,N_13213);
nor U13505 (N_13505,N_13352,N_13218);
nor U13506 (N_13506,N_13356,N_13264);
xor U13507 (N_13507,N_13218,N_13386);
nor U13508 (N_13508,N_13372,N_13358);
and U13509 (N_13509,N_13203,N_13282);
or U13510 (N_13510,N_13249,N_13385);
and U13511 (N_13511,N_13379,N_13325);
nor U13512 (N_13512,N_13332,N_13348);
nand U13513 (N_13513,N_13208,N_13378);
or U13514 (N_13514,N_13303,N_13229);
nand U13515 (N_13515,N_13211,N_13377);
xnor U13516 (N_13516,N_13240,N_13297);
nor U13517 (N_13517,N_13301,N_13342);
xor U13518 (N_13518,N_13222,N_13345);
nor U13519 (N_13519,N_13300,N_13274);
or U13520 (N_13520,N_13217,N_13248);
xor U13521 (N_13521,N_13268,N_13202);
xor U13522 (N_13522,N_13346,N_13308);
nand U13523 (N_13523,N_13241,N_13294);
or U13524 (N_13524,N_13277,N_13320);
or U13525 (N_13525,N_13362,N_13395);
nand U13526 (N_13526,N_13236,N_13268);
xor U13527 (N_13527,N_13229,N_13347);
or U13528 (N_13528,N_13302,N_13330);
or U13529 (N_13529,N_13330,N_13399);
nor U13530 (N_13530,N_13297,N_13214);
xor U13531 (N_13531,N_13399,N_13348);
nor U13532 (N_13532,N_13357,N_13225);
xnor U13533 (N_13533,N_13304,N_13337);
and U13534 (N_13534,N_13258,N_13297);
nor U13535 (N_13535,N_13342,N_13211);
nor U13536 (N_13536,N_13342,N_13341);
nand U13537 (N_13537,N_13207,N_13222);
nand U13538 (N_13538,N_13262,N_13331);
or U13539 (N_13539,N_13385,N_13382);
or U13540 (N_13540,N_13380,N_13218);
nand U13541 (N_13541,N_13379,N_13324);
nand U13542 (N_13542,N_13356,N_13377);
xor U13543 (N_13543,N_13316,N_13280);
nor U13544 (N_13544,N_13347,N_13348);
and U13545 (N_13545,N_13340,N_13388);
nor U13546 (N_13546,N_13236,N_13214);
or U13547 (N_13547,N_13265,N_13384);
nor U13548 (N_13548,N_13252,N_13215);
xnor U13549 (N_13549,N_13273,N_13369);
and U13550 (N_13550,N_13233,N_13283);
xnor U13551 (N_13551,N_13319,N_13316);
or U13552 (N_13552,N_13378,N_13331);
or U13553 (N_13553,N_13228,N_13306);
nand U13554 (N_13554,N_13335,N_13326);
xor U13555 (N_13555,N_13345,N_13234);
and U13556 (N_13556,N_13307,N_13305);
xnor U13557 (N_13557,N_13233,N_13288);
or U13558 (N_13558,N_13203,N_13380);
xor U13559 (N_13559,N_13252,N_13267);
nor U13560 (N_13560,N_13228,N_13330);
and U13561 (N_13561,N_13314,N_13299);
nor U13562 (N_13562,N_13301,N_13360);
xnor U13563 (N_13563,N_13334,N_13266);
nor U13564 (N_13564,N_13207,N_13338);
nand U13565 (N_13565,N_13297,N_13397);
xnor U13566 (N_13566,N_13224,N_13304);
nand U13567 (N_13567,N_13317,N_13341);
nand U13568 (N_13568,N_13256,N_13272);
nand U13569 (N_13569,N_13337,N_13329);
nor U13570 (N_13570,N_13309,N_13316);
xor U13571 (N_13571,N_13301,N_13391);
nand U13572 (N_13572,N_13378,N_13263);
nor U13573 (N_13573,N_13336,N_13204);
nor U13574 (N_13574,N_13325,N_13329);
nand U13575 (N_13575,N_13383,N_13331);
xor U13576 (N_13576,N_13340,N_13334);
or U13577 (N_13577,N_13213,N_13224);
nor U13578 (N_13578,N_13363,N_13325);
xor U13579 (N_13579,N_13254,N_13368);
xnor U13580 (N_13580,N_13225,N_13271);
xnor U13581 (N_13581,N_13275,N_13327);
nor U13582 (N_13582,N_13218,N_13356);
nand U13583 (N_13583,N_13278,N_13313);
or U13584 (N_13584,N_13305,N_13243);
or U13585 (N_13585,N_13389,N_13287);
xor U13586 (N_13586,N_13245,N_13392);
nand U13587 (N_13587,N_13368,N_13397);
and U13588 (N_13588,N_13272,N_13279);
xor U13589 (N_13589,N_13319,N_13356);
xor U13590 (N_13590,N_13356,N_13316);
nor U13591 (N_13591,N_13354,N_13233);
and U13592 (N_13592,N_13297,N_13355);
or U13593 (N_13593,N_13339,N_13231);
or U13594 (N_13594,N_13390,N_13259);
and U13595 (N_13595,N_13325,N_13364);
and U13596 (N_13596,N_13223,N_13319);
and U13597 (N_13597,N_13315,N_13318);
or U13598 (N_13598,N_13210,N_13343);
and U13599 (N_13599,N_13355,N_13255);
xnor U13600 (N_13600,N_13538,N_13598);
or U13601 (N_13601,N_13427,N_13495);
and U13602 (N_13602,N_13555,N_13500);
or U13603 (N_13603,N_13482,N_13515);
nand U13604 (N_13604,N_13573,N_13497);
nor U13605 (N_13605,N_13431,N_13583);
nand U13606 (N_13606,N_13449,N_13422);
nor U13607 (N_13607,N_13432,N_13439);
nor U13608 (N_13608,N_13490,N_13564);
nor U13609 (N_13609,N_13503,N_13484);
or U13610 (N_13610,N_13553,N_13572);
and U13611 (N_13611,N_13400,N_13460);
or U13612 (N_13612,N_13480,N_13464);
xor U13613 (N_13613,N_13409,N_13536);
xnor U13614 (N_13614,N_13471,N_13517);
nor U13615 (N_13615,N_13529,N_13507);
xor U13616 (N_13616,N_13475,N_13445);
nor U13617 (N_13617,N_13588,N_13519);
nand U13618 (N_13618,N_13441,N_13408);
xor U13619 (N_13619,N_13410,N_13566);
or U13620 (N_13620,N_13448,N_13443);
and U13621 (N_13621,N_13590,N_13571);
nand U13622 (N_13622,N_13401,N_13418);
and U13623 (N_13623,N_13499,N_13524);
and U13624 (N_13624,N_13423,N_13550);
nor U13625 (N_13625,N_13470,N_13579);
xor U13626 (N_13626,N_13561,N_13461);
xnor U13627 (N_13627,N_13518,N_13474);
xor U13628 (N_13628,N_13522,N_13521);
and U13629 (N_13629,N_13544,N_13417);
xnor U13630 (N_13630,N_13584,N_13468);
nor U13631 (N_13631,N_13466,N_13446);
xor U13632 (N_13632,N_13543,N_13589);
xor U13633 (N_13633,N_13594,N_13537);
or U13634 (N_13634,N_13540,N_13523);
or U13635 (N_13635,N_13493,N_13514);
nor U13636 (N_13636,N_13508,N_13547);
or U13637 (N_13637,N_13558,N_13557);
nand U13638 (N_13638,N_13597,N_13428);
or U13639 (N_13639,N_13599,N_13509);
nor U13640 (N_13640,N_13429,N_13455);
or U13641 (N_13641,N_13488,N_13592);
nand U13642 (N_13642,N_13534,N_13501);
nand U13643 (N_13643,N_13463,N_13436);
and U13644 (N_13644,N_13494,N_13404);
nor U13645 (N_13645,N_13556,N_13551);
and U13646 (N_13646,N_13420,N_13469);
nor U13647 (N_13647,N_13434,N_13560);
nor U13648 (N_13648,N_13546,N_13442);
nand U13649 (N_13649,N_13402,N_13403);
nor U13650 (N_13650,N_13505,N_13533);
or U13651 (N_13651,N_13415,N_13511);
xor U13652 (N_13652,N_13481,N_13567);
or U13653 (N_13653,N_13438,N_13472);
nor U13654 (N_13654,N_13581,N_13453);
xor U13655 (N_13655,N_13525,N_13435);
nand U13656 (N_13656,N_13582,N_13465);
or U13657 (N_13657,N_13416,N_13548);
or U13658 (N_13658,N_13520,N_13526);
xor U13659 (N_13659,N_13549,N_13502);
or U13660 (N_13660,N_13559,N_13563);
nor U13661 (N_13661,N_13473,N_13596);
nor U13662 (N_13662,N_13447,N_13491);
and U13663 (N_13663,N_13437,N_13577);
and U13664 (N_13664,N_13498,N_13467);
and U13665 (N_13665,N_13462,N_13531);
nor U13666 (N_13666,N_13496,N_13444);
or U13667 (N_13667,N_13578,N_13510);
or U13668 (N_13668,N_13565,N_13430);
and U13669 (N_13669,N_13595,N_13458);
or U13670 (N_13670,N_13562,N_13552);
and U13671 (N_13671,N_13530,N_13414);
or U13672 (N_13672,N_13486,N_13532);
nand U13673 (N_13673,N_13593,N_13585);
and U13674 (N_13674,N_13452,N_13575);
and U13675 (N_13675,N_13411,N_13506);
nand U13676 (N_13676,N_13424,N_13513);
xnor U13677 (N_13677,N_13554,N_13454);
nand U13678 (N_13678,N_13419,N_13450);
and U13679 (N_13679,N_13489,N_13512);
nor U13680 (N_13680,N_13580,N_13492);
or U13681 (N_13681,N_13485,N_13483);
nor U13682 (N_13682,N_13413,N_13479);
xor U13683 (N_13683,N_13407,N_13433);
xor U13684 (N_13684,N_13476,N_13426);
and U13685 (N_13685,N_13478,N_13576);
and U13686 (N_13686,N_13574,N_13459);
nor U13687 (N_13687,N_13528,N_13440);
and U13688 (N_13688,N_13477,N_13504);
xnor U13689 (N_13689,N_13541,N_13457);
and U13690 (N_13690,N_13456,N_13405);
or U13691 (N_13691,N_13568,N_13570);
and U13692 (N_13692,N_13586,N_13587);
nand U13693 (N_13693,N_13421,N_13412);
nor U13694 (N_13694,N_13569,N_13527);
xor U13695 (N_13695,N_13425,N_13487);
xor U13696 (N_13696,N_13406,N_13591);
xnor U13697 (N_13697,N_13545,N_13516);
xor U13698 (N_13698,N_13542,N_13451);
nor U13699 (N_13699,N_13539,N_13535);
or U13700 (N_13700,N_13535,N_13520);
nand U13701 (N_13701,N_13408,N_13524);
nor U13702 (N_13702,N_13584,N_13464);
and U13703 (N_13703,N_13477,N_13454);
or U13704 (N_13704,N_13412,N_13492);
nor U13705 (N_13705,N_13440,N_13552);
and U13706 (N_13706,N_13465,N_13469);
nand U13707 (N_13707,N_13425,N_13548);
nor U13708 (N_13708,N_13522,N_13569);
xor U13709 (N_13709,N_13566,N_13577);
and U13710 (N_13710,N_13536,N_13468);
or U13711 (N_13711,N_13578,N_13473);
nand U13712 (N_13712,N_13508,N_13422);
nor U13713 (N_13713,N_13554,N_13448);
or U13714 (N_13714,N_13419,N_13476);
nor U13715 (N_13715,N_13557,N_13559);
nand U13716 (N_13716,N_13407,N_13515);
xor U13717 (N_13717,N_13582,N_13549);
nand U13718 (N_13718,N_13401,N_13486);
xnor U13719 (N_13719,N_13539,N_13556);
xnor U13720 (N_13720,N_13486,N_13420);
and U13721 (N_13721,N_13433,N_13553);
xor U13722 (N_13722,N_13585,N_13414);
nor U13723 (N_13723,N_13517,N_13503);
xor U13724 (N_13724,N_13577,N_13439);
or U13725 (N_13725,N_13474,N_13411);
nor U13726 (N_13726,N_13591,N_13409);
nor U13727 (N_13727,N_13442,N_13545);
and U13728 (N_13728,N_13578,N_13421);
nand U13729 (N_13729,N_13411,N_13492);
and U13730 (N_13730,N_13508,N_13568);
xor U13731 (N_13731,N_13497,N_13432);
nand U13732 (N_13732,N_13597,N_13429);
nor U13733 (N_13733,N_13407,N_13526);
xnor U13734 (N_13734,N_13572,N_13583);
xnor U13735 (N_13735,N_13520,N_13416);
or U13736 (N_13736,N_13462,N_13401);
nor U13737 (N_13737,N_13439,N_13423);
and U13738 (N_13738,N_13519,N_13584);
nand U13739 (N_13739,N_13462,N_13563);
and U13740 (N_13740,N_13573,N_13561);
nand U13741 (N_13741,N_13548,N_13581);
or U13742 (N_13742,N_13574,N_13439);
xnor U13743 (N_13743,N_13457,N_13504);
nand U13744 (N_13744,N_13417,N_13593);
or U13745 (N_13745,N_13513,N_13490);
nand U13746 (N_13746,N_13429,N_13442);
or U13747 (N_13747,N_13568,N_13582);
xor U13748 (N_13748,N_13505,N_13567);
xor U13749 (N_13749,N_13546,N_13523);
and U13750 (N_13750,N_13544,N_13491);
and U13751 (N_13751,N_13537,N_13576);
nor U13752 (N_13752,N_13456,N_13472);
xor U13753 (N_13753,N_13595,N_13400);
nand U13754 (N_13754,N_13588,N_13576);
xor U13755 (N_13755,N_13519,N_13518);
nor U13756 (N_13756,N_13478,N_13566);
nor U13757 (N_13757,N_13529,N_13427);
and U13758 (N_13758,N_13587,N_13502);
xor U13759 (N_13759,N_13424,N_13448);
nand U13760 (N_13760,N_13567,N_13540);
or U13761 (N_13761,N_13472,N_13548);
xnor U13762 (N_13762,N_13543,N_13459);
or U13763 (N_13763,N_13509,N_13481);
xnor U13764 (N_13764,N_13500,N_13586);
nor U13765 (N_13765,N_13541,N_13419);
or U13766 (N_13766,N_13462,N_13586);
nand U13767 (N_13767,N_13579,N_13474);
nor U13768 (N_13768,N_13507,N_13476);
nor U13769 (N_13769,N_13419,N_13401);
xor U13770 (N_13770,N_13599,N_13421);
and U13771 (N_13771,N_13550,N_13493);
nor U13772 (N_13772,N_13407,N_13484);
and U13773 (N_13773,N_13407,N_13501);
or U13774 (N_13774,N_13431,N_13444);
or U13775 (N_13775,N_13486,N_13572);
xor U13776 (N_13776,N_13492,N_13581);
and U13777 (N_13777,N_13519,N_13477);
or U13778 (N_13778,N_13581,N_13484);
or U13779 (N_13779,N_13430,N_13504);
or U13780 (N_13780,N_13490,N_13587);
nor U13781 (N_13781,N_13594,N_13418);
and U13782 (N_13782,N_13496,N_13495);
xnor U13783 (N_13783,N_13411,N_13531);
or U13784 (N_13784,N_13430,N_13451);
and U13785 (N_13785,N_13500,N_13558);
and U13786 (N_13786,N_13497,N_13587);
nor U13787 (N_13787,N_13456,N_13596);
xnor U13788 (N_13788,N_13521,N_13581);
or U13789 (N_13789,N_13511,N_13472);
xnor U13790 (N_13790,N_13567,N_13522);
nand U13791 (N_13791,N_13417,N_13401);
nor U13792 (N_13792,N_13582,N_13449);
nor U13793 (N_13793,N_13516,N_13510);
or U13794 (N_13794,N_13568,N_13524);
nand U13795 (N_13795,N_13501,N_13540);
and U13796 (N_13796,N_13594,N_13499);
nor U13797 (N_13797,N_13487,N_13571);
nand U13798 (N_13798,N_13501,N_13415);
xor U13799 (N_13799,N_13416,N_13589);
nor U13800 (N_13800,N_13687,N_13745);
or U13801 (N_13801,N_13763,N_13735);
nor U13802 (N_13802,N_13705,N_13636);
or U13803 (N_13803,N_13662,N_13722);
nor U13804 (N_13804,N_13759,N_13625);
and U13805 (N_13805,N_13708,N_13695);
nand U13806 (N_13806,N_13658,N_13781);
or U13807 (N_13807,N_13642,N_13679);
nor U13808 (N_13808,N_13716,N_13664);
nand U13809 (N_13809,N_13707,N_13758);
and U13810 (N_13810,N_13655,N_13721);
xor U13811 (N_13811,N_13739,N_13701);
xor U13812 (N_13812,N_13720,N_13671);
xnor U13813 (N_13813,N_13603,N_13746);
or U13814 (N_13814,N_13730,N_13798);
or U13815 (N_13815,N_13773,N_13681);
nor U13816 (N_13816,N_13756,N_13744);
xor U13817 (N_13817,N_13717,N_13651);
nor U13818 (N_13818,N_13747,N_13646);
and U13819 (N_13819,N_13614,N_13650);
nor U13820 (N_13820,N_13751,N_13620);
nand U13821 (N_13821,N_13616,N_13761);
and U13822 (N_13822,N_13785,N_13666);
and U13823 (N_13823,N_13784,N_13634);
or U13824 (N_13824,N_13704,N_13771);
nand U13825 (N_13825,N_13779,N_13690);
nor U13826 (N_13826,N_13768,N_13649);
xor U13827 (N_13827,N_13731,N_13790);
and U13828 (N_13828,N_13626,N_13633);
nor U13829 (N_13829,N_13733,N_13765);
xnor U13830 (N_13830,N_13712,N_13683);
xnor U13831 (N_13831,N_13602,N_13610);
nand U13832 (N_13832,N_13754,N_13792);
nand U13833 (N_13833,N_13613,N_13667);
or U13834 (N_13834,N_13685,N_13734);
xnor U13835 (N_13835,N_13797,N_13752);
or U13836 (N_13836,N_13622,N_13654);
nand U13837 (N_13837,N_13691,N_13689);
and U13838 (N_13838,N_13749,N_13668);
and U13839 (N_13839,N_13723,N_13778);
nor U13840 (N_13840,N_13680,N_13623);
nor U13841 (N_13841,N_13706,N_13688);
nand U13842 (N_13842,N_13686,N_13760);
nor U13843 (N_13843,N_13600,N_13672);
and U13844 (N_13844,N_13632,N_13630);
nand U13845 (N_13845,N_13656,N_13769);
nand U13846 (N_13846,N_13676,N_13791);
nor U13847 (N_13847,N_13719,N_13729);
nor U13848 (N_13848,N_13727,N_13660);
or U13849 (N_13849,N_13677,N_13608);
and U13850 (N_13850,N_13637,N_13713);
nor U13851 (N_13851,N_13742,N_13659);
nand U13852 (N_13852,N_13641,N_13678);
and U13853 (N_13853,N_13794,N_13640);
nor U13854 (N_13854,N_13710,N_13783);
nand U13855 (N_13855,N_13715,N_13697);
and U13856 (N_13856,N_13775,N_13652);
nor U13857 (N_13857,N_13748,N_13793);
nor U13858 (N_13858,N_13725,N_13601);
nand U13859 (N_13859,N_13682,N_13621);
nor U13860 (N_13860,N_13692,N_13669);
nand U13861 (N_13861,N_13675,N_13750);
nand U13862 (N_13862,N_13615,N_13703);
or U13863 (N_13863,N_13753,N_13770);
nor U13864 (N_13864,N_13766,N_13617);
or U13865 (N_13865,N_13714,N_13787);
or U13866 (N_13866,N_13767,N_13663);
or U13867 (N_13867,N_13743,N_13629);
xnor U13868 (N_13868,N_13631,N_13661);
nor U13869 (N_13869,N_13694,N_13673);
nand U13870 (N_13870,N_13718,N_13627);
or U13871 (N_13871,N_13604,N_13709);
xor U13872 (N_13872,N_13774,N_13657);
and U13873 (N_13873,N_13789,N_13638);
and U13874 (N_13874,N_13740,N_13648);
xnor U13875 (N_13875,N_13788,N_13738);
nor U13876 (N_13876,N_13647,N_13619);
and U13877 (N_13877,N_13635,N_13700);
xor U13878 (N_13878,N_13782,N_13605);
nand U13879 (N_13879,N_13737,N_13757);
nand U13880 (N_13880,N_13776,N_13607);
and U13881 (N_13881,N_13618,N_13777);
and U13882 (N_13882,N_13772,N_13699);
nand U13883 (N_13883,N_13702,N_13670);
nand U13884 (N_13884,N_13780,N_13795);
xnor U13885 (N_13885,N_13732,N_13724);
nand U13886 (N_13886,N_13755,N_13644);
nor U13887 (N_13887,N_13609,N_13628);
nor U13888 (N_13888,N_13786,N_13696);
or U13889 (N_13889,N_13674,N_13796);
xnor U13890 (N_13890,N_13726,N_13611);
and U13891 (N_13891,N_13762,N_13645);
or U13892 (N_13892,N_13643,N_13606);
nand U13893 (N_13893,N_13639,N_13693);
xor U13894 (N_13894,N_13684,N_13764);
xor U13895 (N_13895,N_13728,N_13624);
nand U13896 (N_13896,N_13612,N_13741);
xor U13897 (N_13897,N_13799,N_13665);
xnor U13898 (N_13898,N_13653,N_13736);
and U13899 (N_13899,N_13698,N_13711);
and U13900 (N_13900,N_13719,N_13721);
nor U13901 (N_13901,N_13799,N_13716);
xor U13902 (N_13902,N_13742,N_13698);
nand U13903 (N_13903,N_13774,N_13737);
nand U13904 (N_13904,N_13681,N_13758);
and U13905 (N_13905,N_13602,N_13651);
nor U13906 (N_13906,N_13699,N_13608);
or U13907 (N_13907,N_13659,N_13743);
or U13908 (N_13908,N_13766,N_13676);
nor U13909 (N_13909,N_13761,N_13783);
or U13910 (N_13910,N_13781,N_13729);
or U13911 (N_13911,N_13695,N_13618);
or U13912 (N_13912,N_13697,N_13667);
and U13913 (N_13913,N_13776,N_13773);
nor U13914 (N_13914,N_13660,N_13605);
xnor U13915 (N_13915,N_13603,N_13794);
and U13916 (N_13916,N_13753,N_13740);
and U13917 (N_13917,N_13677,N_13643);
xor U13918 (N_13918,N_13626,N_13795);
and U13919 (N_13919,N_13661,N_13780);
nand U13920 (N_13920,N_13710,N_13612);
xor U13921 (N_13921,N_13724,N_13773);
nand U13922 (N_13922,N_13777,N_13797);
and U13923 (N_13923,N_13671,N_13616);
xor U13924 (N_13924,N_13682,N_13740);
or U13925 (N_13925,N_13669,N_13670);
or U13926 (N_13926,N_13606,N_13641);
nor U13927 (N_13927,N_13726,N_13658);
or U13928 (N_13928,N_13661,N_13641);
xnor U13929 (N_13929,N_13792,N_13657);
or U13930 (N_13930,N_13660,N_13674);
or U13931 (N_13931,N_13636,N_13669);
nand U13932 (N_13932,N_13723,N_13619);
nand U13933 (N_13933,N_13622,N_13749);
nor U13934 (N_13934,N_13792,N_13749);
xnor U13935 (N_13935,N_13687,N_13770);
or U13936 (N_13936,N_13610,N_13744);
xor U13937 (N_13937,N_13698,N_13780);
xnor U13938 (N_13938,N_13769,N_13798);
nor U13939 (N_13939,N_13631,N_13715);
nor U13940 (N_13940,N_13643,N_13621);
and U13941 (N_13941,N_13776,N_13734);
or U13942 (N_13942,N_13673,N_13705);
nand U13943 (N_13943,N_13678,N_13673);
nor U13944 (N_13944,N_13750,N_13718);
and U13945 (N_13945,N_13790,N_13669);
nor U13946 (N_13946,N_13794,N_13605);
nor U13947 (N_13947,N_13663,N_13773);
xnor U13948 (N_13948,N_13607,N_13687);
nand U13949 (N_13949,N_13696,N_13735);
nor U13950 (N_13950,N_13604,N_13793);
or U13951 (N_13951,N_13643,N_13627);
and U13952 (N_13952,N_13621,N_13657);
or U13953 (N_13953,N_13637,N_13686);
or U13954 (N_13954,N_13602,N_13789);
nand U13955 (N_13955,N_13625,N_13638);
nor U13956 (N_13956,N_13622,N_13684);
and U13957 (N_13957,N_13687,N_13612);
nor U13958 (N_13958,N_13649,N_13793);
nor U13959 (N_13959,N_13754,N_13666);
xor U13960 (N_13960,N_13749,N_13604);
nand U13961 (N_13961,N_13633,N_13682);
nand U13962 (N_13962,N_13676,N_13655);
nor U13963 (N_13963,N_13755,N_13785);
xor U13964 (N_13964,N_13679,N_13774);
or U13965 (N_13965,N_13617,N_13670);
and U13966 (N_13966,N_13712,N_13798);
or U13967 (N_13967,N_13793,N_13719);
nor U13968 (N_13968,N_13791,N_13707);
xnor U13969 (N_13969,N_13655,N_13695);
nand U13970 (N_13970,N_13764,N_13695);
nor U13971 (N_13971,N_13766,N_13687);
or U13972 (N_13972,N_13767,N_13706);
nand U13973 (N_13973,N_13639,N_13623);
or U13974 (N_13974,N_13679,N_13751);
xnor U13975 (N_13975,N_13730,N_13789);
nand U13976 (N_13976,N_13662,N_13693);
nor U13977 (N_13977,N_13671,N_13695);
nand U13978 (N_13978,N_13639,N_13713);
and U13979 (N_13979,N_13642,N_13772);
or U13980 (N_13980,N_13748,N_13744);
nand U13981 (N_13981,N_13759,N_13610);
xnor U13982 (N_13982,N_13632,N_13646);
nand U13983 (N_13983,N_13664,N_13623);
or U13984 (N_13984,N_13740,N_13609);
xor U13985 (N_13985,N_13791,N_13793);
and U13986 (N_13986,N_13635,N_13742);
and U13987 (N_13987,N_13723,N_13762);
or U13988 (N_13988,N_13743,N_13763);
xnor U13989 (N_13989,N_13632,N_13662);
or U13990 (N_13990,N_13763,N_13696);
nor U13991 (N_13991,N_13632,N_13675);
nand U13992 (N_13992,N_13699,N_13751);
nand U13993 (N_13993,N_13667,N_13625);
or U13994 (N_13994,N_13697,N_13764);
xnor U13995 (N_13995,N_13664,N_13634);
and U13996 (N_13996,N_13753,N_13687);
nand U13997 (N_13997,N_13722,N_13641);
xnor U13998 (N_13998,N_13701,N_13713);
nand U13999 (N_13999,N_13722,N_13761);
nor U14000 (N_14000,N_13888,N_13851);
and U14001 (N_14001,N_13951,N_13923);
nand U14002 (N_14002,N_13801,N_13901);
nand U14003 (N_14003,N_13973,N_13886);
xnor U14004 (N_14004,N_13814,N_13993);
xnor U14005 (N_14005,N_13980,N_13815);
nor U14006 (N_14006,N_13842,N_13996);
and U14007 (N_14007,N_13865,N_13964);
and U14008 (N_14008,N_13962,N_13843);
xor U14009 (N_14009,N_13957,N_13953);
and U14010 (N_14010,N_13872,N_13885);
xor U14011 (N_14011,N_13868,N_13828);
nor U14012 (N_14012,N_13897,N_13981);
nand U14013 (N_14013,N_13822,N_13864);
nand U14014 (N_14014,N_13956,N_13915);
and U14015 (N_14015,N_13986,N_13803);
xor U14016 (N_14016,N_13987,N_13912);
xnor U14017 (N_14017,N_13858,N_13806);
xnor U14018 (N_14018,N_13892,N_13982);
xnor U14019 (N_14019,N_13989,N_13840);
xnor U14020 (N_14020,N_13808,N_13831);
nand U14021 (N_14021,N_13893,N_13811);
nand U14022 (N_14022,N_13859,N_13926);
nand U14023 (N_14023,N_13807,N_13903);
nand U14024 (N_14024,N_13934,N_13999);
or U14025 (N_14025,N_13940,N_13849);
nor U14026 (N_14026,N_13944,N_13933);
nand U14027 (N_14027,N_13967,N_13873);
nor U14028 (N_14028,N_13970,N_13927);
and U14029 (N_14029,N_13833,N_13832);
and U14030 (N_14030,N_13985,N_13949);
and U14031 (N_14031,N_13917,N_13820);
xnor U14032 (N_14032,N_13984,N_13916);
or U14033 (N_14033,N_13850,N_13979);
or U14034 (N_14034,N_13845,N_13847);
nand U14035 (N_14035,N_13998,N_13939);
and U14036 (N_14036,N_13818,N_13860);
and U14037 (N_14037,N_13961,N_13930);
nor U14038 (N_14038,N_13976,N_13854);
xnor U14039 (N_14039,N_13804,N_13972);
nand U14040 (N_14040,N_13805,N_13846);
or U14041 (N_14041,N_13899,N_13813);
nor U14042 (N_14042,N_13900,N_13884);
or U14043 (N_14043,N_13902,N_13974);
xor U14044 (N_14044,N_13827,N_13932);
or U14045 (N_14045,N_13830,N_13988);
and U14046 (N_14046,N_13906,N_13894);
nor U14047 (N_14047,N_13861,N_13878);
or U14048 (N_14048,N_13817,N_13966);
and U14049 (N_14049,N_13880,N_13834);
and U14050 (N_14050,N_13909,N_13887);
and U14051 (N_14051,N_13852,N_13863);
and U14052 (N_14052,N_13866,N_13836);
and U14053 (N_14053,N_13890,N_13874);
xor U14054 (N_14054,N_13876,N_13826);
and U14055 (N_14055,N_13907,N_13954);
xor U14056 (N_14056,N_13844,N_13918);
nand U14057 (N_14057,N_13875,N_13883);
nor U14058 (N_14058,N_13920,N_13928);
xor U14059 (N_14059,N_13855,N_13881);
nor U14060 (N_14060,N_13889,N_13848);
and U14061 (N_14061,N_13908,N_13945);
and U14062 (N_14062,N_13871,N_13943);
or U14063 (N_14063,N_13877,N_13936);
nor U14064 (N_14064,N_13952,N_13921);
and U14065 (N_14065,N_13810,N_13958);
xor U14066 (N_14066,N_13968,N_13870);
nand U14067 (N_14067,N_13812,N_13965);
and U14068 (N_14068,N_13963,N_13800);
or U14069 (N_14069,N_13839,N_13929);
nand U14070 (N_14070,N_13816,N_13802);
xor U14071 (N_14071,N_13862,N_13857);
xnor U14072 (N_14072,N_13955,N_13819);
or U14073 (N_14073,N_13948,N_13835);
or U14074 (N_14074,N_13910,N_13960);
and U14075 (N_14075,N_13853,N_13925);
nand U14076 (N_14076,N_13838,N_13896);
or U14077 (N_14077,N_13914,N_13895);
nand U14078 (N_14078,N_13942,N_13924);
or U14079 (N_14079,N_13856,N_13931);
or U14080 (N_14080,N_13823,N_13959);
and U14081 (N_14081,N_13992,N_13971);
and U14082 (N_14082,N_13983,N_13829);
nor U14083 (N_14083,N_13990,N_13994);
and U14084 (N_14084,N_13911,N_13950);
nor U14085 (N_14085,N_13904,N_13837);
and U14086 (N_14086,N_13891,N_13997);
nor U14087 (N_14087,N_13869,N_13898);
nand U14088 (N_14088,N_13947,N_13977);
xor U14089 (N_14089,N_13991,N_13935);
xnor U14090 (N_14090,N_13937,N_13975);
nand U14091 (N_14091,N_13913,N_13941);
and U14092 (N_14092,N_13821,N_13922);
or U14093 (N_14093,N_13946,N_13978);
or U14094 (N_14094,N_13825,N_13938);
xor U14095 (N_14095,N_13882,N_13867);
nor U14096 (N_14096,N_13905,N_13841);
or U14097 (N_14097,N_13995,N_13919);
nor U14098 (N_14098,N_13809,N_13824);
nor U14099 (N_14099,N_13879,N_13969);
nor U14100 (N_14100,N_13820,N_13969);
and U14101 (N_14101,N_13931,N_13888);
xnor U14102 (N_14102,N_13855,N_13893);
xor U14103 (N_14103,N_13970,N_13986);
or U14104 (N_14104,N_13863,N_13923);
nand U14105 (N_14105,N_13878,N_13908);
and U14106 (N_14106,N_13834,N_13814);
nand U14107 (N_14107,N_13938,N_13951);
or U14108 (N_14108,N_13898,N_13954);
nor U14109 (N_14109,N_13824,N_13959);
and U14110 (N_14110,N_13925,N_13955);
xor U14111 (N_14111,N_13802,N_13995);
xnor U14112 (N_14112,N_13815,N_13830);
and U14113 (N_14113,N_13851,N_13815);
or U14114 (N_14114,N_13812,N_13886);
xnor U14115 (N_14115,N_13858,N_13992);
nor U14116 (N_14116,N_13806,N_13867);
nand U14117 (N_14117,N_13997,N_13916);
or U14118 (N_14118,N_13914,N_13906);
nor U14119 (N_14119,N_13990,N_13834);
nor U14120 (N_14120,N_13830,N_13819);
xnor U14121 (N_14121,N_13886,N_13877);
nand U14122 (N_14122,N_13887,N_13987);
and U14123 (N_14123,N_13933,N_13826);
or U14124 (N_14124,N_13858,N_13881);
nor U14125 (N_14125,N_13939,N_13827);
or U14126 (N_14126,N_13847,N_13828);
xnor U14127 (N_14127,N_13872,N_13887);
nand U14128 (N_14128,N_13849,N_13824);
nand U14129 (N_14129,N_13969,N_13893);
or U14130 (N_14130,N_13893,N_13966);
nand U14131 (N_14131,N_13998,N_13833);
nor U14132 (N_14132,N_13928,N_13938);
nor U14133 (N_14133,N_13900,N_13808);
xor U14134 (N_14134,N_13964,N_13884);
xnor U14135 (N_14135,N_13922,N_13995);
and U14136 (N_14136,N_13975,N_13821);
nor U14137 (N_14137,N_13897,N_13939);
nor U14138 (N_14138,N_13908,N_13986);
or U14139 (N_14139,N_13855,N_13906);
and U14140 (N_14140,N_13832,N_13810);
nor U14141 (N_14141,N_13887,N_13833);
nand U14142 (N_14142,N_13848,N_13844);
xor U14143 (N_14143,N_13918,N_13851);
xor U14144 (N_14144,N_13915,N_13846);
or U14145 (N_14145,N_13961,N_13907);
or U14146 (N_14146,N_13842,N_13991);
nand U14147 (N_14147,N_13868,N_13921);
and U14148 (N_14148,N_13919,N_13947);
and U14149 (N_14149,N_13964,N_13847);
xnor U14150 (N_14150,N_13931,N_13958);
or U14151 (N_14151,N_13865,N_13912);
nor U14152 (N_14152,N_13963,N_13947);
nand U14153 (N_14153,N_13876,N_13885);
or U14154 (N_14154,N_13979,N_13970);
nand U14155 (N_14155,N_13834,N_13822);
xnor U14156 (N_14156,N_13823,N_13844);
nor U14157 (N_14157,N_13962,N_13936);
nor U14158 (N_14158,N_13948,N_13904);
nor U14159 (N_14159,N_13852,N_13850);
nor U14160 (N_14160,N_13886,N_13874);
and U14161 (N_14161,N_13963,N_13917);
nand U14162 (N_14162,N_13918,N_13826);
nor U14163 (N_14163,N_13842,N_13860);
nand U14164 (N_14164,N_13800,N_13871);
nand U14165 (N_14165,N_13992,N_13901);
nand U14166 (N_14166,N_13856,N_13988);
or U14167 (N_14167,N_13923,N_13885);
nand U14168 (N_14168,N_13898,N_13971);
or U14169 (N_14169,N_13952,N_13856);
xnor U14170 (N_14170,N_13879,N_13884);
nand U14171 (N_14171,N_13825,N_13905);
nand U14172 (N_14172,N_13912,N_13829);
and U14173 (N_14173,N_13857,N_13877);
or U14174 (N_14174,N_13991,N_13807);
xnor U14175 (N_14175,N_13886,N_13808);
nor U14176 (N_14176,N_13991,N_13818);
nand U14177 (N_14177,N_13962,N_13939);
or U14178 (N_14178,N_13935,N_13830);
or U14179 (N_14179,N_13986,N_13848);
nor U14180 (N_14180,N_13979,N_13951);
and U14181 (N_14181,N_13969,N_13831);
and U14182 (N_14182,N_13857,N_13950);
nand U14183 (N_14183,N_13837,N_13809);
and U14184 (N_14184,N_13892,N_13967);
nor U14185 (N_14185,N_13956,N_13947);
xor U14186 (N_14186,N_13929,N_13876);
and U14187 (N_14187,N_13921,N_13859);
or U14188 (N_14188,N_13992,N_13930);
nand U14189 (N_14189,N_13983,N_13984);
nand U14190 (N_14190,N_13859,N_13929);
or U14191 (N_14191,N_13809,N_13828);
and U14192 (N_14192,N_13834,N_13843);
nor U14193 (N_14193,N_13994,N_13835);
or U14194 (N_14194,N_13897,N_13930);
or U14195 (N_14195,N_13923,N_13813);
and U14196 (N_14196,N_13889,N_13976);
nand U14197 (N_14197,N_13816,N_13895);
nor U14198 (N_14198,N_13949,N_13827);
nand U14199 (N_14199,N_13838,N_13982);
nand U14200 (N_14200,N_14116,N_14046);
nor U14201 (N_14201,N_14195,N_14171);
nand U14202 (N_14202,N_14052,N_14061);
xnor U14203 (N_14203,N_14187,N_14117);
nor U14204 (N_14204,N_14142,N_14073);
nand U14205 (N_14205,N_14088,N_14081);
nor U14206 (N_14206,N_14004,N_14023);
nand U14207 (N_14207,N_14125,N_14135);
nand U14208 (N_14208,N_14167,N_14177);
xnor U14209 (N_14209,N_14018,N_14127);
and U14210 (N_14210,N_14038,N_14031);
and U14211 (N_14211,N_14027,N_14013);
and U14212 (N_14212,N_14074,N_14162);
or U14213 (N_14213,N_14030,N_14131);
and U14214 (N_14214,N_14165,N_14179);
xor U14215 (N_14215,N_14028,N_14076);
nor U14216 (N_14216,N_14136,N_14093);
xor U14217 (N_14217,N_14132,N_14160);
or U14218 (N_14218,N_14178,N_14152);
nand U14219 (N_14219,N_14080,N_14095);
nand U14220 (N_14220,N_14140,N_14134);
and U14221 (N_14221,N_14100,N_14158);
xor U14222 (N_14222,N_14128,N_14126);
or U14223 (N_14223,N_14084,N_14077);
nor U14224 (N_14224,N_14112,N_14033);
xor U14225 (N_14225,N_14050,N_14173);
or U14226 (N_14226,N_14041,N_14019);
or U14227 (N_14227,N_14043,N_14198);
nor U14228 (N_14228,N_14035,N_14008);
and U14229 (N_14229,N_14146,N_14096);
nor U14230 (N_14230,N_14109,N_14124);
or U14231 (N_14231,N_14138,N_14054);
nor U14232 (N_14232,N_14098,N_14172);
nand U14233 (N_14233,N_14118,N_14139);
nand U14234 (N_14234,N_14079,N_14067);
xor U14235 (N_14235,N_14087,N_14055);
or U14236 (N_14236,N_14039,N_14101);
and U14237 (N_14237,N_14192,N_14106);
nand U14238 (N_14238,N_14094,N_14047);
xnor U14239 (N_14239,N_14011,N_14194);
or U14240 (N_14240,N_14170,N_14155);
or U14241 (N_14241,N_14032,N_14120);
nor U14242 (N_14242,N_14075,N_14175);
xor U14243 (N_14243,N_14065,N_14196);
and U14244 (N_14244,N_14020,N_14105);
nor U14245 (N_14245,N_14148,N_14154);
nand U14246 (N_14246,N_14062,N_14168);
nor U14247 (N_14247,N_14006,N_14122);
or U14248 (N_14248,N_14010,N_14199);
nand U14249 (N_14249,N_14113,N_14009);
nor U14250 (N_14250,N_14185,N_14149);
xor U14251 (N_14251,N_14082,N_14026);
or U14252 (N_14252,N_14133,N_14029);
nor U14253 (N_14253,N_14048,N_14024);
xor U14254 (N_14254,N_14150,N_14186);
nand U14255 (N_14255,N_14184,N_14053);
xnor U14256 (N_14256,N_14057,N_14130);
nand U14257 (N_14257,N_14111,N_14001);
nand U14258 (N_14258,N_14071,N_14002);
and U14259 (N_14259,N_14072,N_14044);
and U14260 (N_14260,N_14049,N_14083);
xnor U14261 (N_14261,N_14003,N_14137);
nor U14262 (N_14262,N_14091,N_14157);
nor U14263 (N_14263,N_14069,N_14180);
nor U14264 (N_14264,N_14182,N_14090);
nor U14265 (N_14265,N_14007,N_14085);
and U14266 (N_14266,N_14166,N_14036);
or U14267 (N_14267,N_14015,N_14190);
nand U14268 (N_14268,N_14092,N_14108);
nand U14269 (N_14269,N_14115,N_14068);
or U14270 (N_14270,N_14021,N_14089);
xnor U14271 (N_14271,N_14119,N_14056);
nand U14272 (N_14272,N_14051,N_14161);
and U14273 (N_14273,N_14070,N_14012);
xor U14274 (N_14274,N_14121,N_14153);
nand U14275 (N_14275,N_14104,N_14191);
nand U14276 (N_14276,N_14156,N_14014);
nand U14277 (N_14277,N_14097,N_14144);
nor U14278 (N_14278,N_14159,N_14147);
nand U14279 (N_14279,N_14005,N_14016);
and U14280 (N_14280,N_14193,N_14164);
xnor U14281 (N_14281,N_14059,N_14063);
nor U14282 (N_14282,N_14129,N_14058);
nor U14283 (N_14283,N_14042,N_14103);
nor U14284 (N_14284,N_14017,N_14064);
nor U14285 (N_14285,N_14037,N_14107);
nor U14286 (N_14286,N_14086,N_14188);
nand U14287 (N_14287,N_14000,N_14141);
or U14288 (N_14288,N_14110,N_14099);
nor U14289 (N_14289,N_14114,N_14181);
xor U14290 (N_14290,N_14174,N_14169);
nand U14291 (N_14291,N_14022,N_14197);
or U14292 (N_14292,N_14151,N_14123);
or U14293 (N_14293,N_14066,N_14034);
xor U14294 (N_14294,N_14045,N_14145);
or U14295 (N_14295,N_14163,N_14183);
and U14296 (N_14296,N_14143,N_14189);
nand U14297 (N_14297,N_14040,N_14102);
or U14298 (N_14298,N_14025,N_14176);
xnor U14299 (N_14299,N_14078,N_14060);
xor U14300 (N_14300,N_14055,N_14196);
or U14301 (N_14301,N_14014,N_14170);
xnor U14302 (N_14302,N_14006,N_14171);
nand U14303 (N_14303,N_14130,N_14126);
nor U14304 (N_14304,N_14016,N_14073);
and U14305 (N_14305,N_14123,N_14021);
nand U14306 (N_14306,N_14100,N_14160);
nor U14307 (N_14307,N_14113,N_14061);
nand U14308 (N_14308,N_14163,N_14157);
xor U14309 (N_14309,N_14090,N_14128);
nor U14310 (N_14310,N_14183,N_14150);
xor U14311 (N_14311,N_14159,N_14019);
and U14312 (N_14312,N_14188,N_14198);
nor U14313 (N_14313,N_14180,N_14045);
or U14314 (N_14314,N_14022,N_14067);
nor U14315 (N_14315,N_14007,N_14122);
and U14316 (N_14316,N_14081,N_14073);
xor U14317 (N_14317,N_14114,N_14098);
and U14318 (N_14318,N_14052,N_14019);
nor U14319 (N_14319,N_14072,N_14000);
nor U14320 (N_14320,N_14008,N_14061);
and U14321 (N_14321,N_14198,N_14173);
xor U14322 (N_14322,N_14122,N_14167);
nor U14323 (N_14323,N_14077,N_14082);
or U14324 (N_14324,N_14102,N_14043);
nor U14325 (N_14325,N_14146,N_14095);
nor U14326 (N_14326,N_14137,N_14099);
and U14327 (N_14327,N_14167,N_14175);
and U14328 (N_14328,N_14030,N_14005);
xnor U14329 (N_14329,N_14044,N_14037);
and U14330 (N_14330,N_14067,N_14017);
nor U14331 (N_14331,N_14136,N_14091);
nand U14332 (N_14332,N_14031,N_14101);
xor U14333 (N_14333,N_14116,N_14192);
or U14334 (N_14334,N_14173,N_14153);
nor U14335 (N_14335,N_14148,N_14196);
xor U14336 (N_14336,N_14075,N_14023);
nand U14337 (N_14337,N_14081,N_14127);
nor U14338 (N_14338,N_14126,N_14067);
and U14339 (N_14339,N_14165,N_14143);
xor U14340 (N_14340,N_14077,N_14181);
nand U14341 (N_14341,N_14072,N_14131);
nor U14342 (N_14342,N_14049,N_14060);
nor U14343 (N_14343,N_14133,N_14073);
nand U14344 (N_14344,N_14145,N_14190);
xor U14345 (N_14345,N_14095,N_14104);
or U14346 (N_14346,N_14031,N_14110);
nor U14347 (N_14347,N_14049,N_14096);
and U14348 (N_14348,N_14140,N_14049);
nor U14349 (N_14349,N_14029,N_14037);
or U14350 (N_14350,N_14069,N_14153);
nor U14351 (N_14351,N_14080,N_14053);
or U14352 (N_14352,N_14025,N_14010);
or U14353 (N_14353,N_14074,N_14148);
and U14354 (N_14354,N_14097,N_14024);
nand U14355 (N_14355,N_14018,N_14027);
nor U14356 (N_14356,N_14068,N_14140);
xnor U14357 (N_14357,N_14054,N_14112);
nor U14358 (N_14358,N_14170,N_14068);
or U14359 (N_14359,N_14024,N_14030);
nor U14360 (N_14360,N_14000,N_14090);
nor U14361 (N_14361,N_14132,N_14017);
or U14362 (N_14362,N_14190,N_14184);
nand U14363 (N_14363,N_14088,N_14114);
nor U14364 (N_14364,N_14058,N_14068);
xor U14365 (N_14365,N_14020,N_14102);
nor U14366 (N_14366,N_14066,N_14008);
or U14367 (N_14367,N_14159,N_14094);
nand U14368 (N_14368,N_14133,N_14170);
xor U14369 (N_14369,N_14116,N_14078);
and U14370 (N_14370,N_14098,N_14047);
and U14371 (N_14371,N_14142,N_14067);
nand U14372 (N_14372,N_14072,N_14158);
xor U14373 (N_14373,N_14026,N_14169);
and U14374 (N_14374,N_14197,N_14186);
nand U14375 (N_14375,N_14129,N_14021);
nor U14376 (N_14376,N_14079,N_14166);
or U14377 (N_14377,N_14147,N_14146);
xor U14378 (N_14378,N_14078,N_14164);
or U14379 (N_14379,N_14196,N_14064);
and U14380 (N_14380,N_14104,N_14132);
or U14381 (N_14381,N_14117,N_14103);
or U14382 (N_14382,N_14168,N_14144);
nor U14383 (N_14383,N_14141,N_14056);
nor U14384 (N_14384,N_14119,N_14174);
nand U14385 (N_14385,N_14046,N_14017);
and U14386 (N_14386,N_14170,N_14057);
xor U14387 (N_14387,N_14126,N_14194);
and U14388 (N_14388,N_14183,N_14141);
or U14389 (N_14389,N_14184,N_14005);
nand U14390 (N_14390,N_14194,N_14049);
and U14391 (N_14391,N_14165,N_14097);
nor U14392 (N_14392,N_14020,N_14025);
xnor U14393 (N_14393,N_14026,N_14017);
or U14394 (N_14394,N_14154,N_14016);
nor U14395 (N_14395,N_14134,N_14161);
nand U14396 (N_14396,N_14178,N_14010);
nand U14397 (N_14397,N_14161,N_14185);
nor U14398 (N_14398,N_14191,N_14194);
xor U14399 (N_14399,N_14182,N_14065);
xnor U14400 (N_14400,N_14280,N_14389);
nor U14401 (N_14401,N_14218,N_14351);
and U14402 (N_14402,N_14301,N_14226);
xnor U14403 (N_14403,N_14263,N_14333);
nand U14404 (N_14404,N_14233,N_14317);
nand U14405 (N_14405,N_14216,N_14329);
nand U14406 (N_14406,N_14235,N_14270);
and U14407 (N_14407,N_14273,N_14386);
nand U14408 (N_14408,N_14350,N_14369);
nand U14409 (N_14409,N_14376,N_14248);
nand U14410 (N_14410,N_14289,N_14353);
xor U14411 (N_14411,N_14343,N_14236);
xnor U14412 (N_14412,N_14237,N_14272);
nor U14413 (N_14413,N_14340,N_14279);
nor U14414 (N_14414,N_14330,N_14394);
nor U14415 (N_14415,N_14268,N_14311);
xnor U14416 (N_14416,N_14284,N_14336);
or U14417 (N_14417,N_14368,N_14306);
or U14418 (N_14418,N_14282,N_14395);
or U14419 (N_14419,N_14231,N_14359);
nor U14420 (N_14420,N_14243,N_14352);
nand U14421 (N_14421,N_14335,N_14220);
nand U14422 (N_14422,N_14399,N_14206);
or U14423 (N_14423,N_14261,N_14348);
nand U14424 (N_14424,N_14371,N_14259);
nor U14425 (N_14425,N_14288,N_14363);
nand U14426 (N_14426,N_14377,N_14347);
xnor U14427 (N_14427,N_14240,N_14372);
nor U14428 (N_14428,N_14320,N_14360);
nand U14429 (N_14429,N_14365,N_14227);
xor U14430 (N_14430,N_14286,N_14315);
nor U14431 (N_14431,N_14208,N_14275);
and U14432 (N_14432,N_14278,N_14232);
xnor U14433 (N_14433,N_14387,N_14378);
or U14434 (N_14434,N_14205,N_14262);
nand U14435 (N_14435,N_14373,N_14228);
or U14436 (N_14436,N_14341,N_14374);
xor U14437 (N_14437,N_14221,N_14354);
xor U14438 (N_14438,N_14252,N_14287);
xnor U14439 (N_14439,N_14290,N_14210);
and U14440 (N_14440,N_14342,N_14307);
or U14441 (N_14441,N_14277,N_14309);
and U14442 (N_14442,N_14202,N_14222);
nor U14443 (N_14443,N_14382,N_14266);
nand U14444 (N_14444,N_14264,N_14349);
xor U14445 (N_14445,N_14209,N_14364);
nand U14446 (N_14446,N_14274,N_14249);
nand U14447 (N_14447,N_14383,N_14384);
nor U14448 (N_14448,N_14285,N_14283);
xor U14449 (N_14449,N_14267,N_14207);
and U14450 (N_14450,N_14219,N_14291);
xnor U14451 (N_14451,N_14358,N_14324);
and U14452 (N_14452,N_14215,N_14217);
and U14453 (N_14453,N_14246,N_14366);
nor U14454 (N_14454,N_14398,N_14303);
nor U14455 (N_14455,N_14325,N_14379);
xor U14456 (N_14456,N_14338,N_14299);
or U14457 (N_14457,N_14302,N_14362);
xnor U14458 (N_14458,N_14295,N_14388);
nand U14459 (N_14459,N_14241,N_14269);
and U14460 (N_14460,N_14229,N_14203);
xor U14461 (N_14461,N_14250,N_14391);
or U14462 (N_14462,N_14296,N_14213);
and U14463 (N_14463,N_14355,N_14326);
nand U14464 (N_14464,N_14392,N_14276);
xnor U14465 (N_14465,N_14201,N_14211);
nor U14466 (N_14466,N_14242,N_14367);
nand U14467 (N_14467,N_14230,N_14381);
and U14468 (N_14468,N_14223,N_14321);
nand U14469 (N_14469,N_14257,N_14254);
or U14470 (N_14470,N_14260,N_14316);
nor U14471 (N_14471,N_14370,N_14308);
xnor U14472 (N_14472,N_14253,N_14294);
nand U14473 (N_14473,N_14204,N_14298);
and U14474 (N_14474,N_14305,N_14380);
and U14475 (N_14475,N_14361,N_14234);
and U14476 (N_14476,N_14375,N_14281);
or U14477 (N_14477,N_14356,N_14334);
nor U14478 (N_14478,N_14346,N_14212);
or U14479 (N_14479,N_14245,N_14265);
xor U14480 (N_14480,N_14339,N_14393);
xnor U14481 (N_14481,N_14292,N_14297);
xnor U14482 (N_14482,N_14239,N_14323);
and U14483 (N_14483,N_14357,N_14238);
nor U14484 (N_14484,N_14300,N_14319);
or U14485 (N_14485,N_14327,N_14322);
or U14486 (N_14486,N_14214,N_14224);
nor U14487 (N_14487,N_14258,N_14337);
xnor U14488 (N_14488,N_14385,N_14304);
nand U14489 (N_14489,N_14200,N_14271);
xnor U14490 (N_14490,N_14345,N_14332);
and U14491 (N_14491,N_14293,N_14318);
and U14492 (N_14492,N_14314,N_14396);
xnor U14493 (N_14493,N_14225,N_14251);
xnor U14494 (N_14494,N_14255,N_14344);
nor U14495 (N_14495,N_14256,N_14312);
nand U14496 (N_14496,N_14328,N_14397);
xor U14497 (N_14497,N_14247,N_14313);
or U14498 (N_14498,N_14310,N_14390);
nand U14499 (N_14499,N_14331,N_14244);
nor U14500 (N_14500,N_14388,N_14389);
and U14501 (N_14501,N_14311,N_14362);
nand U14502 (N_14502,N_14257,N_14220);
xor U14503 (N_14503,N_14277,N_14221);
or U14504 (N_14504,N_14331,N_14371);
or U14505 (N_14505,N_14366,N_14255);
xor U14506 (N_14506,N_14381,N_14217);
nor U14507 (N_14507,N_14325,N_14262);
and U14508 (N_14508,N_14329,N_14274);
xnor U14509 (N_14509,N_14339,N_14205);
and U14510 (N_14510,N_14396,N_14261);
nand U14511 (N_14511,N_14216,N_14324);
nand U14512 (N_14512,N_14323,N_14367);
xor U14513 (N_14513,N_14351,N_14290);
or U14514 (N_14514,N_14274,N_14209);
or U14515 (N_14515,N_14283,N_14367);
nand U14516 (N_14516,N_14310,N_14328);
or U14517 (N_14517,N_14256,N_14218);
xor U14518 (N_14518,N_14267,N_14209);
and U14519 (N_14519,N_14292,N_14338);
xor U14520 (N_14520,N_14359,N_14216);
or U14521 (N_14521,N_14336,N_14282);
nand U14522 (N_14522,N_14230,N_14333);
or U14523 (N_14523,N_14389,N_14279);
xnor U14524 (N_14524,N_14278,N_14248);
nor U14525 (N_14525,N_14228,N_14279);
nor U14526 (N_14526,N_14363,N_14254);
or U14527 (N_14527,N_14214,N_14389);
xor U14528 (N_14528,N_14257,N_14288);
and U14529 (N_14529,N_14372,N_14324);
nand U14530 (N_14530,N_14369,N_14237);
and U14531 (N_14531,N_14259,N_14387);
xor U14532 (N_14532,N_14343,N_14312);
xor U14533 (N_14533,N_14364,N_14361);
xor U14534 (N_14534,N_14226,N_14251);
xor U14535 (N_14535,N_14268,N_14355);
nor U14536 (N_14536,N_14267,N_14321);
and U14537 (N_14537,N_14266,N_14252);
xnor U14538 (N_14538,N_14259,N_14365);
nand U14539 (N_14539,N_14247,N_14366);
or U14540 (N_14540,N_14335,N_14209);
nor U14541 (N_14541,N_14380,N_14349);
or U14542 (N_14542,N_14350,N_14280);
or U14543 (N_14543,N_14269,N_14395);
and U14544 (N_14544,N_14273,N_14327);
nand U14545 (N_14545,N_14237,N_14341);
or U14546 (N_14546,N_14206,N_14349);
and U14547 (N_14547,N_14251,N_14310);
xnor U14548 (N_14548,N_14246,N_14377);
xor U14549 (N_14549,N_14372,N_14367);
nand U14550 (N_14550,N_14323,N_14328);
nor U14551 (N_14551,N_14380,N_14358);
xnor U14552 (N_14552,N_14206,N_14398);
or U14553 (N_14553,N_14274,N_14206);
and U14554 (N_14554,N_14302,N_14294);
and U14555 (N_14555,N_14272,N_14279);
or U14556 (N_14556,N_14218,N_14241);
nor U14557 (N_14557,N_14344,N_14253);
xnor U14558 (N_14558,N_14302,N_14381);
and U14559 (N_14559,N_14291,N_14325);
or U14560 (N_14560,N_14332,N_14276);
and U14561 (N_14561,N_14232,N_14356);
or U14562 (N_14562,N_14293,N_14316);
xor U14563 (N_14563,N_14302,N_14257);
and U14564 (N_14564,N_14398,N_14346);
nand U14565 (N_14565,N_14241,N_14247);
nor U14566 (N_14566,N_14288,N_14224);
nor U14567 (N_14567,N_14294,N_14318);
and U14568 (N_14568,N_14379,N_14367);
nand U14569 (N_14569,N_14212,N_14303);
xor U14570 (N_14570,N_14253,N_14351);
nor U14571 (N_14571,N_14382,N_14294);
or U14572 (N_14572,N_14394,N_14366);
nand U14573 (N_14573,N_14372,N_14285);
or U14574 (N_14574,N_14381,N_14248);
nand U14575 (N_14575,N_14374,N_14201);
nand U14576 (N_14576,N_14204,N_14295);
and U14577 (N_14577,N_14339,N_14238);
nand U14578 (N_14578,N_14388,N_14270);
nor U14579 (N_14579,N_14372,N_14268);
nor U14580 (N_14580,N_14295,N_14359);
xnor U14581 (N_14581,N_14288,N_14354);
nand U14582 (N_14582,N_14274,N_14382);
and U14583 (N_14583,N_14212,N_14202);
xnor U14584 (N_14584,N_14320,N_14222);
xnor U14585 (N_14585,N_14335,N_14334);
nor U14586 (N_14586,N_14225,N_14299);
xor U14587 (N_14587,N_14209,N_14330);
nand U14588 (N_14588,N_14274,N_14235);
nor U14589 (N_14589,N_14371,N_14277);
xor U14590 (N_14590,N_14340,N_14319);
nand U14591 (N_14591,N_14343,N_14333);
nand U14592 (N_14592,N_14294,N_14224);
xnor U14593 (N_14593,N_14226,N_14259);
or U14594 (N_14594,N_14352,N_14353);
nand U14595 (N_14595,N_14206,N_14216);
nand U14596 (N_14596,N_14357,N_14314);
xnor U14597 (N_14597,N_14218,N_14378);
nor U14598 (N_14598,N_14206,N_14306);
and U14599 (N_14599,N_14345,N_14219);
xor U14600 (N_14600,N_14594,N_14518);
nand U14601 (N_14601,N_14473,N_14572);
xnor U14602 (N_14602,N_14549,N_14402);
or U14603 (N_14603,N_14580,N_14438);
nand U14604 (N_14604,N_14474,N_14581);
xor U14605 (N_14605,N_14552,N_14406);
nor U14606 (N_14606,N_14464,N_14584);
xor U14607 (N_14607,N_14443,N_14528);
xor U14608 (N_14608,N_14453,N_14467);
or U14609 (N_14609,N_14475,N_14423);
or U14610 (N_14610,N_14511,N_14489);
nor U14611 (N_14611,N_14455,N_14405);
nor U14612 (N_14612,N_14400,N_14494);
and U14613 (N_14613,N_14403,N_14483);
and U14614 (N_14614,N_14451,N_14526);
nor U14615 (N_14615,N_14519,N_14414);
nand U14616 (N_14616,N_14424,N_14454);
nand U14617 (N_14617,N_14450,N_14512);
and U14618 (N_14618,N_14431,N_14418);
and U14619 (N_14619,N_14429,N_14478);
nor U14620 (N_14620,N_14509,N_14506);
xor U14621 (N_14621,N_14505,N_14575);
nor U14622 (N_14622,N_14462,N_14415);
nor U14623 (N_14623,N_14550,N_14411);
or U14624 (N_14624,N_14493,N_14485);
xor U14625 (N_14625,N_14576,N_14432);
xor U14626 (N_14626,N_14407,N_14487);
and U14627 (N_14627,N_14466,N_14570);
nand U14628 (N_14628,N_14535,N_14410);
nor U14629 (N_14629,N_14434,N_14554);
or U14630 (N_14630,N_14540,N_14515);
nand U14631 (N_14631,N_14555,N_14579);
nand U14632 (N_14632,N_14520,N_14477);
or U14633 (N_14633,N_14436,N_14404);
and U14634 (N_14634,N_14561,N_14503);
nand U14635 (N_14635,N_14583,N_14481);
nand U14636 (N_14636,N_14521,N_14551);
nand U14637 (N_14637,N_14456,N_14589);
nor U14638 (N_14638,N_14470,N_14445);
nand U14639 (N_14639,N_14504,N_14544);
and U14640 (N_14640,N_14558,N_14452);
or U14641 (N_14641,N_14471,N_14560);
or U14642 (N_14642,N_14476,N_14529);
or U14643 (N_14643,N_14536,N_14537);
or U14644 (N_14644,N_14448,N_14587);
and U14645 (N_14645,N_14413,N_14500);
or U14646 (N_14646,N_14538,N_14440);
or U14647 (N_14647,N_14543,N_14533);
xor U14648 (N_14648,N_14523,N_14495);
or U14649 (N_14649,N_14490,N_14524);
and U14650 (N_14650,N_14590,N_14507);
and U14651 (N_14651,N_14522,N_14428);
xor U14652 (N_14652,N_14530,N_14482);
and U14653 (N_14653,N_14463,N_14565);
xor U14654 (N_14654,N_14573,N_14574);
or U14655 (N_14655,N_14553,N_14421);
nor U14656 (N_14656,N_14510,N_14468);
xor U14657 (N_14657,N_14599,N_14401);
nand U14658 (N_14658,N_14571,N_14567);
and U14659 (N_14659,N_14484,N_14562);
and U14660 (N_14660,N_14514,N_14585);
or U14661 (N_14661,N_14472,N_14556);
nor U14662 (N_14662,N_14559,N_14598);
or U14663 (N_14663,N_14591,N_14525);
or U14664 (N_14664,N_14419,N_14435);
xnor U14665 (N_14665,N_14501,N_14449);
nand U14666 (N_14666,N_14433,N_14508);
nor U14667 (N_14667,N_14460,N_14444);
nor U14668 (N_14668,N_14442,N_14517);
and U14669 (N_14669,N_14568,N_14408);
nor U14670 (N_14670,N_14513,N_14499);
or U14671 (N_14671,N_14595,N_14486);
or U14672 (N_14672,N_14469,N_14465);
nand U14673 (N_14673,N_14479,N_14497);
xor U14674 (N_14674,N_14488,N_14531);
nor U14675 (N_14675,N_14557,N_14546);
or U14676 (N_14676,N_14541,N_14564);
or U14677 (N_14677,N_14545,N_14437);
xor U14678 (N_14678,N_14417,N_14439);
xnor U14679 (N_14679,N_14578,N_14457);
or U14680 (N_14680,N_14597,N_14427);
or U14681 (N_14681,N_14412,N_14548);
or U14682 (N_14682,N_14593,N_14532);
xnor U14683 (N_14683,N_14542,N_14498);
or U14684 (N_14684,N_14592,N_14534);
nand U14685 (N_14685,N_14492,N_14430);
xnor U14686 (N_14686,N_14516,N_14426);
and U14687 (N_14687,N_14447,N_14461);
or U14688 (N_14688,N_14586,N_14420);
nor U14689 (N_14689,N_14416,N_14458);
nand U14690 (N_14690,N_14588,N_14539);
or U14691 (N_14691,N_14502,N_14582);
or U14692 (N_14692,N_14569,N_14566);
nor U14693 (N_14693,N_14425,N_14422);
or U14694 (N_14694,N_14409,N_14547);
or U14695 (N_14695,N_14491,N_14527);
xor U14696 (N_14696,N_14480,N_14496);
nor U14697 (N_14697,N_14563,N_14577);
nor U14698 (N_14698,N_14596,N_14446);
and U14699 (N_14699,N_14441,N_14459);
or U14700 (N_14700,N_14461,N_14561);
and U14701 (N_14701,N_14462,N_14425);
and U14702 (N_14702,N_14525,N_14415);
and U14703 (N_14703,N_14546,N_14441);
nor U14704 (N_14704,N_14444,N_14446);
xnor U14705 (N_14705,N_14542,N_14556);
or U14706 (N_14706,N_14542,N_14503);
xnor U14707 (N_14707,N_14548,N_14476);
xor U14708 (N_14708,N_14425,N_14500);
or U14709 (N_14709,N_14477,N_14542);
nand U14710 (N_14710,N_14426,N_14506);
and U14711 (N_14711,N_14520,N_14459);
or U14712 (N_14712,N_14418,N_14474);
nand U14713 (N_14713,N_14583,N_14448);
or U14714 (N_14714,N_14408,N_14454);
xnor U14715 (N_14715,N_14598,N_14552);
nor U14716 (N_14716,N_14537,N_14409);
and U14717 (N_14717,N_14450,N_14400);
or U14718 (N_14718,N_14469,N_14475);
or U14719 (N_14719,N_14499,N_14542);
nor U14720 (N_14720,N_14465,N_14547);
xor U14721 (N_14721,N_14419,N_14517);
nor U14722 (N_14722,N_14525,N_14489);
or U14723 (N_14723,N_14556,N_14429);
nor U14724 (N_14724,N_14576,N_14457);
nand U14725 (N_14725,N_14559,N_14576);
or U14726 (N_14726,N_14486,N_14446);
and U14727 (N_14727,N_14581,N_14454);
nand U14728 (N_14728,N_14446,N_14532);
nand U14729 (N_14729,N_14578,N_14533);
nor U14730 (N_14730,N_14521,N_14504);
nand U14731 (N_14731,N_14464,N_14403);
nand U14732 (N_14732,N_14532,N_14490);
and U14733 (N_14733,N_14547,N_14430);
or U14734 (N_14734,N_14522,N_14536);
nand U14735 (N_14735,N_14475,N_14559);
nand U14736 (N_14736,N_14438,N_14402);
and U14737 (N_14737,N_14507,N_14500);
or U14738 (N_14738,N_14570,N_14478);
or U14739 (N_14739,N_14441,N_14525);
nor U14740 (N_14740,N_14404,N_14485);
nor U14741 (N_14741,N_14438,N_14458);
xor U14742 (N_14742,N_14468,N_14412);
xor U14743 (N_14743,N_14514,N_14526);
and U14744 (N_14744,N_14406,N_14435);
nand U14745 (N_14745,N_14559,N_14508);
nor U14746 (N_14746,N_14471,N_14443);
nor U14747 (N_14747,N_14448,N_14547);
or U14748 (N_14748,N_14522,N_14434);
or U14749 (N_14749,N_14560,N_14475);
nand U14750 (N_14750,N_14492,N_14459);
nand U14751 (N_14751,N_14562,N_14488);
and U14752 (N_14752,N_14423,N_14507);
nand U14753 (N_14753,N_14484,N_14513);
and U14754 (N_14754,N_14476,N_14588);
or U14755 (N_14755,N_14475,N_14457);
nor U14756 (N_14756,N_14401,N_14422);
nor U14757 (N_14757,N_14513,N_14523);
nor U14758 (N_14758,N_14440,N_14470);
or U14759 (N_14759,N_14420,N_14575);
nor U14760 (N_14760,N_14598,N_14488);
and U14761 (N_14761,N_14511,N_14515);
or U14762 (N_14762,N_14465,N_14558);
nor U14763 (N_14763,N_14535,N_14574);
nor U14764 (N_14764,N_14422,N_14481);
or U14765 (N_14765,N_14584,N_14426);
or U14766 (N_14766,N_14560,N_14586);
nand U14767 (N_14767,N_14522,N_14594);
and U14768 (N_14768,N_14583,N_14534);
nand U14769 (N_14769,N_14438,N_14522);
nor U14770 (N_14770,N_14423,N_14548);
or U14771 (N_14771,N_14593,N_14465);
nand U14772 (N_14772,N_14400,N_14598);
xor U14773 (N_14773,N_14553,N_14489);
or U14774 (N_14774,N_14463,N_14528);
and U14775 (N_14775,N_14458,N_14492);
or U14776 (N_14776,N_14476,N_14519);
or U14777 (N_14777,N_14407,N_14503);
and U14778 (N_14778,N_14560,N_14573);
nand U14779 (N_14779,N_14437,N_14497);
and U14780 (N_14780,N_14545,N_14458);
nand U14781 (N_14781,N_14560,N_14424);
nor U14782 (N_14782,N_14407,N_14526);
nor U14783 (N_14783,N_14414,N_14514);
or U14784 (N_14784,N_14550,N_14532);
and U14785 (N_14785,N_14509,N_14487);
or U14786 (N_14786,N_14543,N_14484);
nand U14787 (N_14787,N_14474,N_14409);
and U14788 (N_14788,N_14594,N_14589);
nand U14789 (N_14789,N_14548,N_14479);
or U14790 (N_14790,N_14442,N_14501);
xor U14791 (N_14791,N_14405,N_14427);
nor U14792 (N_14792,N_14473,N_14598);
xor U14793 (N_14793,N_14437,N_14487);
or U14794 (N_14794,N_14477,N_14447);
nand U14795 (N_14795,N_14549,N_14566);
nor U14796 (N_14796,N_14575,N_14579);
or U14797 (N_14797,N_14594,N_14503);
xor U14798 (N_14798,N_14562,N_14590);
nor U14799 (N_14799,N_14498,N_14463);
or U14800 (N_14800,N_14623,N_14659);
nand U14801 (N_14801,N_14642,N_14680);
nand U14802 (N_14802,N_14649,N_14648);
nand U14803 (N_14803,N_14636,N_14613);
xnor U14804 (N_14804,N_14653,N_14669);
and U14805 (N_14805,N_14717,N_14715);
xor U14806 (N_14806,N_14671,N_14691);
nor U14807 (N_14807,N_14782,N_14673);
and U14808 (N_14808,N_14641,N_14720);
nor U14809 (N_14809,N_14739,N_14651);
nand U14810 (N_14810,N_14703,N_14719);
xnor U14811 (N_14811,N_14606,N_14675);
nand U14812 (N_14812,N_14797,N_14751);
xnor U14813 (N_14813,N_14620,N_14778);
and U14814 (N_14814,N_14652,N_14764);
nor U14815 (N_14815,N_14650,N_14618);
xnor U14816 (N_14816,N_14661,N_14744);
nand U14817 (N_14817,N_14713,N_14707);
xnor U14818 (N_14818,N_14617,N_14645);
or U14819 (N_14819,N_14779,N_14733);
or U14820 (N_14820,N_14616,N_14756);
and U14821 (N_14821,N_14741,N_14759);
and U14822 (N_14822,N_14631,N_14712);
nor U14823 (N_14823,N_14781,N_14604);
or U14824 (N_14824,N_14693,N_14692);
xor U14825 (N_14825,N_14742,N_14683);
and U14826 (N_14826,N_14783,N_14704);
xnor U14827 (N_14827,N_14672,N_14608);
nand U14828 (N_14828,N_14601,N_14714);
nor U14829 (N_14829,N_14646,N_14621);
nor U14830 (N_14830,N_14746,N_14767);
nor U14831 (N_14831,N_14774,N_14619);
nor U14832 (N_14832,N_14789,N_14634);
or U14833 (N_14833,N_14777,N_14793);
or U14834 (N_14834,N_14718,N_14755);
xnor U14835 (N_14835,N_14772,N_14788);
nand U14836 (N_14836,N_14702,N_14644);
nand U14837 (N_14837,N_14635,N_14610);
nor U14838 (N_14838,N_14786,N_14799);
xnor U14839 (N_14839,N_14624,N_14766);
xnor U14840 (N_14840,N_14763,N_14600);
xor U14841 (N_14841,N_14625,N_14709);
or U14842 (N_14842,N_14734,N_14657);
xnor U14843 (N_14843,N_14769,N_14787);
nor U14844 (N_14844,N_14710,N_14681);
nand U14845 (N_14845,N_14666,N_14678);
or U14846 (N_14846,N_14637,N_14773);
and U14847 (N_14847,N_14665,N_14785);
nor U14848 (N_14848,N_14728,N_14761);
nor U14849 (N_14849,N_14706,N_14632);
xnor U14850 (N_14850,N_14737,N_14768);
xnor U14851 (N_14851,N_14726,N_14655);
nor U14852 (N_14852,N_14775,N_14745);
or U14853 (N_14853,N_14663,N_14722);
xor U14854 (N_14854,N_14615,N_14725);
nand U14855 (N_14855,N_14627,N_14750);
and U14856 (N_14856,N_14790,N_14796);
or U14857 (N_14857,N_14607,N_14695);
and U14858 (N_14858,N_14730,N_14727);
nand U14859 (N_14859,N_14694,N_14743);
and U14860 (N_14860,N_14723,N_14614);
xor U14861 (N_14861,N_14740,N_14708);
nor U14862 (N_14862,N_14749,N_14747);
and U14863 (N_14863,N_14667,N_14609);
and U14864 (N_14864,N_14699,N_14762);
nand U14865 (N_14865,N_14753,N_14687);
nor U14866 (N_14866,N_14674,N_14629);
nand U14867 (N_14867,N_14738,N_14690);
xor U14868 (N_14868,N_14603,N_14679);
xnor U14869 (N_14869,N_14705,N_14721);
and U14870 (N_14870,N_14752,N_14792);
and U14871 (N_14871,N_14688,N_14780);
xnor U14872 (N_14872,N_14791,N_14602);
nand U14873 (N_14873,N_14732,N_14628);
nand U14874 (N_14874,N_14622,N_14757);
and U14875 (N_14875,N_14668,N_14731);
nand U14876 (N_14876,N_14689,N_14776);
nand U14877 (N_14877,N_14700,N_14748);
and U14878 (N_14878,N_14660,N_14685);
xor U14879 (N_14879,N_14626,N_14736);
nand U14880 (N_14880,N_14770,N_14771);
nor U14881 (N_14881,N_14638,N_14754);
and U14882 (N_14882,N_14654,N_14729);
xnor U14883 (N_14883,N_14698,N_14765);
nand U14884 (N_14884,N_14611,N_14682);
or U14885 (N_14885,N_14633,N_14670);
nand U14886 (N_14886,N_14664,N_14795);
or U14887 (N_14887,N_14735,N_14784);
or U14888 (N_14888,N_14760,N_14716);
xor U14889 (N_14889,N_14686,N_14630);
nand U14890 (N_14890,N_14758,N_14647);
or U14891 (N_14891,N_14612,N_14639);
and U14892 (N_14892,N_14684,N_14724);
and U14893 (N_14893,N_14658,N_14677);
nand U14894 (N_14894,N_14662,N_14697);
nand U14895 (N_14895,N_14640,N_14656);
nand U14896 (N_14896,N_14643,N_14696);
xnor U14897 (N_14897,N_14711,N_14676);
nand U14898 (N_14898,N_14701,N_14605);
nor U14899 (N_14899,N_14798,N_14794);
and U14900 (N_14900,N_14735,N_14661);
or U14901 (N_14901,N_14659,N_14701);
xor U14902 (N_14902,N_14780,N_14759);
nand U14903 (N_14903,N_14714,N_14672);
xnor U14904 (N_14904,N_14795,N_14628);
or U14905 (N_14905,N_14657,N_14712);
xnor U14906 (N_14906,N_14759,N_14604);
and U14907 (N_14907,N_14774,N_14648);
xor U14908 (N_14908,N_14651,N_14610);
nor U14909 (N_14909,N_14620,N_14630);
nand U14910 (N_14910,N_14618,N_14752);
nand U14911 (N_14911,N_14754,N_14764);
xor U14912 (N_14912,N_14732,N_14784);
nor U14913 (N_14913,N_14639,N_14688);
nand U14914 (N_14914,N_14741,N_14726);
xnor U14915 (N_14915,N_14627,N_14758);
or U14916 (N_14916,N_14620,N_14674);
and U14917 (N_14917,N_14604,N_14621);
xnor U14918 (N_14918,N_14789,N_14651);
and U14919 (N_14919,N_14600,N_14793);
nand U14920 (N_14920,N_14628,N_14624);
xor U14921 (N_14921,N_14639,N_14760);
and U14922 (N_14922,N_14676,N_14607);
and U14923 (N_14923,N_14644,N_14611);
nand U14924 (N_14924,N_14616,N_14691);
nor U14925 (N_14925,N_14643,N_14693);
and U14926 (N_14926,N_14653,N_14773);
nand U14927 (N_14927,N_14635,N_14729);
and U14928 (N_14928,N_14632,N_14736);
nor U14929 (N_14929,N_14641,N_14619);
and U14930 (N_14930,N_14668,N_14606);
nor U14931 (N_14931,N_14787,N_14754);
or U14932 (N_14932,N_14752,N_14757);
nand U14933 (N_14933,N_14785,N_14602);
or U14934 (N_14934,N_14608,N_14658);
and U14935 (N_14935,N_14607,N_14617);
and U14936 (N_14936,N_14636,N_14795);
or U14937 (N_14937,N_14653,N_14687);
xnor U14938 (N_14938,N_14635,N_14659);
nand U14939 (N_14939,N_14615,N_14706);
nand U14940 (N_14940,N_14686,N_14791);
or U14941 (N_14941,N_14655,N_14656);
or U14942 (N_14942,N_14642,N_14638);
or U14943 (N_14943,N_14674,N_14639);
xnor U14944 (N_14944,N_14764,N_14759);
and U14945 (N_14945,N_14652,N_14610);
nor U14946 (N_14946,N_14753,N_14627);
and U14947 (N_14947,N_14628,N_14780);
nor U14948 (N_14948,N_14771,N_14696);
and U14949 (N_14949,N_14608,N_14685);
or U14950 (N_14950,N_14667,N_14691);
nand U14951 (N_14951,N_14617,N_14628);
nor U14952 (N_14952,N_14792,N_14637);
or U14953 (N_14953,N_14661,N_14728);
or U14954 (N_14954,N_14655,N_14611);
and U14955 (N_14955,N_14793,N_14772);
or U14956 (N_14956,N_14667,N_14692);
xnor U14957 (N_14957,N_14787,N_14619);
nor U14958 (N_14958,N_14722,N_14655);
xnor U14959 (N_14959,N_14646,N_14735);
or U14960 (N_14960,N_14692,N_14615);
and U14961 (N_14961,N_14613,N_14626);
nand U14962 (N_14962,N_14782,N_14770);
nor U14963 (N_14963,N_14606,N_14676);
nand U14964 (N_14964,N_14626,N_14776);
nand U14965 (N_14965,N_14767,N_14726);
and U14966 (N_14966,N_14665,N_14685);
nor U14967 (N_14967,N_14699,N_14735);
xor U14968 (N_14968,N_14729,N_14637);
nand U14969 (N_14969,N_14646,N_14669);
nand U14970 (N_14970,N_14638,N_14614);
nand U14971 (N_14971,N_14711,N_14741);
xor U14972 (N_14972,N_14681,N_14768);
nor U14973 (N_14973,N_14716,N_14708);
nand U14974 (N_14974,N_14700,N_14638);
nor U14975 (N_14975,N_14792,N_14751);
xor U14976 (N_14976,N_14609,N_14747);
xnor U14977 (N_14977,N_14731,N_14630);
nand U14978 (N_14978,N_14697,N_14710);
and U14979 (N_14979,N_14731,N_14632);
and U14980 (N_14980,N_14683,N_14685);
nor U14981 (N_14981,N_14608,N_14774);
and U14982 (N_14982,N_14687,N_14738);
nor U14983 (N_14983,N_14797,N_14643);
and U14984 (N_14984,N_14655,N_14721);
nor U14985 (N_14985,N_14683,N_14761);
or U14986 (N_14986,N_14788,N_14787);
or U14987 (N_14987,N_14682,N_14606);
nand U14988 (N_14988,N_14751,N_14609);
xor U14989 (N_14989,N_14668,N_14624);
nor U14990 (N_14990,N_14691,N_14647);
nor U14991 (N_14991,N_14688,N_14774);
or U14992 (N_14992,N_14695,N_14751);
xnor U14993 (N_14993,N_14658,N_14757);
xor U14994 (N_14994,N_14723,N_14703);
xor U14995 (N_14995,N_14621,N_14652);
xor U14996 (N_14996,N_14649,N_14753);
nand U14997 (N_14997,N_14795,N_14730);
xnor U14998 (N_14998,N_14681,N_14786);
xnor U14999 (N_14999,N_14637,N_14655);
xnor UO_0 (O_0,N_14842,N_14830);
or UO_1 (O_1,N_14839,N_14858);
nand UO_2 (O_2,N_14946,N_14992);
or UO_3 (O_3,N_14914,N_14827);
or UO_4 (O_4,N_14998,N_14950);
and UO_5 (O_5,N_14973,N_14818);
nand UO_6 (O_6,N_14942,N_14855);
nand UO_7 (O_7,N_14910,N_14829);
or UO_8 (O_8,N_14989,N_14902);
nor UO_9 (O_9,N_14895,N_14890);
nor UO_10 (O_10,N_14862,N_14817);
nand UO_11 (O_11,N_14835,N_14812);
xor UO_12 (O_12,N_14918,N_14877);
or UO_13 (O_13,N_14800,N_14948);
nand UO_14 (O_14,N_14894,N_14899);
nand UO_15 (O_15,N_14924,N_14898);
or UO_16 (O_16,N_14841,N_14849);
nor UO_17 (O_17,N_14907,N_14937);
and UO_18 (O_18,N_14883,N_14994);
or UO_19 (O_19,N_14867,N_14887);
and UO_20 (O_20,N_14878,N_14853);
nor UO_21 (O_21,N_14923,N_14951);
or UO_22 (O_22,N_14963,N_14856);
or UO_23 (O_23,N_14896,N_14879);
or UO_24 (O_24,N_14947,N_14845);
nand UO_25 (O_25,N_14808,N_14873);
or UO_26 (O_26,N_14881,N_14913);
nand UO_27 (O_27,N_14810,N_14866);
and UO_28 (O_28,N_14997,N_14813);
xor UO_29 (O_29,N_14885,N_14943);
nand UO_30 (O_30,N_14945,N_14995);
or UO_31 (O_31,N_14884,N_14912);
nor UO_32 (O_32,N_14892,N_14931);
nand UO_33 (O_33,N_14876,N_14875);
nand UO_34 (O_34,N_14929,N_14916);
nor UO_35 (O_35,N_14982,N_14964);
nand UO_36 (O_36,N_14968,N_14960);
xnor UO_37 (O_37,N_14903,N_14880);
nand UO_38 (O_38,N_14889,N_14865);
nand UO_39 (O_39,N_14920,N_14906);
or UO_40 (O_40,N_14940,N_14836);
xnor UO_41 (O_41,N_14958,N_14979);
or UO_42 (O_42,N_14847,N_14869);
nand UO_43 (O_43,N_14850,N_14944);
nor UO_44 (O_44,N_14863,N_14868);
and UO_45 (O_45,N_14932,N_14922);
nand UO_46 (O_46,N_14949,N_14915);
nor UO_47 (O_47,N_14919,N_14823);
nand UO_48 (O_48,N_14872,N_14811);
and UO_49 (O_49,N_14807,N_14831);
and UO_50 (O_50,N_14972,N_14983);
nand UO_51 (O_51,N_14926,N_14870);
or UO_52 (O_52,N_14819,N_14956);
and UO_53 (O_53,N_14806,N_14864);
nand UO_54 (O_54,N_14837,N_14952);
nand UO_55 (O_55,N_14985,N_14959);
nand UO_56 (O_56,N_14993,N_14976);
xnor UO_57 (O_57,N_14891,N_14961);
nor UO_58 (O_58,N_14834,N_14996);
or UO_59 (O_59,N_14938,N_14824);
or UO_60 (O_60,N_14802,N_14954);
or UO_61 (O_61,N_14804,N_14861);
nor UO_62 (O_62,N_14953,N_14874);
xnor UO_63 (O_63,N_14848,N_14888);
nor UO_64 (O_64,N_14846,N_14820);
or UO_65 (O_65,N_14816,N_14905);
and UO_66 (O_66,N_14901,N_14822);
and UO_67 (O_67,N_14977,N_14984);
or UO_68 (O_68,N_14809,N_14917);
and UO_69 (O_69,N_14814,N_14854);
and UO_70 (O_70,N_14925,N_14967);
nand UO_71 (O_71,N_14936,N_14978);
and UO_72 (O_72,N_14908,N_14957);
and UO_73 (O_73,N_14962,N_14921);
and UO_74 (O_74,N_14840,N_14999);
or UO_75 (O_75,N_14933,N_14860);
nor UO_76 (O_76,N_14927,N_14990);
nand UO_77 (O_77,N_14904,N_14965);
nand UO_78 (O_78,N_14971,N_14975);
or UO_79 (O_79,N_14871,N_14844);
xor UO_80 (O_80,N_14935,N_14882);
xnor UO_81 (O_81,N_14886,N_14939);
nor UO_82 (O_82,N_14988,N_14930);
nand UO_83 (O_83,N_14851,N_14838);
xor UO_84 (O_84,N_14986,N_14909);
and UO_85 (O_85,N_14826,N_14859);
nand UO_86 (O_86,N_14974,N_14815);
or UO_87 (O_87,N_14928,N_14991);
or UO_88 (O_88,N_14934,N_14828);
xnor UO_89 (O_89,N_14805,N_14900);
or UO_90 (O_90,N_14857,N_14966);
or UO_91 (O_91,N_14832,N_14843);
or UO_92 (O_92,N_14833,N_14801);
and UO_93 (O_93,N_14897,N_14852);
and UO_94 (O_94,N_14825,N_14969);
nand UO_95 (O_95,N_14987,N_14980);
xnor UO_96 (O_96,N_14955,N_14803);
nor UO_97 (O_97,N_14941,N_14911);
or UO_98 (O_98,N_14970,N_14981);
nand UO_99 (O_99,N_14821,N_14893);
or UO_100 (O_100,N_14972,N_14919);
nor UO_101 (O_101,N_14864,N_14926);
nor UO_102 (O_102,N_14854,N_14989);
nand UO_103 (O_103,N_14862,N_14948);
nand UO_104 (O_104,N_14851,N_14819);
nand UO_105 (O_105,N_14810,N_14970);
xnor UO_106 (O_106,N_14906,N_14953);
and UO_107 (O_107,N_14850,N_14864);
nor UO_108 (O_108,N_14901,N_14975);
or UO_109 (O_109,N_14803,N_14976);
nand UO_110 (O_110,N_14940,N_14892);
nor UO_111 (O_111,N_14944,N_14966);
and UO_112 (O_112,N_14990,N_14953);
nand UO_113 (O_113,N_14811,N_14971);
nand UO_114 (O_114,N_14933,N_14996);
xor UO_115 (O_115,N_14977,N_14987);
nor UO_116 (O_116,N_14829,N_14999);
or UO_117 (O_117,N_14935,N_14934);
xor UO_118 (O_118,N_14812,N_14883);
nor UO_119 (O_119,N_14954,N_14817);
nand UO_120 (O_120,N_14865,N_14994);
and UO_121 (O_121,N_14929,N_14812);
or UO_122 (O_122,N_14928,N_14959);
nand UO_123 (O_123,N_14874,N_14999);
xor UO_124 (O_124,N_14852,N_14881);
xor UO_125 (O_125,N_14840,N_14867);
xnor UO_126 (O_126,N_14930,N_14971);
and UO_127 (O_127,N_14960,N_14809);
nand UO_128 (O_128,N_14811,N_14888);
xnor UO_129 (O_129,N_14810,N_14832);
xor UO_130 (O_130,N_14876,N_14936);
nand UO_131 (O_131,N_14845,N_14916);
or UO_132 (O_132,N_14866,N_14946);
nand UO_133 (O_133,N_14885,N_14929);
xnor UO_134 (O_134,N_14912,N_14850);
xnor UO_135 (O_135,N_14989,N_14858);
nand UO_136 (O_136,N_14970,N_14880);
nor UO_137 (O_137,N_14994,N_14885);
and UO_138 (O_138,N_14973,N_14862);
nand UO_139 (O_139,N_14987,N_14862);
nor UO_140 (O_140,N_14906,N_14849);
xor UO_141 (O_141,N_14857,N_14961);
and UO_142 (O_142,N_14802,N_14970);
nand UO_143 (O_143,N_14933,N_14800);
nor UO_144 (O_144,N_14918,N_14819);
nor UO_145 (O_145,N_14877,N_14928);
nand UO_146 (O_146,N_14815,N_14915);
xor UO_147 (O_147,N_14996,N_14995);
nor UO_148 (O_148,N_14898,N_14938);
nand UO_149 (O_149,N_14962,N_14922);
nand UO_150 (O_150,N_14814,N_14862);
nor UO_151 (O_151,N_14927,N_14815);
nand UO_152 (O_152,N_14880,N_14923);
nor UO_153 (O_153,N_14813,N_14973);
and UO_154 (O_154,N_14922,N_14909);
xnor UO_155 (O_155,N_14952,N_14915);
nand UO_156 (O_156,N_14904,N_14910);
nor UO_157 (O_157,N_14993,N_14980);
nor UO_158 (O_158,N_14838,N_14803);
or UO_159 (O_159,N_14808,N_14935);
and UO_160 (O_160,N_14803,N_14866);
xnor UO_161 (O_161,N_14839,N_14826);
or UO_162 (O_162,N_14923,N_14830);
nand UO_163 (O_163,N_14965,N_14858);
or UO_164 (O_164,N_14904,N_14816);
nand UO_165 (O_165,N_14943,N_14944);
and UO_166 (O_166,N_14892,N_14810);
nor UO_167 (O_167,N_14973,N_14841);
nand UO_168 (O_168,N_14979,N_14996);
and UO_169 (O_169,N_14882,N_14861);
or UO_170 (O_170,N_14861,N_14968);
nand UO_171 (O_171,N_14857,N_14831);
xor UO_172 (O_172,N_14800,N_14985);
xnor UO_173 (O_173,N_14981,N_14815);
nor UO_174 (O_174,N_14801,N_14959);
nor UO_175 (O_175,N_14882,N_14808);
nand UO_176 (O_176,N_14830,N_14858);
nor UO_177 (O_177,N_14836,N_14993);
nor UO_178 (O_178,N_14900,N_14982);
nand UO_179 (O_179,N_14835,N_14842);
and UO_180 (O_180,N_14984,N_14908);
and UO_181 (O_181,N_14868,N_14927);
or UO_182 (O_182,N_14891,N_14809);
xor UO_183 (O_183,N_14800,N_14889);
nor UO_184 (O_184,N_14822,N_14993);
xor UO_185 (O_185,N_14836,N_14870);
nor UO_186 (O_186,N_14853,N_14918);
nand UO_187 (O_187,N_14862,N_14811);
nand UO_188 (O_188,N_14899,N_14839);
or UO_189 (O_189,N_14822,N_14882);
and UO_190 (O_190,N_14871,N_14818);
nor UO_191 (O_191,N_14943,N_14863);
xnor UO_192 (O_192,N_14882,N_14972);
nor UO_193 (O_193,N_14881,N_14933);
and UO_194 (O_194,N_14912,N_14878);
or UO_195 (O_195,N_14936,N_14855);
and UO_196 (O_196,N_14847,N_14839);
xor UO_197 (O_197,N_14812,N_14944);
nor UO_198 (O_198,N_14959,N_14927);
or UO_199 (O_199,N_14972,N_14904);
or UO_200 (O_200,N_14909,N_14846);
xor UO_201 (O_201,N_14884,N_14963);
or UO_202 (O_202,N_14822,N_14906);
or UO_203 (O_203,N_14835,N_14825);
or UO_204 (O_204,N_14803,N_14855);
or UO_205 (O_205,N_14877,N_14952);
and UO_206 (O_206,N_14965,N_14897);
nand UO_207 (O_207,N_14852,N_14900);
nor UO_208 (O_208,N_14843,N_14943);
xnor UO_209 (O_209,N_14887,N_14849);
and UO_210 (O_210,N_14948,N_14868);
and UO_211 (O_211,N_14954,N_14984);
or UO_212 (O_212,N_14956,N_14988);
or UO_213 (O_213,N_14976,N_14951);
nand UO_214 (O_214,N_14834,N_14802);
nand UO_215 (O_215,N_14975,N_14849);
and UO_216 (O_216,N_14970,N_14887);
nor UO_217 (O_217,N_14967,N_14841);
nand UO_218 (O_218,N_14885,N_14826);
xnor UO_219 (O_219,N_14988,N_14932);
nand UO_220 (O_220,N_14882,N_14857);
or UO_221 (O_221,N_14813,N_14913);
xor UO_222 (O_222,N_14816,N_14985);
or UO_223 (O_223,N_14981,N_14882);
or UO_224 (O_224,N_14906,N_14889);
nand UO_225 (O_225,N_14952,N_14933);
and UO_226 (O_226,N_14959,N_14846);
nor UO_227 (O_227,N_14966,N_14869);
xnor UO_228 (O_228,N_14845,N_14927);
nor UO_229 (O_229,N_14957,N_14859);
xor UO_230 (O_230,N_14979,N_14929);
xnor UO_231 (O_231,N_14998,N_14886);
xor UO_232 (O_232,N_14906,N_14935);
and UO_233 (O_233,N_14890,N_14851);
xnor UO_234 (O_234,N_14910,N_14832);
nor UO_235 (O_235,N_14970,N_14972);
xor UO_236 (O_236,N_14959,N_14811);
nand UO_237 (O_237,N_14800,N_14961);
and UO_238 (O_238,N_14805,N_14951);
or UO_239 (O_239,N_14865,N_14823);
nand UO_240 (O_240,N_14933,N_14876);
nand UO_241 (O_241,N_14944,N_14846);
or UO_242 (O_242,N_14985,N_14948);
nand UO_243 (O_243,N_14869,N_14989);
or UO_244 (O_244,N_14949,N_14918);
nand UO_245 (O_245,N_14879,N_14971);
xnor UO_246 (O_246,N_14908,N_14829);
and UO_247 (O_247,N_14877,N_14814);
and UO_248 (O_248,N_14926,N_14916);
nor UO_249 (O_249,N_14982,N_14804);
xor UO_250 (O_250,N_14812,N_14924);
and UO_251 (O_251,N_14988,N_14915);
or UO_252 (O_252,N_14911,N_14991);
nor UO_253 (O_253,N_14911,N_14981);
nand UO_254 (O_254,N_14910,N_14972);
and UO_255 (O_255,N_14905,N_14884);
nand UO_256 (O_256,N_14898,N_14975);
nor UO_257 (O_257,N_14837,N_14875);
or UO_258 (O_258,N_14819,N_14991);
nor UO_259 (O_259,N_14835,N_14917);
or UO_260 (O_260,N_14999,N_14808);
and UO_261 (O_261,N_14885,N_14950);
or UO_262 (O_262,N_14963,N_14809);
or UO_263 (O_263,N_14846,N_14869);
and UO_264 (O_264,N_14908,N_14835);
and UO_265 (O_265,N_14849,N_14918);
or UO_266 (O_266,N_14997,N_14981);
nor UO_267 (O_267,N_14909,N_14957);
and UO_268 (O_268,N_14866,N_14847);
xnor UO_269 (O_269,N_14923,N_14858);
xnor UO_270 (O_270,N_14958,N_14963);
or UO_271 (O_271,N_14841,N_14900);
or UO_272 (O_272,N_14898,N_14880);
and UO_273 (O_273,N_14868,N_14987);
or UO_274 (O_274,N_14846,N_14878);
nor UO_275 (O_275,N_14842,N_14966);
or UO_276 (O_276,N_14978,N_14972);
nand UO_277 (O_277,N_14820,N_14993);
xnor UO_278 (O_278,N_14826,N_14996);
nand UO_279 (O_279,N_14816,N_14874);
nor UO_280 (O_280,N_14983,N_14881);
xor UO_281 (O_281,N_14869,N_14967);
or UO_282 (O_282,N_14937,N_14882);
nand UO_283 (O_283,N_14989,N_14840);
xor UO_284 (O_284,N_14814,N_14846);
and UO_285 (O_285,N_14944,N_14911);
nand UO_286 (O_286,N_14952,N_14858);
nand UO_287 (O_287,N_14801,N_14974);
and UO_288 (O_288,N_14808,N_14804);
and UO_289 (O_289,N_14936,N_14949);
nor UO_290 (O_290,N_14909,N_14882);
xnor UO_291 (O_291,N_14921,N_14840);
and UO_292 (O_292,N_14934,N_14844);
nor UO_293 (O_293,N_14903,N_14877);
xor UO_294 (O_294,N_14825,N_14941);
nor UO_295 (O_295,N_14876,N_14994);
and UO_296 (O_296,N_14910,N_14928);
nor UO_297 (O_297,N_14946,N_14994);
and UO_298 (O_298,N_14827,N_14870);
nor UO_299 (O_299,N_14874,N_14837);
xnor UO_300 (O_300,N_14831,N_14805);
and UO_301 (O_301,N_14830,N_14902);
and UO_302 (O_302,N_14978,N_14990);
and UO_303 (O_303,N_14954,N_14929);
nor UO_304 (O_304,N_14925,N_14968);
and UO_305 (O_305,N_14927,N_14891);
nor UO_306 (O_306,N_14874,N_14805);
nor UO_307 (O_307,N_14884,N_14837);
or UO_308 (O_308,N_14916,N_14951);
or UO_309 (O_309,N_14974,N_14963);
or UO_310 (O_310,N_14850,N_14890);
or UO_311 (O_311,N_14943,N_14936);
nand UO_312 (O_312,N_14971,N_14841);
or UO_313 (O_313,N_14829,N_14893);
xnor UO_314 (O_314,N_14883,N_14998);
nor UO_315 (O_315,N_14845,N_14886);
or UO_316 (O_316,N_14955,N_14961);
xor UO_317 (O_317,N_14890,N_14844);
xnor UO_318 (O_318,N_14860,N_14944);
or UO_319 (O_319,N_14857,N_14996);
or UO_320 (O_320,N_14860,N_14817);
or UO_321 (O_321,N_14911,N_14889);
xnor UO_322 (O_322,N_14824,N_14882);
nor UO_323 (O_323,N_14962,N_14959);
xnor UO_324 (O_324,N_14942,N_14813);
or UO_325 (O_325,N_14953,N_14970);
nand UO_326 (O_326,N_14935,N_14999);
xor UO_327 (O_327,N_14825,N_14899);
or UO_328 (O_328,N_14955,N_14890);
and UO_329 (O_329,N_14851,N_14832);
and UO_330 (O_330,N_14931,N_14916);
and UO_331 (O_331,N_14882,N_14978);
and UO_332 (O_332,N_14988,N_14894);
or UO_333 (O_333,N_14999,N_14991);
xnor UO_334 (O_334,N_14939,N_14985);
xor UO_335 (O_335,N_14946,N_14893);
nor UO_336 (O_336,N_14811,N_14880);
nor UO_337 (O_337,N_14939,N_14910);
nor UO_338 (O_338,N_14891,N_14849);
and UO_339 (O_339,N_14801,N_14883);
nor UO_340 (O_340,N_14882,N_14862);
xor UO_341 (O_341,N_14817,N_14992);
and UO_342 (O_342,N_14927,N_14817);
xnor UO_343 (O_343,N_14940,N_14819);
nand UO_344 (O_344,N_14862,N_14820);
nand UO_345 (O_345,N_14832,N_14906);
xnor UO_346 (O_346,N_14842,N_14879);
nand UO_347 (O_347,N_14851,N_14920);
and UO_348 (O_348,N_14902,N_14836);
nand UO_349 (O_349,N_14960,N_14919);
nor UO_350 (O_350,N_14810,N_14948);
nand UO_351 (O_351,N_14931,N_14947);
and UO_352 (O_352,N_14942,N_14814);
nand UO_353 (O_353,N_14925,N_14982);
or UO_354 (O_354,N_14931,N_14849);
or UO_355 (O_355,N_14866,N_14950);
nor UO_356 (O_356,N_14815,N_14866);
or UO_357 (O_357,N_14989,N_14885);
or UO_358 (O_358,N_14964,N_14962);
nor UO_359 (O_359,N_14840,N_14987);
xor UO_360 (O_360,N_14991,N_14808);
and UO_361 (O_361,N_14934,N_14865);
nand UO_362 (O_362,N_14804,N_14955);
nor UO_363 (O_363,N_14994,N_14915);
and UO_364 (O_364,N_14822,N_14987);
xor UO_365 (O_365,N_14956,N_14938);
nand UO_366 (O_366,N_14920,N_14989);
or UO_367 (O_367,N_14850,N_14830);
xor UO_368 (O_368,N_14820,N_14965);
xor UO_369 (O_369,N_14994,N_14852);
xnor UO_370 (O_370,N_14810,N_14883);
nand UO_371 (O_371,N_14814,N_14856);
or UO_372 (O_372,N_14992,N_14898);
xnor UO_373 (O_373,N_14933,N_14845);
nor UO_374 (O_374,N_14944,N_14836);
nor UO_375 (O_375,N_14830,N_14832);
and UO_376 (O_376,N_14819,N_14880);
or UO_377 (O_377,N_14803,N_14990);
nor UO_378 (O_378,N_14942,N_14979);
or UO_379 (O_379,N_14835,N_14932);
or UO_380 (O_380,N_14835,N_14898);
nor UO_381 (O_381,N_14964,N_14802);
nor UO_382 (O_382,N_14856,N_14866);
nand UO_383 (O_383,N_14984,N_14982);
or UO_384 (O_384,N_14940,N_14833);
and UO_385 (O_385,N_14940,N_14817);
nor UO_386 (O_386,N_14832,N_14848);
nor UO_387 (O_387,N_14972,N_14849);
nor UO_388 (O_388,N_14881,N_14828);
xnor UO_389 (O_389,N_14807,N_14948);
xor UO_390 (O_390,N_14903,N_14933);
nor UO_391 (O_391,N_14832,N_14983);
nor UO_392 (O_392,N_14910,N_14982);
and UO_393 (O_393,N_14924,N_14889);
or UO_394 (O_394,N_14937,N_14959);
or UO_395 (O_395,N_14983,N_14984);
nor UO_396 (O_396,N_14802,N_14980);
nor UO_397 (O_397,N_14955,N_14958);
xnor UO_398 (O_398,N_14801,N_14954);
xnor UO_399 (O_399,N_14905,N_14928);
nor UO_400 (O_400,N_14821,N_14827);
nor UO_401 (O_401,N_14922,N_14974);
nand UO_402 (O_402,N_14834,N_14874);
and UO_403 (O_403,N_14975,N_14822);
or UO_404 (O_404,N_14962,N_14987);
nand UO_405 (O_405,N_14897,N_14813);
and UO_406 (O_406,N_14901,N_14808);
or UO_407 (O_407,N_14859,N_14898);
nor UO_408 (O_408,N_14962,N_14840);
xor UO_409 (O_409,N_14911,N_14968);
xnor UO_410 (O_410,N_14824,N_14857);
nor UO_411 (O_411,N_14851,N_14982);
nor UO_412 (O_412,N_14820,N_14897);
nand UO_413 (O_413,N_14938,N_14999);
and UO_414 (O_414,N_14875,N_14895);
or UO_415 (O_415,N_14965,N_14864);
or UO_416 (O_416,N_14931,N_14956);
nand UO_417 (O_417,N_14866,N_14963);
or UO_418 (O_418,N_14993,N_14832);
and UO_419 (O_419,N_14975,N_14832);
nand UO_420 (O_420,N_14956,N_14964);
nand UO_421 (O_421,N_14853,N_14830);
nor UO_422 (O_422,N_14875,N_14939);
xor UO_423 (O_423,N_14830,N_14880);
or UO_424 (O_424,N_14904,N_14885);
and UO_425 (O_425,N_14918,N_14914);
xnor UO_426 (O_426,N_14817,N_14914);
xor UO_427 (O_427,N_14818,N_14890);
and UO_428 (O_428,N_14885,N_14945);
xor UO_429 (O_429,N_14920,N_14965);
and UO_430 (O_430,N_14910,N_14868);
nand UO_431 (O_431,N_14992,N_14904);
nand UO_432 (O_432,N_14843,N_14950);
nand UO_433 (O_433,N_14853,N_14963);
or UO_434 (O_434,N_14867,N_14954);
nand UO_435 (O_435,N_14958,N_14816);
nor UO_436 (O_436,N_14908,N_14818);
or UO_437 (O_437,N_14812,N_14837);
nor UO_438 (O_438,N_14959,N_14816);
nand UO_439 (O_439,N_14941,N_14896);
xnor UO_440 (O_440,N_14924,N_14888);
nand UO_441 (O_441,N_14875,N_14955);
nand UO_442 (O_442,N_14921,N_14936);
or UO_443 (O_443,N_14965,N_14966);
nand UO_444 (O_444,N_14807,N_14815);
nand UO_445 (O_445,N_14872,N_14919);
nor UO_446 (O_446,N_14864,N_14800);
nor UO_447 (O_447,N_14830,N_14962);
and UO_448 (O_448,N_14872,N_14847);
nand UO_449 (O_449,N_14962,N_14904);
and UO_450 (O_450,N_14974,N_14825);
and UO_451 (O_451,N_14867,N_14893);
nor UO_452 (O_452,N_14877,N_14857);
or UO_453 (O_453,N_14887,N_14996);
nand UO_454 (O_454,N_14936,N_14934);
or UO_455 (O_455,N_14926,N_14900);
nand UO_456 (O_456,N_14968,N_14826);
nand UO_457 (O_457,N_14837,N_14900);
and UO_458 (O_458,N_14912,N_14849);
and UO_459 (O_459,N_14823,N_14872);
and UO_460 (O_460,N_14888,N_14926);
xnor UO_461 (O_461,N_14872,N_14962);
nand UO_462 (O_462,N_14989,N_14803);
or UO_463 (O_463,N_14808,N_14803);
or UO_464 (O_464,N_14820,N_14991);
or UO_465 (O_465,N_14811,N_14956);
and UO_466 (O_466,N_14863,N_14889);
nor UO_467 (O_467,N_14825,N_14912);
xnor UO_468 (O_468,N_14922,N_14838);
or UO_469 (O_469,N_14943,N_14949);
xnor UO_470 (O_470,N_14974,N_14951);
and UO_471 (O_471,N_14892,N_14821);
or UO_472 (O_472,N_14935,N_14937);
xor UO_473 (O_473,N_14827,N_14814);
or UO_474 (O_474,N_14881,N_14912);
nand UO_475 (O_475,N_14972,N_14857);
nor UO_476 (O_476,N_14823,N_14887);
xor UO_477 (O_477,N_14836,N_14813);
or UO_478 (O_478,N_14896,N_14830);
nor UO_479 (O_479,N_14849,N_14875);
xnor UO_480 (O_480,N_14970,N_14957);
nand UO_481 (O_481,N_14907,N_14925);
nor UO_482 (O_482,N_14951,N_14942);
or UO_483 (O_483,N_14830,N_14879);
xor UO_484 (O_484,N_14972,N_14899);
nor UO_485 (O_485,N_14998,N_14924);
xnor UO_486 (O_486,N_14995,N_14940);
and UO_487 (O_487,N_14945,N_14870);
or UO_488 (O_488,N_14879,N_14922);
xor UO_489 (O_489,N_14966,N_14825);
and UO_490 (O_490,N_14811,N_14878);
or UO_491 (O_491,N_14964,N_14951);
nor UO_492 (O_492,N_14924,N_14864);
nand UO_493 (O_493,N_14911,N_14925);
xnor UO_494 (O_494,N_14910,N_14967);
nor UO_495 (O_495,N_14937,N_14820);
or UO_496 (O_496,N_14926,N_14936);
or UO_497 (O_497,N_14828,N_14825);
and UO_498 (O_498,N_14985,N_14812);
and UO_499 (O_499,N_14928,N_14887);
xnor UO_500 (O_500,N_14866,N_14988);
and UO_501 (O_501,N_14879,N_14899);
xor UO_502 (O_502,N_14863,N_14941);
or UO_503 (O_503,N_14885,N_14955);
nor UO_504 (O_504,N_14951,N_14837);
xor UO_505 (O_505,N_14841,N_14808);
xnor UO_506 (O_506,N_14949,N_14981);
or UO_507 (O_507,N_14867,N_14945);
nor UO_508 (O_508,N_14946,N_14810);
and UO_509 (O_509,N_14885,N_14875);
xnor UO_510 (O_510,N_14998,N_14923);
nand UO_511 (O_511,N_14839,N_14917);
or UO_512 (O_512,N_14957,N_14968);
nor UO_513 (O_513,N_14894,N_14901);
or UO_514 (O_514,N_14881,N_14942);
and UO_515 (O_515,N_14983,N_14988);
nor UO_516 (O_516,N_14809,N_14925);
or UO_517 (O_517,N_14850,N_14917);
nand UO_518 (O_518,N_14985,N_14912);
or UO_519 (O_519,N_14822,N_14947);
xnor UO_520 (O_520,N_14981,N_14893);
or UO_521 (O_521,N_14877,N_14981);
nor UO_522 (O_522,N_14993,N_14894);
or UO_523 (O_523,N_14905,N_14850);
nor UO_524 (O_524,N_14853,N_14834);
nor UO_525 (O_525,N_14813,N_14984);
xor UO_526 (O_526,N_14833,N_14983);
or UO_527 (O_527,N_14870,N_14829);
nor UO_528 (O_528,N_14924,N_14863);
xor UO_529 (O_529,N_14927,N_14873);
nor UO_530 (O_530,N_14978,N_14876);
nor UO_531 (O_531,N_14947,N_14981);
and UO_532 (O_532,N_14932,N_14969);
and UO_533 (O_533,N_14885,N_14871);
or UO_534 (O_534,N_14978,N_14922);
or UO_535 (O_535,N_14981,N_14956);
xnor UO_536 (O_536,N_14987,N_14900);
nand UO_537 (O_537,N_14904,N_14833);
and UO_538 (O_538,N_14867,N_14896);
or UO_539 (O_539,N_14899,N_14989);
nand UO_540 (O_540,N_14894,N_14835);
and UO_541 (O_541,N_14808,N_14979);
or UO_542 (O_542,N_14916,N_14874);
and UO_543 (O_543,N_14956,N_14998);
nand UO_544 (O_544,N_14939,N_14996);
nand UO_545 (O_545,N_14926,N_14971);
xnor UO_546 (O_546,N_14810,N_14881);
or UO_547 (O_547,N_14963,N_14879);
xnor UO_548 (O_548,N_14966,N_14832);
nand UO_549 (O_549,N_14916,N_14882);
nand UO_550 (O_550,N_14946,N_14859);
or UO_551 (O_551,N_14993,N_14809);
nor UO_552 (O_552,N_14893,N_14887);
nor UO_553 (O_553,N_14909,N_14967);
nor UO_554 (O_554,N_14954,N_14999);
nor UO_555 (O_555,N_14993,N_14869);
and UO_556 (O_556,N_14850,N_14930);
and UO_557 (O_557,N_14931,N_14963);
or UO_558 (O_558,N_14888,N_14931);
xor UO_559 (O_559,N_14861,N_14837);
and UO_560 (O_560,N_14951,N_14920);
and UO_561 (O_561,N_14944,N_14831);
and UO_562 (O_562,N_14870,N_14832);
nand UO_563 (O_563,N_14887,N_14988);
nand UO_564 (O_564,N_14831,N_14887);
nor UO_565 (O_565,N_14856,N_14889);
xnor UO_566 (O_566,N_14976,N_14890);
nand UO_567 (O_567,N_14957,N_14926);
or UO_568 (O_568,N_14800,N_14951);
and UO_569 (O_569,N_14844,N_14975);
xnor UO_570 (O_570,N_14819,N_14826);
xnor UO_571 (O_571,N_14992,N_14808);
nor UO_572 (O_572,N_14803,N_14984);
nor UO_573 (O_573,N_14899,N_14918);
nor UO_574 (O_574,N_14855,N_14825);
xor UO_575 (O_575,N_14889,N_14965);
or UO_576 (O_576,N_14874,N_14872);
and UO_577 (O_577,N_14897,N_14803);
nor UO_578 (O_578,N_14982,N_14877);
nand UO_579 (O_579,N_14840,N_14980);
or UO_580 (O_580,N_14963,N_14959);
nand UO_581 (O_581,N_14986,N_14972);
nor UO_582 (O_582,N_14819,N_14839);
nand UO_583 (O_583,N_14821,N_14816);
nand UO_584 (O_584,N_14921,N_14993);
nand UO_585 (O_585,N_14920,N_14947);
or UO_586 (O_586,N_14854,N_14904);
or UO_587 (O_587,N_14856,N_14807);
nor UO_588 (O_588,N_14912,N_14940);
or UO_589 (O_589,N_14978,N_14833);
nand UO_590 (O_590,N_14959,N_14871);
nor UO_591 (O_591,N_14915,N_14995);
or UO_592 (O_592,N_14973,N_14881);
nand UO_593 (O_593,N_14992,N_14833);
xor UO_594 (O_594,N_14855,N_14944);
nand UO_595 (O_595,N_14910,N_14923);
and UO_596 (O_596,N_14890,N_14900);
xnor UO_597 (O_597,N_14881,N_14883);
and UO_598 (O_598,N_14883,N_14825);
and UO_599 (O_599,N_14868,N_14903);
or UO_600 (O_600,N_14909,N_14847);
nor UO_601 (O_601,N_14966,N_14810);
and UO_602 (O_602,N_14884,N_14812);
nand UO_603 (O_603,N_14895,N_14811);
xor UO_604 (O_604,N_14902,N_14870);
xnor UO_605 (O_605,N_14800,N_14844);
and UO_606 (O_606,N_14875,N_14821);
nand UO_607 (O_607,N_14919,N_14993);
xnor UO_608 (O_608,N_14950,N_14810);
xnor UO_609 (O_609,N_14949,N_14930);
or UO_610 (O_610,N_14864,N_14960);
or UO_611 (O_611,N_14928,N_14974);
nand UO_612 (O_612,N_14985,N_14863);
or UO_613 (O_613,N_14864,N_14941);
nand UO_614 (O_614,N_14959,N_14947);
and UO_615 (O_615,N_14842,N_14819);
nor UO_616 (O_616,N_14814,N_14874);
nor UO_617 (O_617,N_14934,N_14870);
or UO_618 (O_618,N_14898,N_14918);
nor UO_619 (O_619,N_14956,N_14879);
and UO_620 (O_620,N_14839,N_14825);
or UO_621 (O_621,N_14854,N_14818);
or UO_622 (O_622,N_14910,N_14988);
xnor UO_623 (O_623,N_14865,N_14915);
nand UO_624 (O_624,N_14878,N_14857);
and UO_625 (O_625,N_14826,N_14848);
or UO_626 (O_626,N_14804,N_14818);
nand UO_627 (O_627,N_14951,N_14838);
xnor UO_628 (O_628,N_14885,N_14833);
nor UO_629 (O_629,N_14855,N_14878);
and UO_630 (O_630,N_14819,N_14891);
nor UO_631 (O_631,N_14814,N_14994);
nor UO_632 (O_632,N_14871,N_14954);
and UO_633 (O_633,N_14929,N_14844);
nor UO_634 (O_634,N_14880,N_14981);
nor UO_635 (O_635,N_14850,N_14947);
and UO_636 (O_636,N_14811,N_14823);
nor UO_637 (O_637,N_14865,N_14859);
and UO_638 (O_638,N_14962,N_14907);
or UO_639 (O_639,N_14885,N_14944);
nor UO_640 (O_640,N_14854,N_14922);
nand UO_641 (O_641,N_14964,N_14941);
xor UO_642 (O_642,N_14833,N_14909);
or UO_643 (O_643,N_14810,N_14983);
nand UO_644 (O_644,N_14866,N_14928);
nor UO_645 (O_645,N_14814,N_14820);
nand UO_646 (O_646,N_14864,N_14972);
nor UO_647 (O_647,N_14951,N_14929);
nor UO_648 (O_648,N_14983,N_14805);
or UO_649 (O_649,N_14951,N_14967);
and UO_650 (O_650,N_14906,N_14895);
nor UO_651 (O_651,N_14977,N_14998);
and UO_652 (O_652,N_14948,N_14947);
xnor UO_653 (O_653,N_14822,N_14811);
xor UO_654 (O_654,N_14816,N_14892);
nor UO_655 (O_655,N_14816,N_14825);
nand UO_656 (O_656,N_14957,N_14975);
xnor UO_657 (O_657,N_14944,N_14983);
and UO_658 (O_658,N_14846,N_14907);
and UO_659 (O_659,N_14971,N_14935);
nor UO_660 (O_660,N_14988,N_14881);
or UO_661 (O_661,N_14888,N_14865);
or UO_662 (O_662,N_14840,N_14804);
nand UO_663 (O_663,N_14922,N_14835);
and UO_664 (O_664,N_14986,N_14824);
nand UO_665 (O_665,N_14806,N_14942);
or UO_666 (O_666,N_14874,N_14989);
xnor UO_667 (O_667,N_14881,N_14877);
xnor UO_668 (O_668,N_14917,N_14833);
nand UO_669 (O_669,N_14908,N_14995);
xor UO_670 (O_670,N_14903,N_14970);
nand UO_671 (O_671,N_14912,N_14976);
nand UO_672 (O_672,N_14951,N_14919);
nor UO_673 (O_673,N_14941,N_14976);
nor UO_674 (O_674,N_14864,N_14832);
nor UO_675 (O_675,N_14865,N_14849);
and UO_676 (O_676,N_14907,N_14802);
xor UO_677 (O_677,N_14981,N_14819);
and UO_678 (O_678,N_14969,N_14850);
or UO_679 (O_679,N_14818,N_14935);
nor UO_680 (O_680,N_14897,N_14889);
nor UO_681 (O_681,N_14950,N_14996);
nand UO_682 (O_682,N_14927,N_14812);
nor UO_683 (O_683,N_14932,N_14859);
or UO_684 (O_684,N_14931,N_14932);
nand UO_685 (O_685,N_14935,N_14800);
nor UO_686 (O_686,N_14975,N_14871);
and UO_687 (O_687,N_14907,N_14878);
or UO_688 (O_688,N_14805,N_14957);
or UO_689 (O_689,N_14891,N_14949);
or UO_690 (O_690,N_14955,N_14998);
xor UO_691 (O_691,N_14900,N_14980);
or UO_692 (O_692,N_14954,N_14823);
nand UO_693 (O_693,N_14940,N_14874);
or UO_694 (O_694,N_14832,N_14863);
or UO_695 (O_695,N_14807,N_14915);
or UO_696 (O_696,N_14899,N_14916);
or UO_697 (O_697,N_14867,N_14807);
nand UO_698 (O_698,N_14979,N_14840);
and UO_699 (O_699,N_14988,N_14908);
or UO_700 (O_700,N_14882,N_14970);
nand UO_701 (O_701,N_14871,N_14923);
and UO_702 (O_702,N_14913,N_14989);
nand UO_703 (O_703,N_14923,N_14837);
xnor UO_704 (O_704,N_14912,N_14858);
and UO_705 (O_705,N_14948,N_14997);
nor UO_706 (O_706,N_14939,N_14851);
nand UO_707 (O_707,N_14941,N_14872);
and UO_708 (O_708,N_14829,N_14923);
nor UO_709 (O_709,N_14993,N_14911);
and UO_710 (O_710,N_14803,N_14960);
xor UO_711 (O_711,N_14920,N_14827);
nand UO_712 (O_712,N_14922,N_14958);
nor UO_713 (O_713,N_14925,N_14871);
nand UO_714 (O_714,N_14846,N_14996);
nor UO_715 (O_715,N_14938,N_14877);
or UO_716 (O_716,N_14902,N_14954);
nor UO_717 (O_717,N_14814,N_14963);
xor UO_718 (O_718,N_14949,N_14928);
nand UO_719 (O_719,N_14809,N_14845);
nand UO_720 (O_720,N_14893,N_14875);
nor UO_721 (O_721,N_14866,N_14910);
nand UO_722 (O_722,N_14912,N_14930);
nor UO_723 (O_723,N_14975,N_14839);
xnor UO_724 (O_724,N_14828,N_14887);
xor UO_725 (O_725,N_14994,N_14976);
and UO_726 (O_726,N_14978,N_14924);
and UO_727 (O_727,N_14940,N_14866);
xor UO_728 (O_728,N_14883,N_14985);
nand UO_729 (O_729,N_14835,N_14962);
or UO_730 (O_730,N_14825,N_14981);
nand UO_731 (O_731,N_14832,N_14967);
or UO_732 (O_732,N_14829,N_14924);
or UO_733 (O_733,N_14844,N_14991);
nor UO_734 (O_734,N_14931,N_14867);
xor UO_735 (O_735,N_14906,N_14914);
and UO_736 (O_736,N_14898,N_14858);
xor UO_737 (O_737,N_14902,N_14908);
nor UO_738 (O_738,N_14877,N_14905);
nor UO_739 (O_739,N_14862,N_14815);
and UO_740 (O_740,N_14817,N_14966);
nor UO_741 (O_741,N_14889,N_14834);
and UO_742 (O_742,N_14817,N_14815);
nor UO_743 (O_743,N_14955,N_14876);
and UO_744 (O_744,N_14841,N_14806);
nor UO_745 (O_745,N_14950,N_14888);
nor UO_746 (O_746,N_14946,N_14833);
and UO_747 (O_747,N_14842,N_14828);
xor UO_748 (O_748,N_14906,N_14992);
nor UO_749 (O_749,N_14839,N_14978);
or UO_750 (O_750,N_14967,N_14954);
and UO_751 (O_751,N_14927,N_14967);
and UO_752 (O_752,N_14884,N_14861);
and UO_753 (O_753,N_14856,N_14863);
xor UO_754 (O_754,N_14990,N_14845);
or UO_755 (O_755,N_14964,N_14918);
nand UO_756 (O_756,N_14866,N_14832);
or UO_757 (O_757,N_14924,N_14910);
nand UO_758 (O_758,N_14855,N_14949);
and UO_759 (O_759,N_14813,N_14987);
or UO_760 (O_760,N_14992,N_14801);
or UO_761 (O_761,N_14869,N_14863);
or UO_762 (O_762,N_14878,N_14824);
nor UO_763 (O_763,N_14958,N_14835);
nand UO_764 (O_764,N_14907,N_14863);
xnor UO_765 (O_765,N_14892,N_14805);
or UO_766 (O_766,N_14809,N_14944);
or UO_767 (O_767,N_14989,N_14875);
and UO_768 (O_768,N_14883,N_14848);
xnor UO_769 (O_769,N_14862,N_14927);
or UO_770 (O_770,N_14844,N_14928);
or UO_771 (O_771,N_14996,N_14931);
and UO_772 (O_772,N_14873,N_14814);
nor UO_773 (O_773,N_14910,N_14968);
nor UO_774 (O_774,N_14820,N_14835);
nor UO_775 (O_775,N_14851,N_14946);
nand UO_776 (O_776,N_14824,N_14834);
and UO_777 (O_777,N_14936,N_14837);
nor UO_778 (O_778,N_14959,N_14902);
nand UO_779 (O_779,N_14854,N_14861);
xor UO_780 (O_780,N_14998,N_14896);
nand UO_781 (O_781,N_14876,N_14948);
nand UO_782 (O_782,N_14973,N_14809);
nor UO_783 (O_783,N_14867,N_14847);
or UO_784 (O_784,N_14848,N_14814);
or UO_785 (O_785,N_14899,N_14941);
or UO_786 (O_786,N_14951,N_14935);
xor UO_787 (O_787,N_14889,N_14846);
nand UO_788 (O_788,N_14806,N_14881);
nand UO_789 (O_789,N_14963,N_14831);
xnor UO_790 (O_790,N_14957,N_14815);
nand UO_791 (O_791,N_14980,N_14901);
xor UO_792 (O_792,N_14911,N_14964);
xor UO_793 (O_793,N_14949,N_14998);
xnor UO_794 (O_794,N_14800,N_14922);
xnor UO_795 (O_795,N_14897,N_14933);
xor UO_796 (O_796,N_14989,N_14957);
xnor UO_797 (O_797,N_14991,N_14952);
xnor UO_798 (O_798,N_14877,N_14910);
or UO_799 (O_799,N_14912,N_14824);
nor UO_800 (O_800,N_14885,N_14819);
nor UO_801 (O_801,N_14935,N_14911);
nand UO_802 (O_802,N_14938,N_14842);
or UO_803 (O_803,N_14914,N_14984);
nor UO_804 (O_804,N_14950,N_14977);
and UO_805 (O_805,N_14986,N_14997);
nand UO_806 (O_806,N_14892,N_14861);
nor UO_807 (O_807,N_14983,N_14886);
xnor UO_808 (O_808,N_14865,N_14837);
nor UO_809 (O_809,N_14972,N_14839);
xnor UO_810 (O_810,N_14877,N_14813);
nand UO_811 (O_811,N_14999,N_14812);
xnor UO_812 (O_812,N_14988,N_14843);
nand UO_813 (O_813,N_14915,N_14831);
or UO_814 (O_814,N_14964,N_14884);
nand UO_815 (O_815,N_14972,N_14841);
xor UO_816 (O_816,N_14884,N_14865);
and UO_817 (O_817,N_14925,N_14916);
xor UO_818 (O_818,N_14902,N_14868);
and UO_819 (O_819,N_14940,N_14862);
nand UO_820 (O_820,N_14897,N_14884);
or UO_821 (O_821,N_14960,N_14970);
or UO_822 (O_822,N_14888,N_14857);
or UO_823 (O_823,N_14874,N_14906);
and UO_824 (O_824,N_14800,N_14858);
nor UO_825 (O_825,N_14976,N_14834);
and UO_826 (O_826,N_14997,N_14867);
or UO_827 (O_827,N_14883,N_14905);
or UO_828 (O_828,N_14865,N_14913);
or UO_829 (O_829,N_14964,N_14869);
nor UO_830 (O_830,N_14902,N_14827);
or UO_831 (O_831,N_14824,N_14800);
nor UO_832 (O_832,N_14911,N_14955);
or UO_833 (O_833,N_14985,N_14974);
nor UO_834 (O_834,N_14962,N_14989);
nand UO_835 (O_835,N_14846,N_14934);
nor UO_836 (O_836,N_14811,N_14916);
or UO_837 (O_837,N_14897,N_14919);
nand UO_838 (O_838,N_14926,N_14845);
nand UO_839 (O_839,N_14842,N_14856);
xnor UO_840 (O_840,N_14837,N_14827);
or UO_841 (O_841,N_14880,N_14968);
xor UO_842 (O_842,N_14998,N_14803);
xnor UO_843 (O_843,N_14987,N_14932);
xnor UO_844 (O_844,N_14901,N_14973);
nand UO_845 (O_845,N_14872,N_14846);
and UO_846 (O_846,N_14848,N_14935);
and UO_847 (O_847,N_14954,N_14915);
nand UO_848 (O_848,N_14967,N_14813);
nor UO_849 (O_849,N_14857,N_14969);
and UO_850 (O_850,N_14884,N_14830);
nor UO_851 (O_851,N_14905,N_14866);
and UO_852 (O_852,N_14914,N_14924);
nor UO_853 (O_853,N_14879,N_14900);
xnor UO_854 (O_854,N_14947,N_14812);
or UO_855 (O_855,N_14927,N_14913);
nor UO_856 (O_856,N_14903,N_14966);
nand UO_857 (O_857,N_14851,N_14863);
and UO_858 (O_858,N_14922,N_14818);
nor UO_859 (O_859,N_14932,N_14967);
nor UO_860 (O_860,N_14850,N_14892);
xor UO_861 (O_861,N_14869,N_14909);
and UO_862 (O_862,N_14838,N_14945);
and UO_863 (O_863,N_14937,N_14808);
nand UO_864 (O_864,N_14885,N_14952);
xnor UO_865 (O_865,N_14816,N_14814);
xnor UO_866 (O_866,N_14875,N_14965);
nor UO_867 (O_867,N_14895,N_14911);
nor UO_868 (O_868,N_14865,N_14814);
xor UO_869 (O_869,N_14841,N_14852);
and UO_870 (O_870,N_14926,N_14933);
and UO_871 (O_871,N_14990,N_14808);
or UO_872 (O_872,N_14935,N_14905);
or UO_873 (O_873,N_14987,N_14870);
nand UO_874 (O_874,N_14948,N_14863);
xnor UO_875 (O_875,N_14807,N_14885);
nor UO_876 (O_876,N_14802,N_14876);
nand UO_877 (O_877,N_14886,N_14921);
or UO_878 (O_878,N_14859,N_14930);
or UO_879 (O_879,N_14875,N_14807);
and UO_880 (O_880,N_14946,N_14857);
and UO_881 (O_881,N_14835,N_14956);
xor UO_882 (O_882,N_14817,N_14858);
nand UO_883 (O_883,N_14911,N_14997);
xnor UO_884 (O_884,N_14882,N_14896);
or UO_885 (O_885,N_14902,N_14942);
nand UO_886 (O_886,N_14925,N_14805);
xnor UO_887 (O_887,N_14933,N_14858);
and UO_888 (O_888,N_14850,N_14954);
and UO_889 (O_889,N_14938,N_14887);
and UO_890 (O_890,N_14977,N_14988);
or UO_891 (O_891,N_14909,N_14948);
nor UO_892 (O_892,N_14839,N_14824);
xor UO_893 (O_893,N_14944,N_14841);
nor UO_894 (O_894,N_14850,N_14813);
xor UO_895 (O_895,N_14869,N_14990);
nand UO_896 (O_896,N_14915,N_14860);
nor UO_897 (O_897,N_14985,N_14986);
or UO_898 (O_898,N_14984,N_14900);
and UO_899 (O_899,N_14833,N_14824);
nand UO_900 (O_900,N_14970,N_14841);
xnor UO_901 (O_901,N_14985,N_14966);
xnor UO_902 (O_902,N_14831,N_14969);
or UO_903 (O_903,N_14860,N_14971);
nand UO_904 (O_904,N_14945,N_14965);
nand UO_905 (O_905,N_14926,N_14896);
and UO_906 (O_906,N_14973,N_14999);
and UO_907 (O_907,N_14880,N_14877);
nor UO_908 (O_908,N_14807,N_14967);
xnor UO_909 (O_909,N_14950,N_14853);
xor UO_910 (O_910,N_14884,N_14958);
nand UO_911 (O_911,N_14991,N_14841);
or UO_912 (O_912,N_14891,N_14853);
nand UO_913 (O_913,N_14877,N_14988);
xor UO_914 (O_914,N_14935,N_14900);
xor UO_915 (O_915,N_14821,N_14950);
or UO_916 (O_916,N_14840,N_14958);
nand UO_917 (O_917,N_14816,N_14946);
xnor UO_918 (O_918,N_14922,N_14827);
nor UO_919 (O_919,N_14964,N_14886);
nand UO_920 (O_920,N_14933,N_14916);
and UO_921 (O_921,N_14809,N_14847);
nor UO_922 (O_922,N_14966,N_14883);
or UO_923 (O_923,N_14931,N_14909);
nand UO_924 (O_924,N_14824,N_14859);
nand UO_925 (O_925,N_14871,N_14827);
nand UO_926 (O_926,N_14886,N_14999);
or UO_927 (O_927,N_14866,N_14874);
nor UO_928 (O_928,N_14908,N_14909);
nor UO_929 (O_929,N_14816,N_14921);
and UO_930 (O_930,N_14866,N_14872);
nor UO_931 (O_931,N_14962,N_14917);
nand UO_932 (O_932,N_14962,N_14870);
nor UO_933 (O_933,N_14811,N_14955);
nand UO_934 (O_934,N_14831,N_14940);
and UO_935 (O_935,N_14975,N_14886);
xor UO_936 (O_936,N_14989,N_14915);
and UO_937 (O_937,N_14855,N_14954);
or UO_938 (O_938,N_14984,N_14919);
nor UO_939 (O_939,N_14904,N_14938);
nor UO_940 (O_940,N_14854,N_14862);
or UO_941 (O_941,N_14899,N_14960);
nor UO_942 (O_942,N_14952,N_14887);
xnor UO_943 (O_943,N_14984,N_14807);
nand UO_944 (O_944,N_14972,N_14903);
xnor UO_945 (O_945,N_14805,N_14961);
and UO_946 (O_946,N_14874,N_14994);
nand UO_947 (O_947,N_14870,N_14975);
or UO_948 (O_948,N_14905,N_14901);
nor UO_949 (O_949,N_14842,N_14846);
and UO_950 (O_950,N_14841,N_14803);
nand UO_951 (O_951,N_14805,N_14924);
nand UO_952 (O_952,N_14990,N_14887);
nor UO_953 (O_953,N_14969,N_14864);
or UO_954 (O_954,N_14922,N_14892);
nor UO_955 (O_955,N_14865,N_14815);
nand UO_956 (O_956,N_14834,N_14951);
xnor UO_957 (O_957,N_14963,N_14957);
and UO_958 (O_958,N_14975,N_14921);
and UO_959 (O_959,N_14935,N_14806);
and UO_960 (O_960,N_14840,N_14828);
xor UO_961 (O_961,N_14922,N_14820);
xnor UO_962 (O_962,N_14989,N_14993);
or UO_963 (O_963,N_14886,N_14894);
nor UO_964 (O_964,N_14958,N_14925);
or UO_965 (O_965,N_14935,N_14919);
xnor UO_966 (O_966,N_14927,N_14838);
and UO_967 (O_967,N_14832,N_14815);
or UO_968 (O_968,N_14987,N_14845);
and UO_969 (O_969,N_14863,N_14972);
and UO_970 (O_970,N_14950,N_14931);
or UO_971 (O_971,N_14893,N_14965);
and UO_972 (O_972,N_14859,N_14881);
xnor UO_973 (O_973,N_14925,N_14955);
and UO_974 (O_974,N_14944,N_14955);
or UO_975 (O_975,N_14911,N_14967);
nor UO_976 (O_976,N_14884,N_14921);
xnor UO_977 (O_977,N_14994,N_14866);
nor UO_978 (O_978,N_14853,N_14805);
nor UO_979 (O_979,N_14947,N_14877);
and UO_980 (O_980,N_14891,N_14823);
nor UO_981 (O_981,N_14890,N_14918);
xor UO_982 (O_982,N_14995,N_14936);
nor UO_983 (O_983,N_14874,N_14980);
xnor UO_984 (O_984,N_14925,N_14824);
nor UO_985 (O_985,N_14929,N_14804);
nor UO_986 (O_986,N_14975,N_14964);
and UO_987 (O_987,N_14972,N_14871);
and UO_988 (O_988,N_14903,N_14811);
or UO_989 (O_989,N_14889,N_14812);
nand UO_990 (O_990,N_14971,N_14869);
nor UO_991 (O_991,N_14861,N_14908);
or UO_992 (O_992,N_14906,N_14879);
nor UO_993 (O_993,N_14878,N_14885);
nand UO_994 (O_994,N_14952,N_14920);
and UO_995 (O_995,N_14913,N_14897);
or UO_996 (O_996,N_14910,N_14911);
nor UO_997 (O_997,N_14978,N_14932);
and UO_998 (O_998,N_14956,N_14892);
nand UO_999 (O_999,N_14857,N_14805);
nor UO_1000 (O_1000,N_14839,N_14887);
and UO_1001 (O_1001,N_14814,N_14941);
and UO_1002 (O_1002,N_14820,N_14908);
xnor UO_1003 (O_1003,N_14993,N_14981);
and UO_1004 (O_1004,N_14832,N_14985);
nor UO_1005 (O_1005,N_14861,N_14975);
nor UO_1006 (O_1006,N_14944,N_14906);
nand UO_1007 (O_1007,N_14855,N_14950);
or UO_1008 (O_1008,N_14864,N_14978);
xnor UO_1009 (O_1009,N_14817,N_14906);
nor UO_1010 (O_1010,N_14862,N_14962);
nor UO_1011 (O_1011,N_14847,N_14994);
nand UO_1012 (O_1012,N_14945,N_14964);
nor UO_1013 (O_1013,N_14824,N_14990);
nand UO_1014 (O_1014,N_14940,N_14821);
and UO_1015 (O_1015,N_14878,N_14875);
and UO_1016 (O_1016,N_14922,N_14914);
nor UO_1017 (O_1017,N_14951,N_14841);
nand UO_1018 (O_1018,N_14985,N_14993);
or UO_1019 (O_1019,N_14980,N_14916);
xnor UO_1020 (O_1020,N_14957,N_14802);
or UO_1021 (O_1021,N_14873,N_14939);
nor UO_1022 (O_1022,N_14972,N_14925);
nand UO_1023 (O_1023,N_14827,N_14982);
nor UO_1024 (O_1024,N_14803,N_14923);
or UO_1025 (O_1025,N_14929,N_14969);
or UO_1026 (O_1026,N_14878,N_14828);
nor UO_1027 (O_1027,N_14935,N_14825);
nor UO_1028 (O_1028,N_14847,N_14820);
or UO_1029 (O_1029,N_14858,N_14892);
or UO_1030 (O_1030,N_14805,N_14803);
and UO_1031 (O_1031,N_14804,N_14859);
or UO_1032 (O_1032,N_14975,N_14937);
nand UO_1033 (O_1033,N_14810,N_14864);
nand UO_1034 (O_1034,N_14880,N_14982);
and UO_1035 (O_1035,N_14936,N_14972);
nand UO_1036 (O_1036,N_14901,N_14955);
and UO_1037 (O_1037,N_14957,N_14910);
nand UO_1038 (O_1038,N_14866,N_14882);
xor UO_1039 (O_1039,N_14935,N_14932);
nand UO_1040 (O_1040,N_14854,N_14863);
nand UO_1041 (O_1041,N_14934,N_14985);
nor UO_1042 (O_1042,N_14877,N_14873);
or UO_1043 (O_1043,N_14853,N_14864);
nor UO_1044 (O_1044,N_14969,N_14941);
or UO_1045 (O_1045,N_14973,N_14847);
nand UO_1046 (O_1046,N_14880,N_14936);
or UO_1047 (O_1047,N_14903,N_14936);
nand UO_1048 (O_1048,N_14991,N_14961);
xnor UO_1049 (O_1049,N_14985,N_14867);
nor UO_1050 (O_1050,N_14858,N_14874);
nor UO_1051 (O_1051,N_14846,N_14977);
or UO_1052 (O_1052,N_14829,N_14890);
and UO_1053 (O_1053,N_14937,N_14813);
nand UO_1054 (O_1054,N_14836,N_14828);
xnor UO_1055 (O_1055,N_14800,N_14808);
nor UO_1056 (O_1056,N_14957,N_14940);
or UO_1057 (O_1057,N_14963,N_14923);
xor UO_1058 (O_1058,N_14853,N_14803);
xor UO_1059 (O_1059,N_14995,N_14879);
nor UO_1060 (O_1060,N_14854,N_14826);
or UO_1061 (O_1061,N_14909,N_14906);
nand UO_1062 (O_1062,N_14932,N_14899);
or UO_1063 (O_1063,N_14944,N_14941);
xnor UO_1064 (O_1064,N_14895,N_14898);
nor UO_1065 (O_1065,N_14947,N_14833);
nand UO_1066 (O_1066,N_14957,N_14948);
and UO_1067 (O_1067,N_14904,N_14879);
xnor UO_1068 (O_1068,N_14940,N_14992);
and UO_1069 (O_1069,N_14988,N_14882);
nand UO_1070 (O_1070,N_14889,N_14841);
or UO_1071 (O_1071,N_14862,N_14924);
and UO_1072 (O_1072,N_14805,N_14902);
or UO_1073 (O_1073,N_14828,N_14931);
nor UO_1074 (O_1074,N_14968,N_14898);
or UO_1075 (O_1075,N_14834,N_14852);
xor UO_1076 (O_1076,N_14843,N_14926);
xor UO_1077 (O_1077,N_14869,N_14926);
and UO_1078 (O_1078,N_14961,N_14973);
or UO_1079 (O_1079,N_14815,N_14997);
nor UO_1080 (O_1080,N_14843,N_14857);
and UO_1081 (O_1081,N_14877,N_14902);
or UO_1082 (O_1082,N_14889,N_14817);
nor UO_1083 (O_1083,N_14889,N_14842);
nand UO_1084 (O_1084,N_14831,N_14985);
nor UO_1085 (O_1085,N_14827,N_14851);
or UO_1086 (O_1086,N_14937,N_14913);
nor UO_1087 (O_1087,N_14842,N_14987);
nand UO_1088 (O_1088,N_14927,N_14894);
and UO_1089 (O_1089,N_14882,N_14844);
nor UO_1090 (O_1090,N_14807,N_14925);
xor UO_1091 (O_1091,N_14903,N_14844);
xor UO_1092 (O_1092,N_14809,N_14976);
or UO_1093 (O_1093,N_14836,N_14906);
nand UO_1094 (O_1094,N_14995,N_14949);
nor UO_1095 (O_1095,N_14802,N_14868);
or UO_1096 (O_1096,N_14854,N_14919);
nor UO_1097 (O_1097,N_14922,N_14815);
nor UO_1098 (O_1098,N_14905,N_14985);
and UO_1099 (O_1099,N_14872,N_14992);
and UO_1100 (O_1100,N_14825,N_14827);
nor UO_1101 (O_1101,N_14996,N_14890);
nand UO_1102 (O_1102,N_14872,N_14973);
nand UO_1103 (O_1103,N_14860,N_14919);
and UO_1104 (O_1104,N_14916,N_14922);
nor UO_1105 (O_1105,N_14904,N_14967);
nand UO_1106 (O_1106,N_14996,N_14952);
xor UO_1107 (O_1107,N_14889,N_14921);
or UO_1108 (O_1108,N_14823,N_14844);
or UO_1109 (O_1109,N_14813,N_14856);
or UO_1110 (O_1110,N_14956,N_14838);
nor UO_1111 (O_1111,N_14848,N_14964);
and UO_1112 (O_1112,N_14866,N_14889);
nor UO_1113 (O_1113,N_14856,N_14960);
nor UO_1114 (O_1114,N_14878,N_14939);
nand UO_1115 (O_1115,N_14950,N_14944);
nand UO_1116 (O_1116,N_14908,N_14920);
nand UO_1117 (O_1117,N_14997,N_14960);
nand UO_1118 (O_1118,N_14841,N_14945);
or UO_1119 (O_1119,N_14828,N_14877);
xor UO_1120 (O_1120,N_14991,N_14907);
or UO_1121 (O_1121,N_14883,N_14809);
xnor UO_1122 (O_1122,N_14825,N_14859);
or UO_1123 (O_1123,N_14998,N_14903);
nor UO_1124 (O_1124,N_14871,N_14988);
or UO_1125 (O_1125,N_14810,N_14828);
and UO_1126 (O_1126,N_14863,N_14955);
nor UO_1127 (O_1127,N_14910,N_14825);
nor UO_1128 (O_1128,N_14913,N_14908);
xor UO_1129 (O_1129,N_14811,N_14904);
and UO_1130 (O_1130,N_14946,N_14973);
or UO_1131 (O_1131,N_14963,N_14863);
xnor UO_1132 (O_1132,N_14829,N_14997);
and UO_1133 (O_1133,N_14902,N_14973);
or UO_1134 (O_1134,N_14984,N_14800);
or UO_1135 (O_1135,N_14839,N_14880);
nor UO_1136 (O_1136,N_14915,N_14856);
or UO_1137 (O_1137,N_14940,N_14934);
xnor UO_1138 (O_1138,N_14936,N_14916);
and UO_1139 (O_1139,N_14975,N_14923);
xnor UO_1140 (O_1140,N_14954,N_14800);
nor UO_1141 (O_1141,N_14972,N_14853);
xnor UO_1142 (O_1142,N_14908,N_14839);
or UO_1143 (O_1143,N_14897,N_14822);
or UO_1144 (O_1144,N_14937,N_14963);
xnor UO_1145 (O_1145,N_14831,N_14979);
or UO_1146 (O_1146,N_14883,N_14815);
xor UO_1147 (O_1147,N_14800,N_14801);
or UO_1148 (O_1148,N_14853,N_14971);
nor UO_1149 (O_1149,N_14868,N_14919);
and UO_1150 (O_1150,N_14863,N_14841);
nand UO_1151 (O_1151,N_14864,N_14909);
nand UO_1152 (O_1152,N_14817,N_14874);
nor UO_1153 (O_1153,N_14991,N_14840);
and UO_1154 (O_1154,N_14988,N_14999);
or UO_1155 (O_1155,N_14909,N_14995);
and UO_1156 (O_1156,N_14854,N_14868);
nand UO_1157 (O_1157,N_14975,N_14905);
nor UO_1158 (O_1158,N_14890,N_14919);
nand UO_1159 (O_1159,N_14914,N_14844);
or UO_1160 (O_1160,N_14871,N_14807);
nand UO_1161 (O_1161,N_14862,N_14971);
xnor UO_1162 (O_1162,N_14964,N_14976);
and UO_1163 (O_1163,N_14814,N_14976);
and UO_1164 (O_1164,N_14862,N_14872);
and UO_1165 (O_1165,N_14886,N_14882);
nand UO_1166 (O_1166,N_14972,N_14941);
and UO_1167 (O_1167,N_14956,N_14919);
and UO_1168 (O_1168,N_14965,N_14881);
nand UO_1169 (O_1169,N_14829,N_14832);
and UO_1170 (O_1170,N_14902,N_14897);
xor UO_1171 (O_1171,N_14978,N_14835);
xnor UO_1172 (O_1172,N_14921,N_14974);
and UO_1173 (O_1173,N_14989,N_14948);
nand UO_1174 (O_1174,N_14895,N_14809);
nand UO_1175 (O_1175,N_14950,N_14947);
nand UO_1176 (O_1176,N_14826,N_14800);
nor UO_1177 (O_1177,N_14944,N_14894);
and UO_1178 (O_1178,N_14901,N_14824);
and UO_1179 (O_1179,N_14925,N_14847);
or UO_1180 (O_1180,N_14927,N_14866);
xor UO_1181 (O_1181,N_14900,N_14916);
nand UO_1182 (O_1182,N_14838,N_14852);
xnor UO_1183 (O_1183,N_14994,N_14911);
or UO_1184 (O_1184,N_14874,N_14892);
nor UO_1185 (O_1185,N_14850,N_14868);
nor UO_1186 (O_1186,N_14875,N_14975);
nor UO_1187 (O_1187,N_14833,N_14891);
xor UO_1188 (O_1188,N_14882,N_14950);
nand UO_1189 (O_1189,N_14914,N_14841);
nand UO_1190 (O_1190,N_14926,N_14890);
nor UO_1191 (O_1191,N_14888,N_14906);
or UO_1192 (O_1192,N_14954,N_14919);
or UO_1193 (O_1193,N_14841,N_14802);
nor UO_1194 (O_1194,N_14861,N_14863);
xor UO_1195 (O_1195,N_14884,N_14889);
nor UO_1196 (O_1196,N_14874,N_14918);
or UO_1197 (O_1197,N_14933,N_14842);
nor UO_1198 (O_1198,N_14989,N_14800);
or UO_1199 (O_1199,N_14993,N_14847);
nor UO_1200 (O_1200,N_14913,N_14847);
and UO_1201 (O_1201,N_14917,N_14957);
or UO_1202 (O_1202,N_14945,N_14832);
and UO_1203 (O_1203,N_14983,N_14934);
or UO_1204 (O_1204,N_14831,N_14950);
and UO_1205 (O_1205,N_14855,N_14806);
nand UO_1206 (O_1206,N_14803,N_14899);
xor UO_1207 (O_1207,N_14890,N_14812);
nor UO_1208 (O_1208,N_14860,N_14856);
and UO_1209 (O_1209,N_14827,N_14810);
xor UO_1210 (O_1210,N_14921,N_14971);
nor UO_1211 (O_1211,N_14855,N_14890);
xor UO_1212 (O_1212,N_14963,N_14952);
and UO_1213 (O_1213,N_14853,N_14906);
or UO_1214 (O_1214,N_14846,N_14816);
and UO_1215 (O_1215,N_14811,N_14973);
or UO_1216 (O_1216,N_14822,N_14803);
xnor UO_1217 (O_1217,N_14883,N_14962);
and UO_1218 (O_1218,N_14931,N_14874);
and UO_1219 (O_1219,N_14818,N_14812);
nand UO_1220 (O_1220,N_14892,N_14919);
and UO_1221 (O_1221,N_14861,N_14852);
nor UO_1222 (O_1222,N_14831,N_14902);
or UO_1223 (O_1223,N_14874,N_14869);
nand UO_1224 (O_1224,N_14989,N_14852);
nand UO_1225 (O_1225,N_14936,N_14985);
or UO_1226 (O_1226,N_14962,N_14857);
nor UO_1227 (O_1227,N_14820,N_14915);
nor UO_1228 (O_1228,N_14950,N_14849);
and UO_1229 (O_1229,N_14892,N_14934);
and UO_1230 (O_1230,N_14886,N_14895);
or UO_1231 (O_1231,N_14897,N_14866);
xor UO_1232 (O_1232,N_14950,N_14908);
nand UO_1233 (O_1233,N_14937,N_14968);
nor UO_1234 (O_1234,N_14905,N_14922);
nand UO_1235 (O_1235,N_14926,N_14903);
nand UO_1236 (O_1236,N_14875,N_14869);
nand UO_1237 (O_1237,N_14894,N_14924);
and UO_1238 (O_1238,N_14895,N_14851);
xnor UO_1239 (O_1239,N_14925,N_14977);
or UO_1240 (O_1240,N_14946,N_14814);
nand UO_1241 (O_1241,N_14804,N_14952);
or UO_1242 (O_1242,N_14953,N_14928);
and UO_1243 (O_1243,N_14846,N_14884);
or UO_1244 (O_1244,N_14947,N_14938);
nand UO_1245 (O_1245,N_14971,N_14896);
or UO_1246 (O_1246,N_14977,N_14820);
or UO_1247 (O_1247,N_14842,N_14984);
or UO_1248 (O_1248,N_14978,N_14842);
and UO_1249 (O_1249,N_14881,N_14870);
nand UO_1250 (O_1250,N_14972,N_14833);
nand UO_1251 (O_1251,N_14948,N_14852);
or UO_1252 (O_1252,N_14954,N_14805);
and UO_1253 (O_1253,N_14938,N_14965);
nand UO_1254 (O_1254,N_14892,N_14962);
or UO_1255 (O_1255,N_14808,N_14964);
or UO_1256 (O_1256,N_14967,N_14899);
or UO_1257 (O_1257,N_14989,N_14834);
or UO_1258 (O_1258,N_14864,N_14805);
xor UO_1259 (O_1259,N_14966,N_14976);
nand UO_1260 (O_1260,N_14885,N_14931);
and UO_1261 (O_1261,N_14926,N_14997);
or UO_1262 (O_1262,N_14855,N_14852);
nor UO_1263 (O_1263,N_14986,N_14887);
nand UO_1264 (O_1264,N_14828,N_14870);
xnor UO_1265 (O_1265,N_14985,N_14914);
and UO_1266 (O_1266,N_14991,N_14923);
and UO_1267 (O_1267,N_14874,N_14833);
and UO_1268 (O_1268,N_14827,N_14959);
or UO_1269 (O_1269,N_14887,N_14898);
and UO_1270 (O_1270,N_14841,N_14977);
nand UO_1271 (O_1271,N_14888,N_14873);
nor UO_1272 (O_1272,N_14951,N_14952);
xor UO_1273 (O_1273,N_14982,N_14841);
nor UO_1274 (O_1274,N_14961,N_14809);
nor UO_1275 (O_1275,N_14829,N_14949);
and UO_1276 (O_1276,N_14852,N_14895);
or UO_1277 (O_1277,N_14867,N_14972);
and UO_1278 (O_1278,N_14926,N_14830);
and UO_1279 (O_1279,N_14814,N_14978);
or UO_1280 (O_1280,N_14871,N_14946);
nor UO_1281 (O_1281,N_14857,N_14875);
or UO_1282 (O_1282,N_14985,N_14887);
nor UO_1283 (O_1283,N_14963,N_14979);
and UO_1284 (O_1284,N_14938,N_14971);
or UO_1285 (O_1285,N_14938,N_14881);
nor UO_1286 (O_1286,N_14829,N_14823);
nand UO_1287 (O_1287,N_14905,N_14931);
or UO_1288 (O_1288,N_14866,N_14846);
nor UO_1289 (O_1289,N_14905,N_14851);
and UO_1290 (O_1290,N_14992,N_14888);
or UO_1291 (O_1291,N_14850,N_14838);
or UO_1292 (O_1292,N_14885,N_14859);
and UO_1293 (O_1293,N_14880,N_14920);
nor UO_1294 (O_1294,N_14966,N_14994);
and UO_1295 (O_1295,N_14909,N_14803);
nand UO_1296 (O_1296,N_14973,N_14929);
nor UO_1297 (O_1297,N_14950,N_14903);
nor UO_1298 (O_1298,N_14964,N_14930);
or UO_1299 (O_1299,N_14934,N_14894);
nor UO_1300 (O_1300,N_14912,N_14842);
nor UO_1301 (O_1301,N_14818,N_14974);
and UO_1302 (O_1302,N_14935,N_14967);
xnor UO_1303 (O_1303,N_14802,N_14822);
and UO_1304 (O_1304,N_14953,N_14994);
and UO_1305 (O_1305,N_14833,N_14804);
nor UO_1306 (O_1306,N_14978,N_14851);
xnor UO_1307 (O_1307,N_14930,N_14916);
nand UO_1308 (O_1308,N_14833,N_14994);
nor UO_1309 (O_1309,N_14995,N_14961);
nor UO_1310 (O_1310,N_14870,N_14995);
nand UO_1311 (O_1311,N_14935,N_14840);
nor UO_1312 (O_1312,N_14970,N_14995);
and UO_1313 (O_1313,N_14827,N_14964);
nand UO_1314 (O_1314,N_14874,N_14847);
nand UO_1315 (O_1315,N_14922,N_14814);
or UO_1316 (O_1316,N_14874,N_14909);
nor UO_1317 (O_1317,N_14804,N_14979);
nand UO_1318 (O_1318,N_14876,N_14989);
or UO_1319 (O_1319,N_14979,N_14853);
or UO_1320 (O_1320,N_14815,N_14959);
nand UO_1321 (O_1321,N_14925,N_14829);
nand UO_1322 (O_1322,N_14850,N_14910);
nor UO_1323 (O_1323,N_14964,N_14952);
nand UO_1324 (O_1324,N_14918,N_14951);
or UO_1325 (O_1325,N_14831,N_14913);
and UO_1326 (O_1326,N_14905,N_14926);
xnor UO_1327 (O_1327,N_14890,N_14809);
or UO_1328 (O_1328,N_14838,N_14912);
nand UO_1329 (O_1329,N_14991,N_14859);
nor UO_1330 (O_1330,N_14946,N_14832);
and UO_1331 (O_1331,N_14825,N_14936);
xor UO_1332 (O_1332,N_14862,N_14813);
nand UO_1333 (O_1333,N_14873,N_14991);
or UO_1334 (O_1334,N_14889,N_14954);
and UO_1335 (O_1335,N_14825,N_14884);
and UO_1336 (O_1336,N_14874,N_14904);
and UO_1337 (O_1337,N_14945,N_14908);
xor UO_1338 (O_1338,N_14805,N_14820);
nand UO_1339 (O_1339,N_14806,N_14907);
xnor UO_1340 (O_1340,N_14832,N_14856);
xnor UO_1341 (O_1341,N_14868,N_14886);
nor UO_1342 (O_1342,N_14887,N_14917);
nor UO_1343 (O_1343,N_14845,N_14930);
nand UO_1344 (O_1344,N_14979,N_14946);
xor UO_1345 (O_1345,N_14818,N_14964);
xor UO_1346 (O_1346,N_14970,N_14912);
and UO_1347 (O_1347,N_14936,N_14851);
or UO_1348 (O_1348,N_14996,N_14878);
nor UO_1349 (O_1349,N_14977,N_14831);
nor UO_1350 (O_1350,N_14964,N_14810);
nand UO_1351 (O_1351,N_14881,N_14948);
nor UO_1352 (O_1352,N_14996,N_14949);
nand UO_1353 (O_1353,N_14949,N_14934);
or UO_1354 (O_1354,N_14934,N_14868);
xnor UO_1355 (O_1355,N_14970,N_14856);
or UO_1356 (O_1356,N_14944,N_14825);
nor UO_1357 (O_1357,N_14972,N_14902);
and UO_1358 (O_1358,N_14992,N_14895);
xor UO_1359 (O_1359,N_14915,N_14979);
xnor UO_1360 (O_1360,N_14877,N_14971);
and UO_1361 (O_1361,N_14802,N_14844);
nor UO_1362 (O_1362,N_14963,N_14834);
xnor UO_1363 (O_1363,N_14962,N_14977);
xor UO_1364 (O_1364,N_14937,N_14905);
nor UO_1365 (O_1365,N_14922,N_14995);
or UO_1366 (O_1366,N_14970,N_14933);
and UO_1367 (O_1367,N_14927,N_14871);
xor UO_1368 (O_1368,N_14803,N_14864);
xnor UO_1369 (O_1369,N_14966,N_14809);
xor UO_1370 (O_1370,N_14932,N_14866);
nand UO_1371 (O_1371,N_14930,N_14963);
nor UO_1372 (O_1372,N_14929,N_14893);
nor UO_1373 (O_1373,N_14946,N_14862);
or UO_1374 (O_1374,N_14940,N_14867);
nand UO_1375 (O_1375,N_14976,N_14915);
and UO_1376 (O_1376,N_14868,N_14941);
nor UO_1377 (O_1377,N_14856,N_14849);
xnor UO_1378 (O_1378,N_14887,N_14832);
or UO_1379 (O_1379,N_14805,N_14825);
and UO_1380 (O_1380,N_14800,N_14952);
xor UO_1381 (O_1381,N_14958,N_14927);
and UO_1382 (O_1382,N_14980,N_14984);
xor UO_1383 (O_1383,N_14868,N_14968);
nand UO_1384 (O_1384,N_14942,N_14828);
nor UO_1385 (O_1385,N_14902,N_14925);
nor UO_1386 (O_1386,N_14980,N_14986);
or UO_1387 (O_1387,N_14982,N_14873);
xor UO_1388 (O_1388,N_14876,N_14814);
and UO_1389 (O_1389,N_14825,N_14876);
nand UO_1390 (O_1390,N_14806,N_14966);
nand UO_1391 (O_1391,N_14989,N_14971);
nand UO_1392 (O_1392,N_14930,N_14865);
xor UO_1393 (O_1393,N_14871,N_14953);
xnor UO_1394 (O_1394,N_14803,N_14971);
or UO_1395 (O_1395,N_14969,N_14818);
or UO_1396 (O_1396,N_14984,N_14819);
nor UO_1397 (O_1397,N_14906,N_14948);
nor UO_1398 (O_1398,N_14828,N_14893);
or UO_1399 (O_1399,N_14882,N_14865);
or UO_1400 (O_1400,N_14898,N_14956);
nand UO_1401 (O_1401,N_14821,N_14833);
nor UO_1402 (O_1402,N_14815,N_14818);
and UO_1403 (O_1403,N_14948,N_14923);
or UO_1404 (O_1404,N_14969,N_14976);
or UO_1405 (O_1405,N_14975,N_14994);
and UO_1406 (O_1406,N_14946,N_14840);
and UO_1407 (O_1407,N_14996,N_14827);
or UO_1408 (O_1408,N_14875,N_14808);
nand UO_1409 (O_1409,N_14998,N_14854);
nand UO_1410 (O_1410,N_14980,N_14960);
xnor UO_1411 (O_1411,N_14808,N_14886);
and UO_1412 (O_1412,N_14905,N_14972);
or UO_1413 (O_1413,N_14884,N_14994);
or UO_1414 (O_1414,N_14806,N_14810);
xnor UO_1415 (O_1415,N_14947,N_14802);
and UO_1416 (O_1416,N_14870,N_14921);
xor UO_1417 (O_1417,N_14966,N_14831);
nand UO_1418 (O_1418,N_14855,N_14802);
nand UO_1419 (O_1419,N_14961,N_14828);
nand UO_1420 (O_1420,N_14856,N_14958);
nor UO_1421 (O_1421,N_14968,N_14860);
or UO_1422 (O_1422,N_14921,N_14916);
nand UO_1423 (O_1423,N_14999,N_14966);
nand UO_1424 (O_1424,N_14972,N_14932);
xor UO_1425 (O_1425,N_14813,N_14934);
and UO_1426 (O_1426,N_14803,N_14857);
nor UO_1427 (O_1427,N_14853,N_14829);
nor UO_1428 (O_1428,N_14889,N_14882);
and UO_1429 (O_1429,N_14903,N_14918);
xor UO_1430 (O_1430,N_14970,N_14899);
and UO_1431 (O_1431,N_14945,N_14888);
nand UO_1432 (O_1432,N_14959,N_14867);
and UO_1433 (O_1433,N_14923,N_14889);
xnor UO_1434 (O_1434,N_14961,N_14921);
nor UO_1435 (O_1435,N_14803,N_14856);
nor UO_1436 (O_1436,N_14962,N_14914);
or UO_1437 (O_1437,N_14942,N_14851);
and UO_1438 (O_1438,N_14959,N_14964);
nand UO_1439 (O_1439,N_14936,N_14915);
or UO_1440 (O_1440,N_14860,N_14820);
and UO_1441 (O_1441,N_14859,N_14920);
nand UO_1442 (O_1442,N_14903,N_14802);
xnor UO_1443 (O_1443,N_14890,N_14866);
nand UO_1444 (O_1444,N_14896,N_14876);
or UO_1445 (O_1445,N_14977,N_14899);
and UO_1446 (O_1446,N_14820,N_14882);
nor UO_1447 (O_1447,N_14958,N_14863);
xor UO_1448 (O_1448,N_14813,N_14989);
xor UO_1449 (O_1449,N_14987,N_14834);
or UO_1450 (O_1450,N_14916,N_14843);
or UO_1451 (O_1451,N_14853,N_14814);
and UO_1452 (O_1452,N_14800,N_14993);
nor UO_1453 (O_1453,N_14940,N_14962);
or UO_1454 (O_1454,N_14842,N_14848);
or UO_1455 (O_1455,N_14808,N_14883);
or UO_1456 (O_1456,N_14920,N_14939);
nand UO_1457 (O_1457,N_14864,N_14990);
nand UO_1458 (O_1458,N_14956,N_14953);
xnor UO_1459 (O_1459,N_14986,N_14871);
or UO_1460 (O_1460,N_14899,N_14822);
nor UO_1461 (O_1461,N_14976,N_14985);
or UO_1462 (O_1462,N_14993,N_14938);
nor UO_1463 (O_1463,N_14912,N_14882);
nand UO_1464 (O_1464,N_14956,N_14814);
and UO_1465 (O_1465,N_14873,N_14983);
or UO_1466 (O_1466,N_14872,N_14860);
or UO_1467 (O_1467,N_14942,N_14870);
and UO_1468 (O_1468,N_14921,N_14942);
nand UO_1469 (O_1469,N_14965,N_14842);
nor UO_1470 (O_1470,N_14845,N_14830);
nor UO_1471 (O_1471,N_14990,N_14968);
xor UO_1472 (O_1472,N_14942,N_14819);
and UO_1473 (O_1473,N_14812,N_14904);
or UO_1474 (O_1474,N_14834,N_14813);
xor UO_1475 (O_1475,N_14839,N_14893);
nand UO_1476 (O_1476,N_14989,N_14892);
or UO_1477 (O_1477,N_14943,N_14807);
nor UO_1478 (O_1478,N_14875,N_14941);
or UO_1479 (O_1479,N_14851,N_14888);
nor UO_1480 (O_1480,N_14909,N_14884);
or UO_1481 (O_1481,N_14915,N_14937);
xor UO_1482 (O_1482,N_14848,N_14851);
and UO_1483 (O_1483,N_14814,N_14861);
or UO_1484 (O_1484,N_14869,N_14940);
xnor UO_1485 (O_1485,N_14848,N_14960);
nor UO_1486 (O_1486,N_14938,N_14878);
and UO_1487 (O_1487,N_14849,N_14872);
nand UO_1488 (O_1488,N_14955,N_14879);
or UO_1489 (O_1489,N_14981,N_14816);
xnor UO_1490 (O_1490,N_14964,N_14925);
xnor UO_1491 (O_1491,N_14898,N_14926);
nor UO_1492 (O_1492,N_14883,N_14936);
xnor UO_1493 (O_1493,N_14879,N_14948);
xor UO_1494 (O_1494,N_14987,N_14927);
and UO_1495 (O_1495,N_14954,N_14920);
or UO_1496 (O_1496,N_14902,N_14912);
or UO_1497 (O_1497,N_14877,N_14879);
nand UO_1498 (O_1498,N_14939,N_14888);
nand UO_1499 (O_1499,N_14936,N_14889);
and UO_1500 (O_1500,N_14875,N_14889);
nor UO_1501 (O_1501,N_14815,N_14812);
or UO_1502 (O_1502,N_14910,N_14951);
nor UO_1503 (O_1503,N_14811,N_14868);
nor UO_1504 (O_1504,N_14957,N_14855);
or UO_1505 (O_1505,N_14864,N_14862);
nor UO_1506 (O_1506,N_14987,N_14993);
nor UO_1507 (O_1507,N_14942,N_14989);
nand UO_1508 (O_1508,N_14880,N_14856);
xnor UO_1509 (O_1509,N_14832,N_14927);
nand UO_1510 (O_1510,N_14878,N_14982);
and UO_1511 (O_1511,N_14942,N_14933);
and UO_1512 (O_1512,N_14936,N_14930);
nor UO_1513 (O_1513,N_14995,N_14834);
nand UO_1514 (O_1514,N_14816,N_14833);
and UO_1515 (O_1515,N_14873,N_14934);
or UO_1516 (O_1516,N_14974,N_14865);
xnor UO_1517 (O_1517,N_14970,N_14917);
and UO_1518 (O_1518,N_14841,N_14908);
nand UO_1519 (O_1519,N_14933,N_14820);
and UO_1520 (O_1520,N_14853,N_14872);
nand UO_1521 (O_1521,N_14919,N_14801);
xnor UO_1522 (O_1522,N_14814,N_14955);
xnor UO_1523 (O_1523,N_14885,N_14828);
and UO_1524 (O_1524,N_14957,N_14882);
nand UO_1525 (O_1525,N_14984,N_14969);
or UO_1526 (O_1526,N_14891,N_14922);
and UO_1527 (O_1527,N_14975,N_14897);
or UO_1528 (O_1528,N_14999,N_14866);
and UO_1529 (O_1529,N_14996,N_14874);
nand UO_1530 (O_1530,N_14980,N_14853);
nand UO_1531 (O_1531,N_14858,N_14974);
nor UO_1532 (O_1532,N_14915,N_14997);
xnor UO_1533 (O_1533,N_14884,N_14961);
or UO_1534 (O_1534,N_14985,N_14963);
nand UO_1535 (O_1535,N_14898,N_14854);
nand UO_1536 (O_1536,N_14931,N_14945);
xor UO_1537 (O_1537,N_14898,N_14804);
nand UO_1538 (O_1538,N_14864,N_14890);
or UO_1539 (O_1539,N_14904,N_14825);
and UO_1540 (O_1540,N_14915,N_14956);
and UO_1541 (O_1541,N_14939,N_14864);
or UO_1542 (O_1542,N_14826,N_14920);
nand UO_1543 (O_1543,N_14845,N_14984);
xor UO_1544 (O_1544,N_14937,N_14878);
nand UO_1545 (O_1545,N_14821,N_14923);
nor UO_1546 (O_1546,N_14943,N_14965);
or UO_1547 (O_1547,N_14992,N_14919);
and UO_1548 (O_1548,N_14965,N_14985);
and UO_1549 (O_1549,N_14832,N_14923);
and UO_1550 (O_1550,N_14839,N_14988);
or UO_1551 (O_1551,N_14991,N_14901);
nor UO_1552 (O_1552,N_14929,N_14891);
xnor UO_1553 (O_1553,N_14801,N_14847);
nand UO_1554 (O_1554,N_14887,N_14956);
nor UO_1555 (O_1555,N_14920,N_14970);
and UO_1556 (O_1556,N_14996,N_14981);
and UO_1557 (O_1557,N_14944,N_14927);
nor UO_1558 (O_1558,N_14832,N_14992);
nor UO_1559 (O_1559,N_14874,N_14950);
xor UO_1560 (O_1560,N_14864,N_14896);
or UO_1561 (O_1561,N_14825,N_14973);
and UO_1562 (O_1562,N_14807,N_14994);
xor UO_1563 (O_1563,N_14873,N_14834);
xnor UO_1564 (O_1564,N_14895,N_14883);
xor UO_1565 (O_1565,N_14999,N_14970);
nor UO_1566 (O_1566,N_14901,N_14903);
nand UO_1567 (O_1567,N_14930,N_14921);
xor UO_1568 (O_1568,N_14854,N_14907);
and UO_1569 (O_1569,N_14947,N_14983);
nor UO_1570 (O_1570,N_14873,N_14874);
nand UO_1571 (O_1571,N_14958,N_14821);
nor UO_1572 (O_1572,N_14890,N_14889);
xnor UO_1573 (O_1573,N_14942,N_14886);
nand UO_1574 (O_1574,N_14904,N_14943);
and UO_1575 (O_1575,N_14976,N_14999);
xor UO_1576 (O_1576,N_14963,N_14994);
and UO_1577 (O_1577,N_14998,N_14909);
xnor UO_1578 (O_1578,N_14870,N_14979);
xnor UO_1579 (O_1579,N_14874,N_14920);
or UO_1580 (O_1580,N_14950,N_14829);
nand UO_1581 (O_1581,N_14821,N_14933);
xor UO_1582 (O_1582,N_14886,N_14880);
or UO_1583 (O_1583,N_14886,N_14896);
nor UO_1584 (O_1584,N_14887,N_14979);
and UO_1585 (O_1585,N_14961,N_14808);
nand UO_1586 (O_1586,N_14919,N_14834);
nor UO_1587 (O_1587,N_14959,N_14886);
or UO_1588 (O_1588,N_14998,N_14832);
or UO_1589 (O_1589,N_14919,N_14898);
nand UO_1590 (O_1590,N_14890,N_14979);
xnor UO_1591 (O_1591,N_14892,N_14825);
nor UO_1592 (O_1592,N_14832,N_14970);
nand UO_1593 (O_1593,N_14918,N_14881);
nor UO_1594 (O_1594,N_14940,N_14943);
nand UO_1595 (O_1595,N_14877,N_14859);
nand UO_1596 (O_1596,N_14992,N_14814);
nor UO_1597 (O_1597,N_14970,N_14848);
xor UO_1598 (O_1598,N_14829,N_14915);
and UO_1599 (O_1599,N_14802,N_14904);
nor UO_1600 (O_1600,N_14921,N_14904);
xor UO_1601 (O_1601,N_14977,N_14805);
and UO_1602 (O_1602,N_14979,N_14857);
or UO_1603 (O_1603,N_14811,N_14825);
nor UO_1604 (O_1604,N_14984,N_14815);
nor UO_1605 (O_1605,N_14882,N_14920);
and UO_1606 (O_1606,N_14829,N_14888);
xor UO_1607 (O_1607,N_14947,N_14847);
nand UO_1608 (O_1608,N_14977,N_14871);
or UO_1609 (O_1609,N_14839,N_14884);
xnor UO_1610 (O_1610,N_14984,N_14859);
nand UO_1611 (O_1611,N_14816,N_14827);
and UO_1612 (O_1612,N_14820,N_14852);
and UO_1613 (O_1613,N_14932,N_14971);
xnor UO_1614 (O_1614,N_14805,N_14849);
and UO_1615 (O_1615,N_14946,N_14825);
and UO_1616 (O_1616,N_14917,N_14975);
and UO_1617 (O_1617,N_14955,N_14947);
nor UO_1618 (O_1618,N_14862,N_14942);
or UO_1619 (O_1619,N_14856,N_14911);
or UO_1620 (O_1620,N_14826,N_14870);
nand UO_1621 (O_1621,N_14905,N_14940);
xnor UO_1622 (O_1622,N_14819,N_14990);
and UO_1623 (O_1623,N_14826,N_14888);
xnor UO_1624 (O_1624,N_14889,N_14997);
xnor UO_1625 (O_1625,N_14876,N_14943);
nor UO_1626 (O_1626,N_14937,N_14982);
nor UO_1627 (O_1627,N_14987,N_14829);
nor UO_1628 (O_1628,N_14875,N_14970);
or UO_1629 (O_1629,N_14854,N_14808);
nand UO_1630 (O_1630,N_14810,N_14820);
xnor UO_1631 (O_1631,N_14808,N_14860);
nand UO_1632 (O_1632,N_14856,N_14942);
and UO_1633 (O_1633,N_14847,N_14971);
xor UO_1634 (O_1634,N_14919,N_14914);
nor UO_1635 (O_1635,N_14884,N_14823);
nor UO_1636 (O_1636,N_14850,N_14825);
nor UO_1637 (O_1637,N_14835,N_14810);
and UO_1638 (O_1638,N_14984,N_14811);
nand UO_1639 (O_1639,N_14998,N_14964);
and UO_1640 (O_1640,N_14836,N_14838);
or UO_1641 (O_1641,N_14831,N_14835);
nand UO_1642 (O_1642,N_14953,N_14806);
and UO_1643 (O_1643,N_14815,N_14950);
or UO_1644 (O_1644,N_14972,N_14842);
and UO_1645 (O_1645,N_14886,N_14814);
or UO_1646 (O_1646,N_14806,N_14901);
and UO_1647 (O_1647,N_14931,N_14976);
xor UO_1648 (O_1648,N_14830,N_14840);
and UO_1649 (O_1649,N_14940,N_14872);
or UO_1650 (O_1650,N_14813,N_14980);
and UO_1651 (O_1651,N_14847,N_14890);
or UO_1652 (O_1652,N_14962,N_14874);
and UO_1653 (O_1653,N_14986,N_14885);
nand UO_1654 (O_1654,N_14902,N_14861);
nand UO_1655 (O_1655,N_14832,N_14961);
nand UO_1656 (O_1656,N_14822,N_14821);
nand UO_1657 (O_1657,N_14835,N_14948);
or UO_1658 (O_1658,N_14958,N_14839);
nand UO_1659 (O_1659,N_14945,N_14926);
nor UO_1660 (O_1660,N_14859,N_14904);
nor UO_1661 (O_1661,N_14945,N_14977);
and UO_1662 (O_1662,N_14933,N_14988);
xnor UO_1663 (O_1663,N_14881,N_14911);
nor UO_1664 (O_1664,N_14848,N_14993);
and UO_1665 (O_1665,N_14828,N_14806);
nor UO_1666 (O_1666,N_14950,N_14972);
nor UO_1667 (O_1667,N_14888,N_14907);
or UO_1668 (O_1668,N_14974,N_14919);
nand UO_1669 (O_1669,N_14846,N_14849);
xor UO_1670 (O_1670,N_14995,N_14947);
or UO_1671 (O_1671,N_14859,N_14940);
nor UO_1672 (O_1672,N_14846,N_14998);
nand UO_1673 (O_1673,N_14833,N_14985);
xnor UO_1674 (O_1674,N_14953,N_14819);
or UO_1675 (O_1675,N_14939,N_14914);
or UO_1676 (O_1676,N_14982,N_14932);
xnor UO_1677 (O_1677,N_14959,N_14873);
nand UO_1678 (O_1678,N_14866,N_14875);
or UO_1679 (O_1679,N_14874,N_14945);
and UO_1680 (O_1680,N_14811,N_14914);
nor UO_1681 (O_1681,N_14835,N_14970);
xor UO_1682 (O_1682,N_14828,N_14998);
nand UO_1683 (O_1683,N_14909,N_14947);
nand UO_1684 (O_1684,N_14969,N_14889);
nand UO_1685 (O_1685,N_14863,N_14842);
nand UO_1686 (O_1686,N_14861,N_14969);
nand UO_1687 (O_1687,N_14986,N_14888);
nor UO_1688 (O_1688,N_14951,N_14940);
xnor UO_1689 (O_1689,N_14959,N_14952);
nor UO_1690 (O_1690,N_14868,N_14876);
or UO_1691 (O_1691,N_14972,N_14934);
or UO_1692 (O_1692,N_14854,N_14929);
nand UO_1693 (O_1693,N_14941,N_14905);
xnor UO_1694 (O_1694,N_14996,N_14800);
nor UO_1695 (O_1695,N_14899,N_14973);
xor UO_1696 (O_1696,N_14973,N_14952);
or UO_1697 (O_1697,N_14919,N_14884);
or UO_1698 (O_1698,N_14825,N_14907);
nor UO_1699 (O_1699,N_14996,N_14818);
and UO_1700 (O_1700,N_14938,N_14984);
nand UO_1701 (O_1701,N_14917,N_14872);
nor UO_1702 (O_1702,N_14908,N_14870);
or UO_1703 (O_1703,N_14824,N_14942);
or UO_1704 (O_1704,N_14977,N_14813);
nand UO_1705 (O_1705,N_14997,N_14996);
nor UO_1706 (O_1706,N_14979,N_14936);
nor UO_1707 (O_1707,N_14926,N_14918);
or UO_1708 (O_1708,N_14970,N_14837);
nor UO_1709 (O_1709,N_14891,N_14801);
nand UO_1710 (O_1710,N_14879,N_14809);
nand UO_1711 (O_1711,N_14936,N_14964);
nor UO_1712 (O_1712,N_14844,N_14990);
or UO_1713 (O_1713,N_14966,N_14950);
nand UO_1714 (O_1714,N_14810,N_14848);
and UO_1715 (O_1715,N_14838,N_14859);
nor UO_1716 (O_1716,N_14950,N_14911);
or UO_1717 (O_1717,N_14849,N_14834);
nor UO_1718 (O_1718,N_14804,N_14829);
and UO_1719 (O_1719,N_14908,N_14966);
nor UO_1720 (O_1720,N_14990,N_14866);
xnor UO_1721 (O_1721,N_14832,N_14984);
nand UO_1722 (O_1722,N_14892,N_14910);
nor UO_1723 (O_1723,N_14879,N_14859);
or UO_1724 (O_1724,N_14805,N_14811);
nor UO_1725 (O_1725,N_14991,N_14858);
or UO_1726 (O_1726,N_14999,N_14893);
xor UO_1727 (O_1727,N_14902,N_14849);
and UO_1728 (O_1728,N_14921,N_14976);
and UO_1729 (O_1729,N_14806,N_14879);
xor UO_1730 (O_1730,N_14920,N_14978);
or UO_1731 (O_1731,N_14975,N_14893);
nand UO_1732 (O_1732,N_14973,N_14803);
nor UO_1733 (O_1733,N_14875,N_14842);
and UO_1734 (O_1734,N_14816,N_14884);
nand UO_1735 (O_1735,N_14932,N_14897);
and UO_1736 (O_1736,N_14812,N_14856);
xor UO_1737 (O_1737,N_14895,N_14848);
xor UO_1738 (O_1738,N_14894,N_14818);
nand UO_1739 (O_1739,N_14933,N_14816);
and UO_1740 (O_1740,N_14944,N_14904);
or UO_1741 (O_1741,N_14985,N_14842);
and UO_1742 (O_1742,N_14842,N_14926);
and UO_1743 (O_1743,N_14881,N_14945);
and UO_1744 (O_1744,N_14929,N_14932);
and UO_1745 (O_1745,N_14802,N_14993);
xor UO_1746 (O_1746,N_14977,N_14964);
xor UO_1747 (O_1747,N_14860,N_14934);
nor UO_1748 (O_1748,N_14940,N_14860);
nand UO_1749 (O_1749,N_14911,N_14879);
xor UO_1750 (O_1750,N_14802,N_14885);
xor UO_1751 (O_1751,N_14842,N_14990);
nand UO_1752 (O_1752,N_14843,N_14999);
and UO_1753 (O_1753,N_14862,N_14829);
xor UO_1754 (O_1754,N_14839,N_14804);
or UO_1755 (O_1755,N_14899,N_14949);
nand UO_1756 (O_1756,N_14980,N_14978);
nand UO_1757 (O_1757,N_14913,N_14834);
nand UO_1758 (O_1758,N_14817,N_14925);
or UO_1759 (O_1759,N_14926,N_14986);
and UO_1760 (O_1760,N_14883,N_14811);
nand UO_1761 (O_1761,N_14948,N_14814);
and UO_1762 (O_1762,N_14868,N_14989);
xnor UO_1763 (O_1763,N_14893,N_14931);
or UO_1764 (O_1764,N_14862,N_14956);
or UO_1765 (O_1765,N_14957,N_14938);
or UO_1766 (O_1766,N_14930,N_14834);
nand UO_1767 (O_1767,N_14820,N_14833);
xnor UO_1768 (O_1768,N_14893,N_14864);
and UO_1769 (O_1769,N_14863,N_14987);
and UO_1770 (O_1770,N_14882,N_14872);
or UO_1771 (O_1771,N_14810,N_14800);
xnor UO_1772 (O_1772,N_14997,N_14801);
or UO_1773 (O_1773,N_14880,N_14927);
or UO_1774 (O_1774,N_14854,N_14966);
xnor UO_1775 (O_1775,N_14995,N_14984);
nand UO_1776 (O_1776,N_14879,N_14967);
and UO_1777 (O_1777,N_14894,N_14813);
or UO_1778 (O_1778,N_14905,N_14917);
xor UO_1779 (O_1779,N_14808,N_14898);
nor UO_1780 (O_1780,N_14833,N_14807);
and UO_1781 (O_1781,N_14846,N_14982);
and UO_1782 (O_1782,N_14914,N_14885);
nand UO_1783 (O_1783,N_14827,N_14839);
or UO_1784 (O_1784,N_14809,N_14803);
xnor UO_1785 (O_1785,N_14936,N_14865);
nor UO_1786 (O_1786,N_14897,N_14938);
nand UO_1787 (O_1787,N_14804,N_14942);
or UO_1788 (O_1788,N_14910,N_14992);
or UO_1789 (O_1789,N_14852,N_14965);
xor UO_1790 (O_1790,N_14936,N_14871);
nor UO_1791 (O_1791,N_14959,N_14903);
xor UO_1792 (O_1792,N_14815,N_14912);
or UO_1793 (O_1793,N_14960,N_14930);
nor UO_1794 (O_1794,N_14837,N_14941);
nor UO_1795 (O_1795,N_14871,N_14882);
xor UO_1796 (O_1796,N_14945,N_14821);
nand UO_1797 (O_1797,N_14814,N_14919);
xnor UO_1798 (O_1798,N_14951,N_14822);
and UO_1799 (O_1799,N_14831,N_14982);
xor UO_1800 (O_1800,N_14834,N_14991);
nand UO_1801 (O_1801,N_14981,N_14869);
nor UO_1802 (O_1802,N_14933,N_14872);
and UO_1803 (O_1803,N_14930,N_14822);
nand UO_1804 (O_1804,N_14829,N_14816);
xor UO_1805 (O_1805,N_14860,N_14832);
nor UO_1806 (O_1806,N_14902,N_14924);
and UO_1807 (O_1807,N_14946,N_14815);
xnor UO_1808 (O_1808,N_14912,N_14971);
xor UO_1809 (O_1809,N_14818,N_14866);
nor UO_1810 (O_1810,N_14843,N_14838);
nand UO_1811 (O_1811,N_14868,N_14838);
xnor UO_1812 (O_1812,N_14854,N_14948);
xnor UO_1813 (O_1813,N_14876,N_14886);
xor UO_1814 (O_1814,N_14800,N_14856);
nor UO_1815 (O_1815,N_14994,N_14926);
nor UO_1816 (O_1816,N_14996,N_14868);
nor UO_1817 (O_1817,N_14915,N_14832);
xor UO_1818 (O_1818,N_14961,N_14996);
and UO_1819 (O_1819,N_14885,N_14974);
xnor UO_1820 (O_1820,N_14941,N_14884);
and UO_1821 (O_1821,N_14809,N_14939);
nand UO_1822 (O_1822,N_14808,N_14952);
and UO_1823 (O_1823,N_14984,N_14836);
nor UO_1824 (O_1824,N_14937,N_14824);
xnor UO_1825 (O_1825,N_14964,N_14880);
nor UO_1826 (O_1826,N_14914,N_14903);
and UO_1827 (O_1827,N_14956,N_14901);
nand UO_1828 (O_1828,N_14985,N_14838);
nor UO_1829 (O_1829,N_14961,N_14814);
nand UO_1830 (O_1830,N_14917,N_14937);
xnor UO_1831 (O_1831,N_14929,N_14926);
nand UO_1832 (O_1832,N_14855,N_14856);
nor UO_1833 (O_1833,N_14814,N_14832);
nand UO_1834 (O_1834,N_14977,N_14952);
and UO_1835 (O_1835,N_14873,N_14909);
nand UO_1836 (O_1836,N_14837,N_14851);
nand UO_1837 (O_1837,N_14888,N_14959);
nor UO_1838 (O_1838,N_14817,N_14872);
and UO_1839 (O_1839,N_14971,N_14815);
and UO_1840 (O_1840,N_14920,N_14985);
xnor UO_1841 (O_1841,N_14915,N_14891);
nand UO_1842 (O_1842,N_14914,N_14801);
xnor UO_1843 (O_1843,N_14963,N_14939);
and UO_1844 (O_1844,N_14896,N_14990);
nor UO_1845 (O_1845,N_14966,N_14816);
nand UO_1846 (O_1846,N_14883,N_14829);
or UO_1847 (O_1847,N_14958,N_14848);
or UO_1848 (O_1848,N_14812,N_14846);
or UO_1849 (O_1849,N_14952,N_14939);
and UO_1850 (O_1850,N_14947,N_14891);
xor UO_1851 (O_1851,N_14816,N_14881);
xnor UO_1852 (O_1852,N_14989,N_14966);
and UO_1853 (O_1853,N_14857,N_14801);
xor UO_1854 (O_1854,N_14923,N_14955);
xnor UO_1855 (O_1855,N_14993,N_14974);
nor UO_1856 (O_1856,N_14863,N_14951);
xnor UO_1857 (O_1857,N_14804,N_14811);
or UO_1858 (O_1858,N_14954,N_14926);
and UO_1859 (O_1859,N_14828,N_14976);
nor UO_1860 (O_1860,N_14930,N_14934);
and UO_1861 (O_1861,N_14883,N_14996);
and UO_1862 (O_1862,N_14865,N_14911);
or UO_1863 (O_1863,N_14937,N_14877);
xor UO_1864 (O_1864,N_14950,N_14948);
and UO_1865 (O_1865,N_14914,N_14960);
nor UO_1866 (O_1866,N_14871,N_14935);
nor UO_1867 (O_1867,N_14954,N_14862);
and UO_1868 (O_1868,N_14949,N_14875);
and UO_1869 (O_1869,N_14940,N_14812);
xnor UO_1870 (O_1870,N_14956,N_14900);
and UO_1871 (O_1871,N_14899,N_14901);
xor UO_1872 (O_1872,N_14842,N_14910);
xnor UO_1873 (O_1873,N_14964,N_14927);
nor UO_1874 (O_1874,N_14989,N_14804);
nor UO_1875 (O_1875,N_14807,N_14858);
or UO_1876 (O_1876,N_14912,N_14949);
or UO_1877 (O_1877,N_14840,N_14880);
nor UO_1878 (O_1878,N_14966,N_14821);
or UO_1879 (O_1879,N_14869,N_14985);
nor UO_1880 (O_1880,N_14967,N_14886);
nor UO_1881 (O_1881,N_14837,N_14847);
nand UO_1882 (O_1882,N_14996,N_14923);
and UO_1883 (O_1883,N_14811,N_14992);
nor UO_1884 (O_1884,N_14978,N_14944);
or UO_1885 (O_1885,N_14859,N_14808);
nor UO_1886 (O_1886,N_14843,N_14856);
xor UO_1887 (O_1887,N_14935,N_14995);
xor UO_1888 (O_1888,N_14877,N_14848);
nor UO_1889 (O_1889,N_14963,N_14967);
xnor UO_1890 (O_1890,N_14914,N_14909);
or UO_1891 (O_1891,N_14932,N_14893);
nand UO_1892 (O_1892,N_14807,N_14905);
xnor UO_1893 (O_1893,N_14833,N_14828);
or UO_1894 (O_1894,N_14967,N_14929);
or UO_1895 (O_1895,N_14891,N_14980);
and UO_1896 (O_1896,N_14942,N_14953);
or UO_1897 (O_1897,N_14946,N_14966);
or UO_1898 (O_1898,N_14971,N_14948);
nand UO_1899 (O_1899,N_14912,N_14811);
nand UO_1900 (O_1900,N_14867,N_14943);
or UO_1901 (O_1901,N_14947,N_14882);
xor UO_1902 (O_1902,N_14832,N_14827);
nand UO_1903 (O_1903,N_14986,N_14901);
xnor UO_1904 (O_1904,N_14812,N_14898);
nand UO_1905 (O_1905,N_14968,N_14997);
or UO_1906 (O_1906,N_14936,N_14950);
and UO_1907 (O_1907,N_14960,N_14846);
and UO_1908 (O_1908,N_14978,N_14800);
and UO_1909 (O_1909,N_14830,N_14991);
nand UO_1910 (O_1910,N_14932,N_14883);
nand UO_1911 (O_1911,N_14928,N_14987);
and UO_1912 (O_1912,N_14898,N_14892);
xor UO_1913 (O_1913,N_14902,N_14962);
nand UO_1914 (O_1914,N_14939,N_14926);
and UO_1915 (O_1915,N_14919,N_14903);
nor UO_1916 (O_1916,N_14947,N_14901);
nor UO_1917 (O_1917,N_14920,N_14883);
and UO_1918 (O_1918,N_14887,N_14977);
nor UO_1919 (O_1919,N_14809,N_14988);
xnor UO_1920 (O_1920,N_14805,N_14985);
and UO_1921 (O_1921,N_14931,N_14993);
xor UO_1922 (O_1922,N_14895,N_14835);
and UO_1923 (O_1923,N_14970,N_14943);
and UO_1924 (O_1924,N_14824,N_14910);
or UO_1925 (O_1925,N_14942,N_14904);
nand UO_1926 (O_1926,N_14861,N_14940);
and UO_1927 (O_1927,N_14817,N_14934);
xnor UO_1928 (O_1928,N_14882,N_14884);
or UO_1929 (O_1929,N_14855,N_14889);
and UO_1930 (O_1930,N_14934,N_14851);
or UO_1931 (O_1931,N_14824,N_14821);
or UO_1932 (O_1932,N_14936,N_14866);
or UO_1933 (O_1933,N_14892,N_14882);
xor UO_1934 (O_1934,N_14930,N_14872);
nor UO_1935 (O_1935,N_14927,N_14823);
or UO_1936 (O_1936,N_14886,N_14841);
or UO_1937 (O_1937,N_14895,N_14887);
and UO_1938 (O_1938,N_14852,N_14926);
nand UO_1939 (O_1939,N_14821,N_14931);
xnor UO_1940 (O_1940,N_14875,N_14894);
nor UO_1941 (O_1941,N_14852,N_14920);
xnor UO_1942 (O_1942,N_14857,N_14908);
or UO_1943 (O_1943,N_14934,N_14998);
nor UO_1944 (O_1944,N_14969,N_14979);
and UO_1945 (O_1945,N_14890,N_14893);
xnor UO_1946 (O_1946,N_14924,N_14830);
nor UO_1947 (O_1947,N_14865,N_14844);
xor UO_1948 (O_1948,N_14964,N_14833);
nor UO_1949 (O_1949,N_14945,N_14839);
and UO_1950 (O_1950,N_14824,N_14803);
and UO_1951 (O_1951,N_14926,N_14982);
and UO_1952 (O_1952,N_14862,N_14999);
nand UO_1953 (O_1953,N_14969,N_14806);
and UO_1954 (O_1954,N_14952,N_14860);
or UO_1955 (O_1955,N_14859,N_14951);
nor UO_1956 (O_1956,N_14929,N_14953);
nand UO_1957 (O_1957,N_14919,N_14887);
nor UO_1958 (O_1958,N_14983,N_14926);
and UO_1959 (O_1959,N_14823,N_14853);
nand UO_1960 (O_1960,N_14812,N_14996);
nand UO_1961 (O_1961,N_14969,N_14960);
nor UO_1962 (O_1962,N_14979,N_14988);
nand UO_1963 (O_1963,N_14886,N_14818);
xnor UO_1964 (O_1964,N_14888,N_14868);
xnor UO_1965 (O_1965,N_14832,N_14919);
xnor UO_1966 (O_1966,N_14984,N_14857);
nor UO_1967 (O_1967,N_14853,N_14927);
xor UO_1968 (O_1968,N_14823,N_14969);
nand UO_1969 (O_1969,N_14887,N_14907);
nand UO_1970 (O_1970,N_14956,N_14945);
nor UO_1971 (O_1971,N_14999,N_14909);
xnor UO_1972 (O_1972,N_14849,N_14993);
nand UO_1973 (O_1973,N_14913,N_14843);
or UO_1974 (O_1974,N_14874,N_14881);
nand UO_1975 (O_1975,N_14834,N_14932);
xor UO_1976 (O_1976,N_14858,N_14824);
nand UO_1977 (O_1977,N_14989,N_14817);
and UO_1978 (O_1978,N_14948,N_14945);
xnor UO_1979 (O_1979,N_14962,N_14913);
nand UO_1980 (O_1980,N_14829,N_14877);
and UO_1981 (O_1981,N_14900,N_14985);
xnor UO_1982 (O_1982,N_14866,N_14966);
and UO_1983 (O_1983,N_14957,N_14800);
nand UO_1984 (O_1984,N_14873,N_14884);
nor UO_1985 (O_1985,N_14802,N_14831);
xor UO_1986 (O_1986,N_14946,N_14811);
or UO_1987 (O_1987,N_14915,N_14930);
xor UO_1988 (O_1988,N_14828,N_14963);
nor UO_1989 (O_1989,N_14956,N_14886);
xor UO_1990 (O_1990,N_14958,N_14882);
nand UO_1991 (O_1991,N_14821,N_14862);
nand UO_1992 (O_1992,N_14949,N_14873);
xnor UO_1993 (O_1993,N_14963,N_14966);
and UO_1994 (O_1994,N_14918,N_14945);
nor UO_1995 (O_1995,N_14939,N_14860);
nand UO_1996 (O_1996,N_14903,N_14986);
nor UO_1997 (O_1997,N_14818,N_14811);
or UO_1998 (O_1998,N_14805,N_14979);
nor UO_1999 (O_1999,N_14977,N_14900);
endmodule