module basic_1500_15000_2000_60_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_989,In_232);
and U1 (N_1,In_837,In_346);
nor U2 (N_2,In_1030,In_1458);
and U3 (N_3,In_171,In_279);
xnor U4 (N_4,In_1005,In_1400);
or U5 (N_5,In_804,In_391);
nor U6 (N_6,In_277,In_67);
nor U7 (N_7,In_1244,In_927);
nand U8 (N_8,In_1462,In_113);
or U9 (N_9,In_2,In_496);
and U10 (N_10,In_1390,In_302);
nand U11 (N_11,In_883,In_459);
or U12 (N_12,In_271,In_1253);
nand U13 (N_13,In_223,In_1389);
nor U14 (N_14,In_1350,In_506);
xnor U15 (N_15,In_1305,In_153);
or U16 (N_16,In_920,In_123);
and U17 (N_17,In_1054,In_1255);
nor U18 (N_18,In_1203,In_493);
nor U19 (N_19,In_1314,In_1316);
and U20 (N_20,In_1116,In_449);
nor U21 (N_21,In_559,In_889);
and U22 (N_22,In_106,In_1249);
xor U23 (N_23,In_316,In_574);
xnor U24 (N_24,In_1185,In_1242);
or U25 (N_25,In_1236,In_1490);
xnor U26 (N_26,In_761,In_377);
nor U27 (N_27,In_652,In_135);
xor U28 (N_28,In_1359,In_941);
or U29 (N_29,In_1274,In_370);
xnor U30 (N_30,In_1156,In_794);
xnor U31 (N_31,In_251,In_220);
xor U32 (N_32,In_485,In_886);
and U33 (N_33,In_387,In_1263);
xor U34 (N_34,In_1465,In_352);
xnor U35 (N_35,In_748,In_1097);
and U36 (N_36,In_1321,In_473);
nand U37 (N_37,In_210,In_1016);
and U38 (N_38,In_368,In_1167);
nand U39 (N_39,In_1007,In_61);
nor U40 (N_40,In_408,In_1399);
and U41 (N_41,In_772,In_1378);
nand U42 (N_42,In_519,In_914);
nand U43 (N_43,In_584,In_612);
nor U44 (N_44,In_890,In_602);
nor U45 (N_45,In_245,In_747);
and U46 (N_46,In_190,In_1163);
nor U47 (N_47,In_758,In_715);
or U48 (N_48,In_788,In_676);
nor U49 (N_49,In_1320,In_231);
nor U50 (N_50,In_1109,In_207);
and U51 (N_51,In_1260,In_344);
and U52 (N_52,In_1269,In_702);
nor U53 (N_53,In_1094,In_236);
and U54 (N_54,In_32,In_509);
xor U55 (N_55,In_1080,In_563);
or U56 (N_56,In_1391,In_867);
xnor U57 (N_57,In_970,In_1322);
xnor U58 (N_58,In_198,In_813);
or U59 (N_59,In_751,In_1150);
nor U60 (N_60,In_900,In_894);
xnor U61 (N_61,In_1171,In_982);
nor U62 (N_62,In_446,In_1394);
nor U63 (N_63,In_1124,In_1076);
and U64 (N_64,In_875,In_329);
or U65 (N_65,In_1277,In_926);
nor U66 (N_66,In_997,In_293);
or U67 (N_67,In_1198,In_1376);
nor U68 (N_68,In_218,In_1197);
nand U69 (N_69,In_666,In_301);
xnor U70 (N_70,In_1049,In_441);
and U71 (N_71,In_1207,In_439);
xor U72 (N_72,In_1368,In_1216);
and U73 (N_73,In_869,In_505);
nor U74 (N_74,In_242,In_510);
and U75 (N_75,In_540,In_1215);
xor U76 (N_76,In_836,In_1011);
or U77 (N_77,In_925,In_263);
nor U78 (N_78,In_763,In_39);
nor U79 (N_79,In_1132,In_1143);
or U80 (N_80,In_697,In_394);
xnor U81 (N_81,In_1370,In_779);
nor U82 (N_82,In_1302,In_1445);
xor U83 (N_83,In_1038,In_1308);
nand U84 (N_84,In_351,In_206);
and U85 (N_85,In_252,In_1467);
and U86 (N_86,In_1159,In_1276);
or U87 (N_87,In_1023,In_11);
nand U88 (N_88,In_1375,In_1443);
and U89 (N_89,In_572,In_1230);
xnor U90 (N_90,In_60,In_1444);
or U91 (N_91,In_250,In_823);
xnor U92 (N_92,In_1463,In_580);
nor U93 (N_93,In_1258,In_1295);
nand U94 (N_94,In_466,In_1284);
nand U95 (N_95,In_288,In_1093);
nor U96 (N_96,In_1272,In_115);
or U97 (N_97,In_931,In_498);
nor U98 (N_98,In_740,In_627);
nand U99 (N_99,In_332,In_805);
or U100 (N_100,In_91,In_76);
and U101 (N_101,In_303,In_378);
or U102 (N_102,In_756,In_134);
and U103 (N_103,In_281,In_1271);
nor U104 (N_104,In_428,In_735);
nand U105 (N_105,In_599,In_128);
and U106 (N_106,In_561,In_807);
nand U107 (N_107,In_988,In_596);
nor U108 (N_108,In_895,In_1128);
xor U109 (N_109,In_1352,In_1256);
xnor U110 (N_110,In_1142,In_1369);
nor U111 (N_111,In_986,In_284);
or U112 (N_112,In_1425,In_573);
or U113 (N_113,In_484,In_991);
xnor U114 (N_114,In_1144,In_609);
and U115 (N_115,In_624,In_945);
or U116 (N_116,In_582,In_832);
and U117 (N_117,In_347,In_766);
nand U118 (N_118,In_818,In_1432);
or U119 (N_119,In_422,In_1181);
nand U120 (N_120,In_1485,In_354);
xnor U121 (N_121,In_1309,In_814);
xnor U122 (N_122,In_111,In_1092);
nand U123 (N_123,In_307,In_369);
or U124 (N_124,In_732,In_692);
or U125 (N_125,In_1060,In_502);
nand U126 (N_126,In_1146,In_690);
and U127 (N_127,In_99,In_83);
nand U128 (N_128,In_1053,In_500);
and U129 (N_129,In_1015,In_225);
or U130 (N_130,In_166,In_124);
nand U131 (N_131,In_977,In_1491);
or U132 (N_132,In_918,In_825);
xnor U133 (N_133,In_152,In_258);
nor U134 (N_134,In_4,In_226);
and U135 (N_135,In_214,In_170);
nand U136 (N_136,In_736,In_173);
xnor U137 (N_137,In_1211,In_129);
nor U138 (N_138,In_139,In_862);
nand U139 (N_139,In_423,In_642);
nand U140 (N_140,In_37,In_936);
xnor U141 (N_141,In_1127,In_248);
or U142 (N_142,In_1457,In_705);
nor U143 (N_143,In_834,In_1254);
or U144 (N_144,In_546,In_934);
nor U145 (N_145,In_1315,In_1331);
nor U146 (N_146,In_1492,In_97);
and U147 (N_147,In_990,In_1337);
and U148 (N_148,In_186,In_476);
xnor U149 (N_149,In_1017,In_1393);
xor U150 (N_150,In_531,In_784);
nor U151 (N_151,In_217,In_770);
nand U152 (N_152,In_1040,In_1287);
or U153 (N_153,In_1161,In_930);
nor U154 (N_154,In_855,In_512);
xor U155 (N_155,In_1212,In_345);
nor U156 (N_156,In_844,In_744);
xor U157 (N_157,In_554,In_767);
nand U158 (N_158,In_325,In_728);
nand U159 (N_159,In_902,In_1273);
nor U160 (N_160,In_17,In_835);
or U161 (N_161,In_1486,In_939);
or U162 (N_162,In_249,In_1409);
or U163 (N_163,In_1048,In_130);
xor U164 (N_164,In_1362,In_411);
nand U165 (N_165,In_913,In_876);
xnor U166 (N_166,In_237,In_874);
nor U167 (N_167,In_196,In_160);
nand U168 (N_168,In_562,In_730);
nand U169 (N_169,In_363,In_570);
or U170 (N_170,In_843,In_527);
nor U171 (N_171,In_827,In_643);
nor U172 (N_172,In_967,In_731);
or U173 (N_173,In_727,In_1099);
and U174 (N_174,In_1133,In_961);
or U175 (N_175,In_591,In_714);
xnor U176 (N_176,In_1075,In_397);
nand U177 (N_177,In_156,In_853);
or U178 (N_178,In_451,In_219);
xor U179 (N_179,In_655,In_315);
xor U180 (N_180,In_178,In_909);
nor U181 (N_181,In_375,In_838);
or U182 (N_182,In_295,In_707);
nor U183 (N_183,In_188,In_14);
and U184 (N_184,In_791,In_373);
or U185 (N_185,In_713,In_310);
and U186 (N_186,In_850,In_182);
xnor U187 (N_187,In_511,In_318);
xnor U188 (N_188,In_1152,In_1299);
xor U189 (N_189,In_149,In_1396);
or U190 (N_190,In_479,In_65);
and U191 (N_191,In_1147,In_1288);
nand U192 (N_192,In_879,In_132);
nor U193 (N_193,In_659,In_1357);
nand U194 (N_194,In_1317,In_782);
and U195 (N_195,In_1330,In_230);
and U196 (N_196,In_472,In_560);
or U197 (N_197,In_802,In_674);
nor U198 (N_198,In_1329,In_191);
and U199 (N_199,In_739,In_750);
or U200 (N_200,In_975,In_319);
nor U201 (N_201,In_382,In_444);
and U202 (N_202,In_1487,In_1069);
nand U203 (N_203,In_929,In_664);
xor U204 (N_204,In_392,In_1206);
nor U205 (N_205,In_1039,In_1046);
nand U206 (N_206,In_228,In_841);
nand U207 (N_207,In_1424,In_0);
nand U208 (N_208,In_180,In_362);
xnor U209 (N_209,In_424,In_1417);
and U210 (N_210,In_1464,In_916);
and U211 (N_211,In_1103,In_743);
or U212 (N_212,In_1225,In_999);
nand U213 (N_213,In_421,In_172);
or U214 (N_214,In_322,In_443);
nor U215 (N_215,In_1029,In_535);
or U216 (N_216,In_95,In_367);
and U217 (N_217,In_385,In_108);
xor U218 (N_218,In_358,In_434);
or U219 (N_219,In_159,In_1418);
or U220 (N_220,In_670,In_1110);
xor U221 (N_221,In_342,In_523);
nand U222 (N_222,In_854,In_691);
nand U223 (N_223,In_865,In_1345);
xnor U224 (N_224,In_815,In_328);
and U225 (N_225,In_922,In_425);
nand U226 (N_226,In_729,In_826);
xor U227 (N_227,In_43,In_412);
nor U228 (N_228,In_682,In_1192);
nand U229 (N_229,In_175,In_1411);
xor U230 (N_230,In_516,In_901);
xor U231 (N_231,In_1452,In_49);
nand U232 (N_232,In_437,In_515);
xor U233 (N_233,In_278,In_881);
nand U234 (N_234,In_1002,In_458);
nand U235 (N_235,In_1164,In_858);
xnor U236 (N_236,In_304,In_1257);
nor U237 (N_237,In_471,In_287);
nand U238 (N_238,In_1483,In_915);
and U239 (N_239,In_1172,In_1148);
nor U240 (N_240,In_1460,In_1265);
nor U241 (N_241,In_138,In_675);
and U242 (N_242,In_953,In_568);
nand U243 (N_243,In_72,In_786);
nand U244 (N_244,In_845,In_1294);
or U245 (N_245,In_1334,In_107);
xnor U246 (N_246,In_1232,In_100);
xnor U247 (N_247,In_290,In_1442);
nor U248 (N_248,In_384,In_244);
nor U249 (N_249,In_610,In_1414);
and U250 (N_250,In_1416,N_207);
or U251 (N_251,N_205,In_1382);
xnor U252 (N_252,N_241,In_445);
xor U253 (N_253,In_1422,In_882);
nand U254 (N_254,In_492,N_147);
and U255 (N_255,In_109,In_1066);
nor U256 (N_256,In_150,In_985);
nand U257 (N_257,In_131,In_320);
or U258 (N_258,In_1134,In_544);
nor U259 (N_259,N_146,In_1061);
and U260 (N_260,In_1240,In_507);
and U261 (N_261,In_960,In_579);
xor U262 (N_262,In_1484,N_230);
nor U263 (N_263,In_101,In_353);
nand U264 (N_264,In_1246,In_169);
xor U265 (N_265,In_946,N_176);
xnor U266 (N_266,In_615,N_29);
xnor U267 (N_267,In_415,In_298);
and U268 (N_268,In_259,In_904);
or U269 (N_269,In_1307,In_504);
and U270 (N_270,N_24,In_154);
or U271 (N_271,In_616,In_10);
nor U272 (N_272,In_1353,In_1377);
or U273 (N_273,In_557,In_211);
or U274 (N_274,In_828,In_793);
nor U275 (N_275,N_119,In_848);
or U276 (N_276,N_13,In_537);
xor U277 (N_277,In_1243,In_202);
or U278 (N_278,N_156,In_806);
nor U279 (N_279,In_1455,In_1428);
nor U280 (N_280,In_1187,N_79);
and U281 (N_281,In_1182,In_1356);
xor U282 (N_282,N_142,In_1200);
or U283 (N_283,In_403,In_141);
xor U284 (N_284,In_1151,In_1434);
and U285 (N_285,In_1176,In_407);
and U286 (N_286,In_801,In_972);
nor U287 (N_287,In_15,N_60);
xor U288 (N_288,In_571,In_1419);
and U289 (N_289,N_170,N_178);
or U290 (N_290,N_68,In_1250);
nand U291 (N_291,In_1224,In_137);
nand U292 (N_292,In_678,N_93);
nand U293 (N_293,N_231,N_94);
nor U294 (N_294,In_59,In_1031);
nor U295 (N_295,N_150,In_1358);
and U296 (N_296,In_1346,In_654);
nor U297 (N_297,N_51,In_595);
nor U298 (N_298,In_177,N_228);
xor U299 (N_299,In_663,In_117);
nand U300 (N_300,In_1449,In_433);
nor U301 (N_301,In_1494,In_1333);
nand U302 (N_302,In_816,N_35);
or U303 (N_303,In_24,In_1085);
or U304 (N_304,In_1453,In_536);
nor U305 (N_305,In_47,In_955);
nand U306 (N_306,In_63,In_34);
or U307 (N_307,In_777,In_80);
xnor U308 (N_308,In_326,In_121);
or U309 (N_309,In_1383,In_632);
nand U310 (N_310,In_306,In_1415);
xnor U311 (N_311,In_1162,In_1261);
nand U312 (N_312,In_1421,N_57);
nor U313 (N_313,In_905,In_416);
and U314 (N_314,In_868,In_847);
nor U315 (N_315,In_419,In_371);
nor U316 (N_316,In_1427,In_481);
nor U317 (N_317,In_1044,N_118);
xor U318 (N_318,In_253,In_840);
nand U319 (N_319,N_126,In_272);
and U320 (N_320,N_26,N_41);
nand U321 (N_321,In_1006,In_534);
nand U322 (N_322,In_622,In_1482);
or U323 (N_323,N_220,In_77);
nor U324 (N_324,In_760,In_578);
and U325 (N_325,In_619,In_1430);
nand U326 (N_326,In_1480,In_144);
nor U327 (N_327,In_1098,In_647);
and U328 (N_328,In_940,In_822);
xor U329 (N_329,In_265,In_1074);
nand U330 (N_330,In_361,N_227);
nand U331 (N_331,In_402,In_300);
nand U332 (N_332,In_932,In_645);
or U333 (N_333,N_100,In_1130);
xor U334 (N_334,In_1293,In_575);
xor U335 (N_335,In_1210,In_773);
xor U336 (N_336,In_31,In_526);
xor U337 (N_337,In_183,In_737);
and U338 (N_338,N_20,N_203);
nor U339 (N_339,N_243,In_606);
xnor U340 (N_340,In_948,In_1367);
xor U341 (N_341,N_185,N_28);
and U342 (N_342,In_908,In_474);
nor U343 (N_343,In_1096,In_532);
nand U344 (N_344,In_70,In_759);
nand U345 (N_345,N_56,In_1435);
or U346 (N_346,In_613,In_635);
xor U347 (N_347,N_96,In_1471);
nor U348 (N_348,In_508,N_183);
nand U349 (N_349,In_1033,In_824);
or U350 (N_350,In_331,N_85);
nor U351 (N_351,N_22,In_859);
and U352 (N_352,In_398,N_171);
or U353 (N_353,N_65,In_1336);
and U354 (N_354,In_956,In_621);
nor U355 (N_355,In_273,In_482);
nand U356 (N_356,In_725,N_87);
and U357 (N_357,In_1191,In_1328);
or U358 (N_358,In_733,In_216);
nor U359 (N_359,N_86,In_1245);
xnor U360 (N_360,In_1173,In_1045);
nor U361 (N_361,N_131,N_111);
nand U362 (N_362,N_120,In_798);
nand U363 (N_363,In_1498,N_152);
nand U364 (N_364,In_224,In_1115);
nand U365 (N_365,In_565,In_628);
xor U366 (N_366,N_90,In_1499);
and U367 (N_367,In_1009,In_125);
and U368 (N_368,In_120,N_102);
nand U369 (N_369,In_514,In_831);
xor U370 (N_370,In_1466,In_1070);
or U371 (N_371,In_323,In_6);
or U372 (N_372,In_1379,In_435);
and U373 (N_373,In_491,In_477);
nand U374 (N_374,In_1082,In_870);
and U375 (N_375,In_1403,N_158);
xnor U376 (N_376,N_247,In_764);
or U377 (N_377,In_558,In_266);
xnor U378 (N_378,In_992,In_406);
nor U379 (N_379,In_388,In_521);
nand U380 (N_380,In_333,In_528);
or U381 (N_381,N_214,In_350);
nand U382 (N_382,N_181,N_0);
nand U383 (N_383,N_154,N_62);
xor U384 (N_384,In_819,In_312);
xor U385 (N_385,In_1107,In_335);
or U386 (N_386,N_219,N_188);
xnor U387 (N_387,N_91,In_1189);
xor U388 (N_388,In_1041,N_222);
nor U389 (N_389,In_998,In_846);
and U390 (N_390,In_703,In_1063);
xor U391 (N_391,In_860,N_58);
and U392 (N_392,In_1112,In_82);
nor U393 (N_393,In_339,In_85);
nor U394 (N_394,In_762,N_139);
nor U395 (N_395,In_116,In_1489);
and U396 (N_396,In_830,In_1135);
or U397 (N_397,In_1310,In_1429);
or U398 (N_398,In_935,In_1186);
nand U399 (N_399,In_1404,In_899);
or U400 (N_400,In_646,In_530);
and U401 (N_401,In_204,In_23);
or U402 (N_402,In_1248,In_1497);
and U403 (N_403,N_161,In_1062);
and U404 (N_404,N_225,In_969);
nor U405 (N_405,In_753,In_311);
and U406 (N_406,In_1157,In_50);
or U407 (N_407,In_292,In_994);
or U408 (N_408,In_199,In_656);
xor U409 (N_409,In_1153,In_1426);
nor U410 (N_410,N_217,In_399);
or U411 (N_411,In_262,In_455);
and U412 (N_412,In_349,In_1363);
xnor U413 (N_413,In_661,In_1217);
nand U414 (N_414,In_856,N_36);
nand U415 (N_415,In_1222,In_709);
xnor U416 (N_416,In_321,In_1229);
and U417 (N_417,In_381,In_213);
or U418 (N_418,In_952,In_1476);
and U419 (N_419,In_324,In_404);
nor U420 (N_420,In_200,N_2);
and U421 (N_421,N_10,In_1472);
xor U422 (N_422,N_101,In_924);
nor U423 (N_423,In_1496,N_21);
or U424 (N_424,In_1374,In_470);
nor U425 (N_425,In_783,In_667);
nor U426 (N_426,N_18,N_106);
nor U427 (N_427,In_489,In_699);
xor U428 (N_428,N_133,N_59);
or U429 (N_429,In_151,In_1118);
nor U430 (N_430,In_1413,In_1231);
xor U431 (N_431,In_389,N_70);
and U432 (N_432,In_757,In_1234);
and U433 (N_433,N_244,In_420);
or U434 (N_434,In_227,N_12);
and U435 (N_435,In_1433,In_716);
or U436 (N_436,In_712,In_1431);
and U437 (N_437,In_722,In_888);
and U438 (N_438,In_1106,In_1068);
and U439 (N_439,In_73,N_140);
nor U440 (N_440,In_57,In_1251);
nor U441 (N_441,In_8,N_103);
or U442 (N_442,In_282,N_78);
nand U443 (N_443,In_710,In_147);
or U444 (N_444,In_1477,In_55);
nor U445 (N_445,In_1121,In_280);
nand U446 (N_446,In_440,In_58);
nor U447 (N_447,In_1020,In_114);
nand U448 (N_448,In_1026,In_1032);
xor U449 (N_449,In_677,N_55);
nor U450 (N_450,In_567,In_1101);
nand U451 (N_451,In_69,In_222);
or U452 (N_452,In_1055,In_1291);
nand U453 (N_453,N_135,In_1169);
xor U454 (N_454,N_160,In_605);
nand U455 (N_455,In_539,In_1338);
xnor U456 (N_456,N_155,In_396);
or U457 (N_457,In_66,In_765);
nand U458 (N_458,In_1117,In_1102);
and U459 (N_459,In_741,In_1301);
xor U460 (N_460,In_517,In_463);
xnor U461 (N_461,In_181,In_780);
nand U462 (N_462,In_653,In_708);
xor U463 (N_463,In_48,N_149);
and U464 (N_464,In_81,In_7);
and U465 (N_465,N_84,In_1004);
nor U466 (N_466,In_274,In_1351);
and U467 (N_467,In_299,In_1126);
xnor U468 (N_468,N_184,In_1120);
and U469 (N_469,In_254,In_1057);
and U470 (N_470,In_94,In_209);
nor U471 (N_471,In_1077,N_136);
nor U472 (N_472,N_166,In_238);
nor U473 (N_473,In_1154,In_861);
nand U474 (N_474,In_194,N_8);
or U475 (N_475,In_973,In_197);
and U476 (N_476,In_592,In_1059);
nand U477 (N_477,In_745,In_928);
nor U478 (N_478,In_136,In_623);
nor U479 (N_479,In_1084,N_107);
and U480 (N_480,In_1235,In_639);
or U481 (N_481,In_92,In_658);
and U482 (N_482,In_1332,In_1348);
and U483 (N_483,In_51,N_248);
nor U484 (N_484,N_71,In_820);
and U485 (N_485,In_1019,In_33);
nor U486 (N_486,In_852,In_545);
xor U487 (N_487,In_450,N_27);
xnor U488 (N_488,N_211,N_99);
xor U489 (N_489,In_501,In_978);
xor U490 (N_490,N_141,In_787);
nand U491 (N_491,In_790,In_942);
and U492 (N_492,In_192,In_93);
xnor U493 (N_493,In_987,N_123);
nand U494 (N_494,In_296,In_538);
nand U495 (N_495,In_696,In_688);
or U496 (N_496,In_480,In_809);
nand U497 (N_497,N_53,In_462);
and U498 (N_498,In_1241,In_617);
nor U499 (N_499,In_984,N_235);
and U500 (N_500,In_803,In_309);
nor U501 (N_501,In_884,In_651);
nand U502 (N_502,In_1104,In_1282);
nor U503 (N_503,N_208,In_752);
nand U504 (N_504,In_1129,In_965);
xnor U505 (N_505,In_261,N_432);
xor U506 (N_506,N_306,N_232);
or U507 (N_507,In_933,N_484);
nor U508 (N_508,N_48,In_1108);
and U509 (N_509,In_556,In_1086);
nor U510 (N_510,N_467,N_359);
nor U511 (N_511,In_1021,In_457);
nand U512 (N_512,In_811,N_404);
xor U513 (N_513,In_205,In_781);
xnor U514 (N_514,In_638,In_673);
xor U515 (N_515,N_462,N_399);
nand U516 (N_516,N_237,N_421);
and U517 (N_517,In_755,N_288);
or U518 (N_518,N_76,In_962);
and U519 (N_519,In_162,In_1223);
nor U520 (N_520,N_312,In_155);
or U521 (N_521,N_393,In_1325);
nor U522 (N_522,In_851,N_448);
or U523 (N_523,N_173,N_67);
xor U524 (N_524,In_400,N_290);
and U525 (N_525,N_381,In_785);
or U526 (N_526,N_309,In_1423);
nor U527 (N_527,N_296,N_145);
and U528 (N_528,In_1311,In_499);
nand U529 (N_529,In_1456,N_5);
and U530 (N_530,N_481,N_471);
and U531 (N_531,In_586,N_256);
xor U532 (N_532,In_13,In_1014);
and U533 (N_533,In_842,In_1372);
or U534 (N_534,N_356,N_77);
and U535 (N_535,N_271,In_548);
and U536 (N_536,N_425,N_43);
or U537 (N_537,In_308,N_199);
and U538 (N_538,In_839,In_1355);
or U539 (N_539,N_320,In_1050);
nand U540 (N_540,In_44,In_566);
and U541 (N_541,In_903,N_114);
and U542 (N_542,In_1475,In_468);
or U543 (N_543,In_161,In_1072);
nand U544 (N_544,In_717,In_721);
nand U545 (N_545,In_630,In_821);
nor U546 (N_546,In_1131,In_104);
xor U547 (N_547,N_283,In_695);
or U548 (N_548,In_1035,In_1286);
xnor U549 (N_549,In_1193,In_800);
nand U550 (N_550,In_46,In_1136);
or U551 (N_551,In_1140,In_896);
nor U552 (N_552,In_260,N_451);
and U553 (N_553,In_1125,In_409);
xnor U554 (N_554,N_423,N_485);
and U555 (N_555,In_475,In_1196);
or U556 (N_556,N_117,In_167);
or U557 (N_557,N_483,In_799);
and U558 (N_558,In_1205,N_303);
and U559 (N_559,N_479,In_1347);
xnor U560 (N_560,In_812,N_264);
nor U561 (N_561,N_206,N_74);
or U562 (N_562,In_919,N_162);
nor U563 (N_563,N_349,N_213);
xor U564 (N_564,In_1384,In_634);
and U565 (N_565,In_1385,In_1028);
nor U566 (N_566,In_1473,N_165);
nand U567 (N_567,In_778,In_541);
nand U568 (N_568,N_115,N_229);
xnor U569 (N_569,N_493,N_72);
nand U570 (N_570,N_352,In_993);
xnor U571 (N_571,In_460,N_439);
and U572 (N_572,In_581,In_810);
xor U573 (N_573,In_56,In_465);
nand U574 (N_574,In_553,N_191);
xnor U575 (N_575,N_454,N_478);
nand U576 (N_576,N_435,N_322);
nor U577 (N_577,In_453,In_1281);
or U578 (N_578,N_417,In_906);
and U579 (N_579,In_1214,In_430);
and U580 (N_580,In_122,In_1407);
and U581 (N_581,N_371,N_44);
nand U582 (N_582,In_317,In_379);
nand U583 (N_583,N_365,N_3);
nand U584 (N_584,In_631,N_195);
or U585 (N_585,In_1034,N_169);
nor U586 (N_586,In_341,In_16);
or U587 (N_587,N_50,N_212);
and U588 (N_588,In_1474,In_1037);
nor U589 (N_589,In_660,N_105);
or U590 (N_590,In_5,N_382);
or U591 (N_591,In_949,In_1324);
nand U592 (N_592,In_486,N_148);
xnor U593 (N_593,In_355,In_1233);
and U594 (N_594,N_457,N_186);
and U595 (N_595,In_796,In_143);
or U596 (N_596,In_1469,In_817);
and U597 (N_597,In_386,In_68);
xor U598 (N_598,In_1071,N_285);
nand U599 (N_599,N_438,In_518);
or U600 (N_600,In_614,In_21);
or U601 (N_601,In_1270,N_440);
nor U602 (N_602,N_487,N_238);
nand U603 (N_603,In_376,N_446);
and U604 (N_604,In_1298,N_298);
nor U605 (N_605,In_221,N_325);
nand U606 (N_606,In_1285,In_693);
or U607 (N_607,In_1067,In_185);
nor U608 (N_608,N_318,N_326);
nor U609 (N_609,N_476,In_380);
and U610 (N_610,In_1247,In_442);
or U611 (N_611,In_1113,N_11);
xor U612 (N_612,In_1079,In_542);
xor U613 (N_613,In_1354,In_1137);
or U614 (N_614,N_19,In_165);
and U615 (N_615,N_144,N_204);
and U616 (N_616,In_849,N_1);
xor U617 (N_617,In_1111,N_128);
nand U618 (N_618,N_151,N_308);
xnor U619 (N_619,N_347,In_1027);
nor U620 (N_620,In_1008,N_299);
nor U621 (N_621,N_127,N_321);
xnor U622 (N_622,In_410,N_384);
nor U623 (N_623,In_148,In_1051);
nor U624 (N_624,In_795,In_669);
and U625 (N_625,N_374,In_246);
nand U626 (N_626,In_1412,In_833);
or U627 (N_627,N_268,N_402);
xnor U628 (N_628,In_686,N_202);
nor U629 (N_629,N_258,N_323);
and U630 (N_630,In_12,N_474);
and U631 (N_631,In_1252,In_163);
and U632 (N_632,N_267,N_338);
and U633 (N_633,In_464,In_103);
and U634 (N_634,N_98,In_390);
nand U635 (N_635,In_1454,N_431);
and U636 (N_636,In_1339,In_334);
nand U637 (N_637,In_797,In_684);
nor U638 (N_638,In_957,N_469);
or U639 (N_639,In_887,In_1047);
nand U640 (N_640,N_282,In_598);
nand U641 (N_641,In_1221,In_589);
or U642 (N_642,In_52,In_996);
and U643 (N_643,In_1174,N_427);
xnor U644 (N_644,N_63,In_478);
and U645 (N_645,N_346,N_66);
xor U646 (N_646,N_234,In_1209);
nand U647 (N_647,In_1220,In_1083);
nand U648 (N_648,In_427,N_354);
nand U649 (N_649,In_1364,N_433);
nor U650 (N_650,In_637,In_28);
or U651 (N_651,In_1279,N_366);
xor U652 (N_652,In_1387,N_104);
and U653 (N_653,N_249,In_947);
xnor U654 (N_654,N_276,In_338);
and U655 (N_655,In_1448,In_1090);
and U656 (N_656,In_1141,In_897);
xor U657 (N_657,In_1300,N_112);
nor U658 (N_658,N_486,In_979);
or U659 (N_659,In_683,N_443);
and U660 (N_660,In_1297,In_1175);
nor U661 (N_661,In_364,In_467);
xor U662 (N_662,N_167,N_341);
xnor U663 (N_663,In_176,N_121);
nor U664 (N_664,N_460,In_665);
nor U665 (N_665,N_302,In_283);
and U666 (N_666,N_426,In_340);
xnor U667 (N_667,In_1160,In_1095);
or U668 (N_668,In_348,In_88);
xor U669 (N_669,N_429,In_891);
nor U670 (N_670,N_293,In_1266);
or U671 (N_671,In_873,In_938);
nand U672 (N_672,N_116,In_269);
nand U673 (N_673,N_464,In_119);
xor U674 (N_674,N_109,In_40);
and U675 (N_675,N_345,N_31);
or U676 (N_676,N_69,N_215);
and U677 (N_677,In_775,N_442);
xnor U678 (N_678,N_122,In_438);
nor U679 (N_679,N_34,In_36);
or U680 (N_680,In_633,N_348);
nor U681 (N_681,N_329,In_704);
nand U682 (N_682,N_239,In_878);
nor U683 (N_683,In_954,N_193);
and U684 (N_684,N_40,N_180);
and U685 (N_685,In_604,N_450);
and U686 (N_686,In_1478,In_808);
xnor U687 (N_687,In_529,N_251);
nand U688 (N_688,N_47,N_378);
nor U689 (N_689,N_319,In_503);
nor U690 (N_690,In_356,N_465);
or U691 (N_691,In_1401,N_373);
nor U692 (N_692,In_555,N_16);
xnor U693 (N_693,N_130,N_436);
nand U694 (N_694,N_380,In_911);
and U695 (N_695,N_459,N_23);
nand U696 (N_696,In_907,In_618);
nor U697 (N_697,In_174,In_383);
xnor U698 (N_698,N_344,In_255);
nor U699 (N_699,N_38,In_871);
nor U700 (N_700,In_487,In_365);
and U701 (N_701,N_108,In_1344);
or U702 (N_702,In_1438,In_1488);
and U703 (N_703,N_278,In_29);
and U704 (N_704,N_88,In_234);
or U705 (N_705,N_333,N_377);
nand U706 (N_706,N_447,N_250);
and U707 (N_707,N_406,In_724);
nand U708 (N_708,In_1078,In_212);
nor U709 (N_709,N_492,N_7);
and U710 (N_710,N_335,In_87);
nand U711 (N_711,In_1420,In_1000);
nor U712 (N_712,N_407,N_82);
nand U713 (N_713,N_89,In_1);
xnor U714 (N_714,In_146,In_1446);
xnor U715 (N_715,In_189,N_233);
xnor U716 (N_716,N_9,In_576);
nor U717 (N_717,N_192,In_776);
xnor U718 (N_718,In_96,In_681);
and U719 (N_719,In_607,N_274);
nand U720 (N_720,In_42,In_20);
nor U721 (N_721,N_375,In_454);
or U722 (N_722,In_524,In_629);
and U723 (N_723,In_1341,In_600);
and U724 (N_724,In_1459,N_75);
nor U725 (N_725,In_45,N_390);
nor U726 (N_726,N_386,In_241);
and U727 (N_727,In_593,In_366);
nand U728 (N_728,In_1327,In_662);
xnor U729 (N_729,In_330,N_209);
xor U730 (N_730,N_125,In_1227);
nor U731 (N_731,In_1342,In_872);
and U732 (N_732,N_263,N_339);
xnor U733 (N_733,N_301,N_200);
and U734 (N_734,N_242,N_279);
nor U735 (N_735,In_1036,In_687);
nor U736 (N_736,In_1138,In_594);
and U737 (N_737,In_981,In_1058);
xnor U738 (N_738,N_189,In_1052);
nor U739 (N_739,In_1349,In_689);
or U740 (N_740,In_1340,In_640);
nand U741 (N_741,In_1259,In_1395);
nor U742 (N_742,In_289,In_964);
and U743 (N_743,N_281,In_1208);
nor U744 (N_744,In_585,N_414);
nor U745 (N_745,In_86,N_472);
or U746 (N_746,N_434,N_64);
xnor U747 (N_747,In_285,In_1155);
and U748 (N_748,In_1380,In_429);
xor U749 (N_749,In_513,In_201);
xnor U750 (N_750,N_661,N_275);
and U751 (N_751,N_505,N_674);
or U752 (N_752,N_387,N_453);
xnor U753 (N_753,N_332,N_670);
nor U754 (N_754,N_580,In_275);
and U755 (N_755,In_1018,In_549);
nor U756 (N_756,In_1461,In_774);
xnor U757 (N_757,In_1481,In_679);
and U758 (N_758,N_337,N_664);
nand U759 (N_759,In_1149,N_685);
and U760 (N_760,In_203,In_286);
xnor U761 (N_761,N_681,N_260);
xor U762 (N_762,In_1366,In_723);
nor U763 (N_763,In_734,In_432);
or U764 (N_764,In_140,N_182);
or U765 (N_765,N_675,N_292);
nand U766 (N_766,N_546,N_177);
or U767 (N_767,N_360,N_662);
nor U768 (N_768,N_697,N_273);
nor U769 (N_769,N_695,N_223);
nand U770 (N_770,In_19,In_1237);
or U771 (N_771,N_372,In_1166);
xor U772 (N_772,N_124,N_196);
or U773 (N_773,N_668,N_590);
and U774 (N_774,In_483,N_642);
nand U775 (N_775,In_720,N_718);
xnor U776 (N_776,N_596,N_413);
nand U777 (N_777,In_313,In_1013);
nand U778 (N_778,N_527,In_1398);
nand U779 (N_779,In_1406,N_284);
or U780 (N_780,In_126,N_515);
nand U781 (N_781,In_79,N_514);
nor U782 (N_782,N_691,N_54);
nor U783 (N_783,In_1180,N_143);
or U784 (N_784,In_701,In_1043);
or U785 (N_785,In_1025,In_1089);
or U786 (N_786,N_400,N_530);
nor U787 (N_787,N_683,In_112);
or U788 (N_788,In_583,N_621);
or U789 (N_789,N_327,N_52);
nand U790 (N_790,N_466,N_497);
xnor U791 (N_791,N_437,N_617);
nor U792 (N_792,N_401,N_584);
xnor U793 (N_793,In_374,In_644);
xnor U794 (N_794,N_653,In_921);
nor U795 (N_795,In_1168,N_595);
and U796 (N_796,N_536,In_62);
or U797 (N_797,N_672,In_127);
xnor U798 (N_798,In_1012,N_194);
xor U799 (N_799,In_700,N_571);
xnor U800 (N_800,In_657,N_490);
nand U801 (N_801,N_576,In_336);
nand U802 (N_802,In_168,In_719);
and U803 (N_803,In_268,N_30);
and U804 (N_804,In_1105,N_640);
nand U805 (N_805,N_502,N_179);
and U806 (N_806,N_575,N_747);
xnor U807 (N_807,In_966,N_741);
nand U808 (N_808,N_286,In_1195);
or U809 (N_809,N_369,N_644);
nand U810 (N_810,In_1312,N_313);
and U811 (N_811,N_686,In_426);
xor U812 (N_812,N_579,N_245);
nand U813 (N_813,In_864,In_577);
or U814 (N_814,N_594,N_509);
xnor U815 (N_815,N_508,N_690);
or U816 (N_816,In_1064,In_256);
nor U817 (N_817,N_395,In_1100);
or U818 (N_818,In_923,In_193);
or U819 (N_819,N_428,In_1087);
nor U820 (N_820,N_523,N_592);
xnor U821 (N_821,N_604,N_164);
xnor U822 (N_822,N_396,In_257);
xor U823 (N_823,In_1410,In_863);
or U824 (N_824,N_328,N_562);
nand U825 (N_825,In_431,In_958);
nor U826 (N_826,N_455,In_636);
xor U827 (N_827,In_1361,N_743);
and U828 (N_828,N_295,N_733);
and U829 (N_829,In_983,In_1213);
or U830 (N_830,N_616,N_444);
nor U831 (N_831,In_587,N_37);
or U832 (N_832,N_506,N_236);
xnor U833 (N_833,N_641,N_376);
nand U834 (N_834,N_618,N_602);
or U835 (N_835,N_539,N_168);
xor U836 (N_836,In_395,N_706);
nand U837 (N_837,N_370,N_629);
and U838 (N_838,N_615,N_518);
xor U839 (N_839,N_627,N_39);
or U840 (N_840,In_452,N_628);
xnor U841 (N_841,In_680,N_463);
or U842 (N_842,In_1088,N_702);
xnor U843 (N_843,N_409,In_1437);
nor U844 (N_844,N_277,In_1278);
xor U845 (N_845,In_792,N_529);
xor U846 (N_846,N_666,N_398);
xor U847 (N_847,In_405,In_943);
or U848 (N_848,N_651,N_216);
or U849 (N_849,N_408,N_315);
and U850 (N_850,In_469,N_737);
nand U851 (N_851,N_367,In_267);
nor U852 (N_852,In_944,N_555);
nand U853 (N_853,In_649,In_950);
nand U854 (N_854,N_353,N_613);
xor U855 (N_855,N_291,In_229);
or U856 (N_856,N_415,N_533);
or U857 (N_857,In_917,N_684);
or U858 (N_858,In_1290,N_699);
nand U859 (N_859,N_532,In_337);
nor U860 (N_860,In_1493,N_707);
nand U861 (N_861,N_416,N_726);
or U862 (N_862,N_727,In_98);
nand U863 (N_863,In_1081,N_605);
xor U864 (N_864,In_898,N_468);
nand U865 (N_865,In_569,N_620);
nand U866 (N_866,In_738,N_673);
or U867 (N_867,N_42,N_45);
xnor U868 (N_868,N_520,N_569);
nor U869 (N_869,N_714,N_389);
or U870 (N_870,N_588,In_436);
or U871 (N_871,In_1145,N_449);
xnor U872 (N_872,In_294,N_494);
nand U873 (N_873,N_418,In_1402);
nand U874 (N_874,N_495,In_1065);
or U875 (N_875,In_184,N_740);
nor U876 (N_876,In_1194,N_224);
xnor U877 (N_877,In_1439,N_15);
and U878 (N_878,N_607,In_768);
or U879 (N_879,N_97,In_235);
xor U880 (N_880,In_233,In_1170);
or U881 (N_881,N_624,N_526);
xor U882 (N_882,N_570,In_1292);
or U883 (N_883,N_175,In_264);
or U884 (N_884,N_92,In_1343);
or U885 (N_885,In_590,In_1177);
nor U886 (N_886,N_657,N_132);
xor U887 (N_887,In_551,N_547);
nand U888 (N_888,N_512,N_324);
nand U889 (N_889,N_300,N_541);
nor U890 (N_890,N_157,In_1091);
xnor U891 (N_891,In_243,N_259);
or U892 (N_892,N_197,N_358);
nor U893 (N_893,In_1470,N_33);
and U894 (N_894,In_601,N_713);
or U895 (N_895,N_262,N_410);
nor U896 (N_896,N_261,N_174);
or U897 (N_897,In_754,In_829);
nand U898 (N_898,In_1495,N_420);
or U899 (N_899,In_359,In_698);
or U900 (N_900,N_637,In_789);
nand U901 (N_901,N_383,N_491);
or U902 (N_902,In_1056,N_716);
or U903 (N_903,N_379,In_1381);
xnor U904 (N_904,N_330,N_163);
xor U905 (N_905,N_456,N_310);
or U906 (N_906,N_210,In_494);
and U907 (N_907,In_1268,N_477);
or U908 (N_908,N_599,In_239);
nor U909 (N_909,N_659,N_679);
and U910 (N_910,In_54,N_500);
xor U911 (N_911,N_110,In_885);
nor U912 (N_912,In_22,In_522);
or U913 (N_913,In_1001,In_1386);
nor U914 (N_914,N_687,N_734);
or U915 (N_915,N_565,N_357);
nor U916 (N_916,N_287,N_542);
nand U917 (N_917,In_620,N_680);
nand U918 (N_918,N_452,N_445);
and U919 (N_919,N_671,N_631);
xor U920 (N_920,In_974,N_696);
or U921 (N_921,N_458,N_622);
xor U922 (N_922,N_504,N_645);
nand U923 (N_923,In_1405,N_531);
nor U924 (N_924,N_566,N_265);
and U925 (N_925,N_461,In_648);
xor U926 (N_926,N_589,In_35);
xor U927 (N_927,In_357,In_1373);
nand U928 (N_928,N_488,N_559);
nor U929 (N_929,N_568,In_490);
or U930 (N_930,N_655,In_1303);
nor U931 (N_931,N_711,In_1123);
nor U932 (N_932,In_1440,N_660);
nand U933 (N_933,In_625,In_769);
nand U934 (N_934,In_1392,N_350);
nand U935 (N_935,In_1238,In_1122);
xnor U936 (N_936,In_1264,In_297);
xnor U937 (N_937,N_676,In_9);
nor U938 (N_938,In_414,N_138);
xor U939 (N_939,N_688,In_1323);
xor U940 (N_940,N_201,In_1451);
and U941 (N_941,In_1280,In_118);
and U942 (N_942,N_257,In_742);
or U943 (N_943,N_609,N_81);
nor U944 (N_944,In_164,N_709);
and U945 (N_945,N_610,N_693);
nor U946 (N_946,In_1239,In_71);
and U947 (N_947,N_730,N_650);
xnor U948 (N_948,N_581,N_503);
and U949 (N_949,N_665,N_639);
xnor U950 (N_950,In_543,N_403);
or U951 (N_951,In_1365,In_671);
or U952 (N_952,In_110,In_1184);
nor U953 (N_953,In_417,In_393);
nor U954 (N_954,N_397,In_1304);
nor U955 (N_955,In_547,In_588);
nor U956 (N_956,N_722,N_270);
and U957 (N_957,N_652,N_95);
xor U958 (N_958,In_1262,N_704);
nand U959 (N_959,N_316,In_133);
and U960 (N_960,In_327,In_343);
or U961 (N_961,N_545,N_6);
or U962 (N_962,N_742,N_317);
or U963 (N_963,N_725,N_412);
nand U964 (N_964,In_74,N_475);
nand U965 (N_965,In_968,N_489);
or U966 (N_966,In_75,N_705);
nor U967 (N_967,N_535,N_521);
nand U968 (N_968,In_89,In_550);
nor U969 (N_969,N_698,N_305);
nand U970 (N_970,N_654,N_424);
and U971 (N_971,N_46,N_507);
nand U972 (N_972,N_614,In_495);
nor U973 (N_973,In_771,N_331);
nor U974 (N_974,N_510,N_744);
or U975 (N_975,N_619,In_1436);
xor U976 (N_976,N_611,In_1179);
nor U977 (N_977,N_113,In_1165);
or U978 (N_978,In_1024,N_538);
or U979 (N_979,In_1408,N_717);
and U980 (N_980,In_694,In_30);
or U981 (N_981,In_187,In_1289);
and U982 (N_982,N_362,In_401);
nor U983 (N_983,N_511,N_626);
or U984 (N_984,N_351,N_269);
or U985 (N_985,N_551,N_544);
and U986 (N_986,In_910,In_208);
and U987 (N_987,In_1360,N_534);
and U988 (N_988,In_305,In_597);
xor U989 (N_989,N_388,N_405);
nor U990 (N_990,N_501,In_179);
nand U991 (N_991,N_643,N_636);
or U992 (N_992,In_27,N_297);
or U993 (N_993,N_561,N_630);
nor U994 (N_994,N_633,N_391);
nor U995 (N_995,In_893,N_255);
and U996 (N_996,N_658,N_625);
nor U997 (N_997,N_603,N_710);
or U998 (N_998,N_669,In_564);
or U999 (N_999,N_392,In_685);
xor U1000 (N_1000,N_899,N_480);
nand U1001 (N_1001,N_656,N_612);
nand U1002 (N_1002,N_870,N_582);
or U1003 (N_1003,N_554,N_779);
nand U1004 (N_1004,In_1073,N_826);
and U1005 (N_1005,N_955,In_866);
and U1006 (N_1006,N_788,N_731);
nand U1007 (N_1007,N_938,N_549);
nor U1008 (N_1008,In_1450,N_947);
xnor U1009 (N_1009,N_915,N_363);
nand U1010 (N_1010,N_159,N_187);
or U1011 (N_1011,N_762,N_519);
or U1012 (N_1012,In_1202,N_969);
nand U1013 (N_1013,In_980,N_809);
nor U1014 (N_1014,In_25,N_825);
nor U1015 (N_1015,N_851,In_959);
nor U1016 (N_1016,In_276,N_982);
nor U1017 (N_1017,N_935,N_820);
xnor U1018 (N_1018,N_844,N_364);
or U1019 (N_1019,N_951,N_865);
nor U1020 (N_1020,In_650,N_422);
or U1021 (N_1021,N_782,N_597);
nor U1022 (N_1022,In_976,N_824);
xor U1023 (N_1023,N_990,N_962);
nand U1024 (N_1024,N_829,N_897);
nand U1025 (N_1025,In_102,N_49);
or U1026 (N_1026,N_560,N_226);
or U1027 (N_1027,N_723,N_758);
or U1028 (N_1028,N_606,In_552);
nor U1029 (N_1029,N_516,N_266);
or U1030 (N_1030,N_995,N_783);
xnor U1031 (N_1031,N_701,N_781);
xor U1032 (N_1032,N_868,In_497);
nor U1033 (N_1033,N_941,N_394);
and U1034 (N_1034,In_608,N_355);
nor U1035 (N_1035,N_797,N_792);
xnor U1036 (N_1036,N_739,N_874);
or U1037 (N_1037,In_718,N_736);
xnor U1038 (N_1038,N_803,N_866);
and U1039 (N_1039,N_756,N_932);
or U1040 (N_1040,N_957,N_905);
and U1041 (N_1041,In_746,N_837);
or U1042 (N_1042,N_522,N_473);
and U1043 (N_1043,In_360,N_419);
nor U1044 (N_1044,N_996,N_921);
xnor U1045 (N_1045,N_891,N_766);
nand U1046 (N_1046,In_215,N_895);
xor U1047 (N_1047,N_877,In_1114);
nand U1048 (N_1048,In_1188,N_850);
nand U1049 (N_1049,In_1204,N_912);
xnor U1050 (N_1050,In_1003,In_158);
and U1051 (N_1051,N_540,N_61);
or U1052 (N_1052,N_931,N_774);
nor U1053 (N_1053,In_448,N_920);
nand U1054 (N_1054,N_361,In_749);
nor U1055 (N_1055,N_967,In_1190);
nand U1056 (N_1056,N_901,N_908);
xnor U1057 (N_1057,N_720,N_153);
nand U1058 (N_1058,N_719,In_1306);
nand U1059 (N_1059,N_735,N_913);
nand U1060 (N_1060,N_909,N_838);
or U1061 (N_1061,N_14,N_849);
or U1062 (N_1062,N_875,In_1388);
xor U1063 (N_1063,N_583,N_635);
xor U1064 (N_1064,In_1119,N_761);
or U1065 (N_1065,N_172,N_751);
nor U1066 (N_1066,N_757,N_985);
nand U1067 (N_1067,N_928,In_1042);
nand U1068 (N_1068,In_1296,N_942);
xor U1069 (N_1069,N_854,N_971);
and U1070 (N_1070,N_198,N_896);
or U1071 (N_1071,N_304,N_598);
xnor U1072 (N_1072,In_1022,N_648);
and U1073 (N_1073,N_649,N_25);
nor U1074 (N_1074,N_855,N_703);
or U1075 (N_1075,N_772,N_773);
and U1076 (N_1076,N_903,N_787);
nor U1077 (N_1077,N_712,N_600);
nand U1078 (N_1078,N_916,In_26);
nand U1079 (N_1079,N_80,In_461);
nand U1080 (N_1080,In_603,In_611);
or U1081 (N_1081,N_548,N_944);
nand U1082 (N_1082,N_853,N_822);
or U1083 (N_1083,In_1468,N_917);
or U1084 (N_1084,In_726,N_927);
or U1085 (N_1085,N_801,N_632);
nand U1086 (N_1086,N_933,N_470);
nand U1087 (N_1087,N_368,N_775);
xnor U1088 (N_1088,In_447,N_989);
or U1089 (N_1089,N_795,N_754);
or U1090 (N_1090,In_1319,In_1397);
nand U1091 (N_1091,N_663,N_949);
nor U1092 (N_1092,N_988,N_799);
or U1093 (N_1093,N_567,N_898);
xor U1094 (N_1094,N_943,N_922);
and U1095 (N_1095,N_623,In_84);
and U1096 (N_1096,In_672,N_914);
or U1097 (N_1097,N_812,N_252);
xnor U1098 (N_1098,In_1228,N_860);
nor U1099 (N_1099,N_983,In_157);
nand U1100 (N_1100,N_482,In_877);
xnor U1101 (N_1101,N_700,N_959);
nand U1102 (N_1102,N_946,N_558);
nand U1103 (N_1103,N_190,N_73);
or U1104 (N_1104,N_970,N_498);
and U1105 (N_1105,In_1283,N_577);
nor U1106 (N_1106,N_790,N_246);
and U1107 (N_1107,N_694,N_889);
or U1108 (N_1108,N_963,In_951);
nor U1109 (N_1109,In_937,N_524);
or U1110 (N_1110,In_291,N_647);
nor U1111 (N_1111,N_134,N_441);
nand U1112 (N_1112,N_593,N_738);
or U1113 (N_1113,N_776,In_520);
or U1114 (N_1114,N_980,N_682);
nand U1115 (N_1115,N_768,In_641);
nand U1116 (N_1116,In_525,In_1371);
and U1117 (N_1117,In_892,N_667);
nand U1118 (N_1118,N_843,N_385);
or U1119 (N_1119,N_311,N_608);
nand U1120 (N_1120,N_586,N_819);
and U1121 (N_1121,N_32,N_221);
and U1122 (N_1122,N_828,N_430);
or U1123 (N_1123,N_834,N_879);
nand U1124 (N_1124,In_1447,N_998);
nand U1125 (N_1125,N_882,N_770);
and U1126 (N_1126,N_975,N_755);
nand U1127 (N_1127,N_981,In_1158);
or U1128 (N_1128,N_563,N_954);
or U1129 (N_1129,N_748,N_930);
or U1130 (N_1130,In_372,N_767);
xnor U1131 (N_1131,N_883,N_574);
nor U1132 (N_1132,N_517,N_815);
xor U1133 (N_1133,N_972,N_794);
and U1134 (N_1134,N_878,N_808);
xnor U1135 (N_1135,N_796,N_553);
nor U1136 (N_1136,N_752,N_968);
and U1137 (N_1137,N_557,In_456);
nor U1138 (N_1138,In_1218,N_862);
nand U1139 (N_1139,N_918,N_272);
or U1140 (N_1140,N_777,N_902);
nand U1141 (N_1141,N_689,N_678);
nor U1142 (N_1142,In_1199,In_1335);
xor U1143 (N_1143,N_585,In_995);
xnor U1144 (N_1144,N_564,N_218);
or U1145 (N_1145,N_858,N_17);
or U1146 (N_1146,N_552,N_994);
and U1147 (N_1147,N_923,In_195);
nor U1148 (N_1148,In_1178,In_1318);
xnor U1149 (N_1149,N_786,N_827);
and U1150 (N_1150,In_1479,N_893);
or U1151 (N_1151,In_626,N_769);
nand U1152 (N_1152,In_971,N_840);
xor U1153 (N_1153,N_342,N_806);
or U1154 (N_1154,N_869,N_280);
nand U1155 (N_1155,In_1139,N_894);
nand U1156 (N_1156,N_802,N_867);
xor U1157 (N_1157,In_1267,N_784);
nor U1158 (N_1158,N_992,N_817);
xnor U1159 (N_1159,In_1010,N_811);
or U1160 (N_1160,N_960,N_785);
and U1161 (N_1161,N_572,N_993);
nor U1162 (N_1162,In_706,In_38);
xnor U1163 (N_1163,N_578,N_646);
nand U1164 (N_1164,N_979,N_692);
nand U1165 (N_1165,In_1326,In_1441);
and U1166 (N_1166,N_953,N_496);
nand U1167 (N_1167,N_289,N_925);
and U1168 (N_1168,N_852,N_746);
nand U1169 (N_1169,N_892,N_778);
nand U1170 (N_1170,N_876,N_842);
nor U1171 (N_1171,N_638,In_78);
or U1172 (N_1172,N_499,In_1313);
xor U1173 (N_1173,N_771,N_724);
or U1174 (N_1174,N_810,N_888);
and U1175 (N_1175,N_984,N_750);
nor U1176 (N_1176,N_871,N_715);
and U1177 (N_1177,N_861,N_728);
and U1178 (N_1178,N_856,N_818);
xnor U1179 (N_1179,In_240,N_924);
or U1180 (N_1180,N_831,N_550);
xor U1181 (N_1181,N_753,In_1219);
nor U1182 (N_1182,In_668,N_591);
or U1183 (N_1183,N_936,N_823);
or U1184 (N_1184,N_997,N_587);
and U1185 (N_1185,N_978,N_847);
xnor U1186 (N_1186,N_800,N_987);
nor U1187 (N_1187,In_18,N_765);
or U1188 (N_1188,N_846,N_340);
and U1189 (N_1189,N_745,In_711);
nand U1190 (N_1190,N_961,N_904);
xor U1191 (N_1191,N_872,N_816);
or U1192 (N_1192,N_859,N_343);
or U1193 (N_1193,In_1275,N_934);
xor U1194 (N_1194,In_3,N_965);
nor U1195 (N_1195,In_53,N_708);
or U1196 (N_1196,N_863,N_814);
nor U1197 (N_1197,N_793,N_830);
nor U1198 (N_1198,N_845,N_759);
xnor U1199 (N_1199,N_910,N_4);
and U1200 (N_1200,N_907,N_881);
nand U1201 (N_1201,N_841,In_880);
and U1202 (N_1202,N_839,N_805);
or U1203 (N_1203,N_254,N_832);
xor U1204 (N_1204,In_912,N_977);
xor U1205 (N_1205,N_253,N_528);
xor U1206 (N_1206,N_974,N_807);
and U1207 (N_1207,N_857,N_886);
nand U1208 (N_1208,N_732,N_900);
xnor U1209 (N_1209,N_864,N_129);
nand U1210 (N_1210,In_270,N_780);
nand U1211 (N_1211,In_314,In_1183);
nor U1212 (N_1212,N_940,N_890);
and U1213 (N_1213,N_945,N_721);
and U1214 (N_1214,N_986,N_833);
nand U1215 (N_1215,N_911,In_41);
nor U1216 (N_1216,N_926,N_791);
or U1217 (N_1217,N_789,N_763);
or U1218 (N_1218,N_513,N_760);
and U1219 (N_1219,N_543,In_145);
or U1220 (N_1220,N_973,N_573);
xor U1221 (N_1221,N_749,In_857);
and U1222 (N_1222,N_835,N_556);
nor U1223 (N_1223,In_963,N_729);
xor U1224 (N_1224,N_634,N_956);
or U1225 (N_1225,N_601,In_142);
nand U1226 (N_1226,N_999,N_240);
nor U1227 (N_1227,N_887,N_948);
or U1228 (N_1228,N_939,N_976);
xnor U1229 (N_1229,N_950,N_314);
nand U1230 (N_1230,N_336,In_90);
nor U1231 (N_1231,In_64,N_764);
nor U1232 (N_1232,N_919,N_880);
nand U1233 (N_1233,N_952,N_929);
and U1234 (N_1234,In_418,In_105);
and U1235 (N_1235,N_137,In_1226);
xnor U1236 (N_1236,N_958,N_525);
and U1237 (N_1237,N_885,In_488);
xor U1238 (N_1238,N_884,N_836);
xnor U1239 (N_1239,N_966,N_873);
nor U1240 (N_1240,In_1201,N_937);
and U1241 (N_1241,N_411,N_848);
or U1242 (N_1242,N_83,N_677);
or U1243 (N_1243,In_533,N_991);
and U1244 (N_1244,N_294,N_798);
nor U1245 (N_1245,N_804,N_964);
or U1246 (N_1246,N_813,In_413);
or U1247 (N_1247,N_906,N_537);
xnor U1248 (N_1248,N_821,N_334);
nor U1249 (N_1249,N_307,In_247);
nand U1250 (N_1250,N_1248,N_1229);
and U1251 (N_1251,N_1218,N_1152);
or U1252 (N_1252,N_1214,N_1038);
nand U1253 (N_1253,N_1025,N_1132);
and U1254 (N_1254,N_1070,N_1130);
nor U1255 (N_1255,N_1180,N_1129);
or U1256 (N_1256,N_1193,N_1029);
nand U1257 (N_1257,N_1014,N_1222);
xnor U1258 (N_1258,N_1153,N_1237);
nor U1259 (N_1259,N_1177,N_1047);
xor U1260 (N_1260,N_1035,N_1210);
and U1261 (N_1261,N_1186,N_1164);
nor U1262 (N_1262,N_1023,N_1046);
and U1263 (N_1263,N_1149,N_1227);
xor U1264 (N_1264,N_1206,N_1207);
nand U1265 (N_1265,N_1127,N_1201);
nor U1266 (N_1266,N_1240,N_1109);
and U1267 (N_1267,N_1044,N_1169);
and U1268 (N_1268,N_1054,N_1209);
nor U1269 (N_1269,N_1083,N_1133);
nor U1270 (N_1270,N_1112,N_1000);
nor U1271 (N_1271,N_1002,N_1092);
or U1272 (N_1272,N_1102,N_1148);
or U1273 (N_1273,N_1233,N_1163);
nor U1274 (N_1274,N_1062,N_1121);
nor U1275 (N_1275,N_1188,N_1232);
and U1276 (N_1276,N_1008,N_1236);
nor U1277 (N_1277,N_1042,N_1151);
or U1278 (N_1278,N_1128,N_1137);
xor U1279 (N_1279,N_1077,N_1215);
or U1280 (N_1280,N_1199,N_1108);
nand U1281 (N_1281,N_1067,N_1024);
nor U1282 (N_1282,N_1093,N_1058);
or U1283 (N_1283,N_1018,N_1141);
or U1284 (N_1284,N_1099,N_1150);
or U1285 (N_1285,N_1145,N_1053);
nand U1286 (N_1286,N_1016,N_1195);
and U1287 (N_1287,N_1175,N_1246);
and U1288 (N_1288,N_1106,N_1079);
or U1289 (N_1289,N_1087,N_1080);
or U1290 (N_1290,N_1005,N_1213);
and U1291 (N_1291,N_1073,N_1049);
and U1292 (N_1292,N_1006,N_1168);
nor U1293 (N_1293,N_1146,N_1198);
or U1294 (N_1294,N_1172,N_1007);
or U1295 (N_1295,N_1069,N_1082);
xnor U1296 (N_1296,N_1212,N_1182);
and U1297 (N_1297,N_1096,N_1174);
nor U1298 (N_1298,N_1004,N_1230);
nand U1299 (N_1299,N_1244,N_1140);
nand U1300 (N_1300,N_1001,N_1032);
nor U1301 (N_1301,N_1239,N_1245);
nor U1302 (N_1302,N_1139,N_1187);
and U1303 (N_1303,N_1157,N_1134);
and U1304 (N_1304,N_1131,N_1166);
nor U1305 (N_1305,N_1097,N_1194);
or U1306 (N_1306,N_1089,N_1235);
and U1307 (N_1307,N_1221,N_1011);
and U1308 (N_1308,N_1040,N_1033);
xnor U1309 (N_1309,N_1015,N_1242);
or U1310 (N_1310,N_1124,N_1105);
xor U1311 (N_1311,N_1185,N_1111);
and U1312 (N_1312,N_1101,N_1078);
and U1313 (N_1313,N_1165,N_1211);
or U1314 (N_1314,N_1113,N_1216);
and U1315 (N_1315,N_1068,N_1071);
nor U1316 (N_1316,N_1100,N_1200);
xnor U1317 (N_1317,N_1027,N_1085);
nand U1318 (N_1318,N_1118,N_1039);
nor U1319 (N_1319,N_1051,N_1138);
and U1320 (N_1320,N_1190,N_1116);
nand U1321 (N_1321,N_1136,N_1143);
xor U1322 (N_1322,N_1017,N_1013);
xnor U1323 (N_1323,N_1159,N_1224);
or U1324 (N_1324,N_1022,N_1158);
nor U1325 (N_1325,N_1061,N_1126);
nor U1326 (N_1326,N_1037,N_1135);
and U1327 (N_1327,N_1205,N_1088);
or U1328 (N_1328,N_1203,N_1104);
xor U1329 (N_1329,N_1228,N_1019);
nor U1330 (N_1330,N_1090,N_1156);
nor U1331 (N_1331,N_1197,N_1110);
nor U1332 (N_1332,N_1026,N_1010);
xor U1333 (N_1333,N_1050,N_1220);
xor U1334 (N_1334,N_1120,N_1231);
nand U1335 (N_1335,N_1030,N_1036);
xor U1336 (N_1336,N_1147,N_1041);
nor U1337 (N_1337,N_1249,N_1107);
nand U1338 (N_1338,N_1217,N_1155);
nor U1339 (N_1339,N_1184,N_1119);
nand U1340 (N_1340,N_1055,N_1167);
xor U1341 (N_1341,N_1066,N_1192);
or U1342 (N_1342,N_1219,N_1065);
nor U1343 (N_1343,N_1064,N_1142);
or U1344 (N_1344,N_1202,N_1238);
or U1345 (N_1345,N_1204,N_1021);
nor U1346 (N_1346,N_1115,N_1226);
nor U1347 (N_1347,N_1074,N_1176);
nor U1348 (N_1348,N_1103,N_1098);
nor U1349 (N_1349,N_1048,N_1243);
or U1350 (N_1350,N_1063,N_1012);
or U1351 (N_1351,N_1084,N_1171);
nor U1352 (N_1352,N_1170,N_1034);
nor U1353 (N_1353,N_1114,N_1003);
xnor U1354 (N_1354,N_1162,N_1052);
and U1355 (N_1355,N_1056,N_1072);
and U1356 (N_1356,N_1043,N_1091);
or U1357 (N_1357,N_1179,N_1045);
xnor U1358 (N_1358,N_1060,N_1086);
nor U1359 (N_1359,N_1076,N_1161);
xor U1360 (N_1360,N_1009,N_1123);
nor U1361 (N_1361,N_1247,N_1081);
or U1362 (N_1362,N_1223,N_1057);
xnor U1363 (N_1363,N_1183,N_1189);
nor U1364 (N_1364,N_1178,N_1095);
and U1365 (N_1365,N_1208,N_1160);
nor U1366 (N_1366,N_1191,N_1075);
or U1367 (N_1367,N_1122,N_1196);
xnor U1368 (N_1368,N_1154,N_1225);
and U1369 (N_1369,N_1028,N_1173);
or U1370 (N_1370,N_1020,N_1031);
nor U1371 (N_1371,N_1117,N_1125);
xor U1372 (N_1372,N_1144,N_1059);
nor U1373 (N_1373,N_1094,N_1241);
xnor U1374 (N_1374,N_1181,N_1234);
and U1375 (N_1375,N_1150,N_1170);
nand U1376 (N_1376,N_1121,N_1161);
xnor U1377 (N_1377,N_1032,N_1228);
nor U1378 (N_1378,N_1142,N_1184);
xor U1379 (N_1379,N_1146,N_1230);
nor U1380 (N_1380,N_1203,N_1108);
xnor U1381 (N_1381,N_1188,N_1011);
nand U1382 (N_1382,N_1094,N_1028);
and U1383 (N_1383,N_1125,N_1113);
nand U1384 (N_1384,N_1025,N_1153);
nand U1385 (N_1385,N_1212,N_1102);
or U1386 (N_1386,N_1044,N_1087);
nor U1387 (N_1387,N_1090,N_1045);
nor U1388 (N_1388,N_1032,N_1222);
and U1389 (N_1389,N_1212,N_1040);
nand U1390 (N_1390,N_1077,N_1134);
xnor U1391 (N_1391,N_1059,N_1062);
xnor U1392 (N_1392,N_1031,N_1032);
xor U1393 (N_1393,N_1000,N_1162);
nor U1394 (N_1394,N_1217,N_1215);
nand U1395 (N_1395,N_1246,N_1104);
nor U1396 (N_1396,N_1042,N_1136);
xnor U1397 (N_1397,N_1068,N_1063);
nand U1398 (N_1398,N_1103,N_1085);
xnor U1399 (N_1399,N_1011,N_1133);
or U1400 (N_1400,N_1111,N_1053);
or U1401 (N_1401,N_1090,N_1185);
xnor U1402 (N_1402,N_1141,N_1166);
and U1403 (N_1403,N_1190,N_1186);
or U1404 (N_1404,N_1161,N_1242);
nand U1405 (N_1405,N_1076,N_1036);
and U1406 (N_1406,N_1090,N_1231);
nand U1407 (N_1407,N_1052,N_1218);
or U1408 (N_1408,N_1080,N_1093);
and U1409 (N_1409,N_1229,N_1201);
and U1410 (N_1410,N_1030,N_1249);
nor U1411 (N_1411,N_1061,N_1070);
nor U1412 (N_1412,N_1179,N_1088);
or U1413 (N_1413,N_1058,N_1202);
xor U1414 (N_1414,N_1091,N_1086);
xor U1415 (N_1415,N_1061,N_1118);
nand U1416 (N_1416,N_1194,N_1013);
and U1417 (N_1417,N_1017,N_1200);
or U1418 (N_1418,N_1075,N_1152);
or U1419 (N_1419,N_1028,N_1022);
xor U1420 (N_1420,N_1184,N_1077);
and U1421 (N_1421,N_1077,N_1145);
nor U1422 (N_1422,N_1174,N_1162);
and U1423 (N_1423,N_1018,N_1068);
nor U1424 (N_1424,N_1105,N_1008);
nand U1425 (N_1425,N_1216,N_1172);
nor U1426 (N_1426,N_1173,N_1179);
nor U1427 (N_1427,N_1186,N_1139);
nor U1428 (N_1428,N_1167,N_1163);
or U1429 (N_1429,N_1055,N_1064);
xnor U1430 (N_1430,N_1141,N_1198);
xnor U1431 (N_1431,N_1037,N_1234);
or U1432 (N_1432,N_1248,N_1179);
nand U1433 (N_1433,N_1152,N_1044);
and U1434 (N_1434,N_1152,N_1146);
xnor U1435 (N_1435,N_1080,N_1060);
and U1436 (N_1436,N_1059,N_1156);
nand U1437 (N_1437,N_1000,N_1233);
nand U1438 (N_1438,N_1236,N_1084);
and U1439 (N_1439,N_1040,N_1139);
nor U1440 (N_1440,N_1135,N_1036);
nor U1441 (N_1441,N_1070,N_1092);
or U1442 (N_1442,N_1155,N_1005);
nor U1443 (N_1443,N_1097,N_1106);
nand U1444 (N_1444,N_1003,N_1138);
and U1445 (N_1445,N_1026,N_1152);
nor U1446 (N_1446,N_1009,N_1118);
nor U1447 (N_1447,N_1126,N_1073);
xnor U1448 (N_1448,N_1028,N_1016);
nor U1449 (N_1449,N_1020,N_1199);
xor U1450 (N_1450,N_1186,N_1044);
nand U1451 (N_1451,N_1175,N_1055);
nor U1452 (N_1452,N_1231,N_1042);
nor U1453 (N_1453,N_1029,N_1212);
or U1454 (N_1454,N_1056,N_1203);
or U1455 (N_1455,N_1211,N_1215);
nand U1456 (N_1456,N_1219,N_1008);
or U1457 (N_1457,N_1151,N_1247);
or U1458 (N_1458,N_1030,N_1020);
nor U1459 (N_1459,N_1028,N_1197);
and U1460 (N_1460,N_1025,N_1076);
xnor U1461 (N_1461,N_1211,N_1060);
xor U1462 (N_1462,N_1024,N_1134);
xor U1463 (N_1463,N_1133,N_1196);
nand U1464 (N_1464,N_1099,N_1190);
xnor U1465 (N_1465,N_1133,N_1053);
or U1466 (N_1466,N_1249,N_1181);
xor U1467 (N_1467,N_1094,N_1044);
nor U1468 (N_1468,N_1218,N_1204);
or U1469 (N_1469,N_1159,N_1137);
and U1470 (N_1470,N_1112,N_1223);
nor U1471 (N_1471,N_1147,N_1152);
xor U1472 (N_1472,N_1067,N_1159);
or U1473 (N_1473,N_1183,N_1044);
and U1474 (N_1474,N_1058,N_1246);
and U1475 (N_1475,N_1148,N_1208);
or U1476 (N_1476,N_1131,N_1223);
nor U1477 (N_1477,N_1230,N_1137);
nor U1478 (N_1478,N_1040,N_1246);
nand U1479 (N_1479,N_1097,N_1214);
and U1480 (N_1480,N_1129,N_1114);
nor U1481 (N_1481,N_1031,N_1024);
and U1482 (N_1482,N_1100,N_1114);
nor U1483 (N_1483,N_1173,N_1016);
or U1484 (N_1484,N_1080,N_1085);
or U1485 (N_1485,N_1209,N_1125);
xnor U1486 (N_1486,N_1183,N_1088);
nor U1487 (N_1487,N_1157,N_1168);
or U1488 (N_1488,N_1079,N_1103);
nand U1489 (N_1489,N_1154,N_1176);
nor U1490 (N_1490,N_1205,N_1238);
nor U1491 (N_1491,N_1198,N_1186);
nand U1492 (N_1492,N_1147,N_1013);
nand U1493 (N_1493,N_1081,N_1166);
nor U1494 (N_1494,N_1077,N_1216);
nor U1495 (N_1495,N_1154,N_1184);
nand U1496 (N_1496,N_1102,N_1161);
nand U1497 (N_1497,N_1159,N_1107);
xnor U1498 (N_1498,N_1002,N_1124);
nand U1499 (N_1499,N_1230,N_1091);
nor U1500 (N_1500,N_1429,N_1489);
nor U1501 (N_1501,N_1348,N_1441);
nor U1502 (N_1502,N_1405,N_1303);
xnor U1503 (N_1503,N_1326,N_1327);
and U1504 (N_1504,N_1490,N_1262);
and U1505 (N_1505,N_1382,N_1274);
and U1506 (N_1506,N_1428,N_1250);
xor U1507 (N_1507,N_1313,N_1469);
xor U1508 (N_1508,N_1440,N_1307);
or U1509 (N_1509,N_1390,N_1496);
nor U1510 (N_1510,N_1318,N_1331);
nand U1511 (N_1511,N_1290,N_1450);
nor U1512 (N_1512,N_1254,N_1251);
xor U1513 (N_1513,N_1430,N_1386);
and U1514 (N_1514,N_1477,N_1314);
xnor U1515 (N_1515,N_1433,N_1470);
and U1516 (N_1516,N_1361,N_1462);
and U1517 (N_1517,N_1264,N_1445);
nor U1518 (N_1518,N_1420,N_1465);
nor U1519 (N_1519,N_1474,N_1360);
xnor U1520 (N_1520,N_1292,N_1442);
nand U1521 (N_1521,N_1404,N_1350);
xor U1522 (N_1522,N_1460,N_1367);
and U1523 (N_1523,N_1328,N_1396);
or U1524 (N_1524,N_1362,N_1392);
and U1525 (N_1525,N_1457,N_1286);
xnor U1526 (N_1526,N_1497,N_1342);
nor U1527 (N_1527,N_1495,N_1463);
or U1528 (N_1528,N_1373,N_1426);
and U1529 (N_1529,N_1330,N_1446);
xor U1530 (N_1530,N_1343,N_1352);
nor U1531 (N_1531,N_1260,N_1322);
xnor U1532 (N_1532,N_1376,N_1395);
nor U1533 (N_1533,N_1434,N_1493);
nand U1534 (N_1534,N_1499,N_1273);
xnor U1535 (N_1535,N_1263,N_1271);
xor U1536 (N_1536,N_1458,N_1443);
nor U1537 (N_1537,N_1280,N_1391);
nand U1538 (N_1538,N_1431,N_1275);
nand U1539 (N_1539,N_1349,N_1380);
or U1540 (N_1540,N_1436,N_1482);
xnor U1541 (N_1541,N_1253,N_1291);
or U1542 (N_1542,N_1265,N_1488);
and U1543 (N_1543,N_1425,N_1401);
xor U1544 (N_1544,N_1410,N_1494);
nor U1545 (N_1545,N_1485,N_1289);
nor U1546 (N_1546,N_1277,N_1379);
xor U1547 (N_1547,N_1288,N_1483);
nand U1548 (N_1548,N_1365,N_1407);
nor U1549 (N_1549,N_1296,N_1298);
nor U1550 (N_1550,N_1339,N_1356);
nor U1551 (N_1551,N_1403,N_1359);
nand U1552 (N_1552,N_1370,N_1484);
or U1553 (N_1553,N_1269,N_1408);
and U1554 (N_1554,N_1284,N_1372);
and U1555 (N_1555,N_1475,N_1293);
nand U1556 (N_1556,N_1294,N_1419);
nor U1557 (N_1557,N_1398,N_1416);
nor U1558 (N_1558,N_1498,N_1451);
or U1559 (N_1559,N_1304,N_1325);
nor U1560 (N_1560,N_1389,N_1335);
nor U1561 (N_1561,N_1492,N_1385);
xor U1562 (N_1562,N_1406,N_1347);
or U1563 (N_1563,N_1388,N_1472);
nor U1564 (N_1564,N_1479,N_1423);
or U1565 (N_1565,N_1368,N_1394);
or U1566 (N_1566,N_1444,N_1378);
and U1567 (N_1567,N_1334,N_1299);
nand U1568 (N_1568,N_1256,N_1259);
or U1569 (N_1569,N_1383,N_1267);
nand U1570 (N_1570,N_1438,N_1305);
and U1571 (N_1571,N_1437,N_1351);
nor U1572 (N_1572,N_1261,N_1413);
or U1573 (N_1573,N_1338,N_1272);
nand U1574 (N_1574,N_1336,N_1308);
and U1575 (N_1575,N_1309,N_1355);
nor U1576 (N_1576,N_1480,N_1266);
nand U1577 (N_1577,N_1455,N_1393);
nand U1578 (N_1578,N_1366,N_1473);
xor U1579 (N_1579,N_1375,N_1302);
nor U1580 (N_1580,N_1315,N_1464);
or U1581 (N_1581,N_1358,N_1345);
or U1582 (N_1582,N_1258,N_1397);
or U1583 (N_1583,N_1461,N_1279);
and U1584 (N_1584,N_1377,N_1468);
nand U1585 (N_1585,N_1487,N_1449);
nand U1586 (N_1586,N_1417,N_1287);
and U1587 (N_1587,N_1387,N_1456);
nor U1588 (N_1588,N_1297,N_1424);
or U1589 (N_1589,N_1317,N_1270);
nor U1590 (N_1590,N_1276,N_1301);
xnor U1591 (N_1591,N_1459,N_1337);
and U1592 (N_1592,N_1412,N_1283);
nand U1593 (N_1593,N_1422,N_1316);
nand U1594 (N_1594,N_1471,N_1306);
and U1595 (N_1595,N_1402,N_1491);
and U1596 (N_1596,N_1415,N_1252);
xor U1597 (N_1597,N_1300,N_1369);
nor U1598 (N_1598,N_1255,N_1374);
nor U1599 (N_1599,N_1323,N_1363);
xnor U1600 (N_1600,N_1353,N_1371);
nand U1601 (N_1601,N_1467,N_1400);
nand U1602 (N_1602,N_1295,N_1344);
nor U1603 (N_1603,N_1281,N_1448);
and U1604 (N_1604,N_1320,N_1354);
and U1605 (N_1605,N_1357,N_1332);
and U1606 (N_1606,N_1414,N_1409);
and U1607 (N_1607,N_1340,N_1321);
or U1608 (N_1608,N_1435,N_1411);
nor U1609 (N_1609,N_1329,N_1452);
and U1610 (N_1610,N_1418,N_1399);
nor U1611 (N_1611,N_1285,N_1333);
xor U1612 (N_1612,N_1476,N_1384);
xor U1613 (N_1613,N_1346,N_1432);
xor U1614 (N_1614,N_1282,N_1278);
nor U1615 (N_1615,N_1324,N_1439);
and U1616 (N_1616,N_1312,N_1310);
xnor U1617 (N_1617,N_1311,N_1257);
nor U1618 (N_1618,N_1364,N_1478);
or U1619 (N_1619,N_1454,N_1268);
nor U1620 (N_1620,N_1486,N_1481);
nand U1621 (N_1621,N_1319,N_1466);
and U1622 (N_1622,N_1447,N_1453);
nor U1623 (N_1623,N_1427,N_1421);
and U1624 (N_1624,N_1381,N_1341);
and U1625 (N_1625,N_1475,N_1433);
xnor U1626 (N_1626,N_1397,N_1322);
or U1627 (N_1627,N_1355,N_1299);
and U1628 (N_1628,N_1428,N_1419);
nand U1629 (N_1629,N_1434,N_1308);
nand U1630 (N_1630,N_1441,N_1375);
and U1631 (N_1631,N_1483,N_1361);
nor U1632 (N_1632,N_1323,N_1297);
nand U1633 (N_1633,N_1464,N_1469);
xor U1634 (N_1634,N_1309,N_1392);
nand U1635 (N_1635,N_1377,N_1476);
nor U1636 (N_1636,N_1388,N_1383);
nor U1637 (N_1637,N_1306,N_1272);
xnor U1638 (N_1638,N_1440,N_1454);
nor U1639 (N_1639,N_1315,N_1444);
or U1640 (N_1640,N_1323,N_1423);
or U1641 (N_1641,N_1372,N_1317);
xor U1642 (N_1642,N_1433,N_1357);
or U1643 (N_1643,N_1290,N_1312);
nor U1644 (N_1644,N_1387,N_1330);
xnor U1645 (N_1645,N_1296,N_1433);
or U1646 (N_1646,N_1492,N_1286);
nand U1647 (N_1647,N_1275,N_1276);
xnor U1648 (N_1648,N_1368,N_1364);
or U1649 (N_1649,N_1473,N_1306);
nor U1650 (N_1650,N_1398,N_1456);
or U1651 (N_1651,N_1262,N_1427);
nand U1652 (N_1652,N_1254,N_1416);
nor U1653 (N_1653,N_1271,N_1342);
and U1654 (N_1654,N_1453,N_1284);
xor U1655 (N_1655,N_1460,N_1451);
nor U1656 (N_1656,N_1364,N_1299);
xnor U1657 (N_1657,N_1410,N_1294);
and U1658 (N_1658,N_1473,N_1328);
and U1659 (N_1659,N_1377,N_1471);
xnor U1660 (N_1660,N_1440,N_1350);
or U1661 (N_1661,N_1391,N_1460);
nor U1662 (N_1662,N_1278,N_1468);
xor U1663 (N_1663,N_1491,N_1319);
nand U1664 (N_1664,N_1286,N_1392);
xor U1665 (N_1665,N_1265,N_1453);
xor U1666 (N_1666,N_1403,N_1300);
xor U1667 (N_1667,N_1420,N_1411);
or U1668 (N_1668,N_1385,N_1291);
nor U1669 (N_1669,N_1426,N_1353);
and U1670 (N_1670,N_1421,N_1428);
nor U1671 (N_1671,N_1264,N_1352);
nand U1672 (N_1672,N_1393,N_1288);
nor U1673 (N_1673,N_1422,N_1437);
nor U1674 (N_1674,N_1302,N_1258);
or U1675 (N_1675,N_1284,N_1496);
nand U1676 (N_1676,N_1252,N_1294);
and U1677 (N_1677,N_1377,N_1338);
xnor U1678 (N_1678,N_1498,N_1287);
and U1679 (N_1679,N_1311,N_1252);
nand U1680 (N_1680,N_1265,N_1418);
nor U1681 (N_1681,N_1307,N_1302);
and U1682 (N_1682,N_1320,N_1460);
and U1683 (N_1683,N_1253,N_1440);
nor U1684 (N_1684,N_1486,N_1373);
xor U1685 (N_1685,N_1461,N_1415);
nor U1686 (N_1686,N_1473,N_1337);
nor U1687 (N_1687,N_1259,N_1346);
xnor U1688 (N_1688,N_1257,N_1376);
nor U1689 (N_1689,N_1425,N_1468);
and U1690 (N_1690,N_1335,N_1364);
and U1691 (N_1691,N_1421,N_1269);
or U1692 (N_1692,N_1484,N_1300);
nand U1693 (N_1693,N_1253,N_1323);
xor U1694 (N_1694,N_1475,N_1429);
and U1695 (N_1695,N_1406,N_1304);
or U1696 (N_1696,N_1295,N_1448);
xor U1697 (N_1697,N_1320,N_1400);
xor U1698 (N_1698,N_1439,N_1474);
xnor U1699 (N_1699,N_1385,N_1275);
or U1700 (N_1700,N_1327,N_1370);
and U1701 (N_1701,N_1396,N_1353);
or U1702 (N_1702,N_1487,N_1321);
and U1703 (N_1703,N_1468,N_1443);
nand U1704 (N_1704,N_1401,N_1488);
or U1705 (N_1705,N_1322,N_1495);
nand U1706 (N_1706,N_1455,N_1422);
and U1707 (N_1707,N_1435,N_1366);
xnor U1708 (N_1708,N_1309,N_1296);
or U1709 (N_1709,N_1251,N_1268);
or U1710 (N_1710,N_1408,N_1379);
and U1711 (N_1711,N_1476,N_1338);
or U1712 (N_1712,N_1469,N_1479);
nor U1713 (N_1713,N_1433,N_1314);
xnor U1714 (N_1714,N_1446,N_1343);
and U1715 (N_1715,N_1414,N_1426);
nand U1716 (N_1716,N_1291,N_1339);
xor U1717 (N_1717,N_1378,N_1261);
and U1718 (N_1718,N_1495,N_1420);
or U1719 (N_1719,N_1294,N_1292);
or U1720 (N_1720,N_1364,N_1265);
and U1721 (N_1721,N_1390,N_1354);
xnor U1722 (N_1722,N_1440,N_1442);
xor U1723 (N_1723,N_1372,N_1422);
xnor U1724 (N_1724,N_1251,N_1278);
nand U1725 (N_1725,N_1318,N_1484);
xnor U1726 (N_1726,N_1307,N_1468);
nor U1727 (N_1727,N_1418,N_1331);
nand U1728 (N_1728,N_1252,N_1291);
nor U1729 (N_1729,N_1447,N_1353);
or U1730 (N_1730,N_1354,N_1449);
nand U1731 (N_1731,N_1408,N_1354);
nor U1732 (N_1732,N_1490,N_1405);
xnor U1733 (N_1733,N_1250,N_1266);
and U1734 (N_1734,N_1411,N_1302);
nor U1735 (N_1735,N_1257,N_1252);
nand U1736 (N_1736,N_1344,N_1409);
xor U1737 (N_1737,N_1346,N_1357);
and U1738 (N_1738,N_1479,N_1340);
or U1739 (N_1739,N_1329,N_1284);
xor U1740 (N_1740,N_1468,N_1436);
and U1741 (N_1741,N_1415,N_1449);
xnor U1742 (N_1742,N_1432,N_1436);
nor U1743 (N_1743,N_1307,N_1429);
xnor U1744 (N_1744,N_1490,N_1269);
or U1745 (N_1745,N_1317,N_1304);
nor U1746 (N_1746,N_1398,N_1465);
nor U1747 (N_1747,N_1452,N_1382);
nand U1748 (N_1748,N_1262,N_1341);
nor U1749 (N_1749,N_1310,N_1471);
and U1750 (N_1750,N_1500,N_1623);
nand U1751 (N_1751,N_1624,N_1613);
nor U1752 (N_1752,N_1636,N_1568);
and U1753 (N_1753,N_1720,N_1687);
and U1754 (N_1754,N_1610,N_1630);
nand U1755 (N_1755,N_1546,N_1554);
nand U1756 (N_1756,N_1596,N_1682);
or U1757 (N_1757,N_1559,N_1525);
nor U1758 (N_1758,N_1659,N_1694);
xor U1759 (N_1759,N_1701,N_1523);
xnor U1760 (N_1760,N_1593,N_1529);
nand U1761 (N_1761,N_1521,N_1735);
or U1762 (N_1762,N_1717,N_1697);
nor U1763 (N_1763,N_1567,N_1738);
nand U1764 (N_1764,N_1732,N_1584);
nor U1765 (N_1765,N_1619,N_1668);
nand U1766 (N_1766,N_1536,N_1511);
nand U1767 (N_1767,N_1696,N_1582);
or U1768 (N_1768,N_1604,N_1565);
and U1769 (N_1769,N_1503,N_1628);
xnor U1770 (N_1770,N_1540,N_1736);
or U1771 (N_1771,N_1541,N_1656);
nand U1772 (N_1772,N_1716,N_1742);
nor U1773 (N_1773,N_1626,N_1555);
nor U1774 (N_1774,N_1556,N_1722);
nand U1775 (N_1775,N_1648,N_1739);
nand U1776 (N_1776,N_1657,N_1572);
and U1777 (N_1777,N_1614,N_1514);
nor U1778 (N_1778,N_1641,N_1598);
xnor U1779 (N_1779,N_1534,N_1527);
xor U1780 (N_1780,N_1689,N_1562);
nand U1781 (N_1781,N_1729,N_1719);
nand U1782 (N_1782,N_1745,N_1666);
xor U1783 (N_1783,N_1590,N_1520);
nand U1784 (N_1784,N_1714,N_1606);
nand U1785 (N_1785,N_1603,N_1658);
and U1786 (N_1786,N_1721,N_1634);
and U1787 (N_1787,N_1539,N_1519);
nand U1788 (N_1788,N_1600,N_1609);
nor U1789 (N_1789,N_1535,N_1671);
or U1790 (N_1790,N_1505,N_1607);
and U1791 (N_1791,N_1728,N_1680);
nand U1792 (N_1792,N_1618,N_1605);
nand U1793 (N_1793,N_1678,N_1727);
nand U1794 (N_1794,N_1578,N_1509);
or U1795 (N_1795,N_1670,N_1652);
xnor U1796 (N_1796,N_1744,N_1617);
nor U1797 (N_1797,N_1653,N_1686);
nor U1798 (N_1798,N_1608,N_1583);
xor U1799 (N_1799,N_1643,N_1580);
nand U1800 (N_1800,N_1508,N_1507);
or U1801 (N_1801,N_1734,N_1573);
or U1802 (N_1802,N_1704,N_1691);
nor U1803 (N_1803,N_1677,N_1601);
nand U1804 (N_1804,N_1703,N_1602);
nand U1805 (N_1805,N_1698,N_1581);
or U1806 (N_1806,N_1522,N_1551);
nand U1807 (N_1807,N_1501,N_1661);
xor U1808 (N_1808,N_1595,N_1599);
or U1809 (N_1809,N_1748,N_1547);
and U1810 (N_1810,N_1564,N_1663);
nand U1811 (N_1811,N_1635,N_1557);
nand U1812 (N_1812,N_1673,N_1640);
and U1813 (N_1813,N_1711,N_1611);
or U1814 (N_1814,N_1639,N_1589);
nand U1815 (N_1815,N_1528,N_1526);
or U1816 (N_1816,N_1705,N_1684);
xnor U1817 (N_1817,N_1708,N_1615);
xor U1818 (N_1818,N_1749,N_1622);
or U1819 (N_1819,N_1741,N_1740);
nor U1820 (N_1820,N_1518,N_1669);
or U1821 (N_1821,N_1588,N_1594);
or U1822 (N_1822,N_1538,N_1621);
xnor U1823 (N_1823,N_1700,N_1627);
xor U1824 (N_1824,N_1570,N_1707);
nor U1825 (N_1825,N_1517,N_1649);
nor U1826 (N_1826,N_1625,N_1654);
nor U1827 (N_1827,N_1537,N_1549);
or U1828 (N_1828,N_1706,N_1664);
nand U1829 (N_1829,N_1579,N_1510);
and U1830 (N_1830,N_1515,N_1699);
nor U1831 (N_1831,N_1672,N_1662);
nor U1832 (N_1832,N_1548,N_1545);
nand U1833 (N_1833,N_1633,N_1660);
xnor U1834 (N_1834,N_1731,N_1747);
or U1835 (N_1835,N_1576,N_1544);
nor U1836 (N_1836,N_1569,N_1550);
or U1837 (N_1837,N_1693,N_1560);
nor U1838 (N_1838,N_1533,N_1710);
nor U1839 (N_1839,N_1552,N_1644);
or U1840 (N_1840,N_1531,N_1718);
nor U1841 (N_1841,N_1530,N_1692);
or U1842 (N_1842,N_1638,N_1616);
nand U1843 (N_1843,N_1712,N_1577);
and U1844 (N_1844,N_1512,N_1685);
nand U1845 (N_1845,N_1506,N_1504);
and U1846 (N_1846,N_1637,N_1746);
nand U1847 (N_1847,N_1702,N_1502);
nor U1848 (N_1848,N_1715,N_1725);
nor U1849 (N_1849,N_1674,N_1651);
and U1850 (N_1850,N_1713,N_1683);
xor U1851 (N_1851,N_1558,N_1655);
or U1852 (N_1852,N_1646,N_1586);
or U1853 (N_1853,N_1575,N_1730);
or U1854 (N_1854,N_1709,N_1681);
xor U1855 (N_1855,N_1612,N_1690);
nand U1856 (N_1856,N_1543,N_1532);
and U1857 (N_1857,N_1585,N_1733);
or U1858 (N_1858,N_1645,N_1566);
or U1859 (N_1859,N_1676,N_1675);
nand U1860 (N_1860,N_1516,N_1724);
and U1861 (N_1861,N_1688,N_1667);
xnor U1862 (N_1862,N_1542,N_1665);
xnor U1863 (N_1863,N_1524,N_1574);
or U1864 (N_1864,N_1587,N_1650);
nand U1865 (N_1865,N_1632,N_1631);
xnor U1866 (N_1866,N_1726,N_1597);
xor U1867 (N_1867,N_1737,N_1561);
nand U1868 (N_1868,N_1513,N_1647);
and U1869 (N_1869,N_1591,N_1695);
and U1870 (N_1870,N_1679,N_1571);
and U1871 (N_1871,N_1743,N_1629);
and U1872 (N_1872,N_1723,N_1620);
or U1873 (N_1873,N_1563,N_1553);
nand U1874 (N_1874,N_1592,N_1642);
or U1875 (N_1875,N_1551,N_1707);
xnor U1876 (N_1876,N_1515,N_1693);
xnor U1877 (N_1877,N_1569,N_1595);
and U1878 (N_1878,N_1724,N_1727);
nand U1879 (N_1879,N_1505,N_1693);
nand U1880 (N_1880,N_1615,N_1546);
and U1881 (N_1881,N_1562,N_1735);
nor U1882 (N_1882,N_1651,N_1576);
nand U1883 (N_1883,N_1575,N_1528);
nor U1884 (N_1884,N_1534,N_1579);
or U1885 (N_1885,N_1631,N_1516);
or U1886 (N_1886,N_1530,N_1543);
xor U1887 (N_1887,N_1666,N_1691);
and U1888 (N_1888,N_1723,N_1739);
nand U1889 (N_1889,N_1650,N_1733);
nand U1890 (N_1890,N_1566,N_1680);
or U1891 (N_1891,N_1528,N_1518);
and U1892 (N_1892,N_1535,N_1580);
xor U1893 (N_1893,N_1719,N_1732);
and U1894 (N_1894,N_1575,N_1731);
or U1895 (N_1895,N_1588,N_1685);
and U1896 (N_1896,N_1706,N_1715);
xnor U1897 (N_1897,N_1600,N_1551);
nor U1898 (N_1898,N_1704,N_1673);
xnor U1899 (N_1899,N_1708,N_1709);
or U1900 (N_1900,N_1502,N_1740);
and U1901 (N_1901,N_1544,N_1599);
or U1902 (N_1902,N_1571,N_1553);
xor U1903 (N_1903,N_1509,N_1613);
nand U1904 (N_1904,N_1534,N_1531);
nand U1905 (N_1905,N_1629,N_1547);
nor U1906 (N_1906,N_1624,N_1712);
nand U1907 (N_1907,N_1710,N_1566);
or U1908 (N_1908,N_1507,N_1693);
nand U1909 (N_1909,N_1522,N_1685);
nor U1910 (N_1910,N_1680,N_1557);
and U1911 (N_1911,N_1739,N_1649);
or U1912 (N_1912,N_1551,N_1678);
and U1913 (N_1913,N_1655,N_1639);
nand U1914 (N_1914,N_1538,N_1552);
xor U1915 (N_1915,N_1748,N_1648);
nand U1916 (N_1916,N_1655,N_1625);
nor U1917 (N_1917,N_1667,N_1558);
xnor U1918 (N_1918,N_1741,N_1551);
xor U1919 (N_1919,N_1690,N_1735);
nor U1920 (N_1920,N_1735,N_1530);
or U1921 (N_1921,N_1672,N_1528);
nand U1922 (N_1922,N_1589,N_1534);
nor U1923 (N_1923,N_1560,N_1712);
and U1924 (N_1924,N_1542,N_1623);
xor U1925 (N_1925,N_1578,N_1719);
and U1926 (N_1926,N_1729,N_1541);
xnor U1927 (N_1927,N_1733,N_1747);
nor U1928 (N_1928,N_1734,N_1556);
or U1929 (N_1929,N_1709,N_1661);
nor U1930 (N_1930,N_1658,N_1709);
and U1931 (N_1931,N_1533,N_1666);
and U1932 (N_1932,N_1689,N_1534);
or U1933 (N_1933,N_1594,N_1724);
xor U1934 (N_1934,N_1513,N_1638);
xor U1935 (N_1935,N_1536,N_1643);
nand U1936 (N_1936,N_1521,N_1602);
nand U1937 (N_1937,N_1617,N_1559);
nand U1938 (N_1938,N_1632,N_1530);
nor U1939 (N_1939,N_1668,N_1630);
nand U1940 (N_1940,N_1592,N_1604);
nand U1941 (N_1941,N_1625,N_1662);
nor U1942 (N_1942,N_1690,N_1604);
nor U1943 (N_1943,N_1698,N_1621);
nand U1944 (N_1944,N_1697,N_1613);
and U1945 (N_1945,N_1517,N_1729);
and U1946 (N_1946,N_1649,N_1718);
nor U1947 (N_1947,N_1734,N_1553);
xnor U1948 (N_1948,N_1653,N_1588);
nor U1949 (N_1949,N_1539,N_1525);
or U1950 (N_1950,N_1721,N_1548);
and U1951 (N_1951,N_1570,N_1672);
nand U1952 (N_1952,N_1557,N_1568);
and U1953 (N_1953,N_1570,N_1657);
nor U1954 (N_1954,N_1547,N_1529);
nand U1955 (N_1955,N_1666,N_1633);
nand U1956 (N_1956,N_1545,N_1735);
xor U1957 (N_1957,N_1659,N_1624);
and U1958 (N_1958,N_1536,N_1675);
xnor U1959 (N_1959,N_1530,N_1625);
and U1960 (N_1960,N_1582,N_1655);
and U1961 (N_1961,N_1510,N_1697);
and U1962 (N_1962,N_1556,N_1547);
nor U1963 (N_1963,N_1709,N_1536);
xor U1964 (N_1964,N_1549,N_1558);
and U1965 (N_1965,N_1656,N_1533);
and U1966 (N_1966,N_1528,N_1602);
nor U1967 (N_1967,N_1567,N_1599);
or U1968 (N_1968,N_1501,N_1704);
nand U1969 (N_1969,N_1567,N_1604);
nor U1970 (N_1970,N_1595,N_1637);
or U1971 (N_1971,N_1571,N_1620);
or U1972 (N_1972,N_1564,N_1735);
nor U1973 (N_1973,N_1603,N_1711);
or U1974 (N_1974,N_1553,N_1539);
nor U1975 (N_1975,N_1536,N_1732);
or U1976 (N_1976,N_1654,N_1586);
xor U1977 (N_1977,N_1714,N_1664);
nor U1978 (N_1978,N_1678,N_1681);
xor U1979 (N_1979,N_1635,N_1583);
or U1980 (N_1980,N_1623,N_1724);
nand U1981 (N_1981,N_1522,N_1595);
nand U1982 (N_1982,N_1550,N_1626);
and U1983 (N_1983,N_1530,N_1516);
and U1984 (N_1984,N_1662,N_1653);
nand U1985 (N_1985,N_1614,N_1707);
xnor U1986 (N_1986,N_1543,N_1616);
xnor U1987 (N_1987,N_1642,N_1580);
nand U1988 (N_1988,N_1507,N_1655);
xnor U1989 (N_1989,N_1633,N_1749);
nor U1990 (N_1990,N_1502,N_1728);
xor U1991 (N_1991,N_1516,N_1609);
xor U1992 (N_1992,N_1569,N_1656);
xor U1993 (N_1993,N_1509,N_1646);
nor U1994 (N_1994,N_1685,N_1636);
and U1995 (N_1995,N_1665,N_1727);
nor U1996 (N_1996,N_1562,N_1724);
nor U1997 (N_1997,N_1615,N_1730);
or U1998 (N_1998,N_1724,N_1661);
nand U1999 (N_1999,N_1640,N_1679);
or U2000 (N_2000,N_1825,N_1827);
or U2001 (N_2001,N_1776,N_1979);
nor U2002 (N_2002,N_1759,N_1910);
nor U2003 (N_2003,N_1922,N_1750);
and U2004 (N_2004,N_1977,N_1796);
or U2005 (N_2005,N_1804,N_1945);
nor U2006 (N_2006,N_1915,N_1960);
xor U2007 (N_2007,N_1807,N_1919);
nor U2008 (N_2008,N_1940,N_1912);
nor U2009 (N_2009,N_1898,N_1846);
and U2010 (N_2010,N_1782,N_1947);
xor U2011 (N_2011,N_1793,N_1978);
and U2012 (N_2012,N_1891,N_1791);
and U2013 (N_2013,N_1802,N_1789);
nand U2014 (N_2014,N_1808,N_1973);
or U2015 (N_2015,N_1805,N_1844);
or U2016 (N_2016,N_1989,N_1943);
nor U2017 (N_2017,N_1905,N_1930);
or U2018 (N_2018,N_1830,N_1834);
xnor U2019 (N_2019,N_1974,N_1786);
nor U2020 (N_2020,N_1816,N_1884);
xor U2021 (N_2021,N_1933,N_1887);
nand U2022 (N_2022,N_1769,N_1963);
xnor U2023 (N_2023,N_1758,N_1794);
nand U2024 (N_2024,N_1843,N_1941);
or U2025 (N_2025,N_1764,N_1765);
or U2026 (N_2026,N_1952,N_1932);
nand U2027 (N_2027,N_1909,N_1861);
nor U2028 (N_2028,N_1926,N_1876);
nand U2029 (N_2029,N_1879,N_1913);
or U2030 (N_2030,N_1781,N_1775);
nor U2031 (N_2031,N_1835,N_1972);
or U2032 (N_2032,N_1936,N_1755);
nor U2033 (N_2033,N_1761,N_1931);
nand U2034 (N_2034,N_1833,N_1837);
or U2035 (N_2035,N_1859,N_1815);
or U2036 (N_2036,N_1824,N_1939);
and U2037 (N_2037,N_1895,N_1823);
and U2038 (N_2038,N_1868,N_1871);
nand U2039 (N_2039,N_1799,N_1787);
nor U2040 (N_2040,N_1928,N_1961);
nor U2041 (N_2041,N_1773,N_1997);
or U2042 (N_2042,N_1867,N_1770);
and U2043 (N_2043,N_1903,N_1965);
nor U2044 (N_2044,N_1756,N_1763);
nand U2045 (N_2045,N_1766,N_1831);
or U2046 (N_2046,N_1762,N_1858);
nor U2047 (N_2047,N_1829,N_1784);
nand U2048 (N_2048,N_1872,N_1814);
and U2049 (N_2049,N_1991,N_1818);
and U2050 (N_2050,N_1955,N_1878);
xor U2051 (N_2051,N_1800,N_1757);
and U2052 (N_2052,N_1969,N_1767);
xnor U2053 (N_2053,N_1754,N_1962);
nand U2054 (N_2054,N_1987,N_1803);
xnor U2055 (N_2055,N_1988,N_1946);
or U2056 (N_2056,N_1995,N_1981);
and U2057 (N_2057,N_1953,N_1900);
nand U2058 (N_2058,N_1854,N_1883);
or U2059 (N_2059,N_1964,N_1990);
xnor U2060 (N_2060,N_1821,N_1798);
or U2061 (N_2061,N_1893,N_1849);
nand U2062 (N_2062,N_1848,N_1958);
nand U2063 (N_2063,N_1842,N_1840);
nand U2064 (N_2064,N_1896,N_1966);
nand U2065 (N_2065,N_1869,N_1795);
nand U2066 (N_2066,N_1812,N_1771);
xor U2067 (N_2067,N_1968,N_1957);
and U2068 (N_2068,N_1820,N_1847);
and U2069 (N_2069,N_1850,N_1942);
nor U2070 (N_2070,N_1866,N_1918);
or U2071 (N_2071,N_1870,N_1982);
xnor U2072 (N_2072,N_1772,N_1778);
and U2073 (N_2073,N_1934,N_1841);
nor U2074 (N_2074,N_1954,N_1901);
or U2075 (N_2075,N_1992,N_1873);
nand U2076 (N_2076,N_1894,N_1851);
or U2077 (N_2077,N_1863,N_1852);
nor U2078 (N_2078,N_1949,N_1985);
and U2079 (N_2079,N_1886,N_1788);
and U2080 (N_2080,N_1984,N_1865);
nand U2081 (N_2081,N_1785,N_1986);
xnor U2082 (N_2082,N_1881,N_1906);
and U2083 (N_2083,N_1864,N_1888);
nand U2084 (N_2084,N_1811,N_1853);
and U2085 (N_2085,N_1937,N_1828);
and U2086 (N_2086,N_1790,N_1976);
xor U2087 (N_2087,N_1877,N_1938);
xor U2088 (N_2088,N_1845,N_1819);
and U2089 (N_2089,N_1809,N_1857);
xnor U2090 (N_2090,N_1917,N_1999);
nor U2091 (N_2091,N_1924,N_1929);
nand U2092 (N_2092,N_1993,N_1806);
xor U2093 (N_2093,N_1760,N_1907);
nor U2094 (N_2094,N_1948,N_1792);
nand U2095 (N_2095,N_1882,N_1914);
or U2096 (N_2096,N_1921,N_1768);
nor U2097 (N_2097,N_1855,N_1959);
xnor U2098 (N_2098,N_1810,N_1890);
and U2099 (N_2099,N_1874,N_1862);
or U2100 (N_2100,N_1885,N_1801);
or U2101 (N_2101,N_1899,N_1994);
and U2102 (N_2102,N_1980,N_1975);
xor U2103 (N_2103,N_1783,N_1780);
or U2104 (N_2104,N_1967,N_1897);
and U2105 (N_2105,N_1860,N_1777);
nor U2106 (N_2106,N_1970,N_1779);
and U2107 (N_2107,N_1856,N_1889);
or U2108 (N_2108,N_1817,N_1832);
and U2109 (N_2109,N_1998,N_1797);
and U2110 (N_2110,N_1927,N_1902);
and U2111 (N_2111,N_1951,N_1983);
xnor U2112 (N_2112,N_1956,N_1923);
or U2113 (N_2113,N_1751,N_1908);
nor U2114 (N_2114,N_1822,N_1904);
or U2115 (N_2115,N_1880,N_1838);
and U2116 (N_2116,N_1996,N_1925);
or U2117 (N_2117,N_1892,N_1774);
nor U2118 (N_2118,N_1875,N_1950);
nand U2119 (N_2119,N_1911,N_1935);
nor U2120 (N_2120,N_1971,N_1839);
or U2121 (N_2121,N_1836,N_1753);
xor U2122 (N_2122,N_1826,N_1944);
and U2123 (N_2123,N_1916,N_1752);
and U2124 (N_2124,N_1920,N_1813);
or U2125 (N_2125,N_1779,N_1806);
xor U2126 (N_2126,N_1761,N_1992);
xor U2127 (N_2127,N_1936,N_1758);
or U2128 (N_2128,N_1902,N_1897);
or U2129 (N_2129,N_1971,N_1809);
xnor U2130 (N_2130,N_1834,N_1972);
or U2131 (N_2131,N_1853,N_1820);
nor U2132 (N_2132,N_1912,N_1933);
nand U2133 (N_2133,N_1944,N_1905);
xor U2134 (N_2134,N_1817,N_1807);
or U2135 (N_2135,N_1772,N_1904);
and U2136 (N_2136,N_1942,N_1959);
xor U2137 (N_2137,N_1783,N_1927);
nor U2138 (N_2138,N_1986,N_1845);
or U2139 (N_2139,N_1814,N_1787);
and U2140 (N_2140,N_1778,N_1768);
nor U2141 (N_2141,N_1922,N_1883);
nor U2142 (N_2142,N_1760,N_1950);
and U2143 (N_2143,N_1780,N_1852);
and U2144 (N_2144,N_1926,N_1809);
xnor U2145 (N_2145,N_1881,N_1803);
or U2146 (N_2146,N_1860,N_1932);
xnor U2147 (N_2147,N_1797,N_1773);
or U2148 (N_2148,N_1920,N_1833);
nand U2149 (N_2149,N_1945,N_1879);
nor U2150 (N_2150,N_1851,N_1771);
nand U2151 (N_2151,N_1927,N_1986);
nor U2152 (N_2152,N_1890,N_1886);
or U2153 (N_2153,N_1851,N_1827);
nand U2154 (N_2154,N_1837,N_1804);
xnor U2155 (N_2155,N_1857,N_1814);
or U2156 (N_2156,N_1839,N_1944);
and U2157 (N_2157,N_1887,N_1824);
and U2158 (N_2158,N_1996,N_1851);
and U2159 (N_2159,N_1965,N_1960);
xnor U2160 (N_2160,N_1908,N_1874);
nor U2161 (N_2161,N_1759,N_1940);
xor U2162 (N_2162,N_1955,N_1997);
or U2163 (N_2163,N_1893,N_1915);
and U2164 (N_2164,N_1928,N_1973);
nor U2165 (N_2165,N_1928,N_1984);
nor U2166 (N_2166,N_1825,N_1899);
nor U2167 (N_2167,N_1822,N_1854);
and U2168 (N_2168,N_1895,N_1808);
or U2169 (N_2169,N_1826,N_1857);
nand U2170 (N_2170,N_1982,N_1782);
or U2171 (N_2171,N_1884,N_1838);
or U2172 (N_2172,N_1931,N_1870);
nor U2173 (N_2173,N_1952,N_1973);
or U2174 (N_2174,N_1758,N_1945);
or U2175 (N_2175,N_1783,N_1826);
nor U2176 (N_2176,N_1987,N_1851);
nand U2177 (N_2177,N_1777,N_1804);
and U2178 (N_2178,N_1940,N_1798);
xnor U2179 (N_2179,N_1898,N_1978);
nand U2180 (N_2180,N_1923,N_1938);
nand U2181 (N_2181,N_1855,N_1990);
or U2182 (N_2182,N_1753,N_1961);
xnor U2183 (N_2183,N_1790,N_1995);
and U2184 (N_2184,N_1968,N_1838);
nor U2185 (N_2185,N_1826,N_1862);
nor U2186 (N_2186,N_1991,N_1836);
or U2187 (N_2187,N_1950,N_1818);
xor U2188 (N_2188,N_1815,N_1877);
nor U2189 (N_2189,N_1888,N_1857);
or U2190 (N_2190,N_1813,N_1941);
or U2191 (N_2191,N_1830,N_1990);
or U2192 (N_2192,N_1800,N_1917);
or U2193 (N_2193,N_1911,N_1940);
nor U2194 (N_2194,N_1787,N_1955);
nand U2195 (N_2195,N_1790,N_1905);
nand U2196 (N_2196,N_1779,N_1975);
and U2197 (N_2197,N_1908,N_1970);
nand U2198 (N_2198,N_1760,N_1863);
or U2199 (N_2199,N_1805,N_1883);
or U2200 (N_2200,N_1908,N_1850);
nor U2201 (N_2201,N_1964,N_1815);
and U2202 (N_2202,N_1972,N_1802);
or U2203 (N_2203,N_1933,N_1876);
and U2204 (N_2204,N_1910,N_1765);
xnor U2205 (N_2205,N_1877,N_1882);
and U2206 (N_2206,N_1991,N_1822);
nor U2207 (N_2207,N_1879,N_1914);
xor U2208 (N_2208,N_1892,N_1783);
and U2209 (N_2209,N_1761,N_1965);
and U2210 (N_2210,N_1930,N_1966);
xnor U2211 (N_2211,N_1840,N_1935);
and U2212 (N_2212,N_1855,N_1802);
or U2213 (N_2213,N_1905,N_1872);
nor U2214 (N_2214,N_1861,N_1907);
xnor U2215 (N_2215,N_1902,N_1992);
xor U2216 (N_2216,N_1997,N_1996);
nand U2217 (N_2217,N_1807,N_1921);
and U2218 (N_2218,N_1866,N_1846);
nor U2219 (N_2219,N_1918,N_1991);
nor U2220 (N_2220,N_1949,N_1800);
or U2221 (N_2221,N_1816,N_1929);
xor U2222 (N_2222,N_1759,N_1907);
xor U2223 (N_2223,N_1863,N_1934);
nand U2224 (N_2224,N_1841,N_1835);
nor U2225 (N_2225,N_1986,N_1759);
xor U2226 (N_2226,N_1768,N_1905);
or U2227 (N_2227,N_1908,N_1760);
or U2228 (N_2228,N_1890,N_1763);
or U2229 (N_2229,N_1763,N_1787);
or U2230 (N_2230,N_1913,N_1899);
nor U2231 (N_2231,N_1761,N_1849);
and U2232 (N_2232,N_1956,N_1907);
nand U2233 (N_2233,N_1803,N_1815);
xor U2234 (N_2234,N_1752,N_1956);
xor U2235 (N_2235,N_1811,N_1863);
and U2236 (N_2236,N_1880,N_1969);
nand U2237 (N_2237,N_1873,N_1915);
xnor U2238 (N_2238,N_1914,N_1791);
xnor U2239 (N_2239,N_1996,N_1918);
nand U2240 (N_2240,N_1863,N_1796);
nor U2241 (N_2241,N_1959,N_1883);
nand U2242 (N_2242,N_1804,N_1861);
xor U2243 (N_2243,N_1822,N_1785);
nand U2244 (N_2244,N_1910,N_1907);
nor U2245 (N_2245,N_1935,N_1946);
xnor U2246 (N_2246,N_1877,N_1976);
and U2247 (N_2247,N_1975,N_1938);
and U2248 (N_2248,N_1928,N_1896);
nand U2249 (N_2249,N_1928,N_1999);
nand U2250 (N_2250,N_2101,N_2245);
xnor U2251 (N_2251,N_2048,N_2131);
xnor U2252 (N_2252,N_2188,N_2097);
nand U2253 (N_2253,N_2029,N_2244);
nand U2254 (N_2254,N_2104,N_2110);
and U2255 (N_2255,N_2064,N_2023);
nor U2256 (N_2256,N_2020,N_2147);
nand U2257 (N_2257,N_2070,N_2229);
nor U2258 (N_2258,N_2067,N_2167);
xor U2259 (N_2259,N_2010,N_2166);
or U2260 (N_2260,N_2021,N_2078);
xnor U2261 (N_2261,N_2124,N_2194);
nand U2262 (N_2262,N_2084,N_2115);
and U2263 (N_2263,N_2180,N_2211);
nand U2264 (N_2264,N_2226,N_2044);
and U2265 (N_2265,N_2246,N_2248);
or U2266 (N_2266,N_2090,N_2050);
and U2267 (N_2267,N_2122,N_2007);
xnor U2268 (N_2268,N_2158,N_2231);
xnor U2269 (N_2269,N_2154,N_2125);
nor U2270 (N_2270,N_2111,N_2149);
and U2271 (N_2271,N_2026,N_2198);
nor U2272 (N_2272,N_2016,N_2212);
xnor U2273 (N_2273,N_2195,N_2039);
xnor U2274 (N_2274,N_2144,N_2162);
nor U2275 (N_2275,N_2199,N_2132);
or U2276 (N_2276,N_2060,N_2200);
or U2277 (N_2277,N_2213,N_2241);
or U2278 (N_2278,N_2099,N_2221);
xnor U2279 (N_2279,N_2076,N_2160);
nand U2280 (N_2280,N_2164,N_2031);
nor U2281 (N_2281,N_2170,N_2127);
and U2282 (N_2282,N_2239,N_2201);
or U2283 (N_2283,N_2156,N_2142);
or U2284 (N_2284,N_2152,N_2175);
nand U2285 (N_2285,N_2037,N_2063);
and U2286 (N_2286,N_2208,N_2151);
nor U2287 (N_2287,N_2035,N_2058);
and U2288 (N_2288,N_2045,N_2014);
or U2289 (N_2289,N_2069,N_2103);
xnor U2290 (N_2290,N_2001,N_2011);
nand U2291 (N_2291,N_2171,N_2242);
or U2292 (N_2292,N_2236,N_2006);
nand U2293 (N_2293,N_2193,N_2109);
nand U2294 (N_2294,N_2140,N_2093);
and U2295 (N_2295,N_2049,N_2249);
nand U2296 (N_2296,N_2214,N_2012);
nor U2297 (N_2297,N_2190,N_2185);
nand U2298 (N_2298,N_2098,N_2008);
nand U2299 (N_2299,N_2187,N_2106);
nor U2300 (N_2300,N_2203,N_2182);
nor U2301 (N_2301,N_2159,N_2080);
or U2302 (N_2302,N_2136,N_2230);
nor U2303 (N_2303,N_2222,N_2041);
and U2304 (N_2304,N_2072,N_2161);
nand U2305 (N_2305,N_2218,N_2219);
or U2306 (N_2306,N_2217,N_2032);
xnor U2307 (N_2307,N_2234,N_2054);
xnor U2308 (N_2308,N_2105,N_2100);
nor U2309 (N_2309,N_2243,N_2112);
nand U2310 (N_2310,N_2224,N_2068);
nor U2311 (N_2311,N_2247,N_2220);
or U2312 (N_2312,N_2184,N_2138);
xnor U2313 (N_2313,N_2133,N_2077);
or U2314 (N_2314,N_2204,N_2233);
or U2315 (N_2315,N_2191,N_2118);
nand U2316 (N_2316,N_2134,N_2150);
nand U2317 (N_2317,N_2196,N_2225);
nand U2318 (N_2318,N_2096,N_2024);
nor U2319 (N_2319,N_2197,N_2051);
xor U2320 (N_2320,N_2177,N_2013);
and U2321 (N_2321,N_2000,N_2108);
and U2322 (N_2322,N_2209,N_2227);
or U2323 (N_2323,N_2181,N_2082);
nor U2324 (N_2324,N_2206,N_2216);
xnor U2325 (N_2325,N_2085,N_2176);
xnor U2326 (N_2326,N_2129,N_2215);
or U2327 (N_2327,N_2119,N_2179);
and U2328 (N_2328,N_2030,N_2043);
nor U2329 (N_2329,N_2040,N_2089);
xnor U2330 (N_2330,N_2065,N_2107);
nor U2331 (N_2331,N_2192,N_2086);
or U2332 (N_2332,N_2172,N_2141);
nor U2333 (N_2333,N_2126,N_2033);
xor U2334 (N_2334,N_2052,N_2128);
and U2335 (N_2335,N_2153,N_2235);
nor U2336 (N_2336,N_2120,N_2117);
nand U2337 (N_2337,N_2146,N_2036);
xnor U2338 (N_2338,N_2238,N_2083);
xor U2339 (N_2339,N_2228,N_2074);
xnor U2340 (N_2340,N_2165,N_2057);
nand U2341 (N_2341,N_2075,N_2205);
xnor U2342 (N_2342,N_2237,N_2062);
nand U2343 (N_2343,N_2116,N_2202);
xor U2344 (N_2344,N_2059,N_2114);
or U2345 (N_2345,N_2079,N_2027);
xnor U2346 (N_2346,N_2092,N_2137);
nand U2347 (N_2347,N_2002,N_2143);
nand U2348 (N_2348,N_2113,N_2022);
xnor U2349 (N_2349,N_2157,N_2130);
and U2350 (N_2350,N_2148,N_2163);
xnor U2351 (N_2351,N_2210,N_2056);
xnor U2352 (N_2352,N_2028,N_2017);
xnor U2353 (N_2353,N_2061,N_2088);
and U2354 (N_2354,N_2055,N_2025);
nor U2355 (N_2355,N_2240,N_2174);
nor U2356 (N_2356,N_2189,N_2094);
or U2357 (N_2357,N_2071,N_2066);
or U2358 (N_2358,N_2073,N_2169);
nand U2359 (N_2359,N_2042,N_2183);
nor U2360 (N_2360,N_2038,N_2015);
xor U2361 (N_2361,N_2123,N_2095);
and U2362 (N_2362,N_2121,N_2019);
xnor U2363 (N_2363,N_2091,N_2173);
nand U2364 (N_2364,N_2053,N_2145);
nor U2365 (N_2365,N_2186,N_2223);
nor U2366 (N_2366,N_2207,N_2005);
nand U2367 (N_2367,N_2081,N_2034);
nor U2368 (N_2368,N_2046,N_2003);
xor U2369 (N_2369,N_2178,N_2232);
and U2370 (N_2370,N_2102,N_2139);
nand U2371 (N_2371,N_2155,N_2018);
nand U2372 (N_2372,N_2087,N_2004);
or U2373 (N_2373,N_2168,N_2009);
xor U2374 (N_2374,N_2047,N_2135);
or U2375 (N_2375,N_2228,N_2078);
nor U2376 (N_2376,N_2155,N_2242);
and U2377 (N_2377,N_2032,N_2243);
nor U2378 (N_2378,N_2207,N_2191);
xor U2379 (N_2379,N_2213,N_2087);
xnor U2380 (N_2380,N_2033,N_2112);
or U2381 (N_2381,N_2023,N_2140);
nor U2382 (N_2382,N_2095,N_2112);
nand U2383 (N_2383,N_2030,N_2146);
and U2384 (N_2384,N_2109,N_2192);
nor U2385 (N_2385,N_2139,N_2045);
nand U2386 (N_2386,N_2116,N_2195);
nor U2387 (N_2387,N_2063,N_2175);
xnor U2388 (N_2388,N_2080,N_2003);
nand U2389 (N_2389,N_2149,N_2060);
xnor U2390 (N_2390,N_2050,N_2146);
nor U2391 (N_2391,N_2020,N_2207);
and U2392 (N_2392,N_2185,N_2114);
and U2393 (N_2393,N_2085,N_2043);
xnor U2394 (N_2394,N_2154,N_2213);
and U2395 (N_2395,N_2139,N_2228);
nor U2396 (N_2396,N_2208,N_2038);
or U2397 (N_2397,N_2129,N_2154);
nor U2398 (N_2398,N_2181,N_2217);
xor U2399 (N_2399,N_2139,N_2198);
nand U2400 (N_2400,N_2204,N_2062);
and U2401 (N_2401,N_2057,N_2229);
xor U2402 (N_2402,N_2041,N_2179);
and U2403 (N_2403,N_2200,N_2231);
nor U2404 (N_2404,N_2085,N_2047);
nor U2405 (N_2405,N_2211,N_2245);
nand U2406 (N_2406,N_2058,N_2109);
nor U2407 (N_2407,N_2001,N_2014);
and U2408 (N_2408,N_2025,N_2119);
xor U2409 (N_2409,N_2011,N_2009);
xor U2410 (N_2410,N_2009,N_2160);
and U2411 (N_2411,N_2224,N_2216);
nand U2412 (N_2412,N_2087,N_2110);
xor U2413 (N_2413,N_2204,N_2007);
nor U2414 (N_2414,N_2045,N_2127);
nor U2415 (N_2415,N_2079,N_2003);
and U2416 (N_2416,N_2033,N_2034);
nor U2417 (N_2417,N_2247,N_2245);
nand U2418 (N_2418,N_2206,N_2219);
nand U2419 (N_2419,N_2090,N_2156);
and U2420 (N_2420,N_2002,N_2182);
or U2421 (N_2421,N_2162,N_2066);
nor U2422 (N_2422,N_2220,N_2173);
and U2423 (N_2423,N_2087,N_2172);
or U2424 (N_2424,N_2232,N_2038);
nand U2425 (N_2425,N_2051,N_2108);
nor U2426 (N_2426,N_2181,N_2225);
nor U2427 (N_2427,N_2220,N_2170);
or U2428 (N_2428,N_2198,N_2101);
xnor U2429 (N_2429,N_2029,N_2095);
xor U2430 (N_2430,N_2212,N_2243);
nand U2431 (N_2431,N_2013,N_2108);
or U2432 (N_2432,N_2127,N_2204);
or U2433 (N_2433,N_2146,N_2168);
nand U2434 (N_2434,N_2236,N_2031);
nand U2435 (N_2435,N_2091,N_2126);
and U2436 (N_2436,N_2133,N_2050);
and U2437 (N_2437,N_2088,N_2192);
nor U2438 (N_2438,N_2128,N_2196);
xor U2439 (N_2439,N_2007,N_2209);
nand U2440 (N_2440,N_2053,N_2035);
or U2441 (N_2441,N_2210,N_2193);
or U2442 (N_2442,N_2178,N_2169);
nor U2443 (N_2443,N_2050,N_2060);
or U2444 (N_2444,N_2019,N_2220);
nand U2445 (N_2445,N_2120,N_2162);
xnor U2446 (N_2446,N_2115,N_2130);
or U2447 (N_2447,N_2208,N_2214);
nor U2448 (N_2448,N_2039,N_2103);
nand U2449 (N_2449,N_2051,N_2061);
or U2450 (N_2450,N_2023,N_2145);
nor U2451 (N_2451,N_2092,N_2232);
nand U2452 (N_2452,N_2157,N_2225);
and U2453 (N_2453,N_2203,N_2150);
and U2454 (N_2454,N_2187,N_2052);
nor U2455 (N_2455,N_2196,N_2247);
xor U2456 (N_2456,N_2019,N_2016);
nand U2457 (N_2457,N_2060,N_2040);
and U2458 (N_2458,N_2019,N_2138);
nor U2459 (N_2459,N_2002,N_2139);
nor U2460 (N_2460,N_2146,N_2024);
xnor U2461 (N_2461,N_2129,N_2010);
nor U2462 (N_2462,N_2058,N_2249);
xor U2463 (N_2463,N_2210,N_2179);
xor U2464 (N_2464,N_2092,N_2149);
and U2465 (N_2465,N_2034,N_2055);
nor U2466 (N_2466,N_2121,N_2248);
and U2467 (N_2467,N_2131,N_2013);
xor U2468 (N_2468,N_2145,N_2144);
nand U2469 (N_2469,N_2170,N_2096);
nand U2470 (N_2470,N_2095,N_2012);
xnor U2471 (N_2471,N_2020,N_2242);
xor U2472 (N_2472,N_2119,N_2174);
nor U2473 (N_2473,N_2216,N_2032);
or U2474 (N_2474,N_2054,N_2020);
nand U2475 (N_2475,N_2153,N_2050);
nor U2476 (N_2476,N_2113,N_2024);
nand U2477 (N_2477,N_2236,N_2018);
nand U2478 (N_2478,N_2127,N_2118);
and U2479 (N_2479,N_2074,N_2009);
and U2480 (N_2480,N_2207,N_2212);
nand U2481 (N_2481,N_2161,N_2013);
nand U2482 (N_2482,N_2105,N_2124);
xnor U2483 (N_2483,N_2156,N_2125);
nand U2484 (N_2484,N_2088,N_2028);
nand U2485 (N_2485,N_2102,N_2076);
or U2486 (N_2486,N_2174,N_2243);
and U2487 (N_2487,N_2138,N_2100);
xor U2488 (N_2488,N_2148,N_2192);
or U2489 (N_2489,N_2155,N_2136);
or U2490 (N_2490,N_2153,N_2005);
nor U2491 (N_2491,N_2121,N_2032);
xnor U2492 (N_2492,N_2042,N_2188);
and U2493 (N_2493,N_2088,N_2209);
xnor U2494 (N_2494,N_2174,N_2008);
and U2495 (N_2495,N_2005,N_2196);
and U2496 (N_2496,N_2184,N_2238);
xor U2497 (N_2497,N_2167,N_2086);
xnor U2498 (N_2498,N_2238,N_2224);
or U2499 (N_2499,N_2247,N_2103);
or U2500 (N_2500,N_2405,N_2271);
nand U2501 (N_2501,N_2392,N_2364);
or U2502 (N_2502,N_2346,N_2289);
nor U2503 (N_2503,N_2439,N_2295);
and U2504 (N_2504,N_2250,N_2393);
nand U2505 (N_2505,N_2461,N_2363);
nor U2506 (N_2506,N_2314,N_2324);
nor U2507 (N_2507,N_2328,N_2491);
xnor U2508 (N_2508,N_2373,N_2469);
and U2509 (N_2509,N_2350,N_2272);
nand U2510 (N_2510,N_2296,N_2338);
nand U2511 (N_2511,N_2420,N_2342);
nor U2512 (N_2512,N_2336,N_2431);
or U2513 (N_2513,N_2395,N_2367);
xor U2514 (N_2514,N_2413,N_2270);
nand U2515 (N_2515,N_2378,N_2467);
or U2516 (N_2516,N_2290,N_2438);
and U2517 (N_2517,N_2279,N_2316);
xnor U2518 (N_2518,N_2497,N_2282);
and U2519 (N_2519,N_2425,N_2401);
and U2520 (N_2520,N_2376,N_2382);
and U2521 (N_2521,N_2479,N_2404);
or U2522 (N_2522,N_2307,N_2472);
or U2523 (N_2523,N_2453,N_2298);
and U2524 (N_2524,N_2317,N_2322);
and U2525 (N_2525,N_2487,N_2368);
nor U2526 (N_2526,N_2371,N_2285);
xor U2527 (N_2527,N_2352,N_2456);
and U2528 (N_2528,N_2441,N_2495);
nand U2529 (N_2529,N_2255,N_2449);
nand U2530 (N_2530,N_2494,N_2468);
or U2531 (N_2531,N_2433,N_2356);
nor U2532 (N_2532,N_2308,N_2471);
and U2533 (N_2533,N_2435,N_2379);
and U2534 (N_2534,N_2417,N_2277);
nor U2535 (N_2535,N_2304,N_2424);
or U2536 (N_2536,N_2349,N_2490);
or U2537 (N_2537,N_2260,N_2310);
nand U2538 (N_2538,N_2302,N_2327);
nor U2539 (N_2539,N_2443,N_2434);
and U2540 (N_2540,N_2488,N_2269);
and U2541 (N_2541,N_2278,N_2444);
nor U2542 (N_2542,N_2276,N_2403);
or U2543 (N_2543,N_2256,N_2432);
and U2544 (N_2544,N_2463,N_2442);
nand U2545 (N_2545,N_2398,N_2411);
nand U2546 (N_2546,N_2496,N_2428);
or U2547 (N_2547,N_2331,N_2418);
or U2548 (N_2548,N_2415,N_2460);
xnor U2549 (N_2549,N_2389,N_2273);
nand U2550 (N_2550,N_2281,N_2485);
xnor U2551 (N_2551,N_2450,N_2320);
and U2552 (N_2552,N_2347,N_2312);
nand U2553 (N_2553,N_2258,N_2390);
xnor U2554 (N_2554,N_2422,N_2259);
and U2555 (N_2555,N_2333,N_2429);
and U2556 (N_2556,N_2489,N_2306);
xnor U2557 (N_2557,N_2303,N_2360);
nor U2558 (N_2558,N_2459,N_2284);
and U2559 (N_2559,N_2318,N_2383);
nand U2560 (N_2560,N_2386,N_2288);
nor U2561 (N_2561,N_2266,N_2251);
nor U2562 (N_2562,N_2466,N_2354);
xor U2563 (N_2563,N_2291,N_2437);
nor U2564 (N_2564,N_2301,N_2416);
nor U2565 (N_2565,N_2447,N_2375);
or U2566 (N_2566,N_2478,N_2311);
nand U2567 (N_2567,N_2267,N_2464);
nand U2568 (N_2568,N_2355,N_2465);
or U2569 (N_2569,N_2366,N_2305);
nor U2570 (N_2570,N_2262,N_2399);
and U2571 (N_2571,N_2254,N_2365);
nand U2572 (N_2572,N_2326,N_2283);
nor U2573 (N_2573,N_2300,N_2261);
nor U2574 (N_2574,N_2387,N_2426);
and U2575 (N_2575,N_2374,N_2412);
and U2576 (N_2576,N_2483,N_2339);
nor U2577 (N_2577,N_2274,N_2293);
nand U2578 (N_2578,N_2414,N_2470);
and U2579 (N_2579,N_2323,N_2400);
nor U2580 (N_2580,N_2257,N_2391);
nand U2581 (N_2581,N_2335,N_2430);
nand U2582 (N_2582,N_2313,N_2286);
or U2583 (N_2583,N_2476,N_2292);
or U2584 (N_2584,N_2396,N_2343);
xnor U2585 (N_2585,N_2402,N_2440);
or U2586 (N_2586,N_2474,N_2407);
and U2587 (N_2587,N_2275,N_2265);
or U2588 (N_2588,N_2297,N_2340);
nand U2589 (N_2589,N_2357,N_2423);
or U2590 (N_2590,N_2280,N_2397);
and U2591 (N_2591,N_2315,N_2462);
nor U2592 (N_2592,N_2455,N_2362);
nand U2593 (N_2593,N_2330,N_2446);
and U2594 (N_2594,N_2381,N_2268);
nor U2595 (N_2595,N_2385,N_2344);
xor U2596 (N_2596,N_2345,N_2419);
nor U2597 (N_2597,N_2325,N_2406);
and U2598 (N_2598,N_2299,N_2451);
xnor U2599 (N_2599,N_2409,N_2457);
nand U2600 (N_2600,N_2499,N_2480);
and U2601 (N_2601,N_2408,N_2294);
xor U2602 (N_2602,N_2287,N_2482);
xor U2603 (N_2603,N_2337,N_2370);
and U2604 (N_2604,N_2427,N_2477);
or U2605 (N_2605,N_2394,N_2486);
xor U2606 (N_2606,N_2492,N_2380);
or U2607 (N_2607,N_2358,N_2452);
nor U2608 (N_2608,N_2372,N_2475);
nor U2609 (N_2609,N_2341,N_2484);
or U2610 (N_2610,N_2454,N_2369);
or U2611 (N_2611,N_2498,N_2253);
nand U2612 (N_2612,N_2384,N_2481);
nand U2613 (N_2613,N_2351,N_2436);
and U2614 (N_2614,N_2448,N_2263);
and U2615 (N_2615,N_2348,N_2321);
nand U2616 (N_2616,N_2421,N_2377);
and U2617 (N_2617,N_2334,N_2473);
nor U2618 (N_2618,N_2319,N_2458);
nand U2619 (N_2619,N_2329,N_2359);
and U2620 (N_2620,N_2388,N_2361);
nor U2621 (N_2621,N_2445,N_2309);
nand U2622 (N_2622,N_2252,N_2353);
nor U2623 (N_2623,N_2410,N_2332);
and U2624 (N_2624,N_2264,N_2493);
nand U2625 (N_2625,N_2406,N_2345);
and U2626 (N_2626,N_2271,N_2417);
nor U2627 (N_2627,N_2396,N_2327);
xnor U2628 (N_2628,N_2276,N_2331);
or U2629 (N_2629,N_2287,N_2494);
xnor U2630 (N_2630,N_2288,N_2470);
and U2631 (N_2631,N_2277,N_2335);
and U2632 (N_2632,N_2335,N_2320);
and U2633 (N_2633,N_2454,N_2421);
and U2634 (N_2634,N_2447,N_2320);
xnor U2635 (N_2635,N_2446,N_2374);
and U2636 (N_2636,N_2268,N_2279);
nor U2637 (N_2637,N_2393,N_2467);
xnor U2638 (N_2638,N_2294,N_2297);
or U2639 (N_2639,N_2360,N_2299);
and U2640 (N_2640,N_2417,N_2285);
nand U2641 (N_2641,N_2326,N_2381);
nor U2642 (N_2642,N_2498,N_2380);
nand U2643 (N_2643,N_2318,N_2312);
nor U2644 (N_2644,N_2286,N_2478);
nor U2645 (N_2645,N_2374,N_2369);
or U2646 (N_2646,N_2480,N_2369);
nand U2647 (N_2647,N_2269,N_2271);
xnor U2648 (N_2648,N_2487,N_2378);
nor U2649 (N_2649,N_2311,N_2464);
nor U2650 (N_2650,N_2492,N_2446);
xnor U2651 (N_2651,N_2376,N_2273);
xnor U2652 (N_2652,N_2296,N_2381);
or U2653 (N_2653,N_2277,N_2435);
nor U2654 (N_2654,N_2296,N_2452);
nand U2655 (N_2655,N_2332,N_2256);
or U2656 (N_2656,N_2492,N_2332);
and U2657 (N_2657,N_2372,N_2358);
xnor U2658 (N_2658,N_2433,N_2316);
nand U2659 (N_2659,N_2317,N_2302);
xor U2660 (N_2660,N_2336,N_2448);
nand U2661 (N_2661,N_2329,N_2270);
xnor U2662 (N_2662,N_2460,N_2319);
and U2663 (N_2663,N_2422,N_2483);
or U2664 (N_2664,N_2410,N_2370);
nor U2665 (N_2665,N_2345,N_2295);
nor U2666 (N_2666,N_2269,N_2466);
nor U2667 (N_2667,N_2471,N_2429);
nor U2668 (N_2668,N_2272,N_2389);
nand U2669 (N_2669,N_2394,N_2342);
nor U2670 (N_2670,N_2484,N_2319);
xor U2671 (N_2671,N_2440,N_2467);
xnor U2672 (N_2672,N_2254,N_2318);
nor U2673 (N_2673,N_2292,N_2428);
and U2674 (N_2674,N_2281,N_2434);
nand U2675 (N_2675,N_2468,N_2369);
nand U2676 (N_2676,N_2495,N_2420);
nand U2677 (N_2677,N_2297,N_2400);
and U2678 (N_2678,N_2340,N_2410);
nor U2679 (N_2679,N_2279,N_2307);
nand U2680 (N_2680,N_2333,N_2285);
nor U2681 (N_2681,N_2403,N_2421);
nand U2682 (N_2682,N_2456,N_2285);
nor U2683 (N_2683,N_2306,N_2483);
nor U2684 (N_2684,N_2493,N_2387);
and U2685 (N_2685,N_2366,N_2337);
xnor U2686 (N_2686,N_2433,N_2311);
nand U2687 (N_2687,N_2432,N_2469);
nand U2688 (N_2688,N_2301,N_2255);
xnor U2689 (N_2689,N_2458,N_2352);
nand U2690 (N_2690,N_2457,N_2338);
nand U2691 (N_2691,N_2423,N_2475);
xor U2692 (N_2692,N_2368,N_2291);
xor U2693 (N_2693,N_2434,N_2268);
xor U2694 (N_2694,N_2356,N_2296);
xnor U2695 (N_2695,N_2375,N_2431);
xor U2696 (N_2696,N_2297,N_2492);
nand U2697 (N_2697,N_2415,N_2280);
and U2698 (N_2698,N_2373,N_2256);
and U2699 (N_2699,N_2398,N_2287);
nand U2700 (N_2700,N_2302,N_2439);
xor U2701 (N_2701,N_2498,N_2376);
xor U2702 (N_2702,N_2298,N_2365);
xnor U2703 (N_2703,N_2269,N_2291);
nand U2704 (N_2704,N_2463,N_2415);
nand U2705 (N_2705,N_2317,N_2415);
xnor U2706 (N_2706,N_2361,N_2426);
xnor U2707 (N_2707,N_2278,N_2300);
xnor U2708 (N_2708,N_2302,N_2487);
or U2709 (N_2709,N_2480,N_2470);
and U2710 (N_2710,N_2263,N_2390);
and U2711 (N_2711,N_2459,N_2339);
xor U2712 (N_2712,N_2353,N_2457);
nor U2713 (N_2713,N_2286,N_2268);
xor U2714 (N_2714,N_2295,N_2493);
xnor U2715 (N_2715,N_2333,N_2308);
and U2716 (N_2716,N_2474,N_2469);
or U2717 (N_2717,N_2260,N_2359);
nand U2718 (N_2718,N_2326,N_2333);
nand U2719 (N_2719,N_2277,N_2481);
and U2720 (N_2720,N_2376,N_2445);
nor U2721 (N_2721,N_2495,N_2404);
nor U2722 (N_2722,N_2496,N_2284);
or U2723 (N_2723,N_2269,N_2394);
nor U2724 (N_2724,N_2278,N_2408);
and U2725 (N_2725,N_2397,N_2348);
nand U2726 (N_2726,N_2349,N_2399);
and U2727 (N_2727,N_2410,N_2278);
nand U2728 (N_2728,N_2441,N_2462);
nand U2729 (N_2729,N_2452,N_2409);
or U2730 (N_2730,N_2282,N_2350);
xor U2731 (N_2731,N_2419,N_2471);
nor U2732 (N_2732,N_2482,N_2258);
nor U2733 (N_2733,N_2338,N_2399);
or U2734 (N_2734,N_2331,N_2498);
or U2735 (N_2735,N_2354,N_2395);
or U2736 (N_2736,N_2262,N_2349);
xnor U2737 (N_2737,N_2374,N_2496);
nor U2738 (N_2738,N_2260,N_2482);
xor U2739 (N_2739,N_2265,N_2351);
xor U2740 (N_2740,N_2279,N_2254);
or U2741 (N_2741,N_2307,N_2453);
or U2742 (N_2742,N_2366,N_2313);
and U2743 (N_2743,N_2349,N_2364);
nor U2744 (N_2744,N_2285,N_2418);
or U2745 (N_2745,N_2416,N_2367);
nand U2746 (N_2746,N_2264,N_2407);
and U2747 (N_2747,N_2422,N_2489);
nand U2748 (N_2748,N_2272,N_2417);
and U2749 (N_2749,N_2350,N_2312);
nand U2750 (N_2750,N_2677,N_2518);
or U2751 (N_2751,N_2532,N_2602);
or U2752 (N_2752,N_2684,N_2541);
or U2753 (N_2753,N_2556,N_2721);
and U2754 (N_2754,N_2698,N_2676);
nand U2755 (N_2755,N_2515,N_2617);
nor U2756 (N_2756,N_2507,N_2533);
nor U2757 (N_2757,N_2582,N_2585);
xnor U2758 (N_2758,N_2706,N_2718);
nor U2759 (N_2759,N_2600,N_2615);
and U2760 (N_2760,N_2563,N_2548);
nor U2761 (N_2761,N_2737,N_2635);
nand U2762 (N_2762,N_2566,N_2593);
nand U2763 (N_2763,N_2669,N_2517);
and U2764 (N_2764,N_2705,N_2579);
nand U2765 (N_2765,N_2661,N_2637);
or U2766 (N_2766,N_2643,N_2638);
or U2767 (N_2767,N_2622,N_2506);
nand U2768 (N_2768,N_2687,N_2731);
xor U2769 (N_2769,N_2512,N_2538);
nor U2770 (N_2770,N_2690,N_2630);
and U2771 (N_2771,N_2508,N_2722);
xnor U2772 (N_2772,N_2584,N_2658);
or U2773 (N_2773,N_2739,N_2636);
and U2774 (N_2774,N_2713,N_2699);
or U2775 (N_2775,N_2632,N_2589);
nor U2776 (N_2776,N_2645,N_2605);
nor U2777 (N_2777,N_2686,N_2730);
or U2778 (N_2778,N_2570,N_2604);
nand U2779 (N_2779,N_2609,N_2560);
and U2780 (N_2780,N_2550,N_2559);
nor U2781 (N_2781,N_2621,N_2552);
xnor U2782 (N_2782,N_2665,N_2704);
nor U2783 (N_2783,N_2514,N_2701);
and U2784 (N_2784,N_2598,N_2673);
or U2785 (N_2785,N_2539,N_2520);
and U2786 (N_2786,N_2640,N_2671);
xor U2787 (N_2787,N_2562,N_2743);
and U2788 (N_2788,N_2664,N_2742);
nand U2789 (N_2789,N_2537,N_2619);
nand U2790 (N_2790,N_2711,N_2714);
and U2791 (N_2791,N_2680,N_2736);
or U2792 (N_2792,N_2522,N_2688);
xor U2793 (N_2793,N_2513,N_2685);
and U2794 (N_2794,N_2555,N_2712);
nor U2795 (N_2795,N_2717,N_2702);
and U2796 (N_2796,N_2504,N_2573);
xnor U2797 (N_2797,N_2568,N_2709);
nand U2798 (N_2798,N_2672,N_2592);
and U2799 (N_2799,N_2576,N_2577);
xor U2800 (N_2800,N_2603,N_2564);
nor U2801 (N_2801,N_2614,N_2683);
or U2802 (N_2802,N_2659,N_2528);
or U2803 (N_2803,N_2728,N_2501);
or U2804 (N_2804,N_2639,N_2557);
or U2805 (N_2805,N_2623,N_2707);
and U2806 (N_2806,N_2525,N_2543);
nand U2807 (N_2807,N_2748,N_2625);
nand U2808 (N_2808,N_2653,N_2678);
nand U2809 (N_2809,N_2652,N_2608);
nand U2810 (N_2810,N_2535,N_2611);
nand U2811 (N_2811,N_2726,N_2667);
nand U2812 (N_2812,N_2547,N_2519);
and U2813 (N_2813,N_2629,N_2575);
and U2814 (N_2814,N_2590,N_2746);
nor U2815 (N_2815,N_2660,N_2542);
and U2816 (N_2816,N_2612,N_2580);
xnor U2817 (N_2817,N_2679,N_2516);
and U2818 (N_2818,N_2681,N_2618);
xor U2819 (N_2819,N_2654,N_2663);
and U2820 (N_2820,N_2620,N_2567);
and U2821 (N_2821,N_2733,N_2697);
xnor U2822 (N_2822,N_2628,N_2526);
nand U2823 (N_2823,N_2500,N_2720);
nand U2824 (N_2824,N_2633,N_2523);
xnor U2825 (N_2825,N_2641,N_2530);
or U2826 (N_2826,N_2583,N_2651);
and U2827 (N_2827,N_2723,N_2572);
nand U2828 (N_2828,N_2591,N_2505);
and U2829 (N_2829,N_2527,N_2536);
nor U2830 (N_2830,N_2646,N_2719);
nor U2831 (N_2831,N_2695,N_2627);
or U2832 (N_2832,N_2521,N_2740);
or U2833 (N_2833,N_2666,N_2700);
nor U2834 (N_2834,N_2553,N_2561);
and U2835 (N_2835,N_2509,N_2578);
or U2836 (N_2836,N_2696,N_2581);
nand U2837 (N_2837,N_2693,N_2544);
nand U2838 (N_2838,N_2574,N_2569);
nand U2839 (N_2839,N_2727,N_2747);
nor U2840 (N_2840,N_2503,N_2510);
or U2841 (N_2841,N_2644,N_2524);
xnor U2842 (N_2842,N_2708,N_2586);
and U2843 (N_2843,N_2655,N_2648);
nor U2844 (N_2844,N_2703,N_2682);
nand U2845 (N_2845,N_2545,N_2511);
nor U2846 (N_2846,N_2601,N_2670);
nor U2847 (N_2847,N_2694,N_2597);
or U2848 (N_2848,N_2626,N_2715);
and U2849 (N_2849,N_2571,N_2599);
nand U2850 (N_2850,N_2675,N_2546);
xor U2851 (N_2851,N_2657,N_2656);
and U2852 (N_2852,N_2551,N_2531);
and U2853 (N_2853,N_2624,N_2540);
or U2854 (N_2854,N_2725,N_2554);
nand U2855 (N_2855,N_2741,N_2565);
nand U2856 (N_2856,N_2502,N_2691);
and U2857 (N_2857,N_2749,N_2729);
nor U2858 (N_2858,N_2606,N_2734);
and U2859 (N_2859,N_2724,N_2745);
or U2860 (N_2860,N_2647,N_2650);
or U2861 (N_2861,N_2558,N_2631);
nor U2862 (N_2862,N_2689,N_2596);
nand U2863 (N_2863,N_2529,N_2668);
nand U2864 (N_2864,N_2674,N_2613);
and U2865 (N_2865,N_2549,N_2595);
or U2866 (N_2866,N_2607,N_2649);
xor U2867 (N_2867,N_2692,N_2616);
xnor U2868 (N_2868,N_2716,N_2732);
nor U2869 (N_2869,N_2534,N_2735);
nor U2870 (N_2870,N_2594,N_2587);
xnor U2871 (N_2871,N_2588,N_2642);
xor U2872 (N_2872,N_2710,N_2738);
xnor U2873 (N_2873,N_2610,N_2634);
or U2874 (N_2874,N_2662,N_2744);
xor U2875 (N_2875,N_2652,N_2667);
and U2876 (N_2876,N_2557,N_2665);
and U2877 (N_2877,N_2691,N_2570);
xor U2878 (N_2878,N_2678,N_2688);
nand U2879 (N_2879,N_2665,N_2598);
nor U2880 (N_2880,N_2502,N_2737);
nand U2881 (N_2881,N_2550,N_2558);
nand U2882 (N_2882,N_2644,N_2603);
or U2883 (N_2883,N_2502,N_2728);
or U2884 (N_2884,N_2677,N_2546);
xor U2885 (N_2885,N_2556,N_2684);
and U2886 (N_2886,N_2640,N_2608);
or U2887 (N_2887,N_2514,N_2726);
and U2888 (N_2888,N_2554,N_2719);
nand U2889 (N_2889,N_2668,N_2503);
and U2890 (N_2890,N_2641,N_2637);
xnor U2891 (N_2891,N_2529,N_2558);
nand U2892 (N_2892,N_2535,N_2701);
and U2893 (N_2893,N_2732,N_2560);
or U2894 (N_2894,N_2547,N_2539);
or U2895 (N_2895,N_2550,N_2681);
nand U2896 (N_2896,N_2703,N_2670);
nand U2897 (N_2897,N_2523,N_2682);
or U2898 (N_2898,N_2508,N_2569);
nand U2899 (N_2899,N_2549,N_2618);
nor U2900 (N_2900,N_2645,N_2655);
xnor U2901 (N_2901,N_2681,N_2515);
nand U2902 (N_2902,N_2721,N_2660);
nand U2903 (N_2903,N_2634,N_2691);
and U2904 (N_2904,N_2505,N_2657);
and U2905 (N_2905,N_2557,N_2574);
or U2906 (N_2906,N_2575,N_2624);
nand U2907 (N_2907,N_2552,N_2643);
and U2908 (N_2908,N_2611,N_2703);
and U2909 (N_2909,N_2502,N_2538);
nand U2910 (N_2910,N_2635,N_2552);
or U2911 (N_2911,N_2517,N_2728);
xor U2912 (N_2912,N_2706,N_2606);
xor U2913 (N_2913,N_2628,N_2623);
nand U2914 (N_2914,N_2717,N_2520);
xor U2915 (N_2915,N_2503,N_2644);
xnor U2916 (N_2916,N_2565,N_2526);
nor U2917 (N_2917,N_2662,N_2518);
nand U2918 (N_2918,N_2504,N_2506);
nand U2919 (N_2919,N_2658,N_2655);
or U2920 (N_2920,N_2520,N_2738);
and U2921 (N_2921,N_2514,N_2563);
or U2922 (N_2922,N_2729,N_2662);
xnor U2923 (N_2923,N_2592,N_2681);
nor U2924 (N_2924,N_2638,N_2547);
nor U2925 (N_2925,N_2594,N_2668);
nand U2926 (N_2926,N_2724,N_2579);
xnor U2927 (N_2927,N_2577,N_2694);
nand U2928 (N_2928,N_2670,N_2534);
and U2929 (N_2929,N_2694,N_2697);
and U2930 (N_2930,N_2735,N_2561);
nand U2931 (N_2931,N_2713,N_2617);
and U2932 (N_2932,N_2668,N_2703);
nand U2933 (N_2933,N_2647,N_2504);
and U2934 (N_2934,N_2561,N_2513);
nand U2935 (N_2935,N_2713,N_2625);
nand U2936 (N_2936,N_2534,N_2629);
and U2937 (N_2937,N_2732,N_2584);
nor U2938 (N_2938,N_2587,N_2584);
xnor U2939 (N_2939,N_2720,N_2738);
nand U2940 (N_2940,N_2550,N_2557);
nor U2941 (N_2941,N_2645,N_2611);
or U2942 (N_2942,N_2653,N_2688);
nand U2943 (N_2943,N_2728,N_2716);
or U2944 (N_2944,N_2736,N_2735);
nand U2945 (N_2945,N_2518,N_2652);
nand U2946 (N_2946,N_2615,N_2691);
nand U2947 (N_2947,N_2621,N_2632);
nand U2948 (N_2948,N_2664,N_2707);
or U2949 (N_2949,N_2502,N_2577);
or U2950 (N_2950,N_2617,N_2627);
nor U2951 (N_2951,N_2693,N_2723);
or U2952 (N_2952,N_2587,N_2655);
nor U2953 (N_2953,N_2541,N_2542);
and U2954 (N_2954,N_2618,N_2564);
nand U2955 (N_2955,N_2591,N_2536);
nand U2956 (N_2956,N_2730,N_2742);
nand U2957 (N_2957,N_2721,N_2509);
xor U2958 (N_2958,N_2561,N_2504);
nand U2959 (N_2959,N_2573,N_2727);
xnor U2960 (N_2960,N_2546,N_2548);
xor U2961 (N_2961,N_2699,N_2591);
xor U2962 (N_2962,N_2748,N_2566);
xor U2963 (N_2963,N_2673,N_2679);
xnor U2964 (N_2964,N_2684,N_2713);
nand U2965 (N_2965,N_2609,N_2557);
or U2966 (N_2966,N_2514,N_2548);
and U2967 (N_2967,N_2645,N_2648);
nor U2968 (N_2968,N_2607,N_2532);
nand U2969 (N_2969,N_2645,N_2530);
and U2970 (N_2970,N_2636,N_2542);
nand U2971 (N_2971,N_2718,N_2705);
and U2972 (N_2972,N_2694,N_2711);
nor U2973 (N_2973,N_2600,N_2714);
xor U2974 (N_2974,N_2657,N_2551);
and U2975 (N_2975,N_2522,N_2728);
nand U2976 (N_2976,N_2536,N_2511);
or U2977 (N_2977,N_2662,N_2686);
and U2978 (N_2978,N_2741,N_2595);
xor U2979 (N_2979,N_2576,N_2527);
nor U2980 (N_2980,N_2738,N_2641);
nand U2981 (N_2981,N_2559,N_2573);
nand U2982 (N_2982,N_2552,N_2564);
and U2983 (N_2983,N_2742,N_2557);
nor U2984 (N_2984,N_2562,N_2731);
or U2985 (N_2985,N_2730,N_2729);
xnor U2986 (N_2986,N_2647,N_2673);
nand U2987 (N_2987,N_2639,N_2672);
and U2988 (N_2988,N_2570,N_2535);
or U2989 (N_2989,N_2501,N_2608);
nand U2990 (N_2990,N_2586,N_2640);
nand U2991 (N_2991,N_2561,N_2682);
xor U2992 (N_2992,N_2693,N_2608);
xnor U2993 (N_2993,N_2512,N_2565);
nor U2994 (N_2994,N_2676,N_2580);
nand U2995 (N_2995,N_2611,N_2738);
and U2996 (N_2996,N_2501,N_2552);
nand U2997 (N_2997,N_2689,N_2675);
nand U2998 (N_2998,N_2551,N_2708);
nor U2999 (N_2999,N_2589,N_2749);
xnor U3000 (N_3000,N_2828,N_2897);
nor U3001 (N_3001,N_2776,N_2868);
or U3002 (N_3002,N_2975,N_2819);
nand U3003 (N_3003,N_2851,N_2763);
or U3004 (N_3004,N_2931,N_2770);
xor U3005 (N_3005,N_2905,N_2944);
or U3006 (N_3006,N_2854,N_2938);
xnor U3007 (N_3007,N_2812,N_2907);
or U3008 (N_3008,N_2987,N_2867);
or U3009 (N_3009,N_2857,N_2864);
nand U3010 (N_3010,N_2875,N_2895);
xor U3011 (N_3011,N_2943,N_2872);
xnor U3012 (N_3012,N_2996,N_2818);
xnor U3013 (N_3013,N_2891,N_2824);
or U3014 (N_3014,N_2984,N_2928);
nand U3015 (N_3015,N_2848,N_2758);
xnor U3016 (N_3016,N_2925,N_2752);
and U3017 (N_3017,N_2783,N_2918);
xnor U3018 (N_3018,N_2871,N_2821);
or U3019 (N_3019,N_2795,N_2835);
nand U3020 (N_3020,N_2954,N_2865);
nand U3021 (N_3021,N_2849,N_2986);
or U3022 (N_3022,N_2947,N_2978);
nand U3023 (N_3023,N_2760,N_2814);
nand U3024 (N_3024,N_2946,N_2870);
and U3025 (N_3025,N_2962,N_2908);
nand U3026 (N_3026,N_2993,N_2959);
nor U3027 (N_3027,N_2941,N_2757);
nand U3028 (N_3028,N_2764,N_2916);
nand U3029 (N_3029,N_2973,N_2945);
or U3030 (N_3030,N_2919,N_2934);
xnor U3031 (N_3031,N_2898,N_2989);
and U3032 (N_3032,N_2904,N_2914);
xor U3033 (N_3033,N_2968,N_2917);
nand U3034 (N_3034,N_2811,N_2920);
xnor U3035 (N_3035,N_2910,N_2964);
and U3036 (N_3036,N_2772,N_2892);
or U3037 (N_3037,N_2789,N_2785);
nor U3038 (N_3038,N_2886,N_2845);
xor U3039 (N_3039,N_2823,N_2970);
and U3040 (N_3040,N_2782,N_2999);
xnor U3041 (N_3041,N_2903,N_2769);
nand U3042 (N_3042,N_2957,N_2827);
or U3043 (N_3043,N_2816,N_2784);
nor U3044 (N_3044,N_2939,N_2915);
nor U3045 (N_3045,N_2882,N_2767);
xor U3046 (N_3046,N_2974,N_2877);
and U3047 (N_3047,N_2836,N_2766);
nand U3048 (N_3048,N_2806,N_2759);
nand U3049 (N_3049,N_2900,N_2817);
or U3050 (N_3050,N_2955,N_2929);
nor U3051 (N_3051,N_2977,N_2774);
nor U3052 (N_3052,N_2949,N_2855);
nor U3053 (N_3053,N_2873,N_2804);
and U3054 (N_3054,N_2860,N_2801);
and U3055 (N_3055,N_2762,N_2988);
or U3056 (N_3056,N_2960,N_2768);
nand U3057 (N_3057,N_2899,N_2952);
nand U3058 (N_3058,N_2820,N_2844);
nor U3059 (N_3059,N_2961,N_2888);
or U3060 (N_3060,N_2884,N_2756);
or U3061 (N_3061,N_2972,N_2951);
xnor U3062 (N_3062,N_2771,N_2994);
nor U3063 (N_3063,N_2901,N_2773);
and U3064 (N_3064,N_2885,N_2825);
nand U3065 (N_3065,N_2859,N_2788);
and U3066 (N_3066,N_2921,N_2803);
xor U3067 (N_3067,N_2927,N_2936);
nand U3068 (N_3068,N_2922,N_2981);
nor U3069 (N_3069,N_2995,N_2781);
and U3070 (N_3070,N_2894,N_2858);
nand U3071 (N_3071,N_2850,N_2982);
or U3072 (N_3072,N_2880,N_2753);
nand U3073 (N_3073,N_2805,N_2976);
nor U3074 (N_3074,N_2826,N_2791);
nor U3075 (N_3075,N_2906,N_2798);
xnor U3076 (N_3076,N_2809,N_2846);
nand U3077 (N_3077,N_2775,N_2793);
nor U3078 (N_3078,N_2940,N_2985);
and U3079 (N_3079,N_2778,N_2800);
xor U3080 (N_3080,N_2832,N_2862);
or U3081 (N_3081,N_2790,N_2998);
or U3082 (N_3082,N_2843,N_2869);
nor U3083 (N_3083,N_2822,N_2966);
or U3084 (N_3084,N_2815,N_2958);
nand U3085 (N_3085,N_2983,N_2847);
nand U3086 (N_3086,N_2889,N_2838);
or U3087 (N_3087,N_2937,N_2794);
nand U3088 (N_3088,N_2874,N_2878);
and U3089 (N_3089,N_2924,N_2786);
nor U3090 (N_3090,N_2950,N_2853);
or U3091 (N_3091,N_2979,N_2840);
xor U3092 (N_3092,N_2953,N_2807);
xor U3093 (N_3093,N_2881,N_2755);
xnor U3094 (N_3094,N_2969,N_2799);
nor U3095 (N_3095,N_2956,N_2810);
or U3096 (N_3096,N_2856,N_2852);
nand U3097 (N_3097,N_2893,N_2909);
and U3098 (N_3098,N_2887,N_2933);
xor U3099 (N_3099,N_2842,N_2765);
xor U3100 (N_3100,N_2750,N_2813);
xnor U3101 (N_3101,N_2890,N_2839);
or U3102 (N_3102,N_2935,N_2792);
nand U3103 (N_3103,N_2780,N_2883);
and U3104 (N_3104,N_2808,N_2997);
xnor U3105 (N_3105,N_2896,N_2930);
nand U3106 (N_3106,N_2963,N_2992);
or U3107 (N_3107,N_2990,N_2829);
xor U3108 (N_3108,N_2923,N_2902);
xnor U3109 (N_3109,N_2967,N_2754);
and U3110 (N_3110,N_2802,N_2833);
or U3111 (N_3111,N_2911,N_2779);
nor U3112 (N_3112,N_2797,N_2866);
and U3113 (N_3113,N_2761,N_2926);
nor U3114 (N_3114,N_2841,N_2980);
or U3115 (N_3115,N_2912,N_2863);
and U3116 (N_3116,N_2942,N_2837);
xor U3117 (N_3117,N_2965,N_2796);
nand U3118 (N_3118,N_2751,N_2932);
or U3119 (N_3119,N_2948,N_2834);
xnor U3120 (N_3120,N_2787,N_2777);
and U3121 (N_3121,N_2830,N_2831);
or U3122 (N_3122,N_2991,N_2861);
nand U3123 (N_3123,N_2913,N_2876);
xor U3124 (N_3124,N_2879,N_2971);
nand U3125 (N_3125,N_2897,N_2753);
nand U3126 (N_3126,N_2770,N_2862);
and U3127 (N_3127,N_2765,N_2854);
and U3128 (N_3128,N_2838,N_2804);
xnor U3129 (N_3129,N_2759,N_2907);
xor U3130 (N_3130,N_2993,N_2997);
and U3131 (N_3131,N_2819,N_2942);
xnor U3132 (N_3132,N_2981,N_2908);
xor U3133 (N_3133,N_2867,N_2994);
and U3134 (N_3134,N_2890,N_2779);
and U3135 (N_3135,N_2978,N_2864);
xor U3136 (N_3136,N_2997,N_2856);
or U3137 (N_3137,N_2808,N_2929);
nand U3138 (N_3138,N_2915,N_2837);
xor U3139 (N_3139,N_2752,N_2950);
nor U3140 (N_3140,N_2792,N_2807);
nand U3141 (N_3141,N_2871,N_2986);
or U3142 (N_3142,N_2795,N_2811);
nor U3143 (N_3143,N_2915,N_2929);
and U3144 (N_3144,N_2785,N_2919);
xor U3145 (N_3145,N_2883,N_2925);
or U3146 (N_3146,N_2985,N_2804);
and U3147 (N_3147,N_2897,N_2756);
and U3148 (N_3148,N_2899,N_2951);
and U3149 (N_3149,N_2800,N_2950);
nor U3150 (N_3150,N_2838,N_2910);
nor U3151 (N_3151,N_2817,N_2845);
nor U3152 (N_3152,N_2804,N_2881);
nor U3153 (N_3153,N_2998,N_2807);
nor U3154 (N_3154,N_2895,N_2826);
nor U3155 (N_3155,N_2772,N_2886);
or U3156 (N_3156,N_2827,N_2940);
xor U3157 (N_3157,N_2870,N_2907);
nand U3158 (N_3158,N_2892,N_2846);
xor U3159 (N_3159,N_2986,N_2829);
or U3160 (N_3160,N_2833,N_2950);
nor U3161 (N_3161,N_2945,N_2851);
xor U3162 (N_3162,N_2787,N_2945);
nand U3163 (N_3163,N_2782,N_2829);
and U3164 (N_3164,N_2908,N_2992);
or U3165 (N_3165,N_2989,N_2976);
nor U3166 (N_3166,N_2887,N_2846);
nand U3167 (N_3167,N_2851,N_2777);
nand U3168 (N_3168,N_2890,N_2986);
nor U3169 (N_3169,N_2794,N_2960);
nand U3170 (N_3170,N_2887,N_2818);
or U3171 (N_3171,N_2875,N_2857);
xnor U3172 (N_3172,N_2837,N_2918);
nor U3173 (N_3173,N_2915,N_2769);
nor U3174 (N_3174,N_2823,N_2816);
nand U3175 (N_3175,N_2931,N_2833);
nor U3176 (N_3176,N_2885,N_2765);
nor U3177 (N_3177,N_2935,N_2910);
nor U3178 (N_3178,N_2933,N_2915);
xnor U3179 (N_3179,N_2878,N_2998);
nand U3180 (N_3180,N_2998,N_2769);
xor U3181 (N_3181,N_2955,N_2857);
xor U3182 (N_3182,N_2992,N_2757);
or U3183 (N_3183,N_2771,N_2836);
nand U3184 (N_3184,N_2773,N_2940);
nand U3185 (N_3185,N_2779,N_2910);
and U3186 (N_3186,N_2825,N_2886);
nand U3187 (N_3187,N_2881,N_2999);
nand U3188 (N_3188,N_2889,N_2950);
nor U3189 (N_3189,N_2830,N_2856);
xor U3190 (N_3190,N_2971,N_2926);
xnor U3191 (N_3191,N_2880,N_2950);
nor U3192 (N_3192,N_2876,N_2947);
nor U3193 (N_3193,N_2928,N_2978);
nor U3194 (N_3194,N_2808,N_2824);
nand U3195 (N_3195,N_2781,N_2773);
and U3196 (N_3196,N_2948,N_2813);
nand U3197 (N_3197,N_2823,N_2812);
or U3198 (N_3198,N_2760,N_2813);
and U3199 (N_3199,N_2917,N_2873);
nand U3200 (N_3200,N_2837,N_2768);
xor U3201 (N_3201,N_2847,N_2932);
xnor U3202 (N_3202,N_2950,N_2844);
xor U3203 (N_3203,N_2888,N_2924);
nor U3204 (N_3204,N_2781,N_2760);
nand U3205 (N_3205,N_2813,N_2905);
and U3206 (N_3206,N_2880,N_2837);
nand U3207 (N_3207,N_2883,N_2870);
xor U3208 (N_3208,N_2853,N_2868);
xnor U3209 (N_3209,N_2954,N_2909);
nand U3210 (N_3210,N_2805,N_2966);
and U3211 (N_3211,N_2888,N_2894);
nand U3212 (N_3212,N_2923,N_2808);
xnor U3213 (N_3213,N_2921,N_2836);
and U3214 (N_3214,N_2909,N_2784);
nand U3215 (N_3215,N_2945,N_2760);
and U3216 (N_3216,N_2909,N_2925);
nor U3217 (N_3217,N_2824,N_2817);
or U3218 (N_3218,N_2872,N_2754);
or U3219 (N_3219,N_2980,N_2797);
and U3220 (N_3220,N_2760,N_2983);
xnor U3221 (N_3221,N_2779,N_2880);
and U3222 (N_3222,N_2941,N_2852);
or U3223 (N_3223,N_2924,N_2918);
nand U3224 (N_3224,N_2943,N_2966);
nor U3225 (N_3225,N_2894,N_2972);
xor U3226 (N_3226,N_2824,N_2983);
xor U3227 (N_3227,N_2750,N_2834);
nand U3228 (N_3228,N_2931,N_2914);
nor U3229 (N_3229,N_2969,N_2759);
nand U3230 (N_3230,N_2945,N_2772);
nand U3231 (N_3231,N_2953,N_2832);
nand U3232 (N_3232,N_2878,N_2938);
nand U3233 (N_3233,N_2837,N_2813);
nand U3234 (N_3234,N_2928,N_2956);
and U3235 (N_3235,N_2788,N_2762);
and U3236 (N_3236,N_2798,N_2802);
xnor U3237 (N_3237,N_2860,N_2971);
xor U3238 (N_3238,N_2930,N_2981);
xor U3239 (N_3239,N_2752,N_2890);
and U3240 (N_3240,N_2880,N_2913);
or U3241 (N_3241,N_2768,N_2926);
or U3242 (N_3242,N_2770,N_2919);
nor U3243 (N_3243,N_2956,N_2921);
or U3244 (N_3244,N_2861,N_2951);
nor U3245 (N_3245,N_2985,N_2980);
nand U3246 (N_3246,N_2950,N_2904);
nor U3247 (N_3247,N_2967,N_2828);
nor U3248 (N_3248,N_2824,N_2996);
nor U3249 (N_3249,N_2981,N_2822);
xnor U3250 (N_3250,N_3241,N_3188);
or U3251 (N_3251,N_3039,N_3162);
and U3252 (N_3252,N_3075,N_3036);
xor U3253 (N_3253,N_3115,N_3072);
or U3254 (N_3254,N_3144,N_3041);
xnor U3255 (N_3255,N_3062,N_3027);
xor U3256 (N_3256,N_3223,N_3086);
xor U3257 (N_3257,N_3205,N_3110);
and U3258 (N_3258,N_3228,N_3201);
or U3259 (N_3259,N_3200,N_3180);
nand U3260 (N_3260,N_3168,N_3203);
or U3261 (N_3261,N_3038,N_3147);
or U3262 (N_3262,N_3129,N_3152);
or U3263 (N_3263,N_3211,N_3149);
xor U3264 (N_3264,N_3239,N_3021);
nor U3265 (N_3265,N_3113,N_3237);
or U3266 (N_3266,N_3068,N_3190);
and U3267 (N_3267,N_3109,N_3153);
nand U3268 (N_3268,N_3159,N_3081);
nand U3269 (N_3269,N_3161,N_3225);
nand U3270 (N_3270,N_3032,N_3163);
or U3271 (N_3271,N_3112,N_3236);
xor U3272 (N_3272,N_3215,N_3006);
nor U3273 (N_3273,N_3216,N_3126);
nand U3274 (N_3274,N_3091,N_3146);
nand U3275 (N_3275,N_3060,N_3092);
and U3276 (N_3276,N_3076,N_3231);
nand U3277 (N_3277,N_3071,N_3196);
xnor U3278 (N_3278,N_3151,N_3098);
or U3279 (N_3279,N_3234,N_3247);
and U3280 (N_3280,N_3089,N_3170);
xnor U3281 (N_3281,N_3002,N_3173);
xor U3282 (N_3282,N_3179,N_3244);
or U3283 (N_3283,N_3059,N_3212);
nand U3284 (N_3284,N_3045,N_3087);
or U3285 (N_3285,N_3101,N_3130);
nor U3286 (N_3286,N_3198,N_3171);
xnor U3287 (N_3287,N_3095,N_3116);
and U3288 (N_3288,N_3028,N_3033);
and U3289 (N_3289,N_3169,N_3102);
or U3290 (N_3290,N_3233,N_3174);
nor U3291 (N_3291,N_3016,N_3013);
nand U3292 (N_3292,N_3084,N_3105);
or U3293 (N_3293,N_3066,N_3132);
or U3294 (N_3294,N_3030,N_3053);
nand U3295 (N_3295,N_3048,N_3154);
nor U3296 (N_3296,N_3108,N_3145);
and U3297 (N_3297,N_3097,N_3056);
or U3298 (N_3298,N_3150,N_3083);
or U3299 (N_3299,N_3227,N_3243);
nor U3300 (N_3300,N_3090,N_3121);
xor U3301 (N_3301,N_3000,N_3197);
xnor U3302 (N_3302,N_3015,N_3235);
or U3303 (N_3303,N_3044,N_3177);
and U3304 (N_3304,N_3019,N_3049);
xnor U3305 (N_3305,N_3052,N_3057);
and U3306 (N_3306,N_3106,N_3224);
nand U3307 (N_3307,N_3134,N_3183);
nand U3308 (N_3308,N_3080,N_3008);
or U3309 (N_3309,N_3073,N_3140);
and U3310 (N_3310,N_3131,N_3001);
nor U3311 (N_3311,N_3047,N_3054);
nand U3312 (N_3312,N_3158,N_3012);
nand U3313 (N_3313,N_3208,N_3156);
or U3314 (N_3314,N_3128,N_3202);
or U3315 (N_3315,N_3164,N_3182);
nand U3316 (N_3316,N_3166,N_3245);
and U3317 (N_3317,N_3118,N_3242);
nand U3318 (N_3318,N_3031,N_3069);
or U3319 (N_3319,N_3024,N_3037);
nor U3320 (N_3320,N_3005,N_3014);
xor U3321 (N_3321,N_3194,N_3042);
and U3322 (N_3322,N_3067,N_3219);
or U3323 (N_3323,N_3077,N_3155);
and U3324 (N_3324,N_3018,N_3122);
nor U3325 (N_3325,N_3046,N_3240);
xnor U3326 (N_3326,N_3074,N_3213);
and U3327 (N_3327,N_3230,N_3022);
and U3328 (N_3328,N_3193,N_3085);
xnor U3329 (N_3329,N_3189,N_3204);
nor U3330 (N_3330,N_3160,N_3186);
and U3331 (N_3331,N_3093,N_3139);
nand U3332 (N_3332,N_3172,N_3133);
or U3333 (N_3333,N_3127,N_3111);
nor U3334 (N_3334,N_3079,N_3207);
or U3335 (N_3335,N_3020,N_3209);
nand U3336 (N_3336,N_3026,N_3232);
nor U3337 (N_3337,N_3119,N_3023);
nor U3338 (N_3338,N_3229,N_3055);
nor U3339 (N_3339,N_3103,N_3218);
or U3340 (N_3340,N_3199,N_3120);
nand U3341 (N_3341,N_3061,N_3010);
xor U3342 (N_3342,N_3070,N_3249);
nor U3343 (N_3343,N_3003,N_3078);
and U3344 (N_3344,N_3191,N_3124);
and U3345 (N_3345,N_3167,N_3043);
xnor U3346 (N_3346,N_3136,N_3226);
xnor U3347 (N_3347,N_3148,N_3135);
nor U3348 (N_3348,N_3157,N_3187);
and U3349 (N_3349,N_3175,N_3104);
and U3350 (N_3350,N_3063,N_3206);
xor U3351 (N_3351,N_3246,N_3050);
nor U3352 (N_3352,N_3137,N_3222);
nand U3353 (N_3353,N_3125,N_3096);
nor U3354 (N_3354,N_3178,N_3248);
nand U3355 (N_3355,N_3107,N_3114);
nor U3356 (N_3356,N_3029,N_3035);
nor U3357 (N_3357,N_3195,N_3123);
and U3358 (N_3358,N_3138,N_3181);
or U3359 (N_3359,N_3088,N_3184);
xnor U3360 (N_3360,N_3165,N_3176);
nand U3361 (N_3361,N_3217,N_3221);
and U3362 (N_3362,N_3214,N_3117);
nor U3363 (N_3363,N_3210,N_3034);
nand U3364 (N_3364,N_3051,N_3011);
xnor U3365 (N_3365,N_3238,N_3040);
nor U3366 (N_3366,N_3094,N_3192);
and U3367 (N_3367,N_3007,N_3099);
nand U3368 (N_3368,N_3004,N_3017);
nand U3369 (N_3369,N_3025,N_3065);
nor U3370 (N_3370,N_3141,N_3058);
xor U3371 (N_3371,N_3142,N_3009);
xor U3372 (N_3372,N_3220,N_3064);
nor U3373 (N_3373,N_3143,N_3082);
nand U3374 (N_3374,N_3100,N_3185);
nor U3375 (N_3375,N_3138,N_3043);
and U3376 (N_3376,N_3039,N_3114);
and U3377 (N_3377,N_3005,N_3079);
nor U3378 (N_3378,N_3193,N_3131);
nand U3379 (N_3379,N_3006,N_3086);
nand U3380 (N_3380,N_3142,N_3173);
nor U3381 (N_3381,N_3076,N_3050);
nor U3382 (N_3382,N_3197,N_3176);
nor U3383 (N_3383,N_3102,N_3149);
nor U3384 (N_3384,N_3194,N_3226);
or U3385 (N_3385,N_3139,N_3087);
and U3386 (N_3386,N_3019,N_3178);
xor U3387 (N_3387,N_3097,N_3103);
nand U3388 (N_3388,N_3085,N_3126);
and U3389 (N_3389,N_3068,N_3159);
nor U3390 (N_3390,N_3053,N_3050);
xor U3391 (N_3391,N_3115,N_3000);
and U3392 (N_3392,N_3188,N_3189);
or U3393 (N_3393,N_3012,N_3110);
and U3394 (N_3394,N_3231,N_3186);
and U3395 (N_3395,N_3123,N_3055);
or U3396 (N_3396,N_3079,N_3046);
nand U3397 (N_3397,N_3004,N_3050);
nand U3398 (N_3398,N_3222,N_3159);
and U3399 (N_3399,N_3186,N_3243);
nand U3400 (N_3400,N_3091,N_3237);
nor U3401 (N_3401,N_3188,N_3069);
nor U3402 (N_3402,N_3029,N_3212);
or U3403 (N_3403,N_3124,N_3155);
nand U3404 (N_3404,N_3018,N_3082);
nor U3405 (N_3405,N_3159,N_3212);
xor U3406 (N_3406,N_3086,N_3049);
nor U3407 (N_3407,N_3104,N_3102);
nor U3408 (N_3408,N_3044,N_3010);
nand U3409 (N_3409,N_3096,N_3181);
xor U3410 (N_3410,N_3141,N_3244);
nand U3411 (N_3411,N_3204,N_3003);
and U3412 (N_3412,N_3247,N_3081);
xnor U3413 (N_3413,N_3179,N_3192);
xor U3414 (N_3414,N_3072,N_3143);
or U3415 (N_3415,N_3060,N_3175);
and U3416 (N_3416,N_3118,N_3170);
nor U3417 (N_3417,N_3077,N_3194);
or U3418 (N_3418,N_3010,N_3213);
and U3419 (N_3419,N_3128,N_3026);
xnor U3420 (N_3420,N_3230,N_3200);
and U3421 (N_3421,N_3012,N_3169);
nor U3422 (N_3422,N_3217,N_3175);
xnor U3423 (N_3423,N_3210,N_3083);
xor U3424 (N_3424,N_3193,N_3125);
and U3425 (N_3425,N_3077,N_3172);
or U3426 (N_3426,N_3112,N_3162);
and U3427 (N_3427,N_3043,N_3075);
nand U3428 (N_3428,N_3057,N_3037);
nor U3429 (N_3429,N_3168,N_3130);
or U3430 (N_3430,N_3226,N_3212);
or U3431 (N_3431,N_3107,N_3057);
and U3432 (N_3432,N_3230,N_3126);
nor U3433 (N_3433,N_3130,N_3036);
or U3434 (N_3434,N_3051,N_3164);
xor U3435 (N_3435,N_3213,N_3050);
nor U3436 (N_3436,N_3080,N_3039);
or U3437 (N_3437,N_3202,N_3233);
nor U3438 (N_3438,N_3118,N_3214);
nand U3439 (N_3439,N_3008,N_3205);
or U3440 (N_3440,N_3203,N_3034);
nor U3441 (N_3441,N_3239,N_3164);
or U3442 (N_3442,N_3227,N_3031);
nor U3443 (N_3443,N_3002,N_3199);
nand U3444 (N_3444,N_3004,N_3104);
nand U3445 (N_3445,N_3103,N_3066);
xor U3446 (N_3446,N_3090,N_3036);
nor U3447 (N_3447,N_3063,N_3174);
nand U3448 (N_3448,N_3008,N_3216);
xnor U3449 (N_3449,N_3153,N_3106);
nor U3450 (N_3450,N_3022,N_3056);
xnor U3451 (N_3451,N_3003,N_3035);
xnor U3452 (N_3452,N_3138,N_3045);
nor U3453 (N_3453,N_3028,N_3088);
nand U3454 (N_3454,N_3159,N_3045);
and U3455 (N_3455,N_3238,N_3114);
nand U3456 (N_3456,N_3026,N_3049);
and U3457 (N_3457,N_3064,N_3083);
nand U3458 (N_3458,N_3049,N_3152);
and U3459 (N_3459,N_3105,N_3003);
and U3460 (N_3460,N_3138,N_3063);
xnor U3461 (N_3461,N_3041,N_3018);
and U3462 (N_3462,N_3197,N_3241);
xnor U3463 (N_3463,N_3227,N_3024);
nor U3464 (N_3464,N_3062,N_3215);
nor U3465 (N_3465,N_3108,N_3085);
xnor U3466 (N_3466,N_3107,N_3167);
xnor U3467 (N_3467,N_3208,N_3139);
nand U3468 (N_3468,N_3166,N_3065);
xnor U3469 (N_3469,N_3161,N_3230);
xnor U3470 (N_3470,N_3181,N_3132);
xor U3471 (N_3471,N_3048,N_3168);
xnor U3472 (N_3472,N_3023,N_3184);
nor U3473 (N_3473,N_3231,N_3148);
and U3474 (N_3474,N_3166,N_3226);
and U3475 (N_3475,N_3172,N_3225);
or U3476 (N_3476,N_3196,N_3123);
and U3477 (N_3477,N_3191,N_3178);
xnor U3478 (N_3478,N_3202,N_3243);
nor U3479 (N_3479,N_3218,N_3112);
nand U3480 (N_3480,N_3193,N_3212);
and U3481 (N_3481,N_3040,N_3192);
nand U3482 (N_3482,N_3183,N_3062);
nor U3483 (N_3483,N_3179,N_3177);
xnor U3484 (N_3484,N_3067,N_3101);
nor U3485 (N_3485,N_3021,N_3047);
and U3486 (N_3486,N_3059,N_3104);
and U3487 (N_3487,N_3184,N_3094);
or U3488 (N_3488,N_3125,N_3030);
or U3489 (N_3489,N_3148,N_3056);
xor U3490 (N_3490,N_3141,N_3153);
nand U3491 (N_3491,N_3089,N_3194);
nor U3492 (N_3492,N_3008,N_3159);
nor U3493 (N_3493,N_3015,N_3171);
nor U3494 (N_3494,N_3172,N_3014);
nor U3495 (N_3495,N_3117,N_3215);
nand U3496 (N_3496,N_3040,N_3128);
nor U3497 (N_3497,N_3121,N_3176);
nor U3498 (N_3498,N_3184,N_3177);
and U3499 (N_3499,N_3035,N_3019);
nor U3500 (N_3500,N_3421,N_3490);
xor U3501 (N_3501,N_3491,N_3371);
xor U3502 (N_3502,N_3300,N_3486);
and U3503 (N_3503,N_3348,N_3352);
or U3504 (N_3504,N_3426,N_3487);
and U3505 (N_3505,N_3461,N_3329);
nand U3506 (N_3506,N_3281,N_3435);
xor U3507 (N_3507,N_3287,N_3289);
and U3508 (N_3508,N_3332,N_3375);
and U3509 (N_3509,N_3390,N_3312);
or U3510 (N_3510,N_3481,N_3358);
nand U3511 (N_3511,N_3293,N_3464);
and U3512 (N_3512,N_3389,N_3456);
and U3513 (N_3513,N_3410,N_3424);
or U3514 (N_3514,N_3369,N_3261);
nand U3515 (N_3515,N_3394,N_3498);
nor U3516 (N_3516,N_3323,N_3460);
xor U3517 (N_3517,N_3342,N_3473);
nand U3518 (N_3518,N_3262,N_3445);
and U3519 (N_3519,N_3429,N_3275);
and U3520 (N_3520,N_3427,N_3434);
and U3521 (N_3521,N_3299,N_3260);
nor U3522 (N_3522,N_3320,N_3319);
or U3523 (N_3523,N_3428,N_3471);
and U3524 (N_3524,N_3399,N_3422);
nor U3525 (N_3525,N_3310,N_3432);
xnor U3526 (N_3526,N_3452,N_3376);
nor U3527 (N_3527,N_3340,N_3370);
xnor U3528 (N_3528,N_3356,N_3400);
nand U3529 (N_3529,N_3386,N_3318);
nand U3530 (N_3530,N_3405,N_3465);
nand U3531 (N_3531,N_3387,N_3349);
and U3532 (N_3532,N_3475,N_3493);
nor U3533 (N_3533,N_3457,N_3447);
xor U3534 (N_3534,N_3333,N_3357);
xnor U3535 (N_3535,N_3346,N_3401);
or U3536 (N_3536,N_3309,N_3413);
nand U3537 (N_3537,N_3302,N_3466);
and U3538 (N_3538,N_3360,N_3344);
nor U3539 (N_3539,N_3336,N_3458);
nand U3540 (N_3540,N_3315,N_3367);
nand U3541 (N_3541,N_3363,N_3317);
xor U3542 (N_3542,N_3290,N_3303);
nand U3543 (N_3543,N_3372,N_3451);
and U3544 (N_3544,N_3269,N_3404);
nor U3545 (N_3545,N_3377,N_3362);
xnor U3546 (N_3546,N_3469,N_3325);
nor U3547 (N_3547,N_3252,N_3392);
or U3548 (N_3548,N_3365,N_3297);
and U3549 (N_3549,N_3316,N_3470);
or U3550 (N_3550,N_3418,N_3304);
nor U3551 (N_3551,N_3483,N_3351);
or U3552 (N_3552,N_3272,N_3384);
or U3553 (N_3553,N_3324,N_3436);
and U3554 (N_3554,N_3288,N_3301);
nand U3555 (N_3555,N_3373,N_3326);
nor U3556 (N_3556,N_3431,N_3391);
or U3557 (N_3557,N_3403,N_3414);
or U3558 (N_3558,N_3257,N_3472);
xnor U3559 (N_3559,N_3485,N_3368);
or U3560 (N_3560,N_3379,N_3468);
xor U3561 (N_3561,N_3415,N_3416);
nand U3562 (N_3562,N_3495,N_3321);
or U3563 (N_3563,N_3296,N_3378);
or U3564 (N_3564,N_3489,N_3382);
nor U3565 (N_3565,N_3354,N_3254);
nand U3566 (N_3566,N_3353,N_3339);
or U3567 (N_3567,N_3430,N_3420);
nand U3568 (N_3568,N_3406,N_3446);
or U3569 (N_3569,N_3345,N_3278);
or U3570 (N_3570,N_3343,N_3388);
nand U3571 (N_3571,N_3327,N_3282);
nand U3572 (N_3572,N_3480,N_3341);
and U3573 (N_3573,N_3409,N_3338);
xnor U3574 (N_3574,N_3250,N_3273);
nand U3575 (N_3575,N_3494,N_3359);
nand U3576 (N_3576,N_3374,N_3467);
or U3577 (N_3577,N_3393,N_3441);
xor U3578 (N_3578,N_3294,N_3264);
or U3579 (N_3579,N_3361,N_3270);
nor U3580 (N_3580,N_3263,N_3484);
nand U3581 (N_3581,N_3277,N_3337);
or U3582 (N_3582,N_3397,N_3253);
xor U3583 (N_3583,N_3308,N_3463);
xnor U3584 (N_3584,N_3306,N_3444);
and U3585 (N_3585,N_3311,N_3462);
and U3586 (N_3586,N_3331,N_3423);
and U3587 (N_3587,N_3283,N_3285);
and U3588 (N_3588,N_3482,N_3476);
nor U3589 (N_3589,N_3448,N_3478);
nand U3590 (N_3590,N_3412,N_3271);
or U3591 (N_3591,N_3477,N_3381);
nand U3592 (N_3592,N_3347,N_3328);
or U3593 (N_3593,N_3366,N_3267);
and U3594 (N_3594,N_3255,N_3459);
xnor U3595 (N_3595,N_3279,N_3355);
nand U3596 (N_3596,N_3425,N_3335);
xnor U3597 (N_3597,N_3268,N_3298);
or U3598 (N_3598,N_3402,N_3497);
nand U3599 (N_3599,N_3455,N_3433);
and U3600 (N_3600,N_3479,N_3305);
and U3601 (N_3601,N_3419,N_3450);
and U3602 (N_3602,N_3380,N_3265);
nor U3603 (N_3603,N_3286,N_3449);
xor U3604 (N_3604,N_3256,N_3258);
or U3605 (N_3605,N_3266,N_3395);
or U3606 (N_3606,N_3438,N_3291);
nor U3607 (N_3607,N_3350,N_3280);
xnor U3608 (N_3608,N_3396,N_3314);
or U3609 (N_3609,N_3307,N_3440);
xnor U3610 (N_3610,N_3274,N_3499);
nor U3611 (N_3611,N_3443,N_3454);
nor U3612 (N_3612,N_3407,N_3408);
nand U3613 (N_3613,N_3398,N_3385);
xnor U3614 (N_3614,N_3251,N_3292);
xnor U3615 (N_3615,N_3334,N_3276);
nand U3616 (N_3616,N_3437,N_3295);
nand U3617 (N_3617,N_3313,N_3474);
or U3618 (N_3618,N_3492,N_3488);
nand U3619 (N_3619,N_3259,N_3411);
nand U3620 (N_3620,N_3322,N_3439);
nand U3621 (N_3621,N_3442,N_3364);
and U3622 (N_3622,N_3496,N_3284);
or U3623 (N_3623,N_3330,N_3417);
xnor U3624 (N_3624,N_3383,N_3453);
and U3625 (N_3625,N_3479,N_3361);
nand U3626 (N_3626,N_3493,N_3378);
or U3627 (N_3627,N_3256,N_3350);
xnor U3628 (N_3628,N_3263,N_3267);
nand U3629 (N_3629,N_3453,N_3405);
xor U3630 (N_3630,N_3416,N_3315);
nand U3631 (N_3631,N_3395,N_3458);
xnor U3632 (N_3632,N_3282,N_3411);
or U3633 (N_3633,N_3489,N_3324);
or U3634 (N_3634,N_3301,N_3338);
xnor U3635 (N_3635,N_3296,N_3253);
nor U3636 (N_3636,N_3436,N_3286);
or U3637 (N_3637,N_3403,N_3419);
nand U3638 (N_3638,N_3488,N_3321);
nand U3639 (N_3639,N_3469,N_3314);
or U3640 (N_3640,N_3385,N_3395);
and U3641 (N_3641,N_3464,N_3367);
nor U3642 (N_3642,N_3323,N_3498);
or U3643 (N_3643,N_3478,N_3348);
nand U3644 (N_3644,N_3442,N_3339);
and U3645 (N_3645,N_3353,N_3432);
and U3646 (N_3646,N_3442,N_3476);
xnor U3647 (N_3647,N_3348,N_3428);
and U3648 (N_3648,N_3308,N_3262);
or U3649 (N_3649,N_3409,N_3419);
and U3650 (N_3650,N_3392,N_3494);
nand U3651 (N_3651,N_3403,N_3325);
xnor U3652 (N_3652,N_3423,N_3381);
or U3653 (N_3653,N_3298,N_3283);
nand U3654 (N_3654,N_3373,N_3490);
or U3655 (N_3655,N_3262,N_3411);
and U3656 (N_3656,N_3355,N_3318);
and U3657 (N_3657,N_3469,N_3315);
nor U3658 (N_3658,N_3451,N_3307);
nor U3659 (N_3659,N_3394,N_3409);
and U3660 (N_3660,N_3301,N_3436);
nor U3661 (N_3661,N_3332,N_3420);
and U3662 (N_3662,N_3463,N_3303);
and U3663 (N_3663,N_3258,N_3487);
nand U3664 (N_3664,N_3480,N_3460);
xnor U3665 (N_3665,N_3301,N_3409);
or U3666 (N_3666,N_3288,N_3356);
or U3667 (N_3667,N_3445,N_3443);
and U3668 (N_3668,N_3395,N_3417);
and U3669 (N_3669,N_3300,N_3344);
xnor U3670 (N_3670,N_3475,N_3458);
xnor U3671 (N_3671,N_3294,N_3257);
nand U3672 (N_3672,N_3283,N_3494);
and U3673 (N_3673,N_3426,N_3480);
and U3674 (N_3674,N_3496,N_3359);
xnor U3675 (N_3675,N_3356,N_3432);
and U3676 (N_3676,N_3326,N_3457);
xor U3677 (N_3677,N_3471,N_3348);
or U3678 (N_3678,N_3256,N_3474);
nor U3679 (N_3679,N_3283,N_3325);
nand U3680 (N_3680,N_3282,N_3294);
nand U3681 (N_3681,N_3332,N_3468);
xor U3682 (N_3682,N_3427,N_3372);
nor U3683 (N_3683,N_3348,N_3291);
or U3684 (N_3684,N_3379,N_3452);
and U3685 (N_3685,N_3354,N_3274);
nor U3686 (N_3686,N_3497,N_3300);
xnor U3687 (N_3687,N_3307,N_3377);
nand U3688 (N_3688,N_3414,N_3442);
nor U3689 (N_3689,N_3436,N_3345);
xor U3690 (N_3690,N_3291,N_3264);
nand U3691 (N_3691,N_3490,N_3480);
or U3692 (N_3692,N_3346,N_3400);
and U3693 (N_3693,N_3273,N_3333);
and U3694 (N_3694,N_3440,N_3383);
or U3695 (N_3695,N_3315,N_3497);
and U3696 (N_3696,N_3335,N_3348);
and U3697 (N_3697,N_3373,N_3482);
nand U3698 (N_3698,N_3446,N_3491);
xnor U3699 (N_3699,N_3362,N_3372);
nor U3700 (N_3700,N_3417,N_3335);
nand U3701 (N_3701,N_3345,N_3384);
and U3702 (N_3702,N_3359,N_3406);
nand U3703 (N_3703,N_3369,N_3334);
nor U3704 (N_3704,N_3310,N_3448);
or U3705 (N_3705,N_3253,N_3332);
nand U3706 (N_3706,N_3295,N_3499);
xor U3707 (N_3707,N_3306,N_3379);
nand U3708 (N_3708,N_3489,N_3368);
nand U3709 (N_3709,N_3441,N_3274);
and U3710 (N_3710,N_3293,N_3480);
or U3711 (N_3711,N_3442,N_3489);
xor U3712 (N_3712,N_3426,N_3434);
xnor U3713 (N_3713,N_3455,N_3427);
and U3714 (N_3714,N_3284,N_3357);
xnor U3715 (N_3715,N_3472,N_3284);
and U3716 (N_3716,N_3400,N_3367);
or U3717 (N_3717,N_3263,N_3346);
xnor U3718 (N_3718,N_3273,N_3434);
and U3719 (N_3719,N_3366,N_3361);
nor U3720 (N_3720,N_3398,N_3372);
or U3721 (N_3721,N_3332,N_3280);
nor U3722 (N_3722,N_3368,N_3358);
nor U3723 (N_3723,N_3458,N_3414);
nor U3724 (N_3724,N_3393,N_3310);
or U3725 (N_3725,N_3457,N_3408);
and U3726 (N_3726,N_3338,N_3488);
xnor U3727 (N_3727,N_3339,N_3366);
nand U3728 (N_3728,N_3392,N_3440);
and U3729 (N_3729,N_3365,N_3423);
nand U3730 (N_3730,N_3436,N_3261);
and U3731 (N_3731,N_3408,N_3496);
xnor U3732 (N_3732,N_3380,N_3259);
or U3733 (N_3733,N_3284,N_3267);
or U3734 (N_3734,N_3375,N_3438);
xnor U3735 (N_3735,N_3438,N_3259);
and U3736 (N_3736,N_3363,N_3456);
xnor U3737 (N_3737,N_3292,N_3324);
xor U3738 (N_3738,N_3470,N_3462);
nand U3739 (N_3739,N_3475,N_3346);
xor U3740 (N_3740,N_3263,N_3402);
xor U3741 (N_3741,N_3260,N_3301);
xnor U3742 (N_3742,N_3269,N_3388);
nand U3743 (N_3743,N_3484,N_3437);
and U3744 (N_3744,N_3296,N_3346);
and U3745 (N_3745,N_3414,N_3305);
nor U3746 (N_3746,N_3326,N_3444);
and U3747 (N_3747,N_3355,N_3493);
nand U3748 (N_3748,N_3421,N_3430);
or U3749 (N_3749,N_3282,N_3447);
xnor U3750 (N_3750,N_3641,N_3705);
nand U3751 (N_3751,N_3548,N_3557);
xor U3752 (N_3752,N_3608,N_3675);
nor U3753 (N_3753,N_3525,N_3592);
and U3754 (N_3754,N_3537,N_3604);
nand U3755 (N_3755,N_3731,N_3720);
or U3756 (N_3756,N_3544,N_3617);
xor U3757 (N_3757,N_3569,N_3615);
nand U3758 (N_3758,N_3578,N_3530);
and U3759 (N_3759,N_3621,N_3695);
nand U3760 (N_3760,N_3724,N_3741);
or U3761 (N_3761,N_3676,N_3550);
and U3762 (N_3762,N_3523,N_3736);
nand U3763 (N_3763,N_3712,N_3650);
nand U3764 (N_3764,N_3703,N_3568);
xor U3765 (N_3765,N_3664,N_3536);
nand U3766 (N_3766,N_3609,N_3593);
nor U3767 (N_3767,N_3691,N_3574);
nor U3768 (N_3768,N_3631,N_3648);
and U3769 (N_3769,N_3502,N_3554);
xor U3770 (N_3770,N_3743,N_3605);
nor U3771 (N_3771,N_3545,N_3505);
and U3772 (N_3772,N_3588,N_3589);
nor U3773 (N_3773,N_3566,N_3531);
and U3774 (N_3774,N_3688,N_3672);
and U3775 (N_3775,N_3749,N_3694);
and U3776 (N_3776,N_3516,N_3561);
or U3777 (N_3777,N_3696,N_3522);
xor U3778 (N_3778,N_3682,N_3614);
nor U3779 (N_3779,N_3628,N_3541);
xnor U3780 (N_3780,N_3529,N_3580);
nand U3781 (N_3781,N_3700,N_3619);
nor U3782 (N_3782,N_3528,N_3713);
xor U3783 (N_3783,N_3680,N_3507);
and U3784 (N_3784,N_3501,N_3655);
or U3785 (N_3785,N_3627,N_3598);
and U3786 (N_3786,N_3629,N_3666);
nand U3787 (N_3787,N_3500,N_3727);
and U3788 (N_3788,N_3660,N_3504);
xor U3789 (N_3789,N_3607,N_3564);
nor U3790 (N_3790,N_3622,N_3624);
nor U3791 (N_3791,N_3526,N_3517);
or U3792 (N_3792,N_3725,N_3678);
nor U3793 (N_3793,N_3715,N_3726);
nor U3794 (N_3794,N_3613,N_3611);
or U3795 (N_3795,N_3563,N_3709);
xnor U3796 (N_3796,N_3527,N_3639);
nor U3797 (N_3797,N_3534,N_3584);
nand U3798 (N_3798,N_3706,N_3535);
nand U3799 (N_3799,N_3538,N_3539);
nor U3800 (N_3800,N_3571,N_3735);
or U3801 (N_3801,N_3555,N_3646);
xnor U3802 (N_3802,N_3596,N_3633);
nor U3803 (N_3803,N_3677,N_3728);
xnor U3804 (N_3804,N_3625,N_3603);
or U3805 (N_3805,N_3684,N_3644);
nor U3806 (N_3806,N_3637,N_3708);
nand U3807 (N_3807,N_3734,N_3690);
xor U3808 (N_3808,N_3693,N_3573);
nor U3809 (N_3809,N_3626,N_3674);
xnor U3810 (N_3810,N_3582,N_3740);
xnor U3811 (N_3811,N_3746,N_3689);
nand U3812 (N_3812,N_3657,N_3547);
or U3813 (N_3813,N_3585,N_3583);
and U3814 (N_3814,N_3510,N_3513);
nor U3815 (N_3815,N_3509,N_3623);
nor U3816 (N_3816,N_3699,N_3685);
xor U3817 (N_3817,N_3612,N_3524);
xor U3818 (N_3818,N_3601,N_3640);
xnor U3819 (N_3819,N_3519,N_3521);
nor U3820 (N_3820,N_3681,N_3662);
or U3821 (N_3821,N_3514,N_3667);
or U3822 (N_3822,N_3653,N_3591);
or U3823 (N_3823,N_3745,N_3506);
nand U3824 (N_3824,N_3618,N_3656);
nand U3825 (N_3825,N_3575,N_3630);
and U3826 (N_3826,N_3565,N_3542);
nor U3827 (N_3827,N_3707,N_3553);
or U3828 (N_3828,N_3632,N_3665);
nor U3829 (N_3829,N_3503,N_3616);
or U3830 (N_3830,N_3711,N_3649);
and U3831 (N_3831,N_3645,N_3562);
or U3832 (N_3832,N_3532,N_3661);
nand U3833 (N_3833,N_3737,N_3581);
nand U3834 (N_3834,N_3635,N_3739);
nor U3835 (N_3835,N_3552,N_3597);
nand U3836 (N_3836,N_3654,N_3520);
and U3837 (N_3837,N_3549,N_3747);
nand U3838 (N_3838,N_3668,N_3663);
nand U3839 (N_3839,N_3511,N_3733);
xnor U3840 (N_3840,N_3669,N_3560);
and U3841 (N_3841,N_3698,N_3687);
xnor U3842 (N_3842,N_3742,N_3556);
nand U3843 (N_3843,N_3732,N_3738);
nor U3844 (N_3844,N_3697,N_3679);
and U3845 (N_3845,N_3659,N_3647);
nor U3846 (N_3846,N_3610,N_3518);
xnor U3847 (N_3847,N_3594,N_3587);
xor U3848 (N_3848,N_3652,N_3658);
nor U3849 (N_3849,N_3686,N_3606);
and U3850 (N_3850,N_3638,N_3692);
xnor U3851 (N_3851,N_3671,N_3718);
nand U3852 (N_3852,N_3651,N_3577);
nand U3853 (N_3853,N_3634,N_3620);
nand U3854 (N_3854,N_3717,N_3602);
nor U3855 (N_3855,N_3559,N_3636);
xor U3856 (N_3856,N_3533,N_3512);
and U3857 (N_3857,N_3558,N_3714);
xor U3858 (N_3858,N_3719,N_3543);
and U3859 (N_3859,N_3730,N_3670);
or U3860 (N_3860,N_3551,N_3683);
nor U3861 (N_3861,N_3723,N_3590);
and U3862 (N_3862,N_3673,N_3744);
nor U3863 (N_3863,N_3595,N_3546);
nand U3864 (N_3864,N_3722,N_3579);
nor U3865 (N_3865,N_3567,N_3572);
nor U3866 (N_3866,N_3586,N_3515);
nand U3867 (N_3867,N_3508,N_3716);
nand U3868 (N_3868,N_3570,N_3540);
nand U3869 (N_3869,N_3710,N_3701);
xnor U3870 (N_3870,N_3576,N_3721);
or U3871 (N_3871,N_3600,N_3704);
xnor U3872 (N_3872,N_3729,N_3642);
xnor U3873 (N_3873,N_3643,N_3748);
nor U3874 (N_3874,N_3599,N_3702);
nor U3875 (N_3875,N_3651,N_3609);
nand U3876 (N_3876,N_3542,N_3592);
xor U3877 (N_3877,N_3603,N_3589);
or U3878 (N_3878,N_3584,N_3607);
and U3879 (N_3879,N_3660,N_3619);
nand U3880 (N_3880,N_3633,N_3748);
xor U3881 (N_3881,N_3658,N_3592);
nor U3882 (N_3882,N_3678,N_3611);
xnor U3883 (N_3883,N_3602,N_3707);
or U3884 (N_3884,N_3746,N_3541);
nor U3885 (N_3885,N_3749,N_3741);
nand U3886 (N_3886,N_3508,N_3736);
nor U3887 (N_3887,N_3586,N_3548);
nor U3888 (N_3888,N_3724,N_3728);
nor U3889 (N_3889,N_3657,N_3512);
and U3890 (N_3890,N_3703,N_3635);
nand U3891 (N_3891,N_3603,N_3504);
or U3892 (N_3892,N_3548,N_3606);
and U3893 (N_3893,N_3525,N_3506);
or U3894 (N_3894,N_3671,N_3532);
nand U3895 (N_3895,N_3620,N_3740);
and U3896 (N_3896,N_3573,N_3699);
and U3897 (N_3897,N_3683,N_3619);
nor U3898 (N_3898,N_3671,N_3716);
nand U3899 (N_3899,N_3609,N_3662);
nor U3900 (N_3900,N_3584,N_3679);
nand U3901 (N_3901,N_3628,N_3516);
xnor U3902 (N_3902,N_3620,N_3643);
and U3903 (N_3903,N_3626,N_3654);
nand U3904 (N_3904,N_3674,N_3525);
nand U3905 (N_3905,N_3547,N_3676);
nor U3906 (N_3906,N_3718,N_3689);
nor U3907 (N_3907,N_3512,N_3683);
and U3908 (N_3908,N_3733,N_3683);
nand U3909 (N_3909,N_3627,N_3729);
xor U3910 (N_3910,N_3638,N_3666);
or U3911 (N_3911,N_3559,N_3689);
nand U3912 (N_3912,N_3749,N_3701);
nor U3913 (N_3913,N_3588,N_3551);
xor U3914 (N_3914,N_3641,N_3582);
xor U3915 (N_3915,N_3737,N_3552);
and U3916 (N_3916,N_3546,N_3543);
or U3917 (N_3917,N_3749,N_3613);
xnor U3918 (N_3918,N_3647,N_3652);
or U3919 (N_3919,N_3671,N_3502);
and U3920 (N_3920,N_3533,N_3579);
nand U3921 (N_3921,N_3725,N_3552);
nand U3922 (N_3922,N_3671,N_3747);
xnor U3923 (N_3923,N_3615,N_3735);
nand U3924 (N_3924,N_3738,N_3681);
xnor U3925 (N_3925,N_3638,N_3644);
and U3926 (N_3926,N_3524,N_3575);
xor U3927 (N_3927,N_3517,N_3694);
nor U3928 (N_3928,N_3749,N_3508);
nor U3929 (N_3929,N_3572,N_3651);
and U3930 (N_3930,N_3557,N_3678);
or U3931 (N_3931,N_3676,N_3576);
xor U3932 (N_3932,N_3683,N_3686);
nor U3933 (N_3933,N_3612,N_3631);
nand U3934 (N_3934,N_3700,N_3685);
nand U3935 (N_3935,N_3533,N_3703);
nand U3936 (N_3936,N_3512,N_3612);
and U3937 (N_3937,N_3716,N_3653);
and U3938 (N_3938,N_3538,N_3748);
nand U3939 (N_3939,N_3704,N_3691);
and U3940 (N_3940,N_3520,N_3661);
nand U3941 (N_3941,N_3732,N_3688);
xor U3942 (N_3942,N_3507,N_3584);
and U3943 (N_3943,N_3740,N_3722);
xor U3944 (N_3944,N_3728,N_3699);
or U3945 (N_3945,N_3726,N_3519);
nor U3946 (N_3946,N_3748,N_3608);
or U3947 (N_3947,N_3653,N_3703);
nand U3948 (N_3948,N_3659,N_3542);
xnor U3949 (N_3949,N_3652,N_3523);
nand U3950 (N_3950,N_3651,N_3509);
xor U3951 (N_3951,N_3516,N_3684);
and U3952 (N_3952,N_3747,N_3617);
nand U3953 (N_3953,N_3533,N_3585);
nand U3954 (N_3954,N_3680,N_3555);
nand U3955 (N_3955,N_3526,N_3505);
and U3956 (N_3956,N_3702,N_3650);
nand U3957 (N_3957,N_3693,N_3506);
nor U3958 (N_3958,N_3577,N_3593);
or U3959 (N_3959,N_3638,N_3654);
or U3960 (N_3960,N_3711,N_3674);
nand U3961 (N_3961,N_3693,N_3646);
nor U3962 (N_3962,N_3605,N_3614);
or U3963 (N_3963,N_3605,N_3666);
nand U3964 (N_3964,N_3587,N_3713);
and U3965 (N_3965,N_3607,N_3582);
or U3966 (N_3966,N_3568,N_3745);
or U3967 (N_3967,N_3516,N_3545);
and U3968 (N_3968,N_3552,N_3702);
nand U3969 (N_3969,N_3657,N_3694);
nand U3970 (N_3970,N_3683,N_3742);
or U3971 (N_3971,N_3646,N_3543);
and U3972 (N_3972,N_3575,N_3642);
nor U3973 (N_3973,N_3680,N_3570);
nor U3974 (N_3974,N_3704,N_3638);
or U3975 (N_3975,N_3613,N_3616);
nor U3976 (N_3976,N_3525,N_3737);
nand U3977 (N_3977,N_3661,N_3549);
and U3978 (N_3978,N_3666,N_3606);
nand U3979 (N_3979,N_3722,N_3605);
xnor U3980 (N_3980,N_3646,N_3583);
xor U3981 (N_3981,N_3569,N_3583);
xnor U3982 (N_3982,N_3552,N_3731);
xnor U3983 (N_3983,N_3512,N_3510);
xor U3984 (N_3984,N_3720,N_3540);
or U3985 (N_3985,N_3658,N_3630);
or U3986 (N_3986,N_3603,N_3544);
nor U3987 (N_3987,N_3641,N_3749);
xor U3988 (N_3988,N_3546,N_3530);
and U3989 (N_3989,N_3597,N_3680);
or U3990 (N_3990,N_3503,N_3594);
or U3991 (N_3991,N_3731,N_3687);
or U3992 (N_3992,N_3533,N_3641);
nand U3993 (N_3993,N_3678,N_3656);
nor U3994 (N_3994,N_3652,N_3507);
nand U3995 (N_3995,N_3623,N_3748);
xor U3996 (N_3996,N_3605,N_3664);
nor U3997 (N_3997,N_3629,N_3602);
xnor U3998 (N_3998,N_3603,N_3506);
and U3999 (N_3999,N_3600,N_3534);
nand U4000 (N_4000,N_3811,N_3923);
xor U4001 (N_4001,N_3793,N_3761);
nor U4002 (N_4002,N_3905,N_3920);
xnor U4003 (N_4003,N_3967,N_3791);
and U4004 (N_4004,N_3868,N_3778);
nor U4005 (N_4005,N_3823,N_3827);
nand U4006 (N_4006,N_3938,N_3973);
and U4007 (N_4007,N_3825,N_3805);
xnor U4008 (N_4008,N_3919,N_3990);
xor U4009 (N_4009,N_3871,N_3776);
xor U4010 (N_4010,N_3894,N_3829);
xnor U4011 (N_4011,N_3928,N_3876);
nor U4012 (N_4012,N_3820,N_3880);
nor U4013 (N_4013,N_3888,N_3951);
xor U4014 (N_4014,N_3981,N_3937);
and U4015 (N_4015,N_3863,N_3770);
nand U4016 (N_4016,N_3949,N_3918);
and U4017 (N_4017,N_3874,N_3872);
or U4018 (N_4018,N_3842,N_3786);
and U4019 (N_4019,N_3802,N_3760);
and U4020 (N_4020,N_3980,N_3921);
and U4021 (N_4021,N_3839,N_3883);
nor U4022 (N_4022,N_3979,N_3816);
and U4023 (N_4023,N_3843,N_3881);
nand U4024 (N_4024,N_3867,N_3817);
or U4025 (N_4025,N_3806,N_3754);
xor U4026 (N_4026,N_3808,N_3859);
xor U4027 (N_4027,N_3952,N_3984);
or U4028 (N_4028,N_3790,N_3769);
or U4029 (N_4029,N_3813,N_3877);
xnor U4030 (N_4030,N_3955,N_3753);
or U4031 (N_4031,N_3957,N_3785);
nand U4032 (N_4032,N_3902,N_3857);
xor U4033 (N_4033,N_3762,N_3815);
or U4034 (N_4034,N_3986,N_3914);
and U4035 (N_4035,N_3798,N_3830);
nand U4036 (N_4036,N_3828,N_3862);
xor U4037 (N_4037,N_3916,N_3978);
xnor U4038 (N_4038,N_3934,N_3757);
xor U4039 (N_4039,N_3908,N_3925);
xor U4040 (N_4040,N_3822,N_3800);
and U4041 (N_4041,N_3909,N_3755);
xor U4042 (N_4042,N_3807,N_3895);
xor U4043 (N_4043,N_3959,N_3852);
and U4044 (N_4044,N_3963,N_3898);
nor U4045 (N_4045,N_3782,N_3960);
nand U4046 (N_4046,N_3885,N_3958);
nor U4047 (N_4047,N_3787,N_3801);
xor U4048 (N_4048,N_3858,N_3904);
nor U4049 (N_4049,N_3795,N_3911);
and U4050 (N_4050,N_3932,N_3993);
nand U4051 (N_4051,N_3953,N_3861);
nand U4052 (N_4052,N_3936,N_3974);
nand U4053 (N_4053,N_3943,N_3985);
and U4054 (N_4054,N_3869,N_3882);
or U4055 (N_4055,N_3939,N_3834);
xor U4056 (N_4056,N_3948,N_3915);
or U4057 (N_4057,N_3995,N_3835);
nor U4058 (N_4058,N_3794,N_3996);
or U4059 (N_4059,N_3906,N_3983);
or U4060 (N_4060,N_3899,N_3781);
xnor U4061 (N_4061,N_3853,N_3796);
nor U4062 (N_4062,N_3977,N_3931);
nor U4063 (N_4063,N_3961,N_3879);
nand U4064 (N_4064,N_3950,N_3933);
and U4065 (N_4065,N_3774,N_3803);
and U4066 (N_4066,N_3972,N_3942);
and U4067 (N_4067,N_3768,N_3849);
nand U4068 (N_4068,N_3964,N_3892);
nand U4069 (N_4069,N_3897,N_3884);
nand U4070 (N_4070,N_3836,N_3821);
xor U4071 (N_4071,N_3900,N_3818);
or U4072 (N_4072,N_3850,N_3889);
xor U4073 (N_4073,N_3941,N_3992);
nand U4074 (N_4074,N_3779,N_3875);
xnor U4075 (N_4075,N_3763,N_3926);
xnor U4076 (N_4076,N_3772,N_3930);
or U4077 (N_4077,N_3789,N_3890);
or U4078 (N_4078,N_3841,N_3994);
nand U4079 (N_4079,N_3771,N_3809);
nor U4080 (N_4080,N_3860,N_3944);
xnor U4081 (N_4081,N_3780,N_3854);
xnor U4082 (N_4082,N_3976,N_3764);
xnor U4083 (N_4083,N_3924,N_3962);
and U4084 (N_4084,N_3812,N_3997);
xnor U4085 (N_4085,N_3856,N_3917);
nand U4086 (N_4086,N_3999,N_3956);
and U4087 (N_4087,N_3756,N_3975);
nor U4088 (N_4088,N_3965,N_3947);
nand U4089 (N_4089,N_3846,N_3766);
nor U4090 (N_4090,N_3844,N_3824);
xor U4091 (N_4091,N_3946,N_3750);
nand U4092 (N_4092,N_3797,N_3873);
and U4093 (N_4093,N_3752,N_3893);
nand U4094 (N_4094,N_3913,N_3840);
and U4095 (N_4095,N_3988,N_3991);
xor U4096 (N_4096,N_3777,N_3826);
or U4097 (N_4097,N_3788,N_3773);
or U4098 (N_4098,N_3751,N_3784);
nor U4099 (N_4099,N_3982,N_3969);
xor U4100 (N_4100,N_3833,N_3940);
nand U4101 (N_4101,N_3935,N_3971);
nand U4102 (N_4102,N_3765,N_3847);
or U4103 (N_4103,N_3855,N_3891);
nand U4104 (N_4104,N_3954,N_3896);
xnor U4105 (N_4105,N_3831,N_3927);
xor U4106 (N_4106,N_3945,N_3912);
or U4107 (N_4107,N_3783,N_3845);
and U4108 (N_4108,N_3758,N_3887);
or U4109 (N_4109,N_3966,N_3998);
nor U4110 (N_4110,N_3819,N_3837);
nand U4111 (N_4111,N_3804,N_3864);
or U4112 (N_4112,N_3989,N_3759);
or U4113 (N_4113,N_3968,N_3799);
nand U4114 (N_4114,N_3987,N_3848);
or U4115 (N_4115,N_3775,N_3922);
or U4116 (N_4116,N_3886,N_3870);
xor U4117 (N_4117,N_3903,N_3838);
and U4118 (N_4118,N_3865,N_3901);
xor U4119 (N_4119,N_3810,N_3851);
nor U4120 (N_4120,N_3970,N_3832);
or U4121 (N_4121,N_3792,N_3907);
nor U4122 (N_4122,N_3767,N_3910);
and U4123 (N_4123,N_3929,N_3878);
or U4124 (N_4124,N_3866,N_3814);
nor U4125 (N_4125,N_3973,N_3760);
xor U4126 (N_4126,N_3945,N_3957);
or U4127 (N_4127,N_3955,N_3822);
nor U4128 (N_4128,N_3849,N_3769);
nor U4129 (N_4129,N_3778,N_3912);
or U4130 (N_4130,N_3767,N_3978);
nor U4131 (N_4131,N_3870,N_3759);
nand U4132 (N_4132,N_3813,N_3872);
nor U4133 (N_4133,N_3779,N_3898);
nand U4134 (N_4134,N_3964,N_3893);
nand U4135 (N_4135,N_3824,N_3945);
xor U4136 (N_4136,N_3924,N_3810);
and U4137 (N_4137,N_3882,N_3892);
xor U4138 (N_4138,N_3930,N_3890);
nand U4139 (N_4139,N_3969,N_3953);
and U4140 (N_4140,N_3998,N_3901);
nor U4141 (N_4141,N_3762,N_3811);
and U4142 (N_4142,N_3772,N_3868);
xor U4143 (N_4143,N_3982,N_3971);
nand U4144 (N_4144,N_3885,N_3812);
xnor U4145 (N_4145,N_3873,N_3778);
nand U4146 (N_4146,N_3814,N_3968);
nand U4147 (N_4147,N_3788,N_3986);
and U4148 (N_4148,N_3816,N_3982);
nand U4149 (N_4149,N_3915,N_3938);
or U4150 (N_4150,N_3859,N_3809);
and U4151 (N_4151,N_3846,N_3839);
xor U4152 (N_4152,N_3986,N_3770);
nand U4153 (N_4153,N_3935,N_3947);
or U4154 (N_4154,N_3921,N_3899);
and U4155 (N_4155,N_3866,N_3751);
xnor U4156 (N_4156,N_3780,N_3943);
xnor U4157 (N_4157,N_3846,N_3840);
nand U4158 (N_4158,N_3784,N_3987);
xnor U4159 (N_4159,N_3938,N_3806);
and U4160 (N_4160,N_3817,N_3945);
and U4161 (N_4161,N_3783,N_3997);
xnor U4162 (N_4162,N_3758,N_3978);
xor U4163 (N_4163,N_3811,N_3847);
or U4164 (N_4164,N_3818,N_3980);
and U4165 (N_4165,N_3811,N_3851);
xnor U4166 (N_4166,N_3959,N_3866);
and U4167 (N_4167,N_3961,N_3928);
and U4168 (N_4168,N_3782,N_3834);
and U4169 (N_4169,N_3788,N_3906);
xor U4170 (N_4170,N_3790,N_3988);
and U4171 (N_4171,N_3783,N_3795);
nor U4172 (N_4172,N_3993,N_3959);
or U4173 (N_4173,N_3803,N_3979);
nand U4174 (N_4174,N_3963,N_3974);
nand U4175 (N_4175,N_3965,N_3928);
or U4176 (N_4176,N_3820,N_3879);
nand U4177 (N_4177,N_3793,N_3992);
and U4178 (N_4178,N_3989,N_3937);
or U4179 (N_4179,N_3860,N_3779);
or U4180 (N_4180,N_3789,N_3823);
nand U4181 (N_4181,N_3951,N_3935);
nor U4182 (N_4182,N_3842,N_3810);
or U4183 (N_4183,N_3968,N_3912);
nand U4184 (N_4184,N_3907,N_3834);
xor U4185 (N_4185,N_3848,N_3855);
or U4186 (N_4186,N_3891,N_3991);
or U4187 (N_4187,N_3997,N_3770);
nor U4188 (N_4188,N_3912,N_3884);
nand U4189 (N_4189,N_3779,N_3809);
or U4190 (N_4190,N_3957,N_3860);
and U4191 (N_4191,N_3931,N_3988);
xnor U4192 (N_4192,N_3820,N_3806);
nand U4193 (N_4193,N_3914,N_3766);
and U4194 (N_4194,N_3752,N_3830);
or U4195 (N_4195,N_3978,N_3814);
nor U4196 (N_4196,N_3781,N_3991);
xor U4197 (N_4197,N_3817,N_3953);
or U4198 (N_4198,N_3928,N_3758);
nand U4199 (N_4199,N_3991,N_3966);
and U4200 (N_4200,N_3768,N_3921);
nand U4201 (N_4201,N_3973,N_3922);
and U4202 (N_4202,N_3846,N_3848);
or U4203 (N_4203,N_3802,N_3916);
xnor U4204 (N_4204,N_3830,N_3928);
nand U4205 (N_4205,N_3827,N_3783);
or U4206 (N_4206,N_3832,N_3883);
and U4207 (N_4207,N_3835,N_3866);
nor U4208 (N_4208,N_3784,N_3985);
or U4209 (N_4209,N_3752,N_3855);
xor U4210 (N_4210,N_3905,N_3815);
and U4211 (N_4211,N_3811,N_3934);
or U4212 (N_4212,N_3908,N_3778);
nor U4213 (N_4213,N_3893,N_3792);
nor U4214 (N_4214,N_3900,N_3752);
or U4215 (N_4215,N_3785,N_3895);
or U4216 (N_4216,N_3930,N_3806);
or U4217 (N_4217,N_3800,N_3912);
and U4218 (N_4218,N_3950,N_3806);
nand U4219 (N_4219,N_3886,N_3854);
nand U4220 (N_4220,N_3940,N_3821);
xor U4221 (N_4221,N_3890,N_3856);
nand U4222 (N_4222,N_3784,N_3925);
xnor U4223 (N_4223,N_3993,N_3826);
xnor U4224 (N_4224,N_3966,N_3944);
nand U4225 (N_4225,N_3921,N_3853);
xnor U4226 (N_4226,N_3905,N_3913);
or U4227 (N_4227,N_3759,N_3792);
and U4228 (N_4228,N_3889,N_3899);
nand U4229 (N_4229,N_3779,N_3768);
xor U4230 (N_4230,N_3764,N_3967);
or U4231 (N_4231,N_3980,N_3967);
and U4232 (N_4232,N_3966,N_3759);
or U4233 (N_4233,N_3947,N_3759);
or U4234 (N_4234,N_3986,N_3882);
nor U4235 (N_4235,N_3967,N_3867);
nand U4236 (N_4236,N_3802,N_3766);
xor U4237 (N_4237,N_3965,N_3938);
nand U4238 (N_4238,N_3934,N_3971);
nor U4239 (N_4239,N_3906,N_3839);
or U4240 (N_4240,N_3780,N_3843);
nand U4241 (N_4241,N_3976,N_3884);
nand U4242 (N_4242,N_3851,N_3899);
nand U4243 (N_4243,N_3818,N_3889);
or U4244 (N_4244,N_3929,N_3910);
xnor U4245 (N_4245,N_3947,N_3757);
or U4246 (N_4246,N_3856,N_3777);
nor U4247 (N_4247,N_3998,N_3782);
xor U4248 (N_4248,N_3986,N_3841);
nand U4249 (N_4249,N_3922,N_3863);
nand U4250 (N_4250,N_4074,N_4011);
and U4251 (N_4251,N_4036,N_4043);
nor U4252 (N_4252,N_4207,N_4001);
and U4253 (N_4253,N_4159,N_4116);
or U4254 (N_4254,N_4086,N_4137);
xor U4255 (N_4255,N_4205,N_4242);
xor U4256 (N_4256,N_4190,N_4044);
or U4257 (N_4257,N_4025,N_4161);
and U4258 (N_4258,N_4021,N_4217);
and U4259 (N_4259,N_4175,N_4248);
or U4260 (N_4260,N_4123,N_4164);
and U4261 (N_4261,N_4249,N_4100);
nand U4262 (N_4262,N_4122,N_4096);
nand U4263 (N_4263,N_4085,N_4053);
or U4264 (N_4264,N_4196,N_4223);
or U4265 (N_4265,N_4117,N_4002);
nand U4266 (N_4266,N_4212,N_4041);
xnor U4267 (N_4267,N_4170,N_4058);
nor U4268 (N_4268,N_4181,N_4174);
nand U4269 (N_4269,N_4227,N_4082);
nand U4270 (N_4270,N_4120,N_4062);
nand U4271 (N_4271,N_4066,N_4047);
and U4272 (N_4272,N_4108,N_4158);
nor U4273 (N_4273,N_4237,N_4125);
or U4274 (N_4274,N_4195,N_4073);
nor U4275 (N_4275,N_4072,N_4202);
xnor U4276 (N_4276,N_4075,N_4176);
or U4277 (N_4277,N_4135,N_4013);
nand U4278 (N_4278,N_4228,N_4214);
xor U4279 (N_4279,N_4152,N_4008);
nand U4280 (N_4280,N_4051,N_4199);
nor U4281 (N_4281,N_4055,N_4247);
or U4282 (N_4282,N_4084,N_4203);
or U4283 (N_4283,N_4092,N_4143);
nor U4284 (N_4284,N_4064,N_4213);
nor U4285 (N_4285,N_4099,N_4048);
nand U4286 (N_4286,N_4229,N_4091);
and U4287 (N_4287,N_4139,N_4179);
and U4288 (N_4288,N_4140,N_4095);
nand U4289 (N_4289,N_4057,N_4198);
or U4290 (N_4290,N_4016,N_4192);
nor U4291 (N_4291,N_4010,N_4151);
xnor U4292 (N_4292,N_4018,N_4093);
or U4293 (N_4293,N_4065,N_4194);
nor U4294 (N_4294,N_4206,N_4184);
or U4295 (N_4295,N_4241,N_4101);
nand U4296 (N_4296,N_4070,N_4201);
and U4297 (N_4297,N_4127,N_4218);
or U4298 (N_4298,N_4208,N_4146);
xor U4299 (N_4299,N_4149,N_4054);
nor U4300 (N_4300,N_4006,N_4186);
xor U4301 (N_4301,N_4165,N_4019);
nor U4302 (N_4302,N_4180,N_4023);
xor U4303 (N_4303,N_4193,N_4235);
or U4304 (N_4304,N_4160,N_4130);
or U4305 (N_4305,N_4003,N_4124);
nor U4306 (N_4306,N_4168,N_4222);
xor U4307 (N_4307,N_4244,N_4067);
or U4308 (N_4308,N_4077,N_4121);
nand U4309 (N_4309,N_4210,N_4114);
or U4310 (N_4310,N_4076,N_4009);
xor U4311 (N_4311,N_4209,N_4060);
and U4312 (N_4312,N_4182,N_4046);
and U4313 (N_4313,N_4224,N_4232);
xor U4314 (N_4314,N_4071,N_4132);
or U4315 (N_4315,N_4061,N_4173);
xor U4316 (N_4316,N_4191,N_4220);
or U4317 (N_4317,N_4200,N_4156);
nor U4318 (N_4318,N_4236,N_4131);
or U4319 (N_4319,N_4040,N_4211);
nand U4320 (N_4320,N_4017,N_4088);
nor U4321 (N_4321,N_4221,N_4035);
and U4322 (N_4322,N_4144,N_4078);
nand U4323 (N_4323,N_4015,N_4104);
and U4324 (N_4324,N_4038,N_4090);
nor U4325 (N_4325,N_4039,N_4056);
and U4326 (N_4326,N_4037,N_4109);
nand U4327 (N_4327,N_4225,N_4240);
and U4328 (N_4328,N_4231,N_4094);
nand U4329 (N_4329,N_4153,N_4079);
and U4330 (N_4330,N_4172,N_4069);
or U4331 (N_4331,N_4107,N_4042);
xor U4332 (N_4332,N_4183,N_4028);
xor U4333 (N_4333,N_4106,N_4097);
and U4334 (N_4334,N_4012,N_4029);
or U4335 (N_4335,N_4119,N_4063);
or U4336 (N_4336,N_4189,N_4163);
xor U4337 (N_4337,N_4052,N_4014);
or U4338 (N_4338,N_4032,N_4103);
or U4339 (N_4339,N_4031,N_4007);
and U4340 (N_4340,N_4216,N_4081);
and U4341 (N_4341,N_4111,N_4000);
or U4342 (N_4342,N_4020,N_4136);
and U4343 (N_4343,N_4154,N_4234);
and U4344 (N_4344,N_4215,N_4245);
and U4345 (N_4345,N_4049,N_4141);
nor U4346 (N_4346,N_4155,N_4118);
nand U4347 (N_4347,N_4185,N_4134);
xor U4348 (N_4348,N_4239,N_4050);
and U4349 (N_4349,N_4148,N_4150);
nor U4350 (N_4350,N_4033,N_4187);
nand U4351 (N_4351,N_4230,N_4089);
nand U4352 (N_4352,N_4027,N_4059);
nor U4353 (N_4353,N_4098,N_4129);
or U4354 (N_4354,N_4126,N_4045);
or U4355 (N_4355,N_4219,N_4238);
nand U4356 (N_4356,N_4110,N_4022);
xnor U4357 (N_4357,N_4246,N_4171);
nor U4358 (N_4358,N_4026,N_4004);
xor U4359 (N_4359,N_4226,N_4243);
and U4360 (N_4360,N_4087,N_4005);
or U4361 (N_4361,N_4128,N_4147);
nand U4362 (N_4362,N_4167,N_4142);
nand U4363 (N_4363,N_4083,N_4115);
nor U4364 (N_4364,N_4145,N_4105);
nand U4365 (N_4365,N_4169,N_4162);
or U4366 (N_4366,N_4178,N_4157);
xnor U4367 (N_4367,N_4102,N_4197);
nor U4368 (N_4368,N_4204,N_4030);
nor U4369 (N_4369,N_4113,N_4188);
nand U4370 (N_4370,N_4177,N_4166);
nand U4371 (N_4371,N_4034,N_4080);
and U4372 (N_4372,N_4138,N_4233);
or U4373 (N_4373,N_4024,N_4112);
or U4374 (N_4374,N_4133,N_4068);
and U4375 (N_4375,N_4096,N_4146);
nor U4376 (N_4376,N_4005,N_4119);
or U4377 (N_4377,N_4061,N_4068);
nor U4378 (N_4378,N_4244,N_4203);
nand U4379 (N_4379,N_4131,N_4108);
xor U4380 (N_4380,N_4140,N_4078);
or U4381 (N_4381,N_4001,N_4086);
and U4382 (N_4382,N_4026,N_4179);
xnor U4383 (N_4383,N_4229,N_4092);
nand U4384 (N_4384,N_4141,N_4231);
and U4385 (N_4385,N_4011,N_4091);
nor U4386 (N_4386,N_4069,N_4175);
and U4387 (N_4387,N_4093,N_4050);
nand U4388 (N_4388,N_4002,N_4209);
or U4389 (N_4389,N_4067,N_4128);
nand U4390 (N_4390,N_4187,N_4035);
nor U4391 (N_4391,N_4177,N_4016);
nor U4392 (N_4392,N_4085,N_4113);
xnor U4393 (N_4393,N_4233,N_4189);
xnor U4394 (N_4394,N_4172,N_4039);
and U4395 (N_4395,N_4053,N_4178);
nor U4396 (N_4396,N_4221,N_4127);
xnor U4397 (N_4397,N_4126,N_4012);
or U4398 (N_4398,N_4116,N_4088);
xnor U4399 (N_4399,N_4065,N_4057);
nor U4400 (N_4400,N_4032,N_4118);
and U4401 (N_4401,N_4015,N_4223);
nor U4402 (N_4402,N_4182,N_4105);
nand U4403 (N_4403,N_4180,N_4237);
nor U4404 (N_4404,N_4130,N_4194);
or U4405 (N_4405,N_4098,N_4202);
nor U4406 (N_4406,N_4214,N_4217);
xnor U4407 (N_4407,N_4132,N_4243);
or U4408 (N_4408,N_4170,N_4171);
nor U4409 (N_4409,N_4049,N_4183);
or U4410 (N_4410,N_4066,N_4180);
and U4411 (N_4411,N_4201,N_4182);
and U4412 (N_4412,N_4005,N_4011);
nand U4413 (N_4413,N_4014,N_4018);
or U4414 (N_4414,N_4073,N_4081);
and U4415 (N_4415,N_4232,N_4177);
xor U4416 (N_4416,N_4208,N_4230);
and U4417 (N_4417,N_4245,N_4055);
nor U4418 (N_4418,N_4098,N_4154);
nor U4419 (N_4419,N_4154,N_4001);
nor U4420 (N_4420,N_4218,N_4199);
nor U4421 (N_4421,N_4083,N_4236);
nor U4422 (N_4422,N_4013,N_4231);
and U4423 (N_4423,N_4236,N_4144);
nor U4424 (N_4424,N_4216,N_4134);
nand U4425 (N_4425,N_4199,N_4059);
or U4426 (N_4426,N_4243,N_4124);
or U4427 (N_4427,N_4010,N_4097);
nand U4428 (N_4428,N_4073,N_4141);
nor U4429 (N_4429,N_4217,N_4052);
nand U4430 (N_4430,N_4170,N_4221);
nand U4431 (N_4431,N_4010,N_4000);
or U4432 (N_4432,N_4110,N_4078);
nor U4433 (N_4433,N_4143,N_4222);
or U4434 (N_4434,N_4056,N_4150);
nor U4435 (N_4435,N_4140,N_4168);
xnor U4436 (N_4436,N_4169,N_4001);
nand U4437 (N_4437,N_4024,N_4139);
or U4438 (N_4438,N_4055,N_4058);
or U4439 (N_4439,N_4083,N_4239);
xnor U4440 (N_4440,N_4163,N_4055);
or U4441 (N_4441,N_4132,N_4162);
or U4442 (N_4442,N_4204,N_4156);
or U4443 (N_4443,N_4236,N_4170);
nor U4444 (N_4444,N_4105,N_4042);
or U4445 (N_4445,N_4203,N_4110);
and U4446 (N_4446,N_4062,N_4121);
nor U4447 (N_4447,N_4120,N_4097);
xnor U4448 (N_4448,N_4043,N_4146);
nor U4449 (N_4449,N_4195,N_4245);
xor U4450 (N_4450,N_4033,N_4199);
nor U4451 (N_4451,N_4181,N_4141);
or U4452 (N_4452,N_4183,N_4156);
nor U4453 (N_4453,N_4219,N_4073);
nand U4454 (N_4454,N_4074,N_4235);
xor U4455 (N_4455,N_4000,N_4147);
or U4456 (N_4456,N_4198,N_4133);
xnor U4457 (N_4457,N_4209,N_4142);
or U4458 (N_4458,N_4044,N_4079);
xnor U4459 (N_4459,N_4085,N_4032);
or U4460 (N_4460,N_4144,N_4142);
or U4461 (N_4461,N_4014,N_4207);
and U4462 (N_4462,N_4097,N_4028);
xor U4463 (N_4463,N_4102,N_4108);
nor U4464 (N_4464,N_4191,N_4003);
and U4465 (N_4465,N_4208,N_4104);
nand U4466 (N_4466,N_4242,N_4211);
and U4467 (N_4467,N_4034,N_4130);
xnor U4468 (N_4468,N_4041,N_4117);
nand U4469 (N_4469,N_4004,N_4007);
and U4470 (N_4470,N_4126,N_4087);
nor U4471 (N_4471,N_4242,N_4193);
nor U4472 (N_4472,N_4136,N_4220);
nor U4473 (N_4473,N_4066,N_4120);
xor U4474 (N_4474,N_4090,N_4078);
or U4475 (N_4475,N_4176,N_4136);
xor U4476 (N_4476,N_4185,N_4066);
and U4477 (N_4477,N_4026,N_4029);
and U4478 (N_4478,N_4177,N_4098);
xor U4479 (N_4479,N_4203,N_4181);
or U4480 (N_4480,N_4073,N_4049);
nor U4481 (N_4481,N_4202,N_4119);
nand U4482 (N_4482,N_4075,N_4126);
nand U4483 (N_4483,N_4022,N_4241);
nor U4484 (N_4484,N_4011,N_4201);
nand U4485 (N_4485,N_4094,N_4222);
nand U4486 (N_4486,N_4135,N_4081);
nand U4487 (N_4487,N_4063,N_4055);
xor U4488 (N_4488,N_4120,N_4169);
nand U4489 (N_4489,N_4069,N_4084);
and U4490 (N_4490,N_4214,N_4180);
or U4491 (N_4491,N_4211,N_4202);
xor U4492 (N_4492,N_4057,N_4085);
nor U4493 (N_4493,N_4120,N_4214);
xnor U4494 (N_4494,N_4233,N_4083);
xnor U4495 (N_4495,N_4152,N_4144);
nor U4496 (N_4496,N_4201,N_4185);
or U4497 (N_4497,N_4136,N_4096);
nor U4498 (N_4498,N_4073,N_4020);
or U4499 (N_4499,N_4037,N_4098);
or U4500 (N_4500,N_4462,N_4259);
nand U4501 (N_4501,N_4386,N_4449);
or U4502 (N_4502,N_4305,N_4454);
nor U4503 (N_4503,N_4392,N_4297);
xor U4504 (N_4504,N_4254,N_4266);
xnor U4505 (N_4505,N_4471,N_4495);
nor U4506 (N_4506,N_4265,N_4430);
and U4507 (N_4507,N_4269,N_4274);
nand U4508 (N_4508,N_4380,N_4339);
nand U4509 (N_4509,N_4250,N_4442);
nor U4510 (N_4510,N_4286,N_4330);
and U4511 (N_4511,N_4289,N_4448);
or U4512 (N_4512,N_4489,N_4368);
and U4513 (N_4513,N_4315,N_4325);
xnor U4514 (N_4514,N_4393,N_4439);
or U4515 (N_4515,N_4362,N_4318);
xnor U4516 (N_4516,N_4374,N_4497);
nor U4517 (N_4517,N_4252,N_4329);
and U4518 (N_4518,N_4270,N_4264);
or U4519 (N_4519,N_4321,N_4314);
nand U4520 (N_4520,N_4405,N_4320);
nand U4521 (N_4521,N_4415,N_4313);
or U4522 (N_4522,N_4290,N_4378);
xor U4523 (N_4523,N_4451,N_4420);
xnor U4524 (N_4524,N_4434,N_4348);
nand U4525 (N_4525,N_4391,N_4444);
xnor U4526 (N_4526,N_4492,N_4465);
or U4527 (N_4527,N_4429,N_4326);
nand U4528 (N_4528,N_4372,N_4371);
and U4529 (N_4529,N_4369,N_4376);
or U4530 (N_4530,N_4436,N_4255);
nor U4531 (N_4531,N_4328,N_4364);
nand U4532 (N_4532,N_4475,N_4431);
nand U4533 (N_4533,N_4291,N_4417);
xor U4534 (N_4534,N_4443,N_4479);
xnor U4535 (N_4535,N_4384,N_4377);
nor U4536 (N_4536,N_4261,N_4394);
xor U4537 (N_4537,N_4385,N_4404);
xor U4538 (N_4538,N_4312,N_4477);
nand U4539 (N_4539,N_4301,N_4427);
xnor U4540 (N_4540,N_4402,N_4487);
nand U4541 (N_4541,N_4340,N_4423);
xnor U4542 (N_4542,N_4458,N_4303);
xnor U4543 (N_4543,N_4445,N_4310);
xor U4544 (N_4544,N_4282,N_4353);
nand U4545 (N_4545,N_4363,N_4493);
xor U4546 (N_4546,N_4316,N_4300);
xnor U4547 (N_4547,N_4412,N_4260);
and U4548 (N_4548,N_4311,N_4287);
and U4549 (N_4549,N_4324,N_4347);
and U4550 (N_4550,N_4360,N_4411);
nand U4551 (N_4551,N_4272,N_4323);
nand U4552 (N_4552,N_4466,N_4267);
and U4553 (N_4553,N_4499,N_4478);
nor U4554 (N_4554,N_4327,N_4395);
and U4555 (N_4555,N_4295,N_4370);
nand U4556 (N_4556,N_4414,N_4390);
xor U4557 (N_4557,N_4382,N_4467);
nand U4558 (N_4558,N_4284,N_4299);
nor U4559 (N_4559,N_4358,N_4413);
nand U4560 (N_4560,N_4472,N_4361);
nand U4561 (N_4561,N_4468,N_4351);
and U4562 (N_4562,N_4460,N_4331);
and U4563 (N_4563,N_4359,N_4435);
and U4564 (N_4564,N_4332,N_4432);
nor U4565 (N_4565,N_4277,N_4446);
or U4566 (N_4566,N_4279,N_4488);
nand U4567 (N_4567,N_4251,N_4426);
or U4568 (N_4568,N_4419,N_4288);
nor U4569 (N_4569,N_4438,N_4425);
nand U4570 (N_4570,N_4280,N_4457);
or U4571 (N_4571,N_4407,N_4292);
xnor U4572 (N_4572,N_4281,N_4344);
nor U4573 (N_4573,N_4498,N_4257);
nor U4574 (N_4574,N_4253,N_4268);
nand U4575 (N_4575,N_4343,N_4341);
nand U4576 (N_4576,N_4296,N_4346);
nand U4577 (N_4577,N_4470,N_4441);
nand U4578 (N_4578,N_4459,N_4456);
nor U4579 (N_4579,N_4335,N_4357);
xor U4580 (N_4580,N_4401,N_4317);
nand U4581 (N_4581,N_4271,N_4409);
xor U4582 (N_4582,N_4319,N_4480);
or U4583 (N_4583,N_4433,N_4399);
and U4584 (N_4584,N_4387,N_4494);
xor U4585 (N_4585,N_4437,N_4258);
nand U4586 (N_4586,N_4342,N_4333);
or U4587 (N_4587,N_4485,N_4388);
nor U4588 (N_4588,N_4418,N_4396);
nand U4589 (N_4589,N_4410,N_4403);
nor U4590 (N_4590,N_4476,N_4452);
or U4591 (N_4591,N_4302,N_4262);
and U4592 (N_4592,N_4322,N_4482);
nand U4593 (N_4593,N_4473,N_4496);
nor U4594 (N_4594,N_4421,N_4428);
nor U4595 (N_4595,N_4345,N_4336);
nand U4596 (N_4596,N_4307,N_4464);
xor U4597 (N_4597,N_4484,N_4440);
nor U4598 (N_4598,N_4490,N_4285);
and U4599 (N_4599,N_4453,N_4338);
and U4600 (N_4600,N_4293,N_4356);
xor U4601 (N_4601,N_4461,N_4474);
nor U4602 (N_4602,N_4354,N_4298);
xnor U4603 (N_4603,N_4416,N_4424);
nand U4604 (N_4604,N_4306,N_4400);
xnor U4605 (N_4605,N_4383,N_4469);
xor U4606 (N_4606,N_4397,N_4455);
nand U4607 (N_4607,N_4350,N_4481);
nor U4608 (N_4608,N_4447,N_4406);
nand U4609 (N_4609,N_4379,N_4275);
nand U4610 (N_4610,N_4304,N_4256);
nor U4611 (N_4611,N_4373,N_4486);
and U4612 (N_4612,N_4367,N_4463);
and U4613 (N_4613,N_4294,N_4334);
or U4614 (N_4614,N_4273,N_4491);
and U4615 (N_4615,N_4309,N_4398);
nor U4616 (N_4616,N_4381,N_4450);
xor U4617 (N_4617,N_4366,N_4355);
nor U4618 (N_4618,N_4483,N_4408);
nand U4619 (N_4619,N_4283,N_4278);
xnor U4620 (N_4620,N_4375,N_4337);
xor U4621 (N_4621,N_4308,N_4422);
nor U4622 (N_4622,N_4263,N_4389);
and U4623 (N_4623,N_4349,N_4276);
nand U4624 (N_4624,N_4365,N_4352);
or U4625 (N_4625,N_4496,N_4404);
nor U4626 (N_4626,N_4491,N_4387);
xnor U4627 (N_4627,N_4316,N_4270);
nor U4628 (N_4628,N_4358,N_4405);
nor U4629 (N_4629,N_4250,N_4295);
and U4630 (N_4630,N_4259,N_4424);
and U4631 (N_4631,N_4260,N_4362);
or U4632 (N_4632,N_4461,N_4294);
and U4633 (N_4633,N_4312,N_4486);
nand U4634 (N_4634,N_4332,N_4489);
or U4635 (N_4635,N_4257,N_4382);
xnor U4636 (N_4636,N_4452,N_4372);
nor U4637 (N_4637,N_4494,N_4331);
xnor U4638 (N_4638,N_4496,N_4260);
and U4639 (N_4639,N_4301,N_4365);
xor U4640 (N_4640,N_4296,N_4442);
nand U4641 (N_4641,N_4325,N_4473);
nor U4642 (N_4642,N_4481,N_4427);
nor U4643 (N_4643,N_4286,N_4392);
xor U4644 (N_4644,N_4376,N_4325);
nor U4645 (N_4645,N_4297,N_4488);
nand U4646 (N_4646,N_4381,N_4479);
and U4647 (N_4647,N_4281,N_4393);
and U4648 (N_4648,N_4275,N_4380);
and U4649 (N_4649,N_4325,N_4416);
nand U4650 (N_4650,N_4362,N_4290);
or U4651 (N_4651,N_4375,N_4432);
xor U4652 (N_4652,N_4470,N_4273);
nor U4653 (N_4653,N_4255,N_4378);
nor U4654 (N_4654,N_4270,N_4423);
xor U4655 (N_4655,N_4352,N_4410);
nor U4656 (N_4656,N_4416,N_4354);
and U4657 (N_4657,N_4326,N_4275);
nand U4658 (N_4658,N_4266,N_4390);
xor U4659 (N_4659,N_4294,N_4345);
or U4660 (N_4660,N_4383,N_4477);
or U4661 (N_4661,N_4373,N_4364);
xor U4662 (N_4662,N_4493,N_4330);
and U4663 (N_4663,N_4429,N_4434);
nor U4664 (N_4664,N_4253,N_4383);
xnor U4665 (N_4665,N_4253,N_4407);
nor U4666 (N_4666,N_4341,N_4495);
xor U4667 (N_4667,N_4280,N_4452);
xnor U4668 (N_4668,N_4470,N_4453);
nor U4669 (N_4669,N_4436,N_4487);
xnor U4670 (N_4670,N_4453,N_4457);
nand U4671 (N_4671,N_4328,N_4421);
xor U4672 (N_4672,N_4458,N_4343);
or U4673 (N_4673,N_4372,N_4483);
nor U4674 (N_4674,N_4281,N_4456);
xnor U4675 (N_4675,N_4325,N_4432);
or U4676 (N_4676,N_4272,N_4471);
and U4677 (N_4677,N_4481,N_4319);
xor U4678 (N_4678,N_4317,N_4297);
nand U4679 (N_4679,N_4271,N_4438);
nand U4680 (N_4680,N_4305,N_4355);
and U4681 (N_4681,N_4335,N_4399);
nand U4682 (N_4682,N_4462,N_4268);
and U4683 (N_4683,N_4258,N_4309);
or U4684 (N_4684,N_4349,N_4473);
or U4685 (N_4685,N_4263,N_4354);
or U4686 (N_4686,N_4439,N_4437);
xor U4687 (N_4687,N_4252,N_4346);
nor U4688 (N_4688,N_4264,N_4282);
and U4689 (N_4689,N_4283,N_4319);
xnor U4690 (N_4690,N_4279,N_4299);
nor U4691 (N_4691,N_4485,N_4483);
and U4692 (N_4692,N_4289,N_4406);
xnor U4693 (N_4693,N_4282,N_4344);
nand U4694 (N_4694,N_4306,N_4262);
xnor U4695 (N_4695,N_4450,N_4369);
xor U4696 (N_4696,N_4280,N_4464);
nor U4697 (N_4697,N_4342,N_4421);
nand U4698 (N_4698,N_4464,N_4385);
or U4699 (N_4699,N_4254,N_4426);
xnor U4700 (N_4700,N_4495,N_4267);
nor U4701 (N_4701,N_4397,N_4488);
nand U4702 (N_4702,N_4458,N_4262);
and U4703 (N_4703,N_4357,N_4451);
nor U4704 (N_4704,N_4382,N_4253);
nor U4705 (N_4705,N_4362,N_4375);
or U4706 (N_4706,N_4293,N_4286);
xnor U4707 (N_4707,N_4405,N_4396);
nand U4708 (N_4708,N_4320,N_4427);
or U4709 (N_4709,N_4354,N_4326);
nor U4710 (N_4710,N_4394,N_4304);
or U4711 (N_4711,N_4419,N_4385);
nor U4712 (N_4712,N_4356,N_4438);
or U4713 (N_4713,N_4273,N_4289);
or U4714 (N_4714,N_4378,N_4259);
and U4715 (N_4715,N_4281,N_4285);
nor U4716 (N_4716,N_4463,N_4459);
nor U4717 (N_4717,N_4262,N_4477);
nor U4718 (N_4718,N_4339,N_4330);
and U4719 (N_4719,N_4474,N_4329);
nor U4720 (N_4720,N_4486,N_4468);
or U4721 (N_4721,N_4409,N_4324);
nor U4722 (N_4722,N_4464,N_4277);
xor U4723 (N_4723,N_4453,N_4374);
or U4724 (N_4724,N_4290,N_4305);
nor U4725 (N_4725,N_4452,N_4315);
xor U4726 (N_4726,N_4453,N_4380);
nor U4727 (N_4727,N_4274,N_4359);
xnor U4728 (N_4728,N_4454,N_4385);
or U4729 (N_4729,N_4352,N_4367);
nand U4730 (N_4730,N_4428,N_4407);
nand U4731 (N_4731,N_4440,N_4434);
nor U4732 (N_4732,N_4310,N_4383);
and U4733 (N_4733,N_4264,N_4463);
and U4734 (N_4734,N_4424,N_4254);
and U4735 (N_4735,N_4441,N_4300);
xor U4736 (N_4736,N_4331,N_4372);
nand U4737 (N_4737,N_4493,N_4333);
nand U4738 (N_4738,N_4378,N_4425);
nand U4739 (N_4739,N_4268,N_4394);
and U4740 (N_4740,N_4300,N_4375);
and U4741 (N_4741,N_4491,N_4469);
nand U4742 (N_4742,N_4370,N_4405);
and U4743 (N_4743,N_4436,N_4316);
nor U4744 (N_4744,N_4285,N_4433);
and U4745 (N_4745,N_4328,N_4300);
and U4746 (N_4746,N_4275,N_4384);
and U4747 (N_4747,N_4495,N_4433);
and U4748 (N_4748,N_4274,N_4351);
and U4749 (N_4749,N_4437,N_4401);
and U4750 (N_4750,N_4743,N_4655);
and U4751 (N_4751,N_4611,N_4543);
xor U4752 (N_4752,N_4689,N_4568);
nand U4753 (N_4753,N_4511,N_4713);
or U4754 (N_4754,N_4656,N_4719);
nor U4755 (N_4755,N_4506,N_4583);
or U4756 (N_4756,N_4605,N_4650);
xor U4757 (N_4757,N_4678,N_4571);
and U4758 (N_4758,N_4704,N_4594);
nor U4759 (N_4759,N_4586,N_4654);
or U4760 (N_4760,N_4521,N_4552);
or U4761 (N_4761,N_4556,N_4562);
and U4762 (N_4762,N_4544,N_4675);
xnor U4763 (N_4763,N_4684,N_4693);
nor U4764 (N_4764,N_4739,N_4537);
and U4765 (N_4765,N_4580,N_4603);
and U4766 (N_4766,N_4697,N_4664);
or U4767 (N_4767,N_4634,N_4748);
xor U4768 (N_4768,N_4732,N_4618);
xor U4769 (N_4769,N_4519,N_4627);
nor U4770 (N_4770,N_4642,N_4516);
nor U4771 (N_4771,N_4557,N_4622);
and U4772 (N_4772,N_4589,N_4679);
and U4773 (N_4773,N_4645,N_4542);
and U4774 (N_4774,N_4631,N_4529);
and U4775 (N_4775,N_4724,N_4710);
xor U4776 (N_4776,N_4698,N_4527);
and U4777 (N_4777,N_4620,N_4610);
nor U4778 (N_4778,N_4700,N_4660);
nor U4779 (N_4779,N_4503,N_4615);
nand U4780 (N_4780,N_4716,N_4646);
nand U4781 (N_4781,N_4598,N_4595);
nor U4782 (N_4782,N_4515,N_4626);
nor U4783 (N_4783,N_4613,N_4590);
nand U4784 (N_4784,N_4721,N_4623);
nor U4785 (N_4785,N_4676,N_4549);
or U4786 (N_4786,N_4674,N_4536);
nor U4787 (N_4787,N_4741,N_4601);
and U4788 (N_4788,N_4538,N_4709);
xor U4789 (N_4789,N_4682,N_4535);
nand U4790 (N_4790,N_4600,N_4517);
and U4791 (N_4791,N_4602,N_4747);
xnor U4792 (N_4792,N_4670,N_4680);
xnor U4793 (N_4793,N_4632,N_4541);
xor U4794 (N_4794,N_4746,N_4728);
nand U4795 (N_4795,N_4523,N_4577);
or U4796 (N_4796,N_4720,N_4696);
nor U4797 (N_4797,N_4560,N_4559);
xor U4798 (N_4798,N_4702,N_4635);
xnor U4799 (N_4799,N_4715,N_4637);
xnor U4800 (N_4800,N_4553,N_4566);
nor U4801 (N_4801,N_4729,N_4666);
or U4802 (N_4802,N_4578,N_4653);
nor U4803 (N_4803,N_4596,N_4640);
and U4804 (N_4804,N_4539,N_4639);
or U4805 (N_4805,N_4735,N_4591);
nand U4806 (N_4806,N_4722,N_4652);
nor U4807 (N_4807,N_4636,N_4737);
nor U4808 (N_4808,N_4687,N_4545);
xnor U4809 (N_4809,N_4727,N_4744);
nor U4810 (N_4810,N_4692,N_4621);
and U4811 (N_4811,N_4688,N_4582);
nor U4812 (N_4812,N_4712,N_4708);
nand U4813 (N_4813,N_4749,N_4649);
xnor U4814 (N_4814,N_4567,N_4573);
or U4815 (N_4815,N_4657,N_4608);
or U4816 (N_4816,N_4604,N_4561);
nand U4817 (N_4817,N_4592,N_4619);
and U4818 (N_4818,N_4624,N_4528);
and U4819 (N_4819,N_4504,N_4644);
nor U4820 (N_4820,N_4683,N_4555);
nand U4821 (N_4821,N_4699,N_4677);
and U4822 (N_4822,N_4514,N_4659);
or U4823 (N_4823,N_4671,N_4612);
nand U4824 (N_4824,N_4548,N_4706);
and U4825 (N_4825,N_4707,N_4672);
nor U4826 (N_4826,N_4616,N_4597);
or U4827 (N_4827,N_4518,N_4738);
and U4828 (N_4828,N_4701,N_4507);
and U4829 (N_4829,N_4647,N_4530);
nor U4830 (N_4830,N_4574,N_4584);
xnor U4831 (N_4831,N_4651,N_4691);
nor U4832 (N_4832,N_4673,N_4726);
nor U4833 (N_4833,N_4547,N_4725);
xnor U4834 (N_4834,N_4513,N_4588);
or U4835 (N_4835,N_4581,N_4551);
nand U4836 (N_4836,N_4563,N_4531);
xnor U4837 (N_4837,N_4662,N_4607);
nand U4838 (N_4838,N_4525,N_4606);
xnor U4839 (N_4839,N_4711,N_4694);
and U4840 (N_4840,N_4730,N_4629);
or U4841 (N_4841,N_4564,N_4714);
nand U4842 (N_4842,N_4695,N_4512);
xnor U4843 (N_4843,N_4500,N_4630);
and U4844 (N_4844,N_4643,N_4576);
xnor U4845 (N_4845,N_4508,N_4731);
xnor U4846 (N_4846,N_4740,N_4572);
nor U4847 (N_4847,N_4501,N_4593);
or U4848 (N_4848,N_4742,N_4703);
nor U4849 (N_4849,N_4718,N_4625);
and U4850 (N_4850,N_4579,N_4641);
nor U4851 (N_4851,N_4690,N_4505);
nor U4852 (N_4852,N_4587,N_4705);
or U4853 (N_4853,N_4734,N_4736);
xnor U4854 (N_4854,N_4524,N_4546);
xor U4855 (N_4855,N_4658,N_4575);
nor U4856 (N_4856,N_4520,N_4614);
nor U4857 (N_4857,N_4526,N_4522);
or U4858 (N_4858,N_4628,N_4509);
xor U4859 (N_4859,N_4633,N_4558);
and U4860 (N_4860,N_4668,N_4617);
xnor U4861 (N_4861,N_4599,N_4745);
or U4862 (N_4862,N_4533,N_4685);
nor U4863 (N_4863,N_4665,N_4540);
nor U4864 (N_4864,N_4554,N_4585);
nand U4865 (N_4865,N_4723,N_4550);
and U4866 (N_4866,N_4502,N_4565);
nor U4867 (N_4867,N_4570,N_4686);
xnor U4868 (N_4868,N_4681,N_4733);
xor U4869 (N_4869,N_4534,N_4532);
xor U4870 (N_4870,N_4667,N_4510);
nor U4871 (N_4871,N_4638,N_4669);
xnor U4872 (N_4872,N_4717,N_4609);
or U4873 (N_4873,N_4661,N_4569);
nand U4874 (N_4874,N_4663,N_4648);
or U4875 (N_4875,N_4639,N_4631);
xor U4876 (N_4876,N_4657,N_4730);
and U4877 (N_4877,N_4748,N_4722);
and U4878 (N_4878,N_4674,N_4518);
and U4879 (N_4879,N_4527,N_4507);
or U4880 (N_4880,N_4698,N_4505);
and U4881 (N_4881,N_4733,N_4584);
or U4882 (N_4882,N_4549,N_4503);
and U4883 (N_4883,N_4630,N_4685);
or U4884 (N_4884,N_4572,N_4558);
or U4885 (N_4885,N_4603,N_4737);
and U4886 (N_4886,N_4519,N_4621);
nor U4887 (N_4887,N_4680,N_4666);
xor U4888 (N_4888,N_4655,N_4578);
or U4889 (N_4889,N_4614,N_4506);
or U4890 (N_4890,N_4525,N_4580);
nand U4891 (N_4891,N_4587,N_4573);
and U4892 (N_4892,N_4567,N_4743);
nor U4893 (N_4893,N_4711,N_4598);
or U4894 (N_4894,N_4639,N_4714);
nor U4895 (N_4895,N_4620,N_4561);
xnor U4896 (N_4896,N_4567,N_4683);
or U4897 (N_4897,N_4633,N_4666);
nor U4898 (N_4898,N_4634,N_4696);
and U4899 (N_4899,N_4531,N_4513);
nand U4900 (N_4900,N_4504,N_4678);
and U4901 (N_4901,N_4620,N_4654);
nor U4902 (N_4902,N_4596,N_4579);
xor U4903 (N_4903,N_4502,N_4558);
nand U4904 (N_4904,N_4733,N_4641);
xor U4905 (N_4905,N_4661,N_4662);
and U4906 (N_4906,N_4745,N_4554);
nor U4907 (N_4907,N_4642,N_4733);
nand U4908 (N_4908,N_4523,N_4654);
nand U4909 (N_4909,N_4510,N_4542);
and U4910 (N_4910,N_4653,N_4609);
nor U4911 (N_4911,N_4696,N_4673);
and U4912 (N_4912,N_4692,N_4609);
nand U4913 (N_4913,N_4654,N_4573);
nor U4914 (N_4914,N_4519,N_4561);
nand U4915 (N_4915,N_4731,N_4741);
and U4916 (N_4916,N_4749,N_4569);
or U4917 (N_4917,N_4703,N_4626);
xor U4918 (N_4918,N_4599,N_4636);
xnor U4919 (N_4919,N_4710,N_4613);
xnor U4920 (N_4920,N_4577,N_4592);
nor U4921 (N_4921,N_4698,N_4738);
or U4922 (N_4922,N_4677,N_4604);
and U4923 (N_4923,N_4639,N_4548);
nor U4924 (N_4924,N_4714,N_4589);
and U4925 (N_4925,N_4514,N_4641);
xor U4926 (N_4926,N_4542,N_4703);
nand U4927 (N_4927,N_4614,N_4552);
nor U4928 (N_4928,N_4512,N_4745);
nor U4929 (N_4929,N_4740,N_4570);
nand U4930 (N_4930,N_4588,N_4681);
or U4931 (N_4931,N_4611,N_4549);
or U4932 (N_4932,N_4738,N_4719);
or U4933 (N_4933,N_4691,N_4519);
nor U4934 (N_4934,N_4733,N_4614);
xnor U4935 (N_4935,N_4545,N_4505);
nor U4936 (N_4936,N_4569,N_4622);
and U4937 (N_4937,N_4695,N_4727);
nand U4938 (N_4938,N_4541,N_4742);
or U4939 (N_4939,N_4730,N_4553);
nand U4940 (N_4940,N_4715,N_4515);
and U4941 (N_4941,N_4704,N_4730);
nor U4942 (N_4942,N_4713,N_4728);
nor U4943 (N_4943,N_4654,N_4707);
nor U4944 (N_4944,N_4571,N_4745);
and U4945 (N_4945,N_4602,N_4619);
and U4946 (N_4946,N_4707,N_4699);
nand U4947 (N_4947,N_4570,N_4607);
or U4948 (N_4948,N_4588,N_4662);
nand U4949 (N_4949,N_4700,N_4626);
and U4950 (N_4950,N_4741,N_4621);
or U4951 (N_4951,N_4707,N_4568);
or U4952 (N_4952,N_4721,N_4643);
and U4953 (N_4953,N_4656,N_4660);
nor U4954 (N_4954,N_4531,N_4705);
nand U4955 (N_4955,N_4700,N_4683);
and U4956 (N_4956,N_4740,N_4580);
xnor U4957 (N_4957,N_4747,N_4625);
and U4958 (N_4958,N_4739,N_4595);
xor U4959 (N_4959,N_4665,N_4594);
nand U4960 (N_4960,N_4514,N_4597);
nor U4961 (N_4961,N_4537,N_4705);
and U4962 (N_4962,N_4673,N_4560);
and U4963 (N_4963,N_4620,N_4670);
and U4964 (N_4964,N_4566,N_4568);
xnor U4965 (N_4965,N_4659,N_4619);
xnor U4966 (N_4966,N_4708,N_4536);
nor U4967 (N_4967,N_4593,N_4646);
nor U4968 (N_4968,N_4629,N_4508);
or U4969 (N_4969,N_4673,N_4559);
xor U4970 (N_4970,N_4541,N_4723);
or U4971 (N_4971,N_4583,N_4607);
and U4972 (N_4972,N_4517,N_4665);
or U4973 (N_4973,N_4559,N_4579);
or U4974 (N_4974,N_4556,N_4702);
xnor U4975 (N_4975,N_4658,N_4724);
or U4976 (N_4976,N_4733,N_4599);
nand U4977 (N_4977,N_4616,N_4705);
nand U4978 (N_4978,N_4718,N_4586);
xor U4979 (N_4979,N_4725,N_4501);
nor U4980 (N_4980,N_4651,N_4504);
and U4981 (N_4981,N_4655,N_4523);
nand U4982 (N_4982,N_4554,N_4647);
nand U4983 (N_4983,N_4674,N_4641);
and U4984 (N_4984,N_4728,N_4597);
nand U4985 (N_4985,N_4728,N_4565);
and U4986 (N_4986,N_4596,N_4700);
or U4987 (N_4987,N_4540,N_4668);
nor U4988 (N_4988,N_4717,N_4561);
nand U4989 (N_4989,N_4697,N_4685);
and U4990 (N_4990,N_4657,N_4721);
xor U4991 (N_4991,N_4549,N_4661);
and U4992 (N_4992,N_4667,N_4719);
nor U4993 (N_4993,N_4738,N_4617);
and U4994 (N_4994,N_4615,N_4561);
xnor U4995 (N_4995,N_4574,N_4536);
xnor U4996 (N_4996,N_4664,N_4693);
and U4997 (N_4997,N_4579,N_4707);
or U4998 (N_4998,N_4549,N_4586);
xnor U4999 (N_4999,N_4634,N_4653);
xor U5000 (N_5000,N_4937,N_4958);
nor U5001 (N_5001,N_4809,N_4798);
xnor U5002 (N_5002,N_4842,N_4818);
and U5003 (N_5003,N_4873,N_4918);
and U5004 (N_5004,N_4835,N_4976);
nor U5005 (N_5005,N_4804,N_4952);
nor U5006 (N_5006,N_4778,N_4864);
nand U5007 (N_5007,N_4853,N_4838);
nand U5008 (N_5008,N_4961,N_4896);
and U5009 (N_5009,N_4993,N_4841);
xor U5010 (N_5010,N_4762,N_4765);
nand U5011 (N_5011,N_4985,N_4795);
nand U5012 (N_5012,N_4845,N_4895);
nand U5013 (N_5013,N_4783,N_4999);
or U5014 (N_5014,N_4874,N_4965);
or U5015 (N_5015,N_4865,N_4862);
nor U5016 (N_5016,N_4801,N_4988);
xnor U5017 (N_5017,N_4764,N_4870);
xnor U5018 (N_5018,N_4849,N_4806);
nand U5019 (N_5019,N_4984,N_4911);
nand U5020 (N_5020,N_4854,N_4954);
nor U5021 (N_5021,N_4970,N_4782);
or U5022 (N_5022,N_4951,N_4772);
xor U5023 (N_5023,N_4855,N_4940);
nand U5024 (N_5024,N_4850,N_4894);
or U5025 (N_5025,N_4755,N_4964);
xnor U5026 (N_5026,N_4812,N_4750);
xor U5027 (N_5027,N_4761,N_4968);
xnor U5028 (N_5028,N_4959,N_4935);
or U5029 (N_5029,N_4792,N_4986);
nor U5030 (N_5030,N_4876,N_4929);
nor U5031 (N_5031,N_4846,N_4878);
nand U5032 (N_5032,N_4899,N_4913);
and U5033 (N_5033,N_4791,N_4903);
xnor U5034 (N_5034,N_4919,N_4973);
or U5035 (N_5035,N_4826,N_4828);
nor U5036 (N_5036,N_4852,N_4774);
nor U5037 (N_5037,N_4957,N_4861);
xor U5038 (N_5038,N_4816,N_4923);
and U5039 (N_5039,N_4763,N_4824);
nor U5040 (N_5040,N_4757,N_4910);
or U5041 (N_5041,N_4875,N_4802);
and U5042 (N_5042,N_4770,N_4981);
and U5043 (N_5043,N_4920,N_4889);
xor U5044 (N_5044,N_4946,N_4904);
or U5045 (N_5045,N_4839,N_4863);
xnor U5046 (N_5046,N_4837,N_4921);
nor U5047 (N_5047,N_4989,N_4974);
nand U5048 (N_5048,N_4814,N_4925);
and U5049 (N_5049,N_4934,N_4956);
nor U5050 (N_5050,N_4942,N_4827);
nor U5051 (N_5051,N_4927,N_4833);
xnor U5052 (N_5052,N_4858,N_4786);
nor U5053 (N_5053,N_4893,N_4847);
or U5054 (N_5054,N_4992,N_4982);
nor U5055 (N_5055,N_4898,N_4867);
nand U5056 (N_5056,N_4800,N_4758);
and U5057 (N_5057,N_4796,N_4787);
nor U5058 (N_5058,N_4978,N_4836);
nand U5059 (N_5059,N_4781,N_4834);
nand U5060 (N_5060,N_4779,N_4752);
xor U5061 (N_5061,N_4759,N_4817);
nand U5062 (N_5062,N_4784,N_4953);
or U5063 (N_5063,N_4944,N_4912);
nor U5064 (N_5064,N_4820,N_4883);
nand U5065 (N_5065,N_4829,N_4901);
and U5066 (N_5066,N_4995,N_4859);
nor U5067 (N_5067,N_4907,N_4790);
nor U5068 (N_5068,N_4780,N_4971);
xnor U5069 (N_5069,N_4805,N_4897);
nand U5070 (N_5070,N_4821,N_4939);
nand U5071 (N_5071,N_4926,N_4916);
nor U5072 (N_5072,N_4872,N_4905);
nand U5073 (N_5073,N_4928,N_4768);
nor U5074 (N_5074,N_4866,N_4868);
xnor U5075 (N_5075,N_4983,N_4808);
nor U5076 (N_5076,N_4793,N_4760);
or U5077 (N_5077,N_4980,N_4998);
and U5078 (N_5078,N_4769,N_4877);
nor U5079 (N_5079,N_4949,N_4888);
and U5080 (N_5080,N_4825,N_4831);
nor U5081 (N_5081,N_4963,N_4788);
nor U5082 (N_5082,N_4914,N_4902);
nand U5083 (N_5083,N_4766,N_4931);
nor U5084 (N_5084,N_4991,N_4811);
and U5085 (N_5085,N_4856,N_4892);
and U5086 (N_5086,N_4884,N_4810);
nand U5087 (N_5087,N_4936,N_4751);
nand U5088 (N_5088,N_4881,N_4794);
and U5089 (N_5089,N_4922,N_4756);
and U5090 (N_5090,N_4987,N_4930);
or U5091 (N_5091,N_4979,N_4832);
nand U5092 (N_5092,N_4933,N_4945);
xor U5093 (N_5093,N_4917,N_4823);
and U5094 (N_5094,N_4785,N_4767);
and U5095 (N_5095,N_4947,N_4773);
xnor U5096 (N_5096,N_4789,N_4776);
xnor U5097 (N_5097,N_4955,N_4819);
and U5098 (N_5098,N_4799,N_4880);
nand U5099 (N_5099,N_4891,N_4851);
and U5100 (N_5100,N_4950,N_4822);
nor U5101 (N_5101,N_4777,N_4924);
or U5102 (N_5102,N_4960,N_4938);
nor U5103 (N_5103,N_4885,N_4797);
nor U5104 (N_5104,N_4994,N_4909);
nand U5105 (N_5105,N_4857,N_4943);
and U5106 (N_5106,N_4879,N_4807);
and U5107 (N_5107,N_4860,N_4886);
xor U5108 (N_5108,N_4915,N_4941);
xnor U5109 (N_5109,N_4900,N_4813);
nand U5110 (N_5110,N_4753,N_4887);
or U5111 (N_5111,N_4948,N_4869);
nor U5112 (N_5112,N_4962,N_4932);
and U5113 (N_5113,N_4890,N_4966);
or U5114 (N_5114,N_4754,N_4997);
xor U5115 (N_5115,N_4990,N_4969);
and U5116 (N_5116,N_4972,N_4803);
nand U5117 (N_5117,N_4871,N_4830);
nor U5118 (N_5118,N_4996,N_4906);
or U5119 (N_5119,N_4848,N_4775);
nand U5120 (N_5120,N_4967,N_4975);
or U5121 (N_5121,N_4815,N_4908);
nand U5122 (N_5122,N_4977,N_4882);
nor U5123 (N_5123,N_4843,N_4771);
xor U5124 (N_5124,N_4840,N_4844);
nor U5125 (N_5125,N_4972,N_4966);
nor U5126 (N_5126,N_4854,N_4994);
xor U5127 (N_5127,N_4977,N_4815);
nor U5128 (N_5128,N_4878,N_4763);
xor U5129 (N_5129,N_4876,N_4978);
and U5130 (N_5130,N_4815,N_4768);
or U5131 (N_5131,N_4896,N_4765);
and U5132 (N_5132,N_4832,N_4957);
and U5133 (N_5133,N_4751,N_4759);
xor U5134 (N_5134,N_4843,N_4755);
xor U5135 (N_5135,N_4853,N_4768);
nor U5136 (N_5136,N_4757,N_4783);
nor U5137 (N_5137,N_4946,N_4755);
nand U5138 (N_5138,N_4889,N_4859);
nand U5139 (N_5139,N_4865,N_4853);
xor U5140 (N_5140,N_4840,N_4786);
nor U5141 (N_5141,N_4925,N_4897);
xnor U5142 (N_5142,N_4998,N_4972);
and U5143 (N_5143,N_4859,N_4756);
and U5144 (N_5144,N_4976,N_4836);
nand U5145 (N_5145,N_4803,N_4805);
nor U5146 (N_5146,N_4776,N_4801);
xor U5147 (N_5147,N_4832,N_4934);
nor U5148 (N_5148,N_4860,N_4760);
and U5149 (N_5149,N_4967,N_4855);
and U5150 (N_5150,N_4781,N_4800);
xor U5151 (N_5151,N_4901,N_4993);
nor U5152 (N_5152,N_4872,N_4775);
nand U5153 (N_5153,N_4882,N_4862);
nand U5154 (N_5154,N_4878,N_4830);
xor U5155 (N_5155,N_4923,N_4832);
xor U5156 (N_5156,N_4887,N_4807);
nor U5157 (N_5157,N_4755,N_4771);
or U5158 (N_5158,N_4967,N_4795);
nor U5159 (N_5159,N_4778,N_4904);
or U5160 (N_5160,N_4860,N_4905);
xor U5161 (N_5161,N_4961,N_4768);
or U5162 (N_5162,N_4942,N_4851);
xor U5163 (N_5163,N_4966,N_4813);
or U5164 (N_5164,N_4968,N_4869);
nor U5165 (N_5165,N_4850,N_4805);
and U5166 (N_5166,N_4921,N_4754);
nand U5167 (N_5167,N_4759,N_4782);
nor U5168 (N_5168,N_4999,N_4934);
and U5169 (N_5169,N_4986,N_4800);
and U5170 (N_5170,N_4894,N_4769);
or U5171 (N_5171,N_4830,N_4815);
nand U5172 (N_5172,N_4752,N_4941);
xor U5173 (N_5173,N_4819,N_4805);
or U5174 (N_5174,N_4848,N_4900);
or U5175 (N_5175,N_4847,N_4940);
and U5176 (N_5176,N_4830,N_4963);
xor U5177 (N_5177,N_4764,N_4938);
or U5178 (N_5178,N_4863,N_4898);
or U5179 (N_5179,N_4821,N_4990);
nor U5180 (N_5180,N_4873,N_4989);
or U5181 (N_5181,N_4979,N_4850);
xor U5182 (N_5182,N_4779,N_4871);
or U5183 (N_5183,N_4812,N_4797);
nand U5184 (N_5184,N_4874,N_4993);
xor U5185 (N_5185,N_4834,N_4803);
and U5186 (N_5186,N_4939,N_4767);
xor U5187 (N_5187,N_4959,N_4846);
and U5188 (N_5188,N_4869,N_4895);
xnor U5189 (N_5189,N_4865,N_4795);
xnor U5190 (N_5190,N_4836,N_4817);
nor U5191 (N_5191,N_4878,N_4923);
nand U5192 (N_5192,N_4906,N_4806);
nand U5193 (N_5193,N_4762,N_4948);
and U5194 (N_5194,N_4815,N_4970);
nand U5195 (N_5195,N_4814,N_4828);
and U5196 (N_5196,N_4997,N_4917);
nand U5197 (N_5197,N_4847,N_4777);
or U5198 (N_5198,N_4988,N_4778);
nor U5199 (N_5199,N_4811,N_4910);
nand U5200 (N_5200,N_4854,N_4937);
and U5201 (N_5201,N_4919,N_4776);
or U5202 (N_5202,N_4779,N_4781);
or U5203 (N_5203,N_4863,N_4923);
and U5204 (N_5204,N_4870,N_4791);
and U5205 (N_5205,N_4875,N_4765);
xnor U5206 (N_5206,N_4754,N_4913);
nor U5207 (N_5207,N_4872,N_4898);
nand U5208 (N_5208,N_4934,N_4812);
nand U5209 (N_5209,N_4892,N_4979);
xnor U5210 (N_5210,N_4941,N_4788);
nand U5211 (N_5211,N_4822,N_4881);
and U5212 (N_5212,N_4845,N_4810);
nor U5213 (N_5213,N_4953,N_4816);
xor U5214 (N_5214,N_4930,N_4801);
or U5215 (N_5215,N_4964,N_4842);
or U5216 (N_5216,N_4941,N_4810);
and U5217 (N_5217,N_4963,N_4942);
xnor U5218 (N_5218,N_4918,N_4909);
nor U5219 (N_5219,N_4794,N_4861);
nor U5220 (N_5220,N_4871,N_4784);
xor U5221 (N_5221,N_4781,N_4952);
nand U5222 (N_5222,N_4858,N_4803);
xor U5223 (N_5223,N_4962,N_4792);
or U5224 (N_5224,N_4781,N_4757);
xor U5225 (N_5225,N_4886,N_4985);
or U5226 (N_5226,N_4929,N_4931);
or U5227 (N_5227,N_4930,N_4838);
nand U5228 (N_5228,N_4814,N_4847);
or U5229 (N_5229,N_4916,N_4998);
and U5230 (N_5230,N_4900,N_4795);
and U5231 (N_5231,N_4953,N_4945);
and U5232 (N_5232,N_4926,N_4958);
xor U5233 (N_5233,N_4901,N_4974);
xnor U5234 (N_5234,N_4914,N_4814);
and U5235 (N_5235,N_4936,N_4795);
and U5236 (N_5236,N_4978,N_4822);
and U5237 (N_5237,N_4838,N_4924);
xor U5238 (N_5238,N_4890,N_4987);
nand U5239 (N_5239,N_4881,N_4833);
and U5240 (N_5240,N_4939,N_4831);
xor U5241 (N_5241,N_4861,N_4808);
nor U5242 (N_5242,N_4881,N_4933);
nor U5243 (N_5243,N_4768,N_4761);
and U5244 (N_5244,N_4906,N_4892);
and U5245 (N_5245,N_4792,N_4808);
or U5246 (N_5246,N_4841,N_4934);
nand U5247 (N_5247,N_4931,N_4856);
xnor U5248 (N_5248,N_4812,N_4874);
nand U5249 (N_5249,N_4760,N_4823);
or U5250 (N_5250,N_5064,N_5192);
xor U5251 (N_5251,N_5068,N_5241);
nand U5252 (N_5252,N_5066,N_5073);
nor U5253 (N_5253,N_5223,N_5188);
or U5254 (N_5254,N_5141,N_5246);
nand U5255 (N_5255,N_5139,N_5119);
and U5256 (N_5256,N_5009,N_5130);
xor U5257 (N_5257,N_5194,N_5098);
nor U5258 (N_5258,N_5206,N_5146);
xor U5259 (N_5259,N_5237,N_5214);
nand U5260 (N_5260,N_5031,N_5048);
nand U5261 (N_5261,N_5035,N_5080);
or U5262 (N_5262,N_5091,N_5097);
and U5263 (N_5263,N_5109,N_5126);
xnor U5264 (N_5264,N_5199,N_5037);
xor U5265 (N_5265,N_5079,N_5221);
xnor U5266 (N_5266,N_5142,N_5202);
or U5267 (N_5267,N_5195,N_5220);
xnor U5268 (N_5268,N_5183,N_5002);
and U5269 (N_5269,N_5108,N_5170);
and U5270 (N_5270,N_5049,N_5036);
xnor U5271 (N_5271,N_5018,N_5124);
and U5272 (N_5272,N_5205,N_5051);
and U5273 (N_5273,N_5081,N_5006);
nor U5274 (N_5274,N_5065,N_5063);
and U5275 (N_5275,N_5084,N_5076);
or U5276 (N_5276,N_5129,N_5060);
xnor U5277 (N_5277,N_5157,N_5112);
and U5278 (N_5278,N_5054,N_5083);
xor U5279 (N_5279,N_5182,N_5247);
or U5280 (N_5280,N_5026,N_5125);
or U5281 (N_5281,N_5238,N_5216);
nor U5282 (N_5282,N_5011,N_5229);
nand U5283 (N_5283,N_5045,N_5093);
and U5284 (N_5284,N_5027,N_5184);
xor U5285 (N_5285,N_5209,N_5160);
xor U5286 (N_5286,N_5143,N_5193);
xnor U5287 (N_5287,N_5069,N_5210);
nor U5288 (N_5288,N_5015,N_5168);
nand U5289 (N_5289,N_5057,N_5075);
and U5290 (N_5290,N_5133,N_5029);
nor U5291 (N_5291,N_5013,N_5189);
nor U5292 (N_5292,N_5245,N_5115);
and U5293 (N_5293,N_5165,N_5152);
and U5294 (N_5294,N_5086,N_5092);
xor U5295 (N_5295,N_5070,N_5175);
or U5296 (N_5296,N_5116,N_5138);
and U5297 (N_5297,N_5173,N_5236);
and U5298 (N_5298,N_5020,N_5059);
or U5299 (N_5299,N_5094,N_5044);
and U5300 (N_5300,N_5019,N_5024);
or U5301 (N_5301,N_5185,N_5101);
xnor U5302 (N_5302,N_5230,N_5196);
or U5303 (N_5303,N_5147,N_5227);
nand U5304 (N_5304,N_5067,N_5095);
xnor U5305 (N_5305,N_5226,N_5163);
nand U5306 (N_5306,N_5181,N_5178);
nor U5307 (N_5307,N_5113,N_5131);
and U5308 (N_5308,N_5132,N_5148);
and U5309 (N_5309,N_5151,N_5034);
xor U5310 (N_5310,N_5077,N_5100);
xor U5311 (N_5311,N_5212,N_5204);
and U5312 (N_5312,N_5121,N_5243);
nand U5313 (N_5313,N_5104,N_5242);
xnor U5314 (N_5314,N_5117,N_5174);
nor U5315 (N_5315,N_5200,N_5222);
xor U5316 (N_5316,N_5235,N_5047);
xnor U5317 (N_5317,N_5127,N_5040);
nor U5318 (N_5318,N_5128,N_5158);
nor U5319 (N_5319,N_5111,N_5078);
xnor U5320 (N_5320,N_5213,N_5118);
xnor U5321 (N_5321,N_5023,N_5218);
xnor U5322 (N_5322,N_5180,N_5089);
or U5323 (N_5323,N_5203,N_5231);
and U5324 (N_5324,N_5186,N_5215);
or U5325 (N_5325,N_5233,N_5198);
nand U5326 (N_5326,N_5055,N_5032);
or U5327 (N_5327,N_5149,N_5058);
and U5328 (N_5328,N_5176,N_5038);
nor U5329 (N_5329,N_5062,N_5150);
and U5330 (N_5330,N_5000,N_5155);
xor U5331 (N_5331,N_5219,N_5021);
nor U5332 (N_5332,N_5012,N_5056);
or U5333 (N_5333,N_5052,N_5106);
and U5334 (N_5334,N_5022,N_5033);
xor U5335 (N_5335,N_5122,N_5090);
xnor U5336 (N_5336,N_5102,N_5234);
nor U5337 (N_5337,N_5136,N_5211);
nand U5338 (N_5338,N_5053,N_5010);
xor U5339 (N_5339,N_5028,N_5166);
or U5340 (N_5340,N_5004,N_5161);
nand U5341 (N_5341,N_5082,N_5096);
nor U5342 (N_5342,N_5114,N_5046);
or U5343 (N_5343,N_5003,N_5014);
xor U5344 (N_5344,N_5249,N_5187);
or U5345 (N_5345,N_5041,N_5232);
xor U5346 (N_5346,N_5007,N_5153);
nor U5347 (N_5347,N_5072,N_5074);
xnor U5348 (N_5348,N_5179,N_5201);
nand U5349 (N_5349,N_5123,N_5239);
and U5350 (N_5350,N_5008,N_5061);
nand U5351 (N_5351,N_5087,N_5099);
and U5352 (N_5352,N_5167,N_5154);
or U5353 (N_5353,N_5144,N_5164);
and U5354 (N_5354,N_5197,N_5145);
and U5355 (N_5355,N_5207,N_5191);
xor U5356 (N_5356,N_5025,N_5172);
xnor U5357 (N_5357,N_5171,N_5085);
and U5358 (N_5358,N_5042,N_5244);
or U5359 (N_5359,N_5224,N_5162);
or U5360 (N_5360,N_5016,N_5071);
nand U5361 (N_5361,N_5169,N_5248);
and U5362 (N_5362,N_5043,N_5225);
and U5363 (N_5363,N_5039,N_5005);
and U5364 (N_5364,N_5228,N_5159);
xnor U5365 (N_5365,N_5190,N_5140);
nand U5366 (N_5366,N_5134,N_5001);
or U5367 (N_5367,N_5217,N_5120);
or U5368 (N_5368,N_5103,N_5088);
or U5369 (N_5369,N_5030,N_5208);
and U5370 (N_5370,N_5107,N_5177);
or U5371 (N_5371,N_5137,N_5017);
xnor U5372 (N_5372,N_5110,N_5156);
nand U5373 (N_5373,N_5135,N_5105);
and U5374 (N_5374,N_5050,N_5240);
nor U5375 (N_5375,N_5016,N_5022);
xnor U5376 (N_5376,N_5022,N_5115);
and U5377 (N_5377,N_5174,N_5100);
or U5378 (N_5378,N_5199,N_5177);
nor U5379 (N_5379,N_5024,N_5080);
xor U5380 (N_5380,N_5034,N_5017);
nand U5381 (N_5381,N_5057,N_5064);
xor U5382 (N_5382,N_5051,N_5092);
or U5383 (N_5383,N_5006,N_5164);
nor U5384 (N_5384,N_5096,N_5190);
or U5385 (N_5385,N_5211,N_5207);
nand U5386 (N_5386,N_5170,N_5029);
and U5387 (N_5387,N_5105,N_5197);
nor U5388 (N_5388,N_5000,N_5248);
nor U5389 (N_5389,N_5114,N_5045);
and U5390 (N_5390,N_5081,N_5157);
nor U5391 (N_5391,N_5039,N_5226);
nor U5392 (N_5392,N_5089,N_5025);
nor U5393 (N_5393,N_5060,N_5226);
nand U5394 (N_5394,N_5095,N_5136);
nor U5395 (N_5395,N_5091,N_5013);
or U5396 (N_5396,N_5097,N_5200);
nand U5397 (N_5397,N_5043,N_5246);
and U5398 (N_5398,N_5218,N_5030);
nor U5399 (N_5399,N_5000,N_5224);
xnor U5400 (N_5400,N_5004,N_5121);
xor U5401 (N_5401,N_5151,N_5165);
xnor U5402 (N_5402,N_5163,N_5141);
or U5403 (N_5403,N_5128,N_5245);
nor U5404 (N_5404,N_5168,N_5066);
nand U5405 (N_5405,N_5142,N_5013);
and U5406 (N_5406,N_5055,N_5050);
or U5407 (N_5407,N_5221,N_5061);
nor U5408 (N_5408,N_5243,N_5164);
nor U5409 (N_5409,N_5099,N_5178);
nor U5410 (N_5410,N_5021,N_5236);
nor U5411 (N_5411,N_5052,N_5138);
and U5412 (N_5412,N_5236,N_5024);
nand U5413 (N_5413,N_5238,N_5136);
nor U5414 (N_5414,N_5235,N_5066);
and U5415 (N_5415,N_5053,N_5197);
or U5416 (N_5416,N_5161,N_5186);
and U5417 (N_5417,N_5081,N_5248);
or U5418 (N_5418,N_5222,N_5137);
xnor U5419 (N_5419,N_5156,N_5207);
nand U5420 (N_5420,N_5085,N_5155);
nor U5421 (N_5421,N_5151,N_5171);
or U5422 (N_5422,N_5034,N_5140);
xnor U5423 (N_5423,N_5136,N_5150);
nor U5424 (N_5424,N_5093,N_5213);
xnor U5425 (N_5425,N_5087,N_5212);
nand U5426 (N_5426,N_5021,N_5100);
and U5427 (N_5427,N_5171,N_5058);
or U5428 (N_5428,N_5226,N_5011);
and U5429 (N_5429,N_5125,N_5130);
xnor U5430 (N_5430,N_5168,N_5046);
and U5431 (N_5431,N_5023,N_5206);
or U5432 (N_5432,N_5094,N_5229);
and U5433 (N_5433,N_5074,N_5055);
or U5434 (N_5434,N_5146,N_5065);
nand U5435 (N_5435,N_5212,N_5232);
nor U5436 (N_5436,N_5191,N_5173);
and U5437 (N_5437,N_5121,N_5241);
nor U5438 (N_5438,N_5226,N_5149);
or U5439 (N_5439,N_5001,N_5242);
nor U5440 (N_5440,N_5180,N_5162);
and U5441 (N_5441,N_5195,N_5033);
xnor U5442 (N_5442,N_5083,N_5226);
nor U5443 (N_5443,N_5151,N_5044);
xor U5444 (N_5444,N_5183,N_5065);
or U5445 (N_5445,N_5079,N_5066);
or U5446 (N_5446,N_5107,N_5198);
nor U5447 (N_5447,N_5082,N_5210);
and U5448 (N_5448,N_5051,N_5241);
xnor U5449 (N_5449,N_5094,N_5002);
xnor U5450 (N_5450,N_5200,N_5190);
or U5451 (N_5451,N_5039,N_5125);
xnor U5452 (N_5452,N_5164,N_5027);
xor U5453 (N_5453,N_5062,N_5159);
or U5454 (N_5454,N_5014,N_5204);
nor U5455 (N_5455,N_5052,N_5222);
xor U5456 (N_5456,N_5200,N_5036);
or U5457 (N_5457,N_5065,N_5040);
xnor U5458 (N_5458,N_5082,N_5120);
nand U5459 (N_5459,N_5214,N_5181);
nor U5460 (N_5460,N_5043,N_5006);
nor U5461 (N_5461,N_5167,N_5140);
and U5462 (N_5462,N_5221,N_5228);
and U5463 (N_5463,N_5070,N_5221);
or U5464 (N_5464,N_5143,N_5137);
or U5465 (N_5465,N_5028,N_5033);
nor U5466 (N_5466,N_5122,N_5093);
nor U5467 (N_5467,N_5094,N_5195);
nand U5468 (N_5468,N_5230,N_5092);
and U5469 (N_5469,N_5029,N_5070);
and U5470 (N_5470,N_5196,N_5099);
and U5471 (N_5471,N_5074,N_5191);
and U5472 (N_5472,N_5210,N_5010);
and U5473 (N_5473,N_5245,N_5132);
and U5474 (N_5474,N_5123,N_5189);
xnor U5475 (N_5475,N_5046,N_5120);
nand U5476 (N_5476,N_5049,N_5105);
xnor U5477 (N_5477,N_5042,N_5233);
nor U5478 (N_5478,N_5249,N_5202);
and U5479 (N_5479,N_5127,N_5068);
and U5480 (N_5480,N_5020,N_5218);
or U5481 (N_5481,N_5079,N_5228);
and U5482 (N_5482,N_5126,N_5188);
or U5483 (N_5483,N_5144,N_5036);
and U5484 (N_5484,N_5140,N_5135);
or U5485 (N_5485,N_5026,N_5054);
or U5486 (N_5486,N_5047,N_5131);
and U5487 (N_5487,N_5231,N_5066);
xnor U5488 (N_5488,N_5230,N_5021);
xnor U5489 (N_5489,N_5180,N_5219);
and U5490 (N_5490,N_5233,N_5000);
or U5491 (N_5491,N_5015,N_5002);
or U5492 (N_5492,N_5158,N_5028);
and U5493 (N_5493,N_5139,N_5007);
nor U5494 (N_5494,N_5150,N_5196);
nand U5495 (N_5495,N_5135,N_5008);
or U5496 (N_5496,N_5012,N_5126);
or U5497 (N_5497,N_5089,N_5037);
nand U5498 (N_5498,N_5123,N_5032);
and U5499 (N_5499,N_5242,N_5248);
nand U5500 (N_5500,N_5370,N_5495);
xnor U5501 (N_5501,N_5444,N_5350);
nand U5502 (N_5502,N_5428,N_5386);
nand U5503 (N_5503,N_5306,N_5315);
nor U5504 (N_5504,N_5299,N_5333);
nand U5505 (N_5505,N_5390,N_5295);
and U5506 (N_5506,N_5323,N_5363);
or U5507 (N_5507,N_5381,N_5309);
or U5508 (N_5508,N_5492,N_5282);
nand U5509 (N_5509,N_5341,N_5255);
xnor U5510 (N_5510,N_5259,N_5313);
and U5511 (N_5511,N_5317,N_5278);
nor U5512 (N_5512,N_5280,N_5451);
nor U5513 (N_5513,N_5485,N_5483);
nor U5514 (N_5514,N_5368,N_5472);
nor U5515 (N_5515,N_5369,N_5404);
xor U5516 (N_5516,N_5437,N_5332);
xnor U5517 (N_5517,N_5427,N_5430);
nand U5518 (N_5518,N_5499,N_5277);
xnor U5519 (N_5519,N_5486,N_5318);
and U5520 (N_5520,N_5345,N_5416);
or U5521 (N_5521,N_5392,N_5407);
nor U5522 (N_5522,N_5302,N_5300);
xor U5523 (N_5523,N_5424,N_5384);
nand U5524 (N_5524,N_5325,N_5462);
and U5525 (N_5525,N_5425,N_5401);
nor U5526 (N_5526,N_5391,N_5445);
nor U5527 (N_5527,N_5402,N_5376);
xor U5528 (N_5528,N_5324,N_5264);
or U5529 (N_5529,N_5423,N_5467);
xor U5530 (N_5530,N_5343,N_5403);
or U5531 (N_5531,N_5422,N_5463);
nand U5532 (N_5532,N_5491,N_5454);
xnor U5533 (N_5533,N_5353,N_5498);
nand U5534 (N_5534,N_5272,N_5305);
xnor U5535 (N_5535,N_5421,N_5253);
and U5536 (N_5536,N_5352,N_5387);
nor U5537 (N_5537,N_5357,N_5434);
and U5538 (N_5538,N_5348,N_5304);
xnor U5539 (N_5539,N_5456,N_5452);
or U5540 (N_5540,N_5419,N_5408);
nand U5541 (N_5541,N_5261,N_5412);
and U5542 (N_5542,N_5360,N_5258);
xor U5543 (N_5543,N_5479,N_5399);
xor U5544 (N_5544,N_5470,N_5426);
and U5545 (N_5545,N_5312,N_5383);
xor U5546 (N_5546,N_5334,N_5335);
or U5547 (N_5547,N_5320,N_5385);
nor U5548 (N_5548,N_5373,N_5254);
nor U5549 (N_5549,N_5337,N_5339);
or U5550 (N_5550,N_5417,N_5297);
or U5551 (N_5551,N_5367,N_5276);
xor U5552 (N_5552,N_5414,N_5303);
and U5553 (N_5553,N_5466,N_5393);
or U5554 (N_5554,N_5371,N_5374);
or U5555 (N_5555,N_5398,N_5265);
nor U5556 (N_5556,N_5490,N_5395);
and U5557 (N_5557,N_5308,N_5286);
nor U5558 (N_5558,N_5497,N_5394);
and U5559 (N_5559,N_5442,N_5257);
xor U5560 (N_5560,N_5358,N_5418);
and U5561 (N_5561,N_5436,N_5478);
nor U5562 (N_5562,N_5330,N_5275);
or U5563 (N_5563,N_5397,N_5327);
or U5564 (N_5564,N_5291,N_5459);
or U5565 (N_5565,N_5406,N_5362);
and U5566 (N_5566,N_5443,N_5326);
nand U5567 (N_5567,N_5356,N_5439);
and U5568 (N_5568,N_5410,N_5477);
xor U5569 (N_5569,N_5482,N_5450);
and U5570 (N_5570,N_5471,N_5484);
nor U5571 (N_5571,N_5344,N_5328);
nor U5572 (N_5572,N_5266,N_5473);
xor U5573 (N_5573,N_5365,N_5378);
or U5574 (N_5574,N_5413,N_5380);
xor U5575 (N_5575,N_5449,N_5488);
and U5576 (N_5576,N_5331,N_5429);
xor U5577 (N_5577,N_5440,N_5489);
xor U5578 (N_5578,N_5438,N_5447);
nand U5579 (N_5579,N_5342,N_5441);
or U5580 (N_5580,N_5396,N_5354);
or U5581 (N_5581,N_5355,N_5340);
nand U5582 (N_5582,N_5329,N_5379);
or U5583 (N_5583,N_5420,N_5336);
or U5584 (N_5584,N_5260,N_5349);
or U5585 (N_5585,N_5267,N_5446);
nand U5586 (N_5586,N_5263,N_5366);
or U5587 (N_5587,N_5296,N_5415);
nor U5588 (N_5588,N_5274,N_5475);
nand U5589 (N_5589,N_5314,N_5359);
xor U5590 (N_5590,N_5476,N_5310);
xor U5591 (N_5591,N_5262,N_5270);
or U5592 (N_5592,N_5411,N_5465);
or U5593 (N_5593,N_5292,N_5298);
and U5594 (N_5594,N_5287,N_5283);
nor U5595 (N_5595,N_5400,N_5448);
or U5596 (N_5596,N_5351,N_5435);
nor U5597 (N_5597,N_5377,N_5432);
nor U5598 (N_5598,N_5468,N_5284);
nor U5599 (N_5599,N_5474,N_5301);
nand U5600 (N_5600,N_5285,N_5372);
xor U5601 (N_5601,N_5290,N_5480);
nor U5602 (N_5602,N_5455,N_5347);
and U5603 (N_5603,N_5458,N_5322);
nand U5604 (N_5604,N_5268,N_5273);
nor U5605 (N_5605,N_5289,N_5389);
and U5606 (N_5606,N_5271,N_5294);
nor U5607 (N_5607,N_5279,N_5251);
nand U5608 (N_5608,N_5361,N_5321);
xnor U5609 (N_5609,N_5364,N_5388);
xor U5610 (N_5610,N_5288,N_5311);
and U5611 (N_5611,N_5461,N_5405);
nor U5612 (N_5612,N_5469,N_5453);
nor U5613 (N_5613,N_5409,N_5457);
or U5614 (N_5614,N_5496,N_5494);
and U5615 (N_5615,N_5487,N_5319);
and U5616 (N_5616,N_5256,N_5338);
nor U5617 (N_5617,N_5464,N_5481);
and U5618 (N_5618,N_5281,N_5431);
nand U5619 (N_5619,N_5375,N_5382);
or U5620 (N_5620,N_5307,N_5433);
and U5621 (N_5621,N_5250,N_5316);
and U5622 (N_5622,N_5346,N_5493);
and U5623 (N_5623,N_5252,N_5460);
nor U5624 (N_5624,N_5269,N_5293);
and U5625 (N_5625,N_5263,N_5295);
or U5626 (N_5626,N_5354,N_5303);
and U5627 (N_5627,N_5252,N_5270);
and U5628 (N_5628,N_5379,N_5312);
xor U5629 (N_5629,N_5452,N_5378);
or U5630 (N_5630,N_5471,N_5499);
nand U5631 (N_5631,N_5492,N_5496);
nand U5632 (N_5632,N_5442,N_5253);
and U5633 (N_5633,N_5462,N_5302);
or U5634 (N_5634,N_5475,N_5438);
xor U5635 (N_5635,N_5292,N_5431);
and U5636 (N_5636,N_5413,N_5303);
xnor U5637 (N_5637,N_5391,N_5488);
nor U5638 (N_5638,N_5381,N_5279);
xor U5639 (N_5639,N_5292,N_5464);
nor U5640 (N_5640,N_5308,N_5413);
and U5641 (N_5641,N_5322,N_5488);
xnor U5642 (N_5642,N_5291,N_5303);
xor U5643 (N_5643,N_5346,N_5315);
nor U5644 (N_5644,N_5303,N_5310);
nand U5645 (N_5645,N_5360,N_5408);
nor U5646 (N_5646,N_5276,N_5460);
and U5647 (N_5647,N_5253,N_5487);
or U5648 (N_5648,N_5265,N_5358);
nor U5649 (N_5649,N_5479,N_5289);
nand U5650 (N_5650,N_5305,N_5496);
nand U5651 (N_5651,N_5304,N_5372);
nor U5652 (N_5652,N_5404,N_5343);
nand U5653 (N_5653,N_5358,N_5258);
or U5654 (N_5654,N_5324,N_5357);
nor U5655 (N_5655,N_5296,N_5364);
or U5656 (N_5656,N_5466,N_5310);
nor U5657 (N_5657,N_5380,N_5373);
or U5658 (N_5658,N_5455,N_5471);
nor U5659 (N_5659,N_5343,N_5327);
and U5660 (N_5660,N_5430,N_5332);
or U5661 (N_5661,N_5348,N_5390);
nand U5662 (N_5662,N_5466,N_5304);
or U5663 (N_5663,N_5445,N_5333);
or U5664 (N_5664,N_5414,N_5307);
nor U5665 (N_5665,N_5436,N_5266);
nand U5666 (N_5666,N_5467,N_5262);
and U5667 (N_5667,N_5471,N_5385);
or U5668 (N_5668,N_5294,N_5410);
and U5669 (N_5669,N_5292,N_5289);
or U5670 (N_5670,N_5467,N_5301);
and U5671 (N_5671,N_5494,N_5488);
or U5672 (N_5672,N_5379,N_5377);
xnor U5673 (N_5673,N_5464,N_5465);
nand U5674 (N_5674,N_5328,N_5406);
or U5675 (N_5675,N_5318,N_5302);
nor U5676 (N_5676,N_5459,N_5420);
xnor U5677 (N_5677,N_5356,N_5486);
xnor U5678 (N_5678,N_5324,N_5393);
xnor U5679 (N_5679,N_5309,N_5448);
nor U5680 (N_5680,N_5441,N_5403);
nand U5681 (N_5681,N_5253,N_5469);
or U5682 (N_5682,N_5455,N_5403);
and U5683 (N_5683,N_5426,N_5254);
or U5684 (N_5684,N_5263,N_5461);
nor U5685 (N_5685,N_5375,N_5486);
nor U5686 (N_5686,N_5461,N_5335);
nor U5687 (N_5687,N_5354,N_5380);
and U5688 (N_5688,N_5448,N_5494);
and U5689 (N_5689,N_5399,N_5328);
or U5690 (N_5690,N_5270,N_5369);
xnor U5691 (N_5691,N_5250,N_5390);
nand U5692 (N_5692,N_5410,N_5443);
nand U5693 (N_5693,N_5300,N_5429);
or U5694 (N_5694,N_5266,N_5345);
nor U5695 (N_5695,N_5262,N_5351);
nand U5696 (N_5696,N_5291,N_5412);
and U5697 (N_5697,N_5455,N_5342);
or U5698 (N_5698,N_5357,N_5360);
and U5699 (N_5699,N_5283,N_5436);
nor U5700 (N_5700,N_5395,N_5480);
nor U5701 (N_5701,N_5354,N_5479);
xor U5702 (N_5702,N_5348,N_5424);
xnor U5703 (N_5703,N_5257,N_5400);
xor U5704 (N_5704,N_5374,N_5345);
nor U5705 (N_5705,N_5391,N_5307);
nor U5706 (N_5706,N_5261,N_5313);
and U5707 (N_5707,N_5495,N_5343);
and U5708 (N_5708,N_5261,N_5498);
or U5709 (N_5709,N_5272,N_5395);
nor U5710 (N_5710,N_5256,N_5327);
or U5711 (N_5711,N_5414,N_5482);
or U5712 (N_5712,N_5357,N_5368);
or U5713 (N_5713,N_5442,N_5401);
xnor U5714 (N_5714,N_5256,N_5373);
nor U5715 (N_5715,N_5377,N_5406);
nor U5716 (N_5716,N_5425,N_5456);
and U5717 (N_5717,N_5283,N_5310);
xnor U5718 (N_5718,N_5320,N_5457);
and U5719 (N_5719,N_5354,N_5299);
xnor U5720 (N_5720,N_5368,N_5351);
xor U5721 (N_5721,N_5379,N_5494);
and U5722 (N_5722,N_5386,N_5492);
nand U5723 (N_5723,N_5442,N_5416);
nor U5724 (N_5724,N_5436,N_5298);
nand U5725 (N_5725,N_5324,N_5346);
and U5726 (N_5726,N_5407,N_5397);
nand U5727 (N_5727,N_5453,N_5364);
nand U5728 (N_5728,N_5494,N_5311);
nand U5729 (N_5729,N_5373,N_5363);
nand U5730 (N_5730,N_5499,N_5397);
and U5731 (N_5731,N_5385,N_5313);
xor U5732 (N_5732,N_5478,N_5325);
nor U5733 (N_5733,N_5452,N_5477);
xnor U5734 (N_5734,N_5340,N_5339);
nor U5735 (N_5735,N_5433,N_5265);
nor U5736 (N_5736,N_5342,N_5336);
nor U5737 (N_5737,N_5335,N_5419);
and U5738 (N_5738,N_5434,N_5451);
nand U5739 (N_5739,N_5496,N_5432);
nor U5740 (N_5740,N_5284,N_5452);
xor U5741 (N_5741,N_5283,N_5323);
nand U5742 (N_5742,N_5250,N_5347);
and U5743 (N_5743,N_5455,N_5363);
xnor U5744 (N_5744,N_5409,N_5459);
nor U5745 (N_5745,N_5388,N_5288);
or U5746 (N_5746,N_5486,N_5497);
xnor U5747 (N_5747,N_5298,N_5422);
nor U5748 (N_5748,N_5465,N_5468);
or U5749 (N_5749,N_5447,N_5374);
nor U5750 (N_5750,N_5701,N_5714);
nor U5751 (N_5751,N_5508,N_5741);
xnor U5752 (N_5752,N_5626,N_5562);
or U5753 (N_5753,N_5623,N_5549);
and U5754 (N_5754,N_5646,N_5579);
xor U5755 (N_5755,N_5734,N_5721);
nor U5756 (N_5756,N_5689,N_5572);
nand U5757 (N_5757,N_5633,N_5516);
nor U5758 (N_5758,N_5592,N_5690);
xor U5759 (N_5759,N_5695,N_5618);
or U5760 (N_5760,N_5547,N_5660);
xor U5761 (N_5761,N_5621,N_5539);
or U5762 (N_5762,N_5566,N_5733);
and U5763 (N_5763,N_5569,N_5712);
xor U5764 (N_5764,N_5598,N_5573);
or U5765 (N_5765,N_5532,N_5672);
and U5766 (N_5766,N_5608,N_5629);
nor U5767 (N_5767,N_5518,N_5698);
xor U5768 (N_5768,N_5713,N_5552);
xor U5769 (N_5769,N_5700,N_5590);
xnor U5770 (N_5770,N_5649,N_5648);
or U5771 (N_5771,N_5591,N_5513);
nor U5772 (N_5772,N_5725,N_5595);
and U5773 (N_5773,N_5600,N_5686);
or U5774 (N_5774,N_5528,N_5517);
nand U5775 (N_5775,N_5571,N_5650);
nor U5776 (N_5776,N_5682,N_5670);
or U5777 (N_5777,N_5638,N_5577);
and U5778 (N_5778,N_5745,N_5548);
or U5779 (N_5779,N_5643,N_5617);
nand U5780 (N_5780,N_5716,N_5519);
or U5781 (N_5781,N_5564,N_5653);
nand U5782 (N_5782,N_5535,N_5722);
nor U5783 (N_5783,N_5503,N_5647);
nand U5784 (N_5784,N_5523,N_5550);
xnor U5785 (N_5785,N_5597,N_5639);
nand U5786 (N_5786,N_5560,N_5706);
nand U5787 (N_5787,N_5537,N_5509);
and U5788 (N_5788,N_5681,N_5510);
xnor U5789 (N_5789,N_5616,N_5624);
and U5790 (N_5790,N_5568,N_5585);
nor U5791 (N_5791,N_5628,N_5589);
xnor U5792 (N_5792,N_5651,N_5538);
nor U5793 (N_5793,N_5738,N_5609);
nand U5794 (N_5794,N_5731,N_5630);
and U5795 (N_5795,N_5520,N_5501);
nand U5796 (N_5796,N_5744,N_5669);
and U5797 (N_5797,N_5603,N_5557);
and U5798 (N_5798,N_5574,N_5614);
or U5799 (N_5799,N_5511,N_5704);
and U5800 (N_5800,N_5615,N_5656);
nand U5801 (N_5801,N_5556,N_5610);
and U5802 (N_5802,N_5663,N_5596);
and U5803 (N_5803,N_5746,N_5551);
nor U5804 (N_5804,N_5534,N_5594);
or U5805 (N_5805,N_5540,N_5505);
and U5806 (N_5806,N_5729,N_5662);
nor U5807 (N_5807,N_5743,N_5652);
and U5808 (N_5808,N_5545,N_5696);
xor U5809 (N_5809,N_5593,N_5588);
or U5810 (N_5810,N_5697,N_5730);
nor U5811 (N_5811,N_5739,N_5708);
xor U5812 (N_5812,N_5536,N_5687);
nand U5813 (N_5813,N_5674,N_5507);
nand U5814 (N_5814,N_5654,N_5680);
nor U5815 (N_5815,N_5586,N_5567);
nor U5816 (N_5816,N_5737,N_5602);
xnor U5817 (N_5817,N_5673,N_5635);
and U5818 (N_5818,N_5620,N_5742);
or U5819 (N_5819,N_5658,N_5748);
nor U5820 (N_5820,N_5522,N_5699);
or U5821 (N_5821,N_5605,N_5718);
or U5822 (N_5822,N_5740,N_5559);
xnor U5823 (N_5823,N_5606,N_5504);
xnor U5824 (N_5824,N_5724,N_5715);
and U5825 (N_5825,N_5612,N_5703);
and U5826 (N_5826,N_5688,N_5521);
and U5827 (N_5827,N_5717,N_5720);
or U5828 (N_5828,N_5529,N_5645);
nor U5829 (N_5829,N_5531,N_5702);
or U5830 (N_5830,N_5710,N_5691);
xnor U5831 (N_5831,N_5644,N_5580);
nand U5832 (N_5832,N_5683,N_5506);
nand U5833 (N_5833,N_5627,N_5541);
xor U5834 (N_5834,N_5530,N_5533);
xor U5835 (N_5835,N_5705,N_5728);
nor U5836 (N_5836,N_5640,N_5524);
or U5837 (N_5837,N_5694,N_5671);
xor U5838 (N_5838,N_5634,N_5607);
or U5839 (N_5839,N_5665,N_5668);
and U5840 (N_5840,N_5719,N_5676);
and U5841 (N_5841,N_5514,N_5526);
xor U5842 (N_5842,N_5723,N_5625);
nor U5843 (N_5843,N_5684,N_5692);
or U5844 (N_5844,N_5636,N_5619);
or U5845 (N_5845,N_5711,N_5677);
nor U5846 (N_5846,N_5563,N_5576);
nand U5847 (N_5847,N_5747,N_5575);
and U5848 (N_5848,N_5502,N_5611);
nand U5849 (N_5849,N_5655,N_5749);
xnor U5850 (N_5850,N_5546,N_5599);
xnor U5851 (N_5851,N_5527,N_5561);
and U5852 (N_5852,N_5587,N_5500);
xnor U5853 (N_5853,N_5637,N_5582);
and U5854 (N_5854,N_5641,N_5707);
nand U5855 (N_5855,N_5657,N_5736);
and U5856 (N_5856,N_5679,N_5555);
or U5857 (N_5857,N_5632,N_5675);
xor U5858 (N_5858,N_5583,N_5578);
or U5859 (N_5859,N_5678,N_5565);
or U5860 (N_5860,N_5515,N_5581);
and U5861 (N_5861,N_5554,N_5659);
nor U5862 (N_5862,N_5553,N_5570);
xor U5863 (N_5863,N_5558,N_5664);
xnor U5864 (N_5864,N_5726,N_5693);
xor U5865 (N_5865,N_5666,N_5525);
nor U5866 (N_5866,N_5542,N_5642);
or U5867 (N_5867,N_5709,N_5601);
or U5868 (N_5868,N_5727,N_5543);
xor U5869 (N_5869,N_5512,N_5544);
xnor U5870 (N_5870,N_5622,N_5613);
nand U5871 (N_5871,N_5685,N_5661);
xnor U5872 (N_5872,N_5735,N_5584);
nor U5873 (N_5873,N_5732,N_5631);
nor U5874 (N_5874,N_5667,N_5604);
nand U5875 (N_5875,N_5506,N_5615);
nand U5876 (N_5876,N_5681,N_5684);
nor U5877 (N_5877,N_5671,N_5532);
nand U5878 (N_5878,N_5647,N_5592);
nor U5879 (N_5879,N_5624,N_5561);
and U5880 (N_5880,N_5546,N_5664);
nand U5881 (N_5881,N_5581,N_5593);
nand U5882 (N_5882,N_5655,N_5593);
and U5883 (N_5883,N_5515,N_5502);
nor U5884 (N_5884,N_5574,N_5591);
nor U5885 (N_5885,N_5637,N_5602);
or U5886 (N_5886,N_5551,N_5661);
nand U5887 (N_5887,N_5719,N_5697);
nor U5888 (N_5888,N_5705,N_5625);
nand U5889 (N_5889,N_5528,N_5621);
or U5890 (N_5890,N_5539,N_5716);
or U5891 (N_5891,N_5744,N_5665);
nor U5892 (N_5892,N_5714,N_5684);
nor U5893 (N_5893,N_5507,N_5732);
and U5894 (N_5894,N_5662,N_5556);
nor U5895 (N_5895,N_5532,N_5571);
and U5896 (N_5896,N_5611,N_5707);
xnor U5897 (N_5897,N_5718,N_5545);
or U5898 (N_5898,N_5557,N_5577);
and U5899 (N_5899,N_5567,N_5712);
and U5900 (N_5900,N_5699,N_5605);
or U5901 (N_5901,N_5678,N_5692);
and U5902 (N_5902,N_5574,N_5650);
nor U5903 (N_5903,N_5564,N_5659);
xnor U5904 (N_5904,N_5561,N_5525);
nor U5905 (N_5905,N_5530,N_5707);
or U5906 (N_5906,N_5510,N_5685);
xnor U5907 (N_5907,N_5529,N_5670);
xnor U5908 (N_5908,N_5540,N_5571);
xor U5909 (N_5909,N_5564,N_5707);
nor U5910 (N_5910,N_5500,N_5689);
xor U5911 (N_5911,N_5530,N_5681);
or U5912 (N_5912,N_5540,N_5555);
and U5913 (N_5913,N_5638,N_5743);
xnor U5914 (N_5914,N_5691,N_5527);
nand U5915 (N_5915,N_5639,N_5586);
or U5916 (N_5916,N_5684,N_5532);
nand U5917 (N_5917,N_5690,N_5579);
or U5918 (N_5918,N_5728,N_5721);
nand U5919 (N_5919,N_5646,N_5621);
or U5920 (N_5920,N_5701,N_5619);
and U5921 (N_5921,N_5505,N_5680);
nand U5922 (N_5922,N_5664,N_5713);
xnor U5923 (N_5923,N_5543,N_5571);
or U5924 (N_5924,N_5526,N_5592);
or U5925 (N_5925,N_5675,N_5644);
and U5926 (N_5926,N_5505,N_5639);
xnor U5927 (N_5927,N_5727,N_5514);
and U5928 (N_5928,N_5653,N_5643);
nand U5929 (N_5929,N_5701,N_5657);
nor U5930 (N_5930,N_5579,N_5561);
nand U5931 (N_5931,N_5532,N_5633);
xor U5932 (N_5932,N_5629,N_5638);
nor U5933 (N_5933,N_5513,N_5576);
nand U5934 (N_5934,N_5547,N_5575);
xor U5935 (N_5935,N_5596,N_5579);
or U5936 (N_5936,N_5677,N_5628);
or U5937 (N_5937,N_5620,N_5663);
and U5938 (N_5938,N_5532,N_5600);
nand U5939 (N_5939,N_5581,N_5510);
nor U5940 (N_5940,N_5509,N_5628);
nand U5941 (N_5941,N_5615,N_5735);
and U5942 (N_5942,N_5689,N_5654);
and U5943 (N_5943,N_5737,N_5688);
or U5944 (N_5944,N_5606,N_5528);
or U5945 (N_5945,N_5689,N_5631);
nor U5946 (N_5946,N_5589,N_5733);
or U5947 (N_5947,N_5584,N_5621);
nor U5948 (N_5948,N_5562,N_5731);
or U5949 (N_5949,N_5503,N_5520);
and U5950 (N_5950,N_5686,N_5593);
nand U5951 (N_5951,N_5551,N_5575);
and U5952 (N_5952,N_5738,N_5564);
nand U5953 (N_5953,N_5733,N_5666);
xor U5954 (N_5954,N_5589,N_5632);
nor U5955 (N_5955,N_5685,N_5684);
nand U5956 (N_5956,N_5537,N_5576);
nor U5957 (N_5957,N_5696,N_5706);
xnor U5958 (N_5958,N_5644,N_5550);
nor U5959 (N_5959,N_5637,N_5691);
nor U5960 (N_5960,N_5539,N_5737);
nor U5961 (N_5961,N_5606,N_5715);
or U5962 (N_5962,N_5724,N_5603);
and U5963 (N_5963,N_5567,N_5664);
xor U5964 (N_5964,N_5546,N_5563);
nor U5965 (N_5965,N_5650,N_5500);
nor U5966 (N_5966,N_5584,N_5656);
nor U5967 (N_5967,N_5543,N_5518);
xor U5968 (N_5968,N_5564,N_5740);
nand U5969 (N_5969,N_5611,N_5554);
or U5970 (N_5970,N_5558,N_5542);
xnor U5971 (N_5971,N_5725,N_5593);
or U5972 (N_5972,N_5632,N_5594);
and U5973 (N_5973,N_5740,N_5606);
xor U5974 (N_5974,N_5699,N_5653);
xnor U5975 (N_5975,N_5620,N_5599);
and U5976 (N_5976,N_5538,N_5613);
nor U5977 (N_5977,N_5542,N_5721);
and U5978 (N_5978,N_5704,N_5669);
nor U5979 (N_5979,N_5722,N_5613);
xnor U5980 (N_5980,N_5644,N_5693);
or U5981 (N_5981,N_5687,N_5691);
and U5982 (N_5982,N_5720,N_5638);
and U5983 (N_5983,N_5595,N_5703);
or U5984 (N_5984,N_5592,N_5666);
or U5985 (N_5985,N_5552,N_5515);
nand U5986 (N_5986,N_5642,N_5555);
xnor U5987 (N_5987,N_5619,N_5608);
xor U5988 (N_5988,N_5680,N_5705);
and U5989 (N_5989,N_5636,N_5685);
nand U5990 (N_5990,N_5564,N_5579);
and U5991 (N_5991,N_5536,N_5637);
xor U5992 (N_5992,N_5534,N_5616);
nor U5993 (N_5993,N_5679,N_5614);
nor U5994 (N_5994,N_5683,N_5660);
or U5995 (N_5995,N_5711,N_5568);
nand U5996 (N_5996,N_5646,N_5602);
and U5997 (N_5997,N_5580,N_5625);
nor U5998 (N_5998,N_5575,N_5634);
and U5999 (N_5999,N_5594,N_5667);
xor U6000 (N_6000,N_5787,N_5859);
or U6001 (N_6001,N_5751,N_5888);
nor U6002 (N_6002,N_5912,N_5898);
xor U6003 (N_6003,N_5798,N_5869);
and U6004 (N_6004,N_5939,N_5764);
and U6005 (N_6005,N_5935,N_5796);
nor U6006 (N_6006,N_5802,N_5767);
or U6007 (N_6007,N_5877,N_5933);
xor U6008 (N_6008,N_5913,N_5766);
and U6009 (N_6009,N_5980,N_5856);
and U6010 (N_6010,N_5792,N_5806);
xor U6011 (N_6011,N_5837,N_5942);
nor U6012 (N_6012,N_5899,N_5931);
and U6013 (N_6013,N_5985,N_5968);
nand U6014 (N_6014,N_5927,N_5814);
nand U6015 (N_6015,N_5872,N_5768);
or U6016 (N_6016,N_5844,N_5848);
and U6017 (N_6017,N_5956,N_5760);
or U6018 (N_6018,N_5833,N_5772);
xor U6019 (N_6019,N_5762,N_5831);
nor U6020 (N_6020,N_5753,N_5780);
or U6021 (N_6021,N_5979,N_5897);
xor U6022 (N_6022,N_5785,N_5917);
or U6023 (N_6023,N_5819,N_5828);
xnor U6024 (N_6024,N_5786,N_5907);
nand U6025 (N_6025,N_5902,N_5884);
or U6026 (N_6026,N_5915,N_5955);
or U6027 (N_6027,N_5822,N_5783);
or U6028 (N_6028,N_5776,N_5769);
nand U6029 (N_6029,N_5824,N_5826);
nor U6030 (N_6030,N_5839,N_5977);
or U6031 (N_6031,N_5845,N_5949);
nand U6032 (N_6032,N_5849,N_5975);
xnor U6033 (N_6033,N_5882,N_5952);
xnor U6034 (N_6034,N_5922,N_5960);
nor U6035 (N_6035,N_5934,N_5823);
nor U6036 (N_6036,N_5862,N_5843);
or U6037 (N_6037,N_5857,N_5782);
or U6038 (N_6038,N_5873,N_5870);
xor U6039 (N_6039,N_5801,N_5860);
nand U6040 (N_6040,N_5797,N_5793);
and U6041 (N_6041,N_5761,N_5815);
nand U6042 (N_6042,N_5970,N_5791);
and U6043 (N_6043,N_5863,N_5887);
or U6044 (N_6044,N_5832,N_5983);
nand U6045 (N_6045,N_5986,N_5976);
nand U6046 (N_6046,N_5842,N_5966);
xnor U6047 (N_6047,N_5808,N_5900);
nor U6048 (N_6048,N_5962,N_5805);
nand U6049 (N_6049,N_5908,N_5892);
xnor U6050 (N_6050,N_5759,N_5840);
and U6051 (N_6051,N_5846,N_5940);
and U6052 (N_6052,N_5971,N_5829);
and U6053 (N_6053,N_5771,N_5795);
xor U6054 (N_6054,N_5896,N_5804);
xor U6055 (N_6055,N_5958,N_5957);
nand U6056 (N_6056,N_5923,N_5944);
or U6057 (N_6057,N_5946,N_5984);
and U6058 (N_6058,N_5918,N_5936);
nor U6059 (N_6059,N_5969,N_5964);
xor U6060 (N_6060,N_5868,N_5865);
and U6061 (N_6061,N_5929,N_5879);
nor U6062 (N_6062,N_5779,N_5991);
nand U6063 (N_6063,N_5997,N_5850);
nand U6064 (N_6064,N_5864,N_5853);
or U6065 (N_6065,N_5995,N_5827);
or U6066 (N_6066,N_5885,N_5799);
nor U6067 (N_6067,N_5999,N_5794);
and U6068 (N_6068,N_5881,N_5961);
and U6069 (N_6069,N_5932,N_5954);
and U6070 (N_6070,N_5750,N_5874);
nand U6071 (N_6071,N_5994,N_5996);
nand U6072 (N_6072,N_5998,N_5972);
nand U6073 (N_6073,N_5943,N_5758);
or U6074 (N_6074,N_5901,N_5851);
xnor U6075 (N_6075,N_5945,N_5880);
or U6076 (N_6076,N_5925,N_5889);
or U6077 (N_6077,N_5947,N_5965);
xor U6078 (N_6078,N_5921,N_5990);
nor U6079 (N_6079,N_5982,N_5973);
xnor U6080 (N_6080,N_5941,N_5810);
and U6081 (N_6081,N_5963,N_5992);
and U6082 (N_6082,N_5855,N_5930);
nand U6083 (N_6083,N_5773,N_5948);
xor U6084 (N_6084,N_5904,N_5763);
or U6085 (N_6085,N_5988,N_5770);
nand U6086 (N_6086,N_5838,N_5765);
xnor U6087 (N_6087,N_5950,N_5878);
xor U6088 (N_6088,N_5754,N_5895);
and U6089 (N_6089,N_5867,N_5928);
and U6090 (N_6090,N_5910,N_5938);
and U6091 (N_6091,N_5978,N_5911);
nand U6092 (N_6092,N_5919,N_5951);
and U6093 (N_6093,N_5886,N_5893);
and U6094 (N_6094,N_5852,N_5812);
nand U6095 (N_6095,N_5858,N_5784);
and U6096 (N_6096,N_5757,N_5752);
or U6097 (N_6097,N_5835,N_5816);
xnor U6098 (N_6098,N_5905,N_5774);
nand U6099 (N_6099,N_5789,N_5813);
xor U6100 (N_6100,N_5830,N_5926);
nand U6101 (N_6101,N_5967,N_5817);
and U6102 (N_6102,N_5974,N_5909);
xnor U6103 (N_6103,N_5890,N_5989);
and U6104 (N_6104,N_5836,N_5803);
and U6105 (N_6105,N_5788,N_5778);
or U6106 (N_6106,N_5820,N_5903);
or U6107 (N_6107,N_5937,N_5809);
nand U6108 (N_6108,N_5807,N_5854);
nand U6109 (N_6109,N_5818,N_5924);
xnor U6110 (N_6110,N_5914,N_5790);
or U6111 (N_6111,N_5821,N_5775);
or U6112 (N_6112,N_5993,N_5825);
nor U6113 (N_6113,N_5777,N_5953);
and U6114 (N_6114,N_5834,N_5866);
and U6115 (N_6115,N_5756,N_5906);
nand U6116 (N_6116,N_5959,N_5781);
nor U6117 (N_6117,N_5841,N_5987);
xor U6118 (N_6118,N_5916,N_5981);
and U6119 (N_6119,N_5811,N_5800);
nand U6120 (N_6120,N_5883,N_5920);
nand U6121 (N_6121,N_5861,N_5894);
nand U6122 (N_6122,N_5875,N_5891);
nand U6123 (N_6123,N_5755,N_5847);
xnor U6124 (N_6124,N_5876,N_5871);
xor U6125 (N_6125,N_5822,N_5929);
xor U6126 (N_6126,N_5975,N_5880);
xnor U6127 (N_6127,N_5935,N_5941);
or U6128 (N_6128,N_5851,N_5882);
nor U6129 (N_6129,N_5821,N_5985);
or U6130 (N_6130,N_5904,N_5794);
nor U6131 (N_6131,N_5989,N_5944);
nand U6132 (N_6132,N_5907,N_5802);
xor U6133 (N_6133,N_5850,N_5822);
or U6134 (N_6134,N_5764,N_5775);
xnor U6135 (N_6135,N_5910,N_5849);
nor U6136 (N_6136,N_5923,N_5930);
nand U6137 (N_6137,N_5947,N_5824);
nor U6138 (N_6138,N_5865,N_5862);
and U6139 (N_6139,N_5859,N_5929);
nand U6140 (N_6140,N_5981,N_5863);
and U6141 (N_6141,N_5940,N_5984);
nor U6142 (N_6142,N_5922,N_5967);
nand U6143 (N_6143,N_5819,N_5971);
and U6144 (N_6144,N_5959,N_5877);
and U6145 (N_6145,N_5946,N_5830);
and U6146 (N_6146,N_5793,N_5788);
nand U6147 (N_6147,N_5791,N_5951);
and U6148 (N_6148,N_5758,N_5898);
and U6149 (N_6149,N_5790,N_5861);
xor U6150 (N_6150,N_5933,N_5858);
xor U6151 (N_6151,N_5910,N_5777);
or U6152 (N_6152,N_5750,N_5969);
or U6153 (N_6153,N_5826,N_5937);
xnor U6154 (N_6154,N_5985,N_5756);
xor U6155 (N_6155,N_5969,N_5844);
nand U6156 (N_6156,N_5986,N_5988);
or U6157 (N_6157,N_5980,N_5897);
and U6158 (N_6158,N_5969,N_5975);
or U6159 (N_6159,N_5770,N_5866);
nand U6160 (N_6160,N_5761,N_5994);
nor U6161 (N_6161,N_5814,N_5865);
or U6162 (N_6162,N_5801,N_5909);
or U6163 (N_6163,N_5985,N_5788);
and U6164 (N_6164,N_5917,N_5816);
xor U6165 (N_6165,N_5787,N_5973);
xnor U6166 (N_6166,N_5768,N_5954);
or U6167 (N_6167,N_5963,N_5833);
or U6168 (N_6168,N_5795,N_5949);
nor U6169 (N_6169,N_5896,N_5930);
and U6170 (N_6170,N_5938,N_5757);
or U6171 (N_6171,N_5858,N_5889);
xor U6172 (N_6172,N_5824,N_5846);
and U6173 (N_6173,N_5985,N_5817);
nor U6174 (N_6174,N_5792,N_5987);
or U6175 (N_6175,N_5795,N_5845);
and U6176 (N_6176,N_5753,N_5928);
xnor U6177 (N_6177,N_5884,N_5821);
xor U6178 (N_6178,N_5908,N_5895);
xor U6179 (N_6179,N_5899,N_5837);
nor U6180 (N_6180,N_5989,N_5955);
nand U6181 (N_6181,N_5837,N_5804);
nand U6182 (N_6182,N_5924,N_5774);
nand U6183 (N_6183,N_5817,N_5933);
nor U6184 (N_6184,N_5939,N_5942);
nor U6185 (N_6185,N_5963,N_5849);
nor U6186 (N_6186,N_5873,N_5983);
nor U6187 (N_6187,N_5873,N_5820);
xnor U6188 (N_6188,N_5990,N_5841);
xor U6189 (N_6189,N_5831,N_5964);
nor U6190 (N_6190,N_5782,N_5935);
xor U6191 (N_6191,N_5797,N_5764);
and U6192 (N_6192,N_5872,N_5902);
nor U6193 (N_6193,N_5947,N_5792);
nand U6194 (N_6194,N_5776,N_5758);
or U6195 (N_6195,N_5840,N_5984);
and U6196 (N_6196,N_5750,N_5972);
nand U6197 (N_6197,N_5958,N_5760);
nand U6198 (N_6198,N_5758,N_5969);
and U6199 (N_6199,N_5756,N_5881);
xor U6200 (N_6200,N_5965,N_5945);
nor U6201 (N_6201,N_5884,N_5984);
nand U6202 (N_6202,N_5879,N_5761);
nand U6203 (N_6203,N_5984,N_5788);
xnor U6204 (N_6204,N_5979,N_5760);
nor U6205 (N_6205,N_5825,N_5892);
or U6206 (N_6206,N_5912,N_5807);
or U6207 (N_6207,N_5831,N_5882);
or U6208 (N_6208,N_5778,N_5800);
nand U6209 (N_6209,N_5920,N_5904);
nand U6210 (N_6210,N_5990,N_5802);
nor U6211 (N_6211,N_5782,N_5860);
nor U6212 (N_6212,N_5825,N_5866);
or U6213 (N_6213,N_5990,N_5900);
nor U6214 (N_6214,N_5812,N_5786);
and U6215 (N_6215,N_5877,N_5872);
and U6216 (N_6216,N_5844,N_5854);
nor U6217 (N_6217,N_5897,N_5907);
or U6218 (N_6218,N_5770,N_5966);
and U6219 (N_6219,N_5760,N_5917);
xor U6220 (N_6220,N_5846,N_5782);
nor U6221 (N_6221,N_5976,N_5794);
xnor U6222 (N_6222,N_5792,N_5932);
xnor U6223 (N_6223,N_5824,N_5981);
xor U6224 (N_6224,N_5910,N_5893);
nand U6225 (N_6225,N_5907,N_5976);
and U6226 (N_6226,N_5843,N_5931);
xnor U6227 (N_6227,N_5794,N_5817);
xor U6228 (N_6228,N_5854,N_5966);
nor U6229 (N_6229,N_5887,N_5862);
xnor U6230 (N_6230,N_5966,N_5887);
nand U6231 (N_6231,N_5809,N_5886);
nor U6232 (N_6232,N_5775,N_5938);
xnor U6233 (N_6233,N_5854,N_5838);
xor U6234 (N_6234,N_5918,N_5767);
xor U6235 (N_6235,N_5840,N_5751);
and U6236 (N_6236,N_5946,N_5959);
nor U6237 (N_6237,N_5986,N_5842);
and U6238 (N_6238,N_5845,N_5805);
xor U6239 (N_6239,N_5945,N_5997);
and U6240 (N_6240,N_5767,N_5964);
and U6241 (N_6241,N_5981,N_5886);
and U6242 (N_6242,N_5918,N_5852);
nor U6243 (N_6243,N_5855,N_5892);
and U6244 (N_6244,N_5984,N_5827);
nand U6245 (N_6245,N_5966,N_5858);
and U6246 (N_6246,N_5809,N_5790);
or U6247 (N_6247,N_5821,N_5861);
and U6248 (N_6248,N_5956,N_5989);
nor U6249 (N_6249,N_5871,N_5869);
or U6250 (N_6250,N_6232,N_6001);
nor U6251 (N_6251,N_6164,N_6078);
and U6252 (N_6252,N_6229,N_6211);
and U6253 (N_6253,N_6194,N_6234);
or U6254 (N_6254,N_6169,N_6070);
xnor U6255 (N_6255,N_6034,N_6107);
and U6256 (N_6256,N_6185,N_6133);
or U6257 (N_6257,N_6080,N_6228);
xnor U6258 (N_6258,N_6157,N_6042);
nand U6259 (N_6259,N_6204,N_6134);
nor U6260 (N_6260,N_6173,N_6071);
and U6261 (N_6261,N_6023,N_6247);
and U6262 (N_6262,N_6111,N_6047);
xnor U6263 (N_6263,N_6206,N_6153);
nor U6264 (N_6264,N_6017,N_6118);
or U6265 (N_6265,N_6127,N_6066);
xor U6266 (N_6266,N_6132,N_6113);
nor U6267 (N_6267,N_6021,N_6140);
nand U6268 (N_6268,N_6245,N_6033);
or U6269 (N_6269,N_6043,N_6156);
nor U6270 (N_6270,N_6090,N_6104);
and U6271 (N_6271,N_6068,N_6233);
or U6272 (N_6272,N_6181,N_6039);
nor U6273 (N_6273,N_6161,N_6190);
nand U6274 (N_6274,N_6005,N_6031);
and U6275 (N_6275,N_6099,N_6209);
or U6276 (N_6276,N_6026,N_6150);
and U6277 (N_6277,N_6231,N_6077);
and U6278 (N_6278,N_6027,N_6130);
nand U6279 (N_6279,N_6041,N_6085);
and U6280 (N_6280,N_6162,N_6167);
or U6281 (N_6281,N_6193,N_6028);
and U6282 (N_6282,N_6019,N_6146);
or U6283 (N_6283,N_6010,N_6094);
or U6284 (N_6284,N_6239,N_6105);
xnor U6285 (N_6285,N_6144,N_6050);
and U6286 (N_6286,N_6192,N_6121);
and U6287 (N_6287,N_6046,N_6060);
xor U6288 (N_6288,N_6037,N_6096);
and U6289 (N_6289,N_6213,N_6240);
nand U6290 (N_6290,N_6131,N_6171);
nor U6291 (N_6291,N_6015,N_6097);
and U6292 (N_6292,N_6135,N_6159);
or U6293 (N_6293,N_6053,N_6124);
and U6294 (N_6294,N_6238,N_6087);
or U6295 (N_6295,N_6125,N_6038);
nor U6296 (N_6296,N_6014,N_6226);
or U6297 (N_6297,N_6221,N_6115);
or U6298 (N_6298,N_6049,N_6222);
xor U6299 (N_6299,N_6016,N_6123);
and U6300 (N_6300,N_6064,N_6139);
xor U6301 (N_6301,N_6095,N_6142);
or U6302 (N_6302,N_6008,N_6235);
xor U6303 (N_6303,N_6110,N_6207);
and U6304 (N_6304,N_6191,N_6086);
nor U6305 (N_6305,N_6128,N_6061);
or U6306 (N_6306,N_6237,N_6227);
nand U6307 (N_6307,N_6083,N_6223);
and U6308 (N_6308,N_6022,N_6197);
nor U6309 (N_6309,N_6116,N_6184);
xnor U6310 (N_6310,N_6241,N_6152);
nor U6311 (N_6311,N_6199,N_6225);
xnor U6312 (N_6312,N_6036,N_6108);
or U6313 (N_6313,N_6189,N_6218);
and U6314 (N_6314,N_6178,N_6112);
nand U6315 (N_6315,N_6003,N_6212);
and U6316 (N_6316,N_6106,N_6126);
nand U6317 (N_6317,N_6081,N_6170);
or U6318 (N_6318,N_6119,N_6089);
nand U6319 (N_6319,N_6129,N_6004);
xnor U6320 (N_6320,N_6155,N_6200);
or U6321 (N_6321,N_6073,N_6098);
and U6322 (N_6322,N_6180,N_6137);
nand U6323 (N_6323,N_6002,N_6051);
or U6324 (N_6324,N_6101,N_6203);
nor U6325 (N_6325,N_6141,N_6214);
nand U6326 (N_6326,N_6122,N_6092);
or U6327 (N_6327,N_6114,N_6032);
or U6328 (N_6328,N_6143,N_6208);
nand U6329 (N_6329,N_6007,N_6147);
xnor U6330 (N_6330,N_6012,N_6198);
nor U6331 (N_6331,N_6058,N_6093);
or U6332 (N_6332,N_6160,N_6244);
or U6333 (N_6333,N_6102,N_6165);
xor U6334 (N_6334,N_6062,N_6236);
nor U6335 (N_6335,N_6056,N_6176);
or U6336 (N_6336,N_6136,N_6151);
nand U6337 (N_6337,N_6243,N_6168);
or U6338 (N_6338,N_6067,N_6020);
or U6339 (N_6339,N_6154,N_6182);
nand U6340 (N_6340,N_6069,N_6065);
nor U6341 (N_6341,N_6075,N_6220);
xnor U6342 (N_6342,N_6187,N_6100);
xor U6343 (N_6343,N_6201,N_6045);
or U6344 (N_6344,N_6084,N_6246);
xnor U6345 (N_6345,N_6048,N_6210);
xor U6346 (N_6346,N_6196,N_6163);
xor U6347 (N_6347,N_6242,N_6158);
and U6348 (N_6348,N_6009,N_6183);
nand U6349 (N_6349,N_6109,N_6074);
or U6350 (N_6350,N_6013,N_6088);
and U6351 (N_6351,N_6216,N_6052);
xor U6352 (N_6352,N_6215,N_6082);
xnor U6353 (N_6353,N_6006,N_6175);
or U6354 (N_6354,N_6195,N_6217);
nor U6355 (N_6355,N_6044,N_6179);
nor U6356 (N_6356,N_6076,N_6249);
xor U6357 (N_6357,N_6063,N_6000);
nand U6358 (N_6358,N_6024,N_6202);
xnor U6359 (N_6359,N_6138,N_6035);
nor U6360 (N_6360,N_6011,N_6172);
nor U6361 (N_6361,N_6230,N_6188);
and U6362 (N_6362,N_6145,N_6059);
xor U6363 (N_6363,N_6103,N_6030);
and U6364 (N_6364,N_6057,N_6040);
nand U6365 (N_6365,N_6018,N_6120);
xnor U6366 (N_6366,N_6054,N_6177);
xnor U6367 (N_6367,N_6148,N_6219);
and U6368 (N_6368,N_6174,N_6029);
or U6369 (N_6369,N_6025,N_6224);
xnor U6370 (N_6370,N_6149,N_6091);
xor U6371 (N_6371,N_6072,N_6055);
or U6372 (N_6372,N_6186,N_6166);
nor U6373 (N_6373,N_6117,N_6205);
nor U6374 (N_6374,N_6079,N_6248);
nand U6375 (N_6375,N_6075,N_6001);
nand U6376 (N_6376,N_6072,N_6243);
and U6377 (N_6377,N_6206,N_6146);
nand U6378 (N_6378,N_6055,N_6018);
nor U6379 (N_6379,N_6138,N_6036);
or U6380 (N_6380,N_6167,N_6064);
and U6381 (N_6381,N_6011,N_6222);
and U6382 (N_6382,N_6104,N_6209);
nor U6383 (N_6383,N_6220,N_6067);
nor U6384 (N_6384,N_6073,N_6081);
xor U6385 (N_6385,N_6249,N_6028);
nor U6386 (N_6386,N_6061,N_6219);
and U6387 (N_6387,N_6015,N_6131);
and U6388 (N_6388,N_6114,N_6102);
xor U6389 (N_6389,N_6076,N_6007);
nor U6390 (N_6390,N_6100,N_6139);
nand U6391 (N_6391,N_6048,N_6155);
nor U6392 (N_6392,N_6222,N_6155);
nand U6393 (N_6393,N_6021,N_6147);
xor U6394 (N_6394,N_6218,N_6035);
or U6395 (N_6395,N_6056,N_6184);
or U6396 (N_6396,N_6050,N_6207);
nand U6397 (N_6397,N_6201,N_6180);
or U6398 (N_6398,N_6052,N_6208);
xnor U6399 (N_6399,N_6044,N_6131);
or U6400 (N_6400,N_6102,N_6038);
xor U6401 (N_6401,N_6032,N_6028);
nor U6402 (N_6402,N_6028,N_6170);
nor U6403 (N_6403,N_6138,N_6068);
and U6404 (N_6404,N_6232,N_6059);
and U6405 (N_6405,N_6135,N_6025);
xnor U6406 (N_6406,N_6221,N_6131);
or U6407 (N_6407,N_6056,N_6134);
or U6408 (N_6408,N_6116,N_6047);
or U6409 (N_6409,N_6048,N_6194);
and U6410 (N_6410,N_6099,N_6117);
or U6411 (N_6411,N_6089,N_6028);
xor U6412 (N_6412,N_6230,N_6025);
nand U6413 (N_6413,N_6078,N_6112);
or U6414 (N_6414,N_6002,N_6034);
or U6415 (N_6415,N_6161,N_6164);
or U6416 (N_6416,N_6188,N_6141);
nand U6417 (N_6417,N_6179,N_6070);
or U6418 (N_6418,N_6215,N_6180);
xnor U6419 (N_6419,N_6203,N_6226);
nand U6420 (N_6420,N_6192,N_6104);
nand U6421 (N_6421,N_6038,N_6215);
xnor U6422 (N_6422,N_6073,N_6210);
or U6423 (N_6423,N_6004,N_6080);
and U6424 (N_6424,N_6201,N_6024);
nand U6425 (N_6425,N_6215,N_6187);
xor U6426 (N_6426,N_6092,N_6043);
and U6427 (N_6427,N_6055,N_6008);
nor U6428 (N_6428,N_6021,N_6245);
xor U6429 (N_6429,N_6022,N_6128);
or U6430 (N_6430,N_6231,N_6214);
nor U6431 (N_6431,N_6207,N_6246);
xnor U6432 (N_6432,N_6060,N_6130);
and U6433 (N_6433,N_6084,N_6030);
nor U6434 (N_6434,N_6127,N_6011);
xnor U6435 (N_6435,N_6108,N_6120);
or U6436 (N_6436,N_6012,N_6115);
nand U6437 (N_6437,N_6122,N_6191);
nand U6438 (N_6438,N_6064,N_6104);
and U6439 (N_6439,N_6234,N_6009);
nor U6440 (N_6440,N_6139,N_6056);
nor U6441 (N_6441,N_6155,N_6104);
and U6442 (N_6442,N_6000,N_6163);
or U6443 (N_6443,N_6050,N_6156);
nor U6444 (N_6444,N_6160,N_6149);
xnor U6445 (N_6445,N_6047,N_6126);
or U6446 (N_6446,N_6078,N_6199);
nand U6447 (N_6447,N_6144,N_6099);
or U6448 (N_6448,N_6207,N_6007);
and U6449 (N_6449,N_6198,N_6024);
or U6450 (N_6450,N_6230,N_6199);
and U6451 (N_6451,N_6140,N_6093);
and U6452 (N_6452,N_6167,N_6042);
and U6453 (N_6453,N_6009,N_6138);
xnor U6454 (N_6454,N_6164,N_6016);
xor U6455 (N_6455,N_6008,N_6190);
or U6456 (N_6456,N_6125,N_6084);
nor U6457 (N_6457,N_6004,N_6196);
or U6458 (N_6458,N_6072,N_6083);
nor U6459 (N_6459,N_6200,N_6237);
or U6460 (N_6460,N_6065,N_6142);
xnor U6461 (N_6461,N_6000,N_6064);
nor U6462 (N_6462,N_6175,N_6247);
and U6463 (N_6463,N_6035,N_6210);
and U6464 (N_6464,N_6087,N_6198);
and U6465 (N_6465,N_6227,N_6127);
and U6466 (N_6466,N_6231,N_6043);
nand U6467 (N_6467,N_6193,N_6144);
nor U6468 (N_6468,N_6110,N_6074);
or U6469 (N_6469,N_6148,N_6067);
and U6470 (N_6470,N_6238,N_6045);
xor U6471 (N_6471,N_6050,N_6026);
or U6472 (N_6472,N_6139,N_6104);
xnor U6473 (N_6473,N_6006,N_6091);
nand U6474 (N_6474,N_6195,N_6024);
nand U6475 (N_6475,N_6201,N_6035);
nor U6476 (N_6476,N_6232,N_6179);
xor U6477 (N_6477,N_6025,N_6054);
and U6478 (N_6478,N_6086,N_6047);
or U6479 (N_6479,N_6097,N_6063);
nand U6480 (N_6480,N_6219,N_6197);
and U6481 (N_6481,N_6097,N_6048);
xor U6482 (N_6482,N_6041,N_6054);
nand U6483 (N_6483,N_6120,N_6096);
nor U6484 (N_6484,N_6111,N_6030);
nor U6485 (N_6485,N_6064,N_6133);
nor U6486 (N_6486,N_6106,N_6232);
nand U6487 (N_6487,N_6101,N_6089);
xnor U6488 (N_6488,N_6018,N_6220);
and U6489 (N_6489,N_6100,N_6073);
or U6490 (N_6490,N_6182,N_6014);
nor U6491 (N_6491,N_6233,N_6225);
and U6492 (N_6492,N_6038,N_6065);
and U6493 (N_6493,N_6146,N_6141);
nand U6494 (N_6494,N_6007,N_6225);
nand U6495 (N_6495,N_6184,N_6099);
nor U6496 (N_6496,N_6023,N_6159);
and U6497 (N_6497,N_6212,N_6048);
nor U6498 (N_6498,N_6018,N_6195);
nand U6499 (N_6499,N_6166,N_6089);
or U6500 (N_6500,N_6416,N_6422);
nand U6501 (N_6501,N_6258,N_6291);
nand U6502 (N_6502,N_6478,N_6482);
or U6503 (N_6503,N_6495,N_6434);
or U6504 (N_6504,N_6448,N_6286);
nor U6505 (N_6505,N_6271,N_6362);
nor U6506 (N_6506,N_6491,N_6488);
and U6507 (N_6507,N_6326,N_6479);
nor U6508 (N_6508,N_6320,N_6367);
and U6509 (N_6509,N_6463,N_6436);
xnor U6510 (N_6510,N_6363,N_6487);
or U6511 (N_6511,N_6441,N_6270);
nand U6512 (N_6512,N_6498,N_6499);
nand U6513 (N_6513,N_6486,N_6267);
nand U6514 (N_6514,N_6398,N_6407);
and U6515 (N_6515,N_6358,N_6254);
and U6516 (N_6516,N_6447,N_6380);
nand U6517 (N_6517,N_6364,N_6366);
nor U6518 (N_6518,N_6266,N_6356);
or U6519 (N_6519,N_6400,N_6328);
xnor U6520 (N_6520,N_6315,N_6283);
nor U6521 (N_6521,N_6449,N_6395);
nand U6522 (N_6522,N_6373,N_6311);
and U6523 (N_6523,N_6327,N_6393);
xor U6524 (N_6524,N_6308,N_6470);
or U6525 (N_6525,N_6300,N_6466);
or U6526 (N_6526,N_6303,N_6494);
nand U6527 (N_6527,N_6288,N_6287);
nor U6528 (N_6528,N_6299,N_6314);
xnor U6529 (N_6529,N_6361,N_6445);
nand U6530 (N_6530,N_6250,N_6438);
nand U6531 (N_6531,N_6337,N_6329);
and U6532 (N_6532,N_6277,N_6483);
or U6533 (N_6533,N_6325,N_6317);
xnor U6534 (N_6534,N_6323,N_6379);
or U6535 (N_6535,N_6489,N_6424);
and U6536 (N_6536,N_6374,N_6289);
xor U6537 (N_6537,N_6340,N_6412);
and U6538 (N_6538,N_6414,N_6342);
or U6539 (N_6539,N_6410,N_6294);
xor U6540 (N_6540,N_6481,N_6349);
or U6541 (N_6541,N_6425,N_6475);
nor U6542 (N_6542,N_6275,N_6420);
and U6543 (N_6543,N_6456,N_6484);
nand U6544 (N_6544,N_6406,N_6344);
or U6545 (N_6545,N_6391,N_6359);
xor U6546 (N_6546,N_6280,N_6397);
nand U6547 (N_6547,N_6457,N_6432);
or U6548 (N_6548,N_6353,N_6492);
xnor U6549 (N_6549,N_6313,N_6474);
xnor U6550 (N_6550,N_6260,N_6357);
nand U6551 (N_6551,N_6490,N_6429);
nand U6552 (N_6552,N_6433,N_6255);
xor U6553 (N_6553,N_6450,N_6351);
xnor U6554 (N_6554,N_6385,N_6465);
nand U6555 (N_6555,N_6252,N_6290);
and U6556 (N_6556,N_6442,N_6348);
nand U6557 (N_6557,N_6335,N_6274);
xor U6558 (N_6558,N_6439,N_6321);
xor U6559 (N_6559,N_6440,N_6467);
xor U6560 (N_6560,N_6316,N_6455);
nand U6561 (N_6561,N_6281,N_6382);
xor U6562 (N_6562,N_6383,N_6346);
or U6563 (N_6563,N_6427,N_6464);
or U6564 (N_6564,N_6411,N_6302);
and U6565 (N_6565,N_6471,N_6403);
nor U6566 (N_6566,N_6417,N_6387);
and U6567 (N_6567,N_6268,N_6339);
or U6568 (N_6568,N_6347,N_6307);
and U6569 (N_6569,N_6437,N_6345);
xor U6570 (N_6570,N_6298,N_6360);
xor U6571 (N_6571,N_6322,N_6409);
xor U6572 (N_6572,N_6381,N_6350);
and U6573 (N_6573,N_6306,N_6384);
xnor U6574 (N_6574,N_6338,N_6333);
nor U6575 (N_6575,N_6369,N_6454);
and U6576 (N_6576,N_6394,N_6423);
and U6577 (N_6577,N_6365,N_6269);
or U6578 (N_6578,N_6278,N_6377);
or U6579 (N_6579,N_6451,N_6485);
or U6580 (N_6580,N_6415,N_6458);
or U6581 (N_6581,N_6336,N_6309);
and U6582 (N_6582,N_6477,N_6405);
nor U6583 (N_6583,N_6392,N_6472);
xor U6584 (N_6584,N_6334,N_6276);
or U6585 (N_6585,N_6324,N_6401);
or U6586 (N_6586,N_6408,N_6459);
nor U6587 (N_6587,N_6284,N_6295);
nand U6588 (N_6588,N_6341,N_6435);
or U6589 (N_6589,N_6476,N_6468);
xnor U6590 (N_6590,N_6431,N_6460);
or U6591 (N_6591,N_6402,N_6305);
xor U6592 (N_6592,N_6388,N_6292);
nand U6593 (N_6593,N_6297,N_6413);
xor U6594 (N_6594,N_6404,N_6396);
or U6595 (N_6595,N_6473,N_6371);
and U6596 (N_6596,N_6426,N_6310);
and U6597 (N_6597,N_6386,N_6462);
or U6598 (N_6598,N_6376,N_6419);
and U6599 (N_6599,N_6272,N_6265);
xor U6600 (N_6600,N_6256,N_6354);
or U6601 (N_6601,N_6319,N_6352);
and U6602 (N_6602,N_6461,N_6452);
nor U6603 (N_6603,N_6261,N_6343);
and U6604 (N_6604,N_6332,N_6262);
and U6605 (N_6605,N_6469,N_6446);
nand U6606 (N_6606,N_6285,N_6331);
and U6607 (N_6607,N_6355,N_6428);
nand U6608 (N_6608,N_6253,N_6330);
nor U6609 (N_6609,N_6421,N_6430);
nand U6610 (N_6610,N_6378,N_6444);
xor U6611 (N_6611,N_6251,N_6318);
and U6612 (N_6612,N_6375,N_6279);
and U6613 (N_6613,N_6312,N_6480);
nor U6614 (N_6614,N_6282,N_6496);
and U6615 (N_6615,N_6273,N_6368);
or U6616 (N_6616,N_6453,N_6257);
xnor U6617 (N_6617,N_6493,N_6443);
nand U6618 (N_6618,N_6264,N_6259);
or U6619 (N_6619,N_6304,N_6418);
or U6620 (N_6620,N_6497,N_6293);
nand U6621 (N_6621,N_6263,N_6399);
or U6622 (N_6622,N_6372,N_6389);
nand U6623 (N_6623,N_6301,N_6370);
nor U6624 (N_6624,N_6296,N_6390);
nor U6625 (N_6625,N_6477,N_6284);
and U6626 (N_6626,N_6323,N_6435);
nor U6627 (N_6627,N_6415,N_6463);
nor U6628 (N_6628,N_6362,N_6477);
nand U6629 (N_6629,N_6262,N_6253);
nor U6630 (N_6630,N_6272,N_6429);
and U6631 (N_6631,N_6356,N_6461);
or U6632 (N_6632,N_6258,N_6377);
nand U6633 (N_6633,N_6345,N_6269);
and U6634 (N_6634,N_6493,N_6408);
nor U6635 (N_6635,N_6397,N_6331);
or U6636 (N_6636,N_6479,N_6366);
nor U6637 (N_6637,N_6483,N_6327);
and U6638 (N_6638,N_6359,N_6283);
xor U6639 (N_6639,N_6396,N_6266);
nor U6640 (N_6640,N_6253,N_6285);
or U6641 (N_6641,N_6333,N_6472);
or U6642 (N_6642,N_6371,N_6376);
nor U6643 (N_6643,N_6403,N_6346);
and U6644 (N_6644,N_6355,N_6388);
nand U6645 (N_6645,N_6298,N_6469);
and U6646 (N_6646,N_6468,N_6275);
and U6647 (N_6647,N_6384,N_6444);
nand U6648 (N_6648,N_6489,N_6444);
xor U6649 (N_6649,N_6299,N_6306);
xor U6650 (N_6650,N_6301,N_6457);
or U6651 (N_6651,N_6495,N_6369);
nand U6652 (N_6652,N_6316,N_6320);
and U6653 (N_6653,N_6384,N_6484);
or U6654 (N_6654,N_6271,N_6406);
and U6655 (N_6655,N_6445,N_6403);
nand U6656 (N_6656,N_6407,N_6336);
and U6657 (N_6657,N_6484,N_6344);
and U6658 (N_6658,N_6474,N_6449);
or U6659 (N_6659,N_6256,N_6260);
nand U6660 (N_6660,N_6464,N_6471);
or U6661 (N_6661,N_6423,N_6430);
xnor U6662 (N_6662,N_6295,N_6390);
or U6663 (N_6663,N_6409,N_6465);
or U6664 (N_6664,N_6271,N_6262);
nand U6665 (N_6665,N_6296,N_6318);
or U6666 (N_6666,N_6480,N_6406);
xor U6667 (N_6667,N_6411,N_6336);
xor U6668 (N_6668,N_6392,N_6354);
or U6669 (N_6669,N_6449,N_6380);
nand U6670 (N_6670,N_6389,N_6349);
or U6671 (N_6671,N_6352,N_6451);
nand U6672 (N_6672,N_6295,N_6341);
xnor U6673 (N_6673,N_6465,N_6332);
nor U6674 (N_6674,N_6496,N_6291);
nor U6675 (N_6675,N_6356,N_6375);
nand U6676 (N_6676,N_6284,N_6413);
nor U6677 (N_6677,N_6466,N_6274);
nand U6678 (N_6678,N_6360,N_6411);
nor U6679 (N_6679,N_6271,N_6358);
and U6680 (N_6680,N_6368,N_6394);
nor U6681 (N_6681,N_6449,N_6340);
nor U6682 (N_6682,N_6297,N_6437);
xor U6683 (N_6683,N_6274,N_6272);
nand U6684 (N_6684,N_6481,N_6493);
or U6685 (N_6685,N_6478,N_6496);
or U6686 (N_6686,N_6275,N_6379);
nand U6687 (N_6687,N_6329,N_6386);
and U6688 (N_6688,N_6479,N_6398);
nand U6689 (N_6689,N_6298,N_6421);
xnor U6690 (N_6690,N_6286,N_6478);
nor U6691 (N_6691,N_6441,N_6305);
xnor U6692 (N_6692,N_6360,N_6459);
xor U6693 (N_6693,N_6334,N_6364);
xnor U6694 (N_6694,N_6309,N_6260);
xnor U6695 (N_6695,N_6262,N_6341);
and U6696 (N_6696,N_6345,N_6311);
and U6697 (N_6697,N_6354,N_6434);
and U6698 (N_6698,N_6482,N_6389);
nor U6699 (N_6699,N_6438,N_6386);
nand U6700 (N_6700,N_6465,N_6429);
and U6701 (N_6701,N_6304,N_6448);
nor U6702 (N_6702,N_6286,N_6272);
or U6703 (N_6703,N_6287,N_6271);
nor U6704 (N_6704,N_6474,N_6323);
or U6705 (N_6705,N_6426,N_6434);
or U6706 (N_6706,N_6332,N_6417);
nor U6707 (N_6707,N_6471,N_6252);
nor U6708 (N_6708,N_6461,N_6312);
xor U6709 (N_6709,N_6277,N_6334);
and U6710 (N_6710,N_6336,N_6354);
nand U6711 (N_6711,N_6301,N_6464);
and U6712 (N_6712,N_6491,N_6266);
xnor U6713 (N_6713,N_6277,N_6274);
nor U6714 (N_6714,N_6481,N_6479);
or U6715 (N_6715,N_6402,N_6288);
or U6716 (N_6716,N_6435,N_6272);
and U6717 (N_6717,N_6277,N_6281);
nor U6718 (N_6718,N_6347,N_6419);
or U6719 (N_6719,N_6464,N_6388);
or U6720 (N_6720,N_6461,N_6487);
nor U6721 (N_6721,N_6422,N_6474);
xor U6722 (N_6722,N_6355,N_6492);
nand U6723 (N_6723,N_6361,N_6268);
xnor U6724 (N_6724,N_6496,N_6464);
or U6725 (N_6725,N_6488,N_6281);
and U6726 (N_6726,N_6445,N_6270);
or U6727 (N_6727,N_6463,N_6337);
xnor U6728 (N_6728,N_6366,N_6430);
and U6729 (N_6729,N_6273,N_6394);
xnor U6730 (N_6730,N_6469,N_6250);
or U6731 (N_6731,N_6387,N_6292);
and U6732 (N_6732,N_6365,N_6416);
and U6733 (N_6733,N_6375,N_6483);
or U6734 (N_6734,N_6397,N_6390);
xnor U6735 (N_6735,N_6309,N_6357);
nand U6736 (N_6736,N_6479,N_6380);
nor U6737 (N_6737,N_6271,N_6378);
nand U6738 (N_6738,N_6343,N_6300);
and U6739 (N_6739,N_6487,N_6315);
or U6740 (N_6740,N_6318,N_6252);
nor U6741 (N_6741,N_6461,N_6311);
or U6742 (N_6742,N_6293,N_6396);
xnor U6743 (N_6743,N_6358,N_6297);
nor U6744 (N_6744,N_6410,N_6375);
or U6745 (N_6745,N_6364,N_6495);
nor U6746 (N_6746,N_6452,N_6446);
nand U6747 (N_6747,N_6369,N_6450);
or U6748 (N_6748,N_6460,N_6450);
nor U6749 (N_6749,N_6352,N_6459);
and U6750 (N_6750,N_6631,N_6645);
and U6751 (N_6751,N_6591,N_6578);
and U6752 (N_6752,N_6512,N_6683);
and U6753 (N_6753,N_6704,N_6731);
xor U6754 (N_6754,N_6722,N_6543);
xnor U6755 (N_6755,N_6650,N_6715);
nand U6756 (N_6756,N_6506,N_6700);
or U6757 (N_6757,N_6596,N_6565);
or U6758 (N_6758,N_6597,N_6570);
nor U6759 (N_6759,N_6706,N_6646);
and U6760 (N_6760,N_6503,N_6576);
and U6761 (N_6761,N_6654,N_6564);
or U6762 (N_6762,N_6699,N_6644);
or U6763 (N_6763,N_6531,N_6516);
nand U6764 (N_6764,N_6648,N_6659);
nand U6765 (N_6765,N_6669,N_6737);
or U6766 (N_6766,N_6628,N_6657);
or U6767 (N_6767,N_6519,N_6729);
nor U6768 (N_6768,N_6745,N_6690);
nand U6769 (N_6769,N_6610,N_6710);
and U6770 (N_6770,N_6664,N_6600);
nand U6771 (N_6771,N_6542,N_6741);
xnor U6772 (N_6772,N_6556,N_6629);
xor U6773 (N_6773,N_6599,N_6685);
nor U6774 (N_6774,N_6551,N_6589);
xor U6775 (N_6775,N_6530,N_6658);
nor U6776 (N_6776,N_6619,N_6637);
and U6777 (N_6777,N_6559,N_6529);
nand U6778 (N_6778,N_6539,N_6705);
xnor U6779 (N_6779,N_6555,N_6712);
nor U6780 (N_6780,N_6742,N_6535);
and U6781 (N_6781,N_6508,N_6566);
or U6782 (N_6782,N_6667,N_6515);
xor U6783 (N_6783,N_6518,N_6688);
and U6784 (N_6784,N_6725,N_6723);
nand U6785 (N_6785,N_6582,N_6560);
nand U6786 (N_6786,N_6744,N_6671);
xor U6787 (N_6787,N_6572,N_6740);
xor U6788 (N_6788,N_6525,N_6602);
nor U6789 (N_6789,N_6623,N_6717);
and U6790 (N_6790,N_6630,N_6580);
and U6791 (N_6791,N_6532,N_6636);
nor U6792 (N_6792,N_6670,N_6672);
nor U6793 (N_6793,N_6677,N_6579);
or U6794 (N_6794,N_6546,N_6714);
nand U6795 (N_6795,N_6733,N_6562);
and U6796 (N_6796,N_6627,N_6513);
and U6797 (N_6797,N_6656,N_6625);
xnor U6798 (N_6798,N_6526,N_6590);
and U6799 (N_6799,N_6703,N_6614);
nor U6800 (N_6800,N_6675,N_6568);
xnor U6801 (N_6801,N_6608,N_6689);
nor U6802 (N_6802,N_6738,N_6621);
nand U6803 (N_6803,N_6514,N_6624);
xor U6804 (N_6804,N_6674,N_6634);
or U6805 (N_6805,N_6702,N_6563);
and U6806 (N_6806,N_6618,N_6713);
xnor U6807 (N_6807,N_6684,N_6523);
or U6808 (N_6808,N_6719,N_6528);
or U6809 (N_6809,N_6524,N_6538);
xnor U6810 (N_6810,N_6598,N_6718);
or U6811 (N_6811,N_6517,N_6541);
xor U6812 (N_6812,N_6651,N_6569);
xor U6813 (N_6813,N_6661,N_6607);
nand U6814 (N_6814,N_6522,N_6653);
nor U6815 (N_6815,N_6584,N_6633);
xor U6816 (N_6816,N_6693,N_6691);
or U6817 (N_6817,N_6509,N_6694);
and U6818 (N_6818,N_6507,N_6680);
nand U6819 (N_6819,N_6743,N_6553);
and U6820 (N_6820,N_6626,N_6749);
nand U6821 (N_6821,N_6652,N_6545);
nor U6822 (N_6822,N_6649,N_6716);
and U6823 (N_6823,N_6534,N_6550);
and U6824 (N_6824,N_6708,N_6615);
nor U6825 (N_6825,N_6587,N_6605);
nand U6826 (N_6826,N_6592,N_6701);
and U6827 (N_6827,N_6662,N_6609);
and U6828 (N_6828,N_6501,N_6593);
or U6829 (N_6829,N_6622,N_6549);
and U6830 (N_6830,N_6696,N_6581);
and U6831 (N_6831,N_6521,N_6594);
nand U6832 (N_6832,N_6660,N_6668);
nand U6833 (N_6833,N_6724,N_6692);
xor U6834 (N_6834,N_6505,N_6574);
xnor U6835 (N_6835,N_6681,N_6611);
and U6836 (N_6836,N_6746,N_6736);
nor U6837 (N_6837,N_6620,N_6616);
and U6838 (N_6838,N_6720,N_6663);
xor U6839 (N_6839,N_6561,N_6732);
or U6840 (N_6840,N_6640,N_6728);
and U6841 (N_6841,N_6540,N_6588);
nor U6842 (N_6842,N_6695,N_6655);
nand U6843 (N_6843,N_6606,N_6638);
or U6844 (N_6844,N_6601,N_6697);
nand U6845 (N_6845,N_6642,N_6604);
nand U6846 (N_6846,N_6726,N_6721);
xor U6847 (N_6847,N_6739,N_6573);
or U6848 (N_6848,N_6504,N_6665);
xor U6849 (N_6849,N_6586,N_6643);
nand U6850 (N_6850,N_6554,N_6500);
and U6851 (N_6851,N_6673,N_6679);
and U6852 (N_6852,N_6635,N_6536);
nand U6853 (N_6853,N_6686,N_6502);
and U6854 (N_6854,N_6547,N_6617);
xnor U6855 (N_6855,N_6577,N_6595);
nor U6856 (N_6856,N_6558,N_6510);
or U6857 (N_6857,N_6612,N_6647);
nand U6858 (N_6858,N_6709,N_6571);
and U6859 (N_6859,N_6698,N_6676);
nand U6860 (N_6860,N_6567,N_6537);
or U6861 (N_6861,N_6552,N_6533);
xor U6862 (N_6862,N_6730,N_6632);
nand U6863 (N_6863,N_6735,N_6585);
or U6864 (N_6864,N_6527,N_6557);
nand U6865 (N_6865,N_6520,N_6548);
xnor U6866 (N_6866,N_6727,N_6613);
nand U6867 (N_6867,N_6666,N_6639);
xor U6868 (N_6868,N_6583,N_6682);
and U6869 (N_6869,N_6511,N_6678);
or U6870 (N_6870,N_6747,N_6748);
and U6871 (N_6871,N_6641,N_6544);
nand U6872 (N_6872,N_6603,N_6711);
or U6873 (N_6873,N_6687,N_6707);
and U6874 (N_6874,N_6734,N_6575);
nor U6875 (N_6875,N_6659,N_6506);
nor U6876 (N_6876,N_6614,N_6671);
and U6877 (N_6877,N_6647,N_6565);
and U6878 (N_6878,N_6530,N_6623);
or U6879 (N_6879,N_6511,N_6667);
xor U6880 (N_6880,N_6744,N_6573);
nand U6881 (N_6881,N_6566,N_6522);
xor U6882 (N_6882,N_6536,N_6647);
xnor U6883 (N_6883,N_6565,N_6700);
nor U6884 (N_6884,N_6529,N_6701);
and U6885 (N_6885,N_6623,N_6512);
nand U6886 (N_6886,N_6719,N_6569);
or U6887 (N_6887,N_6678,N_6594);
xor U6888 (N_6888,N_6655,N_6513);
xor U6889 (N_6889,N_6656,N_6575);
nand U6890 (N_6890,N_6701,N_6717);
xor U6891 (N_6891,N_6508,N_6667);
or U6892 (N_6892,N_6705,N_6657);
or U6893 (N_6893,N_6533,N_6526);
nor U6894 (N_6894,N_6600,N_6670);
or U6895 (N_6895,N_6538,N_6722);
nor U6896 (N_6896,N_6529,N_6682);
nand U6897 (N_6897,N_6695,N_6649);
nor U6898 (N_6898,N_6534,N_6692);
and U6899 (N_6899,N_6642,N_6515);
xor U6900 (N_6900,N_6557,N_6518);
or U6901 (N_6901,N_6524,N_6643);
or U6902 (N_6902,N_6618,N_6506);
and U6903 (N_6903,N_6718,N_6641);
or U6904 (N_6904,N_6701,N_6588);
xor U6905 (N_6905,N_6703,N_6636);
nand U6906 (N_6906,N_6644,N_6555);
nand U6907 (N_6907,N_6659,N_6696);
nand U6908 (N_6908,N_6701,N_6679);
and U6909 (N_6909,N_6539,N_6578);
nand U6910 (N_6910,N_6687,N_6578);
nand U6911 (N_6911,N_6638,N_6637);
nand U6912 (N_6912,N_6682,N_6687);
and U6913 (N_6913,N_6656,N_6619);
nand U6914 (N_6914,N_6546,N_6622);
and U6915 (N_6915,N_6527,N_6697);
nor U6916 (N_6916,N_6599,N_6551);
and U6917 (N_6917,N_6563,N_6741);
nor U6918 (N_6918,N_6579,N_6648);
nand U6919 (N_6919,N_6718,N_6597);
nand U6920 (N_6920,N_6577,N_6503);
or U6921 (N_6921,N_6618,N_6642);
xnor U6922 (N_6922,N_6528,N_6535);
nor U6923 (N_6923,N_6577,N_6730);
and U6924 (N_6924,N_6551,N_6715);
or U6925 (N_6925,N_6590,N_6583);
or U6926 (N_6926,N_6734,N_6563);
xor U6927 (N_6927,N_6578,N_6740);
xnor U6928 (N_6928,N_6518,N_6552);
xor U6929 (N_6929,N_6541,N_6514);
and U6930 (N_6930,N_6661,N_6522);
or U6931 (N_6931,N_6526,N_6695);
or U6932 (N_6932,N_6626,N_6722);
nor U6933 (N_6933,N_6579,N_6620);
xnor U6934 (N_6934,N_6657,N_6510);
or U6935 (N_6935,N_6510,N_6516);
xnor U6936 (N_6936,N_6705,N_6574);
or U6937 (N_6937,N_6539,N_6568);
xnor U6938 (N_6938,N_6635,N_6702);
nor U6939 (N_6939,N_6734,N_6542);
nand U6940 (N_6940,N_6588,N_6599);
nand U6941 (N_6941,N_6597,N_6591);
xnor U6942 (N_6942,N_6694,N_6699);
xnor U6943 (N_6943,N_6565,N_6632);
or U6944 (N_6944,N_6539,N_6585);
nor U6945 (N_6945,N_6666,N_6562);
or U6946 (N_6946,N_6635,N_6737);
or U6947 (N_6947,N_6700,N_6671);
nand U6948 (N_6948,N_6747,N_6722);
nand U6949 (N_6949,N_6653,N_6727);
nand U6950 (N_6950,N_6694,N_6639);
and U6951 (N_6951,N_6662,N_6729);
xnor U6952 (N_6952,N_6607,N_6536);
nor U6953 (N_6953,N_6606,N_6661);
nor U6954 (N_6954,N_6596,N_6563);
or U6955 (N_6955,N_6599,N_6558);
xnor U6956 (N_6956,N_6524,N_6507);
or U6957 (N_6957,N_6524,N_6591);
or U6958 (N_6958,N_6660,N_6532);
nor U6959 (N_6959,N_6579,N_6552);
and U6960 (N_6960,N_6640,N_6543);
xnor U6961 (N_6961,N_6614,N_6691);
and U6962 (N_6962,N_6727,N_6748);
nor U6963 (N_6963,N_6639,N_6543);
or U6964 (N_6964,N_6669,N_6564);
or U6965 (N_6965,N_6629,N_6628);
nand U6966 (N_6966,N_6521,N_6657);
nor U6967 (N_6967,N_6550,N_6692);
nand U6968 (N_6968,N_6716,N_6549);
or U6969 (N_6969,N_6625,N_6626);
nor U6970 (N_6970,N_6699,N_6668);
nor U6971 (N_6971,N_6621,N_6630);
xnor U6972 (N_6972,N_6686,N_6690);
nor U6973 (N_6973,N_6727,N_6517);
nor U6974 (N_6974,N_6527,N_6579);
nor U6975 (N_6975,N_6711,N_6561);
or U6976 (N_6976,N_6583,N_6510);
nand U6977 (N_6977,N_6624,N_6710);
or U6978 (N_6978,N_6606,N_6662);
nand U6979 (N_6979,N_6698,N_6639);
nor U6980 (N_6980,N_6718,N_6653);
nand U6981 (N_6981,N_6581,N_6669);
xnor U6982 (N_6982,N_6543,N_6595);
xor U6983 (N_6983,N_6585,N_6509);
nand U6984 (N_6984,N_6627,N_6568);
nand U6985 (N_6985,N_6652,N_6740);
or U6986 (N_6986,N_6669,N_6552);
nand U6987 (N_6987,N_6607,N_6729);
nor U6988 (N_6988,N_6617,N_6628);
xnor U6989 (N_6989,N_6705,N_6520);
nand U6990 (N_6990,N_6514,N_6671);
or U6991 (N_6991,N_6537,N_6679);
and U6992 (N_6992,N_6590,N_6582);
and U6993 (N_6993,N_6521,N_6578);
and U6994 (N_6994,N_6561,N_6622);
and U6995 (N_6995,N_6706,N_6569);
or U6996 (N_6996,N_6700,N_6536);
xnor U6997 (N_6997,N_6734,N_6654);
xnor U6998 (N_6998,N_6527,N_6637);
or U6999 (N_6999,N_6545,N_6703);
or U7000 (N_7000,N_6814,N_6825);
xnor U7001 (N_7001,N_6781,N_6992);
nand U7002 (N_7002,N_6897,N_6838);
nor U7003 (N_7003,N_6794,N_6760);
and U7004 (N_7004,N_6994,N_6964);
or U7005 (N_7005,N_6753,N_6959);
or U7006 (N_7006,N_6828,N_6792);
xnor U7007 (N_7007,N_6761,N_6784);
or U7008 (N_7008,N_6762,N_6932);
nand U7009 (N_7009,N_6882,N_6770);
nor U7010 (N_7010,N_6970,N_6983);
nor U7011 (N_7011,N_6839,N_6750);
and U7012 (N_7012,N_6955,N_6812);
or U7013 (N_7013,N_6854,N_6914);
and U7014 (N_7014,N_6852,N_6850);
nor U7015 (N_7015,N_6961,N_6858);
or U7016 (N_7016,N_6908,N_6995);
or U7017 (N_7017,N_6796,N_6798);
nor U7018 (N_7018,N_6936,N_6971);
nor U7019 (N_7019,N_6967,N_6901);
and U7020 (N_7020,N_6763,N_6939);
nand U7021 (N_7021,N_6837,N_6900);
nor U7022 (N_7022,N_6870,N_6972);
xor U7023 (N_7023,N_6843,N_6916);
and U7024 (N_7024,N_6980,N_6802);
or U7025 (N_7025,N_6903,N_6787);
nor U7026 (N_7026,N_6960,N_6867);
xnor U7027 (N_7027,N_6944,N_6842);
nand U7028 (N_7028,N_6928,N_6824);
or U7029 (N_7029,N_6772,N_6966);
xor U7030 (N_7030,N_6930,N_6816);
nand U7031 (N_7031,N_6774,N_6764);
or U7032 (N_7032,N_6834,N_6956);
xor U7033 (N_7033,N_6751,N_6769);
nor U7034 (N_7034,N_6889,N_6780);
and U7035 (N_7035,N_6831,N_6855);
nand U7036 (N_7036,N_6880,N_6974);
or U7037 (N_7037,N_6885,N_6946);
or U7038 (N_7038,N_6922,N_6910);
and U7039 (N_7039,N_6847,N_6759);
and U7040 (N_7040,N_6942,N_6976);
xor U7041 (N_7041,N_6913,N_6861);
nand U7042 (N_7042,N_6979,N_6877);
or U7043 (N_7043,N_6921,N_6866);
or U7044 (N_7044,N_6767,N_6795);
and U7045 (N_7045,N_6786,N_6862);
or U7046 (N_7046,N_6904,N_6818);
nand U7047 (N_7047,N_6952,N_6799);
and U7048 (N_7048,N_6841,N_6963);
or U7049 (N_7049,N_6996,N_6776);
xor U7050 (N_7050,N_6895,N_6872);
xor U7051 (N_7051,N_6934,N_6950);
or U7052 (N_7052,N_6815,N_6884);
nor U7053 (N_7053,N_6989,N_6822);
nor U7054 (N_7054,N_6869,N_6782);
nand U7055 (N_7055,N_6832,N_6803);
nor U7056 (N_7056,N_6929,N_6785);
or U7057 (N_7057,N_6986,N_6902);
xor U7058 (N_7058,N_6851,N_6919);
nand U7059 (N_7059,N_6800,N_6982);
and U7060 (N_7060,N_6789,N_6771);
and U7061 (N_7061,N_6819,N_6797);
or U7062 (N_7062,N_6926,N_6990);
and U7063 (N_7063,N_6864,N_6848);
nor U7064 (N_7064,N_6806,N_6933);
and U7065 (N_7065,N_6860,N_6775);
xnor U7066 (N_7066,N_6947,N_6833);
nand U7067 (N_7067,N_6969,N_6925);
nor U7068 (N_7068,N_6788,N_6907);
xor U7069 (N_7069,N_6757,N_6888);
or U7070 (N_7070,N_6845,N_6981);
nand U7071 (N_7071,N_6778,N_6898);
and U7072 (N_7072,N_6840,N_6809);
nor U7073 (N_7073,N_6953,N_6844);
nor U7074 (N_7074,N_6954,N_6937);
xor U7075 (N_7075,N_6958,N_6893);
or U7076 (N_7076,N_6779,N_6951);
or U7077 (N_7077,N_6999,N_6853);
nor U7078 (N_7078,N_6807,N_6755);
nand U7079 (N_7079,N_6924,N_6886);
or U7080 (N_7080,N_6808,N_6856);
xnor U7081 (N_7081,N_6977,N_6873);
nand U7082 (N_7082,N_6957,N_6754);
or U7083 (N_7083,N_6868,N_6909);
and U7084 (N_7084,N_6899,N_6804);
xnor U7085 (N_7085,N_6827,N_6906);
or U7086 (N_7086,N_6810,N_6793);
nor U7087 (N_7087,N_6768,N_6801);
and U7088 (N_7088,N_6859,N_6892);
nand U7089 (N_7089,N_6811,N_6993);
xnor U7090 (N_7090,N_6765,N_6879);
xor U7091 (N_7091,N_6826,N_6766);
and U7092 (N_7092,N_6927,N_6965);
nand U7093 (N_7093,N_6940,N_6985);
xor U7094 (N_7094,N_6871,N_6905);
nor U7095 (N_7095,N_6777,N_6758);
or U7096 (N_7096,N_6987,N_6820);
nand U7097 (N_7097,N_6991,N_6896);
xnor U7098 (N_7098,N_6791,N_6988);
nor U7099 (N_7099,N_6931,N_6783);
and U7100 (N_7100,N_6975,N_6887);
or U7101 (N_7101,N_6876,N_6883);
xor U7102 (N_7102,N_6823,N_6875);
nand U7103 (N_7103,N_6878,N_6849);
and U7104 (N_7104,N_6948,N_6917);
and U7105 (N_7105,N_6923,N_6935);
nor U7106 (N_7106,N_6997,N_6773);
or U7107 (N_7107,N_6821,N_6915);
nor U7108 (N_7108,N_6949,N_6973);
nor U7109 (N_7109,N_6911,N_6920);
xnor U7110 (N_7110,N_6790,N_6756);
and U7111 (N_7111,N_6874,N_6943);
xnor U7112 (N_7112,N_6938,N_6881);
or U7113 (N_7113,N_6945,N_6857);
nand U7114 (N_7114,N_6865,N_6817);
or U7115 (N_7115,N_6912,N_6829);
nand U7116 (N_7116,N_6962,N_6894);
nor U7117 (N_7117,N_6805,N_6941);
nand U7118 (N_7118,N_6890,N_6998);
and U7119 (N_7119,N_6846,N_6918);
and U7120 (N_7120,N_6984,N_6978);
or U7121 (N_7121,N_6891,N_6752);
nor U7122 (N_7122,N_6813,N_6835);
or U7123 (N_7123,N_6863,N_6830);
and U7124 (N_7124,N_6968,N_6836);
and U7125 (N_7125,N_6931,N_6972);
nor U7126 (N_7126,N_6993,N_6871);
and U7127 (N_7127,N_6883,N_6935);
nor U7128 (N_7128,N_6933,N_6751);
xor U7129 (N_7129,N_6818,N_6942);
nand U7130 (N_7130,N_6984,N_6880);
nor U7131 (N_7131,N_6908,N_6827);
and U7132 (N_7132,N_6760,N_6883);
nand U7133 (N_7133,N_6985,N_6757);
nand U7134 (N_7134,N_6890,N_6919);
nand U7135 (N_7135,N_6933,N_6921);
nand U7136 (N_7136,N_6993,N_6971);
nor U7137 (N_7137,N_6969,N_6978);
and U7138 (N_7138,N_6836,N_6762);
nand U7139 (N_7139,N_6804,N_6822);
nand U7140 (N_7140,N_6904,N_6783);
nor U7141 (N_7141,N_6886,N_6860);
or U7142 (N_7142,N_6982,N_6938);
nor U7143 (N_7143,N_6986,N_6966);
nand U7144 (N_7144,N_6943,N_6897);
nand U7145 (N_7145,N_6843,N_6765);
and U7146 (N_7146,N_6922,N_6860);
nor U7147 (N_7147,N_6921,N_6873);
xnor U7148 (N_7148,N_6832,N_6751);
nand U7149 (N_7149,N_6915,N_6904);
and U7150 (N_7150,N_6794,N_6949);
or U7151 (N_7151,N_6860,N_6865);
or U7152 (N_7152,N_6907,N_6753);
nor U7153 (N_7153,N_6915,N_6803);
xor U7154 (N_7154,N_6803,N_6872);
nor U7155 (N_7155,N_6961,N_6846);
nand U7156 (N_7156,N_6847,N_6958);
xor U7157 (N_7157,N_6946,N_6893);
or U7158 (N_7158,N_6871,N_6953);
nor U7159 (N_7159,N_6916,N_6859);
xnor U7160 (N_7160,N_6766,N_6987);
and U7161 (N_7161,N_6873,N_6932);
or U7162 (N_7162,N_6794,N_6942);
and U7163 (N_7163,N_6876,N_6935);
or U7164 (N_7164,N_6779,N_6797);
xnor U7165 (N_7165,N_6787,N_6917);
nor U7166 (N_7166,N_6863,N_6984);
nand U7167 (N_7167,N_6847,N_6912);
and U7168 (N_7168,N_6985,N_6809);
nor U7169 (N_7169,N_6766,N_6863);
xnor U7170 (N_7170,N_6799,N_6786);
or U7171 (N_7171,N_6815,N_6930);
nand U7172 (N_7172,N_6954,N_6863);
xor U7173 (N_7173,N_6786,N_6950);
or U7174 (N_7174,N_6970,N_6974);
nand U7175 (N_7175,N_6905,N_6815);
or U7176 (N_7176,N_6822,N_6887);
or U7177 (N_7177,N_6821,N_6951);
nor U7178 (N_7178,N_6951,N_6828);
nor U7179 (N_7179,N_6776,N_6819);
and U7180 (N_7180,N_6751,N_6994);
nor U7181 (N_7181,N_6804,N_6785);
nand U7182 (N_7182,N_6896,N_6860);
xor U7183 (N_7183,N_6897,N_6953);
nor U7184 (N_7184,N_6933,N_6859);
or U7185 (N_7185,N_6965,N_6860);
nor U7186 (N_7186,N_6977,N_6961);
xnor U7187 (N_7187,N_6841,N_6991);
and U7188 (N_7188,N_6836,N_6830);
nand U7189 (N_7189,N_6871,N_6934);
nand U7190 (N_7190,N_6765,N_6856);
or U7191 (N_7191,N_6926,N_6750);
or U7192 (N_7192,N_6806,N_6759);
nor U7193 (N_7193,N_6821,N_6752);
xnor U7194 (N_7194,N_6922,N_6778);
nor U7195 (N_7195,N_6920,N_6971);
nand U7196 (N_7196,N_6900,N_6915);
nor U7197 (N_7197,N_6823,N_6836);
nand U7198 (N_7198,N_6942,N_6832);
and U7199 (N_7199,N_6797,N_6802);
xor U7200 (N_7200,N_6903,N_6925);
xor U7201 (N_7201,N_6886,N_6775);
and U7202 (N_7202,N_6776,N_6973);
or U7203 (N_7203,N_6883,N_6999);
xor U7204 (N_7204,N_6797,N_6917);
nor U7205 (N_7205,N_6936,N_6828);
nor U7206 (N_7206,N_6799,N_6894);
and U7207 (N_7207,N_6940,N_6986);
and U7208 (N_7208,N_6932,N_6926);
nand U7209 (N_7209,N_6780,N_6868);
nand U7210 (N_7210,N_6959,N_6880);
or U7211 (N_7211,N_6878,N_6975);
nand U7212 (N_7212,N_6980,N_6997);
or U7213 (N_7213,N_6882,N_6802);
or U7214 (N_7214,N_6753,N_6859);
and U7215 (N_7215,N_6982,N_6841);
nor U7216 (N_7216,N_6865,N_6996);
xnor U7217 (N_7217,N_6881,N_6896);
and U7218 (N_7218,N_6783,N_6935);
nor U7219 (N_7219,N_6885,N_6910);
nor U7220 (N_7220,N_6966,N_6859);
nor U7221 (N_7221,N_6815,N_6999);
xnor U7222 (N_7222,N_6861,N_6877);
and U7223 (N_7223,N_6830,N_6944);
and U7224 (N_7224,N_6825,N_6857);
or U7225 (N_7225,N_6766,N_6777);
nand U7226 (N_7226,N_6997,N_6788);
nand U7227 (N_7227,N_6997,N_6927);
nor U7228 (N_7228,N_6932,N_6855);
or U7229 (N_7229,N_6835,N_6918);
nor U7230 (N_7230,N_6899,N_6872);
nor U7231 (N_7231,N_6958,N_6826);
nor U7232 (N_7232,N_6887,N_6957);
nand U7233 (N_7233,N_6833,N_6985);
or U7234 (N_7234,N_6798,N_6876);
nand U7235 (N_7235,N_6755,N_6927);
nor U7236 (N_7236,N_6805,N_6864);
or U7237 (N_7237,N_6865,N_6920);
or U7238 (N_7238,N_6841,N_6886);
xnor U7239 (N_7239,N_6865,N_6963);
xor U7240 (N_7240,N_6760,N_6754);
or U7241 (N_7241,N_6918,N_6951);
xor U7242 (N_7242,N_6766,N_6943);
and U7243 (N_7243,N_6790,N_6917);
and U7244 (N_7244,N_6996,N_6920);
or U7245 (N_7245,N_6936,N_6778);
and U7246 (N_7246,N_6791,N_6768);
or U7247 (N_7247,N_6979,N_6776);
xnor U7248 (N_7248,N_6902,N_6918);
nor U7249 (N_7249,N_6956,N_6779);
nor U7250 (N_7250,N_7073,N_7072);
nand U7251 (N_7251,N_7143,N_7112);
nor U7252 (N_7252,N_7012,N_7148);
and U7253 (N_7253,N_7240,N_7055);
and U7254 (N_7254,N_7115,N_7183);
and U7255 (N_7255,N_7149,N_7002);
or U7256 (N_7256,N_7160,N_7135);
nand U7257 (N_7257,N_7169,N_7178);
nor U7258 (N_7258,N_7232,N_7120);
and U7259 (N_7259,N_7096,N_7039);
nand U7260 (N_7260,N_7062,N_7199);
or U7261 (N_7261,N_7237,N_7031);
and U7262 (N_7262,N_7027,N_7035);
xor U7263 (N_7263,N_7025,N_7090);
xnor U7264 (N_7264,N_7011,N_7059);
nand U7265 (N_7265,N_7197,N_7053);
nand U7266 (N_7266,N_7229,N_7085);
or U7267 (N_7267,N_7164,N_7171);
nor U7268 (N_7268,N_7210,N_7125);
nand U7269 (N_7269,N_7081,N_7185);
xor U7270 (N_7270,N_7168,N_7196);
and U7271 (N_7271,N_7058,N_7216);
xnor U7272 (N_7272,N_7119,N_7167);
or U7273 (N_7273,N_7147,N_7150);
or U7274 (N_7274,N_7067,N_7004);
or U7275 (N_7275,N_7220,N_7079);
nand U7276 (N_7276,N_7241,N_7231);
nand U7277 (N_7277,N_7034,N_7188);
or U7278 (N_7278,N_7044,N_7130);
nor U7279 (N_7279,N_7218,N_7211);
and U7280 (N_7280,N_7245,N_7207);
or U7281 (N_7281,N_7172,N_7091);
nor U7282 (N_7282,N_7138,N_7180);
xor U7283 (N_7283,N_7202,N_7175);
or U7284 (N_7284,N_7032,N_7113);
or U7285 (N_7285,N_7024,N_7152);
xnor U7286 (N_7286,N_7166,N_7097);
nand U7287 (N_7287,N_7092,N_7154);
and U7288 (N_7288,N_7228,N_7206);
xnor U7289 (N_7289,N_7177,N_7005);
nor U7290 (N_7290,N_7007,N_7040);
xor U7291 (N_7291,N_7239,N_7118);
nor U7292 (N_7292,N_7227,N_7129);
or U7293 (N_7293,N_7111,N_7095);
and U7294 (N_7294,N_7158,N_7132);
xor U7295 (N_7295,N_7198,N_7144);
nor U7296 (N_7296,N_7061,N_7023);
xor U7297 (N_7297,N_7139,N_7137);
xor U7298 (N_7298,N_7030,N_7057);
xnor U7299 (N_7299,N_7200,N_7010);
nand U7300 (N_7300,N_7236,N_7161);
nor U7301 (N_7301,N_7056,N_7131);
or U7302 (N_7302,N_7013,N_7190);
and U7303 (N_7303,N_7153,N_7243);
or U7304 (N_7304,N_7181,N_7068);
nor U7305 (N_7305,N_7046,N_7033);
and U7306 (N_7306,N_7234,N_7014);
or U7307 (N_7307,N_7098,N_7075);
and U7308 (N_7308,N_7204,N_7174);
and U7309 (N_7309,N_7176,N_7047);
nor U7310 (N_7310,N_7018,N_7222);
or U7311 (N_7311,N_7116,N_7248);
nor U7312 (N_7312,N_7121,N_7109);
or U7313 (N_7313,N_7224,N_7187);
xnor U7314 (N_7314,N_7063,N_7173);
nor U7315 (N_7315,N_7221,N_7008);
nor U7316 (N_7316,N_7186,N_7117);
and U7317 (N_7317,N_7155,N_7145);
xnor U7318 (N_7318,N_7006,N_7193);
nand U7319 (N_7319,N_7191,N_7105);
xor U7320 (N_7320,N_7069,N_7015);
nand U7321 (N_7321,N_7048,N_7142);
and U7322 (N_7322,N_7163,N_7065);
and U7323 (N_7323,N_7165,N_7212);
nand U7324 (N_7324,N_7123,N_7242);
and U7325 (N_7325,N_7009,N_7026);
xor U7326 (N_7326,N_7028,N_7052);
or U7327 (N_7327,N_7076,N_7208);
or U7328 (N_7328,N_7101,N_7136);
or U7329 (N_7329,N_7214,N_7050);
nor U7330 (N_7330,N_7088,N_7184);
and U7331 (N_7331,N_7080,N_7146);
xor U7332 (N_7332,N_7049,N_7247);
nor U7333 (N_7333,N_7094,N_7107);
nand U7334 (N_7334,N_7084,N_7122);
and U7335 (N_7335,N_7156,N_7003);
xnor U7336 (N_7336,N_7124,N_7205);
and U7337 (N_7337,N_7082,N_7128);
nand U7338 (N_7338,N_7083,N_7189);
xor U7339 (N_7339,N_7041,N_7022);
xnor U7340 (N_7340,N_7110,N_7192);
xnor U7341 (N_7341,N_7230,N_7086);
nor U7342 (N_7342,N_7042,N_7066);
nand U7343 (N_7343,N_7219,N_7246);
and U7344 (N_7344,N_7159,N_7127);
xor U7345 (N_7345,N_7141,N_7064);
nor U7346 (N_7346,N_7104,N_7102);
nand U7347 (N_7347,N_7021,N_7179);
nor U7348 (N_7348,N_7223,N_7060);
and U7349 (N_7349,N_7225,N_7038);
or U7350 (N_7350,N_7249,N_7020);
nor U7351 (N_7351,N_7087,N_7201);
and U7352 (N_7352,N_7213,N_7140);
nor U7353 (N_7353,N_7162,N_7051);
nor U7354 (N_7354,N_7077,N_7233);
nand U7355 (N_7355,N_7203,N_7194);
xnor U7356 (N_7356,N_7114,N_7019);
and U7357 (N_7357,N_7226,N_7235);
nand U7358 (N_7358,N_7215,N_7054);
or U7359 (N_7359,N_7037,N_7103);
and U7360 (N_7360,N_7089,N_7016);
and U7361 (N_7361,N_7182,N_7074);
nand U7362 (N_7362,N_7001,N_7170);
xnor U7363 (N_7363,N_7106,N_7078);
nand U7364 (N_7364,N_7043,N_7244);
or U7365 (N_7365,N_7133,N_7151);
nand U7366 (N_7366,N_7126,N_7070);
xor U7367 (N_7367,N_7238,N_7134);
or U7368 (N_7368,N_7209,N_7195);
nor U7369 (N_7369,N_7093,N_7217);
and U7370 (N_7370,N_7100,N_7029);
xor U7371 (N_7371,N_7071,N_7000);
and U7372 (N_7372,N_7108,N_7157);
xor U7373 (N_7373,N_7099,N_7045);
nor U7374 (N_7374,N_7036,N_7017);
nand U7375 (N_7375,N_7018,N_7242);
nor U7376 (N_7376,N_7112,N_7072);
or U7377 (N_7377,N_7151,N_7225);
and U7378 (N_7378,N_7146,N_7035);
or U7379 (N_7379,N_7008,N_7039);
and U7380 (N_7380,N_7036,N_7080);
nand U7381 (N_7381,N_7095,N_7084);
xor U7382 (N_7382,N_7190,N_7041);
nand U7383 (N_7383,N_7138,N_7143);
nand U7384 (N_7384,N_7112,N_7026);
nor U7385 (N_7385,N_7245,N_7237);
or U7386 (N_7386,N_7218,N_7083);
nand U7387 (N_7387,N_7061,N_7192);
nand U7388 (N_7388,N_7133,N_7134);
nand U7389 (N_7389,N_7148,N_7048);
and U7390 (N_7390,N_7143,N_7073);
nand U7391 (N_7391,N_7055,N_7200);
or U7392 (N_7392,N_7160,N_7053);
and U7393 (N_7393,N_7089,N_7156);
and U7394 (N_7394,N_7063,N_7038);
nand U7395 (N_7395,N_7093,N_7098);
or U7396 (N_7396,N_7142,N_7231);
nand U7397 (N_7397,N_7099,N_7190);
nor U7398 (N_7398,N_7066,N_7057);
and U7399 (N_7399,N_7195,N_7075);
and U7400 (N_7400,N_7199,N_7155);
nor U7401 (N_7401,N_7138,N_7243);
xor U7402 (N_7402,N_7008,N_7111);
xnor U7403 (N_7403,N_7234,N_7138);
nand U7404 (N_7404,N_7227,N_7000);
and U7405 (N_7405,N_7214,N_7197);
nor U7406 (N_7406,N_7234,N_7126);
nor U7407 (N_7407,N_7036,N_7199);
or U7408 (N_7408,N_7133,N_7168);
or U7409 (N_7409,N_7011,N_7079);
or U7410 (N_7410,N_7077,N_7073);
nor U7411 (N_7411,N_7193,N_7153);
xor U7412 (N_7412,N_7196,N_7107);
and U7413 (N_7413,N_7232,N_7172);
xnor U7414 (N_7414,N_7144,N_7040);
nor U7415 (N_7415,N_7170,N_7137);
and U7416 (N_7416,N_7012,N_7230);
and U7417 (N_7417,N_7149,N_7072);
and U7418 (N_7418,N_7016,N_7112);
nor U7419 (N_7419,N_7247,N_7179);
or U7420 (N_7420,N_7017,N_7108);
or U7421 (N_7421,N_7098,N_7084);
or U7422 (N_7422,N_7209,N_7133);
nor U7423 (N_7423,N_7040,N_7032);
and U7424 (N_7424,N_7130,N_7049);
and U7425 (N_7425,N_7065,N_7084);
xor U7426 (N_7426,N_7111,N_7040);
nand U7427 (N_7427,N_7086,N_7060);
nor U7428 (N_7428,N_7043,N_7236);
or U7429 (N_7429,N_7087,N_7107);
xnor U7430 (N_7430,N_7070,N_7031);
nor U7431 (N_7431,N_7219,N_7146);
and U7432 (N_7432,N_7055,N_7249);
xnor U7433 (N_7433,N_7160,N_7203);
nor U7434 (N_7434,N_7014,N_7020);
nor U7435 (N_7435,N_7184,N_7080);
nand U7436 (N_7436,N_7113,N_7188);
and U7437 (N_7437,N_7223,N_7078);
nor U7438 (N_7438,N_7216,N_7229);
xnor U7439 (N_7439,N_7077,N_7201);
nor U7440 (N_7440,N_7248,N_7127);
or U7441 (N_7441,N_7070,N_7124);
xnor U7442 (N_7442,N_7165,N_7137);
and U7443 (N_7443,N_7132,N_7113);
or U7444 (N_7444,N_7164,N_7084);
or U7445 (N_7445,N_7125,N_7113);
or U7446 (N_7446,N_7039,N_7055);
nand U7447 (N_7447,N_7102,N_7118);
and U7448 (N_7448,N_7085,N_7127);
nor U7449 (N_7449,N_7051,N_7057);
nand U7450 (N_7450,N_7241,N_7113);
nor U7451 (N_7451,N_7212,N_7231);
or U7452 (N_7452,N_7190,N_7042);
or U7453 (N_7453,N_7116,N_7049);
xor U7454 (N_7454,N_7083,N_7163);
and U7455 (N_7455,N_7017,N_7000);
xor U7456 (N_7456,N_7214,N_7073);
and U7457 (N_7457,N_7064,N_7107);
nor U7458 (N_7458,N_7146,N_7112);
or U7459 (N_7459,N_7160,N_7210);
nand U7460 (N_7460,N_7165,N_7016);
nor U7461 (N_7461,N_7054,N_7041);
nor U7462 (N_7462,N_7197,N_7060);
xnor U7463 (N_7463,N_7214,N_7081);
and U7464 (N_7464,N_7163,N_7130);
and U7465 (N_7465,N_7014,N_7156);
or U7466 (N_7466,N_7021,N_7147);
nor U7467 (N_7467,N_7152,N_7050);
nor U7468 (N_7468,N_7025,N_7014);
nand U7469 (N_7469,N_7069,N_7112);
nand U7470 (N_7470,N_7071,N_7012);
nor U7471 (N_7471,N_7098,N_7046);
nand U7472 (N_7472,N_7163,N_7156);
nand U7473 (N_7473,N_7051,N_7017);
and U7474 (N_7474,N_7031,N_7047);
nand U7475 (N_7475,N_7044,N_7023);
nor U7476 (N_7476,N_7213,N_7014);
and U7477 (N_7477,N_7144,N_7179);
xnor U7478 (N_7478,N_7184,N_7200);
and U7479 (N_7479,N_7206,N_7010);
nor U7480 (N_7480,N_7131,N_7112);
nand U7481 (N_7481,N_7012,N_7237);
and U7482 (N_7482,N_7108,N_7149);
or U7483 (N_7483,N_7048,N_7032);
or U7484 (N_7484,N_7175,N_7078);
nor U7485 (N_7485,N_7002,N_7168);
or U7486 (N_7486,N_7242,N_7169);
or U7487 (N_7487,N_7046,N_7146);
nand U7488 (N_7488,N_7166,N_7149);
xor U7489 (N_7489,N_7175,N_7047);
and U7490 (N_7490,N_7105,N_7108);
and U7491 (N_7491,N_7073,N_7176);
and U7492 (N_7492,N_7154,N_7144);
xnor U7493 (N_7493,N_7049,N_7119);
xnor U7494 (N_7494,N_7167,N_7117);
or U7495 (N_7495,N_7116,N_7240);
and U7496 (N_7496,N_7175,N_7153);
and U7497 (N_7497,N_7159,N_7014);
and U7498 (N_7498,N_7122,N_7102);
or U7499 (N_7499,N_7019,N_7063);
nor U7500 (N_7500,N_7311,N_7337);
or U7501 (N_7501,N_7358,N_7443);
or U7502 (N_7502,N_7366,N_7411);
or U7503 (N_7503,N_7302,N_7309);
nand U7504 (N_7504,N_7312,N_7439);
nor U7505 (N_7505,N_7371,N_7424);
or U7506 (N_7506,N_7379,N_7414);
xor U7507 (N_7507,N_7347,N_7380);
and U7508 (N_7508,N_7301,N_7343);
or U7509 (N_7509,N_7332,N_7305);
xor U7510 (N_7510,N_7482,N_7421);
nor U7511 (N_7511,N_7369,N_7429);
nor U7512 (N_7512,N_7474,N_7315);
nand U7513 (N_7513,N_7487,N_7267);
xor U7514 (N_7514,N_7316,N_7419);
or U7515 (N_7515,N_7270,N_7405);
and U7516 (N_7516,N_7460,N_7259);
nor U7517 (N_7517,N_7325,N_7485);
and U7518 (N_7518,N_7255,N_7328);
or U7519 (N_7519,N_7333,N_7265);
and U7520 (N_7520,N_7330,N_7375);
nand U7521 (N_7521,N_7374,N_7351);
xnor U7522 (N_7522,N_7490,N_7364);
nor U7523 (N_7523,N_7495,N_7261);
nor U7524 (N_7524,N_7454,N_7393);
nand U7525 (N_7525,N_7395,N_7258);
and U7526 (N_7526,N_7383,N_7339);
and U7527 (N_7527,N_7481,N_7461);
and U7528 (N_7528,N_7370,N_7403);
nor U7529 (N_7529,N_7420,N_7428);
nor U7530 (N_7530,N_7308,N_7476);
nor U7531 (N_7531,N_7299,N_7350);
nor U7532 (N_7532,N_7404,N_7494);
and U7533 (N_7533,N_7441,N_7277);
xor U7534 (N_7534,N_7321,N_7284);
xnor U7535 (N_7535,N_7372,N_7385);
nand U7536 (N_7536,N_7433,N_7342);
or U7537 (N_7537,N_7322,N_7381);
nand U7538 (N_7538,N_7287,N_7348);
or U7539 (N_7539,N_7323,N_7273);
nand U7540 (N_7540,N_7306,N_7264);
and U7541 (N_7541,N_7295,N_7269);
or U7542 (N_7542,N_7477,N_7257);
nand U7543 (N_7543,N_7300,N_7400);
xnor U7544 (N_7544,N_7462,N_7467);
nor U7545 (N_7545,N_7449,N_7263);
nand U7546 (N_7546,N_7448,N_7480);
nor U7547 (N_7547,N_7445,N_7489);
and U7548 (N_7548,N_7499,N_7418);
or U7549 (N_7549,N_7394,N_7341);
nand U7550 (N_7550,N_7359,N_7458);
xnor U7551 (N_7551,N_7484,N_7304);
xor U7552 (N_7552,N_7314,N_7440);
or U7553 (N_7553,N_7470,N_7392);
nor U7554 (N_7554,N_7252,N_7416);
or U7555 (N_7555,N_7473,N_7361);
nand U7556 (N_7556,N_7457,N_7435);
and U7557 (N_7557,N_7413,N_7486);
nor U7558 (N_7558,N_7260,N_7290);
or U7559 (N_7559,N_7437,N_7283);
and U7560 (N_7560,N_7286,N_7459);
xor U7561 (N_7561,N_7297,N_7384);
and U7562 (N_7562,N_7498,N_7310);
and U7563 (N_7563,N_7422,N_7377);
xor U7564 (N_7564,N_7491,N_7397);
xor U7565 (N_7565,N_7373,N_7389);
and U7566 (N_7566,N_7271,N_7291);
and U7567 (N_7567,N_7417,N_7293);
xor U7568 (N_7568,N_7478,N_7340);
nor U7569 (N_7569,N_7285,N_7453);
nor U7570 (N_7570,N_7298,N_7296);
and U7571 (N_7571,N_7497,N_7390);
or U7572 (N_7572,N_7365,N_7307);
xnor U7573 (N_7573,N_7324,N_7319);
and U7574 (N_7574,N_7472,N_7444);
xnor U7575 (N_7575,N_7426,N_7386);
or U7576 (N_7576,N_7496,N_7320);
nor U7577 (N_7577,N_7434,N_7471);
or U7578 (N_7578,N_7391,N_7274);
xnor U7579 (N_7579,N_7250,N_7408);
nor U7580 (N_7580,N_7430,N_7396);
and U7581 (N_7581,N_7446,N_7292);
and U7582 (N_7582,N_7493,N_7407);
or U7583 (N_7583,N_7349,N_7464);
or U7584 (N_7584,N_7336,N_7327);
xor U7585 (N_7585,N_7398,N_7318);
or U7586 (N_7586,N_7368,N_7388);
and U7587 (N_7587,N_7412,N_7266);
or U7588 (N_7588,N_7363,N_7376);
nor U7589 (N_7589,N_7415,N_7367);
xnor U7590 (N_7590,N_7423,N_7329);
or U7591 (N_7591,N_7427,N_7450);
and U7592 (N_7592,N_7469,N_7256);
or U7593 (N_7593,N_7303,N_7317);
xor U7594 (N_7594,N_7346,N_7278);
or U7595 (N_7595,N_7466,N_7338);
nor U7596 (N_7596,N_7279,N_7378);
nand U7597 (N_7597,N_7475,N_7282);
nor U7598 (N_7598,N_7442,N_7288);
nor U7599 (N_7599,N_7253,N_7354);
nand U7600 (N_7600,N_7488,N_7355);
and U7601 (N_7601,N_7401,N_7331);
xor U7602 (N_7602,N_7438,N_7357);
and U7603 (N_7603,N_7251,N_7352);
and U7604 (N_7604,N_7268,N_7289);
nand U7605 (N_7605,N_7410,N_7272);
nand U7606 (N_7606,N_7463,N_7353);
and U7607 (N_7607,N_7387,N_7468);
or U7608 (N_7608,N_7344,N_7275);
xnor U7609 (N_7609,N_7409,N_7455);
nand U7610 (N_7610,N_7294,N_7313);
and U7611 (N_7611,N_7436,N_7483);
nand U7612 (N_7612,N_7452,N_7425);
xnor U7613 (N_7613,N_7262,N_7382);
nor U7614 (N_7614,N_7402,N_7465);
nor U7615 (N_7615,N_7456,N_7447);
nand U7616 (N_7616,N_7451,N_7431);
nor U7617 (N_7617,N_7280,N_7492);
and U7618 (N_7618,N_7335,N_7362);
and U7619 (N_7619,N_7345,N_7432);
or U7620 (N_7620,N_7326,N_7281);
nand U7621 (N_7621,N_7479,N_7334);
or U7622 (N_7622,N_7399,N_7254);
nand U7623 (N_7623,N_7360,N_7356);
or U7624 (N_7624,N_7406,N_7276);
nor U7625 (N_7625,N_7325,N_7468);
xnor U7626 (N_7626,N_7442,N_7383);
nor U7627 (N_7627,N_7484,N_7355);
nand U7628 (N_7628,N_7261,N_7275);
and U7629 (N_7629,N_7477,N_7326);
nor U7630 (N_7630,N_7349,N_7494);
nand U7631 (N_7631,N_7258,N_7474);
and U7632 (N_7632,N_7352,N_7403);
and U7633 (N_7633,N_7478,N_7463);
or U7634 (N_7634,N_7467,N_7376);
or U7635 (N_7635,N_7432,N_7409);
nand U7636 (N_7636,N_7339,N_7259);
nor U7637 (N_7637,N_7364,N_7375);
nand U7638 (N_7638,N_7402,N_7428);
xor U7639 (N_7639,N_7268,N_7314);
and U7640 (N_7640,N_7286,N_7421);
nand U7641 (N_7641,N_7356,N_7359);
nor U7642 (N_7642,N_7298,N_7443);
nand U7643 (N_7643,N_7454,N_7368);
xnor U7644 (N_7644,N_7456,N_7495);
xor U7645 (N_7645,N_7439,N_7449);
or U7646 (N_7646,N_7463,N_7356);
xor U7647 (N_7647,N_7332,N_7342);
or U7648 (N_7648,N_7383,N_7401);
nor U7649 (N_7649,N_7257,N_7417);
nand U7650 (N_7650,N_7400,N_7475);
and U7651 (N_7651,N_7370,N_7463);
and U7652 (N_7652,N_7348,N_7371);
nand U7653 (N_7653,N_7492,N_7366);
nor U7654 (N_7654,N_7490,N_7254);
xnor U7655 (N_7655,N_7411,N_7267);
xnor U7656 (N_7656,N_7252,N_7263);
nor U7657 (N_7657,N_7324,N_7468);
xnor U7658 (N_7658,N_7433,N_7291);
and U7659 (N_7659,N_7382,N_7323);
and U7660 (N_7660,N_7278,N_7315);
xor U7661 (N_7661,N_7419,N_7300);
and U7662 (N_7662,N_7378,N_7341);
or U7663 (N_7663,N_7367,N_7421);
or U7664 (N_7664,N_7419,N_7370);
and U7665 (N_7665,N_7266,N_7471);
or U7666 (N_7666,N_7396,N_7360);
or U7667 (N_7667,N_7334,N_7308);
or U7668 (N_7668,N_7429,N_7254);
nand U7669 (N_7669,N_7348,N_7434);
or U7670 (N_7670,N_7464,N_7306);
or U7671 (N_7671,N_7388,N_7252);
nand U7672 (N_7672,N_7286,N_7301);
and U7673 (N_7673,N_7276,N_7467);
nor U7674 (N_7674,N_7306,N_7379);
nand U7675 (N_7675,N_7377,N_7385);
nand U7676 (N_7676,N_7453,N_7370);
nor U7677 (N_7677,N_7491,N_7356);
nand U7678 (N_7678,N_7310,N_7333);
nor U7679 (N_7679,N_7419,N_7351);
nand U7680 (N_7680,N_7309,N_7293);
nor U7681 (N_7681,N_7358,N_7390);
nor U7682 (N_7682,N_7295,N_7467);
and U7683 (N_7683,N_7414,N_7282);
nand U7684 (N_7684,N_7344,N_7384);
nor U7685 (N_7685,N_7323,N_7271);
or U7686 (N_7686,N_7312,N_7401);
and U7687 (N_7687,N_7447,N_7358);
or U7688 (N_7688,N_7347,N_7325);
or U7689 (N_7689,N_7334,N_7266);
nand U7690 (N_7690,N_7401,N_7298);
nand U7691 (N_7691,N_7463,N_7364);
xor U7692 (N_7692,N_7287,N_7396);
xor U7693 (N_7693,N_7266,N_7440);
or U7694 (N_7694,N_7377,N_7423);
and U7695 (N_7695,N_7357,N_7362);
nand U7696 (N_7696,N_7399,N_7440);
and U7697 (N_7697,N_7256,N_7333);
and U7698 (N_7698,N_7338,N_7305);
or U7699 (N_7699,N_7401,N_7339);
nor U7700 (N_7700,N_7379,N_7476);
xor U7701 (N_7701,N_7283,N_7478);
and U7702 (N_7702,N_7444,N_7407);
nand U7703 (N_7703,N_7269,N_7462);
xor U7704 (N_7704,N_7318,N_7421);
nor U7705 (N_7705,N_7487,N_7299);
and U7706 (N_7706,N_7345,N_7441);
and U7707 (N_7707,N_7479,N_7261);
nor U7708 (N_7708,N_7276,N_7397);
nand U7709 (N_7709,N_7441,N_7451);
or U7710 (N_7710,N_7496,N_7334);
nor U7711 (N_7711,N_7288,N_7355);
nor U7712 (N_7712,N_7388,N_7461);
xor U7713 (N_7713,N_7461,N_7437);
nand U7714 (N_7714,N_7359,N_7370);
or U7715 (N_7715,N_7493,N_7332);
nor U7716 (N_7716,N_7273,N_7462);
nor U7717 (N_7717,N_7444,N_7464);
nand U7718 (N_7718,N_7476,N_7267);
xnor U7719 (N_7719,N_7306,N_7385);
nor U7720 (N_7720,N_7393,N_7444);
nor U7721 (N_7721,N_7274,N_7253);
nor U7722 (N_7722,N_7371,N_7305);
nand U7723 (N_7723,N_7453,N_7475);
nor U7724 (N_7724,N_7484,N_7322);
or U7725 (N_7725,N_7284,N_7280);
and U7726 (N_7726,N_7498,N_7288);
xnor U7727 (N_7727,N_7311,N_7338);
or U7728 (N_7728,N_7349,N_7270);
nor U7729 (N_7729,N_7499,N_7444);
nor U7730 (N_7730,N_7287,N_7353);
or U7731 (N_7731,N_7274,N_7399);
and U7732 (N_7732,N_7356,N_7371);
or U7733 (N_7733,N_7454,N_7450);
xor U7734 (N_7734,N_7321,N_7494);
xor U7735 (N_7735,N_7309,N_7250);
and U7736 (N_7736,N_7320,N_7290);
and U7737 (N_7737,N_7312,N_7294);
or U7738 (N_7738,N_7375,N_7321);
nor U7739 (N_7739,N_7490,N_7262);
xor U7740 (N_7740,N_7378,N_7299);
nor U7741 (N_7741,N_7269,N_7395);
nor U7742 (N_7742,N_7344,N_7353);
nand U7743 (N_7743,N_7456,N_7488);
or U7744 (N_7744,N_7308,N_7250);
or U7745 (N_7745,N_7278,N_7461);
or U7746 (N_7746,N_7416,N_7296);
and U7747 (N_7747,N_7362,N_7496);
and U7748 (N_7748,N_7321,N_7348);
xor U7749 (N_7749,N_7290,N_7460);
nor U7750 (N_7750,N_7743,N_7739);
xnor U7751 (N_7751,N_7503,N_7535);
and U7752 (N_7752,N_7676,N_7628);
nand U7753 (N_7753,N_7749,N_7515);
nand U7754 (N_7754,N_7579,N_7642);
nor U7755 (N_7755,N_7703,N_7592);
or U7756 (N_7756,N_7625,N_7510);
nand U7757 (N_7757,N_7730,N_7683);
nand U7758 (N_7758,N_7558,N_7685);
nor U7759 (N_7759,N_7721,N_7660);
nand U7760 (N_7760,N_7641,N_7598);
xor U7761 (N_7761,N_7742,N_7626);
nor U7762 (N_7762,N_7618,N_7668);
and U7763 (N_7763,N_7632,N_7543);
or U7764 (N_7764,N_7657,N_7663);
nor U7765 (N_7765,N_7575,N_7562);
xnor U7766 (N_7766,N_7700,N_7634);
nand U7767 (N_7767,N_7741,N_7608);
nand U7768 (N_7768,N_7615,N_7527);
xor U7769 (N_7769,N_7710,N_7720);
and U7770 (N_7770,N_7564,N_7737);
xor U7771 (N_7771,N_7689,N_7692);
and U7772 (N_7772,N_7696,N_7709);
and U7773 (N_7773,N_7655,N_7568);
or U7774 (N_7774,N_7553,N_7607);
and U7775 (N_7775,N_7747,N_7697);
nand U7776 (N_7776,N_7640,N_7500);
nand U7777 (N_7777,N_7744,N_7678);
or U7778 (N_7778,N_7735,N_7551);
and U7779 (N_7779,N_7599,N_7719);
nand U7780 (N_7780,N_7586,N_7534);
nor U7781 (N_7781,N_7629,N_7548);
and U7782 (N_7782,N_7630,N_7684);
and U7783 (N_7783,N_7707,N_7662);
nand U7784 (N_7784,N_7601,N_7605);
nand U7785 (N_7785,N_7603,N_7666);
and U7786 (N_7786,N_7638,N_7648);
nand U7787 (N_7787,N_7585,N_7550);
nor U7788 (N_7788,N_7574,N_7529);
or U7789 (N_7789,N_7519,N_7712);
xor U7790 (N_7790,N_7659,N_7573);
or U7791 (N_7791,N_7522,N_7704);
and U7792 (N_7792,N_7612,N_7542);
nor U7793 (N_7793,N_7509,N_7645);
or U7794 (N_7794,N_7688,N_7544);
nor U7795 (N_7795,N_7524,N_7652);
xor U7796 (N_7796,N_7670,N_7555);
or U7797 (N_7797,N_7595,N_7593);
or U7798 (N_7798,N_7517,N_7520);
and U7799 (N_7799,N_7733,N_7722);
and U7800 (N_7800,N_7694,N_7695);
and U7801 (N_7801,N_7606,N_7647);
xnor U7802 (N_7802,N_7745,N_7578);
and U7803 (N_7803,N_7718,N_7506);
or U7804 (N_7804,N_7563,N_7591);
nor U7805 (N_7805,N_7512,N_7508);
nand U7806 (N_7806,N_7746,N_7633);
xnor U7807 (N_7807,N_7693,N_7674);
xor U7808 (N_7808,N_7594,N_7649);
and U7809 (N_7809,N_7617,N_7729);
and U7810 (N_7810,N_7671,N_7682);
xor U7811 (N_7811,N_7538,N_7636);
xnor U7812 (N_7812,N_7566,N_7673);
or U7813 (N_7813,N_7748,N_7651);
nand U7814 (N_7814,N_7654,N_7569);
or U7815 (N_7815,N_7665,N_7672);
or U7816 (N_7816,N_7717,N_7616);
nand U7817 (N_7817,N_7532,N_7570);
and U7818 (N_7818,N_7699,N_7713);
nor U7819 (N_7819,N_7554,N_7716);
nand U7820 (N_7820,N_7540,N_7646);
or U7821 (N_7821,N_7588,N_7726);
nand U7822 (N_7822,N_7518,N_7583);
and U7823 (N_7823,N_7686,N_7623);
xor U7824 (N_7824,N_7631,N_7576);
or U7825 (N_7825,N_7549,N_7675);
nor U7826 (N_7826,N_7637,N_7581);
xnor U7827 (N_7827,N_7582,N_7546);
xor U7828 (N_7828,N_7664,N_7604);
xor U7829 (N_7829,N_7656,N_7723);
nor U7830 (N_7830,N_7702,N_7537);
or U7831 (N_7831,N_7533,N_7501);
or U7832 (N_7832,N_7528,N_7547);
nand U7833 (N_7833,N_7571,N_7590);
and U7834 (N_7834,N_7653,N_7589);
or U7835 (N_7835,N_7610,N_7513);
xnor U7836 (N_7836,N_7516,N_7627);
or U7837 (N_7837,N_7600,N_7661);
xnor U7838 (N_7838,N_7572,N_7502);
and U7839 (N_7839,N_7622,N_7679);
nand U7840 (N_7840,N_7621,N_7514);
nand U7841 (N_7841,N_7687,N_7715);
nand U7842 (N_7842,N_7511,N_7561);
and U7843 (N_7843,N_7724,N_7650);
or U7844 (N_7844,N_7736,N_7680);
nand U7845 (N_7845,N_7624,N_7677);
nor U7846 (N_7846,N_7740,N_7731);
xor U7847 (N_7847,N_7734,N_7728);
and U7848 (N_7848,N_7557,N_7714);
xor U7849 (N_7849,N_7738,N_7505);
or U7850 (N_7850,N_7577,N_7531);
nor U7851 (N_7851,N_7639,N_7706);
nand U7852 (N_7852,N_7523,N_7565);
nor U7853 (N_7853,N_7560,N_7526);
nor U7854 (N_7854,N_7530,N_7635);
and U7855 (N_7855,N_7556,N_7732);
nand U7856 (N_7856,N_7701,N_7613);
nand U7857 (N_7857,N_7609,N_7507);
or U7858 (N_7858,N_7525,N_7619);
xnor U7859 (N_7859,N_7597,N_7681);
nor U7860 (N_7860,N_7698,N_7691);
nand U7861 (N_7861,N_7545,N_7725);
xor U7862 (N_7862,N_7596,N_7611);
nor U7863 (N_7863,N_7708,N_7587);
xor U7864 (N_7864,N_7552,N_7614);
and U7865 (N_7865,N_7727,N_7690);
or U7866 (N_7866,N_7504,N_7521);
nor U7867 (N_7867,N_7559,N_7580);
and U7868 (N_7868,N_7643,N_7620);
and U7869 (N_7869,N_7567,N_7711);
or U7870 (N_7870,N_7602,N_7644);
or U7871 (N_7871,N_7539,N_7658);
and U7872 (N_7872,N_7536,N_7667);
and U7873 (N_7873,N_7584,N_7541);
or U7874 (N_7874,N_7669,N_7705);
nor U7875 (N_7875,N_7521,N_7709);
and U7876 (N_7876,N_7646,N_7523);
nor U7877 (N_7877,N_7547,N_7627);
nor U7878 (N_7878,N_7690,N_7628);
and U7879 (N_7879,N_7595,N_7653);
xor U7880 (N_7880,N_7543,N_7579);
or U7881 (N_7881,N_7641,N_7604);
and U7882 (N_7882,N_7526,N_7592);
nand U7883 (N_7883,N_7522,N_7574);
or U7884 (N_7884,N_7528,N_7639);
nand U7885 (N_7885,N_7660,N_7702);
and U7886 (N_7886,N_7708,N_7659);
and U7887 (N_7887,N_7701,N_7517);
nor U7888 (N_7888,N_7639,N_7510);
nor U7889 (N_7889,N_7544,N_7502);
or U7890 (N_7890,N_7549,N_7619);
xor U7891 (N_7891,N_7513,N_7644);
xor U7892 (N_7892,N_7558,N_7570);
or U7893 (N_7893,N_7610,N_7552);
and U7894 (N_7894,N_7611,N_7642);
and U7895 (N_7895,N_7619,N_7666);
xnor U7896 (N_7896,N_7724,N_7541);
xor U7897 (N_7897,N_7732,N_7713);
xnor U7898 (N_7898,N_7525,N_7667);
xor U7899 (N_7899,N_7529,N_7638);
nor U7900 (N_7900,N_7500,N_7514);
nand U7901 (N_7901,N_7631,N_7507);
or U7902 (N_7902,N_7677,N_7665);
nor U7903 (N_7903,N_7501,N_7586);
nand U7904 (N_7904,N_7536,N_7505);
or U7905 (N_7905,N_7595,N_7604);
and U7906 (N_7906,N_7645,N_7535);
and U7907 (N_7907,N_7500,N_7718);
nand U7908 (N_7908,N_7553,N_7600);
or U7909 (N_7909,N_7740,N_7674);
nand U7910 (N_7910,N_7679,N_7597);
and U7911 (N_7911,N_7661,N_7641);
nor U7912 (N_7912,N_7693,N_7694);
xor U7913 (N_7913,N_7705,N_7638);
or U7914 (N_7914,N_7615,N_7662);
xnor U7915 (N_7915,N_7607,N_7539);
nor U7916 (N_7916,N_7637,N_7553);
and U7917 (N_7917,N_7665,N_7628);
or U7918 (N_7918,N_7580,N_7639);
xnor U7919 (N_7919,N_7733,N_7602);
xnor U7920 (N_7920,N_7735,N_7647);
nor U7921 (N_7921,N_7676,N_7590);
and U7922 (N_7922,N_7653,N_7503);
xor U7923 (N_7923,N_7559,N_7717);
nor U7924 (N_7924,N_7515,N_7580);
nand U7925 (N_7925,N_7545,N_7544);
nor U7926 (N_7926,N_7576,N_7656);
nand U7927 (N_7927,N_7590,N_7656);
or U7928 (N_7928,N_7716,N_7520);
nand U7929 (N_7929,N_7691,N_7643);
or U7930 (N_7930,N_7645,N_7725);
xnor U7931 (N_7931,N_7741,N_7541);
xor U7932 (N_7932,N_7725,N_7563);
nor U7933 (N_7933,N_7720,N_7633);
xnor U7934 (N_7934,N_7745,N_7527);
nand U7935 (N_7935,N_7609,N_7653);
or U7936 (N_7936,N_7552,N_7690);
nor U7937 (N_7937,N_7682,N_7554);
and U7938 (N_7938,N_7592,N_7573);
nor U7939 (N_7939,N_7603,N_7721);
or U7940 (N_7940,N_7524,N_7702);
nor U7941 (N_7941,N_7515,N_7594);
and U7942 (N_7942,N_7745,N_7541);
and U7943 (N_7943,N_7502,N_7521);
and U7944 (N_7944,N_7513,N_7677);
and U7945 (N_7945,N_7657,N_7527);
xor U7946 (N_7946,N_7685,N_7579);
nand U7947 (N_7947,N_7550,N_7602);
nand U7948 (N_7948,N_7528,N_7506);
xnor U7949 (N_7949,N_7594,N_7711);
xnor U7950 (N_7950,N_7568,N_7699);
nor U7951 (N_7951,N_7702,N_7568);
nor U7952 (N_7952,N_7733,N_7606);
and U7953 (N_7953,N_7628,N_7526);
xor U7954 (N_7954,N_7577,N_7685);
and U7955 (N_7955,N_7605,N_7531);
and U7956 (N_7956,N_7523,N_7586);
and U7957 (N_7957,N_7739,N_7662);
and U7958 (N_7958,N_7508,N_7679);
xor U7959 (N_7959,N_7506,N_7571);
xor U7960 (N_7960,N_7673,N_7714);
xor U7961 (N_7961,N_7542,N_7504);
nand U7962 (N_7962,N_7733,N_7737);
nor U7963 (N_7963,N_7541,N_7704);
xnor U7964 (N_7964,N_7547,N_7692);
and U7965 (N_7965,N_7552,N_7730);
xnor U7966 (N_7966,N_7587,N_7681);
xor U7967 (N_7967,N_7616,N_7736);
xnor U7968 (N_7968,N_7694,N_7594);
and U7969 (N_7969,N_7622,N_7510);
and U7970 (N_7970,N_7720,N_7538);
nand U7971 (N_7971,N_7622,N_7707);
or U7972 (N_7972,N_7641,N_7687);
and U7973 (N_7973,N_7687,N_7633);
or U7974 (N_7974,N_7720,N_7525);
and U7975 (N_7975,N_7560,N_7745);
nor U7976 (N_7976,N_7673,N_7600);
and U7977 (N_7977,N_7545,N_7541);
and U7978 (N_7978,N_7600,N_7593);
nor U7979 (N_7979,N_7627,N_7573);
nand U7980 (N_7980,N_7508,N_7626);
xnor U7981 (N_7981,N_7608,N_7605);
or U7982 (N_7982,N_7519,N_7719);
and U7983 (N_7983,N_7681,N_7541);
nand U7984 (N_7984,N_7683,N_7689);
and U7985 (N_7985,N_7605,N_7545);
or U7986 (N_7986,N_7681,N_7526);
and U7987 (N_7987,N_7590,N_7688);
and U7988 (N_7988,N_7687,N_7660);
or U7989 (N_7989,N_7530,N_7725);
or U7990 (N_7990,N_7634,N_7558);
nor U7991 (N_7991,N_7548,N_7527);
and U7992 (N_7992,N_7512,N_7695);
nand U7993 (N_7993,N_7583,N_7650);
xor U7994 (N_7994,N_7685,N_7731);
nand U7995 (N_7995,N_7725,N_7600);
xor U7996 (N_7996,N_7656,N_7652);
nand U7997 (N_7997,N_7573,N_7654);
xor U7998 (N_7998,N_7552,N_7548);
or U7999 (N_7999,N_7546,N_7665);
xnor U8000 (N_8000,N_7920,N_7984);
nand U8001 (N_8001,N_7971,N_7797);
xnor U8002 (N_8002,N_7995,N_7904);
and U8003 (N_8003,N_7838,N_7852);
and U8004 (N_8004,N_7963,N_7927);
and U8005 (N_8005,N_7799,N_7782);
xor U8006 (N_8006,N_7817,N_7946);
and U8007 (N_8007,N_7805,N_7848);
or U8008 (N_8008,N_7827,N_7931);
xnor U8009 (N_8009,N_7826,N_7874);
xor U8010 (N_8010,N_7895,N_7819);
nand U8011 (N_8011,N_7959,N_7947);
xor U8012 (N_8012,N_7944,N_7899);
nor U8013 (N_8013,N_7915,N_7757);
and U8014 (N_8014,N_7996,N_7754);
nand U8015 (N_8015,N_7810,N_7813);
and U8016 (N_8016,N_7993,N_7935);
xor U8017 (N_8017,N_7869,N_7784);
and U8018 (N_8018,N_7901,N_7778);
or U8019 (N_8019,N_7968,N_7948);
and U8020 (N_8020,N_7942,N_7943);
nand U8021 (N_8021,N_7867,N_7921);
nor U8022 (N_8022,N_7977,N_7870);
or U8023 (N_8023,N_7972,N_7928);
xor U8024 (N_8024,N_7910,N_7879);
nand U8025 (N_8025,N_7860,N_7795);
or U8026 (N_8026,N_7936,N_7866);
nand U8027 (N_8027,N_7938,N_7919);
nor U8028 (N_8028,N_7930,N_7834);
nor U8029 (N_8029,N_7951,N_7856);
and U8030 (N_8030,N_7818,N_7824);
or U8031 (N_8031,N_7969,N_7788);
xnor U8032 (N_8032,N_7922,N_7950);
and U8033 (N_8033,N_7823,N_7850);
xnor U8034 (N_8034,N_7937,N_7786);
xnor U8035 (N_8035,N_7976,N_7815);
or U8036 (N_8036,N_7798,N_7892);
xnor U8037 (N_8037,N_7940,N_7780);
and U8038 (N_8038,N_7851,N_7945);
and U8039 (N_8039,N_7752,N_7883);
xor U8040 (N_8040,N_7796,N_7759);
xnor U8041 (N_8041,N_7794,N_7792);
xnor U8042 (N_8042,N_7967,N_7997);
and U8043 (N_8043,N_7821,N_7884);
nand U8044 (N_8044,N_7756,N_7844);
xor U8045 (N_8045,N_7822,N_7955);
and U8046 (N_8046,N_7987,N_7766);
xnor U8047 (N_8047,N_7916,N_7957);
and U8048 (N_8048,N_7917,N_7808);
or U8049 (N_8049,N_7763,N_7982);
or U8050 (N_8050,N_7983,N_7970);
nor U8051 (N_8051,N_7914,N_7835);
or U8052 (N_8052,N_7900,N_7985);
xnor U8053 (N_8053,N_7839,N_7965);
or U8054 (N_8054,N_7776,N_7924);
and U8055 (N_8055,N_7840,N_7990);
nand U8056 (N_8056,N_7836,N_7772);
nor U8057 (N_8057,N_7961,N_7843);
and U8058 (N_8058,N_7986,N_7888);
or U8059 (N_8059,N_7934,N_7956);
or U8060 (N_8060,N_7979,N_7962);
nor U8061 (N_8061,N_7960,N_7994);
and U8062 (N_8062,N_7767,N_7831);
xnor U8063 (N_8063,N_7768,N_7770);
nand U8064 (N_8064,N_7898,N_7829);
and U8065 (N_8065,N_7769,N_7878);
nor U8066 (N_8066,N_7882,N_7923);
and U8067 (N_8067,N_7872,N_7777);
and U8068 (N_8068,N_7953,N_7855);
nand U8069 (N_8069,N_7903,N_7837);
xnor U8070 (N_8070,N_7758,N_7802);
and U8071 (N_8071,N_7761,N_7876);
nor U8072 (N_8072,N_7893,N_7932);
nand U8073 (N_8073,N_7820,N_7966);
nor U8074 (N_8074,N_7871,N_7809);
nand U8075 (N_8075,N_7849,N_7894);
nand U8076 (N_8076,N_7789,N_7830);
and U8077 (N_8077,N_7787,N_7853);
xnor U8078 (N_8078,N_7861,N_7814);
nor U8079 (N_8079,N_7939,N_7862);
xor U8080 (N_8080,N_7751,N_7816);
or U8081 (N_8081,N_7801,N_7998);
nand U8082 (N_8082,N_7964,N_7864);
or U8083 (N_8083,N_7980,N_7885);
xor U8084 (N_8084,N_7873,N_7750);
nor U8085 (N_8085,N_7886,N_7854);
nor U8086 (N_8086,N_7832,N_7877);
nand U8087 (N_8087,N_7896,N_7791);
or U8088 (N_8088,N_7913,N_7858);
xor U8089 (N_8089,N_7865,N_7989);
xor U8090 (N_8090,N_7775,N_7781);
or U8091 (N_8091,N_7793,N_7905);
xor U8092 (N_8092,N_7753,N_7811);
or U8093 (N_8093,N_7857,N_7806);
nor U8094 (N_8094,N_7887,N_7790);
xnor U8095 (N_8095,N_7890,N_7891);
and U8096 (N_8096,N_7897,N_7842);
and U8097 (N_8097,N_7774,N_7875);
or U8098 (N_8098,N_7912,N_7988);
nor U8099 (N_8099,N_7981,N_7779);
xor U8100 (N_8100,N_7771,N_7847);
nor U8101 (N_8101,N_7803,N_7908);
nor U8102 (N_8102,N_7889,N_7949);
and U8103 (N_8103,N_7906,N_7868);
xnor U8104 (N_8104,N_7846,N_7881);
xor U8105 (N_8105,N_7999,N_7941);
nor U8106 (N_8106,N_7762,N_7929);
nand U8107 (N_8107,N_7975,N_7907);
and U8108 (N_8108,N_7952,N_7760);
and U8109 (N_8109,N_7804,N_7845);
xor U8110 (N_8110,N_7807,N_7833);
or U8111 (N_8111,N_7954,N_7958);
nand U8112 (N_8112,N_7909,N_7828);
or U8113 (N_8113,N_7812,N_7863);
nor U8114 (N_8114,N_7785,N_7859);
xor U8115 (N_8115,N_7825,N_7992);
nor U8116 (N_8116,N_7974,N_7800);
and U8117 (N_8117,N_7902,N_7933);
and U8118 (N_8118,N_7991,N_7926);
nand U8119 (N_8119,N_7841,N_7765);
xnor U8120 (N_8120,N_7773,N_7973);
xnor U8121 (N_8121,N_7783,N_7755);
xnor U8122 (N_8122,N_7978,N_7764);
and U8123 (N_8123,N_7911,N_7925);
nand U8124 (N_8124,N_7880,N_7918);
or U8125 (N_8125,N_7834,N_7912);
nor U8126 (N_8126,N_7948,N_7950);
or U8127 (N_8127,N_7827,N_7895);
nand U8128 (N_8128,N_7826,N_7806);
nand U8129 (N_8129,N_7871,N_7834);
or U8130 (N_8130,N_7983,N_7824);
xor U8131 (N_8131,N_7988,N_7807);
xnor U8132 (N_8132,N_7958,N_7794);
nor U8133 (N_8133,N_7863,N_7836);
xor U8134 (N_8134,N_7883,N_7981);
xor U8135 (N_8135,N_7865,N_7858);
nand U8136 (N_8136,N_7938,N_7756);
nor U8137 (N_8137,N_7969,N_7821);
nand U8138 (N_8138,N_7968,N_7910);
nand U8139 (N_8139,N_7939,N_7988);
xor U8140 (N_8140,N_7765,N_7898);
and U8141 (N_8141,N_7911,N_7813);
nand U8142 (N_8142,N_7800,N_7868);
nand U8143 (N_8143,N_7978,N_7779);
nand U8144 (N_8144,N_7883,N_7894);
or U8145 (N_8145,N_7967,N_7962);
and U8146 (N_8146,N_7862,N_7842);
or U8147 (N_8147,N_7808,N_7779);
nor U8148 (N_8148,N_7881,N_7771);
or U8149 (N_8149,N_7917,N_7871);
nand U8150 (N_8150,N_7996,N_7993);
xnor U8151 (N_8151,N_7758,N_7992);
nor U8152 (N_8152,N_7811,N_7967);
or U8153 (N_8153,N_7994,N_7775);
nand U8154 (N_8154,N_7917,N_7919);
or U8155 (N_8155,N_7915,N_7802);
xor U8156 (N_8156,N_7963,N_7980);
nand U8157 (N_8157,N_7817,N_7848);
nand U8158 (N_8158,N_7807,N_7958);
or U8159 (N_8159,N_7958,N_7762);
nor U8160 (N_8160,N_7786,N_7970);
nor U8161 (N_8161,N_7850,N_7777);
nor U8162 (N_8162,N_7849,N_7756);
nor U8163 (N_8163,N_7904,N_7951);
xor U8164 (N_8164,N_7869,N_7761);
or U8165 (N_8165,N_7779,N_7960);
or U8166 (N_8166,N_7765,N_7903);
and U8167 (N_8167,N_7892,N_7837);
nor U8168 (N_8168,N_7990,N_7775);
nor U8169 (N_8169,N_7974,N_7917);
and U8170 (N_8170,N_7821,N_7781);
and U8171 (N_8171,N_7875,N_7772);
and U8172 (N_8172,N_7984,N_7911);
and U8173 (N_8173,N_7941,N_7814);
nor U8174 (N_8174,N_7940,N_7880);
and U8175 (N_8175,N_7922,N_7820);
xor U8176 (N_8176,N_7985,N_7932);
nand U8177 (N_8177,N_7840,N_7798);
nand U8178 (N_8178,N_7841,N_7833);
nor U8179 (N_8179,N_7928,N_7937);
xor U8180 (N_8180,N_7865,N_7823);
xnor U8181 (N_8181,N_7828,N_7770);
xor U8182 (N_8182,N_7904,N_7981);
nand U8183 (N_8183,N_7778,N_7819);
or U8184 (N_8184,N_7922,N_7814);
or U8185 (N_8185,N_7926,N_7895);
and U8186 (N_8186,N_7957,N_7915);
nor U8187 (N_8187,N_7751,N_7833);
or U8188 (N_8188,N_7869,N_7939);
and U8189 (N_8189,N_7819,N_7773);
nor U8190 (N_8190,N_7943,N_7787);
or U8191 (N_8191,N_7935,N_7833);
or U8192 (N_8192,N_7887,N_7966);
or U8193 (N_8193,N_7992,N_7999);
nand U8194 (N_8194,N_7961,N_7905);
or U8195 (N_8195,N_7751,N_7873);
nor U8196 (N_8196,N_7817,N_7950);
nor U8197 (N_8197,N_7828,N_7879);
xor U8198 (N_8198,N_7904,N_7973);
and U8199 (N_8199,N_7793,N_7947);
or U8200 (N_8200,N_7940,N_7978);
or U8201 (N_8201,N_7897,N_7992);
and U8202 (N_8202,N_7755,N_7995);
or U8203 (N_8203,N_7934,N_7816);
nor U8204 (N_8204,N_7995,N_7834);
xnor U8205 (N_8205,N_7984,N_7819);
and U8206 (N_8206,N_7900,N_7853);
and U8207 (N_8207,N_7976,N_7886);
nand U8208 (N_8208,N_7942,N_7858);
or U8209 (N_8209,N_7909,N_7801);
xnor U8210 (N_8210,N_7844,N_7905);
nand U8211 (N_8211,N_7887,N_7841);
and U8212 (N_8212,N_7940,N_7917);
xor U8213 (N_8213,N_7870,N_7764);
nand U8214 (N_8214,N_7817,N_7796);
nor U8215 (N_8215,N_7888,N_7868);
or U8216 (N_8216,N_7894,N_7756);
xnor U8217 (N_8217,N_7825,N_7834);
or U8218 (N_8218,N_7831,N_7900);
and U8219 (N_8219,N_7961,N_7753);
nand U8220 (N_8220,N_7927,N_7976);
xnor U8221 (N_8221,N_7898,N_7937);
nand U8222 (N_8222,N_7936,N_7879);
nor U8223 (N_8223,N_7833,N_7782);
and U8224 (N_8224,N_7757,N_7806);
xor U8225 (N_8225,N_7794,N_7848);
nor U8226 (N_8226,N_7775,N_7932);
xnor U8227 (N_8227,N_7877,N_7980);
nor U8228 (N_8228,N_7829,N_7934);
nor U8229 (N_8229,N_7786,N_7802);
xor U8230 (N_8230,N_7836,N_7887);
nand U8231 (N_8231,N_7895,N_7917);
nand U8232 (N_8232,N_7787,N_7931);
nor U8233 (N_8233,N_7782,N_7911);
and U8234 (N_8234,N_7804,N_7772);
and U8235 (N_8235,N_7789,N_7980);
xnor U8236 (N_8236,N_7937,N_7953);
or U8237 (N_8237,N_7827,N_7885);
or U8238 (N_8238,N_7779,N_7950);
xnor U8239 (N_8239,N_7996,N_7853);
and U8240 (N_8240,N_7828,N_7923);
or U8241 (N_8241,N_7795,N_7919);
nor U8242 (N_8242,N_7831,N_7998);
xnor U8243 (N_8243,N_7814,N_7955);
and U8244 (N_8244,N_7750,N_7875);
nor U8245 (N_8245,N_7752,N_7834);
nor U8246 (N_8246,N_7894,N_7779);
nand U8247 (N_8247,N_7937,N_7842);
nand U8248 (N_8248,N_7803,N_7882);
nor U8249 (N_8249,N_7760,N_7836);
nor U8250 (N_8250,N_8056,N_8162);
nand U8251 (N_8251,N_8188,N_8227);
nor U8252 (N_8252,N_8004,N_8055);
or U8253 (N_8253,N_8212,N_8131);
and U8254 (N_8254,N_8034,N_8161);
nor U8255 (N_8255,N_8017,N_8201);
and U8256 (N_8256,N_8070,N_8148);
or U8257 (N_8257,N_8177,N_8094);
and U8258 (N_8258,N_8120,N_8075);
and U8259 (N_8259,N_8150,N_8208);
xor U8260 (N_8260,N_8012,N_8052);
and U8261 (N_8261,N_8025,N_8013);
nand U8262 (N_8262,N_8061,N_8091);
nand U8263 (N_8263,N_8112,N_8098);
and U8264 (N_8264,N_8171,N_8099);
nor U8265 (N_8265,N_8092,N_8138);
nor U8266 (N_8266,N_8141,N_8249);
nand U8267 (N_8267,N_8226,N_8168);
xnor U8268 (N_8268,N_8031,N_8118);
nand U8269 (N_8269,N_8030,N_8183);
and U8270 (N_8270,N_8076,N_8153);
nand U8271 (N_8271,N_8239,N_8026);
nor U8272 (N_8272,N_8237,N_8119);
or U8273 (N_8273,N_8081,N_8245);
nor U8274 (N_8274,N_8065,N_8116);
or U8275 (N_8275,N_8202,N_8020);
and U8276 (N_8276,N_8014,N_8068);
nor U8277 (N_8277,N_8104,N_8213);
and U8278 (N_8278,N_8051,N_8022);
or U8279 (N_8279,N_8189,N_8028);
xnor U8280 (N_8280,N_8069,N_8160);
nor U8281 (N_8281,N_8199,N_8163);
nand U8282 (N_8282,N_8105,N_8181);
xor U8283 (N_8283,N_8100,N_8097);
nand U8284 (N_8284,N_8035,N_8193);
nand U8285 (N_8285,N_8067,N_8146);
nor U8286 (N_8286,N_8126,N_8063);
and U8287 (N_8287,N_8205,N_8073);
xor U8288 (N_8288,N_8191,N_8077);
and U8289 (N_8289,N_8049,N_8132);
nand U8290 (N_8290,N_8064,N_8087);
or U8291 (N_8291,N_8142,N_8178);
xnor U8292 (N_8292,N_8241,N_8231);
and U8293 (N_8293,N_8102,N_8174);
xnor U8294 (N_8294,N_8050,N_8190);
nor U8295 (N_8295,N_8210,N_8176);
or U8296 (N_8296,N_8243,N_8164);
nor U8297 (N_8297,N_8042,N_8027);
or U8298 (N_8298,N_8007,N_8223);
and U8299 (N_8299,N_8115,N_8235);
xor U8300 (N_8300,N_8085,N_8127);
nor U8301 (N_8301,N_8018,N_8179);
or U8302 (N_8302,N_8159,N_8152);
nor U8303 (N_8303,N_8072,N_8185);
nand U8304 (N_8304,N_8078,N_8023);
xor U8305 (N_8305,N_8157,N_8229);
or U8306 (N_8306,N_8090,N_8140);
xnor U8307 (N_8307,N_8122,N_8167);
or U8308 (N_8308,N_8003,N_8211);
or U8309 (N_8309,N_8151,N_8145);
or U8310 (N_8310,N_8124,N_8033);
nand U8311 (N_8311,N_8123,N_8107);
nor U8312 (N_8312,N_8121,N_8209);
or U8313 (N_8313,N_8173,N_8047);
or U8314 (N_8314,N_8144,N_8165);
nand U8315 (N_8315,N_8010,N_8019);
and U8316 (N_8316,N_8108,N_8093);
and U8317 (N_8317,N_8101,N_8040);
xnor U8318 (N_8318,N_8198,N_8242);
or U8319 (N_8319,N_8113,N_8222);
nand U8320 (N_8320,N_8032,N_8006);
xnor U8321 (N_8321,N_8001,N_8045);
xnor U8322 (N_8322,N_8224,N_8207);
nor U8323 (N_8323,N_8036,N_8156);
and U8324 (N_8324,N_8039,N_8232);
nor U8325 (N_8325,N_8238,N_8247);
and U8326 (N_8326,N_8082,N_8021);
xnor U8327 (N_8327,N_8220,N_8037);
or U8328 (N_8328,N_8194,N_8109);
xnor U8329 (N_8329,N_8096,N_8154);
and U8330 (N_8330,N_8192,N_8057);
nand U8331 (N_8331,N_8244,N_8139);
nand U8332 (N_8332,N_8197,N_8136);
xor U8333 (N_8333,N_8130,N_8015);
or U8334 (N_8334,N_8129,N_8060);
or U8335 (N_8335,N_8103,N_8074);
nand U8336 (N_8336,N_8083,N_8187);
or U8337 (N_8337,N_8029,N_8079);
and U8338 (N_8338,N_8230,N_8240);
and U8339 (N_8339,N_8114,N_8180);
nand U8340 (N_8340,N_8110,N_8038);
nor U8341 (N_8341,N_8184,N_8149);
nand U8342 (N_8342,N_8236,N_8204);
xor U8343 (N_8343,N_8246,N_8200);
and U8344 (N_8344,N_8158,N_8002);
and U8345 (N_8345,N_8084,N_8111);
and U8346 (N_8346,N_8228,N_8134);
nor U8347 (N_8347,N_8170,N_8182);
and U8348 (N_8348,N_8217,N_8024);
and U8349 (N_8349,N_8233,N_8058);
and U8350 (N_8350,N_8137,N_8066);
nand U8351 (N_8351,N_8218,N_8216);
and U8352 (N_8352,N_8234,N_8155);
or U8353 (N_8353,N_8041,N_8080);
nand U8354 (N_8354,N_8172,N_8044);
nor U8355 (N_8355,N_8143,N_8059);
nor U8356 (N_8356,N_8117,N_8166);
nand U8357 (N_8357,N_8175,N_8048);
nand U8358 (N_8358,N_8225,N_8054);
nor U8359 (N_8359,N_8106,N_8008);
xor U8360 (N_8360,N_8071,N_8089);
or U8361 (N_8361,N_8043,N_8214);
xor U8362 (N_8362,N_8046,N_8169);
nor U8363 (N_8363,N_8221,N_8095);
and U8364 (N_8364,N_8186,N_8196);
xor U8365 (N_8365,N_8133,N_8147);
xnor U8366 (N_8366,N_8128,N_8088);
or U8367 (N_8367,N_8248,N_8011);
nor U8368 (N_8368,N_8215,N_8195);
and U8369 (N_8369,N_8086,N_8005);
nor U8370 (N_8370,N_8219,N_8053);
nor U8371 (N_8371,N_8135,N_8062);
and U8372 (N_8372,N_8000,N_8009);
nor U8373 (N_8373,N_8206,N_8203);
and U8374 (N_8374,N_8125,N_8016);
xnor U8375 (N_8375,N_8118,N_8064);
and U8376 (N_8376,N_8004,N_8203);
xor U8377 (N_8377,N_8167,N_8013);
xor U8378 (N_8378,N_8100,N_8113);
or U8379 (N_8379,N_8134,N_8166);
xnor U8380 (N_8380,N_8233,N_8104);
nor U8381 (N_8381,N_8215,N_8091);
and U8382 (N_8382,N_8063,N_8119);
xnor U8383 (N_8383,N_8229,N_8077);
nand U8384 (N_8384,N_8169,N_8041);
nor U8385 (N_8385,N_8247,N_8072);
or U8386 (N_8386,N_8247,N_8199);
and U8387 (N_8387,N_8244,N_8145);
nor U8388 (N_8388,N_8212,N_8232);
nor U8389 (N_8389,N_8099,N_8142);
nand U8390 (N_8390,N_8044,N_8043);
xor U8391 (N_8391,N_8035,N_8223);
xor U8392 (N_8392,N_8190,N_8051);
nor U8393 (N_8393,N_8066,N_8146);
nand U8394 (N_8394,N_8017,N_8040);
or U8395 (N_8395,N_8242,N_8230);
or U8396 (N_8396,N_8063,N_8194);
nor U8397 (N_8397,N_8186,N_8088);
nor U8398 (N_8398,N_8151,N_8103);
xor U8399 (N_8399,N_8132,N_8226);
and U8400 (N_8400,N_8018,N_8120);
nor U8401 (N_8401,N_8105,N_8223);
xor U8402 (N_8402,N_8102,N_8186);
xnor U8403 (N_8403,N_8170,N_8117);
xnor U8404 (N_8404,N_8193,N_8094);
nor U8405 (N_8405,N_8168,N_8140);
and U8406 (N_8406,N_8138,N_8176);
xnor U8407 (N_8407,N_8152,N_8157);
nor U8408 (N_8408,N_8029,N_8128);
nor U8409 (N_8409,N_8218,N_8240);
or U8410 (N_8410,N_8093,N_8243);
or U8411 (N_8411,N_8091,N_8207);
nor U8412 (N_8412,N_8235,N_8010);
nand U8413 (N_8413,N_8086,N_8117);
xor U8414 (N_8414,N_8015,N_8082);
and U8415 (N_8415,N_8234,N_8004);
and U8416 (N_8416,N_8098,N_8100);
xor U8417 (N_8417,N_8245,N_8114);
and U8418 (N_8418,N_8139,N_8206);
xnor U8419 (N_8419,N_8242,N_8036);
nor U8420 (N_8420,N_8242,N_8030);
or U8421 (N_8421,N_8172,N_8062);
xnor U8422 (N_8422,N_8104,N_8076);
xnor U8423 (N_8423,N_8113,N_8115);
nand U8424 (N_8424,N_8015,N_8122);
nor U8425 (N_8425,N_8201,N_8138);
and U8426 (N_8426,N_8205,N_8051);
xor U8427 (N_8427,N_8098,N_8051);
or U8428 (N_8428,N_8152,N_8188);
nand U8429 (N_8429,N_8039,N_8234);
xor U8430 (N_8430,N_8032,N_8005);
nand U8431 (N_8431,N_8011,N_8200);
nor U8432 (N_8432,N_8139,N_8062);
nand U8433 (N_8433,N_8000,N_8197);
and U8434 (N_8434,N_8081,N_8225);
nor U8435 (N_8435,N_8092,N_8015);
xnor U8436 (N_8436,N_8073,N_8237);
xnor U8437 (N_8437,N_8107,N_8051);
or U8438 (N_8438,N_8151,N_8071);
nand U8439 (N_8439,N_8206,N_8196);
xnor U8440 (N_8440,N_8166,N_8193);
nor U8441 (N_8441,N_8140,N_8245);
xor U8442 (N_8442,N_8018,N_8136);
and U8443 (N_8443,N_8038,N_8055);
nor U8444 (N_8444,N_8016,N_8061);
or U8445 (N_8445,N_8121,N_8206);
nor U8446 (N_8446,N_8215,N_8221);
nand U8447 (N_8447,N_8230,N_8090);
and U8448 (N_8448,N_8055,N_8220);
and U8449 (N_8449,N_8204,N_8033);
and U8450 (N_8450,N_8161,N_8234);
nor U8451 (N_8451,N_8100,N_8048);
or U8452 (N_8452,N_8240,N_8098);
or U8453 (N_8453,N_8223,N_8156);
or U8454 (N_8454,N_8105,N_8045);
nand U8455 (N_8455,N_8183,N_8058);
nor U8456 (N_8456,N_8144,N_8247);
nand U8457 (N_8457,N_8237,N_8060);
nor U8458 (N_8458,N_8154,N_8081);
and U8459 (N_8459,N_8010,N_8240);
nand U8460 (N_8460,N_8062,N_8094);
and U8461 (N_8461,N_8096,N_8118);
nand U8462 (N_8462,N_8133,N_8123);
nor U8463 (N_8463,N_8142,N_8214);
xnor U8464 (N_8464,N_8163,N_8248);
nor U8465 (N_8465,N_8180,N_8187);
or U8466 (N_8466,N_8138,N_8061);
or U8467 (N_8467,N_8134,N_8167);
nor U8468 (N_8468,N_8204,N_8029);
xnor U8469 (N_8469,N_8210,N_8193);
and U8470 (N_8470,N_8106,N_8209);
nand U8471 (N_8471,N_8032,N_8186);
nand U8472 (N_8472,N_8158,N_8065);
nand U8473 (N_8473,N_8084,N_8060);
or U8474 (N_8474,N_8243,N_8007);
and U8475 (N_8475,N_8233,N_8025);
or U8476 (N_8476,N_8219,N_8086);
xnor U8477 (N_8477,N_8077,N_8111);
and U8478 (N_8478,N_8070,N_8237);
and U8479 (N_8479,N_8127,N_8021);
xnor U8480 (N_8480,N_8221,N_8050);
xnor U8481 (N_8481,N_8209,N_8176);
xor U8482 (N_8482,N_8187,N_8206);
and U8483 (N_8483,N_8031,N_8075);
and U8484 (N_8484,N_8245,N_8214);
and U8485 (N_8485,N_8104,N_8240);
xor U8486 (N_8486,N_8012,N_8137);
or U8487 (N_8487,N_8225,N_8224);
nor U8488 (N_8488,N_8046,N_8038);
or U8489 (N_8489,N_8152,N_8056);
nand U8490 (N_8490,N_8057,N_8233);
xnor U8491 (N_8491,N_8131,N_8007);
or U8492 (N_8492,N_8229,N_8191);
nand U8493 (N_8493,N_8011,N_8095);
nand U8494 (N_8494,N_8088,N_8009);
xnor U8495 (N_8495,N_8188,N_8157);
nor U8496 (N_8496,N_8004,N_8029);
xnor U8497 (N_8497,N_8160,N_8112);
and U8498 (N_8498,N_8064,N_8169);
nor U8499 (N_8499,N_8214,N_8058);
and U8500 (N_8500,N_8274,N_8401);
or U8501 (N_8501,N_8341,N_8366);
nand U8502 (N_8502,N_8315,N_8310);
or U8503 (N_8503,N_8432,N_8270);
and U8504 (N_8504,N_8464,N_8252);
or U8505 (N_8505,N_8426,N_8457);
nor U8506 (N_8506,N_8290,N_8284);
xor U8507 (N_8507,N_8415,N_8324);
nor U8508 (N_8508,N_8445,N_8463);
and U8509 (N_8509,N_8363,N_8295);
and U8510 (N_8510,N_8377,N_8361);
or U8511 (N_8511,N_8471,N_8384);
xor U8512 (N_8512,N_8387,N_8326);
and U8513 (N_8513,N_8344,N_8298);
and U8514 (N_8514,N_8333,N_8468);
or U8515 (N_8515,N_8487,N_8360);
nor U8516 (N_8516,N_8425,N_8305);
and U8517 (N_8517,N_8261,N_8408);
nand U8518 (N_8518,N_8480,N_8265);
xor U8519 (N_8519,N_8260,N_8450);
xnor U8520 (N_8520,N_8424,N_8482);
nor U8521 (N_8521,N_8257,N_8452);
or U8522 (N_8522,N_8357,N_8379);
nand U8523 (N_8523,N_8419,N_8352);
nand U8524 (N_8524,N_8410,N_8402);
nor U8525 (N_8525,N_8416,N_8411);
xor U8526 (N_8526,N_8393,N_8264);
and U8527 (N_8527,N_8400,N_8335);
xnor U8528 (N_8528,N_8435,N_8311);
nor U8529 (N_8529,N_8291,N_8369);
and U8530 (N_8530,N_8349,N_8476);
nand U8531 (N_8531,N_8413,N_8281);
nand U8532 (N_8532,N_8456,N_8403);
nand U8533 (N_8533,N_8323,N_8484);
or U8534 (N_8534,N_8370,N_8296);
xnor U8535 (N_8535,N_8478,N_8461);
or U8536 (N_8536,N_8327,N_8446);
and U8537 (N_8537,N_8294,N_8286);
nand U8538 (N_8538,N_8331,N_8497);
nand U8539 (N_8539,N_8440,N_8443);
xnor U8540 (N_8540,N_8371,N_8477);
xnor U8541 (N_8541,N_8434,N_8320);
nand U8542 (N_8542,N_8255,N_8263);
nand U8543 (N_8543,N_8251,N_8302);
and U8544 (N_8544,N_8469,N_8351);
or U8545 (N_8545,N_8303,N_8322);
xor U8546 (N_8546,N_8498,N_8427);
xnor U8547 (N_8547,N_8423,N_8297);
or U8548 (N_8548,N_8447,N_8373);
xor U8549 (N_8549,N_8312,N_8466);
xor U8550 (N_8550,N_8438,N_8495);
or U8551 (N_8551,N_8431,N_8396);
and U8552 (N_8552,N_8307,N_8499);
nor U8553 (N_8553,N_8382,N_8383);
or U8554 (N_8554,N_8490,N_8436);
or U8555 (N_8555,N_8395,N_8472);
nand U8556 (N_8556,N_8346,N_8405);
or U8557 (N_8557,N_8451,N_8325);
nand U8558 (N_8558,N_8406,N_8299);
nor U8559 (N_8559,N_8422,N_8287);
or U8560 (N_8560,N_8429,N_8467);
nor U8561 (N_8561,N_8407,N_8386);
nand U8562 (N_8562,N_8288,N_8420);
nor U8563 (N_8563,N_8283,N_8278);
nor U8564 (N_8564,N_8353,N_8367);
xor U8565 (N_8565,N_8273,N_8459);
nand U8566 (N_8566,N_8272,N_8345);
nand U8567 (N_8567,N_8259,N_8317);
or U8568 (N_8568,N_8398,N_8391);
nor U8569 (N_8569,N_8362,N_8330);
or U8570 (N_8570,N_8271,N_8489);
nor U8571 (N_8571,N_8375,N_8376);
nand U8572 (N_8572,N_8474,N_8439);
and U8573 (N_8573,N_8314,N_8268);
and U8574 (N_8574,N_8300,N_8359);
xnor U8575 (N_8575,N_8355,N_8313);
nand U8576 (N_8576,N_8350,N_8292);
or U8577 (N_8577,N_8348,N_8347);
and U8578 (N_8578,N_8491,N_8448);
nand U8579 (N_8579,N_8358,N_8421);
nand U8580 (N_8580,N_8412,N_8365);
nor U8581 (N_8581,N_8397,N_8392);
and U8582 (N_8582,N_8262,N_8343);
or U8583 (N_8583,N_8492,N_8342);
xnor U8584 (N_8584,N_8318,N_8319);
nor U8585 (N_8585,N_8337,N_8496);
nand U8586 (N_8586,N_8404,N_8304);
nor U8587 (N_8587,N_8455,N_8453);
xnor U8588 (N_8588,N_8309,N_8414);
xor U8589 (N_8589,N_8485,N_8254);
nand U8590 (N_8590,N_8329,N_8428);
or U8591 (N_8591,N_8266,N_8444);
xnor U8592 (N_8592,N_8275,N_8293);
nor U8593 (N_8593,N_8364,N_8479);
and U8594 (N_8594,N_8399,N_8418);
nand U8595 (N_8595,N_8289,N_8483);
nand U8596 (N_8596,N_8460,N_8385);
or U8597 (N_8597,N_8256,N_8258);
and U8598 (N_8598,N_8354,N_8473);
xnor U8599 (N_8599,N_8332,N_8437);
nor U8600 (N_8600,N_8417,N_8475);
nor U8601 (N_8601,N_8285,N_8306);
nand U8602 (N_8602,N_8470,N_8308);
and U8603 (N_8603,N_8388,N_8253);
nand U8604 (N_8604,N_8338,N_8394);
nor U8605 (N_8605,N_8339,N_8465);
nor U8606 (N_8606,N_8481,N_8336);
and U8607 (N_8607,N_8321,N_8279);
nand U8608 (N_8608,N_8493,N_8390);
xor U8609 (N_8609,N_8454,N_8494);
xor U8610 (N_8610,N_8462,N_8301);
xor U8611 (N_8611,N_8277,N_8316);
and U8612 (N_8612,N_8250,N_8441);
xnor U8613 (N_8613,N_8409,N_8328);
nand U8614 (N_8614,N_8449,N_8372);
nor U8615 (N_8615,N_8433,N_8356);
nor U8616 (N_8616,N_8280,N_8389);
nor U8617 (N_8617,N_8282,N_8442);
and U8618 (N_8618,N_8380,N_8267);
nand U8619 (N_8619,N_8368,N_8378);
and U8620 (N_8620,N_8374,N_8488);
nand U8621 (N_8621,N_8340,N_8276);
nand U8622 (N_8622,N_8381,N_8334);
xnor U8623 (N_8623,N_8458,N_8486);
nor U8624 (N_8624,N_8430,N_8269);
nor U8625 (N_8625,N_8292,N_8263);
nor U8626 (N_8626,N_8373,N_8455);
or U8627 (N_8627,N_8403,N_8407);
or U8628 (N_8628,N_8472,N_8294);
and U8629 (N_8629,N_8446,N_8365);
nand U8630 (N_8630,N_8487,N_8293);
or U8631 (N_8631,N_8268,N_8482);
or U8632 (N_8632,N_8288,N_8275);
xnor U8633 (N_8633,N_8492,N_8441);
xnor U8634 (N_8634,N_8377,N_8426);
and U8635 (N_8635,N_8422,N_8353);
or U8636 (N_8636,N_8275,N_8491);
nand U8637 (N_8637,N_8362,N_8472);
nor U8638 (N_8638,N_8407,N_8367);
xor U8639 (N_8639,N_8284,N_8408);
nor U8640 (N_8640,N_8487,N_8250);
nand U8641 (N_8641,N_8384,N_8267);
nand U8642 (N_8642,N_8414,N_8331);
nand U8643 (N_8643,N_8303,N_8285);
nor U8644 (N_8644,N_8284,N_8482);
xnor U8645 (N_8645,N_8298,N_8402);
nand U8646 (N_8646,N_8252,N_8354);
nor U8647 (N_8647,N_8459,N_8264);
and U8648 (N_8648,N_8284,N_8467);
or U8649 (N_8649,N_8479,N_8354);
xor U8650 (N_8650,N_8305,N_8422);
or U8651 (N_8651,N_8424,N_8332);
and U8652 (N_8652,N_8381,N_8455);
or U8653 (N_8653,N_8479,N_8340);
or U8654 (N_8654,N_8387,N_8472);
nor U8655 (N_8655,N_8494,N_8372);
xnor U8656 (N_8656,N_8299,N_8396);
or U8657 (N_8657,N_8464,N_8402);
and U8658 (N_8658,N_8410,N_8326);
or U8659 (N_8659,N_8285,N_8372);
and U8660 (N_8660,N_8397,N_8409);
or U8661 (N_8661,N_8464,N_8310);
and U8662 (N_8662,N_8321,N_8435);
nand U8663 (N_8663,N_8353,N_8410);
nand U8664 (N_8664,N_8476,N_8315);
and U8665 (N_8665,N_8330,N_8464);
nand U8666 (N_8666,N_8295,N_8429);
xor U8667 (N_8667,N_8329,N_8495);
nand U8668 (N_8668,N_8445,N_8390);
nor U8669 (N_8669,N_8411,N_8454);
xor U8670 (N_8670,N_8267,N_8332);
or U8671 (N_8671,N_8355,N_8374);
or U8672 (N_8672,N_8451,N_8480);
or U8673 (N_8673,N_8457,N_8497);
or U8674 (N_8674,N_8425,N_8457);
nand U8675 (N_8675,N_8264,N_8470);
nand U8676 (N_8676,N_8492,N_8309);
xor U8677 (N_8677,N_8488,N_8423);
or U8678 (N_8678,N_8288,N_8470);
and U8679 (N_8679,N_8484,N_8410);
nand U8680 (N_8680,N_8354,N_8293);
nor U8681 (N_8681,N_8378,N_8476);
and U8682 (N_8682,N_8272,N_8316);
or U8683 (N_8683,N_8273,N_8447);
or U8684 (N_8684,N_8270,N_8386);
and U8685 (N_8685,N_8413,N_8250);
and U8686 (N_8686,N_8473,N_8399);
or U8687 (N_8687,N_8427,N_8457);
nor U8688 (N_8688,N_8263,N_8332);
nand U8689 (N_8689,N_8462,N_8281);
nor U8690 (N_8690,N_8454,N_8268);
xnor U8691 (N_8691,N_8347,N_8439);
or U8692 (N_8692,N_8345,N_8361);
or U8693 (N_8693,N_8263,N_8377);
nand U8694 (N_8694,N_8480,N_8302);
nand U8695 (N_8695,N_8492,N_8426);
and U8696 (N_8696,N_8495,N_8312);
nand U8697 (N_8697,N_8455,N_8260);
or U8698 (N_8698,N_8470,N_8305);
nand U8699 (N_8699,N_8465,N_8464);
xor U8700 (N_8700,N_8424,N_8430);
or U8701 (N_8701,N_8288,N_8358);
and U8702 (N_8702,N_8476,N_8422);
nand U8703 (N_8703,N_8316,N_8423);
nor U8704 (N_8704,N_8285,N_8431);
and U8705 (N_8705,N_8499,N_8389);
nand U8706 (N_8706,N_8447,N_8453);
xor U8707 (N_8707,N_8487,N_8440);
or U8708 (N_8708,N_8254,N_8264);
nor U8709 (N_8709,N_8416,N_8253);
xor U8710 (N_8710,N_8377,N_8414);
and U8711 (N_8711,N_8418,N_8305);
nand U8712 (N_8712,N_8430,N_8354);
nor U8713 (N_8713,N_8428,N_8268);
and U8714 (N_8714,N_8301,N_8300);
or U8715 (N_8715,N_8402,N_8472);
and U8716 (N_8716,N_8272,N_8480);
or U8717 (N_8717,N_8464,N_8416);
or U8718 (N_8718,N_8270,N_8260);
nor U8719 (N_8719,N_8362,N_8296);
and U8720 (N_8720,N_8351,N_8390);
or U8721 (N_8721,N_8288,N_8464);
and U8722 (N_8722,N_8394,N_8362);
xnor U8723 (N_8723,N_8401,N_8443);
nor U8724 (N_8724,N_8301,N_8358);
or U8725 (N_8725,N_8424,N_8445);
nor U8726 (N_8726,N_8391,N_8264);
nand U8727 (N_8727,N_8425,N_8315);
or U8728 (N_8728,N_8349,N_8435);
nand U8729 (N_8729,N_8331,N_8304);
or U8730 (N_8730,N_8267,N_8383);
nor U8731 (N_8731,N_8290,N_8348);
nand U8732 (N_8732,N_8383,N_8298);
xnor U8733 (N_8733,N_8471,N_8268);
xnor U8734 (N_8734,N_8403,N_8452);
or U8735 (N_8735,N_8338,N_8392);
and U8736 (N_8736,N_8351,N_8472);
xnor U8737 (N_8737,N_8356,N_8492);
or U8738 (N_8738,N_8288,N_8399);
xor U8739 (N_8739,N_8399,N_8453);
or U8740 (N_8740,N_8338,N_8292);
or U8741 (N_8741,N_8316,N_8324);
and U8742 (N_8742,N_8327,N_8331);
xor U8743 (N_8743,N_8303,N_8364);
nor U8744 (N_8744,N_8405,N_8293);
xnor U8745 (N_8745,N_8497,N_8358);
and U8746 (N_8746,N_8281,N_8374);
nand U8747 (N_8747,N_8453,N_8311);
nand U8748 (N_8748,N_8487,N_8423);
or U8749 (N_8749,N_8391,N_8282);
nor U8750 (N_8750,N_8693,N_8675);
xor U8751 (N_8751,N_8612,N_8606);
and U8752 (N_8752,N_8609,N_8709);
xor U8753 (N_8753,N_8558,N_8569);
and U8754 (N_8754,N_8594,N_8692);
or U8755 (N_8755,N_8573,N_8661);
or U8756 (N_8756,N_8629,N_8551);
nand U8757 (N_8757,N_8716,N_8616);
xor U8758 (N_8758,N_8550,N_8581);
nor U8759 (N_8759,N_8740,N_8619);
and U8760 (N_8760,N_8677,N_8605);
nor U8761 (N_8761,N_8528,N_8523);
nand U8762 (N_8762,N_8583,N_8665);
xor U8763 (N_8763,N_8598,N_8597);
or U8764 (N_8764,N_8721,N_8688);
or U8765 (N_8765,N_8504,N_8570);
or U8766 (N_8766,N_8733,N_8516);
nor U8767 (N_8767,N_8503,N_8541);
nor U8768 (N_8768,N_8711,N_8727);
and U8769 (N_8769,N_8662,N_8640);
or U8770 (N_8770,N_8634,N_8552);
and U8771 (N_8771,N_8588,N_8670);
xnor U8772 (N_8772,N_8572,N_8526);
and U8773 (N_8773,N_8561,N_8617);
and U8774 (N_8774,N_8663,N_8743);
xnor U8775 (N_8775,N_8580,N_8600);
nand U8776 (N_8776,N_8669,N_8610);
and U8777 (N_8777,N_8546,N_8672);
or U8778 (N_8778,N_8547,N_8529);
or U8779 (N_8779,N_8674,N_8577);
xor U8780 (N_8780,N_8698,N_8578);
and U8781 (N_8781,N_8739,N_8564);
xnor U8782 (N_8782,N_8565,N_8522);
or U8783 (N_8783,N_8579,N_8625);
nand U8784 (N_8784,N_8585,N_8559);
or U8785 (N_8785,N_8620,N_8699);
xnor U8786 (N_8786,N_8613,N_8681);
nand U8787 (N_8787,N_8695,N_8645);
or U8788 (N_8788,N_8607,N_8706);
and U8789 (N_8789,N_8510,N_8638);
and U8790 (N_8790,N_8708,N_8531);
or U8791 (N_8791,N_8506,N_8647);
nor U8792 (N_8792,N_8734,N_8631);
nor U8793 (N_8793,N_8630,N_8710);
xnor U8794 (N_8794,N_8608,N_8694);
or U8795 (N_8795,N_8686,N_8738);
nor U8796 (N_8796,N_8587,N_8524);
and U8797 (N_8797,N_8595,N_8736);
nand U8798 (N_8798,N_8533,N_8511);
and U8799 (N_8799,N_8514,N_8652);
nor U8800 (N_8800,N_8532,N_8591);
xor U8801 (N_8801,N_8741,N_8660);
nand U8802 (N_8802,N_8623,N_8560);
xor U8803 (N_8803,N_8508,N_8538);
xor U8804 (N_8804,N_8568,N_8725);
and U8805 (N_8805,N_8521,N_8659);
xor U8806 (N_8806,N_8505,N_8539);
xnor U8807 (N_8807,N_8748,N_8542);
nor U8808 (N_8808,N_8745,N_8726);
and U8809 (N_8809,N_8720,N_8527);
or U8810 (N_8810,N_8575,N_8582);
nor U8811 (N_8811,N_8544,N_8685);
or U8812 (N_8812,N_8735,N_8525);
nand U8813 (N_8813,N_8651,N_8601);
xnor U8814 (N_8814,N_8729,N_8684);
nor U8815 (N_8815,N_8548,N_8628);
or U8816 (N_8816,N_8519,N_8515);
and U8817 (N_8817,N_8690,N_8633);
or U8818 (N_8818,N_8705,N_8589);
or U8819 (N_8819,N_8673,N_8641);
nand U8820 (N_8820,N_8650,N_8599);
xor U8821 (N_8821,N_8689,N_8624);
or U8822 (N_8822,N_8728,N_8747);
or U8823 (N_8823,N_8637,N_8507);
or U8824 (N_8824,N_8696,N_8636);
nor U8825 (N_8825,N_8604,N_8622);
nand U8826 (N_8826,N_8537,N_8602);
xnor U8827 (N_8827,N_8520,N_8603);
nor U8828 (N_8828,N_8621,N_8664);
and U8829 (N_8829,N_8702,N_8700);
nor U8830 (N_8830,N_8679,N_8543);
or U8831 (N_8831,N_8680,N_8615);
and U8832 (N_8832,N_8658,N_8549);
nand U8833 (N_8833,N_8567,N_8557);
nand U8834 (N_8834,N_8644,N_8742);
and U8835 (N_8835,N_8749,N_8732);
xor U8836 (N_8836,N_8530,N_8554);
nor U8837 (N_8837,N_8574,N_8712);
or U8838 (N_8838,N_8562,N_8501);
and U8839 (N_8839,N_8707,N_8704);
or U8840 (N_8840,N_8667,N_8714);
or U8841 (N_8841,N_8655,N_8512);
xnor U8842 (N_8842,N_8635,N_8563);
xor U8843 (N_8843,N_8590,N_8553);
xnor U8844 (N_8844,N_8713,N_8671);
nand U8845 (N_8845,N_8687,N_8676);
or U8846 (N_8846,N_8653,N_8648);
or U8847 (N_8847,N_8719,N_8746);
and U8848 (N_8848,N_8683,N_8744);
and U8849 (N_8849,N_8518,N_8540);
and U8850 (N_8850,N_8614,N_8730);
xor U8851 (N_8851,N_8646,N_8571);
nor U8852 (N_8852,N_8534,N_8632);
nand U8853 (N_8853,N_8668,N_8517);
nand U8854 (N_8854,N_8703,N_8639);
and U8855 (N_8855,N_8715,N_8513);
and U8856 (N_8856,N_8718,N_8586);
nand U8857 (N_8857,N_8536,N_8731);
and U8858 (N_8858,N_8697,N_8724);
and U8859 (N_8859,N_8584,N_8682);
or U8860 (N_8860,N_8556,N_8656);
and U8861 (N_8861,N_8701,N_8596);
nor U8862 (N_8862,N_8509,N_8627);
nand U8863 (N_8863,N_8678,N_8500);
or U8864 (N_8864,N_8593,N_8642);
xnor U8865 (N_8865,N_8657,N_8666);
nand U8866 (N_8866,N_8717,N_8535);
or U8867 (N_8867,N_8722,N_8723);
xor U8868 (N_8868,N_8576,N_8649);
nand U8869 (N_8869,N_8643,N_8566);
nor U8870 (N_8870,N_8626,N_8502);
or U8871 (N_8871,N_8654,N_8555);
or U8872 (N_8872,N_8592,N_8611);
and U8873 (N_8873,N_8737,N_8618);
nand U8874 (N_8874,N_8545,N_8691);
and U8875 (N_8875,N_8520,N_8535);
or U8876 (N_8876,N_8583,N_8707);
nand U8877 (N_8877,N_8518,N_8647);
and U8878 (N_8878,N_8595,N_8638);
and U8879 (N_8879,N_8588,N_8739);
xnor U8880 (N_8880,N_8559,N_8620);
and U8881 (N_8881,N_8626,N_8533);
nor U8882 (N_8882,N_8726,N_8594);
nor U8883 (N_8883,N_8655,N_8561);
xnor U8884 (N_8884,N_8701,N_8658);
and U8885 (N_8885,N_8510,N_8521);
xor U8886 (N_8886,N_8521,N_8522);
and U8887 (N_8887,N_8658,N_8573);
or U8888 (N_8888,N_8628,N_8740);
or U8889 (N_8889,N_8664,N_8645);
and U8890 (N_8890,N_8705,N_8655);
xor U8891 (N_8891,N_8566,N_8578);
and U8892 (N_8892,N_8503,N_8740);
nor U8893 (N_8893,N_8581,N_8635);
nor U8894 (N_8894,N_8724,N_8541);
or U8895 (N_8895,N_8603,N_8521);
nor U8896 (N_8896,N_8645,N_8624);
nand U8897 (N_8897,N_8543,N_8745);
or U8898 (N_8898,N_8559,N_8737);
or U8899 (N_8899,N_8639,N_8601);
nand U8900 (N_8900,N_8534,N_8731);
nor U8901 (N_8901,N_8643,N_8551);
nor U8902 (N_8902,N_8692,N_8654);
nand U8903 (N_8903,N_8635,N_8587);
and U8904 (N_8904,N_8671,N_8731);
nor U8905 (N_8905,N_8553,N_8589);
nand U8906 (N_8906,N_8738,N_8560);
and U8907 (N_8907,N_8604,N_8567);
or U8908 (N_8908,N_8636,N_8590);
xor U8909 (N_8909,N_8702,N_8532);
xnor U8910 (N_8910,N_8707,N_8521);
xor U8911 (N_8911,N_8510,N_8739);
and U8912 (N_8912,N_8519,N_8712);
xor U8913 (N_8913,N_8743,N_8748);
xor U8914 (N_8914,N_8618,N_8524);
nand U8915 (N_8915,N_8657,N_8727);
nand U8916 (N_8916,N_8579,N_8627);
or U8917 (N_8917,N_8682,N_8658);
nor U8918 (N_8918,N_8678,N_8518);
nor U8919 (N_8919,N_8688,N_8733);
or U8920 (N_8920,N_8579,N_8519);
or U8921 (N_8921,N_8588,N_8574);
nor U8922 (N_8922,N_8727,N_8590);
nor U8923 (N_8923,N_8589,N_8536);
nor U8924 (N_8924,N_8704,N_8576);
nand U8925 (N_8925,N_8669,N_8677);
and U8926 (N_8926,N_8710,N_8727);
or U8927 (N_8927,N_8614,N_8665);
and U8928 (N_8928,N_8587,N_8666);
nor U8929 (N_8929,N_8675,N_8748);
nor U8930 (N_8930,N_8610,N_8504);
or U8931 (N_8931,N_8729,N_8540);
or U8932 (N_8932,N_8713,N_8582);
nand U8933 (N_8933,N_8612,N_8569);
nor U8934 (N_8934,N_8749,N_8748);
nor U8935 (N_8935,N_8620,N_8589);
nor U8936 (N_8936,N_8723,N_8720);
nand U8937 (N_8937,N_8739,N_8642);
nand U8938 (N_8938,N_8602,N_8714);
xnor U8939 (N_8939,N_8727,N_8540);
and U8940 (N_8940,N_8533,N_8556);
or U8941 (N_8941,N_8686,N_8566);
or U8942 (N_8942,N_8744,N_8611);
or U8943 (N_8943,N_8677,N_8639);
nand U8944 (N_8944,N_8748,N_8559);
nor U8945 (N_8945,N_8543,N_8574);
nand U8946 (N_8946,N_8695,N_8742);
nor U8947 (N_8947,N_8730,N_8563);
xor U8948 (N_8948,N_8585,N_8749);
and U8949 (N_8949,N_8565,N_8552);
nand U8950 (N_8950,N_8555,N_8578);
or U8951 (N_8951,N_8528,N_8711);
xnor U8952 (N_8952,N_8655,N_8646);
and U8953 (N_8953,N_8508,N_8724);
and U8954 (N_8954,N_8518,N_8605);
or U8955 (N_8955,N_8595,N_8577);
or U8956 (N_8956,N_8615,N_8662);
and U8957 (N_8957,N_8706,N_8532);
and U8958 (N_8958,N_8652,N_8681);
nand U8959 (N_8959,N_8605,N_8634);
xor U8960 (N_8960,N_8576,N_8524);
xor U8961 (N_8961,N_8710,N_8601);
and U8962 (N_8962,N_8703,N_8518);
nand U8963 (N_8963,N_8676,N_8732);
nor U8964 (N_8964,N_8637,N_8644);
nand U8965 (N_8965,N_8521,N_8595);
and U8966 (N_8966,N_8596,N_8604);
xnor U8967 (N_8967,N_8521,N_8652);
or U8968 (N_8968,N_8626,N_8662);
or U8969 (N_8969,N_8701,N_8733);
or U8970 (N_8970,N_8559,N_8556);
or U8971 (N_8971,N_8618,N_8677);
and U8972 (N_8972,N_8588,N_8513);
nor U8973 (N_8973,N_8561,N_8559);
nor U8974 (N_8974,N_8685,N_8659);
and U8975 (N_8975,N_8723,N_8696);
and U8976 (N_8976,N_8719,N_8712);
nor U8977 (N_8977,N_8537,N_8527);
nor U8978 (N_8978,N_8502,N_8609);
nor U8979 (N_8979,N_8517,N_8663);
nand U8980 (N_8980,N_8567,N_8505);
nand U8981 (N_8981,N_8711,N_8647);
nor U8982 (N_8982,N_8529,N_8656);
and U8983 (N_8983,N_8545,N_8590);
nor U8984 (N_8984,N_8562,N_8569);
nand U8985 (N_8985,N_8728,N_8551);
and U8986 (N_8986,N_8636,N_8585);
and U8987 (N_8987,N_8522,N_8722);
nor U8988 (N_8988,N_8598,N_8562);
nor U8989 (N_8989,N_8570,N_8737);
or U8990 (N_8990,N_8742,N_8662);
nand U8991 (N_8991,N_8534,N_8568);
or U8992 (N_8992,N_8735,N_8726);
or U8993 (N_8993,N_8636,N_8647);
xor U8994 (N_8994,N_8522,N_8578);
nand U8995 (N_8995,N_8661,N_8562);
nand U8996 (N_8996,N_8595,N_8596);
nor U8997 (N_8997,N_8690,N_8525);
nand U8998 (N_8998,N_8719,N_8501);
and U8999 (N_8999,N_8675,N_8716);
nand U9000 (N_9000,N_8936,N_8881);
and U9001 (N_9001,N_8999,N_8941);
nor U9002 (N_9002,N_8813,N_8998);
nor U9003 (N_9003,N_8844,N_8784);
and U9004 (N_9004,N_8848,N_8995);
xnor U9005 (N_9005,N_8760,N_8960);
or U9006 (N_9006,N_8834,N_8951);
and U9007 (N_9007,N_8772,N_8935);
and U9008 (N_9008,N_8766,N_8798);
xor U9009 (N_9009,N_8815,N_8767);
and U9010 (N_9010,N_8948,N_8873);
or U9011 (N_9011,N_8773,N_8962);
or U9012 (N_9012,N_8909,N_8853);
or U9013 (N_9013,N_8836,N_8879);
nor U9014 (N_9014,N_8870,N_8857);
or U9015 (N_9015,N_8753,N_8988);
nor U9016 (N_9016,N_8794,N_8980);
nand U9017 (N_9017,N_8833,N_8974);
xor U9018 (N_9018,N_8905,N_8968);
nor U9019 (N_9019,N_8750,N_8934);
xnor U9020 (N_9020,N_8929,N_8952);
or U9021 (N_9021,N_8820,N_8824);
nor U9022 (N_9022,N_8886,N_8906);
or U9023 (N_9023,N_8975,N_8961);
nand U9024 (N_9024,N_8907,N_8755);
nand U9025 (N_9025,N_8842,N_8808);
and U9026 (N_9026,N_8875,N_8942);
nor U9027 (N_9027,N_8762,N_8983);
nor U9028 (N_9028,N_8858,N_8845);
or U9029 (N_9029,N_8963,N_8829);
xnor U9030 (N_9030,N_8817,N_8825);
xnor U9031 (N_9031,N_8866,N_8774);
and U9032 (N_9032,N_8758,N_8956);
and U9033 (N_9033,N_8850,N_8976);
or U9034 (N_9034,N_8984,N_8970);
nand U9035 (N_9035,N_8797,N_8795);
nand U9036 (N_9036,N_8869,N_8789);
nor U9037 (N_9037,N_8947,N_8780);
xor U9038 (N_9038,N_8899,N_8943);
and U9039 (N_9039,N_8771,N_8764);
nor U9040 (N_9040,N_8818,N_8959);
xor U9041 (N_9041,N_8990,N_8982);
nor U9042 (N_9042,N_8864,N_8992);
nand U9043 (N_9043,N_8776,N_8954);
and U9044 (N_9044,N_8884,N_8788);
xor U9045 (N_9045,N_8893,N_8861);
and U9046 (N_9046,N_8837,N_8918);
nand U9047 (N_9047,N_8926,N_8826);
or U9048 (N_9048,N_8868,N_8900);
or U9049 (N_9049,N_8991,N_8903);
nor U9050 (N_9050,N_8770,N_8832);
xnor U9051 (N_9051,N_8783,N_8892);
nand U9052 (N_9052,N_8811,N_8969);
nand U9053 (N_9053,N_8887,N_8793);
and U9054 (N_9054,N_8777,N_8840);
and U9055 (N_9055,N_8839,N_8902);
nand U9056 (N_9056,N_8806,N_8920);
nand U9057 (N_9057,N_8927,N_8966);
nand U9058 (N_9058,N_8769,N_8821);
or U9059 (N_9059,N_8989,N_8846);
or U9060 (N_9060,N_8804,N_8928);
nor U9061 (N_9061,N_8812,N_8925);
nor U9062 (N_9062,N_8828,N_8977);
and U9063 (N_9063,N_8872,N_8778);
and U9064 (N_9064,N_8955,N_8919);
nor U9065 (N_9065,N_8831,N_8964);
and U9066 (N_9066,N_8827,N_8807);
nand U9067 (N_9067,N_8997,N_8913);
xor U9068 (N_9068,N_8849,N_8986);
and U9069 (N_9069,N_8931,N_8768);
xor U9070 (N_9070,N_8946,N_8854);
nor U9071 (N_9071,N_8862,N_8852);
or U9072 (N_9072,N_8859,N_8871);
or U9073 (N_9073,N_8930,N_8901);
or U9074 (N_9074,N_8754,N_8916);
nand U9075 (N_9075,N_8908,N_8752);
and U9076 (N_9076,N_8994,N_8809);
xnor U9077 (N_9077,N_8971,N_8933);
xor U9078 (N_9078,N_8957,N_8944);
xor U9079 (N_9079,N_8785,N_8912);
or U9080 (N_9080,N_8958,N_8838);
and U9081 (N_9081,N_8803,N_8787);
and U9082 (N_9082,N_8847,N_8967);
and U9083 (N_9083,N_8835,N_8841);
and U9084 (N_9084,N_8757,N_8792);
and U9085 (N_9085,N_8823,N_8759);
xnor U9086 (N_9086,N_8756,N_8880);
xor U9087 (N_9087,N_8973,N_8765);
or U9088 (N_9088,N_8761,N_8945);
nor U9089 (N_9089,N_8896,N_8898);
xnor U9090 (N_9090,N_8786,N_8791);
nand U9091 (N_9091,N_8796,N_8882);
and U9092 (N_9092,N_8855,N_8816);
xor U9093 (N_9093,N_8978,N_8939);
or U9094 (N_9094,N_8822,N_8922);
nand U9095 (N_9095,N_8779,N_8814);
nand U9096 (N_9096,N_8897,N_8781);
nor U9097 (N_9097,N_8830,N_8877);
and U9098 (N_9098,N_8923,N_8751);
xnor U9099 (N_9099,N_8987,N_8843);
or U9100 (N_9100,N_8885,N_8890);
xnor U9101 (N_9101,N_8904,N_8889);
or U9102 (N_9102,N_8981,N_8883);
xnor U9103 (N_9103,N_8805,N_8865);
xor U9104 (N_9104,N_8895,N_8953);
or U9105 (N_9105,N_8921,N_8938);
nand U9106 (N_9106,N_8993,N_8878);
nand U9107 (N_9107,N_8888,N_8940);
and U9108 (N_9108,N_8996,N_8876);
or U9109 (N_9109,N_8782,N_8894);
xnor U9110 (N_9110,N_8800,N_8863);
nand U9111 (N_9111,N_8965,N_8915);
xnor U9112 (N_9112,N_8932,N_8819);
nand U9113 (N_9113,N_8851,N_8790);
nand U9114 (N_9114,N_8949,N_8867);
and U9115 (N_9115,N_8874,N_8810);
or U9116 (N_9116,N_8937,N_8801);
nor U9117 (N_9117,N_8924,N_8911);
and U9118 (N_9118,N_8802,N_8775);
and U9119 (N_9119,N_8910,N_8917);
and U9120 (N_9120,N_8856,N_8763);
nand U9121 (N_9121,N_8799,N_8985);
or U9122 (N_9122,N_8891,N_8950);
xor U9123 (N_9123,N_8860,N_8972);
and U9124 (N_9124,N_8979,N_8914);
or U9125 (N_9125,N_8796,N_8783);
or U9126 (N_9126,N_8970,N_8836);
and U9127 (N_9127,N_8815,N_8802);
xnor U9128 (N_9128,N_8822,N_8886);
and U9129 (N_9129,N_8777,N_8865);
or U9130 (N_9130,N_8793,N_8753);
nand U9131 (N_9131,N_8885,N_8985);
or U9132 (N_9132,N_8933,N_8787);
nand U9133 (N_9133,N_8858,N_8907);
nor U9134 (N_9134,N_8759,N_8866);
xnor U9135 (N_9135,N_8790,N_8869);
nor U9136 (N_9136,N_8919,N_8996);
or U9137 (N_9137,N_8918,N_8860);
and U9138 (N_9138,N_8983,N_8869);
xnor U9139 (N_9139,N_8751,N_8835);
nand U9140 (N_9140,N_8990,N_8948);
xnor U9141 (N_9141,N_8982,N_8787);
xor U9142 (N_9142,N_8940,N_8918);
or U9143 (N_9143,N_8930,N_8779);
nor U9144 (N_9144,N_8807,N_8774);
or U9145 (N_9145,N_8865,N_8982);
and U9146 (N_9146,N_8825,N_8913);
and U9147 (N_9147,N_8982,N_8827);
or U9148 (N_9148,N_8924,N_8916);
nor U9149 (N_9149,N_8884,N_8765);
or U9150 (N_9150,N_8971,N_8821);
nor U9151 (N_9151,N_8798,N_8924);
or U9152 (N_9152,N_8958,N_8991);
or U9153 (N_9153,N_8916,N_8790);
xnor U9154 (N_9154,N_8891,N_8751);
or U9155 (N_9155,N_8869,N_8948);
nor U9156 (N_9156,N_8853,N_8928);
and U9157 (N_9157,N_8817,N_8964);
and U9158 (N_9158,N_8821,N_8752);
nor U9159 (N_9159,N_8911,N_8756);
nand U9160 (N_9160,N_8945,N_8959);
nor U9161 (N_9161,N_8762,N_8886);
xnor U9162 (N_9162,N_8934,N_8918);
nand U9163 (N_9163,N_8847,N_8845);
xnor U9164 (N_9164,N_8980,N_8828);
nor U9165 (N_9165,N_8980,N_8918);
and U9166 (N_9166,N_8758,N_8982);
nor U9167 (N_9167,N_8929,N_8960);
and U9168 (N_9168,N_8790,N_8894);
and U9169 (N_9169,N_8811,N_8996);
and U9170 (N_9170,N_8778,N_8912);
and U9171 (N_9171,N_8947,N_8918);
or U9172 (N_9172,N_8917,N_8893);
and U9173 (N_9173,N_8861,N_8947);
nand U9174 (N_9174,N_8854,N_8978);
nor U9175 (N_9175,N_8960,N_8774);
nor U9176 (N_9176,N_8769,N_8756);
or U9177 (N_9177,N_8949,N_8763);
and U9178 (N_9178,N_8936,N_8873);
nand U9179 (N_9179,N_8873,N_8961);
and U9180 (N_9180,N_8978,N_8884);
nand U9181 (N_9181,N_8793,N_8976);
nor U9182 (N_9182,N_8786,N_8922);
nor U9183 (N_9183,N_8997,N_8837);
and U9184 (N_9184,N_8983,N_8850);
nand U9185 (N_9185,N_8791,N_8858);
nand U9186 (N_9186,N_8757,N_8878);
nor U9187 (N_9187,N_8898,N_8791);
or U9188 (N_9188,N_8870,N_8992);
or U9189 (N_9189,N_8885,N_8847);
xor U9190 (N_9190,N_8926,N_8940);
xnor U9191 (N_9191,N_8968,N_8852);
nor U9192 (N_9192,N_8817,N_8790);
nor U9193 (N_9193,N_8943,N_8933);
nor U9194 (N_9194,N_8947,N_8806);
and U9195 (N_9195,N_8979,N_8907);
xnor U9196 (N_9196,N_8811,N_8789);
nand U9197 (N_9197,N_8908,N_8848);
xnor U9198 (N_9198,N_8821,N_8923);
xnor U9199 (N_9199,N_8978,N_8766);
xor U9200 (N_9200,N_8840,N_8843);
xor U9201 (N_9201,N_8789,N_8861);
nand U9202 (N_9202,N_8779,N_8928);
or U9203 (N_9203,N_8914,N_8865);
nor U9204 (N_9204,N_8933,N_8806);
nor U9205 (N_9205,N_8928,N_8936);
and U9206 (N_9206,N_8944,N_8833);
xor U9207 (N_9207,N_8962,N_8848);
nand U9208 (N_9208,N_8752,N_8856);
xor U9209 (N_9209,N_8988,N_8966);
or U9210 (N_9210,N_8792,N_8809);
and U9211 (N_9211,N_8873,N_8826);
nor U9212 (N_9212,N_8873,N_8761);
nor U9213 (N_9213,N_8873,N_8782);
nand U9214 (N_9214,N_8950,N_8969);
or U9215 (N_9215,N_8963,N_8761);
nor U9216 (N_9216,N_8960,N_8895);
xor U9217 (N_9217,N_8980,N_8977);
xnor U9218 (N_9218,N_8775,N_8956);
xnor U9219 (N_9219,N_8866,N_8915);
nand U9220 (N_9220,N_8791,N_8987);
nor U9221 (N_9221,N_8941,N_8911);
xnor U9222 (N_9222,N_8794,N_8985);
and U9223 (N_9223,N_8892,N_8984);
or U9224 (N_9224,N_8842,N_8815);
and U9225 (N_9225,N_8949,N_8841);
nand U9226 (N_9226,N_8973,N_8810);
and U9227 (N_9227,N_8770,N_8791);
nor U9228 (N_9228,N_8905,N_8963);
nor U9229 (N_9229,N_8819,N_8843);
nand U9230 (N_9230,N_8904,N_8981);
and U9231 (N_9231,N_8952,N_8967);
nand U9232 (N_9232,N_8808,N_8844);
and U9233 (N_9233,N_8839,N_8812);
and U9234 (N_9234,N_8987,N_8773);
nor U9235 (N_9235,N_8922,N_8911);
nand U9236 (N_9236,N_8848,N_8998);
xnor U9237 (N_9237,N_8769,N_8837);
xnor U9238 (N_9238,N_8803,N_8895);
xor U9239 (N_9239,N_8798,N_8809);
nor U9240 (N_9240,N_8801,N_8837);
and U9241 (N_9241,N_8874,N_8957);
or U9242 (N_9242,N_8957,N_8882);
xor U9243 (N_9243,N_8781,N_8792);
xor U9244 (N_9244,N_8873,N_8891);
xnor U9245 (N_9245,N_8946,N_8771);
or U9246 (N_9246,N_8767,N_8936);
xor U9247 (N_9247,N_8985,N_8756);
nand U9248 (N_9248,N_8797,N_8976);
nor U9249 (N_9249,N_8768,N_8945);
xnor U9250 (N_9250,N_9228,N_9127);
and U9251 (N_9251,N_9012,N_9234);
or U9252 (N_9252,N_9207,N_9033);
or U9253 (N_9253,N_9211,N_9122);
nor U9254 (N_9254,N_9210,N_9105);
nand U9255 (N_9255,N_9133,N_9071);
xor U9256 (N_9256,N_9103,N_9177);
nand U9257 (N_9257,N_9054,N_9028);
or U9258 (N_9258,N_9227,N_9137);
or U9259 (N_9259,N_9040,N_9246);
nand U9260 (N_9260,N_9126,N_9161);
and U9261 (N_9261,N_9092,N_9077);
nand U9262 (N_9262,N_9183,N_9169);
and U9263 (N_9263,N_9166,N_9194);
or U9264 (N_9264,N_9082,N_9235);
and U9265 (N_9265,N_9130,N_9223);
or U9266 (N_9266,N_9044,N_9001);
xor U9267 (N_9267,N_9062,N_9022);
xnor U9268 (N_9268,N_9242,N_9031);
or U9269 (N_9269,N_9099,N_9164);
and U9270 (N_9270,N_9019,N_9025);
xnor U9271 (N_9271,N_9212,N_9060);
nor U9272 (N_9272,N_9072,N_9029);
and U9273 (N_9273,N_9041,N_9155);
and U9274 (N_9274,N_9139,N_9030);
and U9275 (N_9275,N_9148,N_9093);
xor U9276 (N_9276,N_9063,N_9096);
nand U9277 (N_9277,N_9231,N_9004);
and U9278 (N_9278,N_9229,N_9075);
or U9279 (N_9279,N_9061,N_9221);
nand U9280 (N_9280,N_9247,N_9051);
nand U9281 (N_9281,N_9125,N_9083);
or U9282 (N_9282,N_9239,N_9230);
and U9283 (N_9283,N_9015,N_9232);
nor U9284 (N_9284,N_9209,N_9045);
nand U9285 (N_9285,N_9129,N_9185);
nand U9286 (N_9286,N_9032,N_9007);
xor U9287 (N_9287,N_9165,N_9128);
or U9288 (N_9288,N_9167,N_9188);
nor U9289 (N_9289,N_9184,N_9141);
nand U9290 (N_9290,N_9085,N_9248);
and U9291 (N_9291,N_9008,N_9023);
or U9292 (N_9292,N_9198,N_9186);
and U9293 (N_9293,N_9233,N_9024);
or U9294 (N_9294,N_9100,N_9034);
and U9295 (N_9295,N_9055,N_9011);
nor U9296 (N_9296,N_9218,N_9240);
xor U9297 (N_9297,N_9182,N_9190);
nor U9298 (N_9298,N_9238,N_9199);
nor U9299 (N_9299,N_9116,N_9195);
xor U9300 (N_9300,N_9162,N_9157);
nor U9301 (N_9301,N_9170,N_9236);
nor U9302 (N_9302,N_9158,N_9108);
xnor U9303 (N_9303,N_9215,N_9109);
nor U9304 (N_9304,N_9149,N_9081);
nor U9305 (N_9305,N_9089,N_9053);
xnor U9306 (N_9306,N_9136,N_9144);
xnor U9307 (N_9307,N_9104,N_9052);
xnor U9308 (N_9308,N_9039,N_9078);
and U9309 (N_9309,N_9106,N_9244);
nand U9310 (N_9310,N_9097,N_9009);
or U9311 (N_9311,N_9143,N_9115);
xnor U9312 (N_9312,N_9241,N_9005);
or U9313 (N_9313,N_9159,N_9002);
and U9314 (N_9314,N_9135,N_9095);
xor U9315 (N_9315,N_9111,N_9056);
and U9316 (N_9316,N_9204,N_9168);
nand U9317 (N_9317,N_9131,N_9018);
nand U9318 (N_9318,N_9020,N_9213);
nand U9319 (N_9319,N_9064,N_9088);
or U9320 (N_9320,N_9059,N_9147);
nand U9321 (N_9321,N_9079,N_9065);
or U9322 (N_9322,N_9117,N_9171);
or U9323 (N_9323,N_9021,N_9226);
or U9324 (N_9324,N_9132,N_9037);
or U9325 (N_9325,N_9098,N_9140);
and U9326 (N_9326,N_9123,N_9094);
nor U9327 (N_9327,N_9113,N_9026);
xnor U9328 (N_9328,N_9205,N_9118);
and U9329 (N_9329,N_9193,N_9010);
xor U9330 (N_9330,N_9220,N_9181);
and U9331 (N_9331,N_9175,N_9013);
or U9332 (N_9332,N_9016,N_9086);
nor U9333 (N_9333,N_9043,N_9206);
nor U9334 (N_9334,N_9107,N_9202);
xor U9335 (N_9335,N_9042,N_9080);
and U9336 (N_9336,N_9066,N_9102);
and U9337 (N_9337,N_9119,N_9146);
or U9338 (N_9338,N_9057,N_9249);
or U9339 (N_9339,N_9027,N_9237);
and U9340 (N_9340,N_9178,N_9049);
nor U9341 (N_9341,N_9069,N_9067);
or U9342 (N_9342,N_9160,N_9180);
nand U9343 (N_9343,N_9200,N_9224);
nand U9344 (N_9344,N_9038,N_9121);
or U9345 (N_9345,N_9068,N_9191);
or U9346 (N_9346,N_9156,N_9163);
nand U9347 (N_9347,N_9090,N_9035);
or U9348 (N_9348,N_9112,N_9145);
nor U9349 (N_9349,N_9196,N_9172);
nand U9350 (N_9350,N_9087,N_9208);
xnor U9351 (N_9351,N_9217,N_9070);
and U9352 (N_9352,N_9203,N_9074);
or U9353 (N_9353,N_9189,N_9243);
nand U9354 (N_9354,N_9114,N_9214);
nand U9355 (N_9355,N_9222,N_9110);
nor U9356 (N_9356,N_9187,N_9153);
nand U9357 (N_9357,N_9058,N_9216);
nand U9358 (N_9358,N_9046,N_9091);
xor U9359 (N_9359,N_9174,N_9154);
or U9360 (N_9360,N_9047,N_9150);
nand U9361 (N_9361,N_9173,N_9120);
or U9362 (N_9362,N_9197,N_9201);
nor U9363 (N_9363,N_9245,N_9003);
xor U9364 (N_9364,N_9176,N_9138);
nor U9365 (N_9365,N_9124,N_9073);
nor U9366 (N_9366,N_9050,N_9017);
xor U9367 (N_9367,N_9225,N_9036);
nor U9368 (N_9368,N_9076,N_9014);
xnor U9369 (N_9369,N_9192,N_9152);
and U9370 (N_9370,N_9048,N_9219);
xor U9371 (N_9371,N_9084,N_9134);
or U9372 (N_9372,N_9000,N_9006);
xor U9373 (N_9373,N_9101,N_9142);
nand U9374 (N_9374,N_9151,N_9179);
nor U9375 (N_9375,N_9216,N_9111);
nor U9376 (N_9376,N_9127,N_9083);
and U9377 (N_9377,N_9100,N_9080);
or U9378 (N_9378,N_9029,N_9038);
xor U9379 (N_9379,N_9230,N_9035);
xor U9380 (N_9380,N_9130,N_9162);
nand U9381 (N_9381,N_9017,N_9210);
or U9382 (N_9382,N_9098,N_9148);
nand U9383 (N_9383,N_9166,N_9029);
nand U9384 (N_9384,N_9092,N_9010);
nand U9385 (N_9385,N_9149,N_9203);
or U9386 (N_9386,N_9114,N_9044);
xnor U9387 (N_9387,N_9246,N_9161);
nor U9388 (N_9388,N_9018,N_9209);
xnor U9389 (N_9389,N_9040,N_9125);
and U9390 (N_9390,N_9221,N_9112);
and U9391 (N_9391,N_9006,N_9156);
or U9392 (N_9392,N_9133,N_9154);
nor U9393 (N_9393,N_9068,N_9239);
nand U9394 (N_9394,N_9013,N_9039);
or U9395 (N_9395,N_9121,N_9101);
and U9396 (N_9396,N_9130,N_9192);
xnor U9397 (N_9397,N_9221,N_9136);
and U9398 (N_9398,N_9050,N_9190);
xnor U9399 (N_9399,N_9078,N_9142);
nand U9400 (N_9400,N_9213,N_9173);
and U9401 (N_9401,N_9004,N_9211);
nor U9402 (N_9402,N_9100,N_9230);
xor U9403 (N_9403,N_9105,N_9215);
and U9404 (N_9404,N_9246,N_9155);
nor U9405 (N_9405,N_9132,N_9170);
and U9406 (N_9406,N_9138,N_9114);
and U9407 (N_9407,N_9125,N_9220);
xnor U9408 (N_9408,N_9057,N_9019);
or U9409 (N_9409,N_9234,N_9025);
nand U9410 (N_9410,N_9080,N_9235);
xor U9411 (N_9411,N_9029,N_9115);
nor U9412 (N_9412,N_9109,N_9110);
or U9413 (N_9413,N_9197,N_9165);
nor U9414 (N_9414,N_9232,N_9211);
nor U9415 (N_9415,N_9160,N_9017);
nor U9416 (N_9416,N_9023,N_9127);
and U9417 (N_9417,N_9064,N_9243);
xor U9418 (N_9418,N_9178,N_9056);
and U9419 (N_9419,N_9067,N_9008);
or U9420 (N_9420,N_9028,N_9113);
nor U9421 (N_9421,N_9007,N_9041);
nor U9422 (N_9422,N_9042,N_9236);
and U9423 (N_9423,N_9100,N_9009);
xnor U9424 (N_9424,N_9038,N_9112);
nor U9425 (N_9425,N_9156,N_9111);
or U9426 (N_9426,N_9011,N_9015);
nand U9427 (N_9427,N_9118,N_9175);
or U9428 (N_9428,N_9049,N_9081);
and U9429 (N_9429,N_9169,N_9179);
or U9430 (N_9430,N_9130,N_9151);
nand U9431 (N_9431,N_9100,N_9057);
or U9432 (N_9432,N_9018,N_9210);
xor U9433 (N_9433,N_9158,N_9157);
or U9434 (N_9434,N_9070,N_9172);
or U9435 (N_9435,N_9162,N_9007);
or U9436 (N_9436,N_9151,N_9076);
xnor U9437 (N_9437,N_9121,N_9013);
and U9438 (N_9438,N_9032,N_9104);
xnor U9439 (N_9439,N_9070,N_9124);
and U9440 (N_9440,N_9140,N_9072);
or U9441 (N_9441,N_9085,N_9207);
xnor U9442 (N_9442,N_9185,N_9178);
nand U9443 (N_9443,N_9174,N_9143);
and U9444 (N_9444,N_9015,N_9005);
and U9445 (N_9445,N_9037,N_9040);
nor U9446 (N_9446,N_9199,N_9043);
and U9447 (N_9447,N_9008,N_9014);
nand U9448 (N_9448,N_9033,N_9204);
nand U9449 (N_9449,N_9169,N_9135);
or U9450 (N_9450,N_9127,N_9103);
or U9451 (N_9451,N_9023,N_9143);
and U9452 (N_9452,N_9195,N_9151);
or U9453 (N_9453,N_9242,N_9057);
xor U9454 (N_9454,N_9197,N_9143);
or U9455 (N_9455,N_9002,N_9122);
xor U9456 (N_9456,N_9157,N_9138);
nand U9457 (N_9457,N_9139,N_9031);
xnor U9458 (N_9458,N_9143,N_9074);
or U9459 (N_9459,N_9120,N_9116);
nor U9460 (N_9460,N_9176,N_9042);
nand U9461 (N_9461,N_9088,N_9181);
or U9462 (N_9462,N_9231,N_9042);
or U9463 (N_9463,N_9071,N_9096);
nor U9464 (N_9464,N_9108,N_9015);
xnor U9465 (N_9465,N_9157,N_9131);
nor U9466 (N_9466,N_9247,N_9150);
nand U9467 (N_9467,N_9171,N_9237);
nand U9468 (N_9468,N_9226,N_9063);
nand U9469 (N_9469,N_9218,N_9100);
and U9470 (N_9470,N_9185,N_9028);
nor U9471 (N_9471,N_9076,N_9066);
nand U9472 (N_9472,N_9211,N_9152);
xnor U9473 (N_9473,N_9113,N_9139);
xnor U9474 (N_9474,N_9070,N_9094);
or U9475 (N_9475,N_9061,N_9136);
nor U9476 (N_9476,N_9243,N_9138);
and U9477 (N_9477,N_9203,N_9196);
nor U9478 (N_9478,N_9138,N_9194);
nand U9479 (N_9479,N_9170,N_9124);
or U9480 (N_9480,N_9056,N_9113);
nand U9481 (N_9481,N_9147,N_9023);
and U9482 (N_9482,N_9108,N_9183);
nand U9483 (N_9483,N_9247,N_9221);
or U9484 (N_9484,N_9106,N_9074);
xnor U9485 (N_9485,N_9110,N_9067);
or U9486 (N_9486,N_9131,N_9184);
nor U9487 (N_9487,N_9011,N_9135);
xnor U9488 (N_9488,N_9065,N_9153);
nand U9489 (N_9489,N_9015,N_9027);
or U9490 (N_9490,N_9057,N_9004);
or U9491 (N_9491,N_9091,N_9079);
nand U9492 (N_9492,N_9106,N_9142);
and U9493 (N_9493,N_9063,N_9136);
xor U9494 (N_9494,N_9148,N_9116);
nor U9495 (N_9495,N_9021,N_9018);
xor U9496 (N_9496,N_9103,N_9016);
and U9497 (N_9497,N_9056,N_9075);
xor U9498 (N_9498,N_9087,N_9009);
xor U9499 (N_9499,N_9232,N_9066);
or U9500 (N_9500,N_9481,N_9302);
nand U9501 (N_9501,N_9321,N_9398);
nor U9502 (N_9502,N_9389,N_9379);
nor U9503 (N_9503,N_9427,N_9299);
or U9504 (N_9504,N_9315,N_9309);
xnor U9505 (N_9505,N_9323,N_9393);
nand U9506 (N_9506,N_9382,N_9420);
and U9507 (N_9507,N_9395,N_9385);
or U9508 (N_9508,N_9284,N_9347);
or U9509 (N_9509,N_9449,N_9311);
or U9510 (N_9510,N_9308,N_9346);
xnor U9511 (N_9511,N_9350,N_9258);
nor U9512 (N_9512,N_9274,N_9254);
or U9513 (N_9513,N_9403,N_9278);
xnor U9514 (N_9514,N_9328,N_9461);
or U9515 (N_9515,N_9355,N_9300);
or U9516 (N_9516,N_9335,N_9455);
or U9517 (N_9517,N_9307,N_9368);
or U9518 (N_9518,N_9276,N_9338);
or U9519 (N_9519,N_9405,N_9377);
xor U9520 (N_9520,N_9289,N_9447);
nor U9521 (N_9521,N_9467,N_9290);
and U9522 (N_9522,N_9348,N_9264);
nor U9523 (N_9523,N_9418,N_9361);
xnor U9524 (N_9524,N_9486,N_9411);
nand U9525 (N_9525,N_9425,N_9415);
nor U9526 (N_9526,N_9458,N_9330);
nor U9527 (N_9527,N_9400,N_9443);
or U9528 (N_9528,N_9292,N_9497);
nand U9529 (N_9529,N_9325,N_9391);
or U9530 (N_9530,N_9424,N_9466);
nand U9531 (N_9531,N_9305,N_9472);
or U9532 (N_9532,N_9270,N_9439);
nand U9533 (N_9533,N_9375,N_9373);
or U9534 (N_9534,N_9362,N_9257);
or U9535 (N_9535,N_9478,N_9322);
nor U9536 (N_9536,N_9429,N_9293);
nor U9537 (N_9537,N_9468,N_9370);
nor U9538 (N_9538,N_9386,N_9310);
and U9539 (N_9539,N_9487,N_9261);
nor U9540 (N_9540,N_9471,N_9482);
nor U9541 (N_9541,N_9268,N_9477);
nand U9542 (N_9542,N_9301,N_9483);
and U9543 (N_9543,N_9410,N_9263);
xnor U9544 (N_9544,N_9456,N_9314);
nor U9545 (N_9545,N_9374,N_9460);
or U9546 (N_9546,N_9250,N_9402);
nor U9547 (N_9547,N_9446,N_9457);
or U9548 (N_9548,N_9435,N_9383);
nor U9549 (N_9549,N_9272,N_9416);
xnor U9550 (N_9550,N_9291,N_9253);
or U9551 (N_9551,N_9412,N_9488);
nand U9552 (N_9552,N_9354,N_9331);
nand U9553 (N_9553,N_9436,N_9295);
or U9554 (N_9554,N_9332,N_9353);
and U9555 (N_9555,N_9288,N_9495);
xnor U9556 (N_9556,N_9494,N_9359);
and U9557 (N_9557,N_9426,N_9404);
xnor U9558 (N_9558,N_9320,N_9256);
and U9559 (N_9559,N_9365,N_9450);
nor U9560 (N_9560,N_9358,N_9465);
and U9561 (N_9561,N_9452,N_9397);
nand U9562 (N_9562,N_9448,N_9316);
nand U9563 (N_9563,N_9437,N_9409);
or U9564 (N_9564,N_9312,N_9342);
and U9565 (N_9565,N_9419,N_9369);
or U9566 (N_9566,N_9333,N_9399);
nand U9567 (N_9567,N_9485,N_9479);
or U9568 (N_9568,N_9407,N_9378);
or U9569 (N_9569,N_9296,N_9324);
or U9570 (N_9570,N_9297,N_9306);
xor U9571 (N_9571,N_9431,N_9280);
xor U9572 (N_9572,N_9414,N_9489);
xor U9573 (N_9573,N_9387,N_9341);
or U9574 (N_9574,N_9251,N_9493);
or U9575 (N_9575,N_9445,N_9434);
or U9576 (N_9576,N_9262,N_9364);
nor U9577 (N_9577,N_9255,N_9408);
nor U9578 (N_9578,N_9496,N_9396);
and U9579 (N_9579,N_9473,N_9438);
nor U9580 (N_9580,N_9269,N_9340);
nor U9581 (N_9581,N_9421,N_9337);
xor U9582 (N_9582,N_9475,N_9294);
nand U9583 (N_9583,N_9360,N_9454);
nor U9584 (N_9584,N_9286,N_9417);
xor U9585 (N_9585,N_9317,N_9381);
nor U9586 (N_9586,N_9371,N_9499);
nand U9587 (N_9587,N_9336,N_9356);
or U9588 (N_9588,N_9392,N_9480);
nor U9589 (N_9589,N_9376,N_9329);
nor U9590 (N_9590,N_9304,N_9345);
and U9591 (N_9591,N_9351,N_9394);
xnor U9592 (N_9592,N_9444,N_9252);
nand U9593 (N_9593,N_9367,N_9285);
nor U9594 (N_9594,N_9422,N_9287);
or U9595 (N_9595,N_9491,N_9339);
or U9596 (N_9596,N_9343,N_9484);
or U9597 (N_9597,N_9463,N_9462);
nor U9598 (N_9598,N_9459,N_9476);
xnor U9599 (N_9599,N_9453,N_9349);
nand U9600 (N_9600,N_9401,N_9275);
xnor U9601 (N_9601,N_9388,N_9474);
and U9602 (N_9602,N_9366,N_9260);
and U9603 (N_9603,N_9319,N_9464);
and U9604 (N_9604,N_9281,N_9440);
xor U9605 (N_9605,N_9344,N_9273);
or U9606 (N_9606,N_9490,N_9267);
nand U9607 (N_9607,N_9265,N_9492);
and U9608 (N_9608,N_9313,N_9298);
or U9609 (N_9609,N_9326,N_9266);
or U9610 (N_9610,N_9430,N_9259);
nor U9611 (N_9611,N_9372,N_9282);
nor U9612 (N_9612,N_9451,N_9428);
or U9613 (N_9613,N_9432,N_9406);
xnor U9614 (N_9614,N_9334,N_9380);
or U9615 (N_9615,N_9279,N_9327);
or U9616 (N_9616,N_9433,N_9413);
nand U9617 (N_9617,N_9469,N_9318);
xor U9618 (N_9618,N_9283,N_9352);
xor U9619 (N_9619,N_9423,N_9277);
nand U9620 (N_9620,N_9441,N_9357);
nor U9621 (N_9621,N_9442,N_9384);
and U9622 (N_9622,N_9363,N_9498);
or U9623 (N_9623,N_9271,N_9390);
or U9624 (N_9624,N_9470,N_9303);
or U9625 (N_9625,N_9462,N_9469);
nor U9626 (N_9626,N_9300,N_9316);
nor U9627 (N_9627,N_9404,N_9376);
nand U9628 (N_9628,N_9416,N_9470);
nor U9629 (N_9629,N_9384,N_9250);
nand U9630 (N_9630,N_9402,N_9480);
nand U9631 (N_9631,N_9434,N_9453);
xnor U9632 (N_9632,N_9304,N_9328);
nor U9633 (N_9633,N_9266,N_9397);
nand U9634 (N_9634,N_9302,N_9443);
nor U9635 (N_9635,N_9279,N_9407);
xnor U9636 (N_9636,N_9308,N_9376);
and U9637 (N_9637,N_9281,N_9315);
and U9638 (N_9638,N_9302,N_9437);
and U9639 (N_9639,N_9357,N_9320);
or U9640 (N_9640,N_9319,N_9380);
nand U9641 (N_9641,N_9313,N_9476);
and U9642 (N_9642,N_9444,N_9475);
nor U9643 (N_9643,N_9370,N_9343);
nor U9644 (N_9644,N_9259,N_9290);
nand U9645 (N_9645,N_9274,N_9382);
and U9646 (N_9646,N_9465,N_9425);
or U9647 (N_9647,N_9401,N_9287);
nor U9648 (N_9648,N_9493,N_9475);
nand U9649 (N_9649,N_9356,N_9253);
or U9650 (N_9650,N_9253,N_9467);
xnor U9651 (N_9651,N_9368,N_9472);
and U9652 (N_9652,N_9438,N_9268);
and U9653 (N_9653,N_9345,N_9382);
xor U9654 (N_9654,N_9443,N_9317);
and U9655 (N_9655,N_9311,N_9474);
nand U9656 (N_9656,N_9446,N_9404);
and U9657 (N_9657,N_9386,N_9273);
or U9658 (N_9658,N_9479,N_9321);
or U9659 (N_9659,N_9336,N_9477);
or U9660 (N_9660,N_9296,N_9399);
or U9661 (N_9661,N_9263,N_9425);
xor U9662 (N_9662,N_9312,N_9480);
nor U9663 (N_9663,N_9443,N_9331);
or U9664 (N_9664,N_9476,N_9477);
or U9665 (N_9665,N_9370,N_9266);
or U9666 (N_9666,N_9310,N_9316);
xnor U9667 (N_9667,N_9353,N_9374);
nor U9668 (N_9668,N_9453,N_9328);
nor U9669 (N_9669,N_9355,N_9264);
and U9670 (N_9670,N_9472,N_9478);
xor U9671 (N_9671,N_9260,N_9393);
nand U9672 (N_9672,N_9303,N_9471);
and U9673 (N_9673,N_9467,N_9286);
nand U9674 (N_9674,N_9374,N_9282);
or U9675 (N_9675,N_9381,N_9475);
or U9676 (N_9676,N_9340,N_9377);
xnor U9677 (N_9677,N_9347,N_9471);
or U9678 (N_9678,N_9374,N_9457);
and U9679 (N_9679,N_9426,N_9442);
or U9680 (N_9680,N_9293,N_9353);
xnor U9681 (N_9681,N_9435,N_9486);
xor U9682 (N_9682,N_9266,N_9341);
nor U9683 (N_9683,N_9339,N_9356);
or U9684 (N_9684,N_9289,N_9496);
nand U9685 (N_9685,N_9440,N_9292);
xnor U9686 (N_9686,N_9404,N_9311);
and U9687 (N_9687,N_9255,N_9252);
xor U9688 (N_9688,N_9362,N_9296);
and U9689 (N_9689,N_9376,N_9409);
and U9690 (N_9690,N_9360,N_9373);
or U9691 (N_9691,N_9303,N_9359);
and U9692 (N_9692,N_9271,N_9351);
or U9693 (N_9693,N_9347,N_9379);
xor U9694 (N_9694,N_9289,N_9464);
and U9695 (N_9695,N_9448,N_9491);
nor U9696 (N_9696,N_9487,N_9426);
nor U9697 (N_9697,N_9280,N_9359);
xnor U9698 (N_9698,N_9435,N_9401);
or U9699 (N_9699,N_9320,N_9364);
xnor U9700 (N_9700,N_9443,N_9483);
nor U9701 (N_9701,N_9446,N_9456);
and U9702 (N_9702,N_9478,N_9454);
nor U9703 (N_9703,N_9339,N_9255);
or U9704 (N_9704,N_9343,N_9451);
nand U9705 (N_9705,N_9440,N_9252);
and U9706 (N_9706,N_9327,N_9416);
nand U9707 (N_9707,N_9280,N_9409);
or U9708 (N_9708,N_9255,N_9266);
and U9709 (N_9709,N_9258,N_9297);
nand U9710 (N_9710,N_9486,N_9364);
or U9711 (N_9711,N_9484,N_9356);
and U9712 (N_9712,N_9394,N_9471);
and U9713 (N_9713,N_9334,N_9347);
nand U9714 (N_9714,N_9354,N_9469);
and U9715 (N_9715,N_9326,N_9340);
nand U9716 (N_9716,N_9402,N_9306);
or U9717 (N_9717,N_9395,N_9403);
or U9718 (N_9718,N_9267,N_9355);
nand U9719 (N_9719,N_9299,N_9429);
nand U9720 (N_9720,N_9374,N_9391);
nand U9721 (N_9721,N_9455,N_9275);
xnor U9722 (N_9722,N_9480,N_9257);
nand U9723 (N_9723,N_9380,N_9450);
xnor U9724 (N_9724,N_9491,N_9382);
nand U9725 (N_9725,N_9465,N_9468);
nor U9726 (N_9726,N_9487,N_9447);
nand U9727 (N_9727,N_9448,N_9492);
nand U9728 (N_9728,N_9474,N_9437);
nor U9729 (N_9729,N_9335,N_9330);
xor U9730 (N_9730,N_9336,N_9338);
and U9731 (N_9731,N_9371,N_9294);
nand U9732 (N_9732,N_9414,N_9463);
nand U9733 (N_9733,N_9338,N_9467);
xnor U9734 (N_9734,N_9317,N_9491);
or U9735 (N_9735,N_9434,N_9252);
xor U9736 (N_9736,N_9308,N_9419);
or U9737 (N_9737,N_9321,N_9420);
nor U9738 (N_9738,N_9455,N_9409);
and U9739 (N_9739,N_9445,N_9266);
nand U9740 (N_9740,N_9459,N_9274);
nor U9741 (N_9741,N_9480,N_9459);
nand U9742 (N_9742,N_9315,N_9403);
or U9743 (N_9743,N_9327,N_9432);
and U9744 (N_9744,N_9369,N_9451);
nor U9745 (N_9745,N_9477,N_9384);
or U9746 (N_9746,N_9271,N_9414);
xnor U9747 (N_9747,N_9383,N_9388);
xnor U9748 (N_9748,N_9461,N_9462);
nand U9749 (N_9749,N_9330,N_9423);
and U9750 (N_9750,N_9672,N_9607);
nor U9751 (N_9751,N_9601,N_9714);
nor U9752 (N_9752,N_9608,N_9741);
or U9753 (N_9753,N_9550,N_9517);
nand U9754 (N_9754,N_9560,N_9666);
nand U9755 (N_9755,N_9745,N_9726);
nor U9756 (N_9756,N_9724,N_9504);
xnor U9757 (N_9757,N_9589,N_9682);
or U9758 (N_9758,N_9582,N_9588);
and U9759 (N_9759,N_9651,N_9541);
nand U9760 (N_9760,N_9514,N_9639);
nand U9761 (N_9761,N_9580,N_9576);
xnor U9762 (N_9762,N_9667,N_9543);
xor U9763 (N_9763,N_9509,N_9523);
nor U9764 (N_9764,N_9524,N_9681);
nand U9765 (N_9765,N_9697,N_9669);
and U9766 (N_9766,N_9725,N_9644);
nand U9767 (N_9767,N_9605,N_9629);
or U9768 (N_9768,N_9719,N_9620);
and U9769 (N_9769,N_9641,N_9649);
nor U9770 (N_9770,N_9547,N_9612);
nor U9771 (N_9771,N_9567,N_9532);
or U9772 (N_9772,N_9659,N_9510);
xnor U9773 (N_9773,N_9581,N_9674);
nand U9774 (N_9774,N_9687,N_9614);
nand U9775 (N_9775,N_9729,N_9579);
xor U9776 (N_9776,N_9544,N_9522);
and U9777 (N_9777,N_9707,N_9630);
and U9778 (N_9778,N_9652,N_9529);
nor U9779 (N_9779,N_9556,N_9684);
and U9780 (N_9780,N_9631,N_9671);
nand U9781 (N_9781,N_9721,N_9633);
nor U9782 (N_9782,N_9538,N_9548);
nor U9783 (N_9783,N_9638,N_9545);
nand U9784 (N_9784,N_9683,N_9685);
or U9785 (N_9785,N_9731,N_9735);
or U9786 (N_9786,N_9637,N_9564);
nand U9787 (N_9787,N_9695,N_9555);
nand U9788 (N_9788,N_9570,N_9624);
nor U9789 (N_9789,N_9506,N_9699);
xnor U9790 (N_9790,N_9643,N_9655);
nand U9791 (N_9791,N_9645,N_9673);
or U9792 (N_9792,N_9635,N_9518);
xnor U9793 (N_9793,N_9626,N_9646);
and U9794 (N_9794,N_9568,N_9656);
xor U9795 (N_9795,N_9572,N_9573);
nor U9796 (N_9796,N_9705,N_9546);
nor U9797 (N_9797,N_9539,N_9536);
and U9798 (N_9798,N_9647,N_9528);
nand U9799 (N_9799,N_9531,N_9689);
nor U9800 (N_9800,N_9734,N_9521);
nor U9801 (N_9801,N_9599,N_9696);
and U9802 (N_9802,N_9617,N_9593);
or U9803 (N_9803,N_9535,N_9525);
or U9804 (N_9804,N_9636,N_9688);
and U9805 (N_9805,N_9590,N_9500);
nor U9806 (N_9806,N_9618,N_9508);
nand U9807 (N_9807,N_9664,N_9616);
or U9808 (N_9808,N_9584,N_9662);
and U9809 (N_9809,N_9679,N_9716);
xnor U9810 (N_9810,N_9565,N_9507);
nand U9811 (N_9811,N_9686,N_9742);
nand U9812 (N_9812,N_9658,N_9661);
and U9813 (N_9813,N_9732,N_9746);
xor U9814 (N_9814,N_9738,N_9613);
and U9815 (N_9815,N_9516,N_9503);
or U9816 (N_9816,N_9512,N_9712);
or U9817 (N_9817,N_9709,N_9747);
xnor U9818 (N_9818,N_9625,N_9534);
nor U9819 (N_9819,N_9577,N_9602);
nand U9820 (N_9820,N_9553,N_9610);
or U9821 (N_9821,N_9733,N_9693);
nor U9822 (N_9822,N_9520,N_9596);
and U9823 (N_9823,N_9583,N_9603);
xor U9824 (N_9824,N_9744,N_9694);
and U9825 (N_9825,N_9597,N_9549);
xor U9826 (N_9826,N_9670,N_9701);
and U9827 (N_9827,N_9710,N_9749);
nor U9828 (N_9828,N_9628,N_9604);
or U9829 (N_9829,N_9540,N_9530);
xnor U9830 (N_9830,N_9619,N_9598);
or U9831 (N_9831,N_9501,N_9727);
nand U9832 (N_9832,N_9515,N_9702);
nand U9833 (N_9833,N_9723,N_9708);
nor U9834 (N_9834,N_9587,N_9663);
and U9835 (N_9835,N_9640,N_9657);
or U9836 (N_9836,N_9563,N_9527);
nor U9837 (N_9837,N_9703,N_9678);
nand U9838 (N_9838,N_9737,N_9711);
and U9839 (N_9839,N_9706,N_9575);
and U9840 (N_9840,N_9627,N_9542);
nor U9841 (N_9841,N_9648,N_9730);
nor U9842 (N_9842,N_9586,N_9591);
xnor U9843 (N_9843,N_9675,N_9634);
or U9844 (N_9844,N_9718,N_9717);
and U9845 (N_9845,N_9665,N_9704);
nor U9846 (N_9846,N_9622,N_9552);
and U9847 (N_9847,N_9551,N_9505);
and U9848 (N_9848,N_9574,N_9677);
xor U9849 (N_9849,N_9690,N_9680);
xor U9850 (N_9850,N_9740,N_9502);
xnor U9851 (N_9851,N_9592,N_9511);
nand U9852 (N_9852,N_9743,N_9562);
xor U9853 (N_9853,N_9739,N_9611);
or U9854 (N_9854,N_9558,N_9715);
xnor U9855 (N_9855,N_9722,N_9606);
nor U9856 (N_9856,N_9632,N_9728);
nand U9857 (N_9857,N_9615,N_9650);
nor U9858 (N_9858,N_9660,N_9569);
nand U9859 (N_9859,N_9537,N_9557);
or U9860 (N_9860,N_9654,N_9533);
nor U9861 (N_9861,N_9561,N_9691);
nand U9862 (N_9862,N_9642,N_9513);
nand U9863 (N_9863,N_9571,N_9595);
nor U9864 (N_9864,N_9609,N_9585);
nand U9865 (N_9865,N_9600,N_9713);
xnor U9866 (N_9866,N_9621,N_9526);
nor U9867 (N_9867,N_9748,N_9578);
nand U9868 (N_9868,N_9698,N_9668);
nor U9869 (N_9869,N_9594,N_9720);
nand U9870 (N_9870,N_9559,N_9554);
nand U9871 (N_9871,N_9700,N_9692);
xor U9872 (N_9872,N_9623,N_9736);
and U9873 (N_9873,N_9676,N_9519);
and U9874 (N_9874,N_9566,N_9653);
xnor U9875 (N_9875,N_9552,N_9559);
and U9876 (N_9876,N_9610,N_9706);
nor U9877 (N_9877,N_9731,N_9662);
xnor U9878 (N_9878,N_9644,N_9527);
nor U9879 (N_9879,N_9686,N_9547);
nand U9880 (N_9880,N_9622,N_9621);
xor U9881 (N_9881,N_9695,N_9749);
and U9882 (N_9882,N_9724,N_9700);
xor U9883 (N_9883,N_9566,N_9739);
nand U9884 (N_9884,N_9650,N_9711);
nand U9885 (N_9885,N_9580,N_9638);
nor U9886 (N_9886,N_9526,N_9669);
xor U9887 (N_9887,N_9536,N_9720);
or U9888 (N_9888,N_9725,N_9570);
xor U9889 (N_9889,N_9544,N_9621);
and U9890 (N_9890,N_9505,N_9521);
xnor U9891 (N_9891,N_9728,N_9531);
nor U9892 (N_9892,N_9701,N_9567);
or U9893 (N_9893,N_9539,N_9666);
xnor U9894 (N_9894,N_9706,N_9541);
nor U9895 (N_9895,N_9597,N_9732);
and U9896 (N_9896,N_9666,N_9673);
xnor U9897 (N_9897,N_9552,N_9518);
xor U9898 (N_9898,N_9505,N_9734);
nand U9899 (N_9899,N_9748,N_9701);
xnor U9900 (N_9900,N_9546,N_9611);
nand U9901 (N_9901,N_9713,N_9636);
xnor U9902 (N_9902,N_9639,N_9564);
or U9903 (N_9903,N_9504,N_9533);
xnor U9904 (N_9904,N_9588,N_9643);
or U9905 (N_9905,N_9611,N_9713);
or U9906 (N_9906,N_9612,N_9680);
xnor U9907 (N_9907,N_9746,N_9609);
and U9908 (N_9908,N_9740,N_9647);
nor U9909 (N_9909,N_9681,N_9723);
and U9910 (N_9910,N_9712,N_9552);
nor U9911 (N_9911,N_9605,N_9688);
nor U9912 (N_9912,N_9613,N_9576);
xnor U9913 (N_9913,N_9709,N_9504);
or U9914 (N_9914,N_9696,N_9586);
and U9915 (N_9915,N_9707,N_9615);
nand U9916 (N_9916,N_9648,N_9598);
nand U9917 (N_9917,N_9728,N_9611);
nor U9918 (N_9918,N_9590,N_9612);
xnor U9919 (N_9919,N_9589,N_9701);
nor U9920 (N_9920,N_9555,N_9582);
nor U9921 (N_9921,N_9503,N_9601);
nand U9922 (N_9922,N_9742,N_9608);
and U9923 (N_9923,N_9560,N_9699);
and U9924 (N_9924,N_9747,N_9658);
nand U9925 (N_9925,N_9552,N_9575);
nor U9926 (N_9926,N_9731,N_9519);
xor U9927 (N_9927,N_9705,N_9557);
nand U9928 (N_9928,N_9728,N_9679);
nand U9929 (N_9929,N_9511,N_9582);
nor U9930 (N_9930,N_9549,N_9708);
xor U9931 (N_9931,N_9712,N_9746);
xnor U9932 (N_9932,N_9607,N_9657);
nand U9933 (N_9933,N_9656,N_9556);
nor U9934 (N_9934,N_9577,N_9586);
nand U9935 (N_9935,N_9502,N_9701);
or U9936 (N_9936,N_9626,N_9542);
nand U9937 (N_9937,N_9721,N_9593);
and U9938 (N_9938,N_9669,N_9564);
or U9939 (N_9939,N_9668,N_9656);
nand U9940 (N_9940,N_9547,N_9614);
xnor U9941 (N_9941,N_9546,N_9606);
xor U9942 (N_9942,N_9533,N_9643);
or U9943 (N_9943,N_9624,N_9507);
or U9944 (N_9944,N_9592,N_9540);
xnor U9945 (N_9945,N_9630,N_9730);
nor U9946 (N_9946,N_9616,N_9580);
and U9947 (N_9947,N_9619,N_9612);
xnor U9948 (N_9948,N_9722,N_9649);
and U9949 (N_9949,N_9747,N_9503);
nor U9950 (N_9950,N_9664,N_9689);
and U9951 (N_9951,N_9725,N_9745);
xor U9952 (N_9952,N_9543,N_9672);
or U9953 (N_9953,N_9664,N_9575);
or U9954 (N_9954,N_9598,N_9626);
nor U9955 (N_9955,N_9725,N_9661);
nand U9956 (N_9956,N_9502,N_9742);
nand U9957 (N_9957,N_9707,N_9743);
or U9958 (N_9958,N_9743,N_9520);
nand U9959 (N_9959,N_9677,N_9664);
and U9960 (N_9960,N_9672,N_9576);
nand U9961 (N_9961,N_9613,N_9693);
xor U9962 (N_9962,N_9535,N_9546);
nand U9963 (N_9963,N_9664,N_9656);
and U9964 (N_9964,N_9518,N_9625);
nor U9965 (N_9965,N_9553,N_9597);
nor U9966 (N_9966,N_9502,N_9714);
or U9967 (N_9967,N_9714,N_9593);
and U9968 (N_9968,N_9583,N_9507);
and U9969 (N_9969,N_9566,N_9633);
nand U9970 (N_9970,N_9738,N_9620);
and U9971 (N_9971,N_9560,N_9733);
and U9972 (N_9972,N_9626,N_9511);
and U9973 (N_9973,N_9619,N_9534);
nor U9974 (N_9974,N_9506,N_9518);
and U9975 (N_9975,N_9528,N_9582);
and U9976 (N_9976,N_9665,N_9591);
xnor U9977 (N_9977,N_9713,N_9518);
and U9978 (N_9978,N_9552,N_9561);
or U9979 (N_9979,N_9704,N_9571);
or U9980 (N_9980,N_9682,N_9615);
xor U9981 (N_9981,N_9519,N_9539);
nor U9982 (N_9982,N_9703,N_9709);
nand U9983 (N_9983,N_9622,N_9651);
xnor U9984 (N_9984,N_9586,N_9657);
xnor U9985 (N_9985,N_9532,N_9541);
and U9986 (N_9986,N_9591,N_9661);
or U9987 (N_9987,N_9694,N_9613);
and U9988 (N_9988,N_9705,N_9704);
and U9989 (N_9989,N_9567,N_9696);
xnor U9990 (N_9990,N_9683,N_9628);
and U9991 (N_9991,N_9617,N_9729);
nor U9992 (N_9992,N_9674,N_9696);
xnor U9993 (N_9993,N_9565,N_9712);
or U9994 (N_9994,N_9506,N_9679);
xnor U9995 (N_9995,N_9600,N_9698);
xnor U9996 (N_9996,N_9533,N_9644);
nor U9997 (N_9997,N_9592,N_9655);
or U9998 (N_9998,N_9633,N_9502);
xor U9999 (N_9999,N_9652,N_9508);
or U10000 (N_10000,N_9846,N_9893);
or U10001 (N_10001,N_9778,N_9949);
nor U10002 (N_10002,N_9871,N_9892);
xor U10003 (N_10003,N_9944,N_9856);
nand U10004 (N_10004,N_9844,N_9936);
or U10005 (N_10005,N_9837,N_9888);
nand U10006 (N_10006,N_9793,N_9884);
nor U10007 (N_10007,N_9972,N_9809);
and U10008 (N_10008,N_9927,N_9901);
nor U10009 (N_10009,N_9882,N_9783);
xnor U10010 (N_10010,N_9770,N_9920);
nor U10011 (N_10011,N_9833,N_9913);
and U10012 (N_10012,N_9995,N_9762);
and U10013 (N_10013,N_9885,N_9801);
or U10014 (N_10014,N_9996,N_9835);
xnor U10015 (N_10015,N_9953,N_9755);
nand U10016 (N_10016,N_9786,N_9759);
nor U10017 (N_10017,N_9829,N_9946);
nand U10018 (N_10018,N_9758,N_9806);
nor U10019 (N_10019,N_9990,N_9854);
and U10020 (N_10020,N_9814,N_9872);
and U10021 (N_10021,N_9940,N_9779);
and U10022 (N_10022,N_9878,N_9766);
nand U10023 (N_10023,N_9803,N_9942);
and U10024 (N_10024,N_9889,N_9817);
xnor U10025 (N_10025,N_9869,N_9947);
nand U10026 (N_10026,N_9902,N_9794);
nand U10027 (N_10027,N_9954,N_9767);
nor U10028 (N_10028,N_9780,N_9932);
nand U10029 (N_10029,N_9825,N_9973);
nor U10030 (N_10030,N_9977,N_9867);
nand U10031 (N_10031,N_9978,N_9799);
nand U10032 (N_10032,N_9997,N_9836);
nor U10033 (N_10033,N_9800,N_9787);
xnor U10034 (N_10034,N_9841,N_9812);
nand U10035 (N_10035,N_9959,N_9979);
xnor U10036 (N_10036,N_9850,N_9782);
nor U10037 (N_10037,N_9987,N_9811);
and U10038 (N_10038,N_9980,N_9756);
nor U10039 (N_10039,N_9813,N_9776);
and U10040 (N_10040,N_9823,N_9769);
or U10041 (N_10041,N_9914,N_9816);
nor U10042 (N_10042,N_9956,N_9789);
nand U10043 (N_10043,N_9880,N_9802);
and U10044 (N_10044,N_9847,N_9763);
nor U10045 (N_10045,N_9788,N_9858);
or U10046 (N_10046,N_9772,N_9895);
nand U10047 (N_10047,N_9851,N_9752);
and U10048 (N_10048,N_9790,N_9898);
and U10049 (N_10049,N_9815,N_9773);
and U10050 (N_10050,N_9848,N_9921);
nor U10051 (N_10051,N_9900,N_9839);
nand U10052 (N_10052,N_9751,N_9826);
and U10053 (N_10053,N_9899,N_9985);
xnor U10054 (N_10054,N_9834,N_9970);
and U10055 (N_10055,N_9916,N_9988);
or U10056 (N_10056,N_9964,N_9868);
xor U10057 (N_10057,N_9966,N_9943);
xnor U10058 (N_10058,N_9765,N_9984);
xor U10059 (N_10059,N_9863,N_9866);
nand U10060 (N_10060,N_9860,N_9975);
and U10061 (N_10061,N_9937,N_9753);
xor U10062 (N_10062,N_9785,N_9967);
nor U10063 (N_10063,N_9821,N_9935);
or U10064 (N_10064,N_9962,N_9853);
or U10065 (N_10065,N_9781,N_9915);
or U10066 (N_10066,N_9971,N_9929);
and U10067 (N_10067,N_9777,N_9881);
xor U10068 (N_10068,N_9912,N_9931);
nor U10069 (N_10069,N_9883,N_9859);
or U10070 (N_10070,N_9796,N_9930);
or U10071 (N_10071,N_9792,N_9941);
and U10072 (N_10072,N_9819,N_9795);
and U10073 (N_10073,N_9879,N_9831);
or U10074 (N_10074,N_9807,N_9905);
or U10075 (N_10075,N_9952,N_9945);
nor U10076 (N_10076,N_9963,N_9897);
nand U10077 (N_10077,N_9827,N_9857);
nand U10078 (N_10078,N_9986,N_9838);
and U10079 (N_10079,N_9870,N_9958);
and U10080 (N_10080,N_9861,N_9849);
nand U10081 (N_10081,N_9994,N_9993);
nor U10082 (N_10082,N_9976,N_9891);
or U10083 (N_10083,N_9922,N_9761);
and U10084 (N_10084,N_9918,N_9887);
xnor U10085 (N_10085,N_9896,N_9852);
nand U10086 (N_10086,N_9928,N_9910);
xnor U10087 (N_10087,N_9934,N_9804);
or U10088 (N_10088,N_9998,N_9757);
nand U10089 (N_10089,N_9890,N_9864);
and U10090 (N_10090,N_9808,N_9810);
nor U10091 (N_10091,N_9797,N_9775);
or U10092 (N_10092,N_9992,N_9950);
nand U10093 (N_10093,N_9798,N_9760);
and U10094 (N_10094,N_9965,N_9843);
or U10095 (N_10095,N_9768,N_9818);
and U10096 (N_10096,N_9989,N_9906);
nand U10097 (N_10097,N_9924,N_9771);
nand U10098 (N_10098,N_9862,N_9917);
nor U10099 (N_10099,N_9999,N_9982);
or U10100 (N_10100,N_9911,N_9894);
and U10101 (N_10101,N_9832,N_9877);
nor U10102 (N_10102,N_9842,N_9764);
nand U10103 (N_10103,N_9750,N_9991);
xor U10104 (N_10104,N_9907,N_9820);
or U10105 (N_10105,N_9983,N_9754);
nand U10106 (N_10106,N_9865,N_9791);
and U10107 (N_10107,N_9925,N_9908);
or U10108 (N_10108,N_9873,N_9961);
and U10109 (N_10109,N_9969,N_9875);
nor U10110 (N_10110,N_9981,N_9828);
or U10111 (N_10111,N_9830,N_9974);
nand U10112 (N_10112,N_9939,N_9926);
nor U10113 (N_10113,N_9774,N_9886);
xnor U10114 (N_10114,N_9923,N_9968);
nor U10115 (N_10115,N_9903,N_9822);
or U10116 (N_10116,N_9874,N_9840);
and U10117 (N_10117,N_9845,N_9948);
and U10118 (N_10118,N_9938,N_9876);
xnor U10119 (N_10119,N_9904,N_9951);
and U10120 (N_10120,N_9919,N_9784);
nand U10121 (N_10121,N_9955,N_9960);
or U10122 (N_10122,N_9909,N_9824);
and U10123 (N_10123,N_9933,N_9957);
or U10124 (N_10124,N_9805,N_9855);
nor U10125 (N_10125,N_9927,N_9970);
and U10126 (N_10126,N_9991,N_9799);
nand U10127 (N_10127,N_9954,N_9792);
xnor U10128 (N_10128,N_9829,N_9869);
xor U10129 (N_10129,N_9996,N_9838);
or U10130 (N_10130,N_9838,N_9813);
xnor U10131 (N_10131,N_9931,N_9858);
nand U10132 (N_10132,N_9997,N_9835);
nor U10133 (N_10133,N_9776,N_9770);
nand U10134 (N_10134,N_9953,N_9873);
or U10135 (N_10135,N_9775,N_9859);
or U10136 (N_10136,N_9885,N_9921);
nor U10137 (N_10137,N_9894,N_9854);
and U10138 (N_10138,N_9986,N_9866);
xnor U10139 (N_10139,N_9787,N_9892);
nand U10140 (N_10140,N_9753,N_9843);
or U10141 (N_10141,N_9782,N_9940);
or U10142 (N_10142,N_9755,N_9872);
xor U10143 (N_10143,N_9921,N_9980);
and U10144 (N_10144,N_9947,N_9750);
xnor U10145 (N_10145,N_9777,N_9959);
nor U10146 (N_10146,N_9753,N_9839);
or U10147 (N_10147,N_9930,N_9756);
nand U10148 (N_10148,N_9770,N_9805);
nand U10149 (N_10149,N_9993,N_9969);
xor U10150 (N_10150,N_9846,N_9821);
nand U10151 (N_10151,N_9876,N_9881);
or U10152 (N_10152,N_9761,N_9960);
nor U10153 (N_10153,N_9790,N_9888);
nand U10154 (N_10154,N_9861,N_9769);
or U10155 (N_10155,N_9865,N_9969);
and U10156 (N_10156,N_9811,N_9985);
and U10157 (N_10157,N_9797,N_9996);
and U10158 (N_10158,N_9942,N_9974);
or U10159 (N_10159,N_9768,N_9944);
nor U10160 (N_10160,N_9915,N_9892);
nor U10161 (N_10161,N_9878,N_9812);
nand U10162 (N_10162,N_9852,N_9914);
nor U10163 (N_10163,N_9895,N_9969);
xnor U10164 (N_10164,N_9829,N_9944);
nand U10165 (N_10165,N_9846,N_9938);
or U10166 (N_10166,N_9891,N_9793);
nor U10167 (N_10167,N_9773,N_9930);
nand U10168 (N_10168,N_9782,N_9886);
nand U10169 (N_10169,N_9807,N_9788);
nand U10170 (N_10170,N_9960,N_9941);
xor U10171 (N_10171,N_9794,N_9844);
and U10172 (N_10172,N_9897,N_9991);
and U10173 (N_10173,N_9775,N_9968);
nor U10174 (N_10174,N_9997,N_9916);
and U10175 (N_10175,N_9856,N_9934);
or U10176 (N_10176,N_9818,N_9906);
or U10177 (N_10177,N_9759,N_9869);
xor U10178 (N_10178,N_9772,N_9877);
and U10179 (N_10179,N_9778,N_9864);
xnor U10180 (N_10180,N_9816,N_9930);
xnor U10181 (N_10181,N_9934,N_9868);
nor U10182 (N_10182,N_9973,N_9963);
xor U10183 (N_10183,N_9869,N_9930);
xnor U10184 (N_10184,N_9930,N_9782);
or U10185 (N_10185,N_9820,N_9844);
nor U10186 (N_10186,N_9985,N_9789);
xor U10187 (N_10187,N_9940,N_9835);
and U10188 (N_10188,N_9878,N_9991);
and U10189 (N_10189,N_9810,N_9772);
xnor U10190 (N_10190,N_9773,N_9762);
nor U10191 (N_10191,N_9763,N_9807);
xnor U10192 (N_10192,N_9858,N_9755);
nor U10193 (N_10193,N_9985,N_9762);
and U10194 (N_10194,N_9787,N_9921);
or U10195 (N_10195,N_9922,N_9960);
nand U10196 (N_10196,N_9940,N_9978);
xor U10197 (N_10197,N_9807,N_9830);
and U10198 (N_10198,N_9960,N_9927);
and U10199 (N_10199,N_9965,N_9903);
xor U10200 (N_10200,N_9771,N_9825);
xor U10201 (N_10201,N_9956,N_9897);
or U10202 (N_10202,N_9751,N_9930);
nand U10203 (N_10203,N_9775,N_9953);
nand U10204 (N_10204,N_9868,N_9839);
xor U10205 (N_10205,N_9809,N_9926);
nor U10206 (N_10206,N_9842,N_9949);
nand U10207 (N_10207,N_9890,N_9880);
xnor U10208 (N_10208,N_9888,N_9982);
nand U10209 (N_10209,N_9962,N_9862);
nand U10210 (N_10210,N_9974,N_9805);
nor U10211 (N_10211,N_9759,N_9813);
xnor U10212 (N_10212,N_9949,N_9784);
or U10213 (N_10213,N_9884,N_9759);
xnor U10214 (N_10214,N_9837,N_9770);
or U10215 (N_10215,N_9910,N_9878);
nor U10216 (N_10216,N_9934,N_9850);
nand U10217 (N_10217,N_9860,N_9825);
xor U10218 (N_10218,N_9940,N_9753);
nor U10219 (N_10219,N_9762,N_9848);
and U10220 (N_10220,N_9903,N_9802);
nand U10221 (N_10221,N_9855,N_9923);
nor U10222 (N_10222,N_9772,N_9992);
and U10223 (N_10223,N_9966,N_9896);
and U10224 (N_10224,N_9968,N_9951);
nand U10225 (N_10225,N_9885,N_9819);
and U10226 (N_10226,N_9828,N_9956);
nor U10227 (N_10227,N_9955,N_9877);
xnor U10228 (N_10228,N_9782,N_9798);
and U10229 (N_10229,N_9803,N_9994);
nand U10230 (N_10230,N_9954,N_9930);
xnor U10231 (N_10231,N_9986,N_9890);
nand U10232 (N_10232,N_9954,N_9980);
nor U10233 (N_10233,N_9852,N_9880);
nor U10234 (N_10234,N_9927,N_9903);
and U10235 (N_10235,N_9974,N_9877);
nand U10236 (N_10236,N_9898,N_9750);
nand U10237 (N_10237,N_9945,N_9811);
or U10238 (N_10238,N_9914,N_9966);
nor U10239 (N_10239,N_9961,N_9933);
nand U10240 (N_10240,N_9770,N_9778);
and U10241 (N_10241,N_9966,N_9932);
and U10242 (N_10242,N_9858,N_9889);
xnor U10243 (N_10243,N_9858,N_9816);
or U10244 (N_10244,N_9930,N_9993);
or U10245 (N_10245,N_9970,N_9946);
xnor U10246 (N_10246,N_9762,N_9958);
xnor U10247 (N_10247,N_9980,N_9901);
nand U10248 (N_10248,N_9946,N_9969);
or U10249 (N_10249,N_9933,N_9856);
and U10250 (N_10250,N_10235,N_10060);
nand U10251 (N_10251,N_10143,N_10201);
nand U10252 (N_10252,N_10059,N_10030);
xnor U10253 (N_10253,N_10189,N_10109);
and U10254 (N_10254,N_10118,N_10022);
or U10255 (N_10255,N_10131,N_10199);
nor U10256 (N_10256,N_10073,N_10037);
and U10257 (N_10257,N_10188,N_10048);
nand U10258 (N_10258,N_10012,N_10116);
nand U10259 (N_10259,N_10089,N_10176);
xor U10260 (N_10260,N_10168,N_10238);
nor U10261 (N_10261,N_10098,N_10130);
nor U10262 (N_10262,N_10039,N_10181);
nor U10263 (N_10263,N_10107,N_10007);
nand U10264 (N_10264,N_10160,N_10074);
xnor U10265 (N_10265,N_10186,N_10206);
nor U10266 (N_10266,N_10207,N_10113);
nor U10267 (N_10267,N_10018,N_10159);
and U10268 (N_10268,N_10142,N_10240);
nor U10269 (N_10269,N_10080,N_10071);
nand U10270 (N_10270,N_10145,N_10185);
and U10271 (N_10271,N_10121,N_10064);
or U10272 (N_10272,N_10191,N_10173);
xor U10273 (N_10273,N_10163,N_10100);
or U10274 (N_10274,N_10182,N_10213);
or U10275 (N_10275,N_10230,N_10128);
or U10276 (N_10276,N_10090,N_10237);
xor U10277 (N_10277,N_10187,N_10190);
or U10278 (N_10278,N_10157,N_10070);
and U10279 (N_10279,N_10141,N_10239);
xor U10280 (N_10280,N_10097,N_10156);
nand U10281 (N_10281,N_10249,N_10151);
and U10282 (N_10282,N_10148,N_10241);
nand U10283 (N_10283,N_10171,N_10021);
nor U10284 (N_10284,N_10027,N_10177);
xor U10285 (N_10285,N_10219,N_10038);
xnor U10286 (N_10286,N_10132,N_10155);
xnor U10287 (N_10287,N_10029,N_10023);
xor U10288 (N_10288,N_10138,N_10035);
or U10289 (N_10289,N_10224,N_10081);
xnor U10290 (N_10290,N_10125,N_10003);
nand U10291 (N_10291,N_10193,N_10002);
xnor U10292 (N_10292,N_10026,N_10153);
nor U10293 (N_10293,N_10036,N_10056);
nand U10294 (N_10294,N_10149,N_10072);
or U10295 (N_10295,N_10045,N_10229);
nor U10296 (N_10296,N_10042,N_10222);
xor U10297 (N_10297,N_10198,N_10015);
nor U10298 (N_10298,N_10079,N_10046);
nand U10299 (N_10299,N_10167,N_10053);
and U10300 (N_10300,N_10106,N_10008);
and U10301 (N_10301,N_10117,N_10087);
xnor U10302 (N_10302,N_10068,N_10103);
xnor U10303 (N_10303,N_10040,N_10051);
nor U10304 (N_10304,N_10088,N_10127);
or U10305 (N_10305,N_10005,N_10013);
and U10306 (N_10306,N_10172,N_10119);
and U10307 (N_10307,N_10179,N_10228);
or U10308 (N_10308,N_10028,N_10223);
nand U10309 (N_10309,N_10055,N_10178);
and U10310 (N_10310,N_10140,N_10114);
xnor U10311 (N_10311,N_10120,N_10031);
nand U10312 (N_10312,N_10104,N_10184);
nor U10313 (N_10313,N_10204,N_10047);
or U10314 (N_10314,N_10208,N_10244);
or U10315 (N_10315,N_10233,N_10212);
nor U10316 (N_10316,N_10086,N_10075);
xor U10317 (N_10317,N_10112,N_10058);
nor U10318 (N_10318,N_10062,N_10115);
or U10319 (N_10319,N_10209,N_10243);
nand U10320 (N_10320,N_10041,N_10099);
and U10321 (N_10321,N_10033,N_10101);
nor U10322 (N_10322,N_10245,N_10218);
or U10323 (N_10323,N_10225,N_10093);
nor U10324 (N_10324,N_10010,N_10221);
or U10325 (N_10325,N_10226,N_10082);
or U10326 (N_10326,N_10154,N_10247);
nand U10327 (N_10327,N_10017,N_10144);
or U10328 (N_10328,N_10111,N_10078);
nor U10329 (N_10329,N_10236,N_10009);
xor U10330 (N_10330,N_10083,N_10126);
or U10331 (N_10331,N_10217,N_10000);
or U10332 (N_10332,N_10211,N_10183);
nor U10333 (N_10333,N_10020,N_10162);
and U10334 (N_10334,N_10085,N_10246);
xor U10335 (N_10335,N_10076,N_10195);
nor U10336 (N_10336,N_10161,N_10052);
nand U10337 (N_10337,N_10014,N_10050);
nand U10338 (N_10338,N_10006,N_10092);
xnor U10339 (N_10339,N_10066,N_10122);
or U10340 (N_10340,N_10044,N_10049);
and U10341 (N_10341,N_10032,N_10174);
nor U10342 (N_10342,N_10096,N_10166);
xnor U10343 (N_10343,N_10150,N_10242);
xor U10344 (N_10344,N_10108,N_10170);
xor U10345 (N_10345,N_10011,N_10061);
nand U10346 (N_10346,N_10203,N_10210);
nor U10347 (N_10347,N_10063,N_10137);
nor U10348 (N_10348,N_10084,N_10019);
nand U10349 (N_10349,N_10077,N_10110);
nor U10350 (N_10350,N_10133,N_10043);
or U10351 (N_10351,N_10227,N_10102);
and U10352 (N_10352,N_10024,N_10129);
nand U10353 (N_10353,N_10094,N_10069);
nand U10354 (N_10354,N_10146,N_10147);
and U10355 (N_10355,N_10202,N_10123);
nor U10356 (N_10356,N_10091,N_10065);
nand U10357 (N_10357,N_10067,N_10234);
and U10358 (N_10358,N_10025,N_10216);
nor U10359 (N_10359,N_10004,N_10192);
xnor U10360 (N_10360,N_10124,N_10194);
or U10361 (N_10361,N_10016,N_10164);
xnor U10362 (N_10362,N_10214,N_10165);
nand U10363 (N_10363,N_10220,N_10034);
or U10364 (N_10364,N_10232,N_10057);
and U10365 (N_10365,N_10197,N_10135);
or U10366 (N_10366,N_10200,N_10175);
nor U10367 (N_10367,N_10158,N_10095);
nand U10368 (N_10368,N_10180,N_10231);
xnor U10369 (N_10369,N_10105,N_10134);
and U10370 (N_10370,N_10139,N_10205);
nor U10371 (N_10371,N_10196,N_10001);
or U10372 (N_10372,N_10152,N_10215);
or U10373 (N_10373,N_10169,N_10054);
xnor U10374 (N_10374,N_10136,N_10248);
nor U10375 (N_10375,N_10039,N_10192);
and U10376 (N_10376,N_10111,N_10098);
nor U10377 (N_10377,N_10119,N_10098);
and U10378 (N_10378,N_10217,N_10021);
or U10379 (N_10379,N_10146,N_10101);
nor U10380 (N_10380,N_10229,N_10110);
nor U10381 (N_10381,N_10155,N_10038);
nor U10382 (N_10382,N_10223,N_10102);
nand U10383 (N_10383,N_10118,N_10097);
or U10384 (N_10384,N_10170,N_10070);
or U10385 (N_10385,N_10157,N_10159);
nand U10386 (N_10386,N_10113,N_10238);
xor U10387 (N_10387,N_10183,N_10012);
or U10388 (N_10388,N_10144,N_10197);
nor U10389 (N_10389,N_10044,N_10059);
xnor U10390 (N_10390,N_10169,N_10164);
or U10391 (N_10391,N_10048,N_10030);
nand U10392 (N_10392,N_10038,N_10025);
nor U10393 (N_10393,N_10020,N_10219);
xor U10394 (N_10394,N_10185,N_10106);
and U10395 (N_10395,N_10018,N_10191);
or U10396 (N_10396,N_10044,N_10050);
xnor U10397 (N_10397,N_10217,N_10133);
or U10398 (N_10398,N_10226,N_10125);
xnor U10399 (N_10399,N_10038,N_10017);
or U10400 (N_10400,N_10082,N_10053);
and U10401 (N_10401,N_10109,N_10031);
xnor U10402 (N_10402,N_10165,N_10225);
nor U10403 (N_10403,N_10017,N_10101);
nor U10404 (N_10404,N_10039,N_10077);
or U10405 (N_10405,N_10005,N_10194);
nand U10406 (N_10406,N_10215,N_10239);
and U10407 (N_10407,N_10013,N_10245);
or U10408 (N_10408,N_10158,N_10133);
xnor U10409 (N_10409,N_10166,N_10192);
nor U10410 (N_10410,N_10048,N_10005);
or U10411 (N_10411,N_10054,N_10051);
or U10412 (N_10412,N_10232,N_10098);
xnor U10413 (N_10413,N_10060,N_10158);
or U10414 (N_10414,N_10206,N_10038);
nand U10415 (N_10415,N_10105,N_10055);
and U10416 (N_10416,N_10018,N_10068);
and U10417 (N_10417,N_10164,N_10161);
or U10418 (N_10418,N_10002,N_10192);
nor U10419 (N_10419,N_10138,N_10147);
or U10420 (N_10420,N_10070,N_10214);
nand U10421 (N_10421,N_10156,N_10230);
nand U10422 (N_10422,N_10017,N_10060);
xnor U10423 (N_10423,N_10078,N_10053);
xnor U10424 (N_10424,N_10214,N_10140);
nand U10425 (N_10425,N_10248,N_10071);
nor U10426 (N_10426,N_10013,N_10074);
or U10427 (N_10427,N_10085,N_10210);
xnor U10428 (N_10428,N_10185,N_10144);
nor U10429 (N_10429,N_10117,N_10164);
or U10430 (N_10430,N_10230,N_10085);
and U10431 (N_10431,N_10126,N_10091);
or U10432 (N_10432,N_10211,N_10067);
xnor U10433 (N_10433,N_10016,N_10154);
xor U10434 (N_10434,N_10233,N_10077);
xnor U10435 (N_10435,N_10055,N_10248);
xor U10436 (N_10436,N_10200,N_10205);
nor U10437 (N_10437,N_10013,N_10070);
nor U10438 (N_10438,N_10033,N_10202);
or U10439 (N_10439,N_10087,N_10032);
xor U10440 (N_10440,N_10058,N_10070);
nand U10441 (N_10441,N_10101,N_10085);
nand U10442 (N_10442,N_10224,N_10113);
or U10443 (N_10443,N_10087,N_10080);
nand U10444 (N_10444,N_10136,N_10078);
and U10445 (N_10445,N_10003,N_10180);
or U10446 (N_10446,N_10230,N_10018);
xnor U10447 (N_10447,N_10070,N_10100);
nand U10448 (N_10448,N_10157,N_10117);
nand U10449 (N_10449,N_10009,N_10231);
nor U10450 (N_10450,N_10192,N_10213);
nand U10451 (N_10451,N_10182,N_10138);
and U10452 (N_10452,N_10022,N_10081);
and U10453 (N_10453,N_10009,N_10115);
and U10454 (N_10454,N_10007,N_10112);
nor U10455 (N_10455,N_10145,N_10129);
nand U10456 (N_10456,N_10195,N_10012);
and U10457 (N_10457,N_10124,N_10069);
and U10458 (N_10458,N_10055,N_10042);
or U10459 (N_10459,N_10216,N_10190);
nor U10460 (N_10460,N_10245,N_10018);
and U10461 (N_10461,N_10161,N_10224);
xor U10462 (N_10462,N_10074,N_10003);
xnor U10463 (N_10463,N_10018,N_10092);
or U10464 (N_10464,N_10133,N_10237);
or U10465 (N_10465,N_10116,N_10239);
or U10466 (N_10466,N_10144,N_10036);
and U10467 (N_10467,N_10154,N_10028);
or U10468 (N_10468,N_10081,N_10129);
nor U10469 (N_10469,N_10112,N_10167);
nor U10470 (N_10470,N_10242,N_10027);
nand U10471 (N_10471,N_10100,N_10195);
xor U10472 (N_10472,N_10136,N_10243);
nor U10473 (N_10473,N_10111,N_10112);
xnor U10474 (N_10474,N_10141,N_10111);
or U10475 (N_10475,N_10193,N_10234);
nand U10476 (N_10476,N_10045,N_10143);
xor U10477 (N_10477,N_10038,N_10123);
or U10478 (N_10478,N_10163,N_10023);
or U10479 (N_10479,N_10209,N_10157);
nand U10480 (N_10480,N_10023,N_10148);
xor U10481 (N_10481,N_10232,N_10008);
nand U10482 (N_10482,N_10217,N_10190);
and U10483 (N_10483,N_10006,N_10130);
xor U10484 (N_10484,N_10124,N_10026);
and U10485 (N_10485,N_10092,N_10201);
nor U10486 (N_10486,N_10043,N_10027);
or U10487 (N_10487,N_10158,N_10080);
and U10488 (N_10488,N_10143,N_10128);
nor U10489 (N_10489,N_10006,N_10115);
nand U10490 (N_10490,N_10097,N_10088);
or U10491 (N_10491,N_10027,N_10186);
or U10492 (N_10492,N_10013,N_10008);
nor U10493 (N_10493,N_10214,N_10179);
nand U10494 (N_10494,N_10170,N_10118);
and U10495 (N_10495,N_10140,N_10240);
nand U10496 (N_10496,N_10066,N_10162);
or U10497 (N_10497,N_10023,N_10006);
nand U10498 (N_10498,N_10105,N_10139);
or U10499 (N_10499,N_10247,N_10186);
or U10500 (N_10500,N_10379,N_10380);
nand U10501 (N_10501,N_10472,N_10260);
nand U10502 (N_10502,N_10401,N_10368);
or U10503 (N_10503,N_10491,N_10271);
nand U10504 (N_10504,N_10262,N_10376);
nor U10505 (N_10505,N_10484,N_10342);
and U10506 (N_10506,N_10335,N_10453);
nor U10507 (N_10507,N_10256,N_10333);
or U10508 (N_10508,N_10359,N_10433);
nand U10509 (N_10509,N_10413,N_10253);
nand U10510 (N_10510,N_10305,N_10277);
nand U10511 (N_10511,N_10340,N_10264);
xor U10512 (N_10512,N_10479,N_10452);
or U10513 (N_10513,N_10393,N_10279);
and U10514 (N_10514,N_10434,N_10346);
and U10515 (N_10515,N_10411,N_10469);
xor U10516 (N_10516,N_10427,N_10475);
or U10517 (N_10517,N_10307,N_10332);
nand U10518 (N_10518,N_10292,N_10490);
and U10519 (N_10519,N_10323,N_10425);
or U10520 (N_10520,N_10295,N_10441);
or U10521 (N_10521,N_10481,N_10331);
nand U10522 (N_10522,N_10317,N_10275);
and U10523 (N_10523,N_10325,N_10255);
xnor U10524 (N_10524,N_10440,N_10384);
nand U10525 (N_10525,N_10437,N_10254);
xnor U10526 (N_10526,N_10355,N_10352);
nor U10527 (N_10527,N_10451,N_10337);
xnor U10528 (N_10528,N_10497,N_10311);
nand U10529 (N_10529,N_10374,N_10415);
nor U10530 (N_10530,N_10424,N_10477);
nand U10531 (N_10531,N_10408,N_10321);
and U10532 (N_10532,N_10280,N_10308);
nand U10533 (N_10533,N_10349,N_10302);
nor U10534 (N_10534,N_10460,N_10318);
nor U10535 (N_10535,N_10371,N_10465);
nor U10536 (N_10536,N_10285,N_10466);
xor U10537 (N_10537,N_10429,N_10485);
and U10538 (N_10538,N_10357,N_10334);
and U10539 (N_10539,N_10489,N_10320);
or U10540 (N_10540,N_10404,N_10328);
nand U10541 (N_10541,N_10499,N_10467);
and U10542 (N_10542,N_10369,N_10430);
nor U10543 (N_10543,N_10306,N_10496);
or U10544 (N_10544,N_10373,N_10381);
nand U10545 (N_10545,N_10388,N_10417);
xnor U10546 (N_10546,N_10398,N_10399);
xnor U10547 (N_10547,N_10319,N_10382);
and U10548 (N_10548,N_10290,N_10314);
or U10549 (N_10549,N_10468,N_10299);
and U10550 (N_10550,N_10488,N_10310);
nand U10551 (N_10551,N_10351,N_10495);
or U10552 (N_10552,N_10461,N_10397);
or U10553 (N_10553,N_10406,N_10298);
nor U10554 (N_10554,N_10365,N_10400);
or U10555 (N_10555,N_10312,N_10267);
nand U10556 (N_10556,N_10356,N_10487);
or U10557 (N_10557,N_10265,N_10392);
nor U10558 (N_10558,N_10385,N_10478);
nand U10559 (N_10559,N_10421,N_10370);
xor U10560 (N_10560,N_10445,N_10486);
xnor U10561 (N_10561,N_10316,N_10268);
nand U10562 (N_10562,N_10309,N_10284);
nor U10563 (N_10563,N_10471,N_10418);
nand U10564 (N_10564,N_10294,N_10455);
and U10565 (N_10565,N_10446,N_10358);
or U10566 (N_10566,N_10396,N_10444);
or U10567 (N_10567,N_10270,N_10407);
and U10568 (N_10568,N_10426,N_10326);
and U10569 (N_10569,N_10283,N_10322);
and U10570 (N_10570,N_10409,N_10313);
nand U10571 (N_10571,N_10324,N_10339);
xor U10572 (N_10572,N_10329,N_10482);
nand U10573 (N_10573,N_10301,N_10416);
and U10574 (N_10574,N_10344,N_10273);
nor U10575 (N_10575,N_10272,N_10412);
or U10576 (N_10576,N_10443,N_10338);
nand U10577 (N_10577,N_10269,N_10330);
or U10578 (N_10578,N_10493,N_10422);
xor U10579 (N_10579,N_10251,N_10473);
xor U10580 (N_10580,N_10350,N_10442);
xnor U10581 (N_10581,N_10492,N_10304);
xnor U10582 (N_10582,N_10431,N_10456);
and U10583 (N_10583,N_10447,N_10293);
and U10584 (N_10584,N_10390,N_10449);
and U10585 (N_10585,N_10383,N_10367);
or U10586 (N_10586,N_10448,N_10375);
nor U10587 (N_10587,N_10363,N_10439);
or U10588 (N_10588,N_10366,N_10494);
nor U10589 (N_10589,N_10336,N_10347);
nand U10590 (N_10590,N_10303,N_10377);
and U10591 (N_10591,N_10459,N_10389);
nand U10592 (N_10592,N_10345,N_10454);
nand U10593 (N_10593,N_10354,N_10315);
or U10594 (N_10594,N_10257,N_10483);
nand U10595 (N_10595,N_10364,N_10395);
nor U10596 (N_10596,N_10435,N_10378);
nor U10597 (N_10597,N_10361,N_10480);
and U10598 (N_10598,N_10372,N_10348);
xor U10599 (N_10599,N_10281,N_10410);
xnor U10600 (N_10600,N_10464,N_10394);
and U10601 (N_10601,N_10402,N_10438);
nor U10602 (N_10602,N_10450,N_10288);
or U10603 (N_10603,N_10476,N_10414);
or U10604 (N_10604,N_10282,N_10258);
and U10605 (N_10605,N_10498,N_10252);
xnor U10606 (N_10606,N_10250,N_10297);
and U10607 (N_10607,N_10300,N_10462);
nor U10608 (N_10608,N_10353,N_10463);
or U10609 (N_10609,N_10327,N_10405);
nand U10610 (N_10610,N_10432,N_10391);
nor U10611 (N_10611,N_10287,N_10403);
nand U10612 (N_10612,N_10362,N_10263);
xnor U10613 (N_10613,N_10419,N_10289);
nand U10614 (N_10614,N_10458,N_10423);
or U10615 (N_10615,N_10278,N_10387);
or U10616 (N_10616,N_10296,N_10474);
and U10617 (N_10617,N_10436,N_10470);
and U10618 (N_10618,N_10343,N_10360);
or U10619 (N_10619,N_10259,N_10291);
or U10620 (N_10620,N_10276,N_10428);
nand U10621 (N_10621,N_10286,N_10457);
and U10622 (N_10622,N_10386,N_10261);
and U10623 (N_10623,N_10420,N_10274);
nand U10624 (N_10624,N_10341,N_10266);
or U10625 (N_10625,N_10378,N_10452);
or U10626 (N_10626,N_10267,N_10286);
nand U10627 (N_10627,N_10297,N_10290);
or U10628 (N_10628,N_10483,N_10275);
xor U10629 (N_10629,N_10309,N_10461);
or U10630 (N_10630,N_10412,N_10344);
and U10631 (N_10631,N_10379,N_10276);
and U10632 (N_10632,N_10299,N_10362);
or U10633 (N_10633,N_10301,N_10300);
nor U10634 (N_10634,N_10332,N_10309);
xnor U10635 (N_10635,N_10365,N_10464);
nor U10636 (N_10636,N_10298,N_10270);
or U10637 (N_10637,N_10310,N_10332);
and U10638 (N_10638,N_10263,N_10373);
and U10639 (N_10639,N_10460,N_10389);
xnor U10640 (N_10640,N_10311,N_10308);
or U10641 (N_10641,N_10486,N_10281);
nand U10642 (N_10642,N_10397,N_10475);
and U10643 (N_10643,N_10347,N_10448);
nand U10644 (N_10644,N_10304,N_10319);
and U10645 (N_10645,N_10296,N_10441);
nor U10646 (N_10646,N_10485,N_10497);
nor U10647 (N_10647,N_10488,N_10369);
and U10648 (N_10648,N_10374,N_10260);
nor U10649 (N_10649,N_10256,N_10293);
or U10650 (N_10650,N_10485,N_10459);
nor U10651 (N_10651,N_10298,N_10318);
nand U10652 (N_10652,N_10307,N_10348);
xor U10653 (N_10653,N_10306,N_10321);
xnor U10654 (N_10654,N_10473,N_10253);
or U10655 (N_10655,N_10475,N_10388);
and U10656 (N_10656,N_10475,N_10312);
and U10657 (N_10657,N_10407,N_10299);
nand U10658 (N_10658,N_10395,N_10360);
nor U10659 (N_10659,N_10281,N_10266);
and U10660 (N_10660,N_10298,N_10294);
xor U10661 (N_10661,N_10260,N_10332);
and U10662 (N_10662,N_10371,N_10329);
xor U10663 (N_10663,N_10255,N_10482);
or U10664 (N_10664,N_10459,N_10407);
xor U10665 (N_10665,N_10302,N_10435);
nand U10666 (N_10666,N_10492,N_10478);
or U10667 (N_10667,N_10328,N_10385);
or U10668 (N_10668,N_10437,N_10471);
nand U10669 (N_10669,N_10402,N_10342);
xor U10670 (N_10670,N_10454,N_10427);
nor U10671 (N_10671,N_10276,N_10424);
xnor U10672 (N_10672,N_10369,N_10404);
xor U10673 (N_10673,N_10397,N_10316);
xor U10674 (N_10674,N_10262,N_10252);
or U10675 (N_10675,N_10436,N_10325);
or U10676 (N_10676,N_10342,N_10299);
xnor U10677 (N_10677,N_10337,N_10453);
nand U10678 (N_10678,N_10391,N_10270);
nand U10679 (N_10679,N_10274,N_10407);
nand U10680 (N_10680,N_10414,N_10481);
nand U10681 (N_10681,N_10401,N_10329);
nor U10682 (N_10682,N_10382,N_10272);
xnor U10683 (N_10683,N_10265,N_10481);
and U10684 (N_10684,N_10339,N_10409);
nor U10685 (N_10685,N_10436,N_10401);
nand U10686 (N_10686,N_10429,N_10450);
nor U10687 (N_10687,N_10437,N_10334);
nor U10688 (N_10688,N_10283,N_10412);
nand U10689 (N_10689,N_10486,N_10429);
nor U10690 (N_10690,N_10426,N_10338);
nand U10691 (N_10691,N_10304,N_10263);
nor U10692 (N_10692,N_10301,N_10469);
or U10693 (N_10693,N_10338,N_10495);
xnor U10694 (N_10694,N_10277,N_10307);
nor U10695 (N_10695,N_10337,N_10285);
or U10696 (N_10696,N_10363,N_10399);
xor U10697 (N_10697,N_10395,N_10354);
nor U10698 (N_10698,N_10452,N_10484);
xor U10699 (N_10699,N_10463,N_10420);
nor U10700 (N_10700,N_10312,N_10291);
xor U10701 (N_10701,N_10452,N_10466);
nand U10702 (N_10702,N_10424,N_10399);
xor U10703 (N_10703,N_10273,N_10293);
nor U10704 (N_10704,N_10250,N_10328);
or U10705 (N_10705,N_10496,N_10265);
or U10706 (N_10706,N_10389,N_10412);
xor U10707 (N_10707,N_10343,N_10465);
nand U10708 (N_10708,N_10409,N_10327);
nor U10709 (N_10709,N_10440,N_10428);
and U10710 (N_10710,N_10482,N_10352);
and U10711 (N_10711,N_10271,N_10435);
and U10712 (N_10712,N_10298,N_10487);
xor U10713 (N_10713,N_10433,N_10449);
xor U10714 (N_10714,N_10420,N_10465);
or U10715 (N_10715,N_10271,N_10398);
xor U10716 (N_10716,N_10423,N_10297);
nor U10717 (N_10717,N_10337,N_10416);
nand U10718 (N_10718,N_10269,N_10285);
and U10719 (N_10719,N_10467,N_10318);
nand U10720 (N_10720,N_10354,N_10275);
xnor U10721 (N_10721,N_10302,N_10369);
or U10722 (N_10722,N_10407,N_10433);
nor U10723 (N_10723,N_10255,N_10309);
nor U10724 (N_10724,N_10466,N_10258);
nand U10725 (N_10725,N_10316,N_10348);
xor U10726 (N_10726,N_10271,N_10350);
nor U10727 (N_10727,N_10478,N_10479);
nand U10728 (N_10728,N_10279,N_10487);
and U10729 (N_10729,N_10326,N_10352);
xnor U10730 (N_10730,N_10431,N_10454);
or U10731 (N_10731,N_10296,N_10398);
or U10732 (N_10732,N_10291,N_10390);
xnor U10733 (N_10733,N_10368,N_10384);
or U10734 (N_10734,N_10400,N_10480);
or U10735 (N_10735,N_10284,N_10445);
nand U10736 (N_10736,N_10391,N_10464);
nand U10737 (N_10737,N_10429,N_10272);
xnor U10738 (N_10738,N_10324,N_10362);
nor U10739 (N_10739,N_10385,N_10427);
nor U10740 (N_10740,N_10314,N_10302);
nand U10741 (N_10741,N_10358,N_10398);
nor U10742 (N_10742,N_10259,N_10433);
nor U10743 (N_10743,N_10421,N_10488);
or U10744 (N_10744,N_10282,N_10401);
xor U10745 (N_10745,N_10469,N_10433);
or U10746 (N_10746,N_10407,N_10341);
xor U10747 (N_10747,N_10424,N_10371);
and U10748 (N_10748,N_10488,N_10293);
nor U10749 (N_10749,N_10458,N_10330);
or U10750 (N_10750,N_10569,N_10501);
and U10751 (N_10751,N_10676,N_10540);
nand U10752 (N_10752,N_10570,N_10648);
or U10753 (N_10753,N_10673,N_10576);
xor U10754 (N_10754,N_10607,N_10524);
and U10755 (N_10755,N_10675,N_10630);
nand U10756 (N_10756,N_10668,N_10639);
or U10757 (N_10757,N_10691,N_10579);
xor U10758 (N_10758,N_10530,N_10554);
or U10759 (N_10759,N_10637,N_10694);
nand U10760 (N_10760,N_10535,N_10660);
nor U10761 (N_10761,N_10713,N_10533);
or U10762 (N_10762,N_10517,N_10651);
xor U10763 (N_10763,N_10539,N_10584);
nand U10764 (N_10764,N_10697,N_10632);
xor U10765 (N_10765,N_10730,N_10585);
nor U10766 (N_10766,N_10559,N_10596);
nor U10767 (N_10767,N_10729,N_10724);
or U10768 (N_10768,N_10736,N_10598);
and U10769 (N_10769,N_10706,N_10507);
nor U10770 (N_10770,N_10746,N_10709);
nand U10771 (N_10771,N_10518,N_10555);
nand U10772 (N_10772,N_10710,N_10722);
nor U10773 (N_10773,N_10522,N_10695);
xor U10774 (N_10774,N_10642,N_10603);
and U10775 (N_10775,N_10707,N_10574);
xnor U10776 (N_10776,N_10657,N_10726);
and U10777 (N_10777,N_10600,N_10666);
nor U10778 (N_10778,N_10593,N_10728);
nand U10779 (N_10779,N_10635,N_10616);
or U10780 (N_10780,N_10590,N_10514);
nand U10781 (N_10781,N_10725,N_10690);
nor U10782 (N_10782,N_10580,N_10696);
or U10783 (N_10783,N_10638,N_10715);
nand U10784 (N_10784,N_10571,N_10620);
nor U10785 (N_10785,N_10738,N_10688);
nand U10786 (N_10786,N_10528,N_10609);
or U10787 (N_10787,N_10604,N_10739);
xor U10788 (N_10788,N_10625,N_10599);
and U10789 (N_10789,N_10672,N_10536);
or U10790 (N_10790,N_10512,N_10747);
nand U10791 (N_10791,N_10602,N_10653);
xnor U10792 (N_10792,N_10683,N_10506);
xnor U10793 (N_10793,N_10595,N_10669);
xnor U10794 (N_10794,N_10572,N_10526);
and U10795 (N_10795,N_10628,N_10698);
or U10796 (N_10796,N_10741,N_10684);
xor U10797 (N_10797,N_10671,N_10723);
or U10798 (N_10798,N_10640,N_10682);
and U10799 (N_10799,N_10558,N_10742);
and U10800 (N_10800,N_10662,N_10619);
xor U10801 (N_10801,N_10677,N_10568);
nand U10802 (N_10802,N_10613,N_10615);
and U10803 (N_10803,N_10541,N_10537);
xnor U10804 (N_10804,N_10521,N_10550);
nor U10805 (N_10805,N_10745,N_10608);
nor U10806 (N_10806,N_10611,N_10551);
and U10807 (N_10807,N_10655,N_10610);
and U10808 (N_10808,N_10534,N_10678);
or U10809 (N_10809,N_10646,N_10502);
or U10810 (N_10810,N_10544,N_10553);
nor U10811 (N_10811,N_10703,N_10636);
nand U10812 (N_10812,N_10542,N_10546);
nand U10813 (N_10813,N_10622,N_10563);
or U10814 (N_10814,N_10547,N_10699);
or U10815 (N_10815,N_10689,N_10665);
xor U10816 (N_10816,N_10740,N_10661);
xor U10817 (N_10817,N_10508,N_10700);
and U10818 (N_10818,N_10647,N_10679);
and U10819 (N_10819,N_10606,N_10500);
or U10820 (N_10820,N_10548,N_10749);
and U10821 (N_10821,N_10591,N_10721);
and U10822 (N_10822,N_10618,N_10664);
nand U10823 (N_10823,N_10650,N_10531);
and U10824 (N_10824,N_10624,N_10513);
or U10825 (N_10825,N_10523,N_10543);
or U10826 (N_10826,N_10581,N_10589);
nand U10827 (N_10827,N_10538,N_10505);
or U10828 (N_10828,N_10711,N_10532);
and U10829 (N_10829,N_10716,N_10621);
xnor U10830 (N_10830,N_10734,N_10744);
xnor U10831 (N_10831,N_10519,N_10549);
nor U10832 (N_10832,N_10633,N_10614);
or U10833 (N_10833,N_10562,N_10516);
nand U10834 (N_10834,N_10561,N_10634);
or U10835 (N_10835,N_10718,N_10737);
nor U10836 (N_10836,N_10731,N_10708);
nand U10837 (N_10837,N_10605,N_10582);
xnor U10838 (N_10838,N_10556,N_10626);
nand U10839 (N_10839,N_10680,N_10504);
and U10840 (N_10840,N_10681,N_10586);
xnor U10841 (N_10841,N_10617,N_10527);
or U10842 (N_10842,N_10525,N_10674);
nand U10843 (N_10843,N_10503,N_10656);
and U10844 (N_10844,N_10641,N_10667);
nand U10845 (N_10845,N_10601,N_10658);
nand U10846 (N_10846,N_10597,N_10652);
and U10847 (N_10847,N_10645,N_10663);
or U10848 (N_10848,N_10623,N_10631);
nand U10849 (N_10849,N_10727,N_10685);
nor U10850 (N_10850,N_10515,N_10687);
or U10851 (N_10851,N_10545,N_10575);
nand U10852 (N_10852,N_10704,N_10686);
xnor U10853 (N_10853,N_10705,N_10701);
xor U10854 (N_10854,N_10612,N_10567);
or U10855 (N_10855,N_10693,N_10643);
xnor U10856 (N_10856,N_10712,N_10557);
or U10857 (N_10857,N_10654,N_10573);
xor U10858 (N_10858,N_10592,N_10733);
xor U10859 (N_10859,N_10510,N_10529);
and U10860 (N_10860,N_10644,N_10564);
nand U10861 (N_10861,N_10629,N_10748);
nor U10862 (N_10862,N_10649,N_10565);
and U10863 (N_10863,N_10520,N_10587);
or U10864 (N_10864,N_10594,N_10566);
or U10865 (N_10865,N_10743,N_10717);
xor U10866 (N_10866,N_10714,N_10627);
and U10867 (N_10867,N_10732,N_10720);
nand U10868 (N_10868,N_10583,N_10719);
xnor U10869 (N_10869,N_10588,N_10692);
and U10870 (N_10870,N_10578,N_10735);
and U10871 (N_10871,N_10702,N_10552);
nor U10872 (N_10872,N_10511,N_10560);
xnor U10873 (N_10873,N_10509,N_10670);
nor U10874 (N_10874,N_10577,N_10659);
nand U10875 (N_10875,N_10690,N_10737);
and U10876 (N_10876,N_10536,N_10557);
nand U10877 (N_10877,N_10514,N_10743);
or U10878 (N_10878,N_10595,N_10591);
xnor U10879 (N_10879,N_10579,N_10614);
or U10880 (N_10880,N_10516,N_10615);
xor U10881 (N_10881,N_10702,N_10567);
or U10882 (N_10882,N_10538,N_10726);
nor U10883 (N_10883,N_10592,N_10680);
or U10884 (N_10884,N_10530,N_10559);
or U10885 (N_10885,N_10647,N_10584);
nand U10886 (N_10886,N_10692,N_10712);
xor U10887 (N_10887,N_10686,N_10599);
xor U10888 (N_10888,N_10539,N_10609);
nor U10889 (N_10889,N_10704,N_10712);
nor U10890 (N_10890,N_10625,N_10527);
nand U10891 (N_10891,N_10649,N_10712);
xor U10892 (N_10892,N_10572,N_10588);
nor U10893 (N_10893,N_10691,N_10648);
nand U10894 (N_10894,N_10579,N_10625);
nor U10895 (N_10895,N_10671,N_10630);
xnor U10896 (N_10896,N_10571,N_10581);
nand U10897 (N_10897,N_10545,N_10587);
nand U10898 (N_10898,N_10682,N_10716);
or U10899 (N_10899,N_10674,N_10709);
nor U10900 (N_10900,N_10677,N_10659);
xnor U10901 (N_10901,N_10553,N_10719);
or U10902 (N_10902,N_10731,N_10648);
nor U10903 (N_10903,N_10657,N_10737);
or U10904 (N_10904,N_10661,N_10686);
and U10905 (N_10905,N_10704,N_10668);
xor U10906 (N_10906,N_10528,N_10653);
nand U10907 (N_10907,N_10687,N_10567);
xnor U10908 (N_10908,N_10642,N_10626);
nor U10909 (N_10909,N_10721,N_10518);
nor U10910 (N_10910,N_10502,N_10587);
and U10911 (N_10911,N_10624,N_10542);
nand U10912 (N_10912,N_10549,N_10701);
xnor U10913 (N_10913,N_10667,N_10726);
xor U10914 (N_10914,N_10558,N_10581);
nand U10915 (N_10915,N_10664,N_10586);
xnor U10916 (N_10916,N_10526,N_10685);
nor U10917 (N_10917,N_10707,N_10629);
nand U10918 (N_10918,N_10579,N_10617);
or U10919 (N_10919,N_10565,N_10643);
or U10920 (N_10920,N_10653,N_10593);
and U10921 (N_10921,N_10610,N_10617);
nand U10922 (N_10922,N_10507,N_10587);
nand U10923 (N_10923,N_10552,N_10703);
xor U10924 (N_10924,N_10627,N_10550);
nand U10925 (N_10925,N_10635,N_10544);
nand U10926 (N_10926,N_10646,N_10702);
and U10927 (N_10927,N_10664,N_10523);
xor U10928 (N_10928,N_10647,N_10590);
nand U10929 (N_10929,N_10737,N_10709);
and U10930 (N_10930,N_10641,N_10648);
or U10931 (N_10931,N_10540,N_10632);
or U10932 (N_10932,N_10690,N_10592);
nor U10933 (N_10933,N_10711,N_10539);
or U10934 (N_10934,N_10599,N_10698);
and U10935 (N_10935,N_10562,N_10658);
and U10936 (N_10936,N_10717,N_10667);
and U10937 (N_10937,N_10622,N_10707);
nor U10938 (N_10938,N_10514,N_10578);
and U10939 (N_10939,N_10697,N_10504);
xor U10940 (N_10940,N_10526,N_10674);
nor U10941 (N_10941,N_10569,N_10541);
nand U10942 (N_10942,N_10704,N_10577);
xor U10943 (N_10943,N_10562,N_10712);
xor U10944 (N_10944,N_10599,N_10527);
nand U10945 (N_10945,N_10640,N_10510);
xnor U10946 (N_10946,N_10700,N_10686);
nor U10947 (N_10947,N_10543,N_10606);
xnor U10948 (N_10948,N_10571,N_10622);
nand U10949 (N_10949,N_10653,N_10568);
nand U10950 (N_10950,N_10680,N_10510);
or U10951 (N_10951,N_10578,N_10625);
or U10952 (N_10952,N_10697,N_10506);
xor U10953 (N_10953,N_10501,N_10594);
or U10954 (N_10954,N_10701,N_10541);
and U10955 (N_10955,N_10589,N_10683);
xor U10956 (N_10956,N_10649,N_10618);
or U10957 (N_10957,N_10637,N_10677);
or U10958 (N_10958,N_10676,N_10724);
xor U10959 (N_10959,N_10719,N_10710);
and U10960 (N_10960,N_10516,N_10509);
nor U10961 (N_10961,N_10544,N_10581);
nor U10962 (N_10962,N_10687,N_10593);
nand U10963 (N_10963,N_10685,N_10707);
or U10964 (N_10964,N_10609,N_10735);
nand U10965 (N_10965,N_10583,N_10630);
xor U10966 (N_10966,N_10638,N_10713);
xor U10967 (N_10967,N_10507,N_10637);
or U10968 (N_10968,N_10662,N_10715);
xor U10969 (N_10969,N_10725,N_10616);
nand U10970 (N_10970,N_10664,N_10747);
xor U10971 (N_10971,N_10738,N_10675);
nor U10972 (N_10972,N_10697,N_10591);
or U10973 (N_10973,N_10681,N_10656);
nand U10974 (N_10974,N_10661,N_10536);
nor U10975 (N_10975,N_10571,N_10549);
nor U10976 (N_10976,N_10575,N_10607);
xor U10977 (N_10977,N_10741,N_10705);
or U10978 (N_10978,N_10557,N_10595);
or U10979 (N_10979,N_10669,N_10690);
and U10980 (N_10980,N_10567,N_10719);
or U10981 (N_10981,N_10516,N_10603);
or U10982 (N_10982,N_10544,N_10503);
xor U10983 (N_10983,N_10727,N_10745);
nand U10984 (N_10984,N_10717,N_10524);
and U10985 (N_10985,N_10640,N_10591);
and U10986 (N_10986,N_10738,N_10512);
and U10987 (N_10987,N_10560,N_10683);
nor U10988 (N_10988,N_10722,N_10561);
nand U10989 (N_10989,N_10697,N_10736);
xor U10990 (N_10990,N_10653,N_10709);
and U10991 (N_10991,N_10654,N_10720);
nor U10992 (N_10992,N_10681,N_10590);
and U10993 (N_10993,N_10656,N_10550);
nor U10994 (N_10994,N_10741,N_10566);
and U10995 (N_10995,N_10661,N_10726);
or U10996 (N_10996,N_10675,N_10659);
nand U10997 (N_10997,N_10640,N_10632);
or U10998 (N_10998,N_10604,N_10661);
and U10999 (N_10999,N_10532,N_10511);
and U11000 (N_11000,N_10869,N_10878);
nor U11001 (N_11001,N_10818,N_10904);
nand U11002 (N_11002,N_10919,N_10996);
or U11003 (N_11003,N_10935,N_10837);
and U11004 (N_11004,N_10756,N_10801);
xor U11005 (N_11005,N_10841,N_10856);
or U11006 (N_11006,N_10782,N_10967);
and U11007 (N_11007,N_10848,N_10961);
or U11008 (N_11008,N_10951,N_10854);
xnor U11009 (N_11009,N_10865,N_10930);
xor U11010 (N_11010,N_10948,N_10777);
nand U11011 (N_11011,N_10830,N_10914);
nand U11012 (N_11012,N_10866,N_10792);
and U11013 (N_11013,N_10879,N_10763);
and U11014 (N_11014,N_10903,N_10773);
xnor U11015 (N_11015,N_10981,N_10892);
xnor U11016 (N_11016,N_10891,N_10895);
nor U11017 (N_11017,N_10827,N_10889);
and U11018 (N_11018,N_10970,N_10906);
or U11019 (N_11019,N_10885,N_10832);
nor U11020 (N_11020,N_10765,N_10983);
nor U11021 (N_11021,N_10780,N_10882);
xnor U11022 (N_11022,N_10787,N_10873);
nand U11023 (N_11023,N_10993,N_10942);
xnor U11024 (N_11024,N_10809,N_10868);
and U11025 (N_11025,N_10846,N_10950);
or U11026 (N_11026,N_10959,N_10867);
xnor U11027 (N_11027,N_10766,N_10929);
nor U11028 (N_11028,N_10984,N_10875);
xor U11029 (N_11029,N_10994,N_10898);
and U11030 (N_11030,N_10877,N_10933);
or U11031 (N_11031,N_10833,N_10793);
nor U11032 (N_11032,N_10852,N_10907);
nor U11033 (N_11033,N_10938,N_10963);
xor U11034 (N_11034,N_10776,N_10811);
and U11035 (N_11035,N_10843,N_10954);
and U11036 (N_11036,N_10976,N_10971);
and U11037 (N_11037,N_10939,N_10855);
nand U11038 (N_11038,N_10902,N_10824);
or U11039 (N_11039,N_10803,N_10760);
and U11040 (N_11040,N_10778,N_10813);
and U11041 (N_11041,N_10806,N_10952);
nand U11042 (N_11042,N_10761,N_10943);
nor U11043 (N_11043,N_10884,N_10928);
and U11044 (N_11044,N_10800,N_10759);
or U11045 (N_11045,N_10945,N_10853);
and U11046 (N_11046,N_10874,N_10931);
nor U11047 (N_11047,N_10839,N_10913);
nand U11048 (N_11048,N_10962,N_10888);
nand U11049 (N_11049,N_10775,N_10819);
nor U11050 (N_11050,N_10966,N_10815);
nor U11051 (N_11051,N_10774,N_10975);
nand U11052 (N_11052,N_10785,N_10861);
nand U11053 (N_11053,N_10829,N_10847);
nand U11054 (N_11054,N_10956,N_10890);
nand U11055 (N_11055,N_10880,N_10934);
xor U11056 (N_11056,N_10751,N_10754);
nand U11057 (N_11057,N_10864,N_10978);
or U11058 (N_11058,N_10810,N_10923);
nand U11059 (N_11059,N_10937,N_10805);
nor U11060 (N_11060,N_10784,N_10905);
xnor U11061 (N_11061,N_10990,N_10860);
xnor U11062 (N_11062,N_10842,N_10998);
and U11063 (N_11063,N_10767,N_10851);
and U11064 (N_11064,N_10790,N_10821);
and U11065 (N_11065,N_10758,N_10881);
nand U11066 (N_11066,N_10850,N_10883);
nand U11067 (N_11067,N_10953,N_10755);
nor U11068 (N_11068,N_10922,N_10900);
xor U11069 (N_11069,N_10909,N_10828);
or U11070 (N_11070,N_10849,N_10845);
nor U11071 (N_11071,N_10901,N_10831);
and U11072 (N_11072,N_10757,N_10964);
xor U11073 (N_11073,N_10908,N_10958);
nor U11074 (N_11074,N_10858,N_10789);
nor U11075 (N_11075,N_10995,N_10750);
xnor U11076 (N_11076,N_10817,N_10944);
nor U11077 (N_11077,N_10988,N_10791);
or U11078 (N_11078,N_10752,N_10921);
xnor U11079 (N_11079,N_10985,N_10987);
nor U11080 (N_11080,N_10816,N_10910);
xnor U11081 (N_11081,N_10834,N_10764);
nor U11082 (N_11082,N_10808,N_10781);
and U11083 (N_11083,N_10926,N_10917);
xnor U11084 (N_11084,N_10798,N_10822);
xnor U11085 (N_11085,N_10823,N_10783);
nor U11086 (N_11086,N_10974,N_10863);
xor U11087 (N_11087,N_10804,N_10940);
nand U11088 (N_11088,N_10912,N_10826);
nor U11089 (N_11089,N_10941,N_10911);
nand U11090 (N_11090,N_10949,N_10986);
nor U11091 (N_11091,N_10965,N_10980);
nor U11092 (N_11092,N_10899,N_10972);
or U11093 (N_11093,N_10862,N_10968);
and U11094 (N_11094,N_10796,N_10807);
xor U11095 (N_11095,N_10835,N_10871);
and U11096 (N_11096,N_10897,N_10838);
and U11097 (N_11097,N_10957,N_10915);
nor U11098 (N_11098,N_10927,N_10999);
or U11099 (N_11099,N_10870,N_10946);
xor U11100 (N_11100,N_10925,N_10802);
and U11101 (N_11101,N_10947,N_10795);
and U11102 (N_11102,N_10794,N_10893);
nor U11103 (N_11103,N_10812,N_10969);
nor U11104 (N_11104,N_10762,N_10876);
xor U11105 (N_11105,N_10786,N_10857);
nand U11106 (N_11106,N_10779,N_10814);
and U11107 (N_11107,N_10955,N_10887);
xnor U11108 (N_11108,N_10973,N_10894);
and U11109 (N_11109,N_10872,N_10825);
or U11110 (N_11110,N_10753,N_10924);
and U11111 (N_11111,N_10997,N_10992);
nand U11112 (N_11112,N_10836,N_10844);
or U11113 (N_11113,N_10788,N_10982);
or U11114 (N_11114,N_10920,N_10896);
nor U11115 (N_11115,N_10840,N_10771);
nand U11116 (N_11116,N_10979,N_10859);
xor U11117 (N_11117,N_10989,N_10977);
nor U11118 (N_11118,N_10991,N_10918);
nor U11119 (N_11119,N_10820,N_10932);
nand U11120 (N_11120,N_10799,N_10797);
or U11121 (N_11121,N_10960,N_10916);
and U11122 (N_11122,N_10886,N_10769);
nor U11123 (N_11123,N_10768,N_10772);
nand U11124 (N_11124,N_10770,N_10936);
nand U11125 (N_11125,N_10986,N_10787);
nor U11126 (N_11126,N_10783,N_10912);
and U11127 (N_11127,N_10900,N_10934);
xnor U11128 (N_11128,N_10856,N_10978);
nand U11129 (N_11129,N_10840,N_10848);
and U11130 (N_11130,N_10880,N_10878);
and U11131 (N_11131,N_10839,N_10999);
or U11132 (N_11132,N_10980,N_10764);
nand U11133 (N_11133,N_10999,N_10892);
nand U11134 (N_11134,N_10798,N_10907);
nand U11135 (N_11135,N_10905,N_10762);
nor U11136 (N_11136,N_10784,N_10865);
xor U11137 (N_11137,N_10988,N_10803);
nor U11138 (N_11138,N_10899,N_10854);
or U11139 (N_11139,N_10792,N_10779);
xnor U11140 (N_11140,N_10792,N_10827);
nor U11141 (N_11141,N_10830,N_10810);
or U11142 (N_11142,N_10786,N_10908);
and U11143 (N_11143,N_10986,N_10997);
nand U11144 (N_11144,N_10824,N_10949);
nand U11145 (N_11145,N_10996,N_10803);
nand U11146 (N_11146,N_10953,N_10778);
and U11147 (N_11147,N_10987,N_10935);
nand U11148 (N_11148,N_10984,N_10767);
nand U11149 (N_11149,N_10861,N_10940);
or U11150 (N_11150,N_10789,N_10944);
nor U11151 (N_11151,N_10791,N_10910);
nand U11152 (N_11152,N_10936,N_10924);
nor U11153 (N_11153,N_10911,N_10917);
xnor U11154 (N_11154,N_10833,N_10766);
or U11155 (N_11155,N_10750,N_10913);
nand U11156 (N_11156,N_10926,N_10984);
xor U11157 (N_11157,N_10768,N_10975);
and U11158 (N_11158,N_10808,N_10754);
or U11159 (N_11159,N_10766,N_10874);
nand U11160 (N_11160,N_10798,N_10982);
xnor U11161 (N_11161,N_10800,N_10815);
and U11162 (N_11162,N_10981,N_10824);
and U11163 (N_11163,N_10931,N_10886);
xnor U11164 (N_11164,N_10761,N_10930);
nor U11165 (N_11165,N_10990,N_10807);
xor U11166 (N_11166,N_10958,N_10793);
nor U11167 (N_11167,N_10913,N_10842);
xnor U11168 (N_11168,N_10941,N_10874);
and U11169 (N_11169,N_10774,N_10981);
nor U11170 (N_11170,N_10810,N_10796);
and U11171 (N_11171,N_10836,N_10950);
nand U11172 (N_11172,N_10787,N_10779);
nand U11173 (N_11173,N_10932,N_10781);
nor U11174 (N_11174,N_10871,N_10904);
and U11175 (N_11175,N_10859,N_10816);
xor U11176 (N_11176,N_10778,N_10810);
and U11177 (N_11177,N_10807,N_10880);
nand U11178 (N_11178,N_10874,N_10906);
xor U11179 (N_11179,N_10841,N_10798);
or U11180 (N_11180,N_10934,N_10810);
xor U11181 (N_11181,N_10847,N_10921);
nand U11182 (N_11182,N_10952,N_10972);
nand U11183 (N_11183,N_10918,N_10822);
or U11184 (N_11184,N_10758,N_10915);
or U11185 (N_11185,N_10878,N_10930);
nand U11186 (N_11186,N_10752,N_10758);
and U11187 (N_11187,N_10927,N_10888);
or U11188 (N_11188,N_10844,N_10855);
and U11189 (N_11189,N_10808,N_10930);
or U11190 (N_11190,N_10851,N_10754);
or U11191 (N_11191,N_10915,N_10992);
or U11192 (N_11192,N_10940,N_10868);
and U11193 (N_11193,N_10964,N_10865);
and U11194 (N_11194,N_10830,N_10755);
xnor U11195 (N_11195,N_10906,N_10985);
xnor U11196 (N_11196,N_10803,N_10893);
or U11197 (N_11197,N_10851,N_10868);
nand U11198 (N_11198,N_10829,N_10927);
nor U11199 (N_11199,N_10913,N_10948);
nand U11200 (N_11200,N_10910,N_10992);
nand U11201 (N_11201,N_10827,N_10780);
or U11202 (N_11202,N_10956,N_10846);
nand U11203 (N_11203,N_10909,N_10880);
nand U11204 (N_11204,N_10846,N_10840);
and U11205 (N_11205,N_10869,N_10973);
nor U11206 (N_11206,N_10833,N_10843);
nand U11207 (N_11207,N_10905,N_10917);
xnor U11208 (N_11208,N_10945,N_10949);
nor U11209 (N_11209,N_10876,N_10788);
and U11210 (N_11210,N_10952,N_10779);
nor U11211 (N_11211,N_10767,N_10817);
nand U11212 (N_11212,N_10907,N_10809);
or U11213 (N_11213,N_10945,N_10790);
xnor U11214 (N_11214,N_10989,N_10966);
or U11215 (N_11215,N_10781,N_10956);
nor U11216 (N_11216,N_10922,N_10937);
and U11217 (N_11217,N_10750,N_10922);
nor U11218 (N_11218,N_10758,N_10966);
or U11219 (N_11219,N_10808,N_10839);
or U11220 (N_11220,N_10859,N_10949);
nand U11221 (N_11221,N_10855,N_10978);
nand U11222 (N_11222,N_10835,N_10919);
or U11223 (N_11223,N_10951,N_10813);
nand U11224 (N_11224,N_10857,N_10938);
nor U11225 (N_11225,N_10877,N_10884);
or U11226 (N_11226,N_10816,N_10990);
or U11227 (N_11227,N_10836,N_10941);
nand U11228 (N_11228,N_10897,N_10907);
xnor U11229 (N_11229,N_10895,N_10794);
xnor U11230 (N_11230,N_10828,N_10771);
nand U11231 (N_11231,N_10936,N_10766);
or U11232 (N_11232,N_10968,N_10944);
nand U11233 (N_11233,N_10813,N_10994);
and U11234 (N_11234,N_10938,N_10909);
nand U11235 (N_11235,N_10811,N_10928);
nand U11236 (N_11236,N_10858,N_10820);
or U11237 (N_11237,N_10988,N_10917);
nand U11238 (N_11238,N_10804,N_10830);
or U11239 (N_11239,N_10766,N_10786);
or U11240 (N_11240,N_10781,N_10817);
nand U11241 (N_11241,N_10887,N_10961);
nor U11242 (N_11242,N_10926,N_10955);
or U11243 (N_11243,N_10981,N_10791);
or U11244 (N_11244,N_10980,N_10853);
or U11245 (N_11245,N_10946,N_10844);
xnor U11246 (N_11246,N_10978,N_10778);
nor U11247 (N_11247,N_10857,N_10934);
or U11248 (N_11248,N_10807,N_10972);
nor U11249 (N_11249,N_10979,N_10817);
and U11250 (N_11250,N_11010,N_11194);
and U11251 (N_11251,N_11200,N_11238);
nand U11252 (N_11252,N_11123,N_11102);
or U11253 (N_11253,N_11049,N_11180);
xnor U11254 (N_11254,N_11205,N_11091);
and U11255 (N_11255,N_11115,N_11093);
and U11256 (N_11256,N_11177,N_11138);
nand U11257 (N_11257,N_11004,N_11192);
xor U11258 (N_11258,N_11080,N_11121);
nor U11259 (N_11259,N_11236,N_11202);
nor U11260 (N_11260,N_11197,N_11143);
xor U11261 (N_11261,N_11247,N_11246);
or U11262 (N_11262,N_11041,N_11022);
and U11263 (N_11263,N_11181,N_11075);
xnor U11264 (N_11264,N_11030,N_11243);
xnor U11265 (N_11265,N_11153,N_11056);
nor U11266 (N_11266,N_11150,N_11084);
nor U11267 (N_11267,N_11103,N_11191);
nand U11268 (N_11268,N_11064,N_11196);
nor U11269 (N_11269,N_11245,N_11066);
or U11270 (N_11270,N_11241,N_11040);
or U11271 (N_11271,N_11193,N_11171);
xnor U11272 (N_11272,N_11098,N_11059);
xor U11273 (N_11273,N_11104,N_11070);
nand U11274 (N_11274,N_11055,N_11020);
nor U11275 (N_11275,N_11231,N_11139);
nor U11276 (N_11276,N_11184,N_11152);
and U11277 (N_11277,N_11009,N_11097);
nand U11278 (N_11278,N_11134,N_11141);
and U11279 (N_11279,N_11175,N_11149);
nand U11280 (N_11280,N_11212,N_11240);
and U11281 (N_11281,N_11005,N_11229);
xor U11282 (N_11282,N_11248,N_11223);
xor U11283 (N_11283,N_11094,N_11233);
or U11284 (N_11284,N_11224,N_11169);
or U11285 (N_11285,N_11249,N_11081);
or U11286 (N_11286,N_11065,N_11086);
or U11287 (N_11287,N_11026,N_11018);
nor U11288 (N_11288,N_11222,N_11234);
xor U11289 (N_11289,N_11213,N_11237);
and U11290 (N_11290,N_11105,N_11019);
xor U11291 (N_11291,N_11045,N_11166);
and U11292 (N_11292,N_11118,N_11145);
nor U11293 (N_11293,N_11209,N_11101);
or U11294 (N_11294,N_11178,N_11012);
nor U11295 (N_11295,N_11034,N_11052);
nand U11296 (N_11296,N_11195,N_11095);
xor U11297 (N_11297,N_11244,N_11058);
nand U11298 (N_11298,N_11067,N_11179);
nand U11299 (N_11299,N_11161,N_11120);
nor U11300 (N_11300,N_11210,N_11000);
nand U11301 (N_11301,N_11219,N_11013);
nand U11302 (N_11302,N_11051,N_11140);
nor U11303 (N_11303,N_11016,N_11182);
or U11304 (N_11304,N_11111,N_11214);
and U11305 (N_11305,N_11142,N_11076);
nand U11306 (N_11306,N_11015,N_11239);
nand U11307 (N_11307,N_11036,N_11168);
nor U11308 (N_11308,N_11071,N_11227);
xor U11309 (N_11309,N_11176,N_11148);
or U11310 (N_11310,N_11037,N_11235);
nor U11311 (N_11311,N_11160,N_11083);
and U11312 (N_11312,N_11069,N_11156);
and U11313 (N_11313,N_11025,N_11100);
nand U11314 (N_11314,N_11198,N_11029);
and U11315 (N_11315,N_11003,N_11108);
and U11316 (N_11316,N_11035,N_11047);
and U11317 (N_11317,N_11216,N_11023);
or U11318 (N_11318,N_11057,N_11038);
xor U11319 (N_11319,N_11024,N_11014);
nor U11320 (N_11320,N_11221,N_11201);
nor U11321 (N_11321,N_11187,N_11125);
nand U11322 (N_11322,N_11068,N_11124);
or U11323 (N_11323,N_11033,N_11133);
or U11324 (N_11324,N_11131,N_11085);
xor U11325 (N_11325,N_11151,N_11117);
xnor U11326 (N_11326,N_11230,N_11112);
nor U11327 (N_11327,N_11174,N_11072);
and U11328 (N_11328,N_11220,N_11044);
or U11329 (N_11329,N_11113,N_11188);
nand U11330 (N_11330,N_11027,N_11048);
nor U11331 (N_11331,N_11136,N_11147);
or U11332 (N_11332,N_11021,N_11162);
nand U11333 (N_11333,N_11006,N_11031);
xor U11334 (N_11334,N_11228,N_11110);
nor U11335 (N_11335,N_11199,N_11099);
and U11336 (N_11336,N_11096,N_11116);
nor U11337 (N_11337,N_11060,N_11172);
and U11338 (N_11338,N_11167,N_11073);
nand U11339 (N_11339,N_11032,N_11135);
and U11340 (N_11340,N_11146,N_11046);
nand U11341 (N_11341,N_11232,N_11017);
nor U11342 (N_11342,N_11207,N_11144);
or U11343 (N_11343,N_11129,N_11119);
nor U11344 (N_11344,N_11092,N_11173);
xor U11345 (N_11345,N_11054,N_11164);
nor U11346 (N_11346,N_11002,N_11163);
and U11347 (N_11347,N_11225,N_11043);
xnor U11348 (N_11348,N_11215,N_11122);
nand U11349 (N_11349,N_11217,N_11042);
or U11350 (N_11350,N_11078,N_11132);
nand U11351 (N_11351,N_11208,N_11242);
and U11352 (N_11352,N_11206,N_11106);
nand U11353 (N_11353,N_11183,N_11090);
nor U11354 (N_11354,N_11226,N_11028);
xnor U11355 (N_11355,N_11061,N_11001);
xor U11356 (N_11356,N_11159,N_11203);
and U11357 (N_11357,N_11114,N_11082);
and U11358 (N_11358,N_11050,N_11077);
xnor U11359 (N_11359,N_11130,N_11039);
nor U11360 (N_11360,N_11088,N_11158);
xnor U11361 (N_11361,N_11185,N_11127);
or U11362 (N_11362,N_11126,N_11107);
nor U11363 (N_11363,N_11186,N_11011);
nand U11364 (N_11364,N_11074,N_11218);
nand U11365 (N_11365,N_11008,N_11155);
nand U11366 (N_11366,N_11087,N_11165);
xnor U11367 (N_11367,N_11079,N_11137);
and U11368 (N_11368,N_11157,N_11062);
and U11369 (N_11369,N_11204,N_11128);
or U11370 (N_11370,N_11189,N_11190);
or U11371 (N_11371,N_11170,N_11063);
nand U11372 (N_11372,N_11154,N_11089);
or U11373 (N_11373,N_11007,N_11211);
xnor U11374 (N_11374,N_11109,N_11053);
and U11375 (N_11375,N_11116,N_11046);
and U11376 (N_11376,N_11136,N_11052);
nor U11377 (N_11377,N_11010,N_11124);
nor U11378 (N_11378,N_11164,N_11246);
and U11379 (N_11379,N_11088,N_11050);
and U11380 (N_11380,N_11081,N_11027);
nor U11381 (N_11381,N_11134,N_11082);
nor U11382 (N_11382,N_11035,N_11126);
nor U11383 (N_11383,N_11161,N_11240);
nand U11384 (N_11384,N_11232,N_11234);
or U11385 (N_11385,N_11060,N_11167);
nand U11386 (N_11386,N_11227,N_11074);
and U11387 (N_11387,N_11168,N_11075);
nor U11388 (N_11388,N_11093,N_11026);
xnor U11389 (N_11389,N_11001,N_11239);
nor U11390 (N_11390,N_11047,N_11174);
and U11391 (N_11391,N_11065,N_11046);
or U11392 (N_11392,N_11108,N_11158);
xnor U11393 (N_11393,N_11159,N_11039);
or U11394 (N_11394,N_11165,N_11189);
or U11395 (N_11395,N_11047,N_11108);
xor U11396 (N_11396,N_11129,N_11197);
or U11397 (N_11397,N_11001,N_11129);
nand U11398 (N_11398,N_11074,N_11151);
nor U11399 (N_11399,N_11151,N_11034);
nand U11400 (N_11400,N_11034,N_11054);
nand U11401 (N_11401,N_11166,N_11103);
and U11402 (N_11402,N_11108,N_11044);
xor U11403 (N_11403,N_11044,N_11183);
nor U11404 (N_11404,N_11230,N_11152);
nand U11405 (N_11405,N_11040,N_11215);
and U11406 (N_11406,N_11125,N_11009);
xnor U11407 (N_11407,N_11084,N_11232);
nand U11408 (N_11408,N_11134,N_11061);
or U11409 (N_11409,N_11113,N_11128);
and U11410 (N_11410,N_11148,N_11005);
and U11411 (N_11411,N_11170,N_11098);
xnor U11412 (N_11412,N_11011,N_11167);
or U11413 (N_11413,N_11227,N_11142);
xnor U11414 (N_11414,N_11204,N_11150);
nand U11415 (N_11415,N_11244,N_11076);
and U11416 (N_11416,N_11234,N_11083);
and U11417 (N_11417,N_11129,N_11092);
and U11418 (N_11418,N_11042,N_11235);
nor U11419 (N_11419,N_11165,N_11017);
or U11420 (N_11420,N_11233,N_11009);
or U11421 (N_11421,N_11013,N_11143);
nor U11422 (N_11422,N_11030,N_11006);
and U11423 (N_11423,N_11058,N_11105);
nor U11424 (N_11424,N_11219,N_11119);
nand U11425 (N_11425,N_11155,N_11018);
and U11426 (N_11426,N_11136,N_11064);
and U11427 (N_11427,N_11241,N_11166);
nor U11428 (N_11428,N_11195,N_11020);
and U11429 (N_11429,N_11002,N_11020);
nand U11430 (N_11430,N_11074,N_11099);
or U11431 (N_11431,N_11070,N_11212);
or U11432 (N_11432,N_11182,N_11243);
nor U11433 (N_11433,N_11068,N_11130);
nand U11434 (N_11434,N_11006,N_11170);
xnor U11435 (N_11435,N_11040,N_11223);
or U11436 (N_11436,N_11109,N_11202);
and U11437 (N_11437,N_11097,N_11230);
nand U11438 (N_11438,N_11042,N_11141);
nand U11439 (N_11439,N_11131,N_11179);
nand U11440 (N_11440,N_11229,N_11077);
xor U11441 (N_11441,N_11114,N_11048);
and U11442 (N_11442,N_11190,N_11049);
or U11443 (N_11443,N_11213,N_11115);
nand U11444 (N_11444,N_11239,N_11117);
nor U11445 (N_11445,N_11166,N_11109);
xor U11446 (N_11446,N_11062,N_11178);
nand U11447 (N_11447,N_11210,N_11059);
nand U11448 (N_11448,N_11151,N_11146);
or U11449 (N_11449,N_11112,N_11027);
nor U11450 (N_11450,N_11144,N_11058);
nor U11451 (N_11451,N_11078,N_11114);
nand U11452 (N_11452,N_11151,N_11047);
nand U11453 (N_11453,N_11242,N_11222);
nor U11454 (N_11454,N_11013,N_11096);
and U11455 (N_11455,N_11006,N_11208);
or U11456 (N_11456,N_11000,N_11223);
nand U11457 (N_11457,N_11126,N_11147);
and U11458 (N_11458,N_11004,N_11065);
nand U11459 (N_11459,N_11227,N_11119);
nor U11460 (N_11460,N_11190,N_11121);
nor U11461 (N_11461,N_11245,N_11131);
nand U11462 (N_11462,N_11213,N_11203);
or U11463 (N_11463,N_11048,N_11239);
and U11464 (N_11464,N_11200,N_11125);
nand U11465 (N_11465,N_11059,N_11116);
nand U11466 (N_11466,N_11219,N_11017);
nand U11467 (N_11467,N_11096,N_11031);
nor U11468 (N_11468,N_11229,N_11145);
or U11469 (N_11469,N_11040,N_11166);
and U11470 (N_11470,N_11172,N_11232);
or U11471 (N_11471,N_11099,N_11130);
nor U11472 (N_11472,N_11164,N_11199);
or U11473 (N_11473,N_11046,N_11073);
or U11474 (N_11474,N_11201,N_11163);
nand U11475 (N_11475,N_11044,N_11158);
nand U11476 (N_11476,N_11085,N_11028);
xor U11477 (N_11477,N_11224,N_11071);
nand U11478 (N_11478,N_11028,N_11199);
nor U11479 (N_11479,N_11033,N_11231);
xor U11480 (N_11480,N_11225,N_11085);
nand U11481 (N_11481,N_11179,N_11039);
nor U11482 (N_11482,N_11118,N_11101);
or U11483 (N_11483,N_11212,N_11035);
and U11484 (N_11484,N_11208,N_11058);
xnor U11485 (N_11485,N_11097,N_11212);
or U11486 (N_11486,N_11230,N_11148);
xor U11487 (N_11487,N_11037,N_11125);
or U11488 (N_11488,N_11113,N_11085);
nand U11489 (N_11489,N_11197,N_11065);
nor U11490 (N_11490,N_11218,N_11215);
nand U11491 (N_11491,N_11137,N_11149);
and U11492 (N_11492,N_11224,N_11135);
nand U11493 (N_11493,N_11162,N_11201);
or U11494 (N_11494,N_11198,N_11045);
and U11495 (N_11495,N_11134,N_11140);
or U11496 (N_11496,N_11044,N_11067);
or U11497 (N_11497,N_11110,N_11185);
and U11498 (N_11498,N_11151,N_11134);
or U11499 (N_11499,N_11179,N_11114);
xnor U11500 (N_11500,N_11467,N_11313);
and U11501 (N_11501,N_11432,N_11488);
or U11502 (N_11502,N_11438,N_11357);
or U11503 (N_11503,N_11256,N_11382);
xor U11504 (N_11504,N_11307,N_11296);
nand U11505 (N_11505,N_11493,N_11352);
and U11506 (N_11506,N_11359,N_11370);
and U11507 (N_11507,N_11264,N_11287);
xor U11508 (N_11508,N_11441,N_11485);
nand U11509 (N_11509,N_11481,N_11402);
and U11510 (N_11510,N_11332,N_11430);
xnor U11511 (N_11511,N_11321,N_11305);
nor U11512 (N_11512,N_11339,N_11288);
nand U11513 (N_11513,N_11309,N_11335);
and U11514 (N_11514,N_11311,N_11409);
xnor U11515 (N_11515,N_11427,N_11297);
nand U11516 (N_11516,N_11363,N_11388);
nor U11517 (N_11517,N_11405,N_11385);
and U11518 (N_11518,N_11374,N_11389);
and U11519 (N_11519,N_11383,N_11443);
and U11520 (N_11520,N_11492,N_11324);
or U11521 (N_11521,N_11365,N_11487);
or U11522 (N_11522,N_11468,N_11377);
or U11523 (N_11523,N_11278,N_11449);
or U11524 (N_11524,N_11494,N_11428);
or U11525 (N_11525,N_11406,N_11390);
and U11526 (N_11526,N_11458,N_11445);
and U11527 (N_11527,N_11419,N_11403);
or U11528 (N_11528,N_11396,N_11275);
and U11529 (N_11529,N_11362,N_11499);
xor U11530 (N_11530,N_11333,N_11356);
nor U11531 (N_11531,N_11347,N_11379);
xnor U11532 (N_11532,N_11423,N_11341);
and U11533 (N_11533,N_11314,N_11338);
or U11534 (N_11534,N_11461,N_11259);
or U11535 (N_11535,N_11308,N_11282);
and U11536 (N_11536,N_11330,N_11354);
and U11537 (N_11537,N_11442,N_11253);
nor U11538 (N_11538,N_11350,N_11397);
and U11539 (N_11539,N_11398,N_11280);
nor U11540 (N_11540,N_11294,N_11315);
nand U11541 (N_11541,N_11439,N_11448);
nor U11542 (N_11542,N_11454,N_11368);
or U11543 (N_11543,N_11470,N_11444);
or U11544 (N_11544,N_11387,N_11498);
nor U11545 (N_11545,N_11265,N_11304);
or U11546 (N_11546,N_11447,N_11257);
nand U11547 (N_11547,N_11412,N_11465);
and U11548 (N_11548,N_11299,N_11331);
and U11549 (N_11549,N_11415,N_11455);
or U11550 (N_11550,N_11334,N_11285);
nor U11551 (N_11551,N_11399,N_11491);
or U11552 (N_11552,N_11360,N_11416);
nand U11553 (N_11553,N_11340,N_11424);
nor U11554 (N_11554,N_11435,N_11327);
xnor U11555 (N_11555,N_11369,N_11263);
and U11556 (N_11556,N_11462,N_11283);
nor U11557 (N_11557,N_11456,N_11276);
xor U11558 (N_11558,N_11476,N_11293);
and U11559 (N_11559,N_11422,N_11342);
nand U11560 (N_11560,N_11251,N_11351);
nand U11561 (N_11561,N_11425,N_11266);
and U11562 (N_11562,N_11344,N_11393);
nor U11563 (N_11563,N_11436,N_11404);
xor U11564 (N_11564,N_11291,N_11380);
nor U11565 (N_11565,N_11474,N_11483);
nand U11566 (N_11566,N_11429,N_11459);
nor U11567 (N_11567,N_11286,N_11497);
xor U11568 (N_11568,N_11372,N_11421);
and U11569 (N_11569,N_11384,N_11431);
xor U11570 (N_11570,N_11414,N_11250);
xor U11571 (N_11571,N_11320,N_11480);
and U11572 (N_11572,N_11484,N_11298);
xor U11573 (N_11573,N_11348,N_11295);
nor U11574 (N_11574,N_11281,N_11261);
nor U11575 (N_11575,N_11426,N_11254);
xnor U11576 (N_11576,N_11345,N_11411);
and U11577 (N_11577,N_11262,N_11252);
and U11578 (N_11578,N_11329,N_11337);
nor U11579 (N_11579,N_11289,N_11413);
nand U11580 (N_11580,N_11471,N_11272);
nor U11581 (N_11581,N_11452,N_11408);
nor U11582 (N_11582,N_11453,N_11326);
and U11583 (N_11583,N_11418,N_11378);
and U11584 (N_11584,N_11319,N_11284);
nor U11585 (N_11585,N_11395,N_11269);
nand U11586 (N_11586,N_11336,N_11306);
nor U11587 (N_11587,N_11325,N_11437);
nor U11588 (N_11588,N_11328,N_11358);
or U11589 (N_11589,N_11375,N_11279);
nand U11590 (N_11590,N_11302,N_11381);
and U11591 (N_11591,N_11475,N_11391);
xor U11592 (N_11592,N_11361,N_11376);
nor U11593 (N_11593,N_11463,N_11343);
and U11594 (N_11594,N_11366,N_11353);
nor U11595 (N_11595,N_11473,N_11479);
xnor U11596 (N_11596,N_11460,N_11450);
or U11597 (N_11597,N_11310,N_11312);
nor U11598 (N_11598,N_11466,N_11496);
nor U11599 (N_11599,N_11255,N_11371);
and U11600 (N_11600,N_11349,N_11446);
nor U11601 (N_11601,N_11482,N_11469);
nand U11602 (N_11602,N_11433,N_11440);
nor U11603 (N_11603,N_11400,N_11407);
and U11604 (N_11604,N_11392,N_11464);
xor U11605 (N_11605,N_11364,N_11490);
nor U11606 (N_11606,N_11394,N_11367);
xor U11607 (N_11607,N_11386,N_11301);
nor U11608 (N_11608,N_11290,N_11258);
nand U11609 (N_11609,N_11271,N_11273);
or U11610 (N_11610,N_11486,N_11303);
xnor U11611 (N_11611,N_11316,N_11323);
and U11612 (N_11612,N_11355,N_11318);
nor U11613 (N_11613,N_11417,N_11472);
nor U11614 (N_11614,N_11270,N_11434);
or U11615 (N_11615,N_11401,N_11489);
or U11616 (N_11616,N_11346,N_11457);
or U11617 (N_11617,N_11373,N_11317);
or U11618 (N_11618,N_11260,N_11478);
or U11619 (N_11619,N_11322,N_11410);
nand U11620 (N_11620,N_11267,N_11451);
xnor U11621 (N_11621,N_11268,N_11495);
and U11622 (N_11622,N_11477,N_11292);
nor U11623 (N_11623,N_11420,N_11300);
nand U11624 (N_11624,N_11274,N_11277);
xnor U11625 (N_11625,N_11479,N_11454);
or U11626 (N_11626,N_11384,N_11414);
or U11627 (N_11627,N_11488,N_11436);
xnor U11628 (N_11628,N_11413,N_11306);
nand U11629 (N_11629,N_11401,N_11405);
and U11630 (N_11630,N_11326,N_11296);
or U11631 (N_11631,N_11368,N_11476);
nand U11632 (N_11632,N_11319,N_11289);
nor U11633 (N_11633,N_11256,N_11453);
nor U11634 (N_11634,N_11318,N_11266);
and U11635 (N_11635,N_11311,N_11398);
and U11636 (N_11636,N_11275,N_11375);
nand U11637 (N_11637,N_11468,N_11355);
nor U11638 (N_11638,N_11393,N_11273);
or U11639 (N_11639,N_11330,N_11289);
nand U11640 (N_11640,N_11440,N_11347);
nor U11641 (N_11641,N_11421,N_11298);
nor U11642 (N_11642,N_11465,N_11485);
nand U11643 (N_11643,N_11439,N_11289);
xnor U11644 (N_11644,N_11294,N_11448);
nor U11645 (N_11645,N_11498,N_11334);
xnor U11646 (N_11646,N_11391,N_11398);
or U11647 (N_11647,N_11320,N_11325);
nor U11648 (N_11648,N_11466,N_11283);
nand U11649 (N_11649,N_11436,N_11277);
or U11650 (N_11650,N_11439,N_11322);
nand U11651 (N_11651,N_11433,N_11257);
xnor U11652 (N_11652,N_11486,N_11270);
nand U11653 (N_11653,N_11396,N_11457);
nor U11654 (N_11654,N_11254,N_11292);
nand U11655 (N_11655,N_11433,N_11313);
or U11656 (N_11656,N_11494,N_11491);
and U11657 (N_11657,N_11383,N_11386);
or U11658 (N_11658,N_11372,N_11344);
nand U11659 (N_11659,N_11383,N_11332);
or U11660 (N_11660,N_11408,N_11335);
nand U11661 (N_11661,N_11390,N_11302);
nor U11662 (N_11662,N_11271,N_11460);
xor U11663 (N_11663,N_11377,N_11381);
and U11664 (N_11664,N_11372,N_11277);
and U11665 (N_11665,N_11344,N_11440);
and U11666 (N_11666,N_11292,N_11490);
xnor U11667 (N_11667,N_11336,N_11409);
xor U11668 (N_11668,N_11393,N_11386);
nand U11669 (N_11669,N_11409,N_11341);
xnor U11670 (N_11670,N_11294,N_11431);
xor U11671 (N_11671,N_11286,N_11432);
xnor U11672 (N_11672,N_11467,N_11377);
nand U11673 (N_11673,N_11468,N_11484);
nor U11674 (N_11674,N_11462,N_11363);
or U11675 (N_11675,N_11432,N_11329);
xor U11676 (N_11676,N_11404,N_11442);
nand U11677 (N_11677,N_11305,N_11437);
or U11678 (N_11678,N_11499,N_11450);
nand U11679 (N_11679,N_11468,N_11259);
and U11680 (N_11680,N_11336,N_11438);
nor U11681 (N_11681,N_11286,N_11325);
nor U11682 (N_11682,N_11354,N_11407);
nor U11683 (N_11683,N_11251,N_11411);
and U11684 (N_11684,N_11486,N_11370);
xnor U11685 (N_11685,N_11478,N_11361);
nand U11686 (N_11686,N_11463,N_11402);
xor U11687 (N_11687,N_11484,N_11402);
nand U11688 (N_11688,N_11481,N_11413);
nor U11689 (N_11689,N_11299,N_11411);
or U11690 (N_11690,N_11288,N_11375);
or U11691 (N_11691,N_11345,N_11346);
nand U11692 (N_11692,N_11363,N_11420);
nand U11693 (N_11693,N_11260,N_11376);
nand U11694 (N_11694,N_11484,N_11351);
nor U11695 (N_11695,N_11366,N_11316);
nor U11696 (N_11696,N_11356,N_11447);
nand U11697 (N_11697,N_11378,N_11410);
nor U11698 (N_11698,N_11365,N_11295);
or U11699 (N_11699,N_11366,N_11481);
nor U11700 (N_11700,N_11493,N_11291);
and U11701 (N_11701,N_11332,N_11330);
xor U11702 (N_11702,N_11494,N_11467);
nor U11703 (N_11703,N_11323,N_11412);
and U11704 (N_11704,N_11386,N_11419);
nand U11705 (N_11705,N_11448,N_11359);
or U11706 (N_11706,N_11350,N_11457);
nor U11707 (N_11707,N_11253,N_11399);
nand U11708 (N_11708,N_11291,N_11460);
and U11709 (N_11709,N_11257,N_11486);
and U11710 (N_11710,N_11366,N_11359);
and U11711 (N_11711,N_11408,N_11488);
or U11712 (N_11712,N_11480,N_11354);
nor U11713 (N_11713,N_11443,N_11331);
and U11714 (N_11714,N_11271,N_11367);
and U11715 (N_11715,N_11440,N_11427);
nor U11716 (N_11716,N_11472,N_11366);
nand U11717 (N_11717,N_11350,N_11314);
or U11718 (N_11718,N_11433,N_11482);
xor U11719 (N_11719,N_11466,N_11384);
nor U11720 (N_11720,N_11385,N_11292);
nor U11721 (N_11721,N_11356,N_11272);
nor U11722 (N_11722,N_11433,N_11403);
nor U11723 (N_11723,N_11270,N_11411);
xnor U11724 (N_11724,N_11490,N_11429);
nand U11725 (N_11725,N_11473,N_11445);
xor U11726 (N_11726,N_11472,N_11396);
or U11727 (N_11727,N_11301,N_11381);
or U11728 (N_11728,N_11422,N_11489);
nor U11729 (N_11729,N_11335,N_11321);
and U11730 (N_11730,N_11322,N_11424);
nand U11731 (N_11731,N_11494,N_11316);
xor U11732 (N_11732,N_11294,N_11469);
or U11733 (N_11733,N_11459,N_11437);
or U11734 (N_11734,N_11407,N_11280);
and U11735 (N_11735,N_11256,N_11395);
or U11736 (N_11736,N_11331,N_11342);
xor U11737 (N_11737,N_11445,N_11477);
and U11738 (N_11738,N_11422,N_11445);
nand U11739 (N_11739,N_11455,N_11370);
nand U11740 (N_11740,N_11286,N_11361);
nand U11741 (N_11741,N_11326,N_11310);
nor U11742 (N_11742,N_11346,N_11263);
and U11743 (N_11743,N_11306,N_11346);
xor U11744 (N_11744,N_11305,N_11331);
and U11745 (N_11745,N_11265,N_11298);
nor U11746 (N_11746,N_11488,N_11395);
xor U11747 (N_11747,N_11408,N_11456);
and U11748 (N_11748,N_11349,N_11449);
or U11749 (N_11749,N_11493,N_11261);
and U11750 (N_11750,N_11578,N_11712);
xor U11751 (N_11751,N_11739,N_11599);
nor U11752 (N_11752,N_11609,N_11644);
nor U11753 (N_11753,N_11746,N_11553);
xnor U11754 (N_11754,N_11711,N_11501);
nor U11755 (N_11755,N_11659,N_11592);
nand U11756 (N_11756,N_11694,N_11520);
nor U11757 (N_11757,N_11568,N_11745);
nor U11758 (N_11758,N_11575,N_11563);
or U11759 (N_11759,N_11702,N_11582);
or U11760 (N_11760,N_11721,N_11729);
xor U11761 (N_11761,N_11654,N_11671);
and U11762 (N_11762,N_11580,N_11613);
xnor U11763 (N_11763,N_11640,N_11571);
and U11764 (N_11764,N_11519,N_11699);
or U11765 (N_11765,N_11536,N_11572);
and U11766 (N_11766,N_11635,N_11730);
and U11767 (N_11767,N_11638,N_11576);
nor U11768 (N_11768,N_11742,N_11608);
xnor U11769 (N_11769,N_11627,N_11577);
nor U11770 (N_11770,N_11561,N_11688);
or U11771 (N_11771,N_11593,N_11538);
nand U11772 (N_11772,N_11545,N_11612);
and U11773 (N_11773,N_11529,N_11723);
xnor U11774 (N_11774,N_11722,N_11598);
nor U11775 (N_11775,N_11686,N_11676);
nor U11776 (N_11776,N_11685,N_11714);
and U11777 (N_11777,N_11629,N_11567);
and U11778 (N_11778,N_11617,N_11698);
nor U11779 (N_11779,N_11513,N_11621);
or U11780 (N_11780,N_11653,N_11590);
xnor U11781 (N_11781,N_11648,N_11566);
nand U11782 (N_11782,N_11707,N_11517);
or U11783 (N_11783,N_11533,N_11715);
and U11784 (N_11784,N_11646,N_11634);
nand U11785 (N_11785,N_11740,N_11717);
and U11786 (N_11786,N_11547,N_11650);
nor U11787 (N_11787,N_11594,N_11525);
xor U11788 (N_11788,N_11727,N_11583);
xnor U11789 (N_11789,N_11666,N_11546);
nand U11790 (N_11790,N_11663,N_11539);
or U11791 (N_11791,N_11570,N_11726);
and U11792 (N_11792,N_11509,N_11541);
xnor U11793 (N_11793,N_11674,N_11584);
and U11794 (N_11794,N_11589,N_11744);
xnor U11795 (N_11795,N_11511,N_11741);
nor U11796 (N_11796,N_11530,N_11642);
nor U11797 (N_11797,N_11690,N_11696);
and U11798 (N_11798,N_11679,N_11728);
nor U11799 (N_11799,N_11595,N_11619);
and U11800 (N_11800,N_11656,N_11504);
or U11801 (N_11801,N_11558,N_11720);
and U11802 (N_11802,N_11655,N_11573);
nand U11803 (N_11803,N_11625,N_11710);
nand U11804 (N_11804,N_11603,N_11596);
nor U11805 (N_11805,N_11556,N_11719);
nand U11806 (N_11806,N_11660,N_11651);
nor U11807 (N_11807,N_11557,N_11652);
nor U11808 (N_11808,N_11586,N_11531);
xnor U11809 (N_11809,N_11725,N_11591);
nand U11810 (N_11810,N_11647,N_11673);
nand U11811 (N_11811,N_11581,N_11522);
xor U11812 (N_11812,N_11675,N_11678);
nor U11813 (N_11813,N_11551,N_11624);
nand U11814 (N_11814,N_11540,N_11526);
or U11815 (N_11815,N_11701,N_11623);
nand U11816 (N_11816,N_11709,N_11693);
and U11817 (N_11817,N_11555,N_11502);
nand U11818 (N_11818,N_11610,N_11649);
xor U11819 (N_11819,N_11636,N_11512);
nand U11820 (N_11820,N_11639,N_11569);
nor U11821 (N_11821,N_11677,N_11508);
xor U11822 (N_11822,N_11543,N_11631);
nand U11823 (N_11823,N_11606,N_11705);
or U11824 (N_11824,N_11661,N_11667);
nor U11825 (N_11825,N_11645,N_11510);
or U11826 (N_11826,N_11743,N_11534);
or U11827 (N_11827,N_11713,N_11620);
or U11828 (N_11828,N_11664,N_11697);
xor U11829 (N_11829,N_11507,N_11514);
xnor U11830 (N_11830,N_11550,N_11670);
nand U11831 (N_11831,N_11542,N_11518);
nand U11832 (N_11832,N_11658,N_11641);
or U11833 (N_11833,N_11565,N_11515);
nor U11834 (N_11834,N_11616,N_11588);
and U11835 (N_11835,N_11523,N_11749);
nand U11836 (N_11836,N_11718,N_11600);
xnor U11837 (N_11837,N_11632,N_11548);
nand U11838 (N_11838,N_11552,N_11528);
nand U11839 (N_11839,N_11505,N_11732);
nor U11840 (N_11840,N_11503,N_11735);
or U11841 (N_11841,N_11604,N_11682);
or U11842 (N_11842,N_11681,N_11602);
xnor U11843 (N_11843,N_11537,N_11691);
nand U11844 (N_11844,N_11687,N_11549);
and U11845 (N_11845,N_11700,N_11704);
nand U11846 (N_11846,N_11692,N_11657);
or U11847 (N_11847,N_11668,N_11665);
nor U11848 (N_11848,N_11662,N_11500);
nor U11849 (N_11849,N_11607,N_11669);
xnor U11850 (N_11850,N_11532,N_11747);
or U11851 (N_11851,N_11579,N_11618);
nand U11852 (N_11852,N_11703,N_11626);
xnor U11853 (N_11853,N_11587,N_11535);
and U11854 (N_11854,N_11643,N_11684);
nand U11855 (N_11855,N_11516,N_11559);
nor U11856 (N_11856,N_11562,N_11630);
nand U11857 (N_11857,N_11736,N_11521);
and U11858 (N_11858,N_11637,N_11628);
nand U11859 (N_11859,N_11737,N_11544);
xor U11860 (N_11860,N_11689,N_11527);
or U11861 (N_11861,N_11597,N_11601);
and U11862 (N_11862,N_11706,N_11585);
nor U11863 (N_11863,N_11734,N_11574);
and U11864 (N_11864,N_11683,N_11731);
xnor U11865 (N_11865,N_11680,N_11564);
or U11866 (N_11866,N_11605,N_11560);
nor U11867 (N_11867,N_11614,N_11695);
or U11868 (N_11868,N_11615,N_11506);
nand U11869 (N_11869,N_11524,N_11716);
nand U11870 (N_11870,N_11611,N_11724);
nor U11871 (N_11871,N_11672,N_11633);
nand U11872 (N_11872,N_11733,N_11554);
xor U11873 (N_11873,N_11738,N_11708);
xor U11874 (N_11874,N_11748,N_11622);
nor U11875 (N_11875,N_11610,N_11674);
xor U11876 (N_11876,N_11542,N_11717);
nor U11877 (N_11877,N_11576,N_11555);
nand U11878 (N_11878,N_11718,N_11684);
nand U11879 (N_11879,N_11678,N_11520);
xnor U11880 (N_11880,N_11607,N_11748);
xnor U11881 (N_11881,N_11567,N_11645);
or U11882 (N_11882,N_11523,N_11659);
nand U11883 (N_11883,N_11530,N_11688);
and U11884 (N_11884,N_11525,N_11674);
and U11885 (N_11885,N_11552,N_11520);
xor U11886 (N_11886,N_11626,N_11542);
or U11887 (N_11887,N_11653,N_11610);
xnor U11888 (N_11888,N_11551,N_11699);
nand U11889 (N_11889,N_11611,N_11557);
and U11890 (N_11890,N_11685,N_11502);
and U11891 (N_11891,N_11584,N_11642);
or U11892 (N_11892,N_11600,N_11518);
nand U11893 (N_11893,N_11553,N_11532);
nand U11894 (N_11894,N_11651,N_11525);
nor U11895 (N_11895,N_11541,N_11703);
nor U11896 (N_11896,N_11547,N_11605);
xor U11897 (N_11897,N_11714,N_11617);
or U11898 (N_11898,N_11539,N_11634);
or U11899 (N_11899,N_11507,N_11568);
nand U11900 (N_11900,N_11612,N_11503);
and U11901 (N_11901,N_11513,N_11692);
nand U11902 (N_11902,N_11605,N_11503);
nor U11903 (N_11903,N_11739,N_11737);
and U11904 (N_11904,N_11672,N_11742);
nor U11905 (N_11905,N_11540,N_11704);
nand U11906 (N_11906,N_11716,N_11584);
nor U11907 (N_11907,N_11530,N_11514);
nand U11908 (N_11908,N_11701,N_11678);
or U11909 (N_11909,N_11614,N_11696);
and U11910 (N_11910,N_11539,N_11679);
and U11911 (N_11911,N_11624,N_11601);
nand U11912 (N_11912,N_11712,N_11656);
xnor U11913 (N_11913,N_11513,N_11732);
and U11914 (N_11914,N_11677,N_11738);
xnor U11915 (N_11915,N_11572,N_11689);
nor U11916 (N_11916,N_11588,N_11551);
xor U11917 (N_11917,N_11618,N_11646);
or U11918 (N_11918,N_11587,N_11673);
nor U11919 (N_11919,N_11683,N_11601);
and U11920 (N_11920,N_11503,N_11710);
or U11921 (N_11921,N_11749,N_11525);
or U11922 (N_11922,N_11551,N_11512);
or U11923 (N_11923,N_11624,N_11693);
nor U11924 (N_11924,N_11693,N_11655);
nor U11925 (N_11925,N_11691,N_11540);
nor U11926 (N_11926,N_11555,N_11514);
nand U11927 (N_11927,N_11633,N_11502);
nand U11928 (N_11928,N_11604,N_11542);
xnor U11929 (N_11929,N_11666,N_11663);
or U11930 (N_11930,N_11732,N_11644);
nand U11931 (N_11931,N_11572,N_11678);
nor U11932 (N_11932,N_11597,N_11515);
nand U11933 (N_11933,N_11566,N_11603);
xnor U11934 (N_11934,N_11510,N_11614);
and U11935 (N_11935,N_11619,N_11701);
xor U11936 (N_11936,N_11617,N_11621);
nor U11937 (N_11937,N_11643,N_11646);
or U11938 (N_11938,N_11621,N_11733);
and U11939 (N_11939,N_11612,N_11709);
and U11940 (N_11940,N_11749,N_11673);
and U11941 (N_11941,N_11508,N_11697);
and U11942 (N_11942,N_11659,N_11558);
nand U11943 (N_11943,N_11695,N_11512);
xor U11944 (N_11944,N_11616,N_11738);
or U11945 (N_11945,N_11682,N_11677);
xor U11946 (N_11946,N_11723,N_11718);
nand U11947 (N_11947,N_11581,N_11740);
or U11948 (N_11948,N_11522,N_11536);
nand U11949 (N_11949,N_11602,N_11620);
nor U11950 (N_11950,N_11532,N_11588);
and U11951 (N_11951,N_11613,N_11642);
xor U11952 (N_11952,N_11515,N_11649);
or U11953 (N_11953,N_11690,N_11551);
and U11954 (N_11954,N_11704,N_11615);
nand U11955 (N_11955,N_11689,N_11649);
and U11956 (N_11956,N_11643,N_11740);
nand U11957 (N_11957,N_11554,N_11558);
or U11958 (N_11958,N_11637,N_11699);
and U11959 (N_11959,N_11681,N_11679);
and U11960 (N_11960,N_11648,N_11558);
and U11961 (N_11961,N_11640,N_11655);
nor U11962 (N_11962,N_11601,N_11661);
and U11963 (N_11963,N_11706,N_11742);
or U11964 (N_11964,N_11542,N_11685);
xnor U11965 (N_11965,N_11502,N_11643);
or U11966 (N_11966,N_11656,N_11587);
xnor U11967 (N_11967,N_11601,N_11637);
or U11968 (N_11968,N_11529,N_11558);
or U11969 (N_11969,N_11558,N_11737);
or U11970 (N_11970,N_11578,N_11526);
or U11971 (N_11971,N_11613,N_11709);
and U11972 (N_11972,N_11623,N_11575);
nor U11973 (N_11973,N_11731,N_11735);
and U11974 (N_11974,N_11509,N_11574);
or U11975 (N_11975,N_11621,N_11611);
or U11976 (N_11976,N_11619,N_11578);
nor U11977 (N_11977,N_11633,N_11719);
xor U11978 (N_11978,N_11574,N_11693);
nand U11979 (N_11979,N_11598,N_11706);
and U11980 (N_11980,N_11607,N_11650);
nand U11981 (N_11981,N_11552,N_11678);
and U11982 (N_11982,N_11733,N_11631);
or U11983 (N_11983,N_11658,N_11740);
or U11984 (N_11984,N_11663,N_11728);
nand U11985 (N_11985,N_11636,N_11524);
or U11986 (N_11986,N_11527,N_11528);
or U11987 (N_11987,N_11597,N_11613);
xnor U11988 (N_11988,N_11559,N_11615);
and U11989 (N_11989,N_11724,N_11743);
nand U11990 (N_11990,N_11524,N_11712);
xnor U11991 (N_11991,N_11676,N_11590);
nor U11992 (N_11992,N_11689,N_11710);
or U11993 (N_11993,N_11619,N_11625);
and U11994 (N_11994,N_11743,N_11592);
and U11995 (N_11995,N_11502,N_11520);
or U11996 (N_11996,N_11540,N_11687);
xor U11997 (N_11997,N_11524,N_11502);
nor U11998 (N_11998,N_11674,N_11539);
and U11999 (N_11999,N_11555,N_11575);
and U12000 (N_12000,N_11944,N_11801);
nor U12001 (N_12001,N_11909,N_11892);
xor U12002 (N_12002,N_11951,N_11906);
xnor U12003 (N_12003,N_11868,N_11967);
or U12004 (N_12004,N_11936,N_11761);
nor U12005 (N_12005,N_11949,N_11904);
nand U12006 (N_12006,N_11770,N_11966);
xnor U12007 (N_12007,N_11871,N_11958);
or U12008 (N_12008,N_11901,N_11941);
or U12009 (N_12009,N_11907,N_11838);
nor U12010 (N_12010,N_11803,N_11779);
xnor U12011 (N_12011,N_11980,N_11775);
or U12012 (N_12012,N_11865,N_11862);
xnor U12013 (N_12013,N_11792,N_11992);
nor U12014 (N_12014,N_11880,N_11939);
nor U12015 (N_12015,N_11758,N_11886);
xor U12016 (N_12016,N_11935,N_11953);
nor U12017 (N_12017,N_11916,N_11827);
nand U12018 (N_12018,N_11981,N_11898);
nor U12019 (N_12019,N_11993,N_11872);
nand U12020 (N_12020,N_11855,N_11920);
or U12021 (N_12021,N_11791,N_11945);
or U12022 (N_12022,N_11832,N_11963);
nand U12023 (N_12023,N_11969,N_11989);
or U12024 (N_12024,N_11813,N_11790);
and U12025 (N_12025,N_11850,N_11889);
nor U12026 (N_12026,N_11995,N_11783);
nor U12027 (N_12027,N_11768,N_11873);
nor U12028 (N_12028,N_11990,N_11903);
nor U12029 (N_12029,N_11856,N_11879);
nor U12030 (N_12030,N_11883,N_11787);
xnor U12031 (N_12031,N_11986,N_11960);
nand U12032 (N_12032,N_11962,N_11784);
and U12033 (N_12033,N_11917,N_11776);
xor U12034 (N_12034,N_11789,N_11788);
and U12035 (N_12035,N_11817,N_11846);
xnor U12036 (N_12036,N_11965,N_11751);
xor U12037 (N_12037,N_11928,N_11946);
and U12038 (N_12038,N_11837,N_11964);
nor U12039 (N_12039,N_11805,N_11811);
and U12040 (N_12040,N_11825,N_11853);
and U12041 (N_12041,N_11913,N_11753);
or U12042 (N_12042,N_11925,N_11972);
and U12043 (N_12043,N_11999,N_11952);
nor U12044 (N_12044,N_11942,N_11839);
or U12045 (N_12045,N_11826,N_11998);
nand U12046 (N_12046,N_11819,N_11894);
and U12047 (N_12047,N_11971,N_11822);
nor U12048 (N_12048,N_11836,N_11754);
and U12049 (N_12049,N_11984,N_11875);
xnor U12050 (N_12050,N_11785,N_11937);
and U12051 (N_12051,N_11867,N_11897);
or U12052 (N_12052,N_11845,N_11843);
or U12053 (N_12053,N_11834,N_11772);
nand U12054 (N_12054,N_11908,N_11977);
nand U12055 (N_12055,N_11996,N_11888);
or U12056 (N_12056,N_11982,N_11912);
and U12057 (N_12057,N_11929,N_11757);
nand U12058 (N_12058,N_11816,N_11899);
xor U12059 (N_12059,N_11800,N_11764);
or U12060 (N_12060,N_11881,N_11970);
nor U12061 (N_12061,N_11759,N_11896);
xnor U12062 (N_12062,N_11882,N_11885);
nand U12063 (N_12063,N_11915,N_11807);
xor U12064 (N_12064,N_11814,N_11878);
xnor U12065 (N_12065,N_11798,N_11922);
nand U12066 (N_12066,N_11988,N_11927);
xnor U12067 (N_12067,N_11831,N_11760);
and U12068 (N_12068,N_11854,N_11847);
nand U12069 (N_12069,N_11848,N_11808);
xor U12070 (N_12070,N_11812,N_11884);
xor U12071 (N_12071,N_11893,N_11777);
nand U12072 (N_12072,N_11820,N_11786);
and U12073 (N_12073,N_11976,N_11766);
or U12074 (N_12074,N_11959,N_11858);
or U12075 (N_12075,N_11806,N_11752);
or U12076 (N_12076,N_11891,N_11943);
nand U12077 (N_12077,N_11961,N_11940);
nand U12078 (N_12078,N_11973,N_11950);
or U12079 (N_12079,N_11797,N_11974);
and U12080 (N_12080,N_11833,N_11821);
and U12081 (N_12081,N_11934,N_11948);
xor U12082 (N_12082,N_11890,N_11818);
nand U12083 (N_12083,N_11985,N_11956);
or U12084 (N_12084,N_11921,N_11756);
and U12085 (N_12085,N_11923,N_11844);
nor U12086 (N_12086,N_11991,N_11762);
xor U12087 (N_12087,N_11769,N_11810);
nand U12088 (N_12088,N_11851,N_11918);
nand U12089 (N_12089,N_11931,N_11824);
nor U12090 (N_12090,N_11835,N_11849);
xor U12091 (N_12091,N_11947,N_11975);
nand U12092 (N_12092,N_11978,N_11809);
xor U12093 (N_12093,N_11864,N_11910);
nand U12094 (N_12094,N_11804,N_11828);
xor U12095 (N_12095,N_11860,N_11887);
xnor U12096 (N_12096,N_11767,N_11840);
xor U12097 (N_12097,N_11765,N_11780);
and U12098 (N_12098,N_11895,N_11924);
and U12099 (N_12099,N_11938,N_11874);
or U12100 (N_12100,N_11852,N_11930);
and U12101 (N_12101,N_11900,N_11983);
and U12102 (N_12102,N_11782,N_11750);
nor U12103 (N_12103,N_11954,N_11968);
or U12104 (N_12104,N_11876,N_11793);
xnor U12105 (N_12105,N_11933,N_11902);
nand U12106 (N_12106,N_11778,N_11861);
xnor U12107 (N_12107,N_11842,N_11979);
nand U12108 (N_12108,N_11869,N_11911);
nand U12109 (N_12109,N_11870,N_11919);
or U12110 (N_12110,N_11774,N_11794);
nand U12111 (N_12111,N_11781,N_11763);
nor U12112 (N_12112,N_11830,N_11829);
or U12113 (N_12113,N_11866,N_11857);
or U12114 (N_12114,N_11987,N_11877);
nand U12115 (N_12115,N_11957,N_11863);
xnor U12116 (N_12116,N_11955,N_11997);
xor U12117 (N_12117,N_11823,N_11755);
xor U12118 (N_12118,N_11932,N_11905);
or U12119 (N_12119,N_11771,N_11796);
nor U12120 (N_12120,N_11802,N_11841);
nor U12121 (N_12121,N_11926,N_11994);
xnor U12122 (N_12122,N_11815,N_11859);
nand U12123 (N_12123,N_11773,N_11914);
nor U12124 (N_12124,N_11795,N_11799);
and U12125 (N_12125,N_11852,N_11933);
and U12126 (N_12126,N_11876,N_11753);
and U12127 (N_12127,N_11971,N_11834);
xnor U12128 (N_12128,N_11881,N_11923);
and U12129 (N_12129,N_11841,N_11886);
nor U12130 (N_12130,N_11857,N_11931);
or U12131 (N_12131,N_11792,N_11774);
or U12132 (N_12132,N_11982,N_11816);
nor U12133 (N_12133,N_11754,N_11953);
or U12134 (N_12134,N_11913,N_11774);
or U12135 (N_12135,N_11806,N_11961);
and U12136 (N_12136,N_11858,N_11911);
and U12137 (N_12137,N_11816,N_11927);
or U12138 (N_12138,N_11828,N_11897);
xor U12139 (N_12139,N_11914,N_11903);
or U12140 (N_12140,N_11972,N_11990);
or U12141 (N_12141,N_11756,N_11794);
or U12142 (N_12142,N_11797,N_11862);
and U12143 (N_12143,N_11953,N_11776);
nand U12144 (N_12144,N_11768,N_11767);
nor U12145 (N_12145,N_11848,N_11887);
and U12146 (N_12146,N_11994,N_11867);
or U12147 (N_12147,N_11774,N_11963);
xor U12148 (N_12148,N_11779,N_11913);
nand U12149 (N_12149,N_11916,N_11880);
nor U12150 (N_12150,N_11896,N_11958);
xor U12151 (N_12151,N_11791,N_11880);
nand U12152 (N_12152,N_11858,N_11807);
or U12153 (N_12153,N_11833,N_11807);
nor U12154 (N_12154,N_11886,N_11959);
and U12155 (N_12155,N_11972,N_11962);
and U12156 (N_12156,N_11881,N_11806);
or U12157 (N_12157,N_11773,N_11848);
nand U12158 (N_12158,N_11824,N_11797);
nand U12159 (N_12159,N_11824,N_11990);
and U12160 (N_12160,N_11841,N_11894);
nor U12161 (N_12161,N_11848,N_11854);
nor U12162 (N_12162,N_11834,N_11846);
nand U12163 (N_12163,N_11864,N_11792);
or U12164 (N_12164,N_11902,N_11791);
or U12165 (N_12165,N_11798,N_11840);
xnor U12166 (N_12166,N_11773,N_11894);
xor U12167 (N_12167,N_11839,N_11903);
or U12168 (N_12168,N_11994,N_11876);
or U12169 (N_12169,N_11829,N_11819);
nand U12170 (N_12170,N_11809,N_11880);
nand U12171 (N_12171,N_11776,N_11847);
xor U12172 (N_12172,N_11916,N_11970);
nand U12173 (N_12173,N_11849,N_11790);
nor U12174 (N_12174,N_11820,N_11757);
and U12175 (N_12175,N_11975,N_11792);
and U12176 (N_12176,N_11841,N_11752);
xnor U12177 (N_12177,N_11860,N_11946);
or U12178 (N_12178,N_11980,N_11816);
nand U12179 (N_12179,N_11891,N_11907);
and U12180 (N_12180,N_11823,N_11814);
nor U12181 (N_12181,N_11934,N_11886);
or U12182 (N_12182,N_11884,N_11910);
nor U12183 (N_12183,N_11854,N_11793);
nand U12184 (N_12184,N_11958,N_11977);
nor U12185 (N_12185,N_11968,N_11767);
xor U12186 (N_12186,N_11977,N_11998);
or U12187 (N_12187,N_11882,N_11987);
nor U12188 (N_12188,N_11766,N_11998);
and U12189 (N_12189,N_11848,N_11778);
and U12190 (N_12190,N_11835,N_11785);
or U12191 (N_12191,N_11839,N_11961);
nor U12192 (N_12192,N_11981,N_11920);
xor U12193 (N_12193,N_11918,N_11983);
xor U12194 (N_12194,N_11937,N_11776);
nor U12195 (N_12195,N_11847,N_11996);
xor U12196 (N_12196,N_11934,N_11968);
nor U12197 (N_12197,N_11852,N_11963);
nand U12198 (N_12198,N_11759,N_11910);
nor U12199 (N_12199,N_11880,N_11979);
nand U12200 (N_12200,N_11845,N_11817);
xnor U12201 (N_12201,N_11785,N_11820);
and U12202 (N_12202,N_11886,N_11895);
nor U12203 (N_12203,N_11879,N_11987);
nand U12204 (N_12204,N_11969,N_11827);
or U12205 (N_12205,N_11771,N_11996);
xnor U12206 (N_12206,N_11799,N_11874);
nor U12207 (N_12207,N_11970,N_11844);
and U12208 (N_12208,N_11900,N_11762);
or U12209 (N_12209,N_11968,N_11992);
nand U12210 (N_12210,N_11980,N_11812);
or U12211 (N_12211,N_11909,N_11777);
nor U12212 (N_12212,N_11804,N_11934);
nor U12213 (N_12213,N_11884,N_11768);
nand U12214 (N_12214,N_11761,N_11910);
and U12215 (N_12215,N_11980,N_11871);
xnor U12216 (N_12216,N_11753,N_11993);
xor U12217 (N_12217,N_11981,N_11954);
and U12218 (N_12218,N_11841,N_11786);
or U12219 (N_12219,N_11866,N_11884);
or U12220 (N_12220,N_11848,N_11903);
or U12221 (N_12221,N_11899,N_11876);
nor U12222 (N_12222,N_11874,N_11807);
nor U12223 (N_12223,N_11872,N_11768);
or U12224 (N_12224,N_11981,N_11991);
or U12225 (N_12225,N_11865,N_11841);
xor U12226 (N_12226,N_11915,N_11973);
or U12227 (N_12227,N_11752,N_11793);
xor U12228 (N_12228,N_11931,N_11974);
xnor U12229 (N_12229,N_11994,N_11905);
xor U12230 (N_12230,N_11878,N_11976);
nand U12231 (N_12231,N_11921,N_11750);
nor U12232 (N_12232,N_11928,N_11912);
nor U12233 (N_12233,N_11852,N_11799);
and U12234 (N_12234,N_11779,N_11754);
xor U12235 (N_12235,N_11840,N_11856);
xor U12236 (N_12236,N_11911,N_11791);
nor U12237 (N_12237,N_11978,N_11920);
nor U12238 (N_12238,N_11901,N_11816);
xnor U12239 (N_12239,N_11895,N_11846);
nand U12240 (N_12240,N_11915,N_11947);
or U12241 (N_12241,N_11838,N_11827);
nand U12242 (N_12242,N_11868,N_11790);
nand U12243 (N_12243,N_11809,N_11877);
or U12244 (N_12244,N_11882,N_11869);
or U12245 (N_12245,N_11863,N_11934);
and U12246 (N_12246,N_11763,N_11842);
nand U12247 (N_12247,N_11971,N_11828);
nand U12248 (N_12248,N_11873,N_11918);
and U12249 (N_12249,N_11890,N_11986);
and U12250 (N_12250,N_12003,N_12204);
xnor U12251 (N_12251,N_12143,N_12159);
nor U12252 (N_12252,N_12062,N_12208);
xor U12253 (N_12253,N_12076,N_12164);
xor U12254 (N_12254,N_12100,N_12188);
or U12255 (N_12255,N_12184,N_12185);
or U12256 (N_12256,N_12229,N_12104);
and U12257 (N_12257,N_12019,N_12101);
nor U12258 (N_12258,N_12212,N_12218);
nand U12259 (N_12259,N_12079,N_12065);
nand U12260 (N_12260,N_12162,N_12112);
and U12261 (N_12261,N_12141,N_12091);
nand U12262 (N_12262,N_12055,N_12040);
xnor U12263 (N_12263,N_12048,N_12182);
or U12264 (N_12264,N_12024,N_12210);
xor U12265 (N_12265,N_12113,N_12151);
xor U12266 (N_12266,N_12220,N_12221);
nand U12267 (N_12267,N_12150,N_12012);
and U12268 (N_12268,N_12059,N_12034);
or U12269 (N_12269,N_12053,N_12016);
or U12270 (N_12270,N_12197,N_12237);
and U12271 (N_12271,N_12072,N_12032);
nand U12272 (N_12272,N_12145,N_12238);
or U12273 (N_12273,N_12168,N_12010);
and U12274 (N_12274,N_12224,N_12060);
or U12275 (N_12275,N_12014,N_12147);
nand U12276 (N_12276,N_12183,N_12144);
and U12277 (N_12277,N_12152,N_12045);
nor U12278 (N_12278,N_12105,N_12126);
nand U12279 (N_12279,N_12242,N_12037);
nor U12280 (N_12280,N_12022,N_12240);
xnor U12281 (N_12281,N_12249,N_12115);
nor U12282 (N_12282,N_12050,N_12125);
and U12283 (N_12283,N_12200,N_12085);
and U12284 (N_12284,N_12138,N_12146);
and U12285 (N_12285,N_12083,N_12142);
xnor U12286 (N_12286,N_12128,N_12130);
or U12287 (N_12287,N_12047,N_12061);
nand U12288 (N_12288,N_12018,N_12167);
and U12289 (N_12289,N_12219,N_12133);
nand U12290 (N_12290,N_12154,N_12201);
xnor U12291 (N_12291,N_12023,N_12004);
or U12292 (N_12292,N_12231,N_12127);
and U12293 (N_12293,N_12013,N_12225);
xor U12294 (N_12294,N_12025,N_12129);
and U12295 (N_12295,N_12245,N_12118);
nor U12296 (N_12296,N_12235,N_12068);
xor U12297 (N_12297,N_12227,N_12234);
nor U12298 (N_12298,N_12171,N_12187);
and U12299 (N_12299,N_12029,N_12122);
nor U12300 (N_12300,N_12054,N_12078);
or U12301 (N_12301,N_12230,N_12136);
xor U12302 (N_12302,N_12244,N_12156);
nor U12303 (N_12303,N_12058,N_12033);
xor U12304 (N_12304,N_12158,N_12035);
nand U12305 (N_12305,N_12199,N_12228);
or U12306 (N_12306,N_12075,N_12096);
and U12307 (N_12307,N_12193,N_12009);
nor U12308 (N_12308,N_12117,N_12057);
nor U12309 (N_12309,N_12081,N_12216);
nand U12310 (N_12310,N_12198,N_12215);
nor U12311 (N_12311,N_12106,N_12140);
nand U12312 (N_12312,N_12211,N_12008);
or U12313 (N_12313,N_12203,N_12177);
and U12314 (N_12314,N_12002,N_12064);
nand U12315 (N_12315,N_12176,N_12090);
nor U12316 (N_12316,N_12137,N_12073);
nor U12317 (N_12317,N_12042,N_12170);
and U12318 (N_12318,N_12031,N_12087);
nand U12319 (N_12319,N_12036,N_12131);
nor U12320 (N_12320,N_12000,N_12155);
nor U12321 (N_12321,N_12098,N_12194);
nor U12322 (N_12322,N_12189,N_12132);
or U12323 (N_12323,N_12015,N_12056);
nand U12324 (N_12324,N_12069,N_12181);
nand U12325 (N_12325,N_12148,N_12063);
and U12326 (N_12326,N_12174,N_12080);
or U12327 (N_12327,N_12030,N_12214);
nand U12328 (N_12328,N_12052,N_12149);
xor U12329 (N_12329,N_12166,N_12202);
or U12330 (N_12330,N_12094,N_12093);
nor U12331 (N_12331,N_12173,N_12206);
or U12332 (N_12332,N_12049,N_12066);
xor U12333 (N_12333,N_12074,N_12120);
nand U12334 (N_12334,N_12169,N_12051);
xnor U12335 (N_12335,N_12165,N_12089);
nor U12336 (N_12336,N_12239,N_12071);
nor U12337 (N_12337,N_12119,N_12223);
nor U12338 (N_12338,N_12232,N_12135);
or U12339 (N_12339,N_12213,N_12038);
or U12340 (N_12340,N_12180,N_12092);
xor U12341 (N_12341,N_12196,N_12191);
or U12342 (N_12342,N_12028,N_12108);
or U12343 (N_12343,N_12099,N_12190);
or U12344 (N_12344,N_12007,N_12095);
or U12345 (N_12345,N_12192,N_12001);
and U12346 (N_12346,N_12124,N_12041);
and U12347 (N_12347,N_12121,N_12111);
or U12348 (N_12348,N_12044,N_12020);
nor U12349 (N_12349,N_12017,N_12070);
and U12350 (N_12350,N_12161,N_12114);
xor U12351 (N_12351,N_12233,N_12186);
nand U12352 (N_12352,N_12236,N_12043);
or U12353 (N_12353,N_12102,N_12103);
nor U12354 (N_12354,N_12139,N_12021);
nand U12355 (N_12355,N_12246,N_12226);
nand U12356 (N_12356,N_12153,N_12178);
xnor U12357 (N_12357,N_12179,N_12207);
nand U12358 (N_12358,N_12027,N_12172);
nor U12359 (N_12359,N_12082,N_12241);
nand U12360 (N_12360,N_12011,N_12134);
xor U12361 (N_12361,N_12067,N_12086);
nand U12362 (N_12362,N_12205,N_12077);
or U12363 (N_12363,N_12163,N_12175);
xnor U12364 (N_12364,N_12046,N_12006);
xnor U12365 (N_12365,N_12157,N_12217);
nand U12366 (N_12366,N_12243,N_12160);
nand U12367 (N_12367,N_12039,N_12123);
xor U12368 (N_12368,N_12084,N_12088);
nand U12369 (N_12369,N_12109,N_12222);
nor U12370 (N_12370,N_12097,N_12209);
xnor U12371 (N_12371,N_12026,N_12005);
xnor U12372 (N_12372,N_12107,N_12110);
nor U12373 (N_12373,N_12247,N_12195);
and U12374 (N_12374,N_12248,N_12116);
xor U12375 (N_12375,N_12226,N_12017);
and U12376 (N_12376,N_12095,N_12184);
nor U12377 (N_12377,N_12023,N_12090);
nor U12378 (N_12378,N_12133,N_12035);
nor U12379 (N_12379,N_12249,N_12096);
nand U12380 (N_12380,N_12008,N_12044);
or U12381 (N_12381,N_12226,N_12211);
or U12382 (N_12382,N_12207,N_12038);
nor U12383 (N_12383,N_12218,N_12003);
xor U12384 (N_12384,N_12175,N_12180);
nand U12385 (N_12385,N_12211,N_12224);
or U12386 (N_12386,N_12239,N_12160);
or U12387 (N_12387,N_12236,N_12067);
nor U12388 (N_12388,N_12083,N_12100);
nor U12389 (N_12389,N_12171,N_12060);
and U12390 (N_12390,N_12220,N_12127);
or U12391 (N_12391,N_12239,N_12070);
and U12392 (N_12392,N_12119,N_12045);
nor U12393 (N_12393,N_12190,N_12174);
xor U12394 (N_12394,N_12163,N_12210);
nor U12395 (N_12395,N_12053,N_12097);
and U12396 (N_12396,N_12170,N_12109);
or U12397 (N_12397,N_12095,N_12107);
nor U12398 (N_12398,N_12028,N_12194);
and U12399 (N_12399,N_12214,N_12148);
nand U12400 (N_12400,N_12034,N_12112);
or U12401 (N_12401,N_12033,N_12181);
and U12402 (N_12402,N_12193,N_12100);
nand U12403 (N_12403,N_12013,N_12200);
and U12404 (N_12404,N_12124,N_12008);
nand U12405 (N_12405,N_12187,N_12149);
nor U12406 (N_12406,N_12126,N_12216);
nand U12407 (N_12407,N_12193,N_12235);
nand U12408 (N_12408,N_12047,N_12133);
xor U12409 (N_12409,N_12182,N_12112);
nor U12410 (N_12410,N_12240,N_12089);
or U12411 (N_12411,N_12150,N_12206);
nand U12412 (N_12412,N_12223,N_12114);
and U12413 (N_12413,N_12068,N_12094);
or U12414 (N_12414,N_12010,N_12205);
nor U12415 (N_12415,N_12009,N_12064);
and U12416 (N_12416,N_12041,N_12020);
xnor U12417 (N_12417,N_12078,N_12018);
or U12418 (N_12418,N_12015,N_12129);
nor U12419 (N_12419,N_12161,N_12248);
nand U12420 (N_12420,N_12166,N_12048);
nand U12421 (N_12421,N_12101,N_12081);
xnor U12422 (N_12422,N_12036,N_12031);
and U12423 (N_12423,N_12070,N_12122);
and U12424 (N_12424,N_12212,N_12178);
nand U12425 (N_12425,N_12212,N_12063);
nand U12426 (N_12426,N_12023,N_12019);
nand U12427 (N_12427,N_12234,N_12049);
nor U12428 (N_12428,N_12058,N_12102);
xor U12429 (N_12429,N_12216,N_12119);
or U12430 (N_12430,N_12167,N_12096);
and U12431 (N_12431,N_12092,N_12071);
nand U12432 (N_12432,N_12003,N_12229);
and U12433 (N_12433,N_12129,N_12147);
xor U12434 (N_12434,N_12083,N_12163);
or U12435 (N_12435,N_12106,N_12098);
nor U12436 (N_12436,N_12228,N_12076);
nor U12437 (N_12437,N_12153,N_12201);
nand U12438 (N_12438,N_12039,N_12220);
nor U12439 (N_12439,N_12190,N_12240);
nand U12440 (N_12440,N_12169,N_12104);
xor U12441 (N_12441,N_12109,N_12124);
nor U12442 (N_12442,N_12049,N_12051);
nand U12443 (N_12443,N_12168,N_12035);
nand U12444 (N_12444,N_12075,N_12047);
nand U12445 (N_12445,N_12181,N_12121);
xor U12446 (N_12446,N_12034,N_12137);
and U12447 (N_12447,N_12244,N_12177);
and U12448 (N_12448,N_12117,N_12043);
and U12449 (N_12449,N_12042,N_12249);
and U12450 (N_12450,N_12167,N_12166);
and U12451 (N_12451,N_12034,N_12183);
and U12452 (N_12452,N_12138,N_12117);
nand U12453 (N_12453,N_12020,N_12141);
nor U12454 (N_12454,N_12243,N_12069);
or U12455 (N_12455,N_12205,N_12041);
and U12456 (N_12456,N_12154,N_12019);
nand U12457 (N_12457,N_12232,N_12046);
or U12458 (N_12458,N_12081,N_12022);
and U12459 (N_12459,N_12092,N_12100);
or U12460 (N_12460,N_12036,N_12025);
nand U12461 (N_12461,N_12130,N_12065);
nand U12462 (N_12462,N_12214,N_12043);
nand U12463 (N_12463,N_12065,N_12068);
nand U12464 (N_12464,N_12062,N_12090);
and U12465 (N_12465,N_12027,N_12083);
nand U12466 (N_12466,N_12105,N_12006);
nor U12467 (N_12467,N_12205,N_12177);
nor U12468 (N_12468,N_12127,N_12227);
and U12469 (N_12469,N_12156,N_12200);
xor U12470 (N_12470,N_12142,N_12042);
and U12471 (N_12471,N_12029,N_12044);
nor U12472 (N_12472,N_12036,N_12097);
xnor U12473 (N_12473,N_12026,N_12069);
nor U12474 (N_12474,N_12247,N_12194);
nor U12475 (N_12475,N_12079,N_12036);
nor U12476 (N_12476,N_12113,N_12235);
or U12477 (N_12477,N_12182,N_12173);
nor U12478 (N_12478,N_12168,N_12020);
nand U12479 (N_12479,N_12110,N_12190);
or U12480 (N_12480,N_12116,N_12130);
nor U12481 (N_12481,N_12146,N_12212);
and U12482 (N_12482,N_12214,N_12087);
xnor U12483 (N_12483,N_12186,N_12151);
nor U12484 (N_12484,N_12026,N_12131);
nand U12485 (N_12485,N_12007,N_12127);
nor U12486 (N_12486,N_12170,N_12136);
xor U12487 (N_12487,N_12138,N_12209);
and U12488 (N_12488,N_12101,N_12212);
xor U12489 (N_12489,N_12007,N_12010);
nand U12490 (N_12490,N_12156,N_12073);
and U12491 (N_12491,N_12244,N_12235);
nand U12492 (N_12492,N_12080,N_12166);
xor U12493 (N_12493,N_12072,N_12096);
and U12494 (N_12494,N_12173,N_12245);
and U12495 (N_12495,N_12209,N_12034);
nor U12496 (N_12496,N_12181,N_12211);
or U12497 (N_12497,N_12128,N_12244);
xor U12498 (N_12498,N_12071,N_12124);
nand U12499 (N_12499,N_12195,N_12032);
nor U12500 (N_12500,N_12410,N_12341);
or U12501 (N_12501,N_12399,N_12305);
nand U12502 (N_12502,N_12307,N_12395);
or U12503 (N_12503,N_12260,N_12472);
nor U12504 (N_12504,N_12499,N_12487);
nand U12505 (N_12505,N_12477,N_12425);
nand U12506 (N_12506,N_12436,N_12350);
nand U12507 (N_12507,N_12388,N_12417);
or U12508 (N_12508,N_12349,N_12361);
nor U12509 (N_12509,N_12408,N_12476);
and U12510 (N_12510,N_12366,N_12462);
xor U12511 (N_12511,N_12489,N_12494);
xnor U12512 (N_12512,N_12398,N_12413);
nand U12513 (N_12513,N_12383,N_12284);
nor U12514 (N_12514,N_12327,N_12493);
nand U12515 (N_12515,N_12345,N_12274);
and U12516 (N_12516,N_12406,N_12467);
or U12517 (N_12517,N_12365,N_12432);
nor U12518 (N_12518,N_12315,N_12490);
and U12519 (N_12519,N_12459,N_12468);
and U12520 (N_12520,N_12443,N_12278);
nand U12521 (N_12521,N_12266,N_12412);
nand U12522 (N_12522,N_12497,N_12479);
or U12523 (N_12523,N_12452,N_12288);
or U12524 (N_12524,N_12407,N_12294);
and U12525 (N_12525,N_12251,N_12348);
xor U12526 (N_12526,N_12323,N_12470);
nand U12527 (N_12527,N_12358,N_12469);
xnor U12528 (N_12528,N_12279,N_12332);
nor U12529 (N_12529,N_12411,N_12331);
xnor U12530 (N_12530,N_12387,N_12367);
nor U12531 (N_12531,N_12415,N_12391);
nor U12532 (N_12532,N_12324,N_12355);
or U12533 (N_12533,N_12492,N_12280);
or U12534 (N_12534,N_12314,N_12329);
xor U12535 (N_12535,N_12380,N_12440);
xnor U12536 (N_12536,N_12256,N_12491);
and U12537 (N_12537,N_12330,N_12337);
nand U12538 (N_12538,N_12420,N_12351);
xnor U12539 (N_12539,N_12379,N_12306);
nor U12540 (N_12540,N_12453,N_12302);
xnor U12541 (N_12541,N_12297,N_12496);
nor U12542 (N_12542,N_12336,N_12334);
or U12543 (N_12543,N_12363,N_12333);
nor U12544 (N_12544,N_12449,N_12301);
or U12545 (N_12545,N_12498,N_12291);
and U12546 (N_12546,N_12483,N_12360);
or U12547 (N_12547,N_12396,N_12254);
and U12548 (N_12548,N_12326,N_12478);
or U12549 (N_12549,N_12354,N_12255);
xor U12550 (N_12550,N_12343,N_12375);
nor U12551 (N_12551,N_12454,N_12403);
or U12552 (N_12552,N_12438,N_12346);
or U12553 (N_12553,N_12419,N_12313);
nor U12554 (N_12554,N_12441,N_12356);
nor U12555 (N_12555,N_12252,N_12339);
and U12556 (N_12556,N_12290,N_12289);
nor U12557 (N_12557,N_12261,N_12269);
nor U12558 (N_12558,N_12271,N_12299);
xor U12559 (N_12559,N_12482,N_12265);
or U12560 (N_12560,N_12258,N_12286);
and U12561 (N_12561,N_12393,N_12295);
and U12562 (N_12562,N_12404,N_12342);
xnor U12563 (N_12563,N_12485,N_12451);
xor U12564 (N_12564,N_12385,N_12303);
xnor U12565 (N_12565,N_12424,N_12319);
xnor U12566 (N_12566,N_12262,N_12465);
or U12567 (N_12567,N_12296,N_12283);
nand U12568 (N_12568,N_12409,N_12400);
and U12569 (N_12569,N_12448,N_12352);
and U12570 (N_12570,N_12414,N_12422);
and U12571 (N_12571,N_12257,N_12473);
nand U12572 (N_12572,N_12416,N_12372);
or U12573 (N_12573,N_12389,N_12481);
and U12574 (N_12574,N_12357,N_12369);
and U12575 (N_12575,N_12359,N_12430);
xor U12576 (N_12576,N_12457,N_12464);
nand U12577 (N_12577,N_12370,N_12384);
and U12578 (N_12578,N_12486,N_12328);
xor U12579 (N_12579,N_12321,N_12287);
xnor U12580 (N_12580,N_12347,N_12276);
nor U12581 (N_12581,N_12401,N_12427);
or U12582 (N_12582,N_12433,N_12377);
nand U12583 (N_12583,N_12277,N_12405);
or U12584 (N_12584,N_12435,N_12281);
or U12585 (N_12585,N_12471,N_12397);
or U12586 (N_12586,N_12378,N_12312);
or U12587 (N_12587,N_12394,N_12322);
xnor U12588 (N_12588,N_12442,N_12381);
nor U12589 (N_12589,N_12317,N_12371);
xnor U12590 (N_12590,N_12429,N_12318);
nor U12591 (N_12591,N_12418,N_12466);
nor U12592 (N_12592,N_12353,N_12392);
or U12593 (N_12593,N_12364,N_12458);
nand U12594 (N_12594,N_12460,N_12316);
xnor U12595 (N_12595,N_12428,N_12423);
and U12596 (N_12596,N_12495,N_12463);
and U12597 (N_12597,N_12310,N_12444);
nand U12598 (N_12598,N_12386,N_12275);
or U12599 (N_12599,N_12268,N_12376);
nor U12600 (N_12600,N_12285,N_12325);
xor U12601 (N_12601,N_12390,N_12272);
and U12602 (N_12602,N_12270,N_12421);
and U12603 (N_12603,N_12282,N_12344);
nand U12604 (N_12604,N_12308,N_12450);
or U12605 (N_12605,N_12426,N_12446);
nor U12606 (N_12606,N_12304,N_12456);
xnor U12607 (N_12607,N_12488,N_12402);
nand U12608 (N_12608,N_12382,N_12461);
nor U12609 (N_12609,N_12368,N_12480);
nand U12610 (N_12610,N_12338,N_12253);
or U12611 (N_12611,N_12374,N_12259);
nor U12612 (N_12612,N_12439,N_12434);
or U12613 (N_12613,N_12362,N_12335);
xor U12614 (N_12614,N_12431,N_12475);
xnor U12615 (N_12615,N_12311,N_12320);
or U12616 (N_12616,N_12298,N_12373);
and U12617 (N_12617,N_12250,N_12309);
or U12618 (N_12618,N_12263,N_12273);
nand U12619 (N_12619,N_12437,N_12267);
nand U12620 (N_12620,N_12340,N_12264);
nor U12621 (N_12621,N_12484,N_12445);
nand U12622 (N_12622,N_12293,N_12455);
xnor U12623 (N_12623,N_12447,N_12292);
nand U12624 (N_12624,N_12300,N_12474);
nand U12625 (N_12625,N_12294,N_12331);
nand U12626 (N_12626,N_12351,N_12470);
and U12627 (N_12627,N_12355,N_12464);
and U12628 (N_12628,N_12489,N_12482);
nor U12629 (N_12629,N_12485,N_12435);
or U12630 (N_12630,N_12335,N_12424);
and U12631 (N_12631,N_12291,N_12410);
or U12632 (N_12632,N_12355,N_12377);
xor U12633 (N_12633,N_12435,N_12258);
xnor U12634 (N_12634,N_12337,N_12401);
nand U12635 (N_12635,N_12473,N_12471);
nor U12636 (N_12636,N_12279,N_12320);
xnor U12637 (N_12637,N_12345,N_12468);
nor U12638 (N_12638,N_12340,N_12271);
nand U12639 (N_12639,N_12346,N_12419);
xnor U12640 (N_12640,N_12283,N_12267);
nand U12641 (N_12641,N_12309,N_12369);
and U12642 (N_12642,N_12323,N_12326);
nand U12643 (N_12643,N_12422,N_12486);
nor U12644 (N_12644,N_12355,N_12475);
and U12645 (N_12645,N_12470,N_12325);
or U12646 (N_12646,N_12274,N_12313);
nor U12647 (N_12647,N_12431,N_12419);
xor U12648 (N_12648,N_12255,N_12300);
and U12649 (N_12649,N_12340,N_12412);
or U12650 (N_12650,N_12264,N_12315);
nand U12651 (N_12651,N_12334,N_12280);
or U12652 (N_12652,N_12362,N_12320);
and U12653 (N_12653,N_12383,N_12365);
nand U12654 (N_12654,N_12273,N_12426);
and U12655 (N_12655,N_12270,N_12317);
nand U12656 (N_12656,N_12384,N_12257);
and U12657 (N_12657,N_12260,N_12313);
nor U12658 (N_12658,N_12496,N_12483);
or U12659 (N_12659,N_12272,N_12298);
xor U12660 (N_12660,N_12346,N_12372);
nor U12661 (N_12661,N_12292,N_12290);
and U12662 (N_12662,N_12450,N_12283);
or U12663 (N_12663,N_12482,N_12344);
nand U12664 (N_12664,N_12413,N_12310);
and U12665 (N_12665,N_12298,N_12324);
xor U12666 (N_12666,N_12324,N_12323);
xor U12667 (N_12667,N_12370,N_12471);
nor U12668 (N_12668,N_12330,N_12499);
nand U12669 (N_12669,N_12345,N_12333);
or U12670 (N_12670,N_12307,N_12348);
nand U12671 (N_12671,N_12403,N_12451);
and U12672 (N_12672,N_12391,N_12342);
xnor U12673 (N_12673,N_12257,N_12485);
xor U12674 (N_12674,N_12376,N_12437);
and U12675 (N_12675,N_12278,N_12285);
or U12676 (N_12676,N_12411,N_12293);
nand U12677 (N_12677,N_12462,N_12396);
xor U12678 (N_12678,N_12313,N_12489);
nor U12679 (N_12679,N_12382,N_12264);
nand U12680 (N_12680,N_12420,N_12433);
or U12681 (N_12681,N_12487,N_12256);
and U12682 (N_12682,N_12427,N_12302);
nor U12683 (N_12683,N_12484,N_12286);
nor U12684 (N_12684,N_12384,N_12325);
xor U12685 (N_12685,N_12250,N_12452);
nor U12686 (N_12686,N_12311,N_12485);
xnor U12687 (N_12687,N_12310,N_12454);
or U12688 (N_12688,N_12431,N_12344);
or U12689 (N_12689,N_12393,N_12431);
and U12690 (N_12690,N_12441,N_12250);
and U12691 (N_12691,N_12266,N_12414);
xor U12692 (N_12692,N_12320,N_12489);
xnor U12693 (N_12693,N_12417,N_12430);
or U12694 (N_12694,N_12427,N_12310);
nor U12695 (N_12695,N_12417,N_12475);
and U12696 (N_12696,N_12343,N_12319);
or U12697 (N_12697,N_12482,N_12287);
or U12698 (N_12698,N_12451,N_12307);
nand U12699 (N_12699,N_12379,N_12440);
nand U12700 (N_12700,N_12382,N_12488);
and U12701 (N_12701,N_12359,N_12331);
and U12702 (N_12702,N_12471,N_12344);
and U12703 (N_12703,N_12359,N_12305);
or U12704 (N_12704,N_12446,N_12350);
nor U12705 (N_12705,N_12365,N_12450);
nand U12706 (N_12706,N_12440,N_12264);
nand U12707 (N_12707,N_12327,N_12319);
and U12708 (N_12708,N_12447,N_12489);
xor U12709 (N_12709,N_12413,N_12304);
or U12710 (N_12710,N_12289,N_12441);
nor U12711 (N_12711,N_12459,N_12385);
xor U12712 (N_12712,N_12400,N_12405);
or U12713 (N_12713,N_12256,N_12274);
nor U12714 (N_12714,N_12364,N_12483);
nor U12715 (N_12715,N_12460,N_12362);
nor U12716 (N_12716,N_12480,N_12327);
nor U12717 (N_12717,N_12495,N_12379);
nor U12718 (N_12718,N_12488,N_12369);
or U12719 (N_12719,N_12274,N_12322);
or U12720 (N_12720,N_12343,N_12469);
or U12721 (N_12721,N_12378,N_12448);
xor U12722 (N_12722,N_12260,N_12461);
xnor U12723 (N_12723,N_12261,N_12406);
xor U12724 (N_12724,N_12363,N_12257);
nand U12725 (N_12725,N_12438,N_12487);
or U12726 (N_12726,N_12315,N_12275);
xnor U12727 (N_12727,N_12408,N_12299);
nor U12728 (N_12728,N_12320,N_12450);
nand U12729 (N_12729,N_12402,N_12461);
nand U12730 (N_12730,N_12475,N_12353);
nand U12731 (N_12731,N_12484,N_12392);
or U12732 (N_12732,N_12421,N_12456);
nand U12733 (N_12733,N_12355,N_12291);
and U12734 (N_12734,N_12297,N_12393);
xnor U12735 (N_12735,N_12463,N_12355);
nor U12736 (N_12736,N_12388,N_12399);
xnor U12737 (N_12737,N_12478,N_12290);
and U12738 (N_12738,N_12297,N_12356);
xor U12739 (N_12739,N_12432,N_12421);
nor U12740 (N_12740,N_12250,N_12353);
xor U12741 (N_12741,N_12422,N_12344);
xnor U12742 (N_12742,N_12258,N_12379);
xor U12743 (N_12743,N_12272,N_12420);
nor U12744 (N_12744,N_12445,N_12477);
nor U12745 (N_12745,N_12492,N_12309);
nand U12746 (N_12746,N_12374,N_12415);
nand U12747 (N_12747,N_12308,N_12304);
and U12748 (N_12748,N_12431,N_12322);
nand U12749 (N_12749,N_12384,N_12333);
nand U12750 (N_12750,N_12744,N_12510);
nor U12751 (N_12751,N_12600,N_12711);
nand U12752 (N_12752,N_12738,N_12676);
nor U12753 (N_12753,N_12622,N_12748);
nand U12754 (N_12754,N_12616,N_12532);
or U12755 (N_12755,N_12705,N_12728);
or U12756 (N_12756,N_12673,N_12507);
nor U12757 (N_12757,N_12591,N_12652);
or U12758 (N_12758,N_12694,N_12533);
xor U12759 (N_12759,N_12566,N_12597);
and U12760 (N_12760,N_12730,N_12624);
or U12761 (N_12761,N_12679,N_12731);
nor U12762 (N_12762,N_12604,N_12550);
xor U12763 (N_12763,N_12669,N_12675);
nor U12764 (N_12764,N_12564,N_12653);
xor U12765 (N_12765,N_12603,N_12677);
and U12766 (N_12766,N_12658,N_12538);
nand U12767 (N_12767,N_12617,N_12506);
nand U12768 (N_12768,N_12580,N_12723);
or U12769 (N_12769,N_12559,N_12640);
xnor U12770 (N_12770,N_12635,N_12553);
nand U12771 (N_12771,N_12556,N_12722);
xnor U12772 (N_12772,N_12696,N_12557);
nor U12773 (N_12773,N_12554,N_12613);
nor U12774 (N_12774,N_12645,N_12607);
or U12775 (N_12775,N_12671,N_12663);
or U12776 (N_12776,N_12590,N_12701);
xor U12777 (N_12777,N_12601,N_12514);
xnor U12778 (N_12778,N_12724,N_12531);
nor U12779 (N_12779,N_12664,N_12749);
or U12780 (N_12780,N_12593,N_12708);
or U12781 (N_12781,N_12643,N_12560);
and U12782 (N_12782,N_12699,N_12598);
xor U12783 (N_12783,N_12648,N_12636);
nand U12784 (N_12784,N_12715,N_12686);
and U12785 (N_12785,N_12612,N_12546);
nor U12786 (N_12786,N_12570,N_12541);
xor U12787 (N_12787,N_12583,N_12646);
nand U12788 (N_12788,N_12644,N_12615);
or U12789 (N_12789,N_12516,N_12727);
nand U12790 (N_12790,N_12528,N_12621);
xor U12791 (N_12791,N_12618,N_12626);
nor U12792 (N_12792,N_12569,N_12692);
xnor U12793 (N_12793,N_12567,N_12695);
nor U12794 (N_12794,N_12627,N_12513);
xor U12795 (N_12795,N_12501,N_12525);
nand U12796 (N_12796,N_12562,N_12742);
and U12797 (N_12797,N_12691,N_12595);
and U12798 (N_12798,N_12681,N_12561);
and U12799 (N_12799,N_12670,N_12706);
xnor U12800 (N_12800,N_12697,N_12521);
nand U12801 (N_12801,N_12656,N_12734);
xor U12802 (N_12802,N_12629,N_12678);
xor U12803 (N_12803,N_12743,N_12642);
xnor U12804 (N_12804,N_12729,N_12606);
or U12805 (N_12805,N_12707,N_12641);
and U12806 (N_12806,N_12565,N_12548);
xnor U12807 (N_12807,N_12505,N_12737);
and U12808 (N_12808,N_12605,N_12667);
or U12809 (N_12809,N_12526,N_12584);
or U12810 (N_12810,N_12582,N_12746);
or U12811 (N_12811,N_12610,N_12709);
and U12812 (N_12812,N_12578,N_12574);
or U12813 (N_12813,N_12551,N_12623);
nor U12814 (N_12814,N_12575,N_12581);
nor U12815 (N_12815,N_12576,N_12540);
nor U12816 (N_12816,N_12502,N_12745);
xor U12817 (N_12817,N_12589,N_12682);
and U12818 (N_12818,N_12536,N_12572);
or U12819 (N_12819,N_12608,N_12563);
and U12820 (N_12820,N_12573,N_12544);
and U12821 (N_12821,N_12649,N_12545);
or U12822 (N_12822,N_12638,N_12721);
nand U12823 (N_12823,N_12713,N_12614);
or U12824 (N_12824,N_12655,N_12535);
and U12825 (N_12825,N_12518,N_12720);
or U12826 (N_12826,N_12704,N_12587);
xnor U12827 (N_12827,N_12523,N_12647);
nand U12828 (N_12828,N_12555,N_12735);
and U12829 (N_12829,N_12719,N_12579);
xor U12830 (N_12830,N_12500,N_12508);
nor U12831 (N_12831,N_12628,N_12739);
xor U12832 (N_12832,N_12674,N_12586);
xor U12833 (N_12833,N_12637,N_12588);
xnor U12834 (N_12834,N_12710,N_12539);
xor U12835 (N_12835,N_12747,N_12702);
or U12836 (N_12836,N_12680,N_12568);
or U12837 (N_12837,N_12689,N_12650);
xor U12838 (N_12838,N_12602,N_12558);
xnor U12839 (N_12839,N_12661,N_12524);
or U12840 (N_12840,N_12620,N_12662);
and U12841 (N_12841,N_12683,N_12611);
nand U12842 (N_12842,N_12668,N_12741);
and U12843 (N_12843,N_12672,N_12633);
xnor U12844 (N_12844,N_12592,N_12726);
nand U12845 (N_12845,N_12712,N_12527);
xnor U12846 (N_12846,N_12736,N_12740);
xor U12847 (N_12847,N_12690,N_12609);
xnor U12848 (N_12848,N_12549,N_12511);
xor U12849 (N_12849,N_12639,N_12619);
xor U12850 (N_12850,N_12630,N_12543);
and U12851 (N_12851,N_12688,N_12717);
or U12852 (N_12852,N_12529,N_12651);
xor U12853 (N_12853,N_12520,N_12714);
nand U12854 (N_12854,N_12657,N_12504);
nor U12855 (N_12855,N_12517,N_12700);
xnor U12856 (N_12856,N_12732,N_12512);
or U12857 (N_12857,N_12537,N_12665);
nor U12858 (N_12858,N_12733,N_12659);
nor U12859 (N_12859,N_12666,N_12698);
nand U12860 (N_12860,N_12631,N_12634);
xor U12861 (N_12861,N_12522,N_12596);
or U12862 (N_12862,N_12625,N_12684);
and U12863 (N_12863,N_12509,N_12654);
or U12864 (N_12864,N_12534,N_12716);
nor U12865 (N_12865,N_12594,N_12577);
xor U12866 (N_12866,N_12599,N_12660);
and U12867 (N_12867,N_12585,N_12515);
nor U12868 (N_12868,N_12519,N_12687);
nand U12869 (N_12869,N_12547,N_12685);
xnor U12870 (N_12870,N_12725,N_12530);
and U12871 (N_12871,N_12571,N_12503);
nor U12872 (N_12872,N_12552,N_12718);
xor U12873 (N_12873,N_12632,N_12542);
nor U12874 (N_12874,N_12703,N_12693);
or U12875 (N_12875,N_12536,N_12720);
xor U12876 (N_12876,N_12637,N_12530);
or U12877 (N_12877,N_12590,N_12747);
nand U12878 (N_12878,N_12574,N_12736);
and U12879 (N_12879,N_12683,N_12685);
xnor U12880 (N_12880,N_12685,N_12746);
and U12881 (N_12881,N_12641,N_12635);
nand U12882 (N_12882,N_12736,N_12683);
and U12883 (N_12883,N_12645,N_12736);
nor U12884 (N_12884,N_12722,N_12553);
nand U12885 (N_12885,N_12659,N_12690);
and U12886 (N_12886,N_12646,N_12718);
xor U12887 (N_12887,N_12571,N_12583);
xnor U12888 (N_12888,N_12627,N_12653);
or U12889 (N_12889,N_12614,N_12618);
nand U12890 (N_12890,N_12588,N_12585);
and U12891 (N_12891,N_12526,N_12683);
or U12892 (N_12892,N_12609,N_12748);
and U12893 (N_12893,N_12550,N_12573);
and U12894 (N_12894,N_12645,N_12575);
or U12895 (N_12895,N_12676,N_12599);
or U12896 (N_12896,N_12643,N_12527);
and U12897 (N_12897,N_12670,N_12660);
or U12898 (N_12898,N_12705,N_12677);
or U12899 (N_12899,N_12691,N_12630);
and U12900 (N_12900,N_12567,N_12644);
nor U12901 (N_12901,N_12688,N_12537);
nor U12902 (N_12902,N_12542,N_12618);
and U12903 (N_12903,N_12694,N_12500);
or U12904 (N_12904,N_12557,N_12565);
or U12905 (N_12905,N_12541,N_12686);
xnor U12906 (N_12906,N_12711,N_12606);
nand U12907 (N_12907,N_12505,N_12523);
or U12908 (N_12908,N_12709,N_12655);
nor U12909 (N_12909,N_12661,N_12598);
nor U12910 (N_12910,N_12623,N_12715);
nand U12911 (N_12911,N_12553,N_12701);
or U12912 (N_12912,N_12564,N_12701);
and U12913 (N_12913,N_12671,N_12548);
or U12914 (N_12914,N_12591,N_12706);
xor U12915 (N_12915,N_12670,N_12734);
nor U12916 (N_12916,N_12664,N_12701);
or U12917 (N_12917,N_12639,N_12577);
nand U12918 (N_12918,N_12609,N_12636);
nand U12919 (N_12919,N_12687,N_12547);
xnor U12920 (N_12920,N_12730,N_12675);
nand U12921 (N_12921,N_12688,N_12576);
xnor U12922 (N_12922,N_12577,N_12570);
nand U12923 (N_12923,N_12678,N_12554);
or U12924 (N_12924,N_12514,N_12738);
or U12925 (N_12925,N_12702,N_12628);
nand U12926 (N_12926,N_12655,N_12589);
xnor U12927 (N_12927,N_12630,N_12668);
nor U12928 (N_12928,N_12609,N_12618);
nor U12929 (N_12929,N_12578,N_12647);
or U12930 (N_12930,N_12546,N_12600);
and U12931 (N_12931,N_12573,N_12567);
and U12932 (N_12932,N_12608,N_12544);
nand U12933 (N_12933,N_12620,N_12733);
xor U12934 (N_12934,N_12563,N_12722);
or U12935 (N_12935,N_12694,N_12670);
nor U12936 (N_12936,N_12743,N_12737);
and U12937 (N_12937,N_12678,N_12529);
xnor U12938 (N_12938,N_12642,N_12580);
nand U12939 (N_12939,N_12535,N_12716);
nor U12940 (N_12940,N_12684,N_12615);
and U12941 (N_12941,N_12557,N_12502);
and U12942 (N_12942,N_12716,N_12621);
xor U12943 (N_12943,N_12684,N_12705);
nor U12944 (N_12944,N_12538,N_12732);
xor U12945 (N_12945,N_12504,N_12531);
and U12946 (N_12946,N_12691,N_12610);
nor U12947 (N_12947,N_12569,N_12749);
xnor U12948 (N_12948,N_12744,N_12647);
or U12949 (N_12949,N_12581,N_12535);
or U12950 (N_12950,N_12558,N_12648);
xnor U12951 (N_12951,N_12500,N_12538);
or U12952 (N_12952,N_12590,N_12675);
nor U12953 (N_12953,N_12579,N_12706);
xor U12954 (N_12954,N_12600,N_12513);
and U12955 (N_12955,N_12603,N_12651);
or U12956 (N_12956,N_12575,N_12745);
nand U12957 (N_12957,N_12625,N_12673);
nand U12958 (N_12958,N_12721,N_12524);
and U12959 (N_12959,N_12635,N_12709);
or U12960 (N_12960,N_12686,N_12691);
xnor U12961 (N_12961,N_12656,N_12514);
xnor U12962 (N_12962,N_12607,N_12565);
nand U12963 (N_12963,N_12733,N_12691);
nand U12964 (N_12964,N_12680,N_12709);
xor U12965 (N_12965,N_12701,N_12726);
nor U12966 (N_12966,N_12573,N_12520);
nand U12967 (N_12967,N_12654,N_12546);
or U12968 (N_12968,N_12709,N_12708);
nand U12969 (N_12969,N_12627,N_12698);
xor U12970 (N_12970,N_12747,N_12654);
nor U12971 (N_12971,N_12552,N_12730);
xor U12972 (N_12972,N_12667,N_12650);
nand U12973 (N_12973,N_12560,N_12676);
and U12974 (N_12974,N_12668,N_12551);
or U12975 (N_12975,N_12644,N_12620);
or U12976 (N_12976,N_12530,N_12511);
or U12977 (N_12977,N_12533,N_12680);
nor U12978 (N_12978,N_12594,N_12660);
xnor U12979 (N_12979,N_12721,N_12739);
and U12980 (N_12980,N_12556,N_12595);
or U12981 (N_12981,N_12568,N_12606);
xnor U12982 (N_12982,N_12563,N_12596);
nor U12983 (N_12983,N_12623,N_12548);
nor U12984 (N_12984,N_12653,N_12684);
nand U12985 (N_12985,N_12524,N_12588);
and U12986 (N_12986,N_12679,N_12596);
or U12987 (N_12987,N_12603,N_12564);
nor U12988 (N_12988,N_12592,N_12602);
nand U12989 (N_12989,N_12524,N_12693);
and U12990 (N_12990,N_12703,N_12641);
or U12991 (N_12991,N_12524,N_12582);
nand U12992 (N_12992,N_12528,N_12665);
nand U12993 (N_12993,N_12512,N_12602);
xnor U12994 (N_12994,N_12625,N_12550);
nand U12995 (N_12995,N_12599,N_12607);
nand U12996 (N_12996,N_12645,N_12677);
nor U12997 (N_12997,N_12689,N_12725);
nor U12998 (N_12998,N_12631,N_12517);
xor U12999 (N_12999,N_12593,N_12580);
xor U13000 (N_13000,N_12837,N_12964);
or U13001 (N_13001,N_12792,N_12882);
and U13002 (N_13002,N_12914,N_12800);
or U13003 (N_13003,N_12853,N_12993);
or U13004 (N_13004,N_12859,N_12971);
and U13005 (N_13005,N_12954,N_12847);
nor U13006 (N_13006,N_12835,N_12848);
xnor U13007 (N_13007,N_12825,N_12927);
nand U13008 (N_13008,N_12884,N_12981);
nor U13009 (N_13009,N_12929,N_12975);
nor U13010 (N_13010,N_12955,N_12881);
or U13011 (N_13011,N_12987,N_12810);
xnor U13012 (N_13012,N_12811,N_12933);
nor U13013 (N_13013,N_12753,N_12879);
nand U13014 (N_13014,N_12969,N_12889);
nor U13015 (N_13015,N_12928,N_12867);
and U13016 (N_13016,N_12819,N_12963);
nand U13017 (N_13017,N_12911,N_12768);
and U13018 (N_13018,N_12909,N_12766);
and U13019 (N_13019,N_12828,N_12961);
and U13020 (N_13020,N_12874,N_12862);
xor U13021 (N_13021,N_12946,N_12787);
xnor U13022 (N_13022,N_12843,N_12888);
nor U13023 (N_13023,N_12988,N_12842);
xor U13024 (N_13024,N_12932,N_12930);
nand U13025 (N_13025,N_12901,N_12935);
nor U13026 (N_13026,N_12934,N_12892);
nor U13027 (N_13027,N_12827,N_12947);
or U13028 (N_13028,N_12951,N_12856);
nand U13029 (N_13029,N_12801,N_12960);
and U13030 (N_13030,N_12985,N_12878);
or U13031 (N_13031,N_12832,N_12786);
or U13032 (N_13032,N_12940,N_12887);
or U13033 (N_13033,N_12751,N_12922);
xnor U13034 (N_13034,N_12861,N_12994);
xnor U13035 (N_13035,N_12880,N_12770);
nand U13036 (N_13036,N_12841,N_12952);
nand U13037 (N_13037,N_12936,N_12844);
nand U13038 (N_13038,N_12858,N_12808);
and U13039 (N_13039,N_12817,N_12986);
or U13040 (N_13040,N_12802,N_12763);
or U13041 (N_13041,N_12899,N_12760);
and U13042 (N_13042,N_12794,N_12823);
xnor U13043 (N_13043,N_12807,N_12761);
xor U13044 (N_13044,N_12949,N_12815);
xnor U13045 (N_13045,N_12758,N_12915);
or U13046 (N_13046,N_12854,N_12958);
and U13047 (N_13047,N_12957,N_12798);
and U13048 (N_13048,N_12978,N_12972);
nand U13049 (N_13049,N_12764,N_12908);
or U13050 (N_13050,N_12780,N_12883);
nor U13051 (N_13051,N_12891,N_12939);
and U13052 (N_13052,N_12918,N_12829);
and U13053 (N_13053,N_12970,N_12795);
nor U13054 (N_13054,N_12872,N_12974);
or U13055 (N_13055,N_12779,N_12750);
nor U13056 (N_13056,N_12839,N_12793);
nand U13057 (N_13057,N_12845,N_12885);
nor U13058 (N_13058,N_12789,N_12756);
or U13059 (N_13059,N_12991,N_12890);
xnor U13060 (N_13060,N_12776,N_12875);
nand U13061 (N_13061,N_12781,N_12757);
nand U13062 (N_13062,N_12945,N_12864);
nand U13063 (N_13063,N_12996,N_12990);
xor U13064 (N_13064,N_12788,N_12834);
and U13065 (N_13065,N_12809,N_12956);
or U13066 (N_13066,N_12762,N_12923);
xnor U13067 (N_13067,N_12860,N_12796);
nand U13068 (N_13068,N_12775,N_12886);
or U13069 (N_13069,N_12799,N_12919);
xor U13070 (N_13070,N_12850,N_12903);
xnor U13071 (N_13071,N_12950,N_12852);
nor U13072 (N_13072,N_12824,N_12965);
and U13073 (N_13073,N_12962,N_12765);
nor U13074 (N_13074,N_12821,N_12980);
nor U13075 (N_13075,N_12782,N_12912);
nor U13076 (N_13076,N_12998,N_12755);
nor U13077 (N_13077,N_12959,N_12902);
or U13078 (N_13078,N_12921,N_12948);
or U13079 (N_13079,N_12791,N_12797);
or U13080 (N_13080,N_12924,N_12846);
xor U13081 (N_13081,N_12865,N_12943);
and U13082 (N_13082,N_12778,N_12773);
or U13083 (N_13083,N_12966,N_12840);
or U13084 (N_13084,N_12866,N_12941);
or U13085 (N_13085,N_12893,N_12754);
or U13086 (N_13086,N_12830,N_12999);
and U13087 (N_13087,N_12868,N_12905);
or U13088 (N_13088,N_12831,N_12989);
nor U13089 (N_13089,N_12937,N_12752);
nor U13090 (N_13090,N_12806,N_12838);
and U13091 (N_13091,N_12863,N_12805);
nand U13092 (N_13092,N_12979,N_12977);
or U13093 (N_13093,N_12876,N_12820);
nor U13094 (N_13094,N_12995,N_12783);
or U13095 (N_13095,N_12925,N_12976);
nor U13096 (N_13096,N_12897,N_12992);
or U13097 (N_13097,N_12913,N_12772);
and U13098 (N_13098,N_12953,N_12784);
or U13099 (N_13099,N_12833,N_12822);
and U13100 (N_13100,N_12851,N_12869);
or U13101 (N_13101,N_12818,N_12973);
nand U13102 (N_13102,N_12894,N_12898);
xnor U13103 (N_13103,N_12813,N_12931);
and U13104 (N_13104,N_12826,N_12771);
nand U13105 (N_13105,N_12855,N_12871);
or U13106 (N_13106,N_12769,N_12857);
and U13107 (N_13107,N_12836,N_12812);
nor U13108 (N_13108,N_12926,N_12814);
xnor U13109 (N_13109,N_12900,N_12816);
nand U13110 (N_13110,N_12906,N_12849);
and U13111 (N_13111,N_12873,N_12803);
xor U13112 (N_13112,N_12785,N_12920);
xnor U13113 (N_13113,N_12777,N_12997);
or U13114 (N_13114,N_12942,N_12870);
xor U13115 (N_13115,N_12907,N_12904);
xor U13116 (N_13116,N_12917,N_12790);
or U13117 (N_13117,N_12896,N_12910);
nand U13118 (N_13118,N_12916,N_12877);
and U13119 (N_13119,N_12767,N_12774);
and U13120 (N_13120,N_12967,N_12938);
and U13121 (N_13121,N_12944,N_12983);
or U13122 (N_13122,N_12895,N_12968);
nand U13123 (N_13123,N_12804,N_12984);
and U13124 (N_13124,N_12759,N_12982);
nor U13125 (N_13125,N_12798,N_12835);
xor U13126 (N_13126,N_12827,N_12845);
nor U13127 (N_13127,N_12778,N_12900);
or U13128 (N_13128,N_12900,N_12862);
nor U13129 (N_13129,N_12837,N_12792);
nand U13130 (N_13130,N_12884,N_12984);
xor U13131 (N_13131,N_12943,N_12983);
nand U13132 (N_13132,N_12867,N_12750);
nor U13133 (N_13133,N_12843,N_12880);
nor U13134 (N_13134,N_12921,N_12755);
xor U13135 (N_13135,N_12943,N_12805);
and U13136 (N_13136,N_12928,N_12768);
nand U13137 (N_13137,N_12792,N_12902);
nand U13138 (N_13138,N_12823,N_12751);
and U13139 (N_13139,N_12928,N_12955);
nand U13140 (N_13140,N_12835,N_12904);
or U13141 (N_13141,N_12898,N_12791);
or U13142 (N_13142,N_12828,N_12765);
nand U13143 (N_13143,N_12805,N_12971);
or U13144 (N_13144,N_12898,N_12961);
or U13145 (N_13145,N_12842,N_12755);
xnor U13146 (N_13146,N_12793,N_12936);
nor U13147 (N_13147,N_12918,N_12949);
or U13148 (N_13148,N_12956,N_12957);
xor U13149 (N_13149,N_12957,N_12924);
nor U13150 (N_13150,N_12998,N_12845);
xor U13151 (N_13151,N_12943,N_12807);
or U13152 (N_13152,N_12806,N_12832);
xnor U13153 (N_13153,N_12902,N_12894);
xor U13154 (N_13154,N_12914,N_12992);
xnor U13155 (N_13155,N_12933,N_12791);
nor U13156 (N_13156,N_12970,N_12972);
xor U13157 (N_13157,N_12876,N_12765);
xnor U13158 (N_13158,N_12795,N_12804);
or U13159 (N_13159,N_12760,N_12959);
or U13160 (N_13160,N_12802,N_12974);
and U13161 (N_13161,N_12975,N_12985);
xnor U13162 (N_13162,N_12835,N_12884);
xnor U13163 (N_13163,N_12906,N_12851);
nor U13164 (N_13164,N_12837,N_12923);
nand U13165 (N_13165,N_12966,N_12858);
and U13166 (N_13166,N_12866,N_12991);
xnor U13167 (N_13167,N_12879,N_12843);
xnor U13168 (N_13168,N_12786,N_12917);
nand U13169 (N_13169,N_12932,N_12888);
xnor U13170 (N_13170,N_12848,N_12815);
nor U13171 (N_13171,N_12997,N_12839);
or U13172 (N_13172,N_12932,N_12986);
and U13173 (N_13173,N_12813,N_12756);
and U13174 (N_13174,N_12802,N_12928);
xnor U13175 (N_13175,N_12827,N_12946);
nor U13176 (N_13176,N_12885,N_12963);
or U13177 (N_13177,N_12894,N_12760);
or U13178 (N_13178,N_12849,N_12752);
nand U13179 (N_13179,N_12975,N_12890);
or U13180 (N_13180,N_12793,N_12979);
xor U13181 (N_13181,N_12979,N_12780);
and U13182 (N_13182,N_12849,N_12862);
nor U13183 (N_13183,N_12936,N_12788);
nand U13184 (N_13184,N_12854,N_12980);
or U13185 (N_13185,N_12934,N_12875);
or U13186 (N_13186,N_12986,N_12990);
or U13187 (N_13187,N_12971,N_12882);
and U13188 (N_13188,N_12903,N_12930);
or U13189 (N_13189,N_12798,N_12765);
nor U13190 (N_13190,N_12842,N_12946);
nor U13191 (N_13191,N_12857,N_12761);
and U13192 (N_13192,N_12972,N_12808);
nor U13193 (N_13193,N_12861,N_12973);
nand U13194 (N_13194,N_12874,N_12956);
xor U13195 (N_13195,N_12961,N_12842);
and U13196 (N_13196,N_12865,N_12866);
xnor U13197 (N_13197,N_12828,N_12782);
nand U13198 (N_13198,N_12801,N_12812);
and U13199 (N_13199,N_12787,N_12988);
nor U13200 (N_13200,N_12854,N_12772);
and U13201 (N_13201,N_12963,N_12932);
nand U13202 (N_13202,N_12987,N_12885);
nor U13203 (N_13203,N_12875,N_12786);
xnor U13204 (N_13204,N_12791,N_12819);
xnor U13205 (N_13205,N_12757,N_12837);
nor U13206 (N_13206,N_12765,N_12901);
xnor U13207 (N_13207,N_12887,N_12845);
and U13208 (N_13208,N_12837,N_12846);
and U13209 (N_13209,N_12943,N_12904);
and U13210 (N_13210,N_12863,N_12791);
or U13211 (N_13211,N_12954,N_12960);
and U13212 (N_13212,N_12987,N_12904);
nand U13213 (N_13213,N_12824,N_12808);
and U13214 (N_13214,N_12960,N_12820);
or U13215 (N_13215,N_12907,N_12943);
or U13216 (N_13216,N_12820,N_12759);
xnor U13217 (N_13217,N_12916,N_12768);
or U13218 (N_13218,N_12912,N_12784);
nand U13219 (N_13219,N_12956,N_12953);
or U13220 (N_13220,N_12875,N_12822);
nand U13221 (N_13221,N_12829,N_12974);
or U13222 (N_13222,N_12912,N_12805);
and U13223 (N_13223,N_12774,N_12784);
and U13224 (N_13224,N_12965,N_12781);
and U13225 (N_13225,N_12916,N_12813);
xnor U13226 (N_13226,N_12787,N_12838);
and U13227 (N_13227,N_12771,N_12911);
nor U13228 (N_13228,N_12883,N_12871);
nor U13229 (N_13229,N_12833,N_12940);
nand U13230 (N_13230,N_12897,N_12912);
nor U13231 (N_13231,N_12983,N_12848);
and U13232 (N_13232,N_12771,N_12822);
and U13233 (N_13233,N_12915,N_12836);
nand U13234 (N_13234,N_12758,N_12845);
or U13235 (N_13235,N_12798,N_12966);
nor U13236 (N_13236,N_12912,N_12774);
xnor U13237 (N_13237,N_12773,N_12756);
nor U13238 (N_13238,N_12975,N_12761);
nand U13239 (N_13239,N_12812,N_12852);
xnor U13240 (N_13240,N_12930,N_12960);
and U13241 (N_13241,N_12922,N_12924);
or U13242 (N_13242,N_12806,N_12765);
or U13243 (N_13243,N_12881,N_12984);
nor U13244 (N_13244,N_12899,N_12897);
nand U13245 (N_13245,N_12913,N_12849);
nand U13246 (N_13246,N_12889,N_12870);
xor U13247 (N_13247,N_12987,N_12788);
or U13248 (N_13248,N_12992,N_12852);
xnor U13249 (N_13249,N_12774,N_12879);
xor U13250 (N_13250,N_13189,N_13196);
and U13251 (N_13251,N_13129,N_13141);
nor U13252 (N_13252,N_13178,N_13206);
nor U13253 (N_13253,N_13158,N_13138);
and U13254 (N_13254,N_13050,N_13174);
or U13255 (N_13255,N_13053,N_13078);
nand U13256 (N_13256,N_13093,N_13097);
nor U13257 (N_13257,N_13222,N_13022);
and U13258 (N_13258,N_13167,N_13188);
or U13259 (N_13259,N_13100,N_13221);
nand U13260 (N_13260,N_13126,N_13139);
nand U13261 (N_13261,N_13003,N_13197);
nand U13262 (N_13262,N_13185,N_13166);
nor U13263 (N_13263,N_13068,N_13128);
and U13264 (N_13264,N_13148,N_13008);
nand U13265 (N_13265,N_13106,N_13157);
xnor U13266 (N_13266,N_13035,N_13028);
nand U13267 (N_13267,N_13079,N_13193);
and U13268 (N_13268,N_13095,N_13013);
nand U13269 (N_13269,N_13127,N_13020);
and U13270 (N_13270,N_13110,N_13219);
nand U13271 (N_13271,N_13200,N_13123);
or U13272 (N_13272,N_13143,N_13026);
and U13273 (N_13273,N_13137,N_13223);
xor U13274 (N_13274,N_13056,N_13208);
nand U13275 (N_13275,N_13060,N_13118);
xor U13276 (N_13276,N_13045,N_13172);
or U13277 (N_13277,N_13047,N_13227);
nand U13278 (N_13278,N_13096,N_13226);
nand U13279 (N_13279,N_13205,N_13165);
and U13280 (N_13280,N_13150,N_13229);
nor U13281 (N_13281,N_13145,N_13204);
or U13282 (N_13282,N_13051,N_13182);
xor U13283 (N_13283,N_13218,N_13052);
nand U13284 (N_13284,N_13001,N_13034);
nor U13285 (N_13285,N_13090,N_13194);
or U13286 (N_13286,N_13058,N_13023);
nor U13287 (N_13287,N_13173,N_13142);
or U13288 (N_13288,N_13103,N_13216);
nand U13289 (N_13289,N_13109,N_13120);
nand U13290 (N_13290,N_13072,N_13039);
or U13291 (N_13291,N_13246,N_13149);
and U13292 (N_13292,N_13215,N_13159);
xor U13293 (N_13293,N_13241,N_13240);
nand U13294 (N_13294,N_13006,N_13059);
or U13295 (N_13295,N_13073,N_13081);
and U13296 (N_13296,N_13048,N_13085);
xor U13297 (N_13297,N_13232,N_13029);
nand U13298 (N_13298,N_13074,N_13005);
or U13299 (N_13299,N_13086,N_13105);
and U13300 (N_13300,N_13065,N_13163);
or U13301 (N_13301,N_13214,N_13211);
xor U13302 (N_13302,N_13220,N_13024);
and U13303 (N_13303,N_13049,N_13224);
and U13304 (N_13304,N_13154,N_13146);
nand U13305 (N_13305,N_13071,N_13092);
nor U13306 (N_13306,N_13132,N_13153);
xnor U13307 (N_13307,N_13140,N_13108);
nor U13308 (N_13308,N_13187,N_13147);
xor U13309 (N_13309,N_13247,N_13169);
nor U13310 (N_13310,N_13201,N_13007);
nor U13311 (N_13311,N_13055,N_13033);
nand U13312 (N_13312,N_13066,N_13207);
or U13313 (N_13313,N_13113,N_13070);
or U13314 (N_13314,N_13155,N_13179);
and U13315 (N_13315,N_13116,N_13069);
nand U13316 (N_13316,N_13160,N_13195);
and U13317 (N_13317,N_13156,N_13236);
nor U13318 (N_13318,N_13015,N_13170);
nand U13319 (N_13319,N_13230,N_13042);
xor U13320 (N_13320,N_13122,N_13067);
or U13321 (N_13321,N_13115,N_13030);
and U13322 (N_13322,N_13191,N_13234);
and U13323 (N_13323,N_13002,N_13114);
nand U13324 (N_13324,N_13077,N_13184);
nor U13325 (N_13325,N_13019,N_13202);
and U13326 (N_13326,N_13025,N_13054);
nand U13327 (N_13327,N_13044,N_13121);
nor U13328 (N_13328,N_13018,N_13088);
nor U13329 (N_13329,N_13064,N_13027);
nor U13330 (N_13330,N_13124,N_13112);
nand U13331 (N_13331,N_13176,N_13038);
nor U13332 (N_13332,N_13014,N_13119);
or U13333 (N_13333,N_13076,N_13245);
nor U13334 (N_13334,N_13040,N_13011);
and U13335 (N_13335,N_13217,N_13228);
or U13336 (N_13336,N_13199,N_13243);
nand U13337 (N_13337,N_13057,N_13032);
and U13338 (N_13338,N_13102,N_13089);
and U13339 (N_13339,N_13000,N_13212);
or U13340 (N_13340,N_13171,N_13136);
or U13341 (N_13341,N_13061,N_13213);
xnor U13342 (N_13342,N_13152,N_13098);
nand U13343 (N_13343,N_13134,N_13233);
nor U13344 (N_13344,N_13101,N_13131);
nand U13345 (N_13345,N_13239,N_13012);
or U13346 (N_13346,N_13238,N_13180);
nor U13347 (N_13347,N_13164,N_13190);
nand U13348 (N_13348,N_13186,N_13209);
or U13349 (N_13349,N_13062,N_13111);
xnor U13350 (N_13350,N_13080,N_13183);
xor U13351 (N_13351,N_13162,N_13041);
nor U13352 (N_13352,N_13083,N_13135);
or U13353 (N_13353,N_13031,N_13231);
xor U13354 (N_13354,N_13168,N_13091);
and U13355 (N_13355,N_13017,N_13210);
nor U13356 (N_13356,N_13151,N_13242);
and U13357 (N_13357,N_13010,N_13094);
nand U13358 (N_13358,N_13046,N_13107);
nor U13359 (N_13359,N_13021,N_13104);
nand U13360 (N_13360,N_13225,N_13177);
or U13361 (N_13361,N_13235,N_13192);
or U13362 (N_13362,N_13036,N_13009);
xor U13363 (N_13363,N_13175,N_13117);
or U13364 (N_13364,N_13244,N_13016);
or U13365 (N_13365,N_13004,N_13130);
and U13366 (N_13366,N_13125,N_13198);
or U13367 (N_13367,N_13237,N_13248);
nor U13368 (N_13368,N_13181,N_13144);
xnor U13369 (N_13369,N_13084,N_13249);
and U13370 (N_13370,N_13087,N_13133);
and U13371 (N_13371,N_13037,N_13063);
or U13372 (N_13372,N_13082,N_13075);
and U13373 (N_13373,N_13043,N_13203);
nor U13374 (N_13374,N_13099,N_13161);
or U13375 (N_13375,N_13027,N_13044);
and U13376 (N_13376,N_13100,N_13033);
nand U13377 (N_13377,N_13133,N_13175);
and U13378 (N_13378,N_13123,N_13175);
and U13379 (N_13379,N_13192,N_13083);
xnor U13380 (N_13380,N_13112,N_13101);
nor U13381 (N_13381,N_13199,N_13007);
xnor U13382 (N_13382,N_13066,N_13076);
nand U13383 (N_13383,N_13143,N_13116);
xor U13384 (N_13384,N_13188,N_13138);
nor U13385 (N_13385,N_13187,N_13118);
and U13386 (N_13386,N_13025,N_13059);
xnor U13387 (N_13387,N_13151,N_13016);
nand U13388 (N_13388,N_13120,N_13072);
xor U13389 (N_13389,N_13172,N_13102);
xor U13390 (N_13390,N_13118,N_13055);
nand U13391 (N_13391,N_13052,N_13106);
nand U13392 (N_13392,N_13136,N_13134);
nor U13393 (N_13393,N_13164,N_13129);
or U13394 (N_13394,N_13122,N_13229);
and U13395 (N_13395,N_13123,N_13144);
nor U13396 (N_13396,N_13031,N_13220);
nand U13397 (N_13397,N_13046,N_13225);
nand U13398 (N_13398,N_13144,N_13104);
xor U13399 (N_13399,N_13245,N_13075);
and U13400 (N_13400,N_13081,N_13152);
xnor U13401 (N_13401,N_13240,N_13077);
nor U13402 (N_13402,N_13121,N_13002);
nor U13403 (N_13403,N_13071,N_13057);
xor U13404 (N_13404,N_13228,N_13241);
and U13405 (N_13405,N_13160,N_13232);
nand U13406 (N_13406,N_13109,N_13183);
or U13407 (N_13407,N_13024,N_13100);
xnor U13408 (N_13408,N_13021,N_13222);
nor U13409 (N_13409,N_13104,N_13156);
nor U13410 (N_13410,N_13245,N_13206);
xor U13411 (N_13411,N_13183,N_13018);
nand U13412 (N_13412,N_13128,N_13035);
xnor U13413 (N_13413,N_13071,N_13105);
or U13414 (N_13414,N_13049,N_13097);
and U13415 (N_13415,N_13137,N_13032);
nand U13416 (N_13416,N_13052,N_13246);
and U13417 (N_13417,N_13149,N_13103);
nor U13418 (N_13418,N_13001,N_13218);
nor U13419 (N_13419,N_13181,N_13090);
xnor U13420 (N_13420,N_13125,N_13051);
nand U13421 (N_13421,N_13131,N_13066);
nor U13422 (N_13422,N_13041,N_13118);
nand U13423 (N_13423,N_13097,N_13103);
or U13424 (N_13424,N_13173,N_13174);
nand U13425 (N_13425,N_13119,N_13095);
nand U13426 (N_13426,N_13004,N_13098);
nor U13427 (N_13427,N_13246,N_13201);
or U13428 (N_13428,N_13120,N_13235);
xor U13429 (N_13429,N_13012,N_13155);
nand U13430 (N_13430,N_13100,N_13076);
xnor U13431 (N_13431,N_13190,N_13192);
or U13432 (N_13432,N_13144,N_13113);
xor U13433 (N_13433,N_13019,N_13062);
and U13434 (N_13434,N_13042,N_13125);
nand U13435 (N_13435,N_13053,N_13032);
nand U13436 (N_13436,N_13169,N_13214);
xnor U13437 (N_13437,N_13025,N_13246);
xnor U13438 (N_13438,N_13163,N_13000);
and U13439 (N_13439,N_13095,N_13043);
nand U13440 (N_13440,N_13012,N_13032);
and U13441 (N_13441,N_13097,N_13039);
xnor U13442 (N_13442,N_13228,N_13188);
xor U13443 (N_13443,N_13040,N_13125);
or U13444 (N_13444,N_13125,N_13214);
or U13445 (N_13445,N_13151,N_13189);
and U13446 (N_13446,N_13201,N_13086);
nor U13447 (N_13447,N_13220,N_13027);
and U13448 (N_13448,N_13099,N_13196);
xor U13449 (N_13449,N_13075,N_13206);
xor U13450 (N_13450,N_13021,N_13142);
xnor U13451 (N_13451,N_13135,N_13108);
nor U13452 (N_13452,N_13029,N_13068);
nor U13453 (N_13453,N_13032,N_13028);
or U13454 (N_13454,N_13237,N_13135);
xor U13455 (N_13455,N_13075,N_13103);
nand U13456 (N_13456,N_13148,N_13087);
xnor U13457 (N_13457,N_13078,N_13114);
and U13458 (N_13458,N_13010,N_13235);
and U13459 (N_13459,N_13242,N_13097);
and U13460 (N_13460,N_13051,N_13248);
nand U13461 (N_13461,N_13008,N_13161);
and U13462 (N_13462,N_13130,N_13223);
or U13463 (N_13463,N_13194,N_13046);
and U13464 (N_13464,N_13248,N_13164);
and U13465 (N_13465,N_13130,N_13193);
or U13466 (N_13466,N_13154,N_13138);
and U13467 (N_13467,N_13024,N_13015);
nand U13468 (N_13468,N_13042,N_13188);
or U13469 (N_13469,N_13241,N_13039);
xnor U13470 (N_13470,N_13148,N_13159);
or U13471 (N_13471,N_13245,N_13190);
xnor U13472 (N_13472,N_13121,N_13231);
nand U13473 (N_13473,N_13124,N_13050);
nand U13474 (N_13474,N_13003,N_13202);
nand U13475 (N_13475,N_13006,N_13134);
nand U13476 (N_13476,N_13248,N_13076);
or U13477 (N_13477,N_13138,N_13239);
nand U13478 (N_13478,N_13047,N_13101);
xnor U13479 (N_13479,N_13229,N_13046);
xor U13480 (N_13480,N_13205,N_13045);
xor U13481 (N_13481,N_13163,N_13100);
nand U13482 (N_13482,N_13225,N_13202);
nand U13483 (N_13483,N_13105,N_13117);
xor U13484 (N_13484,N_13042,N_13195);
xnor U13485 (N_13485,N_13209,N_13191);
nor U13486 (N_13486,N_13096,N_13205);
xor U13487 (N_13487,N_13222,N_13059);
nor U13488 (N_13488,N_13228,N_13105);
and U13489 (N_13489,N_13158,N_13094);
nand U13490 (N_13490,N_13141,N_13143);
xor U13491 (N_13491,N_13043,N_13155);
and U13492 (N_13492,N_13029,N_13120);
and U13493 (N_13493,N_13247,N_13024);
or U13494 (N_13494,N_13060,N_13200);
and U13495 (N_13495,N_13242,N_13073);
and U13496 (N_13496,N_13213,N_13234);
or U13497 (N_13497,N_13022,N_13211);
xor U13498 (N_13498,N_13063,N_13000);
and U13499 (N_13499,N_13124,N_13141);
nor U13500 (N_13500,N_13494,N_13497);
nand U13501 (N_13501,N_13458,N_13434);
or U13502 (N_13502,N_13369,N_13456);
or U13503 (N_13503,N_13328,N_13417);
or U13504 (N_13504,N_13489,N_13325);
or U13505 (N_13505,N_13476,N_13277);
xnor U13506 (N_13506,N_13350,N_13463);
nand U13507 (N_13507,N_13484,N_13250);
xnor U13508 (N_13508,N_13345,N_13421);
or U13509 (N_13509,N_13354,N_13390);
and U13510 (N_13510,N_13260,N_13399);
nand U13511 (N_13511,N_13286,N_13379);
or U13512 (N_13512,N_13441,N_13486);
xnor U13513 (N_13513,N_13452,N_13424);
nand U13514 (N_13514,N_13437,N_13372);
or U13515 (N_13515,N_13464,N_13301);
xnor U13516 (N_13516,N_13343,N_13349);
nor U13517 (N_13517,N_13447,N_13380);
xnor U13518 (N_13518,N_13377,N_13366);
and U13519 (N_13519,N_13363,N_13318);
xor U13520 (N_13520,N_13423,N_13392);
xnor U13521 (N_13521,N_13308,N_13493);
nand U13522 (N_13522,N_13468,N_13481);
or U13523 (N_13523,N_13382,N_13305);
xnor U13524 (N_13524,N_13393,N_13474);
or U13525 (N_13525,N_13367,N_13443);
xnor U13526 (N_13526,N_13465,N_13322);
nand U13527 (N_13527,N_13394,N_13347);
and U13528 (N_13528,N_13331,N_13285);
and U13529 (N_13529,N_13267,N_13341);
and U13530 (N_13530,N_13386,N_13428);
or U13531 (N_13531,N_13405,N_13453);
nand U13532 (N_13532,N_13413,N_13270);
nor U13533 (N_13533,N_13398,N_13488);
and U13534 (N_13534,N_13491,N_13256);
and U13535 (N_13535,N_13302,N_13287);
and U13536 (N_13536,N_13268,N_13336);
and U13537 (N_13537,N_13492,N_13264);
nand U13538 (N_13538,N_13385,N_13445);
and U13539 (N_13539,N_13338,N_13314);
nand U13540 (N_13540,N_13439,N_13454);
nand U13541 (N_13541,N_13293,N_13298);
nor U13542 (N_13542,N_13255,N_13451);
xor U13543 (N_13543,N_13383,N_13358);
xnor U13544 (N_13544,N_13310,N_13438);
xnor U13545 (N_13545,N_13353,N_13412);
and U13546 (N_13546,N_13401,N_13351);
nor U13547 (N_13547,N_13499,N_13478);
nand U13548 (N_13548,N_13324,N_13356);
or U13549 (N_13549,N_13272,N_13329);
or U13550 (N_13550,N_13279,N_13311);
nand U13551 (N_13551,N_13435,N_13446);
and U13552 (N_13552,N_13389,N_13275);
and U13553 (N_13553,N_13337,N_13333);
nor U13554 (N_13554,N_13496,N_13265);
nor U13555 (N_13555,N_13289,N_13375);
xnor U13556 (N_13556,N_13259,N_13258);
and U13557 (N_13557,N_13257,N_13334);
and U13558 (N_13558,N_13371,N_13422);
nor U13559 (N_13559,N_13319,N_13365);
and U13560 (N_13560,N_13364,N_13404);
or U13561 (N_13561,N_13291,N_13274);
xnor U13562 (N_13562,N_13425,N_13388);
and U13563 (N_13563,N_13473,N_13309);
and U13564 (N_13564,N_13469,N_13471);
or U13565 (N_13565,N_13427,N_13420);
nand U13566 (N_13566,N_13307,N_13407);
xnor U13567 (N_13567,N_13470,N_13408);
xnor U13568 (N_13568,N_13397,N_13282);
nand U13569 (N_13569,N_13327,N_13455);
and U13570 (N_13570,N_13283,N_13460);
and U13571 (N_13571,N_13339,N_13321);
nand U13572 (N_13572,N_13475,N_13376);
and U13573 (N_13573,N_13391,N_13374);
xnor U13574 (N_13574,N_13482,N_13406);
nor U13575 (N_13575,N_13303,N_13403);
or U13576 (N_13576,N_13490,N_13450);
nor U13577 (N_13577,N_13409,N_13348);
nor U13578 (N_13578,N_13462,N_13429);
or U13579 (N_13579,N_13487,N_13295);
or U13580 (N_13580,N_13416,N_13485);
or U13581 (N_13581,N_13432,N_13359);
xnor U13582 (N_13582,N_13332,N_13352);
or U13583 (N_13583,N_13430,N_13269);
or U13584 (N_13584,N_13251,N_13355);
xor U13585 (N_13585,N_13433,N_13395);
xnor U13586 (N_13586,N_13368,N_13297);
nand U13587 (N_13587,N_13396,N_13400);
nor U13588 (N_13588,N_13461,N_13480);
nand U13589 (N_13589,N_13402,N_13317);
nand U13590 (N_13590,N_13418,N_13320);
and U13591 (N_13591,N_13357,N_13483);
nand U13592 (N_13592,N_13323,N_13262);
nand U13593 (N_13593,N_13381,N_13414);
nor U13594 (N_13594,N_13294,N_13457);
nor U13595 (N_13595,N_13362,N_13316);
nor U13596 (N_13596,N_13479,N_13360);
or U13597 (N_13597,N_13370,N_13276);
or U13598 (N_13598,N_13290,N_13495);
nand U13599 (N_13599,N_13300,N_13448);
or U13600 (N_13600,N_13384,N_13281);
xnor U13601 (N_13601,N_13296,N_13436);
and U13602 (N_13602,N_13387,N_13415);
nand U13603 (N_13603,N_13335,N_13340);
or U13604 (N_13604,N_13472,N_13344);
or U13605 (N_13605,N_13449,N_13253);
nor U13606 (N_13606,N_13342,N_13410);
or U13607 (N_13607,N_13466,N_13271);
and U13608 (N_13608,N_13266,N_13498);
nand U13609 (N_13609,N_13288,N_13263);
nor U13610 (N_13610,N_13330,N_13346);
or U13611 (N_13611,N_13440,N_13459);
xor U13612 (N_13612,N_13312,N_13254);
and U13613 (N_13613,N_13306,N_13299);
nand U13614 (N_13614,N_13292,N_13431);
or U13615 (N_13615,N_13426,N_13326);
or U13616 (N_13616,N_13252,N_13411);
xor U13617 (N_13617,N_13467,N_13304);
and U13618 (N_13618,N_13444,N_13313);
or U13619 (N_13619,N_13378,N_13361);
nand U13620 (N_13620,N_13280,N_13273);
and U13621 (N_13621,N_13261,N_13373);
or U13622 (N_13622,N_13419,N_13442);
and U13623 (N_13623,N_13315,N_13477);
xnor U13624 (N_13624,N_13278,N_13284);
nor U13625 (N_13625,N_13321,N_13450);
or U13626 (N_13626,N_13444,N_13426);
nor U13627 (N_13627,N_13306,N_13342);
or U13628 (N_13628,N_13370,N_13268);
nand U13629 (N_13629,N_13420,N_13440);
or U13630 (N_13630,N_13342,N_13385);
or U13631 (N_13631,N_13376,N_13412);
nand U13632 (N_13632,N_13269,N_13378);
xnor U13633 (N_13633,N_13325,N_13411);
nor U13634 (N_13634,N_13413,N_13488);
xnor U13635 (N_13635,N_13456,N_13457);
or U13636 (N_13636,N_13278,N_13362);
nor U13637 (N_13637,N_13422,N_13383);
or U13638 (N_13638,N_13311,N_13375);
xnor U13639 (N_13639,N_13266,N_13336);
and U13640 (N_13640,N_13357,N_13331);
nand U13641 (N_13641,N_13434,N_13492);
nand U13642 (N_13642,N_13258,N_13394);
nor U13643 (N_13643,N_13455,N_13437);
nand U13644 (N_13644,N_13263,N_13321);
nor U13645 (N_13645,N_13417,N_13286);
or U13646 (N_13646,N_13418,N_13413);
or U13647 (N_13647,N_13300,N_13307);
or U13648 (N_13648,N_13438,N_13376);
or U13649 (N_13649,N_13450,N_13312);
xor U13650 (N_13650,N_13397,N_13298);
xor U13651 (N_13651,N_13349,N_13371);
and U13652 (N_13652,N_13465,N_13469);
and U13653 (N_13653,N_13251,N_13336);
and U13654 (N_13654,N_13294,N_13409);
nor U13655 (N_13655,N_13369,N_13404);
and U13656 (N_13656,N_13386,N_13323);
and U13657 (N_13657,N_13431,N_13399);
and U13658 (N_13658,N_13434,N_13381);
xor U13659 (N_13659,N_13349,N_13269);
or U13660 (N_13660,N_13435,N_13418);
nor U13661 (N_13661,N_13382,N_13285);
nor U13662 (N_13662,N_13299,N_13386);
or U13663 (N_13663,N_13464,N_13413);
nand U13664 (N_13664,N_13426,N_13427);
xor U13665 (N_13665,N_13329,N_13260);
nand U13666 (N_13666,N_13450,N_13368);
and U13667 (N_13667,N_13396,N_13478);
or U13668 (N_13668,N_13396,N_13348);
xnor U13669 (N_13669,N_13467,N_13479);
nor U13670 (N_13670,N_13357,N_13272);
nor U13671 (N_13671,N_13323,N_13397);
or U13672 (N_13672,N_13350,N_13410);
nand U13673 (N_13673,N_13297,N_13425);
xor U13674 (N_13674,N_13428,N_13392);
xor U13675 (N_13675,N_13410,N_13351);
nand U13676 (N_13676,N_13360,N_13283);
xor U13677 (N_13677,N_13411,N_13296);
or U13678 (N_13678,N_13363,N_13438);
and U13679 (N_13679,N_13496,N_13315);
and U13680 (N_13680,N_13250,N_13427);
and U13681 (N_13681,N_13334,N_13349);
or U13682 (N_13682,N_13406,N_13330);
nor U13683 (N_13683,N_13343,N_13263);
and U13684 (N_13684,N_13379,N_13499);
or U13685 (N_13685,N_13433,N_13461);
nand U13686 (N_13686,N_13439,N_13451);
nor U13687 (N_13687,N_13466,N_13474);
nor U13688 (N_13688,N_13458,N_13382);
and U13689 (N_13689,N_13401,N_13444);
xnor U13690 (N_13690,N_13433,N_13335);
nand U13691 (N_13691,N_13393,N_13305);
nand U13692 (N_13692,N_13351,N_13417);
xor U13693 (N_13693,N_13494,N_13428);
or U13694 (N_13694,N_13387,N_13385);
and U13695 (N_13695,N_13335,N_13272);
nand U13696 (N_13696,N_13488,N_13496);
or U13697 (N_13697,N_13411,N_13287);
and U13698 (N_13698,N_13360,N_13393);
and U13699 (N_13699,N_13390,N_13343);
nand U13700 (N_13700,N_13473,N_13448);
xnor U13701 (N_13701,N_13255,N_13267);
and U13702 (N_13702,N_13447,N_13436);
nor U13703 (N_13703,N_13334,N_13475);
nand U13704 (N_13704,N_13292,N_13428);
or U13705 (N_13705,N_13254,N_13331);
nand U13706 (N_13706,N_13368,N_13497);
nand U13707 (N_13707,N_13313,N_13383);
or U13708 (N_13708,N_13402,N_13426);
nor U13709 (N_13709,N_13415,N_13368);
nor U13710 (N_13710,N_13291,N_13423);
nand U13711 (N_13711,N_13285,N_13339);
nor U13712 (N_13712,N_13379,N_13437);
nand U13713 (N_13713,N_13442,N_13345);
nor U13714 (N_13714,N_13371,N_13330);
nand U13715 (N_13715,N_13309,N_13358);
and U13716 (N_13716,N_13396,N_13456);
or U13717 (N_13717,N_13392,N_13461);
and U13718 (N_13718,N_13466,N_13471);
nor U13719 (N_13719,N_13416,N_13423);
nand U13720 (N_13720,N_13265,N_13279);
nand U13721 (N_13721,N_13493,N_13312);
and U13722 (N_13722,N_13395,N_13473);
nand U13723 (N_13723,N_13316,N_13341);
nor U13724 (N_13724,N_13478,N_13334);
or U13725 (N_13725,N_13383,N_13328);
nor U13726 (N_13726,N_13351,N_13262);
xor U13727 (N_13727,N_13428,N_13264);
nor U13728 (N_13728,N_13414,N_13446);
nor U13729 (N_13729,N_13368,N_13401);
and U13730 (N_13730,N_13294,N_13273);
nor U13731 (N_13731,N_13381,N_13324);
xnor U13732 (N_13732,N_13318,N_13466);
or U13733 (N_13733,N_13276,N_13491);
nor U13734 (N_13734,N_13317,N_13447);
nand U13735 (N_13735,N_13450,N_13343);
nand U13736 (N_13736,N_13490,N_13477);
nand U13737 (N_13737,N_13379,N_13303);
nand U13738 (N_13738,N_13456,N_13357);
and U13739 (N_13739,N_13368,N_13327);
nand U13740 (N_13740,N_13424,N_13371);
nand U13741 (N_13741,N_13438,N_13275);
and U13742 (N_13742,N_13490,N_13364);
and U13743 (N_13743,N_13342,N_13257);
xnor U13744 (N_13744,N_13415,N_13450);
or U13745 (N_13745,N_13404,N_13465);
nand U13746 (N_13746,N_13305,N_13335);
and U13747 (N_13747,N_13490,N_13488);
and U13748 (N_13748,N_13334,N_13499);
nor U13749 (N_13749,N_13295,N_13428);
and U13750 (N_13750,N_13570,N_13719);
xnor U13751 (N_13751,N_13546,N_13671);
nor U13752 (N_13752,N_13645,N_13640);
and U13753 (N_13753,N_13643,N_13634);
xnor U13754 (N_13754,N_13705,N_13617);
or U13755 (N_13755,N_13748,N_13597);
xor U13756 (N_13756,N_13609,N_13598);
xnor U13757 (N_13757,N_13696,N_13667);
and U13758 (N_13758,N_13620,N_13538);
nand U13759 (N_13759,N_13527,N_13685);
nand U13760 (N_13760,N_13644,N_13679);
nor U13761 (N_13761,N_13575,N_13724);
xnor U13762 (N_13762,N_13602,N_13511);
xnor U13763 (N_13763,N_13506,N_13518);
or U13764 (N_13764,N_13654,N_13545);
xor U13765 (N_13765,N_13700,N_13703);
nor U13766 (N_13766,N_13557,N_13614);
nor U13767 (N_13767,N_13727,N_13728);
nor U13768 (N_13768,N_13539,N_13621);
xnor U13769 (N_13769,N_13655,N_13601);
or U13770 (N_13770,N_13528,N_13682);
nand U13771 (N_13771,N_13571,N_13653);
nand U13772 (N_13772,N_13738,N_13593);
or U13773 (N_13773,N_13549,N_13576);
or U13774 (N_13774,N_13604,N_13581);
and U13775 (N_13775,N_13695,N_13592);
nor U13776 (N_13776,N_13661,N_13600);
or U13777 (N_13777,N_13739,N_13648);
or U13778 (N_13778,N_13716,N_13521);
and U13779 (N_13779,N_13512,N_13606);
or U13780 (N_13780,N_13559,N_13713);
and U13781 (N_13781,N_13689,N_13708);
xnor U13782 (N_13782,N_13647,N_13674);
nand U13783 (N_13783,N_13572,N_13569);
xnor U13784 (N_13784,N_13721,N_13717);
nor U13785 (N_13785,N_13567,N_13725);
or U13786 (N_13786,N_13637,N_13737);
xnor U13787 (N_13787,N_13730,N_13585);
nand U13788 (N_13788,N_13745,N_13690);
and U13789 (N_13789,N_13564,N_13664);
nand U13790 (N_13790,N_13522,N_13687);
and U13791 (N_13791,N_13710,N_13513);
nor U13792 (N_13792,N_13666,N_13623);
or U13793 (N_13793,N_13507,N_13698);
or U13794 (N_13794,N_13616,N_13638);
nand U13795 (N_13795,N_13534,N_13560);
and U13796 (N_13796,N_13732,N_13612);
xor U13797 (N_13797,N_13520,N_13694);
nor U13798 (N_13798,N_13706,N_13740);
nand U13799 (N_13799,N_13625,N_13624);
and U13800 (N_13800,N_13529,N_13747);
nand U13801 (N_13801,N_13544,N_13741);
nand U13802 (N_13802,N_13524,N_13591);
nand U13803 (N_13803,N_13680,N_13726);
nor U13804 (N_13804,N_13526,N_13548);
nand U13805 (N_13805,N_13532,N_13607);
xnor U13806 (N_13806,N_13583,N_13712);
xnor U13807 (N_13807,N_13537,N_13714);
and U13808 (N_13808,N_13540,N_13589);
and U13809 (N_13809,N_13588,N_13563);
nor U13810 (N_13810,N_13519,N_13514);
xnor U13811 (N_13811,N_13641,N_13650);
or U13812 (N_13812,N_13672,N_13579);
or U13813 (N_13813,N_13630,N_13709);
or U13814 (N_13814,N_13743,N_13733);
and U13815 (N_13815,N_13556,N_13692);
and U13816 (N_13816,N_13547,N_13504);
nand U13817 (N_13817,N_13673,N_13586);
and U13818 (N_13818,N_13686,N_13702);
or U13819 (N_13819,N_13558,N_13584);
and U13820 (N_13820,N_13678,N_13676);
or U13821 (N_13821,N_13566,N_13693);
or U13822 (N_13822,N_13632,N_13608);
nand U13823 (N_13823,N_13541,N_13722);
or U13824 (N_13824,N_13502,N_13701);
and U13825 (N_13825,N_13711,N_13599);
xnor U13826 (N_13826,N_13622,N_13552);
and U13827 (N_13827,N_13699,N_13587);
nand U13828 (N_13828,N_13642,N_13508);
or U13829 (N_13829,N_13651,N_13729);
or U13830 (N_13830,N_13627,N_13530);
nor U13831 (N_13831,N_13568,N_13668);
nand U13832 (N_13832,N_13731,N_13691);
and U13833 (N_13833,N_13742,N_13619);
xor U13834 (N_13834,N_13633,N_13574);
xnor U13835 (N_13835,N_13670,N_13578);
or U13836 (N_13836,N_13531,N_13697);
nand U13837 (N_13837,N_13683,N_13649);
nand U13838 (N_13838,N_13631,N_13720);
nor U13839 (N_13839,N_13523,N_13626);
nor U13840 (N_13840,N_13618,N_13543);
or U13841 (N_13841,N_13516,N_13659);
and U13842 (N_13842,N_13510,N_13596);
nor U13843 (N_13843,N_13515,N_13613);
xnor U13844 (N_13844,N_13553,N_13707);
nand U13845 (N_13845,N_13603,N_13542);
nor U13846 (N_13846,N_13665,N_13715);
nor U13847 (N_13847,N_13565,N_13669);
nor U13848 (N_13848,N_13501,N_13503);
and U13849 (N_13849,N_13749,N_13554);
xnor U13850 (N_13850,N_13517,N_13681);
or U13851 (N_13851,N_13580,N_13594);
xnor U13852 (N_13852,N_13615,N_13636);
or U13853 (N_13853,N_13646,N_13652);
xnor U13854 (N_13854,N_13595,N_13657);
xnor U13855 (N_13855,N_13723,N_13639);
xnor U13856 (N_13856,N_13629,N_13663);
nor U13857 (N_13857,N_13677,N_13684);
nor U13858 (N_13858,N_13628,N_13505);
or U13859 (N_13859,N_13675,N_13525);
nand U13860 (N_13860,N_13734,N_13658);
nor U13861 (N_13861,N_13562,N_13551);
xnor U13862 (N_13862,N_13573,N_13536);
and U13863 (N_13863,N_13688,N_13535);
nand U13864 (N_13864,N_13635,N_13555);
xor U13865 (N_13865,N_13582,N_13735);
xor U13866 (N_13866,N_13718,N_13500);
nand U13867 (N_13867,N_13509,N_13605);
nor U13868 (N_13868,N_13610,N_13533);
nor U13869 (N_13869,N_13561,N_13611);
and U13870 (N_13870,N_13660,N_13656);
or U13871 (N_13871,N_13590,N_13550);
nand U13872 (N_13872,N_13577,N_13746);
xor U13873 (N_13873,N_13744,N_13662);
or U13874 (N_13874,N_13704,N_13736);
and U13875 (N_13875,N_13610,N_13683);
xnor U13876 (N_13876,N_13647,N_13537);
nor U13877 (N_13877,N_13672,N_13680);
xor U13878 (N_13878,N_13529,N_13626);
or U13879 (N_13879,N_13720,N_13505);
xor U13880 (N_13880,N_13550,N_13733);
or U13881 (N_13881,N_13575,N_13598);
nor U13882 (N_13882,N_13510,N_13682);
or U13883 (N_13883,N_13689,N_13637);
xor U13884 (N_13884,N_13504,N_13659);
or U13885 (N_13885,N_13721,N_13654);
xor U13886 (N_13886,N_13534,N_13578);
nand U13887 (N_13887,N_13664,N_13675);
nand U13888 (N_13888,N_13518,N_13743);
and U13889 (N_13889,N_13661,N_13696);
nor U13890 (N_13890,N_13729,N_13692);
nand U13891 (N_13891,N_13713,N_13642);
nor U13892 (N_13892,N_13565,N_13549);
and U13893 (N_13893,N_13654,N_13685);
nor U13894 (N_13894,N_13748,N_13665);
nor U13895 (N_13895,N_13644,N_13640);
nor U13896 (N_13896,N_13748,N_13625);
nor U13897 (N_13897,N_13633,N_13609);
nand U13898 (N_13898,N_13629,N_13711);
nor U13899 (N_13899,N_13653,N_13548);
xnor U13900 (N_13900,N_13543,N_13515);
nor U13901 (N_13901,N_13564,N_13596);
or U13902 (N_13902,N_13582,N_13572);
nor U13903 (N_13903,N_13702,N_13701);
or U13904 (N_13904,N_13720,N_13549);
nand U13905 (N_13905,N_13522,N_13717);
or U13906 (N_13906,N_13505,N_13506);
or U13907 (N_13907,N_13671,N_13639);
nor U13908 (N_13908,N_13700,N_13533);
or U13909 (N_13909,N_13531,N_13677);
nor U13910 (N_13910,N_13583,N_13717);
and U13911 (N_13911,N_13545,N_13542);
or U13912 (N_13912,N_13550,N_13518);
and U13913 (N_13913,N_13690,N_13695);
nand U13914 (N_13914,N_13649,N_13625);
nand U13915 (N_13915,N_13648,N_13662);
nand U13916 (N_13916,N_13674,N_13566);
nor U13917 (N_13917,N_13718,N_13742);
xnor U13918 (N_13918,N_13555,N_13539);
nand U13919 (N_13919,N_13533,N_13628);
and U13920 (N_13920,N_13626,N_13692);
or U13921 (N_13921,N_13723,N_13695);
and U13922 (N_13922,N_13659,N_13707);
nand U13923 (N_13923,N_13746,N_13539);
nand U13924 (N_13924,N_13624,N_13686);
xnor U13925 (N_13925,N_13609,N_13503);
or U13926 (N_13926,N_13629,N_13548);
xnor U13927 (N_13927,N_13550,N_13633);
xor U13928 (N_13928,N_13748,N_13553);
or U13929 (N_13929,N_13662,N_13696);
xor U13930 (N_13930,N_13722,N_13564);
and U13931 (N_13931,N_13642,N_13559);
nand U13932 (N_13932,N_13631,N_13703);
xor U13933 (N_13933,N_13569,N_13544);
nand U13934 (N_13934,N_13562,N_13731);
and U13935 (N_13935,N_13545,N_13551);
nand U13936 (N_13936,N_13739,N_13634);
and U13937 (N_13937,N_13659,N_13588);
and U13938 (N_13938,N_13604,N_13608);
and U13939 (N_13939,N_13744,N_13658);
xor U13940 (N_13940,N_13638,N_13736);
nand U13941 (N_13941,N_13701,N_13588);
or U13942 (N_13942,N_13717,N_13640);
or U13943 (N_13943,N_13545,N_13679);
or U13944 (N_13944,N_13547,N_13597);
or U13945 (N_13945,N_13606,N_13609);
xor U13946 (N_13946,N_13503,N_13699);
or U13947 (N_13947,N_13553,N_13520);
or U13948 (N_13948,N_13561,N_13575);
or U13949 (N_13949,N_13675,N_13719);
xor U13950 (N_13950,N_13506,N_13746);
nand U13951 (N_13951,N_13556,N_13652);
nor U13952 (N_13952,N_13575,N_13701);
or U13953 (N_13953,N_13737,N_13630);
xor U13954 (N_13954,N_13642,N_13663);
and U13955 (N_13955,N_13625,N_13568);
and U13956 (N_13956,N_13604,N_13622);
nand U13957 (N_13957,N_13581,N_13672);
nand U13958 (N_13958,N_13604,N_13621);
nor U13959 (N_13959,N_13724,N_13640);
nand U13960 (N_13960,N_13640,N_13744);
xnor U13961 (N_13961,N_13626,N_13694);
nor U13962 (N_13962,N_13665,N_13652);
nor U13963 (N_13963,N_13634,N_13699);
nand U13964 (N_13964,N_13539,N_13670);
or U13965 (N_13965,N_13513,N_13544);
and U13966 (N_13966,N_13674,N_13554);
nor U13967 (N_13967,N_13663,N_13728);
nand U13968 (N_13968,N_13616,N_13740);
nor U13969 (N_13969,N_13720,N_13565);
or U13970 (N_13970,N_13703,N_13736);
nor U13971 (N_13971,N_13501,N_13695);
xor U13972 (N_13972,N_13588,N_13501);
or U13973 (N_13973,N_13719,N_13689);
nand U13974 (N_13974,N_13536,N_13593);
or U13975 (N_13975,N_13748,N_13536);
xor U13976 (N_13976,N_13535,N_13596);
and U13977 (N_13977,N_13548,N_13705);
nand U13978 (N_13978,N_13580,N_13648);
nor U13979 (N_13979,N_13719,N_13730);
or U13980 (N_13980,N_13602,N_13681);
nand U13981 (N_13981,N_13566,N_13585);
nor U13982 (N_13982,N_13625,N_13653);
nor U13983 (N_13983,N_13605,N_13610);
nand U13984 (N_13984,N_13633,N_13638);
xnor U13985 (N_13985,N_13723,N_13609);
nor U13986 (N_13986,N_13560,N_13551);
or U13987 (N_13987,N_13657,N_13510);
or U13988 (N_13988,N_13539,N_13509);
or U13989 (N_13989,N_13701,N_13599);
nor U13990 (N_13990,N_13537,N_13696);
or U13991 (N_13991,N_13703,N_13656);
nor U13992 (N_13992,N_13726,N_13569);
and U13993 (N_13993,N_13565,N_13687);
or U13994 (N_13994,N_13529,N_13526);
and U13995 (N_13995,N_13657,N_13515);
nor U13996 (N_13996,N_13735,N_13741);
xor U13997 (N_13997,N_13620,N_13512);
and U13998 (N_13998,N_13662,N_13572);
or U13999 (N_13999,N_13532,N_13570);
xnor U14000 (N_14000,N_13943,N_13754);
nand U14001 (N_14001,N_13818,N_13970);
nand U14002 (N_14002,N_13867,N_13775);
and U14003 (N_14003,N_13777,N_13962);
nand U14004 (N_14004,N_13892,N_13833);
and U14005 (N_14005,N_13879,N_13787);
xnor U14006 (N_14006,N_13770,N_13919);
nand U14007 (N_14007,N_13819,N_13788);
nor U14008 (N_14008,N_13825,N_13903);
nor U14009 (N_14009,N_13843,N_13849);
nor U14010 (N_14010,N_13969,N_13928);
nor U14011 (N_14011,N_13858,N_13865);
nor U14012 (N_14012,N_13804,N_13923);
nand U14013 (N_14013,N_13757,N_13976);
nor U14014 (N_14014,N_13841,N_13792);
and U14015 (N_14015,N_13940,N_13875);
or U14016 (N_14016,N_13878,N_13881);
nand U14017 (N_14017,N_13988,N_13912);
nand U14018 (N_14018,N_13887,N_13896);
and U14019 (N_14019,N_13760,N_13750);
nand U14020 (N_14020,N_13989,N_13860);
xnor U14021 (N_14021,N_13963,N_13938);
nand U14022 (N_14022,N_13836,N_13955);
nand U14023 (N_14023,N_13886,N_13926);
nand U14024 (N_14024,N_13781,N_13924);
nor U14025 (N_14025,N_13772,N_13764);
or U14026 (N_14026,N_13813,N_13851);
or U14027 (N_14027,N_13884,N_13801);
xor U14028 (N_14028,N_13946,N_13857);
and U14029 (N_14029,N_13800,N_13987);
and U14030 (N_14030,N_13965,N_13799);
xor U14031 (N_14031,N_13806,N_13871);
and U14032 (N_14032,N_13952,N_13933);
nand U14033 (N_14033,N_13961,N_13791);
and U14034 (N_14034,N_13828,N_13809);
nor U14035 (N_14035,N_13883,N_13755);
nor U14036 (N_14036,N_13866,N_13902);
xor U14037 (N_14037,N_13907,N_13789);
and U14038 (N_14038,N_13921,N_13844);
and U14039 (N_14039,N_13774,N_13894);
nor U14040 (N_14040,N_13798,N_13889);
nand U14041 (N_14041,N_13964,N_13888);
xnor U14042 (N_14042,N_13909,N_13853);
or U14043 (N_14043,N_13936,N_13977);
or U14044 (N_14044,N_13765,N_13766);
or U14045 (N_14045,N_13854,N_13868);
or U14046 (N_14046,N_13758,N_13763);
nand U14047 (N_14047,N_13939,N_13824);
or U14048 (N_14048,N_13802,N_13945);
or U14049 (N_14049,N_13949,N_13999);
xnor U14050 (N_14050,N_13918,N_13914);
or U14051 (N_14051,N_13816,N_13899);
or U14052 (N_14052,N_13931,N_13932);
nor U14053 (N_14053,N_13779,N_13823);
and U14054 (N_14054,N_13773,N_13930);
nor U14055 (N_14055,N_13862,N_13771);
nor U14056 (N_14056,N_13897,N_13807);
xor U14057 (N_14057,N_13994,N_13956);
and U14058 (N_14058,N_13925,N_13855);
nor U14059 (N_14059,N_13793,N_13797);
or U14060 (N_14060,N_13873,N_13937);
and U14061 (N_14061,N_13780,N_13861);
or U14062 (N_14062,N_13847,N_13966);
nand U14063 (N_14063,N_13984,N_13814);
nor U14064 (N_14064,N_13882,N_13845);
or U14065 (N_14065,N_13834,N_13954);
xor U14066 (N_14066,N_13794,N_13796);
nand U14067 (N_14067,N_13944,N_13803);
nor U14068 (N_14068,N_13974,N_13986);
or U14069 (N_14069,N_13998,N_13869);
and U14070 (N_14070,N_13885,N_13927);
and U14071 (N_14071,N_13790,N_13784);
nand U14072 (N_14072,N_13753,N_13953);
xor U14073 (N_14073,N_13810,N_13817);
nor U14074 (N_14074,N_13990,N_13975);
nor U14075 (N_14075,N_13795,N_13769);
xnor U14076 (N_14076,N_13959,N_13996);
and U14077 (N_14077,N_13951,N_13876);
and U14078 (N_14078,N_13972,N_13831);
and U14079 (N_14079,N_13830,N_13820);
nor U14080 (N_14080,N_13915,N_13905);
xnor U14081 (N_14081,N_13852,N_13859);
and U14082 (N_14082,N_13985,N_13827);
nor U14083 (N_14083,N_13992,N_13895);
nand U14084 (N_14084,N_13783,N_13826);
nor U14085 (N_14085,N_13993,N_13929);
or U14086 (N_14086,N_13908,N_13948);
or U14087 (N_14087,N_13916,N_13968);
and U14088 (N_14088,N_13767,N_13822);
xor U14089 (N_14089,N_13756,N_13950);
nand U14090 (N_14090,N_13761,N_13759);
and U14091 (N_14091,N_13898,N_13979);
or U14092 (N_14092,N_13837,N_13960);
and U14093 (N_14093,N_13967,N_13983);
xnor U14094 (N_14094,N_13846,N_13971);
or U14095 (N_14095,N_13782,N_13811);
and U14096 (N_14096,N_13864,N_13880);
nand U14097 (N_14097,N_13752,N_13982);
or U14098 (N_14098,N_13911,N_13874);
nand U14099 (N_14099,N_13848,N_13850);
or U14100 (N_14100,N_13973,N_13821);
nor U14101 (N_14101,N_13786,N_13840);
and U14102 (N_14102,N_13877,N_13978);
nand U14103 (N_14103,N_13906,N_13995);
nor U14104 (N_14104,N_13776,N_13890);
xnor U14105 (N_14105,N_13941,N_13839);
and U14106 (N_14106,N_13957,N_13778);
or U14107 (N_14107,N_13997,N_13942);
nor U14108 (N_14108,N_13891,N_13805);
and U14109 (N_14109,N_13901,N_13751);
or U14110 (N_14110,N_13863,N_13785);
and U14111 (N_14111,N_13842,N_13913);
or U14112 (N_14112,N_13893,N_13991);
xor U14113 (N_14113,N_13958,N_13768);
and U14114 (N_14114,N_13980,N_13838);
and U14115 (N_14115,N_13947,N_13904);
and U14116 (N_14116,N_13900,N_13832);
and U14117 (N_14117,N_13922,N_13910);
and U14118 (N_14118,N_13762,N_13935);
and U14119 (N_14119,N_13808,N_13872);
or U14120 (N_14120,N_13812,N_13920);
nand U14121 (N_14121,N_13981,N_13870);
nand U14122 (N_14122,N_13835,N_13815);
xor U14123 (N_14123,N_13917,N_13829);
xnor U14124 (N_14124,N_13934,N_13856);
nor U14125 (N_14125,N_13838,N_13916);
nand U14126 (N_14126,N_13758,N_13994);
or U14127 (N_14127,N_13895,N_13828);
xnor U14128 (N_14128,N_13843,N_13947);
nor U14129 (N_14129,N_13804,N_13881);
and U14130 (N_14130,N_13837,N_13831);
nand U14131 (N_14131,N_13818,N_13796);
nor U14132 (N_14132,N_13831,N_13841);
or U14133 (N_14133,N_13793,N_13822);
xor U14134 (N_14134,N_13970,N_13761);
and U14135 (N_14135,N_13815,N_13877);
or U14136 (N_14136,N_13801,N_13800);
nand U14137 (N_14137,N_13856,N_13976);
xnor U14138 (N_14138,N_13930,N_13986);
nand U14139 (N_14139,N_13801,N_13973);
or U14140 (N_14140,N_13880,N_13961);
nand U14141 (N_14141,N_13890,N_13786);
nand U14142 (N_14142,N_13959,N_13968);
nand U14143 (N_14143,N_13938,N_13951);
xnor U14144 (N_14144,N_13802,N_13946);
nor U14145 (N_14145,N_13832,N_13944);
and U14146 (N_14146,N_13815,N_13889);
or U14147 (N_14147,N_13786,N_13762);
nor U14148 (N_14148,N_13861,N_13860);
nor U14149 (N_14149,N_13843,N_13834);
and U14150 (N_14150,N_13973,N_13778);
nand U14151 (N_14151,N_13920,N_13852);
xor U14152 (N_14152,N_13950,N_13936);
xnor U14153 (N_14153,N_13870,N_13777);
and U14154 (N_14154,N_13855,N_13987);
nor U14155 (N_14155,N_13793,N_13896);
nor U14156 (N_14156,N_13925,N_13757);
or U14157 (N_14157,N_13949,N_13871);
xor U14158 (N_14158,N_13928,N_13789);
and U14159 (N_14159,N_13782,N_13958);
or U14160 (N_14160,N_13851,N_13953);
nor U14161 (N_14161,N_13834,N_13784);
or U14162 (N_14162,N_13785,N_13828);
nand U14163 (N_14163,N_13869,N_13953);
or U14164 (N_14164,N_13845,N_13911);
nand U14165 (N_14165,N_13776,N_13992);
or U14166 (N_14166,N_13757,N_13960);
or U14167 (N_14167,N_13936,N_13988);
nor U14168 (N_14168,N_13886,N_13935);
nand U14169 (N_14169,N_13869,N_13858);
and U14170 (N_14170,N_13929,N_13981);
nor U14171 (N_14171,N_13923,N_13864);
and U14172 (N_14172,N_13843,N_13794);
nor U14173 (N_14173,N_13972,N_13806);
xor U14174 (N_14174,N_13787,N_13987);
nor U14175 (N_14175,N_13751,N_13848);
nand U14176 (N_14176,N_13998,N_13884);
or U14177 (N_14177,N_13783,N_13876);
nand U14178 (N_14178,N_13922,N_13864);
and U14179 (N_14179,N_13774,N_13856);
and U14180 (N_14180,N_13881,N_13832);
and U14181 (N_14181,N_13832,N_13986);
or U14182 (N_14182,N_13842,N_13771);
nand U14183 (N_14183,N_13900,N_13848);
and U14184 (N_14184,N_13991,N_13827);
nand U14185 (N_14185,N_13865,N_13767);
nor U14186 (N_14186,N_13794,N_13940);
nor U14187 (N_14187,N_13812,N_13948);
or U14188 (N_14188,N_13805,N_13799);
and U14189 (N_14189,N_13983,N_13779);
nand U14190 (N_14190,N_13841,N_13883);
xor U14191 (N_14191,N_13949,N_13830);
nor U14192 (N_14192,N_13928,N_13982);
nor U14193 (N_14193,N_13808,N_13834);
nor U14194 (N_14194,N_13813,N_13995);
nor U14195 (N_14195,N_13926,N_13896);
nand U14196 (N_14196,N_13772,N_13955);
xnor U14197 (N_14197,N_13933,N_13973);
nor U14198 (N_14198,N_13868,N_13761);
nor U14199 (N_14199,N_13799,N_13969);
xnor U14200 (N_14200,N_13919,N_13873);
or U14201 (N_14201,N_13824,N_13943);
xor U14202 (N_14202,N_13903,N_13842);
xor U14203 (N_14203,N_13995,N_13994);
nor U14204 (N_14204,N_13914,N_13876);
or U14205 (N_14205,N_13786,N_13969);
or U14206 (N_14206,N_13874,N_13869);
and U14207 (N_14207,N_13886,N_13862);
and U14208 (N_14208,N_13981,N_13799);
or U14209 (N_14209,N_13921,N_13915);
and U14210 (N_14210,N_13793,N_13791);
nand U14211 (N_14211,N_13989,N_13770);
or U14212 (N_14212,N_13854,N_13760);
nand U14213 (N_14213,N_13970,N_13834);
nor U14214 (N_14214,N_13851,N_13753);
xnor U14215 (N_14215,N_13951,N_13829);
xor U14216 (N_14216,N_13851,N_13932);
or U14217 (N_14217,N_13880,N_13898);
xnor U14218 (N_14218,N_13885,N_13953);
nor U14219 (N_14219,N_13758,N_13808);
xnor U14220 (N_14220,N_13832,N_13827);
and U14221 (N_14221,N_13809,N_13918);
nand U14222 (N_14222,N_13909,N_13896);
nand U14223 (N_14223,N_13846,N_13985);
xor U14224 (N_14224,N_13925,N_13960);
or U14225 (N_14225,N_13891,N_13905);
and U14226 (N_14226,N_13919,N_13965);
nor U14227 (N_14227,N_13885,N_13978);
and U14228 (N_14228,N_13955,N_13831);
nand U14229 (N_14229,N_13862,N_13825);
or U14230 (N_14230,N_13845,N_13765);
xor U14231 (N_14231,N_13890,N_13884);
or U14232 (N_14232,N_13916,N_13766);
nand U14233 (N_14233,N_13905,N_13844);
nor U14234 (N_14234,N_13947,N_13869);
xnor U14235 (N_14235,N_13878,N_13816);
xnor U14236 (N_14236,N_13781,N_13826);
or U14237 (N_14237,N_13816,N_13757);
xnor U14238 (N_14238,N_13931,N_13942);
and U14239 (N_14239,N_13892,N_13819);
or U14240 (N_14240,N_13877,N_13819);
xor U14241 (N_14241,N_13961,N_13985);
or U14242 (N_14242,N_13755,N_13911);
xnor U14243 (N_14243,N_13808,N_13979);
xor U14244 (N_14244,N_13869,N_13770);
nor U14245 (N_14245,N_13839,N_13929);
xnor U14246 (N_14246,N_13887,N_13979);
nand U14247 (N_14247,N_13921,N_13940);
xor U14248 (N_14248,N_13924,N_13926);
xor U14249 (N_14249,N_13936,N_13829);
or U14250 (N_14250,N_14052,N_14010);
and U14251 (N_14251,N_14215,N_14129);
and U14252 (N_14252,N_14040,N_14139);
nand U14253 (N_14253,N_14117,N_14028);
nand U14254 (N_14254,N_14152,N_14091);
xnor U14255 (N_14255,N_14160,N_14008);
xor U14256 (N_14256,N_14184,N_14187);
or U14257 (N_14257,N_14212,N_14179);
xnor U14258 (N_14258,N_14136,N_14083);
nand U14259 (N_14259,N_14197,N_14232);
nor U14260 (N_14260,N_14190,N_14219);
or U14261 (N_14261,N_14023,N_14033);
and U14262 (N_14262,N_14162,N_14013);
nor U14263 (N_14263,N_14027,N_14110);
nor U14264 (N_14264,N_14082,N_14238);
and U14265 (N_14265,N_14119,N_14004);
xnor U14266 (N_14266,N_14249,N_14089);
or U14267 (N_14267,N_14041,N_14196);
or U14268 (N_14268,N_14120,N_14243);
nor U14269 (N_14269,N_14032,N_14167);
nor U14270 (N_14270,N_14049,N_14072);
or U14271 (N_14271,N_14054,N_14224);
nand U14272 (N_14272,N_14065,N_14170);
xor U14273 (N_14273,N_14235,N_14036);
xor U14274 (N_14274,N_14019,N_14007);
and U14275 (N_14275,N_14189,N_14199);
nand U14276 (N_14276,N_14188,N_14201);
nand U14277 (N_14277,N_14029,N_14166);
xor U14278 (N_14278,N_14230,N_14221);
nand U14279 (N_14279,N_14090,N_14217);
and U14280 (N_14280,N_14131,N_14046);
and U14281 (N_14281,N_14073,N_14148);
nand U14282 (N_14282,N_14157,N_14181);
nor U14283 (N_14283,N_14210,N_14233);
and U14284 (N_14284,N_14079,N_14084);
and U14285 (N_14285,N_14015,N_14241);
nor U14286 (N_14286,N_14114,N_14132);
or U14287 (N_14287,N_14056,N_14014);
nor U14288 (N_14288,N_14077,N_14005);
nand U14289 (N_14289,N_14145,N_14048);
and U14290 (N_14290,N_14126,N_14016);
or U14291 (N_14291,N_14047,N_14209);
or U14292 (N_14292,N_14053,N_14246);
or U14293 (N_14293,N_14081,N_14130);
or U14294 (N_14294,N_14149,N_14022);
and U14295 (N_14295,N_14085,N_14123);
xnor U14296 (N_14296,N_14024,N_14144);
and U14297 (N_14297,N_14070,N_14099);
nand U14298 (N_14298,N_14218,N_14000);
and U14299 (N_14299,N_14227,N_14002);
xor U14300 (N_14300,N_14192,N_14026);
xnor U14301 (N_14301,N_14071,N_14208);
nor U14302 (N_14302,N_14109,N_14037);
and U14303 (N_14303,N_14133,N_14092);
and U14304 (N_14304,N_14205,N_14061);
xnor U14305 (N_14305,N_14097,N_14102);
xor U14306 (N_14306,N_14135,N_14220);
nand U14307 (N_14307,N_14186,N_14175);
xor U14308 (N_14308,N_14150,N_14017);
xor U14309 (N_14309,N_14159,N_14161);
xnor U14310 (N_14310,N_14011,N_14153);
nand U14311 (N_14311,N_14035,N_14247);
and U14312 (N_14312,N_14095,N_14154);
and U14313 (N_14313,N_14057,N_14198);
nor U14314 (N_14314,N_14080,N_14087);
or U14315 (N_14315,N_14178,N_14088);
nand U14316 (N_14316,N_14234,N_14100);
and U14317 (N_14317,N_14121,N_14169);
xnor U14318 (N_14318,N_14060,N_14158);
nor U14319 (N_14319,N_14108,N_14141);
xnor U14320 (N_14320,N_14193,N_14031);
and U14321 (N_14321,N_14043,N_14059);
xnor U14322 (N_14322,N_14113,N_14006);
xnor U14323 (N_14323,N_14122,N_14143);
and U14324 (N_14324,N_14094,N_14231);
xnor U14325 (N_14325,N_14245,N_14018);
nor U14326 (N_14326,N_14030,N_14244);
and U14327 (N_14327,N_14134,N_14111);
nand U14328 (N_14328,N_14138,N_14204);
nor U14329 (N_14329,N_14177,N_14021);
nand U14330 (N_14330,N_14012,N_14118);
xnor U14331 (N_14331,N_14051,N_14239);
xor U14332 (N_14332,N_14171,N_14174);
nor U14333 (N_14333,N_14214,N_14237);
and U14334 (N_14334,N_14104,N_14063);
xor U14335 (N_14335,N_14001,N_14207);
and U14336 (N_14336,N_14137,N_14222);
nand U14337 (N_14337,N_14206,N_14128);
xnor U14338 (N_14338,N_14168,N_14062);
xor U14339 (N_14339,N_14112,N_14156);
xnor U14340 (N_14340,N_14172,N_14069);
and U14341 (N_14341,N_14101,N_14213);
nand U14342 (N_14342,N_14045,N_14078);
nand U14343 (N_14343,N_14116,N_14140);
and U14344 (N_14344,N_14066,N_14106);
nor U14345 (N_14345,N_14038,N_14127);
and U14346 (N_14346,N_14125,N_14067);
xnor U14347 (N_14347,N_14034,N_14086);
xnor U14348 (N_14348,N_14185,N_14211);
xnor U14349 (N_14349,N_14203,N_14009);
nand U14350 (N_14350,N_14236,N_14075);
xor U14351 (N_14351,N_14225,N_14248);
or U14352 (N_14352,N_14173,N_14093);
or U14353 (N_14353,N_14068,N_14003);
and U14354 (N_14354,N_14076,N_14200);
xor U14355 (N_14355,N_14107,N_14142);
or U14356 (N_14356,N_14025,N_14105);
nor U14357 (N_14357,N_14151,N_14042);
nand U14358 (N_14358,N_14146,N_14229);
and U14359 (N_14359,N_14180,N_14228);
nand U14360 (N_14360,N_14242,N_14020);
nor U14361 (N_14361,N_14165,N_14124);
and U14362 (N_14362,N_14055,N_14098);
nor U14363 (N_14363,N_14039,N_14195);
and U14364 (N_14364,N_14163,N_14223);
or U14365 (N_14365,N_14182,N_14064);
xnor U14366 (N_14366,N_14183,N_14240);
and U14367 (N_14367,N_14226,N_14176);
nand U14368 (N_14368,N_14044,N_14115);
and U14369 (N_14369,N_14164,N_14058);
or U14370 (N_14370,N_14147,N_14096);
or U14371 (N_14371,N_14074,N_14103);
and U14372 (N_14372,N_14050,N_14155);
xor U14373 (N_14373,N_14202,N_14194);
nor U14374 (N_14374,N_14191,N_14216);
nand U14375 (N_14375,N_14093,N_14062);
and U14376 (N_14376,N_14041,N_14145);
nor U14377 (N_14377,N_14233,N_14172);
xnor U14378 (N_14378,N_14242,N_14015);
and U14379 (N_14379,N_14041,N_14048);
xnor U14380 (N_14380,N_14155,N_14148);
or U14381 (N_14381,N_14009,N_14062);
xor U14382 (N_14382,N_14012,N_14203);
and U14383 (N_14383,N_14070,N_14041);
xor U14384 (N_14384,N_14128,N_14088);
xor U14385 (N_14385,N_14109,N_14194);
nor U14386 (N_14386,N_14005,N_14148);
xor U14387 (N_14387,N_14166,N_14176);
xor U14388 (N_14388,N_14105,N_14150);
xnor U14389 (N_14389,N_14190,N_14160);
nor U14390 (N_14390,N_14138,N_14128);
nand U14391 (N_14391,N_14125,N_14224);
or U14392 (N_14392,N_14248,N_14228);
or U14393 (N_14393,N_14239,N_14120);
nor U14394 (N_14394,N_14103,N_14210);
xnor U14395 (N_14395,N_14104,N_14013);
nand U14396 (N_14396,N_14042,N_14075);
nand U14397 (N_14397,N_14173,N_14161);
xnor U14398 (N_14398,N_14239,N_14127);
nand U14399 (N_14399,N_14040,N_14126);
xor U14400 (N_14400,N_14021,N_14110);
nand U14401 (N_14401,N_14186,N_14193);
and U14402 (N_14402,N_14183,N_14037);
and U14403 (N_14403,N_14130,N_14145);
nand U14404 (N_14404,N_14245,N_14086);
nor U14405 (N_14405,N_14066,N_14246);
and U14406 (N_14406,N_14211,N_14051);
and U14407 (N_14407,N_14132,N_14202);
nor U14408 (N_14408,N_14174,N_14038);
and U14409 (N_14409,N_14233,N_14221);
nor U14410 (N_14410,N_14016,N_14048);
xnor U14411 (N_14411,N_14088,N_14202);
xor U14412 (N_14412,N_14103,N_14090);
xor U14413 (N_14413,N_14148,N_14196);
xor U14414 (N_14414,N_14187,N_14007);
and U14415 (N_14415,N_14191,N_14097);
nand U14416 (N_14416,N_14102,N_14014);
xnor U14417 (N_14417,N_14081,N_14144);
nand U14418 (N_14418,N_14225,N_14024);
nand U14419 (N_14419,N_14094,N_14097);
xor U14420 (N_14420,N_14180,N_14240);
nor U14421 (N_14421,N_14192,N_14040);
xor U14422 (N_14422,N_14165,N_14182);
and U14423 (N_14423,N_14100,N_14070);
or U14424 (N_14424,N_14242,N_14007);
xor U14425 (N_14425,N_14103,N_14022);
nor U14426 (N_14426,N_14164,N_14240);
nor U14427 (N_14427,N_14137,N_14027);
xor U14428 (N_14428,N_14055,N_14074);
nand U14429 (N_14429,N_14029,N_14165);
nand U14430 (N_14430,N_14208,N_14137);
nand U14431 (N_14431,N_14086,N_14121);
or U14432 (N_14432,N_14244,N_14164);
and U14433 (N_14433,N_14226,N_14200);
nor U14434 (N_14434,N_14239,N_14219);
and U14435 (N_14435,N_14207,N_14053);
and U14436 (N_14436,N_14095,N_14177);
nand U14437 (N_14437,N_14213,N_14161);
and U14438 (N_14438,N_14073,N_14162);
or U14439 (N_14439,N_14159,N_14186);
nand U14440 (N_14440,N_14077,N_14030);
and U14441 (N_14441,N_14113,N_14119);
xnor U14442 (N_14442,N_14001,N_14049);
or U14443 (N_14443,N_14184,N_14241);
nor U14444 (N_14444,N_14004,N_14058);
or U14445 (N_14445,N_14229,N_14069);
or U14446 (N_14446,N_14081,N_14120);
xnor U14447 (N_14447,N_14089,N_14191);
and U14448 (N_14448,N_14160,N_14156);
and U14449 (N_14449,N_14045,N_14231);
nor U14450 (N_14450,N_14028,N_14061);
or U14451 (N_14451,N_14081,N_14221);
and U14452 (N_14452,N_14108,N_14013);
or U14453 (N_14453,N_14126,N_14195);
or U14454 (N_14454,N_14248,N_14150);
xor U14455 (N_14455,N_14207,N_14045);
xnor U14456 (N_14456,N_14011,N_14152);
nand U14457 (N_14457,N_14243,N_14136);
and U14458 (N_14458,N_14023,N_14042);
xnor U14459 (N_14459,N_14187,N_14074);
nand U14460 (N_14460,N_14226,N_14011);
xor U14461 (N_14461,N_14047,N_14092);
and U14462 (N_14462,N_14062,N_14040);
xor U14463 (N_14463,N_14113,N_14103);
xor U14464 (N_14464,N_14169,N_14219);
nand U14465 (N_14465,N_14197,N_14241);
nand U14466 (N_14466,N_14042,N_14205);
and U14467 (N_14467,N_14009,N_14139);
nand U14468 (N_14468,N_14170,N_14123);
and U14469 (N_14469,N_14101,N_14210);
or U14470 (N_14470,N_14147,N_14193);
and U14471 (N_14471,N_14241,N_14081);
xnor U14472 (N_14472,N_14132,N_14065);
and U14473 (N_14473,N_14008,N_14061);
nand U14474 (N_14474,N_14107,N_14006);
nand U14475 (N_14475,N_14098,N_14089);
and U14476 (N_14476,N_14157,N_14119);
nor U14477 (N_14477,N_14116,N_14236);
xor U14478 (N_14478,N_14094,N_14224);
or U14479 (N_14479,N_14145,N_14095);
nand U14480 (N_14480,N_14094,N_14055);
and U14481 (N_14481,N_14160,N_14080);
nand U14482 (N_14482,N_14091,N_14221);
and U14483 (N_14483,N_14040,N_14140);
nor U14484 (N_14484,N_14229,N_14105);
xnor U14485 (N_14485,N_14036,N_14108);
xor U14486 (N_14486,N_14116,N_14232);
and U14487 (N_14487,N_14194,N_14117);
xor U14488 (N_14488,N_14003,N_14145);
or U14489 (N_14489,N_14125,N_14066);
and U14490 (N_14490,N_14161,N_14210);
nor U14491 (N_14491,N_14137,N_14033);
or U14492 (N_14492,N_14096,N_14226);
or U14493 (N_14493,N_14132,N_14156);
and U14494 (N_14494,N_14055,N_14222);
nand U14495 (N_14495,N_14033,N_14234);
nor U14496 (N_14496,N_14203,N_14208);
and U14497 (N_14497,N_14088,N_14061);
and U14498 (N_14498,N_14214,N_14100);
nand U14499 (N_14499,N_14022,N_14151);
or U14500 (N_14500,N_14348,N_14277);
xor U14501 (N_14501,N_14414,N_14413);
nand U14502 (N_14502,N_14266,N_14465);
and U14503 (N_14503,N_14343,N_14316);
and U14504 (N_14504,N_14353,N_14363);
nand U14505 (N_14505,N_14416,N_14284);
nand U14506 (N_14506,N_14302,N_14368);
nand U14507 (N_14507,N_14419,N_14483);
and U14508 (N_14508,N_14379,N_14369);
nor U14509 (N_14509,N_14443,N_14390);
xnor U14510 (N_14510,N_14377,N_14338);
xor U14511 (N_14511,N_14301,N_14344);
xnor U14512 (N_14512,N_14321,N_14396);
and U14513 (N_14513,N_14424,N_14380);
nand U14514 (N_14514,N_14273,N_14275);
nand U14515 (N_14515,N_14432,N_14361);
xor U14516 (N_14516,N_14337,N_14411);
xnor U14517 (N_14517,N_14331,N_14327);
nor U14518 (N_14518,N_14429,N_14373);
and U14519 (N_14519,N_14255,N_14287);
nor U14520 (N_14520,N_14263,N_14288);
or U14521 (N_14521,N_14276,N_14487);
or U14522 (N_14522,N_14322,N_14422);
xor U14523 (N_14523,N_14289,N_14365);
nand U14524 (N_14524,N_14375,N_14260);
xnor U14525 (N_14525,N_14445,N_14378);
nand U14526 (N_14526,N_14472,N_14261);
and U14527 (N_14527,N_14488,N_14490);
and U14528 (N_14528,N_14399,N_14460);
or U14529 (N_14529,N_14258,N_14270);
nor U14530 (N_14530,N_14433,N_14421);
or U14531 (N_14531,N_14383,N_14423);
and U14532 (N_14532,N_14281,N_14484);
and U14533 (N_14533,N_14468,N_14317);
nand U14534 (N_14534,N_14446,N_14403);
xnor U14535 (N_14535,N_14364,N_14444);
nor U14536 (N_14536,N_14431,N_14496);
xor U14537 (N_14537,N_14485,N_14351);
nand U14538 (N_14538,N_14350,N_14451);
and U14539 (N_14539,N_14358,N_14340);
nand U14540 (N_14540,N_14459,N_14291);
and U14541 (N_14541,N_14372,N_14308);
xnor U14542 (N_14542,N_14286,N_14309);
and U14543 (N_14543,N_14320,N_14314);
or U14544 (N_14544,N_14311,N_14262);
and U14545 (N_14545,N_14486,N_14250);
nor U14546 (N_14546,N_14466,N_14251);
and U14547 (N_14547,N_14271,N_14285);
nand U14548 (N_14548,N_14300,N_14257);
xor U14549 (N_14549,N_14417,N_14282);
xnor U14550 (N_14550,N_14254,N_14323);
and U14551 (N_14551,N_14400,N_14296);
nand U14552 (N_14552,N_14315,N_14440);
and U14553 (N_14553,N_14415,N_14319);
and U14554 (N_14554,N_14359,N_14434);
nor U14555 (N_14555,N_14402,N_14435);
nor U14556 (N_14556,N_14325,N_14332);
or U14557 (N_14557,N_14387,N_14494);
xor U14558 (N_14558,N_14283,N_14326);
xor U14559 (N_14559,N_14398,N_14329);
or U14560 (N_14560,N_14475,N_14253);
nand U14561 (N_14561,N_14409,N_14401);
nor U14562 (N_14562,N_14265,N_14430);
nand U14563 (N_14563,N_14476,N_14469);
or U14564 (N_14564,N_14450,N_14303);
or U14565 (N_14565,N_14385,N_14473);
nor U14566 (N_14566,N_14374,N_14341);
nor U14567 (N_14567,N_14493,N_14252);
nor U14568 (N_14568,N_14464,N_14355);
and U14569 (N_14569,N_14313,N_14357);
and U14570 (N_14570,N_14376,N_14439);
nor U14571 (N_14571,N_14356,N_14442);
and U14572 (N_14572,N_14274,N_14453);
or U14573 (N_14573,N_14426,N_14334);
xnor U14574 (N_14574,N_14272,N_14418);
nor U14575 (N_14575,N_14345,N_14437);
or U14576 (N_14576,N_14389,N_14498);
xor U14577 (N_14577,N_14386,N_14461);
and U14578 (N_14578,N_14290,N_14481);
nand U14579 (N_14579,N_14447,N_14256);
nor U14580 (N_14580,N_14349,N_14278);
nand U14581 (N_14581,N_14299,N_14427);
and U14582 (N_14582,N_14408,N_14449);
xnor U14583 (N_14583,N_14489,N_14480);
and U14584 (N_14584,N_14497,N_14463);
nor U14585 (N_14585,N_14477,N_14333);
or U14586 (N_14586,N_14479,N_14335);
nand U14587 (N_14587,N_14292,N_14412);
nand U14588 (N_14588,N_14499,N_14259);
nand U14589 (N_14589,N_14293,N_14474);
nand U14590 (N_14590,N_14354,N_14407);
nand U14591 (N_14591,N_14482,N_14267);
xnor U14592 (N_14592,N_14393,N_14307);
xor U14593 (N_14593,N_14280,N_14467);
nor U14594 (N_14594,N_14388,N_14428);
or U14595 (N_14595,N_14382,N_14397);
and U14596 (N_14596,N_14452,N_14371);
xor U14597 (N_14597,N_14346,N_14384);
or U14598 (N_14598,N_14438,N_14352);
xnor U14599 (N_14599,N_14366,N_14310);
nor U14600 (N_14600,N_14436,N_14471);
xor U14601 (N_14601,N_14441,N_14339);
nor U14602 (N_14602,N_14448,N_14425);
xnor U14603 (N_14603,N_14297,N_14454);
nor U14604 (N_14604,N_14347,N_14362);
or U14605 (N_14605,N_14470,N_14395);
or U14606 (N_14606,N_14391,N_14462);
or U14607 (N_14607,N_14298,N_14328);
and U14608 (N_14608,N_14294,N_14360);
xor U14609 (N_14609,N_14457,N_14330);
or U14610 (N_14610,N_14405,N_14478);
or U14611 (N_14611,N_14370,N_14342);
and U14612 (N_14612,N_14410,N_14264);
nand U14613 (N_14613,N_14406,N_14394);
nor U14614 (N_14614,N_14456,N_14312);
xnor U14615 (N_14615,N_14336,N_14324);
nand U14616 (N_14616,N_14295,N_14492);
nand U14617 (N_14617,N_14268,N_14381);
nand U14618 (N_14618,N_14306,N_14404);
nand U14619 (N_14619,N_14279,N_14392);
nand U14620 (N_14620,N_14458,N_14269);
xor U14621 (N_14621,N_14420,N_14367);
or U14622 (N_14622,N_14304,N_14305);
and U14623 (N_14623,N_14318,N_14495);
xor U14624 (N_14624,N_14491,N_14455);
and U14625 (N_14625,N_14399,N_14301);
and U14626 (N_14626,N_14381,N_14343);
xor U14627 (N_14627,N_14354,N_14323);
and U14628 (N_14628,N_14399,N_14461);
and U14629 (N_14629,N_14294,N_14372);
or U14630 (N_14630,N_14463,N_14329);
or U14631 (N_14631,N_14301,N_14412);
xnor U14632 (N_14632,N_14348,N_14325);
xor U14633 (N_14633,N_14498,N_14312);
nand U14634 (N_14634,N_14414,N_14279);
and U14635 (N_14635,N_14437,N_14406);
nand U14636 (N_14636,N_14263,N_14254);
nand U14637 (N_14637,N_14343,N_14442);
and U14638 (N_14638,N_14350,N_14347);
or U14639 (N_14639,N_14430,N_14424);
xor U14640 (N_14640,N_14259,N_14377);
nor U14641 (N_14641,N_14435,N_14420);
nand U14642 (N_14642,N_14320,N_14330);
nor U14643 (N_14643,N_14285,N_14436);
and U14644 (N_14644,N_14397,N_14366);
xor U14645 (N_14645,N_14372,N_14410);
xor U14646 (N_14646,N_14383,N_14292);
nand U14647 (N_14647,N_14368,N_14441);
or U14648 (N_14648,N_14267,N_14476);
xnor U14649 (N_14649,N_14383,N_14348);
nand U14650 (N_14650,N_14399,N_14300);
and U14651 (N_14651,N_14404,N_14304);
or U14652 (N_14652,N_14421,N_14344);
or U14653 (N_14653,N_14412,N_14424);
xnor U14654 (N_14654,N_14376,N_14359);
nor U14655 (N_14655,N_14276,N_14259);
or U14656 (N_14656,N_14431,N_14264);
or U14657 (N_14657,N_14463,N_14479);
nor U14658 (N_14658,N_14328,N_14251);
nand U14659 (N_14659,N_14300,N_14329);
xnor U14660 (N_14660,N_14347,N_14295);
xor U14661 (N_14661,N_14480,N_14371);
or U14662 (N_14662,N_14465,N_14392);
and U14663 (N_14663,N_14434,N_14406);
or U14664 (N_14664,N_14300,N_14417);
xnor U14665 (N_14665,N_14458,N_14444);
nor U14666 (N_14666,N_14377,N_14405);
and U14667 (N_14667,N_14477,N_14250);
xnor U14668 (N_14668,N_14331,N_14387);
or U14669 (N_14669,N_14445,N_14460);
nand U14670 (N_14670,N_14423,N_14374);
nor U14671 (N_14671,N_14370,N_14412);
nand U14672 (N_14672,N_14481,N_14321);
xor U14673 (N_14673,N_14446,N_14389);
nand U14674 (N_14674,N_14312,N_14372);
nor U14675 (N_14675,N_14399,N_14490);
nand U14676 (N_14676,N_14466,N_14437);
xor U14677 (N_14677,N_14390,N_14308);
nand U14678 (N_14678,N_14356,N_14381);
and U14679 (N_14679,N_14426,N_14441);
nor U14680 (N_14680,N_14362,N_14281);
or U14681 (N_14681,N_14341,N_14377);
and U14682 (N_14682,N_14430,N_14275);
nor U14683 (N_14683,N_14407,N_14265);
nand U14684 (N_14684,N_14316,N_14441);
and U14685 (N_14685,N_14324,N_14299);
nand U14686 (N_14686,N_14461,N_14490);
or U14687 (N_14687,N_14476,N_14338);
nand U14688 (N_14688,N_14269,N_14444);
nand U14689 (N_14689,N_14354,N_14350);
or U14690 (N_14690,N_14361,N_14333);
nand U14691 (N_14691,N_14473,N_14410);
nor U14692 (N_14692,N_14430,N_14493);
xor U14693 (N_14693,N_14391,N_14299);
or U14694 (N_14694,N_14427,N_14281);
nor U14695 (N_14695,N_14316,N_14295);
or U14696 (N_14696,N_14316,N_14465);
and U14697 (N_14697,N_14435,N_14401);
nor U14698 (N_14698,N_14433,N_14410);
and U14699 (N_14699,N_14456,N_14486);
nand U14700 (N_14700,N_14349,N_14467);
and U14701 (N_14701,N_14364,N_14366);
nand U14702 (N_14702,N_14318,N_14370);
nand U14703 (N_14703,N_14342,N_14413);
or U14704 (N_14704,N_14410,N_14366);
or U14705 (N_14705,N_14441,N_14375);
nand U14706 (N_14706,N_14490,N_14275);
and U14707 (N_14707,N_14331,N_14438);
and U14708 (N_14708,N_14307,N_14408);
nor U14709 (N_14709,N_14373,N_14316);
xnor U14710 (N_14710,N_14374,N_14425);
and U14711 (N_14711,N_14393,N_14296);
or U14712 (N_14712,N_14307,N_14481);
and U14713 (N_14713,N_14261,N_14372);
nor U14714 (N_14714,N_14393,N_14415);
nor U14715 (N_14715,N_14360,N_14285);
nor U14716 (N_14716,N_14471,N_14326);
xor U14717 (N_14717,N_14318,N_14298);
and U14718 (N_14718,N_14302,N_14306);
xor U14719 (N_14719,N_14345,N_14369);
nor U14720 (N_14720,N_14253,N_14415);
xor U14721 (N_14721,N_14277,N_14315);
nor U14722 (N_14722,N_14430,N_14411);
nor U14723 (N_14723,N_14492,N_14434);
nor U14724 (N_14724,N_14298,N_14375);
nand U14725 (N_14725,N_14397,N_14300);
and U14726 (N_14726,N_14256,N_14325);
xor U14727 (N_14727,N_14467,N_14363);
xor U14728 (N_14728,N_14478,N_14386);
and U14729 (N_14729,N_14250,N_14399);
xnor U14730 (N_14730,N_14455,N_14351);
and U14731 (N_14731,N_14390,N_14464);
and U14732 (N_14732,N_14428,N_14411);
xnor U14733 (N_14733,N_14469,N_14474);
nor U14734 (N_14734,N_14309,N_14395);
or U14735 (N_14735,N_14359,N_14328);
nor U14736 (N_14736,N_14375,N_14412);
xor U14737 (N_14737,N_14429,N_14299);
nor U14738 (N_14738,N_14452,N_14489);
nor U14739 (N_14739,N_14397,N_14257);
nor U14740 (N_14740,N_14390,N_14340);
nor U14741 (N_14741,N_14341,N_14434);
xnor U14742 (N_14742,N_14431,N_14471);
nand U14743 (N_14743,N_14253,N_14382);
xor U14744 (N_14744,N_14298,N_14396);
xor U14745 (N_14745,N_14449,N_14387);
xnor U14746 (N_14746,N_14332,N_14324);
nand U14747 (N_14747,N_14321,N_14266);
and U14748 (N_14748,N_14410,N_14280);
xnor U14749 (N_14749,N_14326,N_14426);
nor U14750 (N_14750,N_14593,N_14633);
xor U14751 (N_14751,N_14641,N_14588);
xnor U14752 (N_14752,N_14627,N_14708);
or U14753 (N_14753,N_14591,N_14605);
nor U14754 (N_14754,N_14562,N_14642);
xnor U14755 (N_14755,N_14589,N_14602);
and U14756 (N_14756,N_14636,N_14696);
nor U14757 (N_14757,N_14668,N_14505);
xor U14758 (N_14758,N_14608,N_14666);
and U14759 (N_14759,N_14689,N_14516);
nand U14760 (N_14760,N_14542,N_14652);
and U14761 (N_14761,N_14582,N_14682);
and U14762 (N_14762,N_14670,N_14727);
nand U14763 (N_14763,N_14713,N_14526);
or U14764 (N_14764,N_14658,N_14730);
xor U14765 (N_14765,N_14663,N_14744);
or U14766 (N_14766,N_14679,N_14547);
nor U14767 (N_14767,N_14502,N_14732);
nand U14768 (N_14768,N_14687,N_14628);
nor U14769 (N_14769,N_14657,N_14619);
xnor U14770 (N_14770,N_14699,N_14692);
xnor U14771 (N_14771,N_14726,N_14714);
nor U14772 (N_14772,N_14700,N_14717);
and U14773 (N_14773,N_14614,N_14573);
nor U14774 (N_14774,N_14749,N_14731);
and U14775 (N_14775,N_14674,N_14695);
nand U14776 (N_14776,N_14584,N_14541);
xor U14777 (N_14777,N_14643,N_14523);
and U14778 (N_14778,N_14688,N_14506);
nor U14779 (N_14779,N_14578,N_14653);
nor U14780 (N_14780,N_14722,N_14595);
and U14781 (N_14781,N_14551,N_14651);
and U14782 (N_14782,N_14583,N_14500);
nor U14783 (N_14783,N_14672,N_14587);
nor U14784 (N_14784,N_14634,N_14533);
xor U14785 (N_14785,N_14626,N_14590);
nand U14786 (N_14786,N_14720,N_14599);
nor U14787 (N_14787,N_14579,N_14550);
or U14788 (N_14788,N_14527,N_14733);
or U14789 (N_14789,N_14686,N_14662);
or U14790 (N_14790,N_14685,N_14552);
or U14791 (N_14791,N_14534,N_14748);
or U14792 (N_14792,N_14567,N_14565);
nor U14793 (N_14793,N_14525,N_14510);
nor U14794 (N_14794,N_14564,N_14665);
nor U14795 (N_14795,N_14560,N_14569);
and U14796 (N_14796,N_14716,N_14508);
nor U14797 (N_14797,N_14725,N_14683);
xor U14798 (N_14798,N_14617,N_14677);
or U14799 (N_14799,N_14719,N_14570);
or U14800 (N_14800,N_14639,N_14640);
and U14801 (N_14801,N_14648,N_14566);
nor U14802 (N_14802,N_14721,N_14518);
xor U14803 (N_14803,N_14705,N_14581);
nand U14804 (N_14804,N_14675,N_14586);
or U14805 (N_14805,N_14563,N_14537);
xnor U14806 (N_14806,N_14709,N_14649);
and U14807 (N_14807,N_14735,N_14610);
xnor U14808 (N_14808,N_14654,N_14606);
nor U14809 (N_14809,N_14549,N_14600);
nor U14810 (N_14810,N_14598,N_14742);
and U14811 (N_14811,N_14684,N_14690);
nand U14812 (N_14812,N_14544,N_14637);
xnor U14813 (N_14813,N_14580,N_14535);
nor U14814 (N_14814,N_14554,N_14522);
nor U14815 (N_14815,N_14660,N_14718);
nand U14816 (N_14816,N_14745,N_14507);
and U14817 (N_14817,N_14715,N_14707);
and U14818 (N_14818,N_14511,N_14532);
nand U14819 (N_14819,N_14571,N_14618);
xor U14820 (N_14820,N_14538,N_14555);
or U14821 (N_14821,N_14585,N_14655);
or U14822 (N_14822,N_14738,N_14548);
nor U14823 (N_14823,N_14702,N_14521);
nor U14824 (N_14824,N_14671,N_14531);
nor U14825 (N_14825,N_14712,N_14514);
or U14826 (N_14826,N_14575,N_14728);
xnor U14827 (N_14827,N_14616,N_14604);
xor U14828 (N_14828,N_14734,N_14620);
and U14829 (N_14829,N_14559,N_14529);
nor U14830 (N_14830,N_14646,N_14625);
or U14831 (N_14831,N_14624,N_14609);
nand U14832 (N_14832,N_14729,N_14543);
xor U14833 (N_14833,N_14530,N_14743);
nand U14834 (N_14834,N_14572,N_14659);
nor U14835 (N_14835,N_14644,N_14740);
nor U14836 (N_14836,N_14594,N_14540);
xor U14837 (N_14837,N_14630,N_14524);
nand U14838 (N_14838,N_14694,N_14632);
and U14839 (N_14839,N_14681,N_14710);
and U14840 (N_14840,N_14656,N_14623);
nor U14841 (N_14841,N_14661,N_14706);
nand U14842 (N_14842,N_14723,N_14638);
and U14843 (N_14843,N_14746,N_14701);
nor U14844 (N_14844,N_14676,N_14553);
nand U14845 (N_14845,N_14557,N_14673);
nand U14846 (N_14846,N_14612,N_14647);
xnor U14847 (N_14847,N_14697,N_14503);
or U14848 (N_14848,N_14739,N_14693);
nor U14849 (N_14849,N_14513,N_14546);
nand U14850 (N_14850,N_14635,N_14504);
or U14851 (N_14851,N_14613,N_14577);
nand U14852 (N_14852,N_14703,N_14517);
or U14853 (N_14853,N_14704,N_14737);
and U14854 (N_14854,N_14515,N_14741);
nor U14855 (N_14855,N_14691,N_14678);
nor U14856 (N_14856,N_14736,N_14568);
nor U14857 (N_14857,N_14669,N_14519);
and U14858 (N_14858,N_14747,N_14536);
and U14859 (N_14859,N_14631,N_14576);
nor U14860 (N_14860,N_14596,N_14509);
xor U14861 (N_14861,N_14664,N_14615);
nor U14862 (N_14862,N_14512,N_14556);
or U14863 (N_14863,N_14680,N_14698);
xor U14864 (N_14864,N_14603,N_14545);
nand U14865 (N_14865,N_14622,N_14607);
nand U14866 (N_14866,N_14574,N_14711);
nand U14867 (N_14867,N_14520,N_14645);
nand U14868 (N_14868,N_14539,N_14528);
nand U14869 (N_14869,N_14667,N_14650);
or U14870 (N_14870,N_14501,N_14597);
nor U14871 (N_14871,N_14592,N_14621);
and U14872 (N_14872,N_14561,N_14611);
and U14873 (N_14873,N_14724,N_14629);
nor U14874 (N_14874,N_14601,N_14558);
nor U14875 (N_14875,N_14611,N_14515);
or U14876 (N_14876,N_14609,N_14520);
or U14877 (N_14877,N_14622,N_14597);
and U14878 (N_14878,N_14683,N_14545);
nand U14879 (N_14879,N_14555,N_14723);
and U14880 (N_14880,N_14664,N_14746);
nor U14881 (N_14881,N_14589,N_14632);
xor U14882 (N_14882,N_14710,N_14715);
xnor U14883 (N_14883,N_14628,N_14571);
and U14884 (N_14884,N_14655,N_14620);
or U14885 (N_14885,N_14540,N_14678);
nand U14886 (N_14886,N_14686,N_14595);
nand U14887 (N_14887,N_14576,N_14574);
and U14888 (N_14888,N_14505,N_14593);
and U14889 (N_14889,N_14633,N_14719);
and U14890 (N_14890,N_14602,N_14503);
xnor U14891 (N_14891,N_14501,N_14690);
nand U14892 (N_14892,N_14598,N_14739);
or U14893 (N_14893,N_14546,N_14589);
nand U14894 (N_14894,N_14603,N_14618);
and U14895 (N_14895,N_14550,N_14610);
nor U14896 (N_14896,N_14654,N_14547);
or U14897 (N_14897,N_14500,N_14694);
and U14898 (N_14898,N_14536,N_14524);
nor U14899 (N_14899,N_14675,N_14552);
xor U14900 (N_14900,N_14574,N_14745);
nor U14901 (N_14901,N_14627,N_14659);
and U14902 (N_14902,N_14734,N_14525);
nand U14903 (N_14903,N_14637,N_14595);
nor U14904 (N_14904,N_14727,N_14697);
xor U14905 (N_14905,N_14686,N_14648);
nand U14906 (N_14906,N_14596,N_14658);
nand U14907 (N_14907,N_14556,N_14507);
or U14908 (N_14908,N_14558,N_14723);
nor U14909 (N_14909,N_14551,N_14520);
and U14910 (N_14910,N_14718,N_14709);
nor U14911 (N_14911,N_14557,N_14566);
nand U14912 (N_14912,N_14567,N_14556);
xor U14913 (N_14913,N_14614,N_14663);
nand U14914 (N_14914,N_14675,N_14632);
nand U14915 (N_14915,N_14578,N_14518);
or U14916 (N_14916,N_14563,N_14747);
nor U14917 (N_14917,N_14662,N_14616);
and U14918 (N_14918,N_14595,N_14699);
or U14919 (N_14919,N_14662,N_14526);
nand U14920 (N_14920,N_14740,N_14629);
xnor U14921 (N_14921,N_14548,N_14534);
or U14922 (N_14922,N_14605,N_14538);
nor U14923 (N_14923,N_14599,N_14613);
or U14924 (N_14924,N_14660,N_14741);
or U14925 (N_14925,N_14630,N_14699);
nand U14926 (N_14926,N_14596,N_14603);
nor U14927 (N_14927,N_14748,N_14549);
or U14928 (N_14928,N_14705,N_14655);
or U14929 (N_14929,N_14747,N_14525);
nand U14930 (N_14930,N_14533,N_14733);
nand U14931 (N_14931,N_14634,N_14703);
nand U14932 (N_14932,N_14672,N_14693);
nor U14933 (N_14933,N_14576,N_14732);
and U14934 (N_14934,N_14688,N_14562);
and U14935 (N_14935,N_14589,N_14658);
or U14936 (N_14936,N_14604,N_14701);
and U14937 (N_14937,N_14519,N_14696);
and U14938 (N_14938,N_14603,N_14713);
xor U14939 (N_14939,N_14501,N_14708);
xnor U14940 (N_14940,N_14688,N_14650);
xor U14941 (N_14941,N_14742,N_14687);
xnor U14942 (N_14942,N_14724,N_14680);
or U14943 (N_14943,N_14516,N_14616);
xor U14944 (N_14944,N_14526,N_14532);
xor U14945 (N_14945,N_14682,N_14649);
nand U14946 (N_14946,N_14655,N_14521);
xor U14947 (N_14947,N_14744,N_14695);
xnor U14948 (N_14948,N_14676,N_14704);
nor U14949 (N_14949,N_14564,N_14608);
nor U14950 (N_14950,N_14734,N_14711);
and U14951 (N_14951,N_14597,N_14626);
or U14952 (N_14952,N_14597,N_14589);
xor U14953 (N_14953,N_14551,N_14726);
or U14954 (N_14954,N_14572,N_14730);
nor U14955 (N_14955,N_14575,N_14576);
nand U14956 (N_14956,N_14664,N_14667);
or U14957 (N_14957,N_14570,N_14661);
and U14958 (N_14958,N_14718,N_14707);
xor U14959 (N_14959,N_14634,N_14666);
xor U14960 (N_14960,N_14609,N_14566);
xnor U14961 (N_14961,N_14528,N_14632);
or U14962 (N_14962,N_14701,N_14669);
and U14963 (N_14963,N_14740,N_14697);
nand U14964 (N_14964,N_14689,N_14509);
xor U14965 (N_14965,N_14573,N_14571);
nand U14966 (N_14966,N_14599,N_14742);
and U14967 (N_14967,N_14604,N_14583);
xnor U14968 (N_14968,N_14513,N_14516);
or U14969 (N_14969,N_14673,N_14537);
and U14970 (N_14970,N_14658,N_14524);
nand U14971 (N_14971,N_14609,N_14522);
and U14972 (N_14972,N_14748,N_14733);
or U14973 (N_14973,N_14542,N_14689);
xor U14974 (N_14974,N_14530,N_14558);
nand U14975 (N_14975,N_14558,N_14584);
nand U14976 (N_14976,N_14617,N_14589);
xnor U14977 (N_14977,N_14560,N_14565);
nor U14978 (N_14978,N_14605,N_14723);
xor U14979 (N_14979,N_14538,N_14640);
xor U14980 (N_14980,N_14554,N_14690);
nand U14981 (N_14981,N_14576,N_14647);
nor U14982 (N_14982,N_14642,N_14645);
nand U14983 (N_14983,N_14586,N_14536);
or U14984 (N_14984,N_14706,N_14622);
or U14985 (N_14985,N_14565,N_14720);
and U14986 (N_14986,N_14730,N_14682);
xnor U14987 (N_14987,N_14616,N_14568);
nand U14988 (N_14988,N_14611,N_14649);
nand U14989 (N_14989,N_14551,N_14623);
nand U14990 (N_14990,N_14725,N_14610);
nor U14991 (N_14991,N_14689,N_14606);
xor U14992 (N_14992,N_14575,N_14549);
nor U14993 (N_14993,N_14584,N_14556);
nor U14994 (N_14994,N_14570,N_14622);
and U14995 (N_14995,N_14659,N_14502);
or U14996 (N_14996,N_14673,N_14717);
or U14997 (N_14997,N_14682,N_14523);
nand U14998 (N_14998,N_14521,N_14563);
nand U14999 (N_14999,N_14596,N_14574);
nand UO_0 (O_0,N_14958,N_14833);
nor UO_1 (O_1,N_14901,N_14788);
nor UO_2 (O_2,N_14826,N_14801);
xnor UO_3 (O_3,N_14979,N_14880);
or UO_4 (O_4,N_14997,N_14774);
nor UO_5 (O_5,N_14882,N_14893);
nand UO_6 (O_6,N_14789,N_14797);
nand UO_7 (O_7,N_14839,N_14957);
nor UO_8 (O_8,N_14910,N_14886);
nand UO_9 (O_9,N_14920,N_14761);
or UO_10 (O_10,N_14951,N_14853);
and UO_11 (O_11,N_14806,N_14998);
and UO_12 (O_12,N_14768,N_14929);
nor UO_13 (O_13,N_14778,N_14786);
xnor UO_14 (O_14,N_14887,N_14904);
or UO_15 (O_15,N_14900,N_14837);
or UO_16 (O_16,N_14995,N_14800);
nor UO_17 (O_17,N_14984,N_14857);
nor UO_18 (O_18,N_14969,N_14851);
xnor UO_19 (O_19,N_14828,N_14754);
nand UO_20 (O_20,N_14898,N_14945);
and UO_21 (O_21,N_14803,N_14885);
nor UO_22 (O_22,N_14794,N_14936);
and UO_23 (O_23,N_14988,N_14755);
nand UO_24 (O_24,N_14991,N_14807);
or UO_25 (O_25,N_14975,N_14913);
nand UO_26 (O_26,N_14770,N_14932);
or UO_27 (O_27,N_14869,N_14854);
or UO_28 (O_28,N_14841,N_14883);
or UO_29 (O_29,N_14923,N_14962);
nand UO_30 (O_30,N_14971,N_14859);
xor UO_31 (O_31,N_14934,N_14821);
xnor UO_32 (O_32,N_14863,N_14888);
and UO_33 (O_33,N_14987,N_14909);
or UO_34 (O_34,N_14960,N_14844);
nand UO_35 (O_35,N_14965,N_14889);
xnor UO_36 (O_36,N_14937,N_14915);
nor UO_37 (O_37,N_14750,N_14921);
nand UO_38 (O_38,N_14813,N_14831);
nand UO_39 (O_39,N_14911,N_14875);
and UO_40 (O_40,N_14899,N_14925);
nor UO_41 (O_41,N_14779,N_14842);
xor UO_42 (O_42,N_14762,N_14773);
or UO_43 (O_43,N_14815,N_14798);
or UO_44 (O_44,N_14760,N_14940);
xnor UO_45 (O_45,N_14799,N_14787);
and UO_46 (O_46,N_14771,N_14986);
and UO_47 (O_47,N_14756,N_14766);
xor UO_48 (O_48,N_14825,N_14784);
xor UO_49 (O_49,N_14918,N_14845);
or UO_50 (O_50,N_14823,N_14968);
nor UO_51 (O_51,N_14930,N_14757);
nand UO_52 (O_52,N_14895,N_14878);
or UO_53 (O_53,N_14926,N_14956);
and UO_54 (O_54,N_14812,N_14811);
or UO_55 (O_55,N_14871,N_14941);
nor UO_56 (O_56,N_14783,N_14856);
nor UO_57 (O_57,N_14976,N_14876);
and UO_58 (O_58,N_14974,N_14922);
or UO_59 (O_59,N_14972,N_14892);
xor UO_60 (O_60,N_14805,N_14989);
nor UO_61 (O_61,N_14919,N_14765);
nand UO_62 (O_62,N_14830,N_14793);
nor UO_63 (O_63,N_14785,N_14843);
nand UO_64 (O_64,N_14917,N_14752);
xnor UO_65 (O_65,N_14870,N_14818);
and UO_66 (O_66,N_14817,N_14804);
or UO_67 (O_67,N_14847,N_14903);
xor UO_68 (O_68,N_14967,N_14874);
nor UO_69 (O_69,N_14810,N_14816);
and UO_70 (O_70,N_14855,N_14907);
nor UO_71 (O_71,N_14942,N_14873);
nand UO_72 (O_72,N_14840,N_14890);
and UO_73 (O_73,N_14916,N_14924);
and UO_74 (O_74,N_14795,N_14867);
or UO_75 (O_75,N_14849,N_14781);
or UO_76 (O_76,N_14931,N_14946);
nand UO_77 (O_77,N_14758,N_14767);
nand UO_78 (O_78,N_14834,N_14927);
and UO_79 (O_79,N_14906,N_14964);
and UO_80 (O_80,N_14759,N_14884);
and UO_81 (O_81,N_14829,N_14996);
nand UO_82 (O_82,N_14905,N_14838);
nor UO_83 (O_83,N_14836,N_14792);
and UO_84 (O_84,N_14777,N_14928);
and UO_85 (O_85,N_14999,N_14814);
nand UO_86 (O_86,N_14963,N_14862);
and UO_87 (O_87,N_14990,N_14802);
nand UO_88 (O_88,N_14982,N_14973);
and UO_89 (O_89,N_14808,N_14877);
or UO_90 (O_90,N_14881,N_14978);
xnor UO_91 (O_91,N_14948,N_14981);
xor UO_92 (O_92,N_14866,N_14947);
or UO_93 (O_93,N_14796,N_14912);
or UO_94 (O_94,N_14860,N_14872);
or UO_95 (O_95,N_14902,N_14954);
xor UO_96 (O_96,N_14846,N_14858);
nand UO_97 (O_97,N_14961,N_14776);
xor UO_98 (O_98,N_14955,N_14935);
xor UO_99 (O_99,N_14952,N_14820);
nor UO_100 (O_100,N_14914,N_14850);
or UO_101 (O_101,N_14835,N_14827);
or UO_102 (O_102,N_14751,N_14775);
or UO_103 (O_103,N_14769,N_14943);
or UO_104 (O_104,N_14824,N_14896);
xor UO_105 (O_105,N_14992,N_14966);
and UO_106 (O_106,N_14953,N_14983);
and UO_107 (O_107,N_14891,N_14809);
nor UO_108 (O_108,N_14938,N_14753);
and UO_109 (O_109,N_14861,N_14864);
nand UO_110 (O_110,N_14950,N_14782);
and UO_111 (O_111,N_14832,N_14994);
or UO_112 (O_112,N_14939,N_14879);
xor UO_113 (O_113,N_14897,N_14959);
nor UO_114 (O_114,N_14763,N_14865);
and UO_115 (O_115,N_14933,N_14868);
xnor UO_116 (O_116,N_14852,N_14908);
xnor UO_117 (O_117,N_14993,N_14780);
nor UO_118 (O_118,N_14985,N_14949);
nor UO_119 (O_119,N_14980,N_14944);
or UO_120 (O_120,N_14970,N_14772);
or UO_121 (O_121,N_14791,N_14977);
nand UO_122 (O_122,N_14822,N_14790);
and UO_123 (O_123,N_14848,N_14894);
nor UO_124 (O_124,N_14819,N_14764);
nand UO_125 (O_125,N_14877,N_14845);
or UO_126 (O_126,N_14982,N_14754);
or UO_127 (O_127,N_14992,N_14872);
nand UO_128 (O_128,N_14956,N_14817);
nor UO_129 (O_129,N_14772,N_14819);
or UO_130 (O_130,N_14966,N_14982);
xor UO_131 (O_131,N_14814,N_14837);
and UO_132 (O_132,N_14842,N_14972);
nor UO_133 (O_133,N_14919,N_14831);
nand UO_134 (O_134,N_14947,N_14808);
or UO_135 (O_135,N_14879,N_14770);
and UO_136 (O_136,N_14827,N_14922);
nor UO_137 (O_137,N_14985,N_14759);
or UO_138 (O_138,N_14991,N_14978);
nor UO_139 (O_139,N_14937,N_14850);
xnor UO_140 (O_140,N_14867,N_14851);
and UO_141 (O_141,N_14898,N_14979);
nor UO_142 (O_142,N_14932,N_14813);
nor UO_143 (O_143,N_14776,N_14848);
nor UO_144 (O_144,N_14982,N_14812);
nand UO_145 (O_145,N_14840,N_14810);
or UO_146 (O_146,N_14787,N_14994);
and UO_147 (O_147,N_14920,N_14876);
nor UO_148 (O_148,N_14792,N_14819);
or UO_149 (O_149,N_14799,N_14948);
nor UO_150 (O_150,N_14801,N_14898);
and UO_151 (O_151,N_14753,N_14860);
and UO_152 (O_152,N_14911,N_14863);
or UO_153 (O_153,N_14949,N_14973);
nor UO_154 (O_154,N_14854,N_14950);
and UO_155 (O_155,N_14785,N_14829);
nand UO_156 (O_156,N_14873,N_14893);
or UO_157 (O_157,N_14784,N_14793);
and UO_158 (O_158,N_14956,N_14830);
nand UO_159 (O_159,N_14974,N_14869);
nand UO_160 (O_160,N_14880,N_14844);
nor UO_161 (O_161,N_14858,N_14864);
and UO_162 (O_162,N_14980,N_14989);
nor UO_163 (O_163,N_14986,N_14910);
xor UO_164 (O_164,N_14857,N_14753);
nand UO_165 (O_165,N_14938,N_14922);
xnor UO_166 (O_166,N_14792,N_14988);
xnor UO_167 (O_167,N_14839,N_14878);
nor UO_168 (O_168,N_14846,N_14767);
or UO_169 (O_169,N_14881,N_14975);
and UO_170 (O_170,N_14883,N_14923);
or UO_171 (O_171,N_14986,N_14798);
nor UO_172 (O_172,N_14892,N_14753);
xnor UO_173 (O_173,N_14829,N_14768);
nand UO_174 (O_174,N_14992,N_14969);
nand UO_175 (O_175,N_14926,N_14903);
or UO_176 (O_176,N_14943,N_14782);
nand UO_177 (O_177,N_14880,N_14939);
or UO_178 (O_178,N_14856,N_14778);
nand UO_179 (O_179,N_14947,N_14921);
and UO_180 (O_180,N_14876,N_14779);
xor UO_181 (O_181,N_14983,N_14916);
and UO_182 (O_182,N_14759,N_14914);
and UO_183 (O_183,N_14894,N_14903);
or UO_184 (O_184,N_14852,N_14932);
xor UO_185 (O_185,N_14952,N_14961);
or UO_186 (O_186,N_14781,N_14791);
nor UO_187 (O_187,N_14845,N_14995);
or UO_188 (O_188,N_14785,N_14954);
xor UO_189 (O_189,N_14900,N_14874);
and UO_190 (O_190,N_14981,N_14806);
and UO_191 (O_191,N_14886,N_14917);
and UO_192 (O_192,N_14880,N_14971);
xnor UO_193 (O_193,N_14945,N_14804);
and UO_194 (O_194,N_14893,N_14864);
or UO_195 (O_195,N_14903,N_14885);
or UO_196 (O_196,N_14829,N_14755);
nor UO_197 (O_197,N_14815,N_14929);
and UO_198 (O_198,N_14888,N_14774);
or UO_199 (O_199,N_14811,N_14914);
and UO_200 (O_200,N_14976,N_14809);
nor UO_201 (O_201,N_14904,N_14794);
xor UO_202 (O_202,N_14961,N_14814);
or UO_203 (O_203,N_14964,N_14973);
nor UO_204 (O_204,N_14780,N_14924);
nor UO_205 (O_205,N_14848,N_14881);
and UO_206 (O_206,N_14760,N_14972);
nand UO_207 (O_207,N_14771,N_14837);
nand UO_208 (O_208,N_14950,N_14905);
xor UO_209 (O_209,N_14832,N_14887);
nor UO_210 (O_210,N_14904,N_14962);
nor UO_211 (O_211,N_14967,N_14922);
nand UO_212 (O_212,N_14925,N_14773);
nor UO_213 (O_213,N_14856,N_14900);
and UO_214 (O_214,N_14842,N_14928);
and UO_215 (O_215,N_14983,N_14879);
or UO_216 (O_216,N_14829,N_14808);
and UO_217 (O_217,N_14771,N_14816);
nand UO_218 (O_218,N_14816,N_14821);
nand UO_219 (O_219,N_14894,N_14995);
or UO_220 (O_220,N_14768,N_14877);
or UO_221 (O_221,N_14794,N_14761);
and UO_222 (O_222,N_14767,N_14874);
or UO_223 (O_223,N_14798,N_14926);
nand UO_224 (O_224,N_14818,N_14774);
xnor UO_225 (O_225,N_14906,N_14762);
nor UO_226 (O_226,N_14766,N_14937);
xor UO_227 (O_227,N_14860,N_14776);
xnor UO_228 (O_228,N_14830,N_14995);
or UO_229 (O_229,N_14930,N_14891);
and UO_230 (O_230,N_14895,N_14773);
or UO_231 (O_231,N_14806,N_14883);
nor UO_232 (O_232,N_14997,N_14925);
or UO_233 (O_233,N_14822,N_14890);
nand UO_234 (O_234,N_14963,N_14901);
and UO_235 (O_235,N_14855,N_14863);
or UO_236 (O_236,N_14757,N_14899);
nand UO_237 (O_237,N_14928,N_14818);
nor UO_238 (O_238,N_14942,N_14850);
and UO_239 (O_239,N_14869,N_14804);
xnor UO_240 (O_240,N_14809,N_14933);
and UO_241 (O_241,N_14755,N_14986);
nor UO_242 (O_242,N_14898,N_14928);
nand UO_243 (O_243,N_14973,N_14935);
or UO_244 (O_244,N_14909,N_14935);
and UO_245 (O_245,N_14825,N_14894);
or UO_246 (O_246,N_14958,N_14866);
nor UO_247 (O_247,N_14761,N_14899);
xor UO_248 (O_248,N_14754,N_14890);
and UO_249 (O_249,N_14891,N_14989);
nor UO_250 (O_250,N_14903,N_14782);
or UO_251 (O_251,N_14878,N_14835);
nand UO_252 (O_252,N_14788,N_14821);
nor UO_253 (O_253,N_14881,N_14800);
and UO_254 (O_254,N_14774,N_14939);
nor UO_255 (O_255,N_14829,N_14752);
xnor UO_256 (O_256,N_14947,N_14839);
xnor UO_257 (O_257,N_14980,N_14885);
nand UO_258 (O_258,N_14912,N_14782);
xor UO_259 (O_259,N_14982,N_14939);
and UO_260 (O_260,N_14811,N_14783);
or UO_261 (O_261,N_14996,N_14998);
nor UO_262 (O_262,N_14863,N_14903);
or UO_263 (O_263,N_14824,N_14917);
and UO_264 (O_264,N_14918,N_14939);
xor UO_265 (O_265,N_14842,N_14927);
xnor UO_266 (O_266,N_14763,N_14851);
nand UO_267 (O_267,N_14809,N_14953);
xor UO_268 (O_268,N_14817,N_14939);
and UO_269 (O_269,N_14882,N_14894);
xnor UO_270 (O_270,N_14882,N_14959);
nand UO_271 (O_271,N_14916,N_14895);
nor UO_272 (O_272,N_14901,N_14982);
or UO_273 (O_273,N_14822,N_14805);
nor UO_274 (O_274,N_14855,N_14849);
and UO_275 (O_275,N_14846,N_14785);
or UO_276 (O_276,N_14993,N_14768);
and UO_277 (O_277,N_14783,N_14799);
and UO_278 (O_278,N_14767,N_14870);
xnor UO_279 (O_279,N_14981,N_14807);
or UO_280 (O_280,N_14984,N_14791);
nand UO_281 (O_281,N_14970,N_14761);
xor UO_282 (O_282,N_14927,N_14852);
or UO_283 (O_283,N_14898,N_14896);
xnor UO_284 (O_284,N_14812,N_14971);
and UO_285 (O_285,N_14866,N_14854);
or UO_286 (O_286,N_14903,N_14827);
and UO_287 (O_287,N_14974,N_14970);
or UO_288 (O_288,N_14839,N_14812);
xor UO_289 (O_289,N_14904,N_14958);
or UO_290 (O_290,N_14808,N_14762);
or UO_291 (O_291,N_14940,N_14789);
and UO_292 (O_292,N_14999,N_14861);
and UO_293 (O_293,N_14869,N_14908);
nor UO_294 (O_294,N_14845,N_14914);
xor UO_295 (O_295,N_14860,N_14901);
and UO_296 (O_296,N_14945,N_14845);
nand UO_297 (O_297,N_14938,N_14858);
and UO_298 (O_298,N_14805,N_14976);
or UO_299 (O_299,N_14770,N_14819);
and UO_300 (O_300,N_14908,N_14808);
xnor UO_301 (O_301,N_14955,N_14875);
or UO_302 (O_302,N_14834,N_14760);
nor UO_303 (O_303,N_14850,N_14774);
nand UO_304 (O_304,N_14895,N_14922);
nor UO_305 (O_305,N_14891,N_14963);
and UO_306 (O_306,N_14785,N_14862);
and UO_307 (O_307,N_14888,N_14904);
xor UO_308 (O_308,N_14859,N_14852);
nand UO_309 (O_309,N_14990,N_14946);
nor UO_310 (O_310,N_14820,N_14999);
or UO_311 (O_311,N_14821,N_14914);
xnor UO_312 (O_312,N_14951,N_14859);
xnor UO_313 (O_313,N_14767,N_14916);
nand UO_314 (O_314,N_14753,N_14803);
xor UO_315 (O_315,N_14967,N_14935);
and UO_316 (O_316,N_14984,N_14830);
nand UO_317 (O_317,N_14983,N_14874);
and UO_318 (O_318,N_14804,N_14972);
nand UO_319 (O_319,N_14964,N_14965);
or UO_320 (O_320,N_14827,N_14875);
and UO_321 (O_321,N_14973,N_14905);
and UO_322 (O_322,N_14862,N_14983);
or UO_323 (O_323,N_14849,N_14949);
xor UO_324 (O_324,N_14750,N_14990);
xnor UO_325 (O_325,N_14828,N_14775);
nand UO_326 (O_326,N_14989,N_14825);
nand UO_327 (O_327,N_14872,N_14942);
or UO_328 (O_328,N_14896,N_14751);
or UO_329 (O_329,N_14772,N_14768);
xor UO_330 (O_330,N_14884,N_14928);
nand UO_331 (O_331,N_14757,N_14857);
nor UO_332 (O_332,N_14953,N_14965);
or UO_333 (O_333,N_14935,N_14928);
nor UO_334 (O_334,N_14873,N_14955);
xor UO_335 (O_335,N_14834,N_14900);
or UO_336 (O_336,N_14823,N_14999);
xor UO_337 (O_337,N_14820,N_14937);
nand UO_338 (O_338,N_14782,N_14784);
or UO_339 (O_339,N_14956,N_14789);
nor UO_340 (O_340,N_14889,N_14980);
or UO_341 (O_341,N_14882,N_14924);
xor UO_342 (O_342,N_14829,N_14810);
xnor UO_343 (O_343,N_14908,N_14916);
nand UO_344 (O_344,N_14876,N_14979);
nor UO_345 (O_345,N_14798,N_14865);
and UO_346 (O_346,N_14750,N_14760);
or UO_347 (O_347,N_14891,N_14839);
and UO_348 (O_348,N_14866,N_14884);
xor UO_349 (O_349,N_14905,N_14908);
or UO_350 (O_350,N_14886,N_14982);
nand UO_351 (O_351,N_14885,N_14932);
or UO_352 (O_352,N_14910,N_14871);
or UO_353 (O_353,N_14847,N_14915);
nor UO_354 (O_354,N_14865,N_14774);
nor UO_355 (O_355,N_14871,N_14809);
or UO_356 (O_356,N_14994,N_14846);
nor UO_357 (O_357,N_14887,N_14981);
or UO_358 (O_358,N_14811,N_14807);
or UO_359 (O_359,N_14965,N_14891);
xor UO_360 (O_360,N_14941,N_14913);
nor UO_361 (O_361,N_14752,N_14925);
xnor UO_362 (O_362,N_14925,N_14769);
and UO_363 (O_363,N_14988,N_14974);
or UO_364 (O_364,N_14799,N_14814);
xnor UO_365 (O_365,N_14827,N_14772);
and UO_366 (O_366,N_14890,N_14794);
or UO_367 (O_367,N_14901,N_14876);
or UO_368 (O_368,N_14980,N_14898);
xnor UO_369 (O_369,N_14877,N_14793);
and UO_370 (O_370,N_14994,N_14753);
nor UO_371 (O_371,N_14993,N_14851);
nor UO_372 (O_372,N_14755,N_14871);
nand UO_373 (O_373,N_14890,N_14790);
or UO_374 (O_374,N_14942,N_14800);
nand UO_375 (O_375,N_14817,N_14905);
nor UO_376 (O_376,N_14837,N_14757);
or UO_377 (O_377,N_14943,N_14879);
xnor UO_378 (O_378,N_14890,N_14968);
nor UO_379 (O_379,N_14847,N_14798);
nor UO_380 (O_380,N_14815,N_14960);
xnor UO_381 (O_381,N_14965,N_14868);
and UO_382 (O_382,N_14915,N_14971);
or UO_383 (O_383,N_14883,N_14942);
xnor UO_384 (O_384,N_14758,N_14871);
xnor UO_385 (O_385,N_14973,N_14834);
nand UO_386 (O_386,N_14824,N_14926);
and UO_387 (O_387,N_14994,N_14811);
or UO_388 (O_388,N_14864,N_14875);
nor UO_389 (O_389,N_14776,N_14983);
nor UO_390 (O_390,N_14934,N_14933);
or UO_391 (O_391,N_14768,N_14805);
and UO_392 (O_392,N_14826,N_14889);
nor UO_393 (O_393,N_14943,N_14989);
xor UO_394 (O_394,N_14901,N_14848);
nand UO_395 (O_395,N_14869,N_14970);
nand UO_396 (O_396,N_14879,N_14863);
xnor UO_397 (O_397,N_14904,N_14834);
xor UO_398 (O_398,N_14815,N_14993);
nor UO_399 (O_399,N_14863,N_14894);
nor UO_400 (O_400,N_14830,N_14928);
xnor UO_401 (O_401,N_14810,N_14930);
or UO_402 (O_402,N_14806,N_14923);
and UO_403 (O_403,N_14799,N_14846);
nand UO_404 (O_404,N_14977,N_14883);
or UO_405 (O_405,N_14750,N_14936);
or UO_406 (O_406,N_14882,N_14910);
nor UO_407 (O_407,N_14922,N_14852);
and UO_408 (O_408,N_14990,N_14895);
or UO_409 (O_409,N_14805,N_14953);
xnor UO_410 (O_410,N_14961,N_14803);
nand UO_411 (O_411,N_14799,N_14947);
nor UO_412 (O_412,N_14768,N_14990);
xnor UO_413 (O_413,N_14759,N_14997);
nand UO_414 (O_414,N_14772,N_14938);
xnor UO_415 (O_415,N_14765,N_14850);
nor UO_416 (O_416,N_14872,N_14870);
nor UO_417 (O_417,N_14757,N_14785);
and UO_418 (O_418,N_14964,N_14820);
nor UO_419 (O_419,N_14801,N_14956);
nand UO_420 (O_420,N_14967,N_14893);
and UO_421 (O_421,N_14971,N_14911);
and UO_422 (O_422,N_14869,N_14858);
or UO_423 (O_423,N_14779,N_14820);
xor UO_424 (O_424,N_14882,N_14914);
or UO_425 (O_425,N_14938,N_14774);
xor UO_426 (O_426,N_14983,N_14944);
and UO_427 (O_427,N_14880,N_14976);
nand UO_428 (O_428,N_14912,N_14987);
xnor UO_429 (O_429,N_14828,N_14810);
or UO_430 (O_430,N_14850,N_14794);
or UO_431 (O_431,N_14977,N_14753);
nor UO_432 (O_432,N_14917,N_14813);
and UO_433 (O_433,N_14919,N_14811);
nor UO_434 (O_434,N_14937,N_14980);
nor UO_435 (O_435,N_14915,N_14968);
nor UO_436 (O_436,N_14826,N_14806);
nor UO_437 (O_437,N_14852,N_14874);
and UO_438 (O_438,N_14911,N_14872);
xnor UO_439 (O_439,N_14908,N_14839);
nor UO_440 (O_440,N_14782,N_14955);
or UO_441 (O_441,N_14868,N_14768);
nand UO_442 (O_442,N_14778,N_14999);
and UO_443 (O_443,N_14892,N_14993);
nor UO_444 (O_444,N_14828,N_14902);
nor UO_445 (O_445,N_14968,N_14826);
nand UO_446 (O_446,N_14946,N_14972);
and UO_447 (O_447,N_14981,N_14855);
xor UO_448 (O_448,N_14903,N_14757);
and UO_449 (O_449,N_14798,N_14891);
xor UO_450 (O_450,N_14942,N_14781);
nor UO_451 (O_451,N_14751,N_14845);
nor UO_452 (O_452,N_14980,N_14886);
xnor UO_453 (O_453,N_14762,N_14830);
nor UO_454 (O_454,N_14844,N_14821);
nand UO_455 (O_455,N_14915,N_14890);
nor UO_456 (O_456,N_14882,N_14913);
nand UO_457 (O_457,N_14833,N_14806);
and UO_458 (O_458,N_14924,N_14906);
xnor UO_459 (O_459,N_14907,N_14877);
xnor UO_460 (O_460,N_14984,N_14920);
or UO_461 (O_461,N_14989,N_14924);
xor UO_462 (O_462,N_14908,N_14971);
nor UO_463 (O_463,N_14769,N_14811);
nor UO_464 (O_464,N_14848,N_14948);
xor UO_465 (O_465,N_14896,N_14946);
nor UO_466 (O_466,N_14993,N_14884);
or UO_467 (O_467,N_14998,N_14834);
or UO_468 (O_468,N_14973,N_14943);
xor UO_469 (O_469,N_14894,N_14773);
and UO_470 (O_470,N_14900,N_14860);
nor UO_471 (O_471,N_14875,N_14771);
xnor UO_472 (O_472,N_14893,N_14977);
xor UO_473 (O_473,N_14849,N_14839);
or UO_474 (O_474,N_14919,N_14949);
xnor UO_475 (O_475,N_14772,N_14862);
nor UO_476 (O_476,N_14752,N_14924);
or UO_477 (O_477,N_14942,N_14932);
and UO_478 (O_478,N_14993,N_14875);
and UO_479 (O_479,N_14751,N_14914);
xnor UO_480 (O_480,N_14829,N_14828);
nand UO_481 (O_481,N_14969,N_14973);
and UO_482 (O_482,N_14968,N_14767);
nand UO_483 (O_483,N_14771,N_14898);
and UO_484 (O_484,N_14925,N_14859);
nor UO_485 (O_485,N_14916,N_14925);
or UO_486 (O_486,N_14984,N_14789);
nand UO_487 (O_487,N_14814,N_14769);
xnor UO_488 (O_488,N_14981,N_14960);
or UO_489 (O_489,N_14933,N_14835);
xnor UO_490 (O_490,N_14939,N_14750);
xor UO_491 (O_491,N_14895,N_14821);
nor UO_492 (O_492,N_14944,N_14855);
and UO_493 (O_493,N_14862,N_14858);
nand UO_494 (O_494,N_14873,N_14940);
nor UO_495 (O_495,N_14909,N_14760);
xnor UO_496 (O_496,N_14757,N_14861);
nor UO_497 (O_497,N_14826,N_14807);
xor UO_498 (O_498,N_14983,N_14976);
or UO_499 (O_499,N_14937,N_14810);
or UO_500 (O_500,N_14911,N_14999);
or UO_501 (O_501,N_14940,N_14783);
xnor UO_502 (O_502,N_14981,N_14982);
nand UO_503 (O_503,N_14945,N_14968);
nand UO_504 (O_504,N_14848,N_14996);
xnor UO_505 (O_505,N_14846,N_14896);
and UO_506 (O_506,N_14995,N_14960);
and UO_507 (O_507,N_14760,N_14914);
nor UO_508 (O_508,N_14924,N_14808);
nand UO_509 (O_509,N_14774,N_14821);
and UO_510 (O_510,N_14761,N_14913);
or UO_511 (O_511,N_14891,N_14797);
nand UO_512 (O_512,N_14990,N_14847);
nand UO_513 (O_513,N_14801,N_14839);
nand UO_514 (O_514,N_14997,N_14891);
xnor UO_515 (O_515,N_14838,N_14853);
and UO_516 (O_516,N_14937,N_14913);
or UO_517 (O_517,N_14933,N_14932);
and UO_518 (O_518,N_14888,N_14920);
xnor UO_519 (O_519,N_14890,N_14778);
or UO_520 (O_520,N_14770,N_14823);
or UO_521 (O_521,N_14786,N_14770);
nor UO_522 (O_522,N_14840,N_14891);
and UO_523 (O_523,N_14758,N_14846);
xor UO_524 (O_524,N_14789,N_14931);
xor UO_525 (O_525,N_14909,N_14820);
nand UO_526 (O_526,N_14912,N_14866);
or UO_527 (O_527,N_14852,N_14946);
nor UO_528 (O_528,N_14821,N_14871);
and UO_529 (O_529,N_14932,N_14784);
or UO_530 (O_530,N_14978,N_14822);
and UO_531 (O_531,N_14941,N_14838);
or UO_532 (O_532,N_14842,N_14994);
or UO_533 (O_533,N_14991,N_14928);
and UO_534 (O_534,N_14942,N_14998);
xor UO_535 (O_535,N_14863,N_14967);
nand UO_536 (O_536,N_14836,N_14903);
nor UO_537 (O_537,N_14925,N_14863);
nand UO_538 (O_538,N_14753,N_14871);
nand UO_539 (O_539,N_14834,N_14873);
nor UO_540 (O_540,N_14901,N_14904);
xor UO_541 (O_541,N_14858,N_14779);
xor UO_542 (O_542,N_14756,N_14948);
xor UO_543 (O_543,N_14819,N_14825);
and UO_544 (O_544,N_14942,N_14928);
or UO_545 (O_545,N_14864,N_14879);
or UO_546 (O_546,N_14876,N_14884);
and UO_547 (O_547,N_14969,N_14849);
nor UO_548 (O_548,N_14812,N_14999);
and UO_549 (O_549,N_14916,N_14992);
and UO_550 (O_550,N_14863,N_14849);
nor UO_551 (O_551,N_14763,N_14780);
and UO_552 (O_552,N_14864,N_14910);
xnor UO_553 (O_553,N_14757,N_14838);
or UO_554 (O_554,N_14783,N_14905);
xnor UO_555 (O_555,N_14974,N_14782);
nor UO_556 (O_556,N_14780,N_14922);
and UO_557 (O_557,N_14922,N_14912);
or UO_558 (O_558,N_14985,N_14769);
xor UO_559 (O_559,N_14972,N_14935);
or UO_560 (O_560,N_14855,N_14821);
xor UO_561 (O_561,N_14941,N_14877);
nand UO_562 (O_562,N_14813,N_14993);
nor UO_563 (O_563,N_14827,N_14890);
xor UO_564 (O_564,N_14966,N_14948);
or UO_565 (O_565,N_14803,N_14772);
nor UO_566 (O_566,N_14907,N_14974);
or UO_567 (O_567,N_14995,N_14863);
nor UO_568 (O_568,N_14762,N_14967);
nor UO_569 (O_569,N_14775,N_14832);
and UO_570 (O_570,N_14911,N_14788);
nand UO_571 (O_571,N_14842,N_14987);
or UO_572 (O_572,N_14895,N_14912);
nor UO_573 (O_573,N_14957,N_14964);
nor UO_574 (O_574,N_14766,N_14964);
nor UO_575 (O_575,N_14777,N_14833);
and UO_576 (O_576,N_14859,N_14840);
xor UO_577 (O_577,N_14987,N_14952);
xor UO_578 (O_578,N_14907,N_14900);
xor UO_579 (O_579,N_14985,N_14844);
nor UO_580 (O_580,N_14923,N_14959);
nor UO_581 (O_581,N_14850,N_14928);
and UO_582 (O_582,N_14983,N_14764);
nand UO_583 (O_583,N_14868,N_14855);
or UO_584 (O_584,N_14860,N_14960);
xor UO_585 (O_585,N_14997,N_14869);
or UO_586 (O_586,N_14916,N_14993);
or UO_587 (O_587,N_14921,N_14817);
or UO_588 (O_588,N_14839,N_14808);
or UO_589 (O_589,N_14921,N_14919);
and UO_590 (O_590,N_14893,N_14939);
xnor UO_591 (O_591,N_14908,N_14795);
and UO_592 (O_592,N_14862,N_14807);
nand UO_593 (O_593,N_14864,N_14971);
and UO_594 (O_594,N_14853,N_14831);
nand UO_595 (O_595,N_14855,N_14875);
xnor UO_596 (O_596,N_14824,N_14875);
xor UO_597 (O_597,N_14765,N_14879);
and UO_598 (O_598,N_14945,N_14934);
nand UO_599 (O_599,N_14841,N_14802);
nor UO_600 (O_600,N_14792,N_14960);
or UO_601 (O_601,N_14991,N_14919);
and UO_602 (O_602,N_14796,N_14871);
or UO_603 (O_603,N_14769,N_14998);
xor UO_604 (O_604,N_14900,N_14761);
nand UO_605 (O_605,N_14974,N_14979);
xor UO_606 (O_606,N_14904,N_14902);
xnor UO_607 (O_607,N_14953,N_14836);
nor UO_608 (O_608,N_14943,N_14952);
nand UO_609 (O_609,N_14882,N_14864);
or UO_610 (O_610,N_14795,N_14890);
or UO_611 (O_611,N_14886,N_14810);
xnor UO_612 (O_612,N_14855,N_14977);
nand UO_613 (O_613,N_14771,N_14932);
and UO_614 (O_614,N_14842,N_14887);
and UO_615 (O_615,N_14839,N_14877);
and UO_616 (O_616,N_14978,N_14954);
xnor UO_617 (O_617,N_14938,N_14986);
nor UO_618 (O_618,N_14948,N_14837);
and UO_619 (O_619,N_14864,N_14832);
and UO_620 (O_620,N_14817,N_14865);
nor UO_621 (O_621,N_14881,N_14986);
nand UO_622 (O_622,N_14917,N_14941);
and UO_623 (O_623,N_14954,N_14887);
or UO_624 (O_624,N_14964,N_14781);
xnor UO_625 (O_625,N_14933,N_14921);
xnor UO_626 (O_626,N_14853,N_14805);
xnor UO_627 (O_627,N_14874,N_14810);
or UO_628 (O_628,N_14873,N_14774);
xor UO_629 (O_629,N_14753,N_14906);
or UO_630 (O_630,N_14969,N_14876);
xor UO_631 (O_631,N_14845,N_14757);
nor UO_632 (O_632,N_14764,N_14809);
nor UO_633 (O_633,N_14885,N_14896);
xor UO_634 (O_634,N_14773,N_14929);
and UO_635 (O_635,N_14903,N_14949);
and UO_636 (O_636,N_14985,N_14901);
or UO_637 (O_637,N_14852,N_14775);
or UO_638 (O_638,N_14766,N_14864);
xnor UO_639 (O_639,N_14753,N_14785);
and UO_640 (O_640,N_14751,N_14825);
nand UO_641 (O_641,N_14919,N_14878);
nor UO_642 (O_642,N_14784,N_14830);
and UO_643 (O_643,N_14863,N_14876);
nand UO_644 (O_644,N_14938,N_14878);
nand UO_645 (O_645,N_14780,N_14875);
and UO_646 (O_646,N_14779,N_14808);
and UO_647 (O_647,N_14750,N_14978);
nand UO_648 (O_648,N_14945,N_14933);
nor UO_649 (O_649,N_14934,N_14872);
xnor UO_650 (O_650,N_14979,N_14903);
nand UO_651 (O_651,N_14751,N_14859);
xor UO_652 (O_652,N_14815,N_14920);
or UO_653 (O_653,N_14986,N_14827);
and UO_654 (O_654,N_14944,N_14846);
and UO_655 (O_655,N_14978,N_14887);
nand UO_656 (O_656,N_14756,N_14805);
nand UO_657 (O_657,N_14761,N_14921);
nand UO_658 (O_658,N_14910,N_14775);
nand UO_659 (O_659,N_14821,N_14803);
nor UO_660 (O_660,N_14986,N_14800);
xor UO_661 (O_661,N_14913,N_14899);
xnor UO_662 (O_662,N_14921,N_14870);
and UO_663 (O_663,N_14891,N_14860);
nor UO_664 (O_664,N_14800,N_14926);
or UO_665 (O_665,N_14764,N_14929);
xnor UO_666 (O_666,N_14812,N_14782);
nand UO_667 (O_667,N_14792,N_14798);
nor UO_668 (O_668,N_14841,N_14979);
or UO_669 (O_669,N_14997,N_14999);
and UO_670 (O_670,N_14912,N_14828);
nand UO_671 (O_671,N_14946,N_14815);
xor UO_672 (O_672,N_14792,N_14985);
nand UO_673 (O_673,N_14951,N_14760);
and UO_674 (O_674,N_14997,N_14877);
nand UO_675 (O_675,N_14855,N_14961);
xor UO_676 (O_676,N_14966,N_14863);
nor UO_677 (O_677,N_14977,N_14884);
xor UO_678 (O_678,N_14981,N_14856);
and UO_679 (O_679,N_14928,N_14767);
nand UO_680 (O_680,N_14871,N_14940);
xor UO_681 (O_681,N_14847,N_14959);
or UO_682 (O_682,N_14993,N_14870);
or UO_683 (O_683,N_14805,N_14983);
nor UO_684 (O_684,N_14816,N_14876);
and UO_685 (O_685,N_14833,N_14933);
xnor UO_686 (O_686,N_14815,N_14787);
nand UO_687 (O_687,N_14983,N_14853);
xor UO_688 (O_688,N_14933,N_14828);
xor UO_689 (O_689,N_14912,N_14877);
nor UO_690 (O_690,N_14857,N_14810);
nor UO_691 (O_691,N_14770,N_14812);
nand UO_692 (O_692,N_14773,N_14780);
nor UO_693 (O_693,N_14781,N_14875);
nor UO_694 (O_694,N_14781,N_14865);
nor UO_695 (O_695,N_14779,N_14912);
or UO_696 (O_696,N_14826,N_14927);
nor UO_697 (O_697,N_14759,N_14946);
or UO_698 (O_698,N_14939,N_14833);
or UO_699 (O_699,N_14994,N_14871);
or UO_700 (O_700,N_14827,N_14960);
nor UO_701 (O_701,N_14877,N_14921);
and UO_702 (O_702,N_14767,N_14990);
and UO_703 (O_703,N_14761,N_14843);
nor UO_704 (O_704,N_14755,N_14817);
or UO_705 (O_705,N_14815,N_14965);
nand UO_706 (O_706,N_14996,N_14930);
nor UO_707 (O_707,N_14757,N_14894);
and UO_708 (O_708,N_14790,N_14838);
or UO_709 (O_709,N_14949,N_14873);
nand UO_710 (O_710,N_14813,N_14928);
xor UO_711 (O_711,N_14825,N_14840);
nand UO_712 (O_712,N_14772,N_14791);
and UO_713 (O_713,N_14831,N_14962);
xnor UO_714 (O_714,N_14844,N_14865);
nand UO_715 (O_715,N_14751,N_14940);
xor UO_716 (O_716,N_14817,N_14787);
and UO_717 (O_717,N_14981,N_14983);
or UO_718 (O_718,N_14793,N_14787);
or UO_719 (O_719,N_14956,N_14853);
nor UO_720 (O_720,N_14871,N_14817);
nand UO_721 (O_721,N_14970,N_14888);
xor UO_722 (O_722,N_14823,N_14854);
nand UO_723 (O_723,N_14877,N_14794);
nand UO_724 (O_724,N_14775,N_14767);
nor UO_725 (O_725,N_14762,N_14864);
nor UO_726 (O_726,N_14968,N_14904);
nand UO_727 (O_727,N_14995,N_14912);
xor UO_728 (O_728,N_14841,N_14826);
or UO_729 (O_729,N_14785,N_14780);
or UO_730 (O_730,N_14911,N_14975);
nand UO_731 (O_731,N_14989,N_14777);
xnor UO_732 (O_732,N_14807,N_14868);
nor UO_733 (O_733,N_14815,N_14827);
nor UO_734 (O_734,N_14951,N_14934);
nor UO_735 (O_735,N_14760,N_14832);
or UO_736 (O_736,N_14911,N_14880);
or UO_737 (O_737,N_14778,N_14975);
nor UO_738 (O_738,N_14774,N_14883);
or UO_739 (O_739,N_14798,N_14970);
nor UO_740 (O_740,N_14833,N_14953);
nor UO_741 (O_741,N_14781,N_14965);
and UO_742 (O_742,N_14769,N_14856);
nor UO_743 (O_743,N_14944,N_14813);
and UO_744 (O_744,N_14750,N_14985);
or UO_745 (O_745,N_14763,N_14864);
and UO_746 (O_746,N_14872,N_14950);
xor UO_747 (O_747,N_14913,N_14970);
xnor UO_748 (O_748,N_14974,N_14851);
nand UO_749 (O_749,N_14857,N_14782);
and UO_750 (O_750,N_14937,N_14966);
and UO_751 (O_751,N_14872,N_14810);
or UO_752 (O_752,N_14876,N_14767);
nand UO_753 (O_753,N_14802,N_14772);
nand UO_754 (O_754,N_14949,N_14970);
xor UO_755 (O_755,N_14773,N_14829);
xnor UO_756 (O_756,N_14898,N_14956);
nand UO_757 (O_757,N_14777,N_14901);
nor UO_758 (O_758,N_14997,N_14992);
nand UO_759 (O_759,N_14995,N_14848);
and UO_760 (O_760,N_14998,N_14970);
xnor UO_761 (O_761,N_14937,N_14775);
xnor UO_762 (O_762,N_14768,N_14771);
xnor UO_763 (O_763,N_14801,N_14761);
nand UO_764 (O_764,N_14998,N_14862);
and UO_765 (O_765,N_14850,N_14989);
xnor UO_766 (O_766,N_14845,N_14776);
xor UO_767 (O_767,N_14968,N_14905);
nand UO_768 (O_768,N_14836,N_14769);
and UO_769 (O_769,N_14917,N_14812);
nor UO_770 (O_770,N_14757,N_14893);
nand UO_771 (O_771,N_14968,N_14847);
and UO_772 (O_772,N_14769,N_14917);
or UO_773 (O_773,N_14869,N_14892);
or UO_774 (O_774,N_14853,N_14959);
nand UO_775 (O_775,N_14791,N_14992);
nand UO_776 (O_776,N_14942,N_14980);
nand UO_777 (O_777,N_14857,N_14785);
nand UO_778 (O_778,N_14785,N_14800);
or UO_779 (O_779,N_14896,N_14949);
xor UO_780 (O_780,N_14989,N_14812);
nor UO_781 (O_781,N_14781,N_14891);
or UO_782 (O_782,N_14824,N_14820);
or UO_783 (O_783,N_14973,N_14867);
and UO_784 (O_784,N_14845,N_14885);
xnor UO_785 (O_785,N_14962,N_14927);
xor UO_786 (O_786,N_14838,N_14955);
or UO_787 (O_787,N_14924,N_14995);
nand UO_788 (O_788,N_14938,N_14831);
or UO_789 (O_789,N_14933,N_14787);
nand UO_790 (O_790,N_14897,N_14866);
xor UO_791 (O_791,N_14909,N_14773);
xnor UO_792 (O_792,N_14775,N_14951);
nand UO_793 (O_793,N_14759,N_14776);
and UO_794 (O_794,N_14790,N_14754);
and UO_795 (O_795,N_14797,N_14779);
or UO_796 (O_796,N_14996,N_14851);
and UO_797 (O_797,N_14836,N_14941);
nand UO_798 (O_798,N_14921,N_14942);
and UO_799 (O_799,N_14787,N_14908);
and UO_800 (O_800,N_14947,N_14912);
and UO_801 (O_801,N_14882,N_14828);
xor UO_802 (O_802,N_14937,N_14955);
xor UO_803 (O_803,N_14976,N_14968);
xnor UO_804 (O_804,N_14984,N_14779);
nor UO_805 (O_805,N_14926,N_14855);
and UO_806 (O_806,N_14830,N_14883);
nand UO_807 (O_807,N_14797,N_14935);
nand UO_808 (O_808,N_14813,N_14880);
and UO_809 (O_809,N_14785,N_14940);
or UO_810 (O_810,N_14975,N_14923);
xnor UO_811 (O_811,N_14957,N_14974);
and UO_812 (O_812,N_14912,N_14894);
xnor UO_813 (O_813,N_14905,N_14774);
xnor UO_814 (O_814,N_14973,N_14996);
xnor UO_815 (O_815,N_14778,N_14943);
nand UO_816 (O_816,N_14988,N_14794);
or UO_817 (O_817,N_14976,N_14924);
or UO_818 (O_818,N_14875,N_14784);
xor UO_819 (O_819,N_14920,N_14917);
xor UO_820 (O_820,N_14797,N_14917);
and UO_821 (O_821,N_14968,N_14804);
nand UO_822 (O_822,N_14989,N_14828);
xnor UO_823 (O_823,N_14945,N_14843);
nor UO_824 (O_824,N_14955,N_14832);
xor UO_825 (O_825,N_14831,N_14915);
nor UO_826 (O_826,N_14942,N_14789);
xnor UO_827 (O_827,N_14957,N_14864);
nand UO_828 (O_828,N_14758,N_14888);
or UO_829 (O_829,N_14897,N_14807);
nor UO_830 (O_830,N_14935,N_14969);
nor UO_831 (O_831,N_14843,N_14814);
xnor UO_832 (O_832,N_14967,N_14786);
nor UO_833 (O_833,N_14756,N_14820);
and UO_834 (O_834,N_14831,N_14868);
or UO_835 (O_835,N_14821,N_14963);
nor UO_836 (O_836,N_14845,N_14852);
and UO_837 (O_837,N_14924,N_14753);
nor UO_838 (O_838,N_14979,N_14872);
nand UO_839 (O_839,N_14993,N_14880);
xnor UO_840 (O_840,N_14771,N_14987);
and UO_841 (O_841,N_14913,N_14868);
nor UO_842 (O_842,N_14982,N_14995);
or UO_843 (O_843,N_14811,N_14845);
nor UO_844 (O_844,N_14814,N_14846);
or UO_845 (O_845,N_14840,N_14794);
nor UO_846 (O_846,N_14860,N_14931);
xnor UO_847 (O_847,N_14829,N_14838);
or UO_848 (O_848,N_14847,N_14851);
and UO_849 (O_849,N_14898,N_14818);
nand UO_850 (O_850,N_14924,N_14887);
and UO_851 (O_851,N_14989,N_14768);
nand UO_852 (O_852,N_14874,N_14764);
or UO_853 (O_853,N_14848,N_14993);
or UO_854 (O_854,N_14788,N_14975);
and UO_855 (O_855,N_14970,N_14867);
or UO_856 (O_856,N_14905,N_14891);
or UO_857 (O_857,N_14866,N_14948);
nor UO_858 (O_858,N_14789,N_14758);
nand UO_859 (O_859,N_14821,N_14913);
nor UO_860 (O_860,N_14888,N_14925);
xnor UO_861 (O_861,N_14929,N_14754);
nor UO_862 (O_862,N_14793,N_14812);
or UO_863 (O_863,N_14986,N_14835);
nand UO_864 (O_864,N_14900,N_14946);
nor UO_865 (O_865,N_14914,N_14772);
nand UO_866 (O_866,N_14984,N_14790);
or UO_867 (O_867,N_14751,N_14890);
or UO_868 (O_868,N_14783,N_14766);
and UO_869 (O_869,N_14790,N_14903);
xor UO_870 (O_870,N_14756,N_14841);
nor UO_871 (O_871,N_14764,N_14829);
xor UO_872 (O_872,N_14889,N_14776);
xor UO_873 (O_873,N_14875,N_14867);
and UO_874 (O_874,N_14952,N_14996);
xnor UO_875 (O_875,N_14944,N_14845);
nor UO_876 (O_876,N_14860,N_14966);
and UO_877 (O_877,N_14753,N_14800);
or UO_878 (O_878,N_14788,N_14972);
or UO_879 (O_879,N_14997,N_14928);
xnor UO_880 (O_880,N_14784,N_14816);
nand UO_881 (O_881,N_14765,N_14863);
or UO_882 (O_882,N_14963,N_14953);
xnor UO_883 (O_883,N_14898,N_14888);
or UO_884 (O_884,N_14910,N_14900);
nand UO_885 (O_885,N_14966,N_14865);
or UO_886 (O_886,N_14864,N_14892);
or UO_887 (O_887,N_14955,N_14944);
or UO_888 (O_888,N_14783,N_14900);
xor UO_889 (O_889,N_14833,N_14784);
xor UO_890 (O_890,N_14753,N_14755);
or UO_891 (O_891,N_14849,N_14883);
or UO_892 (O_892,N_14928,N_14858);
nand UO_893 (O_893,N_14889,N_14750);
or UO_894 (O_894,N_14986,N_14920);
nor UO_895 (O_895,N_14752,N_14942);
or UO_896 (O_896,N_14887,N_14824);
nor UO_897 (O_897,N_14804,N_14871);
nand UO_898 (O_898,N_14828,N_14934);
xnor UO_899 (O_899,N_14965,N_14805);
nor UO_900 (O_900,N_14816,N_14970);
xnor UO_901 (O_901,N_14779,N_14776);
and UO_902 (O_902,N_14791,N_14876);
or UO_903 (O_903,N_14892,N_14981);
and UO_904 (O_904,N_14775,N_14811);
or UO_905 (O_905,N_14922,N_14901);
nor UO_906 (O_906,N_14869,N_14825);
xor UO_907 (O_907,N_14941,N_14831);
xnor UO_908 (O_908,N_14898,N_14901);
nor UO_909 (O_909,N_14993,N_14810);
xnor UO_910 (O_910,N_14790,N_14967);
and UO_911 (O_911,N_14861,N_14869);
nand UO_912 (O_912,N_14815,N_14776);
and UO_913 (O_913,N_14818,N_14958);
nor UO_914 (O_914,N_14865,N_14921);
xor UO_915 (O_915,N_14763,N_14841);
or UO_916 (O_916,N_14822,N_14813);
and UO_917 (O_917,N_14772,N_14953);
nand UO_918 (O_918,N_14886,N_14768);
xnor UO_919 (O_919,N_14898,N_14895);
xor UO_920 (O_920,N_14914,N_14919);
nor UO_921 (O_921,N_14917,N_14999);
xnor UO_922 (O_922,N_14858,N_14878);
nor UO_923 (O_923,N_14959,N_14977);
xnor UO_924 (O_924,N_14957,N_14991);
nor UO_925 (O_925,N_14882,N_14896);
xnor UO_926 (O_926,N_14788,N_14764);
or UO_927 (O_927,N_14756,N_14998);
nand UO_928 (O_928,N_14835,N_14832);
and UO_929 (O_929,N_14890,N_14946);
or UO_930 (O_930,N_14878,N_14903);
and UO_931 (O_931,N_14929,N_14974);
nand UO_932 (O_932,N_14943,N_14788);
xnor UO_933 (O_933,N_14873,N_14804);
or UO_934 (O_934,N_14810,N_14912);
nand UO_935 (O_935,N_14821,N_14961);
and UO_936 (O_936,N_14825,N_14931);
nand UO_937 (O_937,N_14907,N_14971);
and UO_938 (O_938,N_14991,N_14797);
and UO_939 (O_939,N_14864,N_14921);
nand UO_940 (O_940,N_14853,N_14835);
nor UO_941 (O_941,N_14836,N_14855);
or UO_942 (O_942,N_14780,N_14752);
and UO_943 (O_943,N_14910,N_14964);
nand UO_944 (O_944,N_14891,N_14918);
or UO_945 (O_945,N_14770,N_14892);
nand UO_946 (O_946,N_14922,N_14876);
nor UO_947 (O_947,N_14997,N_14853);
and UO_948 (O_948,N_14822,N_14862);
xnor UO_949 (O_949,N_14900,N_14773);
and UO_950 (O_950,N_14888,N_14787);
nor UO_951 (O_951,N_14832,N_14762);
or UO_952 (O_952,N_14998,N_14850);
or UO_953 (O_953,N_14902,N_14913);
xnor UO_954 (O_954,N_14828,N_14992);
nor UO_955 (O_955,N_14902,N_14806);
xnor UO_956 (O_956,N_14780,N_14846);
xor UO_957 (O_957,N_14878,N_14989);
nor UO_958 (O_958,N_14834,N_14844);
or UO_959 (O_959,N_14953,N_14956);
nor UO_960 (O_960,N_14890,N_14847);
or UO_961 (O_961,N_14829,N_14945);
nand UO_962 (O_962,N_14928,N_14919);
nor UO_963 (O_963,N_14969,N_14852);
nor UO_964 (O_964,N_14846,N_14755);
nor UO_965 (O_965,N_14864,N_14769);
xor UO_966 (O_966,N_14783,N_14932);
xor UO_967 (O_967,N_14960,N_14885);
xor UO_968 (O_968,N_14988,N_14848);
xor UO_969 (O_969,N_14797,N_14826);
or UO_970 (O_970,N_14847,N_14809);
nor UO_971 (O_971,N_14937,N_14790);
and UO_972 (O_972,N_14757,N_14796);
and UO_973 (O_973,N_14981,N_14843);
and UO_974 (O_974,N_14767,N_14982);
nor UO_975 (O_975,N_14768,N_14806);
or UO_976 (O_976,N_14806,N_14852);
or UO_977 (O_977,N_14989,N_14860);
nor UO_978 (O_978,N_14759,N_14933);
nor UO_979 (O_979,N_14840,N_14775);
nor UO_980 (O_980,N_14794,N_14848);
nor UO_981 (O_981,N_14784,N_14815);
nor UO_982 (O_982,N_14977,N_14992);
xor UO_983 (O_983,N_14997,N_14882);
and UO_984 (O_984,N_14782,N_14827);
or UO_985 (O_985,N_14861,N_14975);
and UO_986 (O_986,N_14810,N_14914);
xor UO_987 (O_987,N_14861,N_14911);
xor UO_988 (O_988,N_14936,N_14779);
nand UO_989 (O_989,N_14813,N_14759);
and UO_990 (O_990,N_14818,N_14905);
or UO_991 (O_991,N_14785,N_14994);
or UO_992 (O_992,N_14829,N_14961);
xnor UO_993 (O_993,N_14756,N_14864);
and UO_994 (O_994,N_14802,N_14909);
nor UO_995 (O_995,N_14976,N_14782);
and UO_996 (O_996,N_14944,N_14927);
nand UO_997 (O_997,N_14760,N_14767);
or UO_998 (O_998,N_14969,N_14764);
or UO_999 (O_999,N_14906,N_14996);
nand UO_1000 (O_1000,N_14990,N_14978);
xor UO_1001 (O_1001,N_14982,N_14787);
nor UO_1002 (O_1002,N_14823,N_14814);
xnor UO_1003 (O_1003,N_14754,N_14857);
or UO_1004 (O_1004,N_14798,N_14878);
xor UO_1005 (O_1005,N_14953,N_14763);
or UO_1006 (O_1006,N_14829,N_14769);
nand UO_1007 (O_1007,N_14792,N_14952);
nor UO_1008 (O_1008,N_14791,N_14767);
nor UO_1009 (O_1009,N_14792,N_14922);
or UO_1010 (O_1010,N_14989,N_14826);
nor UO_1011 (O_1011,N_14775,N_14860);
or UO_1012 (O_1012,N_14821,N_14750);
or UO_1013 (O_1013,N_14984,N_14778);
and UO_1014 (O_1014,N_14850,N_14952);
nand UO_1015 (O_1015,N_14968,N_14845);
or UO_1016 (O_1016,N_14909,N_14794);
nand UO_1017 (O_1017,N_14882,N_14943);
nor UO_1018 (O_1018,N_14912,N_14969);
or UO_1019 (O_1019,N_14808,N_14758);
nor UO_1020 (O_1020,N_14811,N_14825);
nor UO_1021 (O_1021,N_14915,N_14824);
xor UO_1022 (O_1022,N_14997,N_14858);
or UO_1023 (O_1023,N_14827,N_14876);
and UO_1024 (O_1024,N_14950,N_14996);
or UO_1025 (O_1025,N_14977,N_14846);
or UO_1026 (O_1026,N_14980,N_14958);
xor UO_1027 (O_1027,N_14858,N_14939);
xnor UO_1028 (O_1028,N_14969,N_14895);
nand UO_1029 (O_1029,N_14923,N_14826);
or UO_1030 (O_1030,N_14815,N_14832);
and UO_1031 (O_1031,N_14986,N_14795);
or UO_1032 (O_1032,N_14970,N_14971);
and UO_1033 (O_1033,N_14906,N_14848);
and UO_1034 (O_1034,N_14853,N_14842);
nor UO_1035 (O_1035,N_14855,N_14844);
nand UO_1036 (O_1036,N_14812,N_14813);
nor UO_1037 (O_1037,N_14776,N_14822);
and UO_1038 (O_1038,N_14816,N_14926);
xor UO_1039 (O_1039,N_14916,N_14752);
nand UO_1040 (O_1040,N_14834,N_14919);
and UO_1041 (O_1041,N_14892,N_14955);
xor UO_1042 (O_1042,N_14793,N_14796);
nand UO_1043 (O_1043,N_14823,N_14923);
nor UO_1044 (O_1044,N_14933,N_14776);
xor UO_1045 (O_1045,N_14975,N_14949);
nor UO_1046 (O_1046,N_14826,N_14896);
and UO_1047 (O_1047,N_14978,N_14880);
nor UO_1048 (O_1048,N_14928,N_14876);
xnor UO_1049 (O_1049,N_14838,N_14844);
nor UO_1050 (O_1050,N_14782,N_14804);
xor UO_1051 (O_1051,N_14827,N_14831);
xor UO_1052 (O_1052,N_14786,N_14843);
nor UO_1053 (O_1053,N_14752,N_14995);
and UO_1054 (O_1054,N_14764,N_14934);
and UO_1055 (O_1055,N_14751,N_14822);
nor UO_1056 (O_1056,N_14786,N_14974);
nand UO_1057 (O_1057,N_14773,N_14966);
nand UO_1058 (O_1058,N_14759,N_14796);
xnor UO_1059 (O_1059,N_14889,N_14922);
or UO_1060 (O_1060,N_14951,N_14809);
and UO_1061 (O_1061,N_14954,N_14897);
or UO_1062 (O_1062,N_14776,N_14775);
nor UO_1063 (O_1063,N_14843,N_14844);
xor UO_1064 (O_1064,N_14917,N_14968);
and UO_1065 (O_1065,N_14820,N_14850);
or UO_1066 (O_1066,N_14930,N_14935);
nand UO_1067 (O_1067,N_14801,N_14998);
xnor UO_1068 (O_1068,N_14866,N_14785);
and UO_1069 (O_1069,N_14997,N_14970);
xor UO_1070 (O_1070,N_14978,N_14992);
nand UO_1071 (O_1071,N_14908,N_14780);
xor UO_1072 (O_1072,N_14915,N_14954);
or UO_1073 (O_1073,N_14858,N_14842);
xor UO_1074 (O_1074,N_14753,N_14882);
nand UO_1075 (O_1075,N_14991,N_14914);
or UO_1076 (O_1076,N_14782,N_14911);
or UO_1077 (O_1077,N_14779,N_14948);
nand UO_1078 (O_1078,N_14848,N_14921);
xor UO_1079 (O_1079,N_14936,N_14992);
xor UO_1080 (O_1080,N_14836,N_14906);
xor UO_1081 (O_1081,N_14915,N_14814);
nand UO_1082 (O_1082,N_14855,N_14837);
and UO_1083 (O_1083,N_14811,N_14829);
nor UO_1084 (O_1084,N_14777,N_14942);
and UO_1085 (O_1085,N_14827,N_14860);
nand UO_1086 (O_1086,N_14979,N_14882);
or UO_1087 (O_1087,N_14829,N_14821);
xnor UO_1088 (O_1088,N_14973,N_14917);
nand UO_1089 (O_1089,N_14856,N_14985);
xnor UO_1090 (O_1090,N_14760,N_14891);
nand UO_1091 (O_1091,N_14777,N_14878);
nand UO_1092 (O_1092,N_14758,N_14780);
xor UO_1093 (O_1093,N_14804,N_14764);
nand UO_1094 (O_1094,N_14898,N_14784);
nor UO_1095 (O_1095,N_14817,N_14932);
xnor UO_1096 (O_1096,N_14812,N_14935);
and UO_1097 (O_1097,N_14848,N_14768);
or UO_1098 (O_1098,N_14995,N_14778);
and UO_1099 (O_1099,N_14822,N_14899);
and UO_1100 (O_1100,N_14786,N_14792);
or UO_1101 (O_1101,N_14932,N_14807);
and UO_1102 (O_1102,N_14914,N_14886);
or UO_1103 (O_1103,N_14933,N_14832);
nor UO_1104 (O_1104,N_14809,N_14962);
and UO_1105 (O_1105,N_14788,N_14795);
or UO_1106 (O_1106,N_14790,N_14891);
or UO_1107 (O_1107,N_14913,N_14828);
and UO_1108 (O_1108,N_14982,N_14970);
and UO_1109 (O_1109,N_14805,N_14981);
nor UO_1110 (O_1110,N_14867,N_14988);
or UO_1111 (O_1111,N_14755,N_14993);
xor UO_1112 (O_1112,N_14959,N_14768);
xnor UO_1113 (O_1113,N_14962,N_14965);
and UO_1114 (O_1114,N_14985,N_14930);
and UO_1115 (O_1115,N_14885,N_14835);
xnor UO_1116 (O_1116,N_14751,N_14905);
or UO_1117 (O_1117,N_14878,N_14807);
nor UO_1118 (O_1118,N_14975,N_14819);
xor UO_1119 (O_1119,N_14881,N_14810);
and UO_1120 (O_1120,N_14954,N_14759);
and UO_1121 (O_1121,N_14779,N_14802);
or UO_1122 (O_1122,N_14984,N_14835);
or UO_1123 (O_1123,N_14854,N_14808);
xor UO_1124 (O_1124,N_14997,N_14822);
and UO_1125 (O_1125,N_14973,N_14927);
and UO_1126 (O_1126,N_14781,N_14761);
and UO_1127 (O_1127,N_14773,N_14845);
nor UO_1128 (O_1128,N_14901,N_14928);
nor UO_1129 (O_1129,N_14761,N_14977);
and UO_1130 (O_1130,N_14888,N_14838);
xor UO_1131 (O_1131,N_14998,N_14868);
and UO_1132 (O_1132,N_14947,N_14786);
or UO_1133 (O_1133,N_14899,N_14990);
nand UO_1134 (O_1134,N_14807,N_14872);
and UO_1135 (O_1135,N_14792,N_14911);
nand UO_1136 (O_1136,N_14960,N_14952);
or UO_1137 (O_1137,N_14787,N_14871);
or UO_1138 (O_1138,N_14770,N_14904);
xnor UO_1139 (O_1139,N_14893,N_14961);
xor UO_1140 (O_1140,N_14856,N_14819);
nor UO_1141 (O_1141,N_14841,N_14773);
nor UO_1142 (O_1142,N_14796,N_14775);
and UO_1143 (O_1143,N_14788,N_14941);
nand UO_1144 (O_1144,N_14799,N_14750);
nor UO_1145 (O_1145,N_14993,N_14753);
or UO_1146 (O_1146,N_14779,N_14968);
xor UO_1147 (O_1147,N_14779,N_14751);
nand UO_1148 (O_1148,N_14881,N_14960);
xnor UO_1149 (O_1149,N_14814,N_14833);
xnor UO_1150 (O_1150,N_14944,N_14794);
and UO_1151 (O_1151,N_14756,N_14795);
and UO_1152 (O_1152,N_14903,N_14902);
nand UO_1153 (O_1153,N_14992,N_14884);
and UO_1154 (O_1154,N_14837,N_14762);
xnor UO_1155 (O_1155,N_14915,N_14880);
xor UO_1156 (O_1156,N_14962,N_14807);
xnor UO_1157 (O_1157,N_14894,N_14760);
nand UO_1158 (O_1158,N_14858,N_14832);
or UO_1159 (O_1159,N_14944,N_14856);
xor UO_1160 (O_1160,N_14999,N_14912);
and UO_1161 (O_1161,N_14812,N_14942);
nand UO_1162 (O_1162,N_14830,N_14936);
and UO_1163 (O_1163,N_14965,N_14963);
or UO_1164 (O_1164,N_14829,N_14803);
or UO_1165 (O_1165,N_14880,N_14823);
nor UO_1166 (O_1166,N_14792,N_14881);
nor UO_1167 (O_1167,N_14886,N_14958);
nand UO_1168 (O_1168,N_14862,N_14771);
nor UO_1169 (O_1169,N_14754,N_14943);
and UO_1170 (O_1170,N_14793,N_14833);
or UO_1171 (O_1171,N_14999,N_14991);
or UO_1172 (O_1172,N_14750,N_14942);
nor UO_1173 (O_1173,N_14765,N_14763);
and UO_1174 (O_1174,N_14954,N_14999);
xnor UO_1175 (O_1175,N_14881,N_14874);
or UO_1176 (O_1176,N_14943,N_14815);
nor UO_1177 (O_1177,N_14791,N_14893);
nand UO_1178 (O_1178,N_14975,N_14888);
and UO_1179 (O_1179,N_14979,N_14919);
and UO_1180 (O_1180,N_14774,N_14768);
nand UO_1181 (O_1181,N_14846,N_14975);
and UO_1182 (O_1182,N_14813,N_14858);
nand UO_1183 (O_1183,N_14927,N_14845);
xor UO_1184 (O_1184,N_14930,N_14956);
nand UO_1185 (O_1185,N_14775,N_14867);
nor UO_1186 (O_1186,N_14898,N_14996);
and UO_1187 (O_1187,N_14950,N_14851);
or UO_1188 (O_1188,N_14916,N_14804);
and UO_1189 (O_1189,N_14904,N_14967);
nand UO_1190 (O_1190,N_14882,N_14942);
or UO_1191 (O_1191,N_14889,N_14812);
xor UO_1192 (O_1192,N_14841,N_14949);
and UO_1193 (O_1193,N_14767,N_14801);
nor UO_1194 (O_1194,N_14845,N_14750);
xor UO_1195 (O_1195,N_14943,N_14791);
nor UO_1196 (O_1196,N_14990,N_14960);
or UO_1197 (O_1197,N_14906,N_14988);
and UO_1198 (O_1198,N_14774,N_14772);
and UO_1199 (O_1199,N_14978,N_14976);
nor UO_1200 (O_1200,N_14769,N_14817);
and UO_1201 (O_1201,N_14977,N_14754);
and UO_1202 (O_1202,N_14915,N_14784);
or UO_1203 (O_1203,N_14895,N_14897);
nor UO_1204 (O_1204,N_14969,N_14920);
nand UO_1205 (O_1205,N_14894,N_14888);
and UO_1206 (O_1206,N_14915,N_14850);
xnor UO_1207 (O_1207,N_14812,N_14953);
xor UO_1208 (O_1208,N_14971,N_14769);
and UO_1209 (O_1209,N_14996,N_14767);
and UO_1210 (O_1210,N_14814,N_14756);
or UO_1211 (O_1211,N_14872,N_14825);
and UO_1212 (O_1212,N_14822,N_14864);
nor UO_1213 (O_1213,N_14906,N_14983);
xor UO_1214 (O_1214,N_14991,N_14774);
nand UO_1215 (O_1215,N_14991,N_14824);
nor UO_1216 (O_1216,N_14857,N_14935);
xor UO_1217 (O_1217,N_14939,N_14978);
and UO_1218 (O_1218,N_14817,N_14877);
nor UO_1219 (O_1219,N_14990,N_14892);
xor UO_1220 (O_1220,N_14930,N_14905);
nand UO_1221 (O_1221,N_14853,N_14803);
xnor UO_1222 (O_1222,N_14804,N_14974);
or UO_1223 (O_1223,N_14780,N_14912);
nor UO_1224 (O_1224,N_14946,N_14913);
or UO_1225 (O_1225,N_14996,N_14763);
or UO_1226 (O_1226,N_14928,N_14832);
xor UO_1227 (O_1227,N_14844,N_14949);
nor UO_1228 (O_1228,N_14943,N_14845);
nor UO_1229 (O_1229,N_14899,N_14820);
or UO_1230 (O_1230,N_14836,N_14879);
and UO_1231 (O_1231,N_14810,N_14957);
xnor UO_1232 (O_1232,N_14859,N_14973);
nand UO_1233 (O_1233,N_14811,N_14972);
nand UO_1234 (O_1234,N_14863,N_14917);
xor UO_1235 (O_1235,N_14804,N_14938);
nor UO_1236 (O_1236,N_14871,N_14830);
and UO_1237 (O_1237,N_14945,N_14788);
nor UO_1238 (O_1238,N_14760,N_14919);
xnor UO_1239 (O_1239,N_14918,N_14965);
xor UO_1240 (O_1240,N_14987,N_14944);
and UO_1241 (O_1241,N_14820,N_14788);
nand UO_1242 (O_1242,N_14889,N_14877);
or UO_1243 (O_1243,N_14953,N_14858);
and UO_1244 (O_1244,N_14801,N_14920);
or UO_1245 (O_1245,N_14775,N_14920);
nand UO_1246 (O_1246,N_14946,N_14779);
xor UO_1247 (O_1247,N_14883,N_14939);
or UO_1248 (O_1248,N_14770,N_14847);
and UO_1249 (O_1249,N_14912,N_14965);
nand UO_1250 (O_1250,N_14891,N_14761);
and UO_1251 (O_1251,N_14963,N_14958);
or UO_1252 (O_1252,N_14854,N_14929);
and UO_1253 (O_1253,N_14754,N_14807);
nand UO_1254 (O_1254,N_14991,N_14924);
xnor UO_1255 (O_1255,N_14797,N_14807);
xor UO_1256 (O_1256,N_14964,N_14901);
xor UO_1257 (O_1257,N_14956,N_14875);
xor UO_1258 (O_1258,N_14847,N_14850);
or UO_1259 (O_1259,N_14801,N_14787);
or UO_1260 (O_1260,N_14788,N_14903);
or UO_1261 (O_1261,N_14832,N_14795);
nor UO_1262 (O_1262,N_14896,N_14965);
xor UO_1263 (O_1263,N_14911,N_14964);
nand UO_1264 (O_1264,N_14830,N_14764);
xor UO_1265 (O_1265,N_14833,N_14758);
xnor UO_1266 (O_1266,N_14844,N_14811);
nand UO_1267 (O_1267,N_14962,N_14979);
nor UO_1268 (O_1268,N_14800,N_14886);
xnor UO_1269 (O_1269,N_14830,N_14794);
nor UO_1270 (O_1270,N_14948,N_14922);
and UO_1271 (O_1271,N_14856,N_14942);
or UO_1272 (O_1272,N_14983,N_14791);
nand UO_1273 (O_1273,N_14966,N_14813);
and UO_1274 (O_1274,N_14909,N_14799);
nor UO_1275 (O_1275,N_14788,N_14924);
and UO_1276 (O_1276,N_14920,N_14885);
nand UO_1277 (O_1277,N_14841,N_14786);
and UO_1278 (O_1278,N_14845,N_14808);
and UO_1279 (O_1279,N_14883,N_14816);
nor UO_1280 (O_1280,N_14859,N_14804);
or UO_1281 (O_1281,N_14779,N_14895);
nor UO_1282 (O_1282,N_14956,N_14999);
xnor UO_1283 (O_1283,N_14869,N_14905);
and UO_1284 (O_1284,N_14913,N_14871);
xnor UO_1285 (O_1285,N_14992,N_14829);
nand UO_1286 (O_1286,N_14767,N_14858);
nand UO_1287 (O_1287,N_14911,N_14860);
nand UO_1288 (O_1288,N_14948,N_14842);
nor UO_1289 (O_1289,N_14786,N_14773);
nor UO_1290 (O_1290,N_14801,N_14986);
nand UO_1291 (O_1291,N_14943,N_14776);
and UO_1292 (O_1292,N_14963,N_14887);
nand UO_1293 (O_1293,N_14887,N_14817);
or UO_1294 (O_1294,N_14952,N_14918);
nand UO_1295 (O_1295,N_14758,N_14960);
xor UO_1296 (O_1296,N_14872,N_14770);
or UO_1297 (O_1297,N_14872,N_14886);
or UO_1298 (O_1298,N_14751,N_14864);
nor UO_1299 (O_1299,N_14834,N_14896);
xor UO_1300 (O_1300,N_14956,N_14944);
nand UO_1301 (O_1301,N_14912,N_14751);
xnor UO_1302 (O_1302,N_14768,N_14987);
and UO_1303 (O_1303,N_14840,N_14851);
xnor UO_1304 (O_1304,N_14998,N_14946);
or UO_1305 (O_1305,N_14955,N_14799);
nand UO_1306 (O_1306,N_14971,N_14838);
xnor UO_1307 (O_1307,N_14992,N_14881);
xor UO_1308 (O_1308,N_14786,N_14774);
xnor UO_1309 (O_1309,N_14908,N_14875);
xnor UO_1310 (O_1310,N_14953,N_14880);
xor UO_1311 (O_1311,N_14793,N_14890);
and UO_1312 (O_1312,N_14791,N_14823);
nand UO_1313 (O_1313,N_14934,N_14975);
and UO_1314 (O_1314,N_14846,N_14771);
and UO_1315 (O_1315,N_14942,N_14787);
or UO_1316 (O_1316,N_14871,N_14791);
nor UO_1317 (O_1317,N_14878,N_14869);
and UO_1318 (O_1318,N_14864,N_14905);
nor UO_1319 (O_1319,N_14878,N_14788);
xor UO_1320 (O_1320,N_14912,N_14813);
xor UO_1321 (O_1321,N_14911,N_14919);
xnor UO_1322 (O_1322,N_14810,N_14803);
xor UO_1323 (O_1323,N_14785,N_14893);
or UO_1324 (O_1324,N_14914,N_14996);
and UO_1325 (O_1325,N_14783,N_14796);
and UO_1326 (O_1326,N_14944,N_14963);
nand UO_1327 (O_1327,N_14853,N_14943);
and UO_1328 (O_1328,N_14812,N_14950);
xor UO_1329 (O_1329,N_14995,N_14827);
nand UO_1330 (O_1330,N_14809,N_14792);
and UO_1331 (O_1331,N_14830,N_14875);
or UO_1332 (O_1332,N_14777,N_14790);
nor UO_1333 (O_1333,N_14926,N_14911);
nand UO_1334 (O_1334,N_14800,N_14983);
xnor UO_1335 (O_1335,N_14971,N_14869);
and UO_1336 (O_1336,N_14847,N_14991);
nor UO_1337 (O_1337,N_14921,N_14867);
nand UO_1338 (O_1338,N_14761,N_14939);
and UO_1339 (O_1339,N_14811,N_14940);
nor UO_1340 (O_1340,N_14792,N_14781);
and UO_1341 (O_1341,N_14934,N_14778);
nand UO_1342 (O_1342,N_14907,N_14851);
nand UO_1343 (O_1343,N_14798,N_14866);
xnor UO_1344 (O_1344,N_14955,N_14771);
nand UO_1345 (O_1345,N_14804,N_14814);
nand UO_1346 (O_1346,N_14842,N_14914);
or UO_1347 (O_1347,N_14873,N_14953);
nor UO_1348 (O_1348,N_14811,N_14870);
xor UO_1349 (O_1349,N_14956,N_14880);
xor UO_1350 (O_1350,N_14860,N_14936);
and UO_1351 (O_1351,N_14800,N_14980);
nor UO_1352 (O_1352,N_14991,N_14751);
and UO_1353 (O_1353,N_14896,N_14857);
nor UO_1354 (O_1354,N_14757,N_14914);
nor UO_1355 (O_1355,N_14871,N_14880);
and UO_1356 (O_1356,N_14821,N_14984);
or UO_1357 (O_1357,N_14821,N_14928);
xor UO_1358 (O_1358,N_14766,N_14950);
xnor UO_1359 (O_1359,N_14970,N_14822);
nand UO_1360 (O_1360,N_14957,N_14963);
or UO_1361 (O_1361,N_14979,N_14978);
xor UO_1362 (O_1362,N_14964,N_14750);
nand UO_1363 (O_1363,N_14898,N_14859);
nor UO_1364 (O_1364,N_14784,N_14942);
or UO_1365 (O_1365,N_14916,N_14859);
or UO_1366 (O_1366,N_14991,N_14899);
nor UO_1367 (O_1367,N_14959,N_14883);
xnor UO_1368 (O_1368,N_14776,N_14816);
nand UO_1369 (O_1369,N_14882,N_14792);
xor UO_1370 (O_1370,N_14855,N_14856);
and UO_1371 (O_1371,N_14815,N_14973);
and UO_1372 (O_1372,N_14809,N_14894);
or UO_1373 (O_1373,N_14797,N_14874);
xnor UO_1374 (O_1374,N_14818,N_14981);
nand UO_1375 (O_1375,N_14871,N_14854);
xor UO_1376 (O_1376,N_14947,N_14784);
nand UO_1377 (O_1377,N_14967,N_14997);
xnor UO_1378 (O_1378,N_14990,N_14873);
or UO_1379 (O_1379,N_14926,N_14985);
nand UO_1380 (O_1380,N_14970,N_14906);
and UO_1381 (O_1381,N_14826,N_14986);
or UO_1382 (O_1382,N_14941,N_14923);
or UO_1383 (O_1383,N_14987,N_14932);
and UO_1384 (O_1384,N_14876,N_14984);
nand UO_1385 (O_1385,N_14803,N_14970);
xnor UO_1386 (O_1386,N_14797,N_14800);
and UO_1387 (O_1387,N_14943,N_14800);
nand UO_1388 (O_1388,N_14865,N_14964);
or UO_1389 (O_1389,N_14799,N_14864);
or UO_1390 (O_1390,N_14958,N_14938);
nor UO_1391 (O_1391,N_14792,N_14943);
or UO_1392 (O_1392,N_14959,N_14961);
nand UO_1393 (O_1393,N_14868,N_14944);
nand UO_1394 (O_1394,N_14877,N_14760);
nand UO_1395 (O_1395,N_14752,N_14927);
xor UO_1396 (O_1396,N_14851,N_14966);
and UO_1397 (O_1397,N_14761,N_14752);
nor UO_1398 (O_1398,N_14844,N_14754);
nor UO_1399 (O_1399,N_14924,N_14965);
or UO_1400 (O_1400,N_14970,N_14915);
nor UO_1401 (O_1401,N_14820,N_14792);
or UO_1402 (O_1402,N_14828,N_14779);
nand UO_1403 (O_1403,N_14840,N_14836);
or UO_1404 (O_1404,N_14821,N_14752);
xnor UO_1405 (O_1405,N_14873,N_14937);
and UO_1406 (O_1406,N_14887,N_14976);
nor UO_1407 (O_1407,N_14976,N_14863);
xor UO_1408 (O_1408,N_14803,N_14826);
and UO_1409 (O_1409,N_14799,N_14808);
and UO_1410 (O_1410,N_14775,N_14895);
and UO_1411 (O_1411,N_14834,N_14907);
nor UO_1412 (O_1412,N_14969,N_14775);
nor UO_1413 (O_1413,N_14850,N_14843);
nand UO_1414 (O_1414,N_14989,N_14956);
or UO_1415 (O_1415,N_14873,N_14840);
and UO_1416 (O_1416,N_14777,N_14912);
nand UO_1417 (O_1417,N_14832,N_14863);
and UO_1418 (O_1418,N_14994,N_14831);
nor UO_1419 (O_1419,N_14931,N_14982);
or UO_1420 (O_1420,N_14889,N_14802);
or UO_1421 (O_1421,N_14990,N_14868);
and UO_1422 (O_1422,N_14997,N_14922);
or UO_1423 (O_1423,N_14768,N_14799);
xnor UO_1424 (O_1424,N_14963,N_14961);
and UO_1425 (O_1425,N_14846,N_14981);
nor UO_1426 (O_1426,N_14937,N_14884);
and UO_1427 (O_1427,N_14809,N_14875);
nor UO_1428 (O_1428,N_14774,N_14987);
nand UO_1429 (O_1429,N_14954,N_14766);
or UO_1430 (O_1430,N_14753,N_14793);
and UO_1431 (O_1431,N_14753,N_14816);
xor UO_1432 (O_1432,N_14984,N_14945);
and UO_1433 (O_1433,N_14816,N_14830);
xor UO_1434 (O_1434,N_14881,N_14860);
xor UO_1435 (O_1435,N_14998,N_14958);
nand UO_1436 (O_1436,N_14898,N_14906);
nand UO_1437 (O_1437,N_14975,N_14860);
nor UO_1438 (O_1438,N_14997,N_14780);
nor UO_1439 (O_1439,N_14932,N_14831);
nor UO_1440 (O_1440,N_14811,N_14903);
and UO_1441 (O_1441,N_14821,N_14838);
xor UO_1442 (O_1442,N_14793,N_14774);
nor UO_1443 (O_1443,N_14934,N_14972);
or UO_1444 (O_1444,N_14882,N_14796);
nor UO_1445 (O_1445,N_14857,N_14837);
nor UO_1446 (O_1446,N_14863,N_14845);
or UO_1447 (O_1447,N_14889,N_14927);
or UO_1448 (O_1448,N_14806,N_14757);
xnor UO_1449 (O_1449,N_14799,N_14896);
xor UO_1450 (O_1450,N_14903,N_14817);
or UO_1451 (O_1451,N_14848,N_14847);
or UO_1452 (O_1452,N_14995,N_14889);
nor UO_1453 (O_1453,N_14834,N_14995);
nor UO_1454 (O_1454,N_14852,N_14971);
nand UO_1455 (O_1455,N_14850,N_14974);
nor UO_1456 (O_1456,N_14852,N_14759);
xnor UO_1457 (O_1457,N_14907,N_14883);
xnor UO_1458 (O_1458,N_14752,N_14922);
nand UO_1459 (O_1459,N_14909,N_14948);
nand UO_1460 (O_1460,N_14846,N_14918);
nand UO_1461 (O_1461,N_14978,N_14815);
xor UO_1462 (O_1462,N_14776,N_14975);
xor UO_1463 (O_1463,N_14985,N_14773);
nand UO_1464 (O_1464,N_14963,N_14860);
or UO_1465 (O_1465,N_14846,N_14791);
nor UO_1466 (O_1466,N_14786,N_14782);
nor UO_1467 (O_1467,N_14911,N_14805);
and UO_1468 (O_1468,N_14881,N_14764);
xor UO_1469 (O_1469,N_14856,N_14928);
xor UO_1470 (O_1470,N_14922,N_14757);
nand UO_1471 (O_1471,N_14857,N_14996);
xor UO_1472 (O_1472,N_14853,N_14985);
nor UO_1473 (O_1473,N_14990,N_14878);
nand UO_1474 (O_1474,N_14822,N_14779);
or UO_1475 (O_1475,N_14806,N_14904);
or UO_1476 (O_1476,N_14951,N_14816);
xnor UO_1477 (O_1477,N_14967,N_14880);
nor UO_1478 (O_1478,N_14839,N_14760);
or UO_1479 (O_1479,N_14764,N_14961);
and UO_1480 (O_1480,N_14926,N_14819);
and UO_1481 (O_1481,N_14844,N_14921);
nor UO_1482 (O_1482,N_14990,N_14884);
nor UO_1483 (O_1483,N_14904,N_14898);
xnor UO_1484 (O_1484,N_14833,N_14901);
and UO_1485 (O_1485,N_14912,N_14812);
nand UO_1486 (O_1486,N_14896,N_14994);
nand UO_1487 (O_1487,N_14919,N_14931);
xnor UO_1488 (O_1488,N_14908,N_14833);
or UO_1489 (O_1489,N_14954,N_14818);
xnor UO_1490 (O_1490,N_14981,N_14877);
nor UO_1491 (O_1491,N_14928,N_14810);
nand UO_1492 (O_1492,N_14784,N_14804);
nand UO_1493 (O_1493,N_14895,N_14980);
and UO_1494 (O_1494,N_14751,N_14762);
nor UO_1495 (O_1495,N_14795,N_14791);
and UO_1496 (O_1496,N_14880,N_14857);
nor UO_1497 (O_1497,N_14892,N_14914);
or UO_1498 (O_1498,N_14847,N_14751);
or UO_1499 (O_1499,N_14965,N_14937);
nor UO_1500 (O_1500,N_14887,N_14996);
or UO_1501 (O_1501,N_14953,N_14816);
xnor UO_1502 (O_1502,N_14913,N_14762);
nand UO_1503 (O_1503,N_14887,N_14877);
and UO_1504 (O_1504,N_14853,N_14765);
nand UO_1505 (O_1505,N_14752,N_14997);
nor UO_1506 (O_1506,N_14871,N_14921);
and UO_1507 (O_1507,N_14985,N_14774);
and UO_1508 (O_1508,N_14959,N_14819);
xor UO_1509 (O_1509,N_14760,N_14810);
and UO_1510 (O_1510,N_14796,N_14917);
nand UO_1511 (O_1511,N_14930,N_14875);
nand UO_1512 (O_1512,N_14841,N_14996);
or UO_1513 (O_1513,N_14981,N_14886);
nor UO_1514 (O_1514,N_14823,N_14914);
or UO_1515 (O_1515,N_14982,N_14987);
xnor UO_1516 (O_1516,N_14963,N_14999);
or UO_1517 (O_1517,N_14887,N_14965);
nor UO_1518 (O_1518,N_14985,N_14821);
nor UO_1519 (O_1519,N_14804,N_14943);
or UO_1520 (O_1520,N_14792,N_14779);
nor UO_1521 (O_1521,N_14894,N_14761);
xor UO_1522 (O_1522,N_14947,N_14929);
nor UO_1523 (O_1523,N_14750,N_14967);
xor UO_1524 (O_1524,N_14993,N_14921);
xor UO_1525 (O_1525,N_14951,N_14822);
and UO_1526 (O_1526,N_14957,N_14977);
and UO_1527 (O_1527,N_14754,N_14934);
or UO_1528 (O_1528,N_14772,N_14763);
or UO_1529 (O_1529,N_14831,N_14770);
nand UO_1530 (O_1530,N_14853,N_14850);
xor UO_1531 (O_1531,N_14945,N_14825);
or UO_1532 (O_1532,N_14871,N_14857);
nand UO_1533 (O_1533,N_14879,N_14841);
nand UO_1534 (O_1534,N_14886,N_14772);
xor UO_1535 (O_1535,N_14958,N_14995);
nand UO_1536 (O_1536,N_14894,N_14834);
nor UO_1537 (O_1537,N_14828,N_14773);
xnor UO_1538 (O_1538,N_14765,N_14959);
nor UO_1539 (O_1539,N_14910,N_14770);
nand UO_1540 (O_1540,N_14859,N_14765);
nand UO_1541 (O_1541,N_14832,N_14806);
or UO_1542 (O_1542,N_14904,N_14856);
xor UO_1543 (O_1543,N_14972,N_14759);
xor UO_1544 (O_1544,N_14903,N_14818);
xnor UO_1545 (O_1545,N_14778,N_14830);
or UO_1546 (O_1546,N_14767,N_14807);
or UO_1547 (O_1547,N_14970,N_14821);
or UO_1548 (O_1548,N_14912,N_14910);
and UO_1549 (O_1549,N_14811,N_14760);
or UO_1550 (O_1550,N_14775,N_14986);
nand UO_1551 (O_1551,N_14905,N_14932);
and UO_1552 (O_1552,N_14933,N_14796);
nand UO_1553 (O_1553,N_14902,N_14932);
and UO_1554 (O_1554,N_14765,N_14964);
xor UO_1555 (O_1555,N_14923,N_14866);
nand UO_1556 (O_1556,N_14929,N_14828);
or UO_1557 (O_1557,N_14945,N_14787);
xnor UO_1558 (O_1558,N_14986,N_14831);
nand UO_1559 (O_1559,N_14848,N_14895);
or UO_1560 (O_1560,N_14921,N_14938);
xnor UO_1561 (O_1561,N_14984,N_14924);
or UO_1562 (O_1562,N_14916,N_14845);
and UO_1563 (O_1563,N_14896,N_14797);
xnor UO_1564 (O_1564,N_14999,N_14967);
or UO_1565 (O_1565,N_14764,N_14760);
xnor UO_1566 (O_1566,N_14934,N_14961);
xnor UO_1567 (O_1567,N_14802,N_14997);
or UO_1568 (O_1568,N_14767,N_14824);
or UO_1569 (O_1569,N_14953,N_14843);
nor UO_1570 (O_1570,N_14963,N_14844);
nor UO_1571 (O_1571,N_14762,N_14794);
nor UO_1572 (O_1572,N_14823,N_14983);
nand UO_1573 (O_1573,N_14928,N_14872);
nand UO_1574 (O_1574,N_14944,N_14788);
nor UO_1575 (O_1575,N_14772,N_14778);
or UO_1576 (O_1576,N_14819,N_14768);
nor UO_1577 (O_1577,N_14826,N_14974);
xnor UO_1578 (O_1578,N_14983,N_14926);
nand UO_1579 (O_1579,N_14919,N_14970);
or UO_1580 (O_1580,N_14934,N_14879);
and UO_1581 (O_1581,N_14867,N_14756);
and UO_1582 (O_1582,N_14810,N_14926);
nor UO_1583 (O_1583,N_14972,N_14957);
or UO_1584 (O_1584,N_14755,N_14964);
nand UO_1585 (O_1585,N_14907,N_14788);
and UO_1586 (O_1586,N_14890,N_14904);
nor UO_1587 (O_1587,N_14939,N_14909);
xor UO_1588 (O_1588,N_14830,N_14801);
xnor UO_1589 (O_1589,N_14854,N_14933);
and UO_1590 (O_1590,N_14857,N_14906);
or UO_1591 (O_1591,N_14965,N_14810);
or UO_1592 (O_1592,N_14784,N_14884);
or UO_1593 (O_1593,N_14849,N_14841);
xnor UO_1594 (O_1594,N_14832,N_14807);
and UO_1595 (O_1595,N_14835,N_14759);
nor UO_1596 (O_1596,N_14895,N_14750);
or UO_1597 (O_1597,N_14976,N_14898);
xnor UO_1598 (O_1598,N_14787,N_14996);
and UO_1599 (O_1599,N_14993,N_14803);
and UO_1600 (O_1600,N_14940,N_14892);
nand UO_1601 (O_1601,N_14937,N_14857);
or UO_1602 (O_1602,N_14928,N_14841);
nand UO_1603 (O_1603,N_14870,N_14768);
nor UO_1604 (O_1604,N_14768,N_14822);
nand UO_1605 (O_1605,N_14922,N_14851);
and UO_1606 (O_1606,N_14970,N_14890);
nor UO_1607 (O_1607,N_14926,N_14878);
and UO_1608 (O_1608,N_14907,N_14779);
nor UO_1609 (O_1609,N_14939,N_14807);
or UO_1610 (O_1610,N_14866,N_14860);
and UO_1611 (O_1611,N_14849,N_14963);
and UO_1612 (O_1612,N_14868,N_14976);
or UO_1613 (O_1613,N_14860,N_14782);
nor UO_1614 (O_1614,N_14911,N_14952);
or UO_1615 (O_1615,N_14971,N_14980);
nor UO_1616 (O_1616,N_14940,N_14956);
xor UO_1617 (O_1617,N_14827,N_14948);
and UO_1618 (O_1618,N_14896,N_14974);
xnor UO_1619 (O_1619,N_14982,N_14941);
nor UO_1620 (O_1620,N_14980,N_14968);
nor UO_1621 (O_1621,N_14946,N_14801);
and UO_1622 (O_1622,N_14977,N_14797);
xnor UO_1623 (O_1623,N_14910,N_14959);
nand UO_1624 (O_1624,N_14776,N_14915);
nor UO_1625 (O_1625,N_14791,N_14991);
nor UO_1626 (O_1626,N_14791,N_14976);
xnor UO_1627 (O_1627,N_14962,N_14830);
or UO_1628 (O_1628,N_14839,N_14975);
and UO_1629 (O_1629,N_14910,N_14999);
and UO_1630 (O_1630,N_14984,N_14985);
or UO_1631 (O_1631,N_14936,N_14783);
nand UO_1632 (O_1632,N_14988,N_14996);
and UO_1633 (O_1633,N_14831,N_14803);
or UO_1634 (O_1634,N_14818,N_14895);
nand UO_1635 (O_1635,N_14763,N_14817);
nand UO_1636 (O_1636,N_14954,N_14924);
xnor UO_1637 (O_1637,N_14924,N_14867);
nand UO_1638 (O_1638,N_14764,N_14817);
nor UO_1639 (O_1639,N_14859,N_14882);
and UO_1640 (O_1640,N_14952,N_14913);
nor UO_1641 (O_1641,N_14921,N_14873);
or UO_1642 (O_1642,N_14939,N_14838);
xnor UO_1643 (O_1643,N_14945,N_14890);
xnor UO_1644 (O_1644,N_14832,N_14995);
or UO_1645 (O_1645,N_14941,N_14849);
nand UO_1646 (O_1646,N_14961,N_14980);
xnor UO_1647 (O_1647,N_14898,N_14893);
or UO_1648 (O_1648,N_14897,N_14847);
nor UO_1649 (O_1649,N_14881,N_14939);
xor UO_1650 (O_1650,N_14859,N_14911);
nor UO_1651 (O_1651,N_14912,N_14997);
nor UO_1652 (O_1652,N_14870,N_14752);
or UO_1653 (O_1653,N_14948,N_14891);
nor UO_1654 (O_1654,N_14794,N_14756);
or UO_1655 (O_1655,N_14788,N_14965);
xor UO_1656 (O_1656,N_14797,N_14876);
xor UO_1657 (O_1657,N_14949,N_14796);
or UO_1658 (O_1658,N_14842,N_14930);
nand UO_1659 (O_1659,N_14784,N_14759);
nor UO_1660 (O_1660,N_14892,N_14936);
and UO_1661 (O_1661,N_14978,N_14913);
and UO_1662 (O_1662,N_14818,N_14765);
nor UO_1663 (O_1663,N_14784,N_14835);
and UO_1664 (O_1664,N_14893,N_14885);
nor UO_1665 (O_1665,N_14816,N_14962);
and UO_1666 (O_1666,N_14848,N_14916);
and UO_1667 (O_1667,N_14963,N_14867);
and UO_1668 (O_1668,N_14923,N_14901);
and UO_1669 (O_1669,N_14962,N_14943);
or UO_1670 (O_1670,N_14805,N_14884);
and UO_1671 (O_1671,N_14825,N_14886);
or UO_1672 (O_1672,N_14881,N_14819);
or UO_1673 (O_1673,N_14933,N_14818);
xnor UO_1674 (O_1674,N_14984,N_14927);
xnor UO_1675 (O_1675,N_14822,N_14940);
and UO_1676 (O_1676,N_14794,N_14962);
nand UO_1677 (O_1677,N_14820,N_14977);
nand UO_1678 (O_1678,N_14800,N_14984);
xor UO_1679 (O_1679,N_14999,N_14822);
or UO_1680 (O_1680,N_14949,N_14829);
nand UO_1681 (O_1681,N_14813,N_14893);
nand UO_1682 (O_1682,N_14987,N_14793);
nor UO_1683 (O_1683,N_14826,N_14820);
nand UO_1684 (O_1684,N_14989,N_14820);
xor UO_1685 (O_1685,N_14966,N_14942);
nand UO_1686 (O_1686,N_14960,N_14891);
and UO_1687 (O_1687,N_14932,N_14971);
xor UO_1688 (O_1688,N_14919,N_14883);
and UO_1689 (O_1689,N_14833,N_14867);
or UO_1690 (O_1690,N_14960,N_14847);
or UO_1691 (O_1691,N_14905,N_14888);
or UO_1692 (O_1692,N_14752,N_14907);
and UO_1693 (O_1693,N_14907,N_14893);
nor UO_1694 (O_1694,N_14929,N_14970);
nand UO_1695 (O_1695,N_14808,N_14792);
and UO_1696 (O_1696,N_14987,N_14977);
nand UO_1697 (O_1697,N_14764,N_14750);
and UO_1698 (O_1698,N_14766,N_14956);
nor UO_1699 (O_1699,N_14854,N_14983);
and UO_1700 (O_1700,N_14787,N_14921);
nor UO_1701 (O_1701,N_14999,N_14968);
and UO_1702 (O_1702,N_14928,N_14839);
and UO_1703 (O_1703,N_14823,N_14966);
nand UO_1704 (O_1704,N_14851,N_14881);
nand UO_1705 (O_1705,N_14837,N_14970);
xor UO_1706 (O_1706,N_14773,N_14905);
or UO_1707 (O_1707,N_14950,N_14796);
nand UO_1708 (O_1708,N_14862,N_14911);
and UO_1709 (O_1709,N_14793,N_14901);
or UO_1710 (O_1710,N_14907,N_14770);
and UO_1711 (O_1711,N_14988,N_14820);
nand UO_1712 (O_1712,N_14985,N_14992);
and UO_1713 (O_1713,N_14760,N_14981);
nor UO_1714 (O_1714,N_14819,N_14778);
or UO_1715 (O_1715,N_14846,N_14946);
nor UO_1716 (O_1716,N_14834,N_14860);
nand UO_1717 (O_1717,N_14757,N_14967);
xnor UO_1718 (O_1718,N_14834,N_14938);
and UO_1719 (O_1719,N_14790,N_14782);
xor UO_1720 (O_1720,N_14832,N_14913);
and UO_1721 (O_1721,N_14910,N_14824);
and UO_1722 (O_1722,N_14987,N_14763);
nor UO_1723 (O_1723,N_14787,N_14756);
or UO_1724 (O_1724,N_14752,N_14987);
or UO_1725 (O_1725,N_14885,N_14771);
nand UO_1726 (O_1726,N_14836,N_14770);
and UO_1727 (O_1727,N_14958,N_14791);
nor UO_1728 (O_1728,N_14795,N_14806);
or UO_1729 (O_1729,N_14935,N_14902);
and UO_1730 (O_1730,N_14943,N_14983);
or UO_1731 (O_1731,N_14922,N_14906);
and UO_1732 (O_1732,N_14782,N_14762);
xor UO_1733 (O_1733,N_14900,N_14810);
xnor UO_1734 (O_1734,N_14940,N_14854);
xnor UO_1735 (O_1735,N_14922,N_14907);
nand UO_1736 (O_1736,N_14791,N_14856);
nor UO_1737 (O_1737,N_14883,N_14781);
nand UO_1738 (O_1738,N_14961,N_14785);
and UO_1739 (O_1739,N_14989,N_14799);
and UO_1740 (O_1740,N_14908,N_14926);
xor UO_1741 (O_1741,N_14836,N_14874);
nor UO_1742 (O_1742,N_14844,N_14992);
nand UO_1743 (O_1743,N_14976,N_14897);
nand UO_1744 (O_1744,N_14869,N_14940);
or UO_1745 (O_1745,N_14882,N_14861);
nand UO_1746 (O_1746,N_14752,N_14984);
nand UO_1747 (O_1747,N_14839,N_14781);
nand UO_1748 (O_1748,N_14889,N_14953);
or UO_1749 (O_1749,N_14916,N_14937);
or UO_1750 (O_1750,N_14826,N_14980);
nand UO_1751 (O_1751,N_14971,N_14796);
or UO_1752 (O_1752,N_14814,N_14959);
nor UO_1753 (O_1753,N_14819,N_14992);
and UO_1754 (O_1754,N_14815,N_14821);
nand UO_1755 (O_1755,N_14947,N_14766);
and UO_1756 (O_1756,N_14821,N_14786);
and UO_1757 (O_1757,N_14874,N_14951);
and UO_1758 (O_1758,N_14980,N_14775);
xnor UO_1759 (O_1759,N_14778,N_14828);
nor UO_1760 (O_1760,N_14957,N_14971);
nand UO_1761 (O_1761,N_14887,N_14998);
and UO_1762 (O_1762,N_14951,N_14826);
and UO_1763 (O_1763,N_14878,N_14870);
and UO_1764 (O_1764,N_14875,N_14969);
and UO_1765 (O_1765,N_14851,N_14776);
or UO_1766 (O_1766,N_14932,N_14801);
or UO_1767 (O_1767,N_14811,N_14785);
nor UO_1768 (O_1768,N_14916,N_14957);
nor UO_1769 (O_1769,N_14832,N_14867);
and UO_1770 (O_1770,N_14980,N_14819);
nor UO_1771 (O_1771,N_14860,N_14826);
nor UO_1772 (O_1772,N_14845,N_14886);
nor UO_1773 (O_1773,N_14853,N_14763);
nand UO_1774 (O_1774,N_14935,N_14891);
xor UO_1775 (O_1775,N_14890,N_14982);
or UO_1776 (O_1776,N_14947,N_14797);
xnor UO_1777 (O_1777,N_14963,N_14908);
and UO_1778 (O_1778,N_14946,N_14955);
or UO_1779 (O_1779,N_14856,N_14818);
nor UO_1780 (O_1780,N_14948,N_14785);
nor UO_1781 (O_1781,N_14810,N_14866);
or UO_1782 (O_1782,N_14965,N_14977);
or UO_1783 (O_1783,N_14933,N_14866);
or UO_1784 (O_1784,N_14859,N_14848);
xnor UO_1785 (O_1785,N_14915,N_14896);
xnor UO_1786 (O_1786,N_14762,N_14943);
nor UO_1787 (O_1787,N_14796,N_14812);
and UO_1788 (O_1788,N_14936,N_14761);
nand UO_1789 (O_1789,N_14750,N_14994);
xnor UO_1790 (O_1790,N_14758,N_14771);
or UO_1791 (O_1791,N_14907,N_14789);
nand UO_1792 (O_1792,N_14769,N_14988);
nor UO_1793 (O_1793,N_14946,N_14909);
or UO_1794 (O_1794,N_14870,N_14756);
and UO_1795 (O_1795,N_14991,N_14800);
nor UO_1796 (O_1796,N_14835,N_14837);
nand UO_1797 (O_1797,N_14755,N_14872);
nor UO_1798 (O_1798,N_14986,N_14896);
and UO_1799 (O_1799,N_14786,N_14848);
or UO_1800 (O_1800,N_14908,N_14755);
nand UO_1801 (O_1801,N_14984,N_14963);
nand UO_1802 (O_1802,N_14878,N_14792);
xnor UO_1803 (O_1803,N_14952,N_14770);
or UO_1804 (O_1804,N_14989,N_14817);
nand UO_1805 (O_1805,N_14936,N_14901);
nand UO_1806 (O_1806,N_14898,N_14993);
xor UO_1807 (O_1807,N_14859,N_14933);
or UO_1808 (O_1808,N_14996,N_14859);
nand UO_1809 (O_1809,N_14880,N_14897);
nand UO_1810 (O_1810,N_14887,N_14882);
nor UO_1811 (O_1811,N_14981,N_14756);
and UO_1812 (O_1812,N_14966,N_14776);
nor UO_1813 (O_1813,N_14907,N_14884);
nor UO_1814 (O_1814,N_14826,N_14913);
and UO_1815 (O_1815,N_14924,N_14958);
or UO_1816 (O_1816,N_14783,N_14979);
nand UO_1817 (O_1817,N_14868,N_14924);
nor UO_1818 (O_1818,N_14854,N_14898);
and UO_1819 (O_1819,N_14986,N_14898);
xor UO_1820 (O_1820,N_14774,N_14934);
and UO_1821 (O_1821,N_14905,N_14961);
nand UO_1822 (O_1822,N_14799,N_14870);
and UO_1823 (O_1823,N_14952,N_14919);
and UO_1824 (O_1824,N_14759,N_14855);
nand UO_1825 (O_1825,N_14908,N_14759);
xor UO_1826 (O_1826,N_14810,N_14931);
nand UO_1827 (O_1827,N_14760,N_14976);
or UO_1828 (O_1828,N_14993,N_14995);
and UO_1829 (O_1829,N_14927,N_14767);
nand UO_1830 (O_1830,N_14888,N_14866);
and UO_1831 (O_1831,N_14756,N_14817);
nor UO_1832 (O_1832,N_14897,N_14812);
or UO_1833 (O_1833,N_14807,N_14867);
xor UO_1834 (O_1834,N_14948,N_14788);
nand UO_1835 (O_1835,N_14919,N_14893);
or UO_1836 (O_1836,N_14968,N_14806);
nor UO_1837 (O_1837,N_14937,N_14922);
and UO_1838 (O_1838,N_14901,N_14761);
nand UO_1839 (O_1839,N_14873,N_14902);
nand UO_1840 (O_1840,N_14808,N_14827);
nor UO_1841 (O_1841,N_14920,N_14811);
xor UO_1842 (O_1842,N_14956,N_14774);
nor UO_1843 (O_1843,N_14879,N_14778);
nand UO_1844 (O_1844,N_14799,N_14997);
nand UO_1845 (O_1845,N_14880,N_14855);
and UO_1846 (O_1846,N_14935,N_14939);
or UO_1847 (O_1847,N_14802,N_14993);
and UO_1848 (O_1848,N_14975,N_14959);
nand UO_1849 (O_1849,N_14916,N_14834);
nor UO_1850 (O_1850,N_14854,N_14915);
nand UO_1851 (O_1851,N_14831,N_14910);
nor UO_1852 (O_1852,N_14806,N_14900);
nor UO_1853 (O_1853,N_14903,N_14753);
xnor UO_1854 (O_1854,N_14937,N_14801);
xnor UO_1855 (O_1855,N_14972,N_14855);
and UO_1856 (O_1856,N_14878,N_14911);
and UO_1857 (O_1857,N_14841,N_14991);
and UO_1858 (O_1858,N_14868,N_14783);
xnor UO_1859 (O_1859,N_14799,N_14827);
or UO_1860 (O_1860,N_14919,N_14900);
nand UO_1861 (O_1861,N_14898,N_14826);
and UO_1862 (O_1862,N_14842,N_14865);
xor UO_1863 (O_1863,N_14845,N_14962);
nor UO_1864 (O_1864,N_14915,N_14930);
or UO_1865 (O_1865,N_14783,N_14849);
nand UO_1866 (O_1866,N_14827,N_14848);
or UO_1867 (O_1867,N_14985,N_14811);
nand UO_1868 (O_1868,N_14924,N_14846);
nor UO_1869 (O_1869,N_14903,N_14764);
nor UO_1870 (O_1870,N_14892,N_14933);
and UO_1871 (O_1871,N_14949,N_14854);
or UO_1872 (O_1872,N_14763,N_14867);
and UO_1873 (O_1873,N_14942,N_14960);
and UO_1874 (O_1874,N_14809,N_14905);
or UO_1875 (O_1875,N_14886,N_14894);
and UO_1876 (O_1876,N_14818,N_14806);
and UO_1877 (O_1877,N_14983,N_14883);
xor UO_1878 (O_1878,N_14877,N_14978);
nand UO_1879 (O_1879,N_14886,N_14906);
and UO_1880 (O_1880,N_14958,N_14820);
nor UO_1881 (O_1881,N_14788,N_14851);
xor UO_1882 (O_1882,N_14752,N_14921);
or UO_1883 (O_1883,N_14791,N_14834);
xnor UO_1884 (O_1884,N_14783,N_14767);
nor UO_1885 (O_1885,N_14973,N_14951);
xnor UO_1886 (O_1886,N_14875,N_14890);
xor UO_1887 (O_1887,N_14951,N_14845);
and UO_1888 (O_1888,N_14943,N_14783);
nand UO_1889 (O_1889,N_14755,N_14850);
and UO_1890 (O_1890,N_14899,N_14826);
and UO_1891 (O_1891,N_14892,N_14839);
nand UO_1892 (O_1892,N_14793,N_14847);
xor UO_1893 (O_1893,N_14915,N_14840);
xor UO_1894 (O_1894,N_14842,N_14901);
nor UO_1895 (O_1895,N_14971,N_14933);
and UO_1896 (O_1896,N_14856,N_14815);
and UO_1897 (O_1897,N_14952,N_14881);
nor UO_1898 (O_1898,N_14959,N_14820);
nand UO_1899 (O_1899,N_14977,N_14942);
or UO_1900 (O_1900,N_14874,N_14815);
or UO_1901 (O_1901,N_14795,N_14816);
or UO_1902 (O_1902,N_14768,N_14859);
nand UO_1903 (O_1903,N_14815,N_14903);
nand UO_1904 (O_1904,N_14887,N_14837);
and UO_1905 (O_1905,N_14885,N_14897);
nor UO_1906 (O_1906,N_14757,N_14945);
nor UO_1907 (O_1907,N_14940,N_14776);
xor UO_1908 (O_1908,N_14994,N_14771);
nor UO_1909 (O_1909,N_14862,N_14966);
and UO_1910 (O_1910,N_14893,N_14849);
or UO_1911 (O_1911,N_14819,N_14775);
xor UO_1912 (O_1912,N_14914,N_14907);
nand UO_1913 (O_1913,N_14902,N_14976);
nand UO_1914 (O_1914,N_14791,N_14754);
or UO_1915 (O_1915,N_14813,N_14877);
or UO_1916 (O_1916,N_14978,N_14811);
xnor UO_1917 (O_1917,N_14762,N_14829);
and UO_1918 (O_1918,N_14788,N_14923);
or UO_1919 (O_1919,N_14820,N_14996);
and UO_1920 (O_1920,N_14964,N_14764);
and UO_1921 (O_1921,N_14825,N_14810);
xor UO_1922 (O_1922,N_14893,N_14883);
xor UO_1923 (O_1923,N_14894,N_14884);
xor UO_1924 (O_1924,N_14826,N_14983);
xor UO_1925 (O_1925,N_14808,N_14997);
nand UO_1926 (O_1926,N_14915,N_14812);
nor UO_1927 (O_1927,N_14948,N_14840);
xnor UO_1928 (O_1928,N_14879,N_14987);
nor UO_1929 (O_1929,N_14911,N_14843);
and UO_1930 (O_1930,N_14887,N_14970);
or UO_1931 (O_1931,N_14832,N_14914);
or UO_1932 (O_1932,N_14928,N_14793);
or UO_1933 (O_1933,N_14861,N_14872);
nor UO_1934 (O_1934,N_14994,N_14911);
or UO_1935 (O_1935,N_14799,N_14805);
and UO_1936 (O_1936,N_14892,N_14951);
or UO_1937 (O_1937,N_14962,N_14978);
xnor UO_1938 (O_1938,N_14916,N_14826);
xnor UO_1939 (O_1939,N_14944,N_14863);
nand UO_1940 (O_1940,N_14986,N_14958);
or UO_1941 (O_1941,N_14875,N_14766);
nand UO_1942 (O_1942,N_14935,N_14805);
nor UO_1943 (O_1943,N_14996,N_14975);
and UO_1944 (O_1944,N_14840,N_14788);
nor UO_1945 (O_1945,N_14770,N_14789);
and UO_1946 (O_1946,N_14788,N_14771);
nor UO_1947 (O_1947,N_14975,N_14752);
nor UO_1948 (O_1948,N_14806,N_14823);
xnor UO_1949 (O_1949,N_14953,N_14829);
nor UO_1950 (O_1950,N_14980,N_14899);
nor UO_1951 (O_1951,N_14913,N_14822);
nor UO_1952 (O_1952,N_14888,N_14999);
xnor UO_1953 (O_1953,N_14867,N_14847);
xnor UO_1954 (O_1954,N_14982,N_14826);
nor UO_1955 (O_1955,N_14766,N_14978);
xnor UO_1956 (O_1956,N_14930,N_14838);
xor UO_1957 (O_1957,N_14900,N_14935);
and UO_1958 (O_1958,N_14952,N_14903);
or UO_1959 (O_1959,N_14770,N_14834);
and UO_1960 (O_1960,N_14799,N_14931);
and UO_1961 (O_1961,N_14983,N_14807);
xnor UO_1962 (O_1962,N_14884,N_14868);
nor UO_1963 (O_1963,N_14876,N_14988);
or UO_1964 (O_1964,N_14934,N_14962);
nand UO_1965 (O_1965,N_14862,N_14895);
and UO_1966 (O_1966,N_14827,N_14757);
nor UO_1967 (O_1967,N_14762,N_14980);
nand UO_1968 (O_1968,N_14842,N_14869);
and UO_1969 (O_1969,N_14946,N_14894);
xor UO_1970 (O_1970,N_14885,N_14850);
nand UO_1971 (O_1971,N_14787,N_14798);
nand UO_1972 (O_1972,N_14861,N_14905);
xnor UO_1973 (O_1973,N_14958,N_14854);
xor UO_1974 (O_1974,N_14865,N_14938);
xnor UO_1975 (O_1975,N_14835,N_14773);
nor UO_1976 (O_1976,N_14844,N_14836);
nor UO_1977 (O_1977,N_14997,N_14786);
nor UO_1978 (O_1978,N_14805,N_14970);
and UO_1979 (O_1979,N_14858,N_14922);
xor UO_1980 (O_1980,N_14905,N_14992);
nor UO_1981 (O_1981,N_14858,N_14990);
xor UO_1982 (O_1982,N_14934,N_14936);
xnor UO_1983 (O_1983,N_14858,N_14782);
and UO_1984 (O_1984,N_14847,N_14889);
and UO_1985 (O_1985,N_14876,N_14834);
nor UO_1986 (O_1986,N_14876,N_14829);
xor UO_1987 (O_1987,N_14927,N_14873);
or UO_1988 (O_1988,N_14804,N_14856);
and UO_1989 (O_1989,N_14806,N_14930);
xor UO_1990 (O_1990,N_14781,N_14858);
nor UO_1991 (O_1991,N_14941,N_14752);
nor UO_1992 (O_1992,N_14819,N_14783);
xnor UO_1993 (O_1993,N_14854,N_14816);
or UO_1994 (O_1994,N_14781,N_14842);
nand UO_1995 (O_1995,N_14899,N_14912);
nand UO_1996 (O_1996,N_14945,N_14967);
nor UO_1997 (O_1997,N_14932,N_14814);
nor UO_1998 (O_1998,N_14800,N_14917);
and UO_1999 (O_1999,N_14809,N_14941);
endmodule