module basic_750_5000_1000_25_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_587,In_168);
nor U1 (N_1,In_637,In_131);
nor U2 (N_2,In_713,In_583);
or U3 (N_3,In_236,In_731);
nand U4 (N_4,In_262,In_634);
xor U5 (N_5,In_647,In_288);
xor U6 (N_6,In_151,In_567);
nor U7 (N_7,In_163,In_613);
nand U8 (N_8,In_86,In_15);
or U9 (N_9,In_721,In_569);
and U10 (N_10,In_114,In_492);
nor U11 (N_11,In_626,In_242);
nand U12 (N_12,In_271,In_176);
nor U13 (N_13,In_400,In_680);
nor U14 (N_14,In_379,In_574);
nor U15 (N_15,In_497,In_289);
nand U16 (N_16,In_3,In_748);
xor U17 (N_17,In_164,In_211);
nand U18 (N_18,In_710,In_295);
or U19 (N_19,In_93,In_430);
or U20 (N_20,In_505,In_280);
or U21 (N_21,In_432,In_132);
nand U22 (N_22,In_126,In_630);
or U23 (N_23,In_408,In_204);
and U24 (N_24,In_364,In_403);
nor U25 (N_25,In_718,In_150);
nand U26 (N_26,In_40,In_452);
xor U27 (N_27,In_405,In_458);
or U28 (N_28,In_709,In_140);
xnor U29 (N_29,In_217,In_740);
nand U30 (N_30,In_627,In_592);
or U31 (N_31,In_376,In_658);
and U32 (N_32,In_555,In_181);
nor U33 (N_33,In_623,In_621);
nor U34 (N_34,In_120,In_187);
xnor U35 (N_35,In_744,In_27);
nand U36 (N_36,In_87,In_253);
and U37 (N_37,In_322,In_196);
nand U38 (N_38,In_509,In_410);
or U39 (N_39,In_531,In_314);
nand U40 (N_40,In_707,In_213);
or U41 (N_41,In_231,In_661);
nand U42 (N_42,In_708,In_423);
xnor U43 (N_43,In_97,In_160);
and U44 (N_44,In_687,In_536);
xor U45 (N_45,In_340,In_38);
nand U46 (N_46,In_420,In_734);
and U47 (N_47,In_477,In_94);
or U48 (N_48,In_304,In_109);
or U49 (N_49,In_113,In_69);
or U50 (N_50,In_527,In_240);
and U51 (N_51,In_427,In_572);
nand U52 (N_52,In_66,In_673);
xnor U53 (N_53,In_716,In_350);
nor U54 (N_54,In_655,In_538);
xnor U55 (N_55,In_169,In_317);
nand U56 (N_56,In_218,In_115);
nor U57 (N_57,In_232,In_153);
nand U58 (N_58,In_639,In_471);
nand U59 (N_59,In_25,In_101);
and U60 (N_60,In_287,In_476);
and U61 (N_61,In_368,In_679);
nor U62 (N_62,In_186,In_541);
and U63 (N_63,In_83,In_336);
or U64 (N_64,In_89,In_535);
xnor U65 (N_65,In_515,In_136);
xnor U66 (N_66,In_33,In_631);
and U67 (N_67,In_300,In_450);
and U68 (N_68,In_278,In_440);
and U69 (N_69,In_498,In_31);
nor U70 (N_70,In_103,In_216);
xor U71 (N_71,In_202,In_618);
nor U72 (N_72,In_306,In_399);
nand U73 (N_73,In_389,In_17);
and U74 (N_74,In_666,In_124);
nor U75 (N_75,In_699,In_274);
xnor U76 (N_76,In_615,In_585);
or U77 (N_77,In_539,In_270);
and U78 (N_78,In_528,In_434);
or U79 (N_79,In_229,In_469);
xor U80 (N_80,In_199,In_603);
nand U81 (N_81,In_92,In_468);
xor U82 (N_82,In_52,In_155);
nand U83 (N_83,In_127,In_723);
or U84 (N_84,In_313,In_51);
or U85 (N_85,In_294,In_532);
or U86 (N_86,In_510,In_173);
nor U87 (N_87,In_475,In_417);
and U88 (N_88,In_332,In_650);
or U89 (N_89,In_682,In_39);
xor U90 (N_90,In_286,In_425);
xor U91 (N_91,In_501,In_593);
nor U92 (N_92,In_13,In_111);
nand U93 (N_93,In_348,In_674);
nor U94 (N_94,In_544,In_62);
and U95 (N_95,In_586,In_657);
xor U96 (N_96,In_606,In_642);
or U97 (N_97,In_193,In_273);
xor U98 (N_98,In_342,In_506);
and U99 (N_99,In_580,In_261);
or U100 (N_100,In_424,In_326);
xor U101 (N_101,In_435,In_416);
and U102 (N_102,In_523,In_601);
xnor U103 (N_103,In_652,In_0);
nor U104 (N_104,In_148,In_10);
xnor U105 (N_105,In_363,In_610);
and U106 (N_106,In_362,In_293);
xnor U107 (N_107,In_7,In_45);
nor U108 (N_108,In_684,In_547);
xor U109 (N_109,In_341,In_490);
nand U110 (N_110,In_594,In_23);
or U111 (N_111,In_43,In_197);
or U112 (N_112,In_358,In_352);
nand U113 (N_113,In_299,In_693);
and U114 (N_114,In_144,In_59);
or U115 (N_115,In_483,In_503);
xor U116 (N_116,In_398,In_14);
and U117 (N_117,In_701,In_409);
nand U118 (N_118,In_316,In_269);
nor U119 (N_119,In_695,In_455);
xor U120 (N_120,In_486,In_99);
nor U121 (N_121,In_491,In_456);
xor U122 (N_122,In_656,In_5);
nand U123 (N_123,In_102,In_500);
xnor U124 (N_124,In_502,In_129);
and U125 (N_125,In_714,In_577);
and U126 (N_126,In_524,In_525);
or U127 (N_127,In_2,In_234);
xor U128 (N_128,In_225,In_565);
xnor U129 (N_129,In_357,In_275);
and U130 (N_130,In_268,In_690);
or U131 (N_131,In_119,In_104);
or U132 (N_132,In_96,In_643);
nand U133 (N_133,In_54,In_521);
xor U134 (N_134,In_121,In_75);
and U135 (N_135,In_42,In_677);
nand U136 (N_136,In_619,In_488);
xnor U137 (N_137,In_739,In_551);
or U138 (N_138,In_422,In_743);
nand U139 (N_139,In_238,In_404);
and U140 (N_140,In_210,In_382);
nand U141 (N_141,In_412,In_122);
and U142 (N_142,In_720,In_371);
and U143 (N_143,In_214,In_206);
xnor U144 (N_144,In_365,In_705);
or U145 (N_145,In_442,In_493);
nor U146 (N_146,In_198,In_47);
nor U147 (N_147,In_11,In_737);
or U148 (N_148,In_175,In_465);
or U149 (N_149,In_495,In_159);
nor U150 (N_150,In_745,In_448);
xor U151 (N_151,In_641,In_557);
xor U152 (N_152,In_582,In_161);
nor U153 (N_153,In_530,In_243);
or U154 (N_154,In_543,In_685);
nor U155 (N_155,In_715,In_349);
or U156 (N_156,In_29,In_648);
nor U157 (N_157,In_296,In_518);
or U158 (N_158,In_374,In_323);
or U159 (N_159,In_507,In_71);
nor U160 (N_160,In_616,In_562);
nor U161 (N_161,In_381,In_56);
nand U162 (N_162,In_667,In_60);
xor U163 (N_163,In_391,In_135);
xor U164 (N_164,In_254,In_628);
nand U165 (N_165,In_90,In_375);
nor U166 (N_166,In_264,In_325);
and U167 (N_167,In_702,In_34);
and U168 (N_168,In_449,In_252);
xor U169 (N_169,In_522,In_519);
nand U170 (N_170,In_607,In_177);
nor U171 (N_171,In_517,In_479);
nand U172 (N_172,In_653,In_730);
nor U173 (N_173,In_72,In_327);
or U174 (N_174,In_308,In_372);
xnor U175 (N_175,In_474,In_200);
or U176 (N_176,In_73,In_370);
nor U177 (N_177,In_670,In_24);
or U178 (N_178,In_41,In_611);
xnor U179 (N_179,In_233,In_85);
nor U180 (N_180,In_282,In_9);
and U181 (N_181,In_180,In_116);
nand U182 (N_182,In_726,In_549);
or U183 (N_183,In_166,In_152);
and U184 (N_184,In_719,In_665);
or U185 (N_185,In_335,In_575);
or U186 (N_186,In_37,In_227);
or U187 (N_187,In_333,In_478);
nor U188 (N_188,In_76,In_22);
xnor U189 (N_189,In_346,In_383);
xor U190 (N_190,In_138,In_728);
nor U191 (N_191,In_290,In_481);
and U192 (N_192,In_504,In_46);
nor U193 (N_193,In_443,In_499);
nor U194 (N_194,In_30,In_453);
nor U195 (N_195,In_598,In_741);
xnor U196 (N_196,In_185,In_265);
nand U197 (N_197,In_165,In_407);
and U198 (N_198,In_390,In_251);
and U199 (N_199,In_18,In_259);
nand U200 (N_200,N_51,In_188);
xnor U201 (N_201,In_484,In_546);
nand U202 (N_202,N_15,N_180);
and U203 (N_203,In_513,In_386);
nor U204 (N_204,N_111,In_545);
and U205 (N_205,N_98,N_62);
nor U206 (N_206,In_742,N_156);
and U207 (N_207,In_310,In_636);
nand U208 (N_208,N_112,In_8);
and U209 (N_209,N_193,In_605);
and U210 (N_210,In_130,N_66);
xor U211 (N_211,N_13,In_145);
or U212 (N_212,N_90,N_143);
nor U213 (N_213,In_429,In_277);
and U214 (N_214,In_19,In_329);
xor U215 (N_215,N_37,In_201);
nand U216 (N_216,In_260,In_80);
or U217 (N_217,In_624,N_131);
or U218 (N_218,In_339,N_83);
xnor U219 (N_219,N_25,N_91);
and U220 (N_220,In_529,N_142);
or U221 (N_221,In_561,In_170);
or U222 (N_222,N_115,N_113);
nor U223 (N_223,In_651,In_230);
xnor U224 (N_224,N_153,In_550);
and U225 (N_225,In_671,In_117);
or U226 (N_226,In_596,N_157);
and U227 (N_227,N_126,In_344);
and U228 (N_228,In_315,In_589);
and U229 (N_229,In_267,In_467);
nand U230 (N_230,In_88,In_178);
or U231 (N_231,In_65,N_47);
xnor U232 (N_232,N_137,N_54);
nand U233 (N_233,In_182,In_139);
and U234 (N_234,N_163,N_11);
xor U235 (N_235,N_30,N_12);
and U236 (N_236,In_485,In_415);
and U237 (N_237,In_413,In_747);
or U238 (N_238,In_397,In_428);
nand U239 (N_239,In_167,N_16);
or U240 (N_240,In_533,N_110);
and U241 (N_241,N_72,In_172);
nand U242 (N_242,N_123,N_139);
xor U243 (N_243,In_118,In_303);
nor U244 (N_244,In_128,In_209);
xor U245 (N_245,In_353,N_9);
or U246 (N_246,In_645,In_292);
nor U247 (N_247,In_334,In_77);
nor U248 (N_248,In_604,N_70);
nor U249 (N_249,N_71,In_394);
and U250 (N_250,In_402,In_692);
or U251 (N_251,N_128,In_722);
nor U252 (N_252,In_686,In_58);
xnor U253 (N_253,N_102,N_35);
or U254 (N_254,N_175,In_49);
nand U255 (N_255,N_189,In_622);
xnor U256 (N_256,N_26,N_105);
or U257 (N_257,N_162,N_40);
or U258 (N_258,In_222,N_184);
xor U259 (N_259,In_359,In_84);
nand U260 (N_260,N_141,In_662);
or U261 (N_261,In_711,In_570);
xnor U262 (N_262,N_107,N_186);
and U263 (N_263,In_57,In_414);
nand U264 (N_264,N_140,In_307);
nand U265 (N_265,N_183,In_143);
nand U266 (N_266,In_330,N_19);
xor U267 (N_267,In_608,N_65);
nand U268 (N_268,N_196,N_147);
or U269 (N_269,N_22,N_192);
and U270 (N_270,In_257,N_109);
and U271 (N_271,In_612,In_584);
nand U272 (N_272,N_178,N_10);
nand U273 (N_273,N_36,N_172);
xor U274 (N_274,In_331,N_46);
and U275 (N_275,N_58,N_79);
nand U276 (N_276,In_134,N_39);
or U277 (N_277,N_174,N_81);
xnor U278 (N_278,In_411,In_355);
or U279 (N_279,In_560,In_675);
nand U280 (N_280,In_98,In_595);
and U281 (N_281,N_132,N_27);
or U282 (N_282,In_246,In_298);
xnor U283 (N_283,In_746,In_678);
or U284 (N_284,N_76,In_717);
nor U285 (N_285,In_581,In_190);
nor U286 (N_286,In_16,In_324);
nand U287 (N_287,N_38,In_377);
nand U288 (N_288,In_305,In_681);
or U289 (N_289,N_129,N_8);
xor U290 (N_290,N_114,N_138);
or U291 (N_291,In_194,In_276);
or U292 (N_292,In_683,In_573);
nor U293 (N_293,In_633,In_110);
xor U294 (N_294,In_28,N_74);
xor U295 (N_295,N_21,In_157);
or U296 (N_296,In_632,In_179);
nand U297 (N_297,N_50,In_640);
nand U298 (N_298,In_32,N_0);
and U299 (N_299,In_749,In_107);
and U300 (N_300,In_419,N_20);
and U301 (N_301,In_55,N_198);
or U302 (N_302,In_691,In_64);
or U303 (N_303,In_67,In_360);
or U304 (N_304,In_380,N_57);
nor U305 (N_305,In_247,In_571);
nor U306 (N_306,In_318,In_378);
nor U307 (N_307,In_664,In_361);
nor U308 (N_308,In_215,In_149);
nor U309 (N_309,N_146,N_135);
or U310 (N_310,N_101,N_42);
xnor U311 (N_311,In_105,In_660);
nor U312 (N_312,In_301,In_462);
and U313 (N_313,In_508,In_100);
nand U314 (N_314,In_602,In_548);
xnor U315 (N_315,In_609,N_75);
or U316 (N_316,In_736,In_511);
nand U317 (N_317,N_14,In_703);
or U318 (N_318,In_454,In_162);
or U319 (N_319,In_255,N_80);
xor U320 (N_320,N_29,N_95);
xor U321 (N_321,In_466,In_563);
and U322 (N_322,In_487,In_438);
or U323 (N_323,In_635,In_223);
nor U324 (N_324,N_185,N_17);
xnor U325 (N_325,N_1,In_444);
or U326 (N_326,In_226,In_431);
nor U327 (N_327,In_473,In_418);
nand U328 (N_328,N_59,N_168);
or U329 (N_329,N_144,In_646);
xor U330 (N_330,In_644,In_297);
and U331 (N_331,In_396,In_472);
and U332 (N_332,In_228,N_161);
and U333 (N_333,In_63,In_241);
and U334 (N_334,N_195,In_366);
nand U335 (N_335,N_43,N_61);
xor U336 (N_336,In_284,In_512);
nand U337 (N_337,In_320,In_625);
nand U338 (N_338,N_197,N_94);
or U339 (N_339,N_99,In_704);
xor U340 (N_340,N_130,N_23);
nand U341 (N_341,N_45,In_464);
nand U342 (N_342,In_540,In_663);
and U343 (N_343,In_266,N_158);
nor U344 (N_344,N_85,In_516);
xor U345 (N_345,N_34,In_590);
or U346 (N_346,In_537,In_356);
or U347 (N_347,N_69,In_174);
nor U348 (N_348,In_345,In_672);
and U349 (N_349,In_6,In_195);
or U350 (N_350,In_554,In_133);
xor U351 (N_351,In_147,N_119);
or U352 (N_352,In_192,In_369);
and U353 (N_353,N_55,In_496);
nor U354 (N_354,In_171,N_108);
or U355 (N_355,In_12,In_461);
or U356 (N_356,N_7,In_50);
nand U357 (N_357,N_87,In_439);
nand U358 (N_358,In_207,In_183);
or U359 (N_359,N_5,N_24);
and U360 (N_360,In_436,N_41);
xor U361 (N_361,In_649,In_35);
and U362 (N_362,In_597,In_735);
nor U363 (N_363,N_6,In_447);
nor U364 (N_364,N_116,In_48);
and U365 (N_365,N_33,N_78);
and U366 (N_366,In_219,In_347);
nand U367 (N_367,In_319,In_248);
and U368 (N_368,In_244,N_187);
nor U369 (N_369,In_79,In_576);
xnor U370 (N_370,N_165,In_732);
xor U371 (N_371,In_617,In_68);
nand U372 (N_372,N_154,In_588);
nand U373 (N_373,In_82,N_82);
nor U374 (N_374,In_36,In_354);
and U375 (N_375,N_164,In_387);
or U376 (N_376,In_579,N_106);
nor U377 (N_377,In_457,N_151);
xnor U378 (N_378,In_309,In_689);
or U379 (N_379,In_21,In_426);
nand U380 (N_380,N_169,In_599);
and U381 (N_381,N_150,In_514);
nand U382 (N_382,In_250,In_669);
nand U383 (N_383,In_125,N_173);
nor U384 (N_384,N_118,In_433);
nor U385 (N_385,In_558,In_239);
and U386 (N_386,In_106,N_44);
xnor U387 (N_387,In_212,In_385);
xnor U388 (N_388,In_81,In_460);
nor U389 (N_389,In_659,N_60);
and U390 (N_390,N_2,In_312);
and U391 (N_391,In_343,N_159);
nor U392 (N_392,N_122,N_179);
nand U393 (N_393,In_388,In_725);
nor U394 (N_394,In_556,In_534);
nand U395 (N_395,N_73,In_446);
xor U396 (N_396,N_124,In_494);
and U397 (N_397,In_482,N_28);
nand U398 (N_398,In_112,N_56);
xor U399 (N_399,In_245,In_568);
xnor U400 (N_400,N_249,N_379);
or U401 (N_401,In_698,N_191);
xnor U402 (N_402,N_358,N_354);
or U403 (N_403,N_364,N_368);
nand U404 (N_404,N_375,N_32);
nand U405 (N_405,N_171,N_223);
nor U406 (N_406,N_304,N_307);
or U407 (N_407,N_170,N_103);
xor U408 (N_408,N_64,In_373);
or U409 (N_409,N_336,N_255);
xor U410 (N_410,N_286,N_394);
and U411 (N_411,In_189,N_264);
nor U412 (N_412,N_244,N_145);
or U413 (N_413,In_78,N_378);
and U414 (N_414,N_356,N_271);
or U415 (N_415,In_4,In_564);
or U416 (N_416,N_299,In_401);
nand U417 (N_417,N_371,N_353);
xnor U418 (N_418,In_1,N_388);
or U419 (N_419,N_373,In_600);
xnor U420 (N_420,N_332,In_367);
or U421 (N_421,N_369,N_225);
nor U422 (N_422,N_277,N_372);
xor U423 (N_423,In_205,N_351);
and U424 (N_424,N_334,In_142);
or U425 (N_425,In_256,N_231);
nand U426 (N_426,N_265,N_246);
xor U427 (N_427,N_276,N_329);
xnor U428 (N_428,N_216,N_392);
and U429 (N_429,In_395,N_238);
nor U430 (N_430,In_61,N_300);
xor U431 (N_431,N_395,In_351);
nor U432 (N_432,N_120,N_308);
nor U433 (N_433,N_322,In_384);
xor U434 (N_434,In_224,N_218);
nand U435 (N_435,In_141,N_194);
xor U436 (N_436,N_222,N_260);
xor U437 (N_437,N_18,N_261);
nor U438 (N_438,N_200,In_263);
xor U439 (N_439,In_542,N_290);
nand U440 (N_440,In_654,N_287);
and U441 (N_441,N_397,In_237);
nor U442 (N_442,In_393,In_26);
nand U443 (N_443,N_291,N_295);
nand U444 (N_444,N_229,In_337);
and U445 (N_445,In_208,N_166);
and U446 (N_446,N_167,In_552);
or U447 (N_447,N_235,N_391);
nor U448 (N_448,N_311,N_134);
nand U449 (N_449,N_152,N_239);
xnor U450 (N_450,N_279,N_219);
xnor U451 (N_451,N_227,N_202);
and U452 (N_452,N_121,N_365);
nand U453 (N_453,N_315,In_74);
and U454 (N_454,N_338,In_480);
nand U455 (N_455,N_345,N_148);
and U456 (N_456,In_235,In_184);
xor U457 (N_457,N_93,N_190);
nor U458 (N_458,N_355,In_108);
and U459 (N_459,N_263,N_292);
and U460 (N_460,N_232,N_243);
and U461 (N_461,In_489,N_237);
nor U462 (N_462,N_294,N_374);
or U463 (N_463,N_335,N_4);
or U464 (N_464,N_350,N_283);
and U465 (N_465,N_63,N_89);
nand U466 (N_466,N_280,N_204);
nand U467 (N_467,N_213,N_252);
xor U468 (N_468,N_288,N_133);
nor U469 (N_469,N_211,N_362);
xor U470 (N_470,N_262,In_70);
nand U471 (N_471,N_381,N_251);
or U472 (N_472,In_156,In_158);
nor U473 (N_473,In_668,N_313);
nor U474 (N_474,N_228,N_349);
xor U475 (N_475,In_697,N_176);
nor U476 (N_476,N_245,N_127);
or U477 (N_477,N_398,N_297);
and U478 (N_478,In_445,N_393);
and U479 (N_479,N_97,N_317);
nor U480 (N_480,In_620,N_323);
and U481 (N_481,N_319,N_370);
and U482 (N_482,In_559,In_154);
or U483 (N_483,N_390,In_220);
nand U484 (N_484,N_247,N_357);
nand U485 (N_485,N_230,N_49);
nand U486 (N_486,N_256,N_327);
nor U487 (N_487,N_301,N_331);
and U488 (N_488,N_347,N_296);
xor U489 (N_489,N_258,N_399);
xor U490 (N_490,N_330,N_289);
or U491 (N_491,N_272,N_377);
or U492 (N_492,In_520,N_100);
or U493 (N_493,In_459,N_343);
or U494 (N_494,N_155,N_352);
xnor U495 (N_495,N_298,N_53);
nand U496 (N_496,N_266,In_676);
or U497 (N_497,N_31,In_470);
nor U498 (N_498,N_217,N_270);
xnor U499 (N_499,In_302,N_241);
or U500 (N_500,In_137,In_526);
and U501 (N_501,In_700,In_738);
xnor U502 (N_502,In_694,N_253);
or U503 (N_503,N_340,N_383);
or U504 (N_504,In_463,In_123);
nor U505 (N_505,N_233,In_441);
and U506 (N_506,N_281,N_309);
nand U507 (N_507,N_333,N_207);
nand U508 (N_508,N_384,N_77);
xor U509 (N_509,N_376,In_566);
or U510 (N_510,N_48,In_629);
and U511 (N_511,In_191,N_396);
nor U512 (N_512,N_382,N_284);
nand U513 (N_513,N_318,N_341);
xnor U514 (N_514,N_305,In_727);
nand U515 (N_515,N_342,In_578);
nor U516 (N_516,N_250,In_733);
nand U517 (N_517,N_92,N_259);
nor U518 (N_518,In_95,N_306);
xor U519 (N_519,In_392,N_324);
nor U520 (N_520,N_220,N_208);
xnor U521 (N_521,N_267,N_337);
xnor U522 (N_522,N_149,N_386);
nor U523 (N_523,N_312,In_20);
xor U524 (N_524,N_117,In_406);
or U525 (N_525,In_451,N_359);
xnor U526 (N_526,N_366,N_236);
or U527 (N_527,N_86,N_361);
and U528 (N_528,In_258,N_274);
nor U529 (N_529,In_688,N_326);
nor U530 (N_530,N_389,N_104);
or U531 (N_531,In_724,N_385);
xnor U532 (N_532,In_285,N_3);
and U533 (N_533,In_729,N_214);
or U534 (N_534,N_254,N_221);
xnor U535 (N_535,N_282,N_346);
and U536 (N_536,N_215,N_201);
and U537 (N_537,N_363,In_712);
or U538 (N_538,N_181,N_321);
xor U539 (N_539,N_316,N_240);
and U540 (N_540,N_125,In_338);
nand U541 (N_541,In_279,N_206);
xor U542 (N_542,N_275,N_360);
nand U543 (N_543,In_421,N_88);
nor U544 (N_544,N_273,N_348);
nand U545 (N_545,In_553,N_199);
or U546 (N_546,N_303,N_52);
nor U547 (N_547,N_136,N_293);
nand U548 (N_548,N_310,In_283);
nand U549 (N_549,N_212,In_91);
or U550 (N_550,N_387,In_706);
nor U551 (N_551,In_328,N_328);
or U552 (N_552,N_257,In_221);
and U553 (N_553,N_242,N_320);
nand U554 (N_554,N_84,N_367);
and U555 (N_555,N_68,N_248);
xor U556 (N_556,In_311,N_188);
xnor U557 (N_557,N_67,N_380);
xnor U558 (N_558,N_314,In_281);
nand U559 (N_559,N_160,N_344);
xnor U560 (N_560,N_210,N_177);
xor U561 (N_561,In_437,N_224);
nor U562 (N_562,N_182,N_268);
or U563 (N_563,N_234,N_278);
nor U564 (N_564,N_269,In_249);
nand U565 (N_565,In_591,N_96);
nor U566 (N_566,In_614,N_203);
nand U567 (N_567,In_638,N_339);
or U568 (N_568,In_44,In_53);
or U569 (N_569,N_209,N_325);
and U570 (N_570,In_291,In_203);
nor U571 (N_571,N_302,N_226);
and U572 (N_572,In_272,In_146);
nand U573 (N_573,In_696,N_285);
nand U574 (N_574,N_205,In_321);
xor U575 (N_575,N_289,In_263);
and U576 (N_576,N_171,N_243);
nor U577 (N_577,In_729,N_280);
xor U578 (N_578,N_239,In_729);
and U579 (N_579,N_225,N_212);
nor U580 (N_580,In_237,N_351);
or U581 (N_581,N_376,N_231);
xnor U582 (N_582,N_364,In_141);
or U583 (N_583,In_256,N_339);
or U584 (N_584,N_386,N_191);
nor U585 (N_585,N_253,N_52);
or U586 (N_586,In_4,N_63);
or U587 (N_587,N_63,In_733);
or U588 (N_588,N_292,N_231);
nand U589 (N_589,In_26,In_638);
and U590 (N_590,N_272,N_233);
and U591 (N_591,In_4,N_245);
or U592 (N_592,N_270,N_245);
nor U593 (N_593,N_210,N_167);
xor U594 (N_594,N_224,N_225);
xor U595 (N_595,N_370,N_97);
and U596 (N_596,In_249,N_256);
nand U597 (N_597,N_318,N_241);
nand U598 (N_598,In_459,In_395);
and U599 (N_599,N_280,N_316);
xnor U600 (N_600,N_463,N_432);
xnor U601 (N_601,N_457,N_587);
xnor U602 (N_602,N_585,N_532);
or U603 (N_603,N_500,N_571);
nor U604 (N_604,N_558,N_486);
and U605 (N_605,N_570,N_450);
or U606 (N_606,N_595,N_522);
or U607 (N_607,N_519,N_593);
xor U608 (N_608,N_481,N_430);
or U609 (N_609,N_572,N_424);
and U610 (N_610,N_557,N_577);
and U611 (N_611,N_435,N_515);
or U612 (N_612,N_584,N_476);
xnor U613 (N_613,N_573,N_555);
and U614 (N_614,N_434,N_443);
nor U615 (N_615,N_512,N_564);
nor U616 (N_616,N_565,N_483);
xnor U617 (N_617,N_507,N_549);
nand U618 (N_618,N_413,N_469);
nor U619 (N_619,N_464,N_495);
xnor U620 (N_620,N_566,N_465);
nor U621 (N_621,N_436,N_451);
and U622 (N_622,N_520,N_505);
xor U623 (N_623,N_438,N_422);
and U624 (N_624,N_477,N_466);
and U625 (N_625,N_586,N_419);
nor U626 (N_626,N_523,N_485);
nand U627 (N_627,N_411,N_460);
nand U628 (N_628,N_590,N_526);
and U629 (N_629,N_578,N_493);
and U630 (N_630,N_404,N_531);
and U631 (N_631,N_423,N_444);
nand U632 (N_632,N_561,N_579);
nor U633 (N_633,N_554,N_425);
nand U634 (N_634,N_442,N_538);
and U635 (N_635,N_491,N_541);
or U636 (N_636,N_440,N_503);
nor U637 (N_637,N_508,N_528);
or U638 (N_638,N_417,N_458);
and U639 (N_639,N_574,N_498);
xor U640 (N_640,N_518,N_427);
and U641 (N_641,N_475,N_405);
and U642 (N_642,N_494,N_599);
xor U643 (N_643,N_559,N_473);
nor U644 (N_644,N_556,N_445);
and U645 (N_645,N_474,N_418);
and U646 (N_646,N_479,N_537);
xnor U647 (N_647,N_502,N_521);
and U648 (N_648,N_535,N_514);
or U649 (N_649,N_470,N_594);
or U650 (N_650,N_478,N_421);
or U651 (N_651,N_420,N_525);
xnor U652 (N_652,N_441,N_544);
or U653 (N_653,N_488,N_472);
nor U654 (N_654,N_468,N_511);
xor U655 (N_655,N_529,N_575);
nor U656 (N_656,N_553,N_580);
nor U657 (N_657,N_416,N_401);
xnor U658 (N_658,N_533,N_539);
and U659 (N_659,N_552,N_545);
and U660 (N_660,N_426,N_467);
and U661 (N_661,N_524,N_596);
or U662 (N_662,N_516,N_489);
or U663 (N_663,N_414,N_415);
nor U664 (N_664,N_402,N_582);
and U665 (N_665,N_403,N_581);
xnor U666 (N_666,N_499,N_448);
nand U667 (N_667,N_562,N_456);
or U668 (N_668,N_509,N_548);
xnor U669 (N_669,N_409,N_452);
or U670 (N_670,N_510,N_407);
and U671 (N_671,N_563,N_412);
nand U672 (N_672,N_543,N_439);
xor U673 (N_673,N_568,N_597);
xnor U674 (N_674,N_497,N_576);
nor U675 (N_675,N_536,N_547);
nor U676 (N_676,N_408,N_455);
and U677 (N_677,N_501,N_546);
nor U678 (N_678,N_527,N_453);
xnor U679 (N_679,N_569,N_530);
nand U680 (N_680,N_461,N_598);
nor U681 (N_681,N_517,N_462);
and U682 (N_682,N_542,N_567);
nand U683 (N_683,N_487,N_496);
xnor U684 (N_684,N_482,N_560);
or U685 (N_685,N_591,N_410);
xor U686 (N_686,N_513,N_437);
xnor U687 (N_687,N_433,N_400);
and U688 (N_688,N_506,N_588);
and U689 (N_689,N_492,N_583);
nand U690 (N_690,N_406,N_447);
nor U691 (N_691,N_446,N_534);
or U692 (N_692,N_592,N_504);
and U693 (N_693,N_550,N_449);
nor U694 (N_694,N_471,N_429);
and U695 (N_695,N_490,N_589);
xor U696 (N_696,N_428,N_480);
or U697 (N_697,N_484,N_454);
or U698 (N_698,N_540,N_551);
and U699 (N_699,N_431,N_459);
nor U700 (N_700,N_502,N_513);
nor U701 (N_701,N_461,N_536);
xnor U702 (N_702,N_548,N_456);
and U703 (N_703,N_543,N_556);
nand U704 (N_704,N_570,N_494);
or U705 (N_705,N_586,N_517);
nand U706 (N_706,N_457,N_583);
nor U707 (N_707,N_497,N_545);
nor U708 (N_708,N_530,N_513);
and U709 (N_709,N_532,N_507);
nand U710 (N_710,N_591,N_433);
or U711 (N_711,N_533,N_559);
and U712 (N_712,N_457,N_419);
nand U713 (N_713,N_466,N_508);
or U714 (N_714,N_526,N_595);
xor U715 (N_715,N_510,N_597);
and U716 (N_716,N_495,N_435);
and U717 (N_717,N_554,N_464);
nor U718 (N_718,N_455,N_457);
nand U719 (N_719,N_474,N_525);
nor U720 (N_720,N_433,N_544);
and U721 (N_721,N_486,N_561);
xnor U722 (N_722,N_479,N_422);
nor U723 (N_723,N_574,N_495);
nand U724 (N_724,N_572,N_435);
xor U725 (N_725,N_444,N_502);
or U726 (N_726,N_537,N_495);
nand U727 (N_727,N_435,N_590);
nor U728 (N_728,N_426,N_546);
nor U729 (N_729,N_567,N_452);
xor U730 (N_730,N_566,N_448);
xnor U731 (N_731,N_437,N_531);
nand U732 (N_732,N_563,N_595);
nand U733 (N_733,N_578,N_518);
xor U734 (N_734,N_541,N_462);
nand U735 (N_735,N_435,N_473);
nand U736 (N_736,N_426,N_561);
and U737 (N_737,N_450,N_408);
nand U738 (N_738,N_588,N_531);
xor U739 (N_739,N_428,N_424);
nor U740 (N_740,N_517,N_445);
xor U741 (N_741,N_488,N_589);
nand U742 (N_742,N_584,N_526);
nor U743 (N_743,N_450,N_522);
or U744 (N_744,N_465,N_417);
xor U745 (N_745,N_417,N_513);
nand U746 (N_746,N_529,N_487);
or U747 (N_747,N_463,N_539);
nor U748 (N_748,N_492,N_511);
nand U749 (N_749,N_581,N_508);
nand U750 (N_750,N_506,N_471);
or U751 (N_751,N_522,N_591);
and U752 (N_752,N_467,N_515);
nand U753 (N_753,N_434,N_511);
and U754 (N_754,N_452,N_510);
nor U755 (N_755,N_540,N_575);
nand U756 (N_756,N_526,N_554);
and U757 (N_757,N_435,N_552);
nand U758 (N_758,N_401,N_496);
xor U759 (N_759,N_549,N_559);
and U760 (N_760,N_473,N_548);
xor U761 (N_761,N_596,N_575);
and U762 (N_762,N_591,N_551);
nand U763 (N_763,N_573,N_548);
xor U764 (N_764,N_443,N_418);
or U765 (N_765,N_441,N_503);
or U766 (N_766,N_434,N_544);
and U767 (N_767,N_493,N_443);
nand U768 (N_768,N_432,N_483);
nand U769 (N_769,N_459,N_417);
and U770 (N_770,N_553,N_595);
and U771 (N_771,N_477,N_418);
nand U772 (N_772,N_432,N_425);
nand U773 (N_773,N_595,N_439);
or U774 (N_774,N_585,N_521);
or U775 (N_775,N_515,N_408);
nor U776 (N_776,N_589,N_473);
or U777 (N_777,N_443,N_436);
or U778 (N_778,N_492,N_401);
nor U779 (N_779,N_443,N_586);
xor U780 (N_780,N_478,N_511);
and U781 (N_781,N_536,N_565);
or U782 (N_782,N_467,N_562);
or U783 (N_783,N_511,N_499);
and U784 (N_784,N_445,N_413);
nor U785 (N_785,N_441,N_454);
xor U786 (N_786,N_409,N_561);
nand U787 (N_787,N_465,N_510);
xnor U788 (N_788,N_528,N_511);
nor U789 (N_789,N_464,N_538);
and U790 (N_790,N_483,N_522);
nor U791 (N_791,N_480,N_561);
and U792 (N_792,N_466,N_552);
and U793 (N_793,N_433,N_597);
or U794 (N_794,N_586,N_507);
nand U795 (N_795,N_566,N_411);
and U796 (N_796,N_524,N_543);
nor U797 (N_797,N_582,N_410);
or U798 (N_798,N_527,N_533);
or U799 (N_799,N_440,N_568);
nand U800 (N_800,N_712,N_784);
nand U801 (N_801,N_714,N_707);
or U802 (N_802,N_652,N_724);
nor U803 (N_803,N_751,N_680);
or U804 (N_804,N_711,N_689);
nor U805 (N_805,N_630,N_640);
xor U806 (N_806,N_683,N_732);
or U807 (N_807,N_781,N_637);
xor U808 (N_808,N_793,N_603);
or U809 (N_809,N_655,N_795);
nor U810 (N_810,N_700,N_612);
or U811 (N_811,N_686,N_765);
and U812 (N_812,N_694,N_737);
or U813 (N_813,N_750,N_664);
xnor U814 (N_814,N_624,N_696);
nand U815 (N_815,N_709,N_705);
nand U816 (N_816,N_717,N_753);
nor U817 (N_817,N_602,N_657);
and U818 (N_818,N_730,N_727);
and U819 (N_819,N_617,N_739);
xor U820 (N_820,N_605,N_762);
and U821 (N_821,N_744,N_718);
xnor U822 (N_822,N_608,N_676);
xnor U823 (N_823,N_754,N_703);
or U824 (N_824,N_729,N_789);
or U825 (N_825,N_755,N_663);
nor U826 (N_826,N_791,N_759);
nor U827 (N_827,N_644,N_623);
and U828 (N_828,N_685,N_691);
nand U829 (N_829,N_638,N_761);
xor U830 (N_830,N_742,N_797);
or U831 (N_831,N_601,N_662);
nor U832 (N_832,N_756,N_613);
xor U833 (N_833,N_757,N_641);
nand U834 (N_834,N_799,N_632);
xor U835 (N_835,N_758,N_604);
and U836 (N_836,N_635,N_787);
xnor U837 (N_837,N_610,N_658);
or U838 (N_838,N_704,N_738);
xor U839 (N_839,N_687,N_722);
nor U840 (N_840,N_740,N_764);
nand U841 (N_841,N_710,N_769);
and U842 (N_842,N_790,N_779);
nor U843 (N_843,N_780,N_636);
and U844 (N_844,N_618,N_681);
nand U845 (N_845,N_743,N_734);
nor U846 (N_846,N_760,N_621);
or U847 (N_847,N_661,N_788);
or U848 (N_848,N_774,N_611);
xor U849 (N_849,N_713,N_715);
nor U850 (N_850,N_747,N_748);
nor U851 (N_851,N_643,N_682);
and U852 (N_852,N_745,N_665);
and U853 (N_853,N_698,N_666);
nand U854 (N_854,N_653,N_794);
nor U855 (N_855,N_778,N_656);
nor U856 (N_856,N_674,N_792);
or U857 (N_857,N_763,N_673);
and U858 (N_858,N_642,N_725);
nand U859 (N_859,N_798,N_773);
nand U860 (N_860,N_629,N_741);
and U861 (N_861,N_692,N_634);
and U862 (N_862,N_669,N_783);
xor U863 (N_863,N_671,N_633);
and U864 (N_864,N_628,N_719);
and U865 (N_865,N_708,N_667);
xnor U866 (N_866,N_684,N_735);
and U867 (N_867,N_782,N_706);
xnor U868 (N_868,N_723,N_606);
or U869 (N_869,N_619,N_786);
xor U870 (N_870,N_614,N_699);
nand U871 (N_871,N_776,N_631);
nor U872 (N_872,N_693,N_672);
nand U873 (N_873,N_620,N_668);
nand U874 (N_874,N_749,N_615);
nand U875 (N_875,N_695,N_731);
nand U876 (N_876,N_600,N_771);
nor U877 (N_877,N_733,N_702);
nand U878 (N_878,N_625,N_647);
nand U879 (N_879,N_766,N_650);
and U880 (N_880,N_690,N_679);
and U881 (N_881,N_677,N_622);
and U882 (N_882,N_796,N_736);
and U883 (N_883,N_616,N_649);
nand U884 (N_884,N_697,N_770);
xor U885 (N_885,N_772,N_720);
xor U886 (N_886,N_659,N_627);
nor U887 (N_887,N_777,N_639);
or U888 (N_888,N_678,N_651);
and U889 (N_889,N_701,N_609);
nand U890 (N_890,N_607,N_688);
or U891 (N_891,N_646,N_675);
and U892 (N_892,N_716,N_775);
nor U893 (N_893,N_767,N_785);
and U894 (N_894,N_626,N_721);
and U895 (N_895,N_670,N_746);
xnor U896 (N_896,N_645,N_752);
and U897 (N_897,N_726,N_728);
and U898 (N_898,N_660,N_654);
xor U899 (N_899,N_648,N_768);
or U900 (N_900,N_773,N_626);
xnor U901 (N_901,N_788,N_664);
nand U902 (N_902,N_756,N_725);
and U903 (N_903,N_622,N_759);
nor U904 (N_904,N_627,N_793);
xor U905 (N_905,N_689,N_768);
or U906 (N_906,N_747,N_611);
nor U907 (N_907,N_786,N_648);
and U908 (N_908,N_739,N_674);
or U909 (N_909,N_698,N_766);
nor U910 (N_910,N_651,N_693);
nor U911 (N_911,N_798,N_752);
nor U912 (N_912,N_780,N_754);
or U913 (N_913,N_734,N_786);
xor U914 (N_914,N_736,N_723);
xor U915 (N_915,N_746,N_695);
nor U916 (N_916,N_641,N_643);
nor U917 (N_917,N_731,N_692);
nor U918 (N_918,N_684,N_646);
and U919 (N_919,N_681,N_699);
xor U920 (N_920,N_649,N_743);
and U921 (N_921,N_768,N_773);
or U922 (N_922,N_708,N_741);
or U923 (N_923,N_777,N_610);
xor U924 (N_924,N_711,N_702);
and U925 (N_925,N_707,N_745);
nand U926 (N_926,N_680,N_667);
or U927 (N_927,N_713,N_663);
nor U928 (N_928,N_678,N_733);
xnor U929 (N_929,N_734,N_797);
xor U930 (N_930,N_666,N_672);
nand U931 (N_931,N_642,N_786);
or U932 (N_932,N_775,N_615);
nand U933 (N_933,N_735,N_620);
xor U934 (N_934,N_701,N_777);
and U935 (N_935,N_762,N_745);
xnor U936 (N_936,N_770,N_642);
and U937 (N_937,N_746,N_728);
xor U938 (N_938,N_626,N_606);
nor U939 (N_939,N_683,N_783);
nor U940 (N_940,N_717,N_798);
and U941 (N_941,N_681,N_731);
xor U942 (N_942,N_710,N_661);
and U943 (N_943,N_650,N_725);
nor U944 (N_944,N_788,N_689);
xnor U945 (N_945,N_635,N_779);
xor U946 (N_946,N_779,N_789);
nand U947 (N_947,N_720,N_780);
xnor U948 (N_948,N_669,N_736);
nand U949 (N_949,N_739,N_720);
nand U950 (N_950,N_687,N_605);
and U951 (N_951,N_776,N_668);
nand U952 (N_952,N_616,N_792);
nor U953 (N_953,N_677,N_620);
nor U954 (N_954,N_622,N_627);
and U955 (N_955,N_693,N_700);
xor U956 (N_956,N_605,N_656);
and U957 (N_957,N_686,N_697);
xnor U958 (N_958,N_794,N_709);
nor U959 (N_959,N_719,N_782);
or U960 (N_960,N_613,N_631);
xnor U961 (N_961,N_768,N_751);
nand U962 (N_962,N_692,N_625);
nand U963 (N_963,N_661,N_658);
xnor U964 (N_964,N_728,N_785);
or U965 (N_965,N_717,N_621);
and U966 (N_966,N_681,N_711);
xnor U967 (N_967,N_762,N_639);
and U968 (N_968,N_618,N_603);
xor U969 (N_969,N_612,N_630);
nand U970 (N_970,N_794,N_607);
or U971 (N_971,N_779,N_759);
and U972 (N_972,N_642,N_766);
and U973 (N_973,N_797,N_765);
nor U974 (N_974,N_769,N_760);
xor U975 (N_975,N_786,N_672);
and U976 (N_976,N_730,N_782);
nand U977 (N_977,N_767,N_717);
and U978 (N_978,N_611,N_622);
xor U979 (N_979,N_617,N_676);
or U980 (N_980,N_653,N_650);
xnor U981 (N_981,N_601,N_696);
and U982 (N_982,N_761,N_609);
nand U983 (N_983,N_639,N_621);
and U984 (N_984,N_708,N_794);
or U985 (N_985,N_766,N_623);
xor U986 (N_986,N_799,N_672);
nor U987 (N_987,N_716,N_701);
nor U988 (N_988,N_676,N_768);
or U989 (N_989,N_799,N_760);
nand U990 (N_990,N_761,N_791);
nand U991 (N_991,N_781,N_798);
xnor U992 (N_992,N_746,N_686);
nand U993 (N_993,N_675,N_609);
xnor U994 (N_994,N_702,N_739);
nand U995 (N_995,N_668,N_651);
nor U996 (N_996,N_608,N_742);
and U997 (N_997,N_790,N_766);
nor U998 (N_998,N_681,N_691);
xor U999 (N_999,N_708,N_770);
xnor U1000 (N_1000,N_958,N_981);
nor U1001 (N_1001,N_943,N_909);
nor U1002 (N_1002,N_835,N_852);
nand U1003 (N_1003,N_833,N_997);
or U1004 (N_1004,N_834,N_971);
or U1005 (N_1005,N_820,N_865);
or U1006 (N_1006,N_923,N_927);
or U1007 (N_1007,N_914,N_829);
or U1008 (N_1008,N_888,N_851);
and U1009 (N_1009,N_926,N_864);
and U1010 (N_1010,N_845,N_942);
or U1011 (N_1011,N_871,N_973);
xnor U1012 (N_1012,N_964,N_920);
xor U1013 (N_1013,N_897,N_823);
nand U1014 (N_1014,N_875,N_953);
nand U1015 (N_1015,N_990,N_806);
xor U1016 (N_1016,N_966,N_947);
nor U1017 (N_1017,N_838,N_861);
xor U1018 (N_1018,N_885,N_972);
and U1019 (N_1019,N_887,N_841);
xnor U1020 (N_1020,N_881,N_969);
and U1021 (N_1021,N_999,N_828);
and U1022 (N_1022,N_917,N_936);
nor U1023 (N_1023,N_886,N_867);
nor U1024 (N_1024,N_975,N_991);
and U1025 (N_1025,N_814,N_911);
and U1026 (N_1026,N_945,N_980);
nor U1027 (N_1027,N_863,N_915);
nand U1028 (N_1028,N_944,N_815);
xnor U1029 (N_1029,N_860,N_869);
or U1030 (N_1030,N_987,N_978);
xnor U1031 (N_1031,N_818,N_849);
nand U1032 (N_1032,N_949,N_846);
xor U1033 (N_1033,N_982,N_921);
xnor U1034 (N_1034,N_847,N_893);
or U1035 (N_1035,N_819,N_922);
nor U1036 (N_1036,N_933,N_977);
and U1037 (N_1037,N_894,N_935);
nand U1038 (N_1038,N_995,N_952);
or U1039 (N_1039,N_839,N_956);
or U1040 (N_1040,N_919,N_850);
nand U1041 (N_1041,N_872,N_928);
nand U1042 (N_1042,N_963,N_810);
or U1043 (N_1043,N_937,N_824);
nor U1044 (N_1044,N_930,N_892);
nand U1045 (N_1045,N_891,N_889);
or U1046 (N_1046,N_900,N_817);
or U1047 (N_1047,N_950,N_811);
nand U1048 (N_1048,N_836,N_998);
xnor U1049 (N_1049,N_859,N_957);
or U1050 (N_1050,N_932,N_837);
and U1051 (N_1051,N_965,N_844);
and U1052 (N_1052,N_902,N_924);
xnor U1053 (N_1053,N_960,N_858);
and U1054 (N_1054,N_882,N_906);
or U1055 (N_1055,N_989,N_821);
nand U1056 (N_1056,N_985,N_855);
or U1057 (N_1057,N_853,N_948);
xor U1058 (N_1058,N_946,N_951);
and U1059 (N_1059,N_918,N_807);
or U1060 (N_1060,N_874,N_994);
nor U1061 (N_1061,N_938,N_934);
or U1062 (N_1062,N_854,N_802);
or U1063 (N_1063,N_848,N_832);
xnor U1064 (N_1064,N_974,N_840);
nand U1065 (N_1065,N_804,N_876);
and U1066 (N_1066,N_968,N_899);
nor U1067 (N_1067,N_822,N_976);
nor U1068 (N_1068,N_940,N_878);
nand U1069 (N_1069,N_929,N_856);
and U1070 (N_1070,N_983,N_842);
xnor U1071 (N_1071,N_907,N_992);
and U1072 (N_1072,N_961,N_913);
xor U1073 (N_1073,N_805,N_941);
and U1074 (N_1074,N_962,N_866);
nand U1075 (N_1075,N_895,N_905);
xor U1076 (N_1076,N_908,N_988);
and U1077 (N_1077,N_883,N_812);
xor U1078 (N_1078,N_862,N_884);
xnor U1079 (N_1079,N_831,N_910);
xor U1080 (N_1080,N_873,N_984);
or U1081 (N_1081,N_931,N_868);
or U1082 (N_1082,N_986,N_890);
or U1083 (N_1083,N_925,N_916);
xor U1084 (N_1084,N_826,N_880);
nand U1085 (N_1085,N_809,N_896);
and U1086 (N_1086,N_803,N_912);
nand U1087 (N_1087,N_993,N_843);
or U1088 (N_1088,N_901,N_830);
or U1089 (N_1089,N_800,N_801);
nand U1090 (N_1090,N_954,N_939);
nor U1091 (N_1091,N_996,N_898);
xor U1092 (N_1092,N_979,N_959);
nand U1093 (N_1093,N_955,N_870);
nor U1094 (N_1094,N_903,N_857);
or U1095 (N_1095,N_879,N_827);
xnor U1096 (N_1096,N_877,N_967);
or U1097 (N_1097,N_816,N_970);
xnor U1098 (N_1098,N_813,N_904);
xor U1099 (N_1099,N_808,N_825);
xor U1100 (N_1100,N_875,N_840);
xor U1101 (N_1101,N_909,N_991);
or U1102 (N_1102,N_926,N_966);
nor U1103 (N_1103,N_860,N_977);
or U1104 (N_1104,N_967,N_917);
nand U1105 (N_1105,N_901,N_846);
nor U1106 (N_1106,N_899,N_943);
xnor U1107 (N_1107,N_865,N_943);
and U1108 (N_1108,N_826,N_818);
nor U1109 (N_1109,N_876,N_969);
xor U1110 (N_1110,N_897,N_942);
or U1111 (N_1111,N_949,N_936);
nor U1112 (N_1112,N_961,N_821);
or U1113 (N_1113,N_858,N_804);
nor U1114 (N_1114,N_993,N_984);
and U1115 (N_1115,N_835,N_888);
or U1116 (N_1116,N_885,N_985);
nor U1117 (N_1117,N_971,N_993);
nor U1118 (N_1118,N_998,N_996);
nor U1119 (N_1119,N_881,N_874);
or U1120 (N_1120,N_854,N_833);
xnor U1121 (N_1121,N_992,N_856);
and U1122 (N_1122,N_881,N_929);
and U1123 (N_1123,N_852,N_831);
or U1124 (N_1124,N_893,N_979);
nand U1125 (N_1125,N_958,N_882);
nand U1126 (N_1126,N_945,N_935);
xnor U1127 (N_1127,N_948,N_914);
or U1128 (N_1128,N_885,N_990);
xor U1129 (N_1129,N_812,N_866);
xor U1130 (N_1130,N_860,N_948);
and U1131 (N_1131,N_937,N_886);
xor U1132 (N_1132,N_922,N_831);
or U1133 (N_1133,N_803,N_836);
or U1134 (N_1134,N_932,N_834);
and U1135 (N_1135,N_807,N_806);
or U1136 (N_1136,N_967,N_975);
nand U1137 (N_1137,N_852,N_930);
xor U1138 (N_1138,N_856,N_944);
nand U1139 (N_1139,N_828,N_853);
xnor U1140 (N_1140,N_993,N_958);
nor U1141 (N_1141,N_859,N_972);
and U1142 (N_1142,N_988,N_845);
xor U1143 (N_1143,N_888,N_983);
xnor U1144 (N_1144,N_900,N_885);
and U1145 (N_1145,N_944,N_951);
nor U1146 (N_1146,N_877,N_912);
xor U1147 (N_1147,N_874,N_946);
xor U1148 (N_1148,N_946,N_819);
xor U1149 (N_1149,N_953,N_879);
or U1150 (N_1150,N_916,N_896);
xor U1151 (N_1151,N_888,N_892);
nor U1152 (N_1152,N_904,N_931);
and U1153 (N_1153,N_878,N_953);
or U1154 (N_1154,N_806,N_853);
xnor U1155 (N_1155,N_984,N_877);
nand U1156 (N_1156,N_809,N_859);
nand U1157 (N_1157,N_859,N_935);
nand U1158 (N_1158,N_895,N_902);
or U1159 (N_1159,N_935,N_829);
or U1160 (N_1160,N_989,N_948);
xor U1161 (N_1161,N_850,N_842);
nand U1162 (N_1162,N_962,N_956);
and U1163 (N_1163,N_842,N_975);
and U1164 (N_1164,N_906,N_811);
xnor U1165 (N_1165,N_882,N_928);
nand U1166 (N_1166,N_818,N_988);
and U1167 (N_1167,N_956,N_866);
nand U1168 (N_1168,N_852,N_998);
xnor U1169 (N_1169,N_956,N_814);
nor U1170 (N_1170,N_915,N_905);
or U1171 (N_1171,N_822,N_845);
xor U1172 (N_1172,N_829,N_870);
nand U1173 (N_1173,N_840,N_997);
or U1174 (N_1174,N_824,N_983);
xnor U1175 (N_1175,N_819,N_950);
nand U1176 (N_1176,N_887,N_901);
and U1177 (N_1177,N_842,N_902);
nand U1178 (N_1178,N_937,N_830);
xor U1179 (N_1179,N_960,N_833);
nand U1180 (N_1180,N_991,N_920);
nand U1181 (N_1181,N_998,N_811);
nor U1182 (N_1182,N_906,N_838);
xnor U1183 (N_1183,N_801,N_940);
xnor U1184 (N_1184,N_831,N_924);
nand U1185 (N_1185,N_820,N_972);
xor U1186 (N_1186,N_847,N_800);
nand U1187 (N_1187,N_863,N_991);
nand U1188 (N_1188,N_965,N_921);
and U1189 (N_1189,N_999,N_931);
or U1190 (N_1190,N_825,N_887);
xor U1191 (N_1191,N_973,N_878);
nand U1192 (N_1192,N_953,N_955);
nand U1193 (N_1193,N_946,N_828);
and U1194 (N_1194,N_877,N_878);
xnor U1195 (N_1195,N_918,N_813);
xor U1196 (N_1196,N_961,N_867);
nand U1197 (N_1197,N_890,N_942);
or U1198 (N_1198,N_972,N_992);
nor U1199 (N_1199,N_921,N_919);
nand U1200 (N_1200,N_1043,N_1125);
nor U1201 (N_1201,N_1081,N_1029);
and U1202 (N_1202,N_1016,N_1187);
or U1203 (N_1203,N_1090,N_1176);
and U1204 (N_1204,N_1002,N_1059);
or U1205 (N_1205,N_1113,N_1158);
or U1206 (N_1206,N_1127,N_1160);
nand U1207 (N_1207,N_1157,N_1198);
and U1208 (N_1208,N_1131,N_1000);
nor U1209 (N_1209,N_1075,N_1183);
or U1210 (N_1210,N_1173,N_1026);
nand U1211 (N_1211,N_1027,N_1119);
xor U1212 (N_1212,N_1118,N_1012);
nor U1213 (N_1213,N_1124,N_1180);
nand U1214 (N_1214,N_1122,N_1069);
or U1215 (N_1215,N_1150,N_1011);
or U1216 (N_1216,N_1193,N_1047);
or U1217 (N_1217,N_1037,N_1022);
and U1218 (N_1218,N_1162,N_1163);
nand U1219 (N_1219,N_1182,N_1100);
or U1220 (N_1220,N_1007,N_1116);
nor U1221 (N_1221,N_1060,N_1080);
nor U1222 (N_1222,N_1067,N_1136);
nand U1223 (N_1223,N_1003,N_1057);
nor U1224 (N_1224,N_1126,N_1139);
or U1225 (N_1225,N_1021,N_1025);
xor U1226 (N_1226,N_1041,N_1145);
or U1227 (N_1227,N_1018,N_1076);
xnor U1228 (N_1228,N_1086,N_1020);
and U1229 (N_1229,N_1005,N_1087);
nand U1230 (N_1230,N_1149,N_1030);
xnor U1231 (N_1231,N_1107,N_1062);
or U1232 (N_1232,N_1077,N_1121);
nor U1233 (N_1233,N_1013,N_1096);
nor U1234 (N_1234,N_1088,N_1009);
or U1235 (N_1235,N_1102,N_1105);
nand U1236 (N_1236,N_1024,N_1031);
nor U1237 (N_1237,N_1190,N_1054);
or U1238 (N_1238,N_1093,N_1074);
nand U1239 (N_1239,N_1103,N_1159);
nand U1240 (N_1240,N_1109,N_1189);
and U1241 (N_1241,N_1194,N_1161);
and U1242 (N_1242,N_1196,N_1171);
nor U1243 (N_1243,N_1128,N_1165);
nor U1244 (N_1244,N_1199,N_1083);
nor U1245 (N_1245,N_1185,N_1138);
nand U1246 (N_1246,N_1004,N_1104);
nor U1247 (N_1247,N_1046,N_1147);
and U1248 (N_1248,N_1049,N_1058);
xor U1249 (N_1249,N_1073,N_1164);
xor U1250 (N_1250,N_1192,N_1040);
xnor U1251 (N_1251,N_1112,N_1170);
xor U1252 (N_1252,N_1061,N_1068);
or U1253 (N_1253,N_1082,N_1063);
nor U1254 (N_1254,N_1177,N_1108);
and U1255 (N_1255,N_1110,N_1172);
and U1256 (N_1256,N_1035,N_1039);
and U1257 (N_1257,N_1079,N_1174);
nor U1258 (N_1258,N_1015,N_1111);
nor U1259 (N_1259,N_1053,N_1168);
nand U1260 (N_1260,N_1144,N_1028);
or U1261 (N_1261,N_1120,N_1038);
and U1262 (N_1262,N_1132,N_1186);
nand U1263 (N_1263,N_1117,N_1123);
nand U1264 (N_1264,N_1091,N_1175);
and U1265 (N_1265,N_1092,N_1006);
nor U1266 (N_1266,N_1056,N_1085);
and U1267 (N_1267,N_1036,N_1048);
nor U1268 (N_1268,N_1179,N_1064);
or U1269 (N_1269,N_1151,N_1010);
nor U1270 (N_1270,N_1089,N_1001);
xor U1271 (N_1271,N_1014,N_1044);
nand U1272 (N_1272,N_1133,N_1034);
nor U1273 (N_1273,N_1072,N_1141);
nand U1274 (N_1274,N_1106,N_1140);
nand U1275 (N_1275,N_1154,N_1181);
and U1276 (N_1276,N_1033,N_1153);
nand U1277 (N_1277,N_1070,N_1071);
and U1278 (N_1278,N_1152,N_1115);
or U1279 (N_1279,N_1019,N_1130);
or U1280 (N_1280,N_1148,N_1042);
nand U1281 (N_1281,N_1101,N_1134);
nand U1282 (N_1282,N_1167,N_1129);
xnor U1283 (N_1283,N_1169,N_1050);
or U1284 (N_1284,N_1094,N_1032);
and U1285 (N_1285,N_1137,N_1052);
nand U1286 (N_1286,N_1097,N_1095);
xor U1287 (N_1287,N_1045,N_1142);
nor U1288 (N_1288,N_1188,N_1051);
or U1289 (N_1289,N_1166,N_1114);
nor U1290 (N_1290,N_1195,N_1184);
nor U1291 (N_1291,N_1065,N_1099);
nor U1292 (N_1292,N_1155,N_1078);
and U1293 (N_1293,N_1143,N_1191);
or U1294 (N_1294,N_1098,N_1055);
nor U1295 (N_1295,N_1135,N_1066);
or U1296 (N_1296,N_1023,N_1008);
nand U1297 (N_1297,N_1084,N_1197);
xor U1298 (N_1298,N_1146,N_1178);
and U1299 (N_1299,N_1156,N_1017);
xnor U1300 (N_1300,N_1110,N_1145);
nand U1301 (N_1301,N_1028,N_1036);
nand U1302 (N_1302,N_1192,N_1162);
or U1303 (N_1303,N_1164,N_1052);
or U1304 (N_1304,N_1112,N_1016);
and U1305 (N_1305,N_1141,N_1011);
and U1306 (N_1306,N_1017,N_1179);
nand U1307 (N_1307,N_1199,N_1165);
or U1308 (N_1308,N_1197,N_1138);
nor U1309 (N_1309,N_1165,N_1179);
or U1310 (N_1310,N_1099,N_1053);
xor U1311 (N_1311,N_1189,N_1120);
nor U1312 (N_1312,N_1000,N_1197);
nand U1313 (N_1313,N_1037,N_1048);
or U1314 (N_1314,N_1048,N_1061);
nor U1315 (N_1315,N_1146,N_1063);
xor U1316 (N_1316,N_1159,N_1167);
nor U1317 (N_1317,N_1166,N_1121);
nor U1318 (N_1318,N_1016,N_1182);
and U1319 (N_1319,N_1144,N_1176);
nor U1320 (N_1320,N_1066,N_1013);
nor U1321 (N_1321,N_1036,N_1150);
xor U1322 (N_1322,N_1086,N_1128);
nand U1323 (N_1323,N_1036,N_1006);
nor U1324 (N_1324,N_1055,N_1190);
and U1325 (N_1325,N_1046,N_1019);
xnor U1326 (N_1326,N_1098,N_1073);
or U1327 (N_1327,N_1075,N_1035);
and U1328 (N_1328,N_1186,N_1064);
nor U1329 (N_1329,N_1185,N_1085);
or U1330 (N_1330,N_1048,N_1189);
nor U1331 (N_1331,N_1160,N_1018);
nor U1332 (N_1332,N_1098,N_1123);
and U1333 (N_1333,N_1039,N_1189);
nor U1334 (N_1334,N_1070,N_1124);
or U1335 (N_1335,N_1047,N_1030);
or U1336 (N_1336,N_1074,N_1100);
nor U1337 (N_1337,N_1031,N_1089);
xnor U1338 (N_1338,N_1161,N_1111);
xnor U1339 (N_1339,N_1073,N_1050);
nor U1340 (N_1340,N_1084,N_1015);
xnor U1341 (N_1341,N_1162,N_1004);
and U1342 (N_1342,N_1135,N_1008);
nand U1343 (N_1343,N_1053,N_1106);
nor U1344 (N_1344,N_1007,N_1057);
and U1345 (N_1345,N_1047,N_1065);
nor U1346 (N_1346,N_1198,N_1174);
or U1347 (N_1347,N_1070,N_1120);
nor U1348 (N_1348,N_1113,N_1142);
nor U1349 (N_1349,N_1023,N_1103);
and U1350 (N_1350,N_1059,N_1157);
xor U1351 (N_1351,N_1082,N_1170);
and U1352 (N_1352,N_1055,N_1143);
or U1353 (N_1353,N_1076,N_1025);
and U1354 (N_1354,N_1126,N_1180);
or U1355 (N_1355,N_1148,N_1019);
and U1356 (N_1356,N_1022,N_1124);
nand U1357 (N_1357,N_1156,N_1123);
xor U1358 (N_1358,N_1022,N_1173);
xor U1359 (N_1359,N_1102,N_1187);
or U1360 (N_1360,N_1073,N_1153);
nand U1361 (N_1361,N_1087,N_1123);
xnor U1362 (N_1362,N_1199,N_1080);
xnor U1363 (N_1363,N_1199,N_1136);
xor U1364 (N_1364,N_1017,N_1060);
nor U1365 (N_1365,N_1017,N_1039);
or U1366 (N_1366,N_1147,N_1044);
xnor U1367 (N_1367,N_1012,N_1053);
xnor U1368 (N_1368,N_1057,N_1138);
xnor U1369 (N_1369,N_1073,N_1006);
nor U1370 (N_1370,N_1001,N_1145);
nor U1371 (N_1371,N_1004,N_1164);
or U1372 (N_1372,N_1146,N_1104);
xnor U1373 (N_1373,N_1069,N_1170);
nor U1374 (N_1374,N_1065,N_1040);
nor U1375 (N_1375,N_1187,N_1087);
or U1376 (N_1376,N_1056,N_1039);
nor U1377 (N_1377,N_1094,N_1130);
or U1378 (N_1378,N_1137,N_1125);
nor U1379 (N_1379,N_1037,N_1146);
nand U1380 (N_1380,N_1177,N_1039);
and U1381 (N_1381,N_1156,N_1190);
nand U1382 (N_1382,N_1178,N_1103);
nand U1383 (N_1383,N_1131,N_1068);
nand U1384 (N_1384,N_1161,N_1132);
or U1385 (N_1385,N_1067,N_1188);
xnor U1386 (N_1386,N_1097,N_1002);
and U1387 (N_1387,N_1150,N_1180);
xor U1388 (N_1388,N_1034,N_1078);
nand U1389 (N_1389,N_1009,N_1001);
or U1390 (N_1390,N_1052,N_1093);
xor U1391 (N_1391,N_1193,N_1189);
nor U1392 (N_1392,N_1189,N_1157);
nand U1393 (N_1393,N_1189,N_1176);
and U1394 (N_1394,N_1073,N_1015);
and U1395 (N_1395,N_1117,N_1191);
or U1396 (N_1396,N_1057,N_1097);
and U1397 (N_1397,N_1078,N_1086);
nor U1398 (N_1398,N_1138,N_1199);
nor U1399 (N_1399,N_1174,N_1085);
xor U1400 (N_1400,N_1384,N_1201);
nor U1401 (N_1401,N_1369,N_1221);
nand U1402 (N_1402,N_1358,N_1223);
and U1403 (N_1403,N_1374,N_1218);
nand U1404 (N_1404,N_1263,N_1236);
xor U1405 (N_1405,N_1210,N_1319);
xor U1406 (N_1406,N_1379,N_1262);
nand U1407 (N_1407,N_1326,N_1303);
and U1408 (N_1408,N_1288,N_1270);
and U1409 (N_1409,N_1284,N_1363);
nor U1410 (N_1410,N_1233,N_1232);
xnor U1411 (N_1411,N_1225,N_1217);
nor U1412 (N_1412,N_1220,N_1304);
nor U1413 (N_1413,N_1327,N_1311);
xor U1414 (N_1414,N_1275,N_1398);
nand U1415 (N_1415,N_1227,N_1360);
xnor U1416 (N_1416,N_1302,N_1299);
xor U1417 (N_1417,N_1213,N_1243);
nor U1418 (N_1418,N_1377,N_1322);
xnor U1419 (N_1419,N_1387,N_1208);
nor U1420 (N_1420,N_1339,N_1224);
or U1421 (N_1421,N_1317,N_1229);
nor U1422 (N_1422,N_1321,N_1200);
xnor U1423 (N_1423,N_1281,N_1372);
or U1424 (N_1424,N_1340,N_1312);
and U1425 (N_1425,N_1249,N_1235);
nor U1426 (N_1426,N_1378,N_1357);
or U1427 (N_1427,N_1399,N_1366);
and U1428 (N_1428,N_1267,N_1202);
and U1429 (N_1429,N_1226,N_1241);
and U1430 (N_1430,N_1301,N_1308);
nand U1431 (N_1431,N_1314,N_1204);
xor U1432 (N_1432,N_1397,N_1300);
xor U1433 (N_1433,N_1257,N_1274);
nand U1434 (N_1434,N_1355,N_1252);
nand U1435 (N_1435,N_1231,N_1367);
or U1436 (N_1436,N_1348,N_1380);
nand U1437 (N_1437,N_1248,N_1253);
and U1438 (N_1438,N_1328,N_1316);
or U1439 (N_1439,N_1365,N_1386);
and U1440 (N_1440,N_1254,N_1359);
nor U1441 (N_1441,N_1395,N_1370);
nor U1442 (N_1442,N_1362,N_1215);
xor U1443 (N_1443,N_1350,N_1272);
or U1444 (N_1444,N_1255,N_1222);
nor U1445 (N_1445,N_1315,N_1342);
nor U1446 (N_1446,N_1216,N_1290);
nor U1447 (N_1447,N_1245,N_1287);
nand U1448 (N_1448,N_1305,N_1376);
or U1449 (N_1449,N_1318,N_1310);
nand U1450 (N_1450,N_1278,N_1391);
or U1451 (N_1451,N_1298,N_1336);
and U1452 (N_1452,N_1256,N_1246);
xnor U1453 (N_1453,N_1335,N_1371);
xnor U1454 (N_1454,N_1268,N_1283);
xnor U1455 (N_1455,N_1206,N_1341);
or U1456 (N_1456,N_1297,N_1334);
or U1457 (N_1457,N_1291,N_1259);
or U1458 (N_1458,N_1237,N_1203);
or U1459 (N_1459,N_1211,N_1289);
and U1460 (N_1460,N_1207,N_1338);
and U1461 (N_1461,N_1205,N_1295);
and U1462 (N_1462,N_1266,N_1389);
nor U1463 (N_1463,N_1209,N_1329);
xor U1464 (N_1464,N_1234,N_1277);
nor U1465 (N_1465,N_1261,N_1242);
nor U1466 (N_1466,N_1347,N_1351);
nor U1467 (N_1467,N_1247,N_1331);
xor U1468 (N_1468,N_1393,N_1219);
nand U1469 (N_1469,N_1282,N_1346);
xnor U1470 (N_1470,N_1368,N_1265);
nand U1471 (N_1471,N_1212,N_1244);
nand U1472 (N_1472,N_1385,N_1324);
and U1473 (N_1473,N_1333,N_1356);
nand U1474 (N_1474,N_1345,N_1375);
and U1475 (N_1475,N_1388,N_1381);
or U1476 (N_1476,N_1264,N_1323);
and U1477 (N_1477,N_1251,N_1293);
nor U1478 (N_1478,N_1309,N_1330);
and U1479 (N_1479,N_1228,N_1344);
nor U1480 (N_1480,N_1390,N_1349);
or U1481 (N_1481,N_1352,N_1238);
or U1482 (N_1482,N_1354,N_1337);
nand U1483 (N_1483,N_1313,N_1364);
or U1484 (N_1484,N_1296,N_1394);
or U1485 (N_1485,N_1286,N_1392);
xnor U1486 (N_1486,N_1332,N_1373);
xor U1487 (N_1487,N_1361,N_1258);
and U1488 (N_1488,N_1325,N_1273);
nand U1489 (N_1489,N_1239,N_1240);
nor U1490 (N_1490,N_1396,N_1306);
nand U1491 (N_1491,N_1230,N_1214);
and U1492 (N_1492,N_1271,N_1294);
or U1493 (N_1493,N_1285,N_1382);
nand U1494 (N_1494,N_1307,N_1383);
xor U1495 (N_1495,N_1292,N_1260);
and U1496 (N_1496,N_1320,N_1276);
nor U1497 (N_1497,N_1250,N_1343);
xor U1498 (N_1498,N_1269,N_1353);
nand U1499 (N_1499,N_1280,N_1279);
nand U1500 (N_1500,N_1353,N_1222);
nand U1501 (N_1501,N_1200,N_1235);
or U1502 (N_1502,N_1399,N_1215);
nor U1503 (N_1503,N_1280,N_1376);
nor U1504 (N_1504,N_1362,N_1201);
nand U1505 (N_1505,N_1351,N_1319);
xnor U1506 (N_1506,N_1306,N_1218);
nor U1507 (N_1507,N_1284,N_1296);
nand U1508 (N_1508,N_1237,N_1338);
nor U1509 (N_1509,N_1326,N_1298);
nor U1510 (N_1510,N_1311,N_1254);
or U1511 (N_1511,N_1381,N_1298);
xnor U1512 (N_1512,N_1350,N_1359);
xor U1513 (N_1513,N_1346,N_1268);
xor U1514 (N_1514,N_1261,N_1399);
xor U1515 (N_1515,N_1267,N_1280);
or U1516 (N_1516,N_1331,N_1371);
or U1517 (N_1517,N_1355,N_1286);
and U1518 (N_1518,N_1334,N_1352);
and U1519 (N_1519,N_1261,N_1285);
or U1520 (N_1520,N_1279,N_1277);
nor U1521 (N_1521,N_1326,N_1227);
or U1522 (N_1522,N_1236,N_1303);
nand U1523 (N_1523,N_1364,N_1344);
xor U1524 (N_1524,N_1309,N_1285);
xor U1525 (N_1525,N_1284,N_1333);
and U1526 (N_1526,N_1230,N_1307);
nand U1527 (N_1527,N_1392,N_1209);
or U1528 (N_1528,N_1232,N_1301);
xor U1529 (N_1529,N_1382,N_1397);
or U1530 (N_1530,N_1368,N_1207);
nor U1531 (N_1531,N_1386,N_1368);
xor U1532 (N_1532,N_1373,N_1258);
xor U1533 (N_1533,N_1285,N_1334);
xor U1534 (N_1534,N_1210,N_1378);
nor U1535 (N_1535,N_1255,N_1246);
and U1536 (N_1536,N_1360,N_1203);
nor U1537 (N_1537,N_1281,N_1246);
and U1538 (N_1538,N_1200,N_1315);
nand U1539 (N_1539,N_1256,N_1315);
and U1540 (N_1540,N_1214,N_1242);
or U1541 (N_1541,N_1364,N_1302);
nor U1542 (N_1542,N_1265,N_1297);
nor U1543 (N_1543,N_1225,N_1270);
xnor U1544 (N_1544,N_1340,N_1391);
xor U1545 (N_1545,N_1395,N_1288);
or U1546 (N_1546,N_1314,N_1349);
xnor U1547 (N_1547,N_1227,N_1338);
or U1548 (N_1548,N_1202,N_1399);
nor U1549 (N_1549,N_1217,N_1329);
and U1550 (N_1550,N_1229,N_1393);
xnor U1551 (N_1551,N_1298,N_1236);
nand U1552 (N_1552,N_1237,N_1395);
and U1553 (N_1553,N_1292,N_1278);
nand U1554 (N_1554,N_1364,N_1392);
nor U1555 (N_1555,N_1329,N_1241);
nand U1556 (N_1556,N_1337,N_1288);
nand U1557 (N_1557,N_1266,N_1210);
nor U1558 (N_1558,N_1386,N_1322);
or U1559 (N_1559,N_1250,N_1365);
xor U1560 (N_1560,N_1317,N_1340);
or U1561 (N_1561,N_1375,N_1349);
or U1562 (N_1562,N_1289,N_1306);
nor U1563 (N_1563,N_1327,N_1217);
xor U1564 (N_1564,N_1307,N_1276);
and U1565 (N_1565,N_1336,N_1326);
nor U1566 (N_1566,N_1321,N_1389);
or U1567 (N_1567,N_1267,N_1223);
xnor U1568 (N_1568,N_1228,N_1390);
nand U1569 (N_1569,N_1313,N_1214);
xor U1570 (N_1570,N_1395,N_1354);
nand U1571 (N_1571,N_1305,N_1370);
nand U1572 (N_1572,N_1388,N_1319);
nand U1573 (N_1573,N_1332,N_1381);
nor U1574 (N_1574,N_1279,N_1215);
and U1575 (N_1575,N_1288,N_1359);
or U1576 (N_1576,N_1359,N_1335);
or U1577 (N_1577,N_1331,N_1360);
or U1578 (N_1578,N_1396,N_1358);
nor U1579 (N_1579,N_1389,N_1288);
or U1580 (N_1580,N_1203,N_1252);
xnor U1581 (N_1581,N_1358,N_1380);
and U1582 (N_1582,N_1297,N_1214);
xor U1583 (N_1583,N_1205,N_1265);
or U1584 (N_1584,N_1351,N_1299);
nand U1585 (N_1585,N_1340,N_1308);
or U1586 (N_1586,N_1397,N_1316);
or U1587 (N_1587,N_1328,N_1336);
xnor U1588 (N_1588,N_1336,N_1214);
or U1589 (N_1589,N_1339,N_1255);
xor U1590 (N_1590,N_1302,N_1304);
nor U1591 (N_1591,N_1298,N_1366);
or U1592 (N_1592,N_1372,N_1379);
nor U1593 (N_1593,N_1316,N_1391);
nand U1594 (N_1594,N_1375,N_1297);
or U1595 (N_1595,N_1288,N_1380);
nor U1596 (N_1596,N_1337,N_1303);
nor U1597 (N_1597,N_1359,N_1237);
nor U1598 (N_1598,N_1282,N_1221);
nor U1599 (N_1599,N_1279,N_1337);
nor U1600 (N_1600,N_1533,N_1461);
or U1601 (N_1601,N_1580,N_1485);
xor U1602 (N_1602,N_1456,N_1573);
nand U1603 (N_1603,N_1570,N_1509);
or U1604 (N_1604,N_1516,N_1511);
nor U1605 (N_1605,N_1527,N_1530);
xnor U1606 (N_1606,N_1434,N_1486);
nor U1607 (N_1607,N_1577,N_1500);
nor U1608 (N_1608,N_1519,N_1507);
nand U1609 (N_1609,N_1465,N_1437);
xnor U1610 (N_1610,N_1459,N_1477);
nand U1611 (N_1611,N_1471,N_1449);
nor U1612 (N_1612,N_1592,N_1402);
and U1613 (N_1613,N_1403,N_1598);
nor U1614 (N_1614,N_1520,N_1421);
and U1615 (N_1615,N_1554,N_1420);
and U1616 (N_1616,N_1529,N_1467);
or U1617 (N_1617,N_1588,N_1413);
or U1618 (N_1618,N_1593,N_1484);
nor U1619 (N_1619,N_1595,N_1487);
or U1620 (N_1620,N_1584,N_1571);
and U1621 (N_1621,N_1526,N_1512);
and U1622 (N_1622,N_1576,N_1599);
xor U1623 (N_1623,N_1425,N_1581);
and U1624 (N_1624,N_1407,N_1452);
xnor U1625 (N_1625,N_1443,N_1586);
xor U1626 (N_1626,N_1522,N_1596);
nand U1627 (N_1627,N_1439,N_1560);
and U1628 (N_1628,N_1513,N_1433);
xnor U1629 (N_1629,N_1545,N_1451);
and U1630 (N_1630,N_1501,N_1400);
and U1631 (N_1631,N_1542,N_1540);
xnor U1632 (N_1632,N_1565,N_1553);
and U1633 (N_1633,N_1503,N_1401);
and U1634 (N_1634,N_1406,N_1438);
nand U1635 (N_1635,N_1585,N_1404);
or U1636 (N_1636,N_1568,N_1492);
xor U1637 (N_1637,N_1502,N_1475);
nor U1638 (N_1638,N_1523,N_1460);
nor U1639 (N_1639,N_1473,N_1478);
nor U1640 (N_1640,N_1422,N_1564);
xnor U1641 (N_1641,N_1440,N_1508);
or U1642 (N_1642,N_1412,N_1441);
nand U1643 (N_1643,N_1423,N_1538);
nand U1644 (N_1644,N_1578,N_1566);
or U1645 (N_1645,N_1532,N_1575);
nor U1646 (N_1646,N_1506,N_1574);
or U1647 (N_1647,N_1408,N_1496);
xor U1648 (N_1648,N_1589,N_1537);
nand U1649 (N_1649,N_1414,N_1510);
and U1650 (N_1650,N_1494,N_1457);
nor U1651 (N_1651,N_1454,N_1432);
nand U1652 (N_1652,N_1488,N_1498);
and U1653 (N_1653,N_1428,N_1405);
or U1654 (N_1654,N_1557,N_1431);
or U1655 (N_1655,N_1481,N_1430);
nand U1656 (N_1656,N_1536,N_1448);
and U1657 (N_1657,N_1582,N_1483);
xnor U1658 (N_1658,N_1479,N_1491);
and U1659 (N_1659,N_1409,N_1505);
or U1660 (N_1660,N_1579,N_1559);
nand U1661 (N_1661,N_1468,N_1569);
or U1662 (N_1662,N_1551,N_1450);
or U1663 (N_1663,N_1525,N_1435);
xnor U1664 (N_1664,N_1495,N_1427);
or U1665 (N_1665,N_1556,N_1535);
and U1666 (N_1666,N_1531,N_1490);
xnor U1667 (N_1667,N_1558,N_1497);
nand U1668 (N_1668,N_1534,N_1499);
xor U1669 (N_1669,N_1447,N_1562);
xnor U1670 (N_1670,N_1539,N_1544);
xor U1671 (N_1671,N_1436,N_1572);
or U1672 (N_1672,N_1547,N_1594);
nand U1673 (N_1673,N_1470,N_1561);
nor U1674 (N_1674,N_1429,N_1445);
nand U1675 (N_1675,N_1583,N_1543);
or U1676 (N_1676,N_1482,N_1517);
and U1677 (N_1677,N_1549,N_1563);
nor U1678 (N_1678,N_1476,N_1541);
nor U1679 (N_1679,N_1472,N_1518);
or U1680 (N_1680,N_1548,N_1591);
nor U1681 (N_1681,N_1410,N_1504);
xor U1682 (N_1682,N_1466,N_1489);
nor U1683 (N_1683,N_1418,N_1493);
nand U1684 (N_1684,N_1528,N_1555);
and U1685 (N_1685,N_1464,N_1416);
xor U1686 (N_1686,N_1426,N_1453);
and U1687 (N_1687,N_1469,N_1480);
nand U1688 (N_1688,N_1552,N_1411);
xor U1689 (N_1689,N_1567,N_1521);
nor U1690 (N_1690,N_1446,N_1442);
or U1691 (N_1691,N_1474,N_1419);
or U1692 (N_1692,N_1597,N_1550);
and U1693 (N_1693,N_1546,N_1587);
nand U1694 (N_1694,N_1415,N_1590);
nor U1695 (N_1695,N_1462,N_1515);
and U1696 (N_1696,N_1444,N_1524);
nand U1697 (N_1697,N_1417,N_1514);
nand U1698 (N_1698,N_1458,N_1455);
nand U1699 (N_1699,N_1463,N_1424);
or U1700 (N_1700,N_1484,N_1499);
nor U1701 (N_1701,N_1416,N_1415);
nand U1702 (N_1702,N_1414,N_1521);
nand U1703 (N_1703,N_1596,N_1425);
xor U1704 (N_1704,N_1467,N_1490);
nor U1705 (N_1705,N_1576,N_1420);
nor U1706 (N_1706,N_1581,N_1584);
xor U1707 (N_1707,N_1431,N_1462);
nand U1708 (N_1708,N_1549,N_1453);
xnor U1709 (N_1709,N_1429,N_1589);
nand U1710 (N_1710,N_1408,N_1472);
xnor U1711 (N_1711,N_1519,N_1548);
xor U1712 (N_1712,N_1548,N_1477);
nor U1713 (N_1713,N_1496,N_1433);
and U1714 (N_1714,N_1487,N_1529);
nand U1715 (N_1715,N_1517,N_1557);
nor U1716 (N_1716,N_1407,N_1598);
nor U1717 (N_1717,N_1532,N_1404);
xnor U1718 (N_1718,N_1576,N_1586);
nand U1719 (N_1719,N_1411,N_1505);
xnor U1720 (N_1720,N_1560,N_1466);
nand U1721 (N_1721,N_1595,N_1580);
nor U1722 (N_1722,N_1492,N_1589);
and U1723 (N_1723,N_1572,N_1575);
nor U1724 (N_1724,N_1481,N_1508);
nor U1725 (N_1725,N_1550,N_1540);
nor U1726 (N_1726,N_1521,N_1477);
nor U1727 (N_1727,N_1428,N_1484);
nor U1728 (N_1728,N_1465,N_1498);
and U1729 (N_1729,N_1438,N_1419);
xnor U1730 (N_1730,N_1419,N_1565);
or U1731 (N_1731,N_1411,N_1490);
nand U1732 (N_1732,N_1460,N_1587);
xor U1733 (N_1733,N_1577,N_1457);
and U1734 (N_1734,N_1467,N_1408);
nand U1735 (N_1735,N_1553,N_1566);
and U1736 (N_1736,N_1529,N_1426);
or U1737 (N_1737,N_1585,N_1426);
nand U1738 (N_1738,N_1454,N_1470);
or U1739 (N_1739,N_1591,N_1468);
and U1740 (N_1740,N_1400,N_1581);
nand U1741 (N_1741,N_1517,N_1591);
nand U1742 (N_1742,N_1513,N_1515);
nand U1743 (N_1743,N_1479,N_1437);
nor U1744 (N_1744,N_1481,N_1407);
and U1745 (N_1745,N_1450,N_1472);
and U1746 (N_1746,N_1596,N_1554);
nor U1747 (N_1747,N_1476,N_1553);
nor U1748 (N_1748,N_1505,N_1446);
nor U1749 (N_1749,N_1588,N_1498);
and U1750 (N_1750,N_1417,N_1494);
or U1751 (N_1751,N_1411,N_1409);
nand U1752 (N_1752,N_1597,N_1593);
or U1753 (N_1753,N_1549,N_1513);
nor U1754 (N_1754,N_1413,N_1537);
nand U1755 (N_1755,N_1539,N_1510);
nand U1756 (N_1756,N_1421,N_1428);
nand U1757 (N_1757,N_1552,N_1502);
nor U1758 (N_1758,N_1543,N_1489);
nand U1759 (N_1759,N_1495,N_1554);
xor U1760 (N_1760,N_1596,N_1597);
nand U1761 (N_1761,N_1486,N_1584);
nand U1762 (N_1762,N_1554,N_1507);
nand U1763 (N_1763,N_1466,N_1564);
nand U1764 (N_1764,N_1458,N_1401);
xnor U1765 (N_1765,N_1425,N_1421);
xor U1766 (N_1766,N_1473,N_1484);
nand U1767 (N_1767,N_1415,N_1405);
and U1768 (N_1768,N_1451,N_1517);
nand U1769 (N_1769,N_1455,N_1471);
nor U1770 (N_1770,N_1545,N_1417);
nor U1771 (N_1771,N_1552,N_1449);
nor U1772 (N_1772,N_1463,N_1559);
and U1773 (N_1773,N_1586,N_1436);
nor U1774 (N_1774,N_1432,N_1473);
nor U1775 (N_1775,N_1547,N_1595);
nor U1776 (N_1776,N_1424,N_1534);
nor U1777 (N_1777,N_1516,N_1564);
nor U1778 (N_1778,N_1511,N_1507);
nor U1779 (N_1779,N_1539,N_1444);
xor U1780 (N_1780,N_1529,N_1517);
and U1781 (N_1781,N_1492,N_1591);
xnor U1782 (N_1782,N_1580,N_1481);
and U1783 (N_1783,N_1526,N_1410);
or U1784 (N_1784,N_1493,N_1545);
nor U1785 (N_1785,N_1556,N_1446);
nor U1786 (N_1786,N_1427,N_1526);
and U1787 (N_1787,N_1433,N_1477);
or U1788 (N_1788,N_1407,N_1421);
xnor U1789 (N_1789,N_1454,N_1506);
and U1790 (N_1790,N_1504,N_1510);
nand U1791 (N_1791,N_1441,N_1514);
nand U1792 (N_1792,N_1520,N_1536);
nand U1793 (N_1793,N_1566,N_1581);
and U1794 (N_1794,N_1473,N_1411);
or U1795 (N_1795,N_1573,N_1599);
or U1796 (N_1796,N_1494,N_1458);
or U1797 (N_1797,N_1400,N_1576);
and U1798 (N_1798,N_1532,N_1590);
nand U1799 (N_1799,N_1590,N_1459);
xnor U1800 (N_1800,N_1639,N_1784);
or U1801 (N_1801,N_1609,N_1753);
nor U1802 (N_1802,N_1642,N_1603);
or U1803 (N_1803,N_1740,N_1649);
nand U1804 (N_1804,N_1617,N_1636);
and U1805 (N_1805,N_1679,N_1678);
nand U1806 (N_1806,N_1608,N_1602);
and U1807 (N_1807,N_1604,N_1702);
or U1808 (N_1808,N_1681,N_1673);
or U1809 (N_1809,N_1721,N_1668);
nand U1810 (N_1810,N_1682,N_1684);
nor U1811 (N_1811,N_1777,N_1764);
nor U1812 (N_1812,N_1700,N_1719);
nand U1813 (N_1813,N_1762,N_1688);
xnor U1814 (N_1814,N_1621,N_1701);
nor U1815 (N_1815,N_1660,N_1683);
or U1816 (N_1816,N_1637,N_1645);
nand U1817 (N_1817,N_1778,N_1779);
nor U1818 (N_1818,N_1686,N_1692);
xnor U1819 (N_1819,N_1780,N_1693);
and U1820 (N_1820,N_1767,N_1723);
or U1821 (N_1821,N_1793,N_1670);
xor U1822 (N_1822,N_1680,N_1694);
nor U1823 (N_1823,N_1651,N_1631);
xnor U1824 (N_1824,N_1755,N_1640);
nor U1825 (N_1825,N_1771,N_1607);
and U1826 (N_1826,N_1796,N_1785);
or U1827 (N_1827,N_1733,N_1695);
nand U1828 (N_1828,N_1648,N_1606);
nor U1829 (N_1829,N_1710,N_1745);
and U1830 (N_1830,N_1671,N_1708);
nor U1831 (N_1831,N_1610,N_1741);
or U1832 (N_1832,N_1716,N_1709);
nand U1833 (N_1833,N_1768,N_1798);
nand U1834 (N_1834,N_1657,N_1748);
or U1835 (N_1835,N_1739,N_1674);
and U1836 (N_1836,N_1687,N_1672);
and U1837 (N_1837,N_1664,N_1799);
or U1838 (N_1838,N_1773,N_1737);
or U1839 (N_1839,N_1794,N_1791);
nor U1840 (N_1840,N_1667,N_1751);
nand U1841 (N_1841,N_1763,N_1792);
nand U1842 (N_1842,N_1783,N_1646);
or U1843 (N_1843,N_1754,N_1725);
or U1844 (N_1844,N_1758,N_1638);
or U1845 (N_1845,N_1628,N_1720);
nand U1846 (N_1846,N_1776,N_1644);
xnor U1847 (N_1847,N_1766,N_1611);
or U1848 (N_1848,N_1635,N_1736);
nor U1849 (N_1849,N_1662,N_1655);
and U1850 (N_1850,N_1600,N_1714);
or U1851 (N_1851,N_1616,N_1759);
and U1852 (N_1852,N_1728,N_1731);
or U1853 (N_1853,N_1724,N_1772);
nand U1854 (N_1854,N_1706,N_1601);
xnor U1855 (N_1855,N_1698,N_1659);
xnor U1856 (N_1856,N_1605,N_1653);
xnor U1857 (N_1857,N_1712,N_1614);
xnor U1858 (N_1858,N_1717,N_1690);
or U1859 (N_1859,N_1761,N_1620);
xnor U1860 (N_1860,N_1626,N_1788);
nand U1861 (N_1861,N_1743,N_1756);
or U1862 (N_1862,N_1623,N_1744);
nand U1863 (N_1863,N_1774,N_1615);
nor U1864 (N_1864,N_1729,N_1752);
and U1865 (N_1865,N_1795,N_1732);
xor U1866 (N_1866,N_1715,N_1691);
nand U1867 (N_1867,N_1749,N_1634);
nand U1868 (N_1868,N_1726,N_1705);
and U1869 (N_1869,N_1654,N_1797);
and U1870 (N_1870,N_1643,N_1656);
nand U1871 (N_1871,N_1632,N_1622);
nand U1872 (N_1872,N_1612,N_1658);
nor U1873 (N_1873,N_1627,N_1689);
xor U1874 (N_1874,N_1630,N_1677);
and U1875 (N_1875,N_1707,N_1713);
nand U1876 (N_1876,N_1730,N_1633);
xnor U1877 (N_1877,N_1727,N_1742);
and U1878 (N_1878,N_1661,N_1722);
or U1879 (N_1879,N_1734,N_1765);
and U1880 (N_1880,N_1747,N_1625);
xnor U1881 (N_1881,N_1613,N_1704);
nand U1882 (N_1882,N_1735,N_1760);
nor U1883 (N_1883,N_1618,N_1696);
or U1884 (N_1884,N_1750,N_1669);
xnor U1885 (N_1885,N_1675,N_1666);
nand U1886 (N_1886,N_1769,N_1787);
and U1887 (N_1887,N_1663,N_1641);
nand U1888 (N_1888,N_1699,N_1738);
or U1889 (N_1889,N_1703,N_1624);
nand U1890 (N_1890,N_1789,N_1746);
nand U1891 (N_1891,N_1697,N_1711);
or U1892 (N_1892,N_1652,N_1786);
xnor U1893 (N_1893,N_1665,N_1782);
nor U1894 (N_1894,N_1619,N_1781);
nor U1895 (N_1895,N_1650,N_1770);
and U1896 (N_1896,N_1718,N_1647);
nor U1897 (N_1897,N_1790,N_1676);
xnor U1898 (N_1898,N_1629,N_1757);
and U1899 (N_1899,N_1775,N_1685);
or U1900 (N_1900,N_1662,N_1785);
xnor U1901 (N_1901,N_1607,N_1726);
nor U1902 (N_1902,N_1684,N_1678);
xnor U1903 (N_1903,N_1647,N_1651);
xnor U1904 (N_1904,N_1674,N_1724);
or U1905 (N_1905,N_1735,N_1726);
nand U1906 (N_1906,N_1744,N_1792);
or U1907 (N_1907,N_1772,N_1615);
xor U1908 (N_1908,N_1664,N_1668);
xor U1909 (N_1909,N_1746,N_1743);
and U1910 (N_1910,N_1789,N_1676);
and U1911 (N_1911,N_1781,N_1739);
or U1912 (N_1912,N_1796,N_1782);
nand U1913 (N_1913,N_1618,N_1643);
and U1914 (N_1914,N_1654,N_1687);
nor U1915 (N_1915,N_1674,N_1641);
xor U1916 (N_1916,N_1703,N_1603);
xor U1917 (N_1917,N_1617,N_1766);
xnor U1918 (N_1918,N_1692,N_1687);
xor U1919 (N_1919,N_1634,N_1636);
xnor U1920 (N_1920,N_1689,N_1761);
nand U1921 (N_1921,N_1616,N_1634);
nor U1922 (N_1922,N_1658,N_1626);
or U1923 (N_1923,N_1715,N_1605);
nor U1924 (N_1924,N_1689,N_1796);
nor U1925 (N_1925,N_1793,N_1790);
or U1926 (N_1926,N_1713,N_1745);
and U1927 (N_1927,N_1643,N_1688);
or U1928 (N_1928,N_1680,N_1697);
and U1929 (N_1929,N_1689,N_1612);
nor U1930 (N_1930,N_1768,N_1710);
or U1931 (N_1931,N_1606,N_1711);
nand U1932 (N_1932,N_1632,N_1657);
nor U1933 (N_1933,N_1764,N_1603);
and U1934 (N_1934,N_1614,N_1640);
nor U1935 (N_1935,N_1766,N_1700);
and U1936 (N_1936,N_1736,N_1723);
nor U1937 (N_1937,N_1797,N_1662);
or U1938 (N_1938,N_1761,N_1639);
and U1939 (N_1939,N_1711,N_1687);
and U1940 (N_1940,N_1663,N_1771);
and U1941 (N_1941,N_1607,N_1695);
and U1942 (N_1942,N_1717,N_1644);
nor U1943 (N_1943,N_1658,N_1669);
xnor U1944 (N_1944,N_1719,N_1756);
nor U1945 (N_1945,N_1690,N_1751);
and U1946 (N_1946,N_1674,N_1686);
xor U1947 (N_1947,N_1691,N_1664);
and U1948 (N_1948,N_1714,N_1720);
xnor U1949 (N_1949,N_1670,N_1717);
and U1950 (N_1950,N_1763,N_1764);
xor U1951 (N_1951,N_1799,N_1733);
or U1952 (N_1952,N_1745,N_1784);
nand U1953 (N_1953,N_1726,N_1700);
nand U1954 (N_1954,N_1621,N_1763);
nand U1955 (N_1955,N_1730,N_1722);
xor U1956 (N_1956,N_1633,N_1615);
or U1957 (N_1957,N_1780,N_1743);
or U1958 (N_1958,N_1671,N_1631);
xor U1959 (N_1959,N_1663,N_1626);
and U1960 (N_1960,N_1656,N_1700);
or U1961 (N_1961,N_1705,N_1658);
and U1962 (N_1962,N_1718,N_1642);
nor U1963 (N_1963,N_1632,N_1778);
nor U1964 (N_1964,N_1641,N_1766);
xnor U1965 (N_1965,N_1756,N_1792);
xor U1966 (N_1966,N_1698,N_1600);
xnor U1967 (N_1967,N_1610,N_1633);
xnor U1968 (N_1968,N_1740,N_1766);
nand U1969 (N_1969,N_1601,N_1682);
or U1970 (N_1970,N_1660,N_1769);
and U1971 (N_1971,N_1796,N_1676);
or U1972 (N_1972,N_1771,N_1649);
and U1973 (N_1973,N_1691,N_1617);
xnor U1974 (N_1974,N_1763,N_1779);
or U1975 (N_1975,N_1631,N_1763);
or U1976 (N_1976,N_1700,N_1608);
xnor U1977 (N_1977,N_1644,N_1631);
nor U1978 (N_1978,N_1607,N_1693);
nor U1979 (N_1979,N_1742,N_1715);
and U1980 (N_1980,N_1766,N_1747);
or U1981 (N_1981,N_1742,N_1695);
or U1982 (N_1982,N_1746,N_1679);
or U1983 (N_1983,N_1773,N_1700);
xnor U1984 (N_1984,N_1604,N_1619);
nor U1985 (N_1985,N_1608,N_1763);
nand U1986 (N_1986,N_1619,N_1756);
nor U1987 (N_1987,N_1686,N_1625);
nor U1988 (N_1988,N_1685,N_1648);
nand U1989 (N_1989,N_1763,N_1701);
or U1990 (N_1990,N_1764,N_1667);
nand U1991 (N_1991,N_1751,N_1642);
nor U1992 (N_1992,N_1728,N_1698);
nor U1993 (N_1993,N_1641,N_1624);
and U1994 (N_1994,N_1698,N_1662);
xor U1995 (N_1995,N_1756,N_1772);
xor U1996 (N_1996,N_1626,N_1744);
and U1997 (N_1997,N_1620,N_1767);
nand U1998 (N_1998,N_1696,N_1771);
or U1999 (N_1999,N_1741,N_1709);
and U2000 (N_2000,N_1861,N_1967);
and U2001 (N_2001,N_1888,N_1892);
nor U2002 (N_2002,N_1994,N_1896);
or U2003 (N_2003,N_1823,N_1927);
nor U2004 (N_2004,N_1824,N_1807);
xnor U2005 (N_2005,N_1884,N_1985);
nand U2006 (N_2006,N_1870,N_1834);
nor U2007 (N_2007,N_1815,N_1862);
and U2008 (N_2008,N_1812,N_1981);
nand U2009 (N_2009,N_1826,N_1960);
or U2010 (N_2010,N_1804,N_1904);
nor U2011 (N_2011,N_1879,N_1928);
xor U2012 (N_2012,N_1808,N_1856);
nand U2013 (N_2013,N_1833,N_1947);
xor U2014 (N_2014,N_1991,N_1800);
and U2015 (N_2015,N_1929,N_1850);
or U2016 (N_2016,N_1940,N_1851);
or U2017 (N_2017,N_1887,N_1934);
or U2018 (N_2018,N_1962,N_1902);
or U2019 (N_2019,N_1933,N_1853);
and U2020 (N_2020,N_1935,N_1974);
or U2021 (N_2021,N_1939,N_1970);
and U2022 (N_2022,N_1945,N_1980);
nor U2023 (N_2023,N_1891,N_1890);
and U2024 (N_2024,N_1844,N_1911);
xnor U2025 (N_2025,N_1941,N_1839);
nor U2026 (N_2026,N_1880,N_1802);
nor U2027 (N_2027,N_1898,N_1825);
nand U2028 (N_2028,N_1924,N_1801);
and U2029 (N_2029,N_1946,N_1822);
and U2030 (N_2030,N_1901,N_1855);
nand U2031 (N_2031,N_1931,N_1835);
nor U2032 (N_2032,N_1920,N_1916);
or U2033 (N_2033,N_1849,N_1936);
nand U2034 (N_2034,N_1882,N_1841);
and U2035 (N_2035,N_1963,N_1984);
nand U2036 (N_2036,N_1836,N_1872);
xnor U2037 (N_2037,N_1909,N_1968);
xnor U2038 (N_2038,N_1978,N_1910);
xnor U2039 (N_2039,N_1877,N_1948);
xnor U2040 (N_2040,N_1952,N_1996);
and U2041 (N_2041,N_1907,N_1846);
nand U2042 (N_2042,N_1806,N_1873);
and U2043 (N_2043,N_1876,N_1831);
nor U2044 (N_2044,N_1866,N_1937);
and U2045 (N_2045,N_1828,N_1938);
or U2046 (N_2046,N_1814,N_1950);
xor U2047 (N_2047,N_1926,N_1982);
or U2048 (N_2048,N_1987,N_1813);
and U2049 (N_2049,N_1976,N_1949);
nor U2050 (N_2050,N_1859,N_1905);
or U2051 (N_2051,N_1990,N_1838);
xor U2052 (N_2052,N_1897,N_1817);
and U2053 (N_2053,N_1914,N_1875);
and U2054 (N_2054,N_1832,N_1958);
xor U2055 (N_2055,N_1821,N_1864);
and U2056 (N_2056,N_1930,N_1899);
nor U2057 (N_2057,N_1969,N_1829);
and U2058 (N_2058,N_1918,N_1925);
or U2059 (N_2059,N_1863,N_1989);
nor U2060 (N_2060,N_1915,N_1874);
and U2061 (N_2061,N_1820,N_1805);
nor U2062 (N_2062,N_1857,N_1965);
xnor U2063 (N_2063,N_1998,N_1852);
nor U2064 (N_2064,N_1913,N_1883);
or U2065 (N_2065,N_1889,N_1971);
or U2066 (N_2066,N_1973,N_1964);
or U2067 (N_2067,N_1830,N_1840);
or U2068 (N_2068,N_1881,N_1919);
nor U2069 (N_2069,N_1810,N_1858);
nand U2070 (N_2070,N_1988,N_1972);
or U2071 (N_2071,N_1959,N_1819);
and U2072 (N_2072,N_1986,N_1908);
and U2073 (N_2073,N_1977,N_1894);
nor U2074 (N_2074,N_1886,N_1803);
xor U2075 (N_2075,N_1921,N_1893);
or U2076 (N_2076,N_1983,N_1837);
and U2077 (N_2077,N_1956,N_1997);
nand U2078 (N_2078,N_1906,N_1818);
or U2079 (N_2079,N_1843,N_1954);
or U2080 (N_2080,N_1979,N_1885);
and U2081 (N_2081,N_1865,N_1942);
nand U2082 (N_2082,N_1912,N_1923);
nor U2083 (N_2083,N_1999,N_1845);
or U2084 (N_2084,N_1903,N_1869);
xor U2085 (N_2085,N_1944,N_1943);
xor U2086 (N_2086,N_1922,N_1953);
or U2087 (N_2087,N_1878,N_1860);
nor U2088 (N_2088,N_1816,N_1955);
nand U2089 (N_2089,N_1809,N_1995);
nor U2090 (N_2090,N_1854,N_1932);
and U2091 (N_2091,N_1811,N_1961);
xnor U2092 (N_2092,N_1847,N_1993);
and U2093 (N_2093,N_1951,N_1917);
nor U2094 (N_2094,N_1966,N_1895);
or U2095 (N_2095,N_1957,N_1900);
nand U2096 (N_2096,N_1827,N_1992);
nor U2097 (N_2097,N_1868,N_1871);
or U2098 (N_2098,N_1867,N_1848);
nor U2099 (N_2099,N_1975,N_1842);
and U2100 (N_2100,N_1878,N_1800);
or U2101 (N_2101,N_1845,N_1980);
nor U2102 (N_2102,N_1947,N_1866);
nand U2103 (N_2103,N_1995,N_1839);
nand U2104 (N_2104,N_1823,N_1828);
xnor U2105 (N_2105,N_1820,N_1825);
and U2106 (N_2106,N_1815,N_1819);
nand U2107 (N_2107,N_1919,N_1871);
xor U2108 (N_2108,N_1874,N_1946);
nand U2109 (N_2109,N_1860,N_1918);
nor U2110 (N_2110,N_1824,N_1929);
xnor U2111 (N_2111,N_1900,N_1923);
nand U2112 (N_2112,N_1882,N_1923);
xnor U2113 (N_2113,N_1947,N_1931);
xor U2114 (N_2114,N_1846,N_1932);
or U2115 (N_2115,N_1942,N_1952);
or U2116 (N_2116,N_1930,N_1882);
nor U2117 (N_2117,N_1843,N_1923);
xnor U2118 (N_2118,N_1928,N_1883);
and U2119 (N_2119,N_1995,N_1829);
and U2120 (N_2120,N_1994,N_1926);
nor U2121 (N_2121,N_1812,N_1886);
nor U2122 (N_2122,N_1906,N_1991);
xor U2123 (N_2123,N_1990,N_1847);
and U2124 (N_2124,N_1954,N_1919);
nor U2125 (N_2125,N_1867,N_1882);
nor U2126 (N_2126,N_1807,N_1814);
xor U2127 (N_2127,N_1921,N_1830);
nand U2128 (N_2128,N_1921,N_1968);
or U2129 (N_2129,N_1829,N_1976);
nor U2130 (N_2130,N_1983,N_1811);
xor U2131 (N_2131,N_1977,N_1987);
xor U2132 (N_2132,N_1953,N_1989);
and U2133 (N_2133,N_1843,N_1984);
nand U2134 (N_2134,N_1806,N_1993);
nor U2135 (N_2135,N_1980,N_1961);
nand U2136 (N_2136,N_1825,N_1878);
xor U2137 (N_2137,N_1901,N_1915);
or U2138 (N_2138,N_1893,N_1980);
and U2139 (N_2139,N_1871,N_1817);
nand U2140 (N_2140,N_1850,N_1857);
and U2141 (N_2141,N_1815,N_1831);
and U2142 (N_2142,N_1878,N_1850);
nor U2143 (N_2143,N_1813,N_1994);
xnor U2144 (N_2144,N_1969,N_1973);
nor U2145 (N_2145,N_1805,N_1836);
nor U2146 (N_2146,N_1876,N_1808);
xnor U2147 (N_2147,N_1942,N_1934);
nor U2148 (N_2148,N_1903,N_1801);
nand U2149 (N_2149,N_1830,N_1963);
xor U2150 (N_2150,N_1958,N_1968);
xor U2151 (N_2151,N_1879,N_1809);
xnor U2152 (N_2152,N_1844,N_1892);
nand U2153 (N_2153,N_1875,N_1954);
nand U2154 (N_2154,N_1828,N_1966);
nor U2155 (N_2155,N_1925,N_1937);
nor U2156 (N_2156,N_1883,N_1805);
nand U2157 (N_2157,N_1847,N_1975);
or U2158 (N_2158,N_1860,N_1909);
nor U2159 (N_2159,N_1919,N_1879);
xnor U2160 (N_2160,N_1827,N_1983);
xnor U2161 (N_2161,N_1947,N_1938);
xnor U2162 (N_2162,N_1847,N_1901);
and U2163 (N_2163,N_1814,N_1993);
and U2164 (N_2164,N_1881,N_1818);
xor U2165 (N_2165,N_1845,N_1835);
nor U2166 (N_2166,N_1947,N_1954);
and U2167 (N_2167,N_1929,N_1938);
xor U2168 (N_2168,N_1966,N_1913);
xnor U2169 (N_2169,N_1801,N_1961);
xor U2170 (N_2170,N_1863,N_1990);
or U2171 (N_2171,N_1866,N_1974);
xnor U2172 (N_2172,N_1982,N_1929);
and U2173 (N_2173,N_1961,N_1890);
nor U2174 (N_2174,N_1902,N_1954);
nor U2175 (N_2175,N_1889,N_1948);
and U2176 (N_2176,N_1941,N_1855);
or U2177 (N_2177,N_1936,N_1870);
nor U2178 (N_2178,N_1981,N_1836);
nor U2179 (N_2179,N_1927,N_1903);
and U2180 (N_2180,N_1951,N_1870);
and U2181 (N_2181,N_1887,N_1877);
nand U2182 (N_2182,N_1810,N_1928);
nand U2183 (N_2183,N_1926,N_1975);
and U2184 (N_2184,N_1983,N_1975);
xnor U2185 (N_2185,N_1846,N_1959);
nor U2186 (N_2186,N_1838,N_1811);
or U2187 (N_2187,N_1988,N_1872);
xor U2188 (N_2188,N_1996,N_1897);
nand U2189 (N_2189,N_1910,N_1919);
nand U2190 (N_2190,N_1887,N_1923);
nor U2191 (N_2191,N_1885,N_1977);
and U2192 (N_2192,N_1923,N_1951);
or U2193 (N_2193,N_1843,N_1998);
nor U2194 (N_2194,N_1923,N_1841);
nand U2195 (N_2195,N_1991,N_1951);
xnor U2196 (N_2196,N_1834,N_1842);
nor U2197 (N_2197,N_1978,N_1964);
nor U2198 (N_2198,N_1845,N_1816);
or U2199 (N_2199,N_1957,N_1925);
or U2200 (N_2200,N_2040,N_2115);
xor U2201 (N_2201,N_2162,N_2139);
xnor U2202 (N_2202,N_2179,N_2062);
xnor U2203 (N_2203,N_2076,N_2079);
or U2204 (N_2204,N_2019,N_2001);
nand U2205 (N_2205,N_2178,N_2156);
xnor U2206 (N_2206,N_2014,N_2083);
nor U2207 (N_2207,N_2145,N_2080);
nand U2208 (N_2208,N_2068,N_2011);
xor U2209 (N_2209,N_2038,N_2097);
or U2210 (N_2210,N_2118,N_2154);
nand U2211 (N_2211,N_2074,N_2129);
or U2212 (N_2212,N_2007,N_2058);
xnor U2213 (N_2213,N_2050,N_2137);
nor U2214 (N_2214,N_2047,N_2123);
nand U2215 (N_2215,N_2167,N_2177);
nand U2216 (N_2216,N_2067,N_2187);
or U2217 (N_2217,N_2122,N_2142);
or U2218 (N_2218,N_2072,N_2091);
nor U2219 (N_2219,N_2052,N_2146);
or U2220 (N_2220,N_2109,N_2099);
and U2221 (N_2221,N_2121,N_2135);
or U2222 (N_2222,N_2039,N_2075);
or U2223 (N_2223,N_2119,N_2150);
and U2224 (N_2224,N_2073,N_2078);
and U2225 (N_2225,N_2153,N_2087);
and U2226 (N_2226,N_2101,N_2172);
xnor U2227 (N_2227,N_2116,N_2157);
nor U2228 (N_2228,N_2026,N_2031);
and U2229 (N_2229,N_2100,N_2161);
nor U2230 (N_2230,N_2148,N_2042);
nand U2231 (N_2231,N_2029,N_2032);
or U2232 (N_2232,N_2124,N_2034);
and U2233 (N_2233,N_2166,N_2009);
nand U2234 (N_2234,N_2183,N_2090);
nor U2235 (N_2235,N_2192,N_2176);
nand U2236 (N_2236,N_2188,N_2071);
or U2237 (N_2237,N_2095,N_2195);
or U2238 (N_2238,N_2065,N_2094);
or U2239 (N_2239,N_2063,N_2189);
nand U2240 (N_2240,N_2168,N_2184);
and U2241 (N_2241,N_2193,N_2046);
nor U2242 (N_2242,N_2171,N_2117);
xnor U2243 (N_2243,N_2155,N_2030);
or U2244 (N_2244,N_2021,N_2133);
and U2245 (N_2245,N_2023,N_2000);
nand U2246 (N_2246,N_2085,N_2160);
nand U2247 (N_2247,N_2066,N_2015);
and U2248 (N_2248,N_2103,N_2158);
nand U2249 (N_2249,N_2170,N_2060);
nand U2250 (N_2250,N_2084,N_2152);
and U2251 (N_2251,N_2044,N_2131);
nand U2252 (N_2252,N_2104,N_2125);
and U2253 (N_2253,N_2141,N_2092);
and U2254 (N_2254,N_2082,N_2036);
nor U2255 (N_2255,N_2012,N_2182);
nor U2256 (N_2256,N_2081,N_2008);
and U2257 (N_2257,N_2037,N_2165);
and U2258 (N_2258,N_2024,N_2089);
and U2259 (N_2259,N_2173,N_2175);
nand U2260 (N_2260,N_2106,N_2028);
and U2261 (N_2261,N_2169,N_2061);
xnor U2262 (N_2262,N_2136,N_2196);
and U2263 (N_2263,N_2191,N_2113);
nor U2264 (N_2264,N_2102,N_2041);
nor U2265 (N_2265,N_2056,N_2064);
and U2266 (N_2266,N_2017,N_2107);
xor U2267 (N_2267,N_2051,N_2143);
and U2268 (N_2268,N_2186,N_2088);
and U2269 (N_2269,N_2002,N_2004);
nor U2270 (N_2270,N_2053,N_2132);
and U2271 (N_2271,N_2027,N_2174);
or U2272 (N_2272,N_2096,N_2144);
xnor U2273 (N_2273,N_2151,N_2006);
and U2274 (N_2274,N_2098,N_2020);
and U2275 (N_2275,N_2190,N_2126);
nand U2276 (N_2276,N_2057,N_2093);
and U2277 (N_2277,N_2185,N_2045);
xor U2278 (N_2278,N_2110,N_2018);
nand U2279 (N_2279,N_2086,N_2180);
xor U2280 (N_2280,N_2055,N_2069);
xor U2281 (N_2281,N_2105,N_2181);
and U2282 (N_2282,N_2070,N_2159);
nor U2283 (N_2283,N_2049,N_2164);
or U2284 (N_2284,N_2134,N_2003);
nand U2285 (N_2285,N_2043,N_2048);
nand U2286 (N_2286,N_2054,N_2120);
nor U2287 (N_2287,N_2033,N_2077);
nor U2288 (N_2288,N_2140,N_2163);
nor U2289 (N_2289,N_2059,N_2194);
and U2290 (N_2290,N_2013,N_2130);
nor U2291 (N_2291,N_2010,N_2138);
and U2292 (N_2292,N_2149,N_2005);
and U2293 (N_2293,N_2111,N_2112);
nor U2294 (N_2294,N_2114,N_2108);
or U2295 (N_2295,N_2025,N_2035);
xnor U2296 (N_2296,N_2022,N_2198);
and U2297 (N_2297,N_2147,N_2127);
or U2298 (N_2298,N_2128,N_2199);
or U2299 (N_2299,N_2016,N_2197);
or U2300 (N_2300,N_2162,N_2145);
or U2301 (N_2301,N_2120,N_2022);
and U2302 (N_2302,N_2138,N_2089);
xor U2303 (N_2303,N_2098,N_2140);
and U2304 (N_2304,N_2071,N_2041);
or U2305 (N_2305,N_2055,N_2050);
and U2306 (N_2306,N_2113,N_2044);
and U2307 (N_2307,N_2056,N_2083);
and U2308 (N_2308,N_2154,N_2193);
or U2309 (N_2309,N_2064,N_2071);
or U2310 (N_2310,N_2148,N_2068);
and U2311 (N_2311,N_2101,N_2141);
and U2312 (N_2312,N_2188,N_2120);
nand U2313 (N_2313,N_2033,N_2024);
or U2314 (N_2314,N_2145,N_2045);
nand U2315 (N_2315,N_2194,N_2004);
nor U2316 (N_2316,N_2114,N_2124);
nor U2317 (N_2317,N_2196,N_2131);
nor U2318 (N_2318,N_2003,N_2015);
or U2319 (N_2319,N_2086,N_2159);
and U2320 (N_2320,N_2190,N_2176);
xor U2321 (N_2321,N_2059,N_2100);
nor U2322 (N_2322,N_2112,N_2126);
xnor U2323 (N_2323,N_2198,N_2115);
and U2324 (N_2324,N_2034,N_2110);
or U2325 (N_2325,N_2051,N_2108);
nand U2326 (N_2326,N_2160,N_2127);
or U2327 (N_2327,N_2030,N_2047);
nor U2328 (N_2328,N_2114,N_2167);
and U2329 (N_2329,N_2043,N_2037);
and U2330 (N_2330,N_2179,N_2118);
and U2331 (N_2331,N_2073,N_2150);
and U2332 (N_2332,N_2020,N_2162);
and U2333 (N_2333,N_2073,N_2146);
or U2334 (N_2334,N_2101,N_2105);
nor U2335 (N_2335,N_2077,N_2195);
or U2336 (N_2336,N_2161,N_2091);
and U2337 (N_2337,N_2112,N_2002);
or U2338 (N_2338,N_2032,N_2190);
or U2339 (N_2339,N_2175,N_2052);
nor U2340 (N_2340,N_2112,N_2182);
nand U2341 (N_2341,N_2151,N_2145);
or U2342 (N_2342,N_2026,N_2067);
and U2343 (N_2343,N_2054,N_2198);
xor U2344 (N_2344,N_2119,N_2137);
and U2345 (N_2345,N_2197,N_2188);
or U2346 (N_2346,N_2152,N_2194);
nor U2347 (N_2347,N_2010,N_2102);
nor U2348 (N_2348,N_2105,N_2090);
and U2349 (N_2349,N_2130,N_2046);
nand U2350 (N_2350,N_2001,N_2177);
nand U2351 (N_2351,N_2090,N_2157);
nand U2352 (N_2352,N_2102,N_2061);
or U2353 (N_2353,N_2042,N_2179);
or U2354 (N_2354,N_2068,N_2082);
nor U2355 (N_2355,N_2187,N_2100);
or U2356 (N_2356,N_2146,N_2176);
xnor U2357 (N_2357,N_2063,N_2004);
or U2358 (N_2358,N_2011,N_2166);
or U2359 (N_2359,N_2155,N_2121);
nor U2360 (N_2360,N_2010,N_2041);
and U2361 (N_2361,N_2151,N_2175);
nor U2362 (N_2362,N_2168,N_2149);
and U2363 (N_2363,N_2073,N_2076);
and U2364 (N_2364,N_2018,N_2172);
nor U2365 (N_2365,N_2057,N_2129);
or U2366 (N_2366,N_2198,N_2021);
xnor U2367 (N_2367,N_2044,N_2145);
or U2368 (N_2368,N_2119,N_2181);
nand U2369 (N_2369,N_2000,N_2144);
nand U2370 (N_2370,N_2002,N_2150);
nand U2371 (N_2371,N_2052,N_2114);
xnor U2372 (N_2372,N_2173,N_2129);
or U2373 (N_2373,N_2119,N_2067);
xnor U2374 (N_2374,N_2009,N_2099);
or U2375 (N_2375,N_2039,N_2005);
nor U2376 (N_2376,N_2082,N_2014);
nand U2377 (N_2377,N_2167,N_2003);
and U2378 (N_2378,N_2079,N_2026);
nand U2379 (N_2379,N_2170,N_2091);
nor U2380 (N_2380,N_2021,N_2185);
nor U2381 (N_2381,N_2194,N_2032);
and U2382 (N_2382,N_2053,N_2074);
or U2383 (N_2383,N_2003,N_2165);
nand U2384 (N_2384,N_2040,N_2179);
and U2385 (N_2385,N_2182,N_2020);
and U2386 (N_2386,N_2105,N_2133);
nand U2387 (N_2387,N_2098,N_2108);
nor U2388 (N_2388,N_2079,N_2126);
and U2389 (N_2389,N_2134,N_2169);
and U2390 (N_2390,N_2087,N_2143);
or U2391 (N_2391,N_2072,N_2041);
and U2392 (N_2392,N_2010,N_2062);
or U2393 (N_2393,N_2046,N_2191);
or U2394 (N_2394,N_2006,N_2115);
nor U2395 (N_2395,N_2005,N_2115);
and U2396 (N_2396,N_2128,N_2026);
nand U2397 (N_2397,N_2022,N_2034);
xor U2398 (N_2398,N_2112,N_2157);
xnor U2399 (N_2399,N_2128,N_2108);
nand U2400 (N_2400,N_2220,N_2218);
and U2401 (N_2401,N_2270,N_2304);
nand U2402 (N_2402,N_2299,N_2319);
or U2403 (N_2403,N_2374,N_2228);
and U2404 (N_2404,N_2307,N_2350);
and U2405 (N_2405,N_2278,N_2372);
xnor U2406 (N_2406,N_2225,N_2296);
and U2407 (N_2407,N_2236,N_2370);
or U2408 (N_2408,N_2398,N_2366);
nand U2409 (N_2409,N_2262,N_2314);
xnor U2410 (N_2410,N_2362,N_2308);
xnor U2411 (N_2411,N_2338,N_2271);
nand U2412 (N_2412,N_2323,N_2301);
nor U2413 (N_2413,N_2238,N_2223);
and U2414 (N_2414,N_2325,N_2283);
or U2415 (N_2415,N_2332,N_2349);
or U2416 (N_2416,N_2231,N_2356);
xnor U2417 (N_2417,N_2335,N_2254);
or U2418 (N_2418,N_2293,N_2295);
or U2419 (N_2419,N_2294,N_2206);
nand U2420 (N_2420,N_2333,N_2336);
or U2421 (N_2421,N_2290,N_2397);
and U2422 (N_2422,N_2392,N_2240);
and U2423 (N_2423,N_2205,N_2217);
and U2424 (N_2424,N_2352,N_2327);
or U2425 (N_2425,N_2277,N_2306);
xnor U2426 (N_2426,N_2354,N_2367);
or U2427 (N_2427,N_2256,N_2250);
xnor U2428 (N_2428,N_2212,N_2235);
nand U2429 (N_2429,N_2341,N_2221);
or U2430 (N_2430,N_2251,N_2382);
nand U2431 (N_2431,N_2395,N_2259);
nand U2432 (N_2432,N_2275,N_2269);
nand U2433 (N_2433,N_2320,N_2245);
and U2434 (N_2434,N_2313,N_2285);
nor U2435 (N_2435,N_2364,N_2329);
xor U2436 (N_2436,N_2318,N_2234);
or U2437 (N_2437,N_2286,N_2342);
or U2438 (N_2438,N_2331,N_2334);
or U2439 (N_2439,N_2303,N_2317);
nor U2440 (N_2440,N_2389,N_2288);
nor U2441 (N_2441,N_2222,N_2312);
xor U2442 (N_2442,N_2263,N_2207);
nor U2443 (N_2443,N_2209,N_2266);
or U2444 (N_2444,N_2226,N_2339);
nand U2445 (N_2445,N_2261,N_2249);
nor U2446 (N_2446,N_2363,N_2343);
nor U2447 (N_2447,N_2227,N_2388);
nand U2448 (N_2448,N_2345,N_2368);
and U2449 (N_2449,N_2242,N_2369);
xor U2450 (N_2450,N_2280,N_2380);
nand U2451 (N_2451,N_2287,N_2383);
xnor U2452 (N_2452,N_2219,N_2322);
nor U2453 (N_2453,N_2360,N_2276);
or U2454 (N_2454,N_2201,N_2321);
or U2455 (N_2455,N_2361,N_2371);
xor U2456 (N_2456,N_2378,N_2233);
and U2457 (N_2457,N_2381,N_2309);
nor U2458 (N_2458,N_2291,N_2255);
xor U2459 (N_2459,N_2391,N_2272);
xor U2460 (N_2460,N_2365,N_2328);
nand U2461 (N_2461,N_2337,N_2316);
nand U2462 (N_2462,N_2253,N_2340);
nand U2463 (N_2463,N_2359,N_2265);
nand U2464 (N_2464,N_2330,N_2279);
nor U2465 (N_2465,N_2284,N_2292);
nand U2466 (N_2466,N_2200,N_2257);
nand U2467 (N_2467,N_2208,N_2274);
or U2468 (N_2468,N_2230,N_2347);
nand U2469 (N_2469,N_2213,N_2305);
and U2470 (N_2470,N_2224,N_2210);
nor U2471 (N_2471,N_2373,N_2258);
nor U2472 (N_2472,N_2204,N_2282);
xnor U2473 (N_2473,N_2229,N_2300);
and U2474 (N_2474,N_2376,N_2289);
xnor U2475 (N_2475,N_2248,N_2311);
or U2476 (N_2476,N_2241,N_2346);
xor U2477 (N_2477,N_2353,N_2390);
xnor U2478 (N_2478,N_2246,N_2237);
nor U2479 (N_2479,N_2281,N_2232);
and U2480 (N_2480,N_2247,N_2267);
and U2481 (N_2481,N_2244,N_2399);
and U2482 (N_2482,N_2302,N_2252);
and U2483 (N_2483,N_2298,N_2211);
or U2484 (N_2484,N_2351,N_2375);
or U2485 (N_2485,N_2214,N_2387);
and U2486 (N_2486,N_2396,N_2310);
nor U2487 (N_2487,N_2273,N_2324);
or U2488 (N_2488,N_2358,N_2315);
xor U2489 (N_2489,N_2239,N_2384);
nor U2490 (N_2490,N_2377,N_2268);
xnor U2491 (N_2491,N_2348,N_2379);
or U2492 (N_2492,N_2355,N_2326);
or U2493 (N_2493,N_2357,N_2297);
or U2494 (N_2494,N_2394,N_2393);
and U2495 (N_2495,N_2202,N_2203);
nand U2496 (N_2496,N_2264,N_2385);
nand U2497 (N_2497,N_2243,N_2215);
and U2498 (N_2498,N_2344,N_2260);
xnor U2499 (N_2499,N_2216,N_2386);
and U2500 (N_2500,N_2371,N_2341);
nor U2501 (N_2501,N_2313,N_2265);
or U2502 (N_2502,N_2236,N_2376);
or U2503 (N_2503,N_2257,N_2215);
nor U2504 (N_2504,N_2337,N_2365);
nand U2505 (N_2505,N_2229,N_2277);
xor U2506 (N_2506,N_2393,N_2313);
or U2507 (N_2507,N_2397,N_2270);
and U2508 (N_2508,N_2258,N_2328);
nor U2509 (N_2509,N_2398,N_2218);
or U2510 (N_2510,N_2204,N_2260);
and U2511 (N_2511,N_2240,N_2278);
xnor U2512 (N_2512,N_2236,N_2373);
or U2513 (N_2513,N_2398,N_2284);
nor U2514 (N_2514,N_2287,N_2204);
xor U2515 (N_2515,N_2291,N_2387);
xor U2516 (N_2516,N_2368,N_2203);
nor U2517 (N_2517,N_2383,N_2326);
nor U2518 (N_2518,N_2370,N_2302);
xor U2519 (N_2519,N_2399,N_2287);
nand U2520 (N_2520,N_2317,N_2339);
xor U2521 (N_2521,N_2350,N_2265);
xnor U2522 (N_2522,N_2232,N_2296);
and U2523 (N_2523,N_2385,N_2241);
or U2524 (N_2524,N_2275,N_2392);
or U2525 (N_2525,N_2348,N_2367);
or U2526 (N_2526,N_2386,N_2242);
or U2527 (N_2527,N_2256,N_2221);
and U2528 (N_2528,N_2363,N_2288);
xor U2529 (N_2529,N_2396,N_2323);
or U2530 (N_2530,N_2347,N_2273);
nand U2531 (N_2531,N_2378,N_2351);
nor U2532 (N_2532,N_2258,N_2226);
and U2533 (N_2533,N_2325,N_2209);
xor U2534 (N_2534,N_2273,N_2346);
nand U2535 (N_2535,N_2389,N_2280);
and U2536 (N_2536,N_2374,N_2245);
and U2537 (N_2537,N_2346,N_2208);
and U2538 (N_2538,N_2368,N_2282);
or U2539 (N_2539,N_2359,N_2209);
nor U2540 (N_2540,N_2367,N_2369);
nor U2541 (N_2541,N_2357,N_2372);
xor U2542 (N_2542,N_2399,N_2275);
xnor U2543 (N_2543,N_2215,N_2286);
and U2544 (N_2544,N_2384,N_2211);
xor U2545 (N_2545,N_2372,N_2268);
nor U2546 (N_2546,N_2304,N_2303);
xor U2547 (N_2547,N_2350,N_2351);
and U2548 (N_2548,N_2212,N_2256);
nand U2549 (N_2549,N_2354,N_2280);
and U2550 (N_2550,N_2289,N_2353);
nand U2551 (N_2551,N_2323,N_2356);
nor U2552 (N_2552,N_2379,N_2394);
nor U2553 (N_2553,N_2303,N_2232);
or U2554 (N_2554,N_2394,N_2332);
and U2555 (N_2555,N_2294,N_2388);
xnor U2556 (N_2556,N_2285,N_2364);
nand U2557 (N_2557,N_2229,N_2279);
or U2558 (N_2558,N_2283,N_2297);
or U2559 (N_2559,N_2302,N_2301);
nor U2560 (N_2560,N_2200,N_2213);
nor U2561 (N_2561,N_2333,N_2210);
nor U2562 (N_2562,N_2320,N_2219);
xor U2563 (N_2563,N_2214,N_2378);
nor U2564 (N_2564,N_2200,N_2397);
and U2565 (N_2565,N_2294,N_2392);
nand U2566 (N_2566,N_2240,N_2324);
nor U2567 (N_2567,N_2391,N_2364);
and U2568 (N_2568,N_2264,N_2295);
xor U2569 (N_2569,N_2363,N_2284);
xnor U2570 (N_2570,N_2378,N_2213);
and U2571 (N_2571,N_2383,N_2272);
or U2572 (N_2572,N_2303,N_2250);
and U2573 (N_2573,N_2260,N_2371);
and U2574 (N_2574,N_2355,N_2212);
nor U2575 (N_2575,N_2242,N_2285);
or U2576 (N_2576,N_2223,N_2215);
xor U2577 (N_2577,N_2260,N_2298);
and U2578 (N_2578,N_2381,N_2312);
nor U2579 (N_2579,N_2224,N_2226);
nor U2580 (N_2580,N_2325,N_2381);
or U2581 (N_2581,N_2206,N_2299);
nor U2582 (N_2582,N_2360,N_2349);
and U2583 (N_2583,N_2279,N_2336);
and U2584 (N_2584,N_2363,N_2364);
xor U2585 (N_2585,N_2324,N_2369);
and U2586 (N_2586,N_2382,N_2355);
nand U2587 (N_2587,N_2362,N_2241);
xnor U2588 (N_2588,N_2331,N_2207);
xor U2589 (N_2589,N_2215,N_2350);
xor U2590 (N_2590,N_2206,N_2293);
nor U2591 (N_2591,N_2343,N_2315);
xor U2592 (N_2592,N_2355,N_2302);
nor U2593 (N_2593,N_2394,N_2330);
nor U2594 (N_2594,N_2384,N_2344);
nand U2595 (N_2595,N_2307,N_2274);
and U2596 (N_2596,N_2390,N_2221);
or U2597 (N_2597,N_2313,N_2270);
and U2598 (N_2598,N_2387,N_2320);
and U2599 (N_2599,N_2318,N_2389);
and U2600 (N_2600,N_2466,N_2468);
or U2601 (N_2601,N_2498,N_2469);
or U2602 (N_2602,N_2513,N_2594);
nand U2603 (N_2603,N_2534,N_2518);
nor U2604 (N_2604,N_2579,N_2517);
xnor U2605 (N_2605,N_2436,N_2522);
or U2606 (N_2606,N_2561,N_2489);
and U2607 (N_2607,N_2559,N_2543);
and U2608 (N_2608,N_2593,N_2526);
nand U2609 (N_2609,N_2463,N_2500);
nor U2610 (N_2610,N_2512,N_2490);
or U2611 (N_2611,N_2519,N_2524);
xnor U2612 (N_2612,N_2556,N_2516);
nor U2613 (N_2613,N_2442,N_2525);
or U2614 (N_2614,N_2584,N_2426);
and U2615 (N_2615,N_2486,N_2465);
nor U2616 (N_2616,N_2562,N_2434);
nor U2617 (N_2617,N_2550,N_2470);
xnor U2618 (N_2618,N_2406,N_2422);
and U2619 (N_2619,N_2503,N_2440);
nor U2620 (N_2620,N_2402,N_2458);
or U2621 (N_2621,N_2427,N_2464);
nor U2622 (N_2622,N_2551,N_2501);
xnor U2623 (N_2623,N_2557,N_2407);
nand U2624 (N_2624,N_2529,N_2587);
and U2625 (N_2625,N_2541,N_2493);
or U2626 (N_2626,N_2453,N_2497);
nor U2627 (N_2627,N_2438,N_2437);
nand U2628 (N_2628,N_2445,N_2510);
or U2629 (N_2629,N_2549,N_2590);
or U2630 (N_2630,N_2456,N_2571);
xnor U2631 (N_2631,N_2539,N_2449);
or U2632 (N_2632,N_2491,N_2425);
and U2633 (N_2633,N_2573,N_2467);
xor U2634 (N_2634,N_2531,N_2408);
or U2635 (N_2635,N_2574,N_2419);
and U2636 (N_2636,N_2448,N_2570);
or U2637 (N_2637,N_2599,N_2569);
nor U2638 (N_2638,N_2576,N_2568);
xnor U2639 (N_2639,N_2495,N_2589);
and U2640 (N_2640,N_2476,N_2588);
xor U2641 (N_2641,N_2554,N_2401);
or U2642 (N_2642,N_2563,N_2509);
and U2643 (N_2643,N_2454,N_2450);
xor U2644 (N_2644,N_2578,N_2537);
and U2645 (N_2645,N_2462,N_2542);
xnor U2646 (N_2646,N_2403,N_2487);
and U2647 (N_2647,N_2560,N_2591);
and U2648 (N_2648,N_2478,N_2428);
or U2649 (N_2649,N_2443,N_2474);
xnor U2650 (N_2650,N_2553,N_2484);
nand U2651 (N_2651,N_2488,N_2405);
nand U2652 (N_2652,N_2528,N_2548);
nand U2653 (N_2653,N_2429,N_2400);
and U2654 (N_2654,N_2418,N_2496);
and U2655 (N_2655,N_2455,N_2567);
nor U2656 (N_2656,N_2546,N_2430);
nand U2657 (N_2657,N_2439,N_2552);
and U2658 (N_2658,N_2461,N_2414);
and U2659 (N_2659,N_2547,N_2582);
and U2660 (N_2660,N_2592,N_2564);
nand U2661 (N_2661,N_2499,N_2535);
or U2662 (N_2662,N_2451,N_2420);
nor U2663 (N_2663,N_2521,N_2572);
or U2664 (N_2664,N_2480,N_2411);
or U2665 (N_2665,N_2412,N_2515);
nand U2666 (N_2666,N_2502,N_2410);
nor U2667 (N_2667,N_2597,N_2404);
nand U2668 (N_2668,N_2540,N_2417);
and U2669 (N_2669,N_2505,N_2585);
and U2670 (N_2670,N_2504,N_2533);
nor U2671 (N_2671,N_2581,N_2508);
and U2672 (N_2672,N_2506,N_2477);
or U2673 (N_2673,N_2566,N_2536);
and U2674 (N_2674,N_2441,N_2523);
xnor U2675 (N_2675,N_2527,N_2416);
nand U2676 (N_2676,N_2596,N_2479);
xnor U2677 (N_2677,N_2583,N_2424);
and U2678 (N_2678,N_2460,N_2485);
and U2679 (N_2679,N_2409,N_2457);
xnor U2680 (N_2680,N_2575,N_2483);
and U2681 (N_2681,N_2444,N_2514);
nor U2682 (N_2682,N_2447,N_2481);
or U2683 (N_2683,N_2595,N_2482);
or U2684 (N_2684,N_2530,N_2471);
xnor U2685 (N_2685,N_2473,N_2431);
or U2686 (N_2686,N_2492,N_2494);
xor U2687 (N_2687,N_2413,N_2459);
and U2688 (N_2688,N_2520,N_2475);
and U2689 (N_2689,N_2544,N_2586);
nand U2690 (N_2690,N_2580,N_2565);
nor U2691 (N_2691,N_2452,N_2511);
xnor U2692 (N_2692,N_2545,N_2555);
and U2693 (N_2693,N_2507,N_2472);
and U2694 (N_2694,N_2532,N_2446);
and U2695 (N_2695,N_2598,N_2433);
nor U2696 (N_2696,N_2415,N_2558);
nand U2697 (N_2697,N_2577,N_2432);
xnor U2698 (N_2698,N_2435,N_2423);
nand U2699 (N_2699,N_2538,N_2421);
and U2700 (N_2700,N_2590,N_2571);
and U2701 (N_2701,N_2412,N_2466);
nand U2702 (N_2702,N_2439,N_2505);
nor U2703 (N_2703,N_2428,N_2496);
and U2704 (N_2704,N_2445,N_2575);
nor U2705 (N_2705,N_2576,N_2532);
or U2706 (N_2706,N_2495,N_2563);
or U2707 (N_2707,N_2543,N_2592);
and U2708 (N_2708,N_2470,N_2546);
or U2709 (N_2709,N_2400,N_2439);
or U2710 (N_2710,N_2455,N_2554);
or U2711 (N_2711,N_2500,N_2537);
nand U2712 (N_2712,N_2421,N_2597);
nand U2713 (N_2713,N_2598,N_2595);
nand U2714 (N_2714,N_2424,N_2550);
or U2715 (N_2715,N_2518,N_2521);
xnor U2716 (N_2716,N_2506,N_2574);
nand U2717 (N_2717,N_2575,N_2507);
or U2718 (N_2718,N_2405,N_2422);
nand U2719 (N_2719,N_2458,N_2544);
nand U2720 (N_2720,N_2580,N_2540);
xnor U2721 (N_2721,N_2585,N_2550);
nor U2722 (N_2722,N_2585,N_2544);
nor U2723 (N_2723,N_2533,N_2549);
nor U2724 (N_2724,N_2548,N_2507);
or U2725 (N_2725,N_2550,N_2512);
or U2726 (N_2726,N_2414,N_2546);
nand U2727 (N_2727,N_2434,N_2475);
or U2728 (N_2728,N_2405,N_2538);
and U2729 (N_2729,N_2595,N_2538);
xor U2730 (N_2730,N_2548,N_2438);
nor U2731 (N_2731,N_2420,N_2556);
nor U2732 (N_2732,N_2593,N_2497);
and U2733 (N_2733,N_2407,N_2437);
xnor U2734 (N_2734,N_2467,N_2585);
or U2735 (N_2735,N_2520,N_2510);
and U2736 (N_2736,N_2549,N_2456);
and U2737 (N_2737,N_2459,N_2527);
and U2738 (N_2738,N_2469,N_2548);
nand U2739 (N_2739,N_2462,N_2487);
and U2740 (N_2740,N_2472,N_2543);
nor U2741 (N_2741,N_2532,N_2528);
or U2742 (N_2742,N_2549,N_2468);
nand U2743 (N_2743,N_2456,N_2469);
and U2744 (N_2744,N_2547,N_2409);
xor U2745 (N_2745,N_2509,N_2579);
and U2746 (N_2746,N_2403,N_2599);
or U2747 (N_2747,N_2529,N_2423);
xor U2748 (N_2748,N_2511,N_2493);
and U2749 (N_2749,N_2528,N_2407);
nor U2750 (N_2750,N_2454,N_2515);
xnor U2751 (N_2751,N_2509,N_2437);
xor U2752 (N_2752,N_2565,N_2485);
and U2753 (N_2753,N_2591,N_2502);
or U2754 (N_2754,N_2599,N_2425);
xnor U2755 (N_2755,N_2529,N_2482);
nor U2756 (N_2756,N_2475,N_2402);
nor U2757 (N_2757,N_2474,N_2529);
xnor U2758 (N_2758,N_2461,N_2449);
or U2759 (N_2759,N_2433,N_2464);
or U2760 (N_2760,N_2592,N_2578);
nor U2761 (N_2761,N_2429,N_2488);
and U2762 (N_2762,N_2520,N_2413);
xor U2763 (N_2763,N_2557,N_2422);
nand U2764 (N_2764,N_2522,N_2448);
and U2765 (N_2765,N_2504,N_2583);
or U2766 (N_2766,N_2421,N_2446);
nor U2767 (N_2767,N_2532,N_2485);
nand U2768 (N_2768,N_2573,N_2418);
xnor U2769 (N_2769,N_2484,N_2481);
and U2770 (N_2770,N_2413,N_2585);
nor U2771 (N_2771,N_2589,N_2510);
and U2772 (N_2772,N_2578,N_2477);
nand U2773 (N_2773,N_2569,N_2526);
and U2774 (N_2774,N_2408,N_2429);
and U2775 (N_2775,N_2521,N_2411);
nand U2776 (N_2776,N_2415,N_2570);
nand U2777 (N_2777,N_2591,N_2432);
and U2778 (N_2778,N_2502,N_2441);
xnor U2779 (N_2779,N_2404,N_2475);
nor U2780 (N_2780,N_2520,N_2550);
or U2781 (N_2781,N_2473,N_2444);
xnor U2782 (N_2782,N_2502,N_2507);
nor U2783 (N_2783,N_2489,N_2492);
and U2784 (N_2784,N_2476,N_2506);
xor U2785 (N_2785,N_2578,N_2539);
nor U2786 (N_2786,N_2467,N_2412);
nand U2787 (N_2787,N_2551,N_2504);
and U2788 (N_2788,N_2588,N_2596);
or U2789 (N_2789,N_2428,N_2561);
and U2790 (N_2790,N_2554,N_2402);
xor U2791 (N_2791,N_2426,N_2579);
nor U2792 (N_2792,N_2566,N_2455);
or U2793 (N_2793,N_2516,N_2401);
nand U2794 (N_2794,N_2539,N_2494);
nor U2795 (N_2795,N_2413,N_2572);
nor U2796 (N_2796,N_2442,N_2477);
and U2797 (N_2797,N_2437,N_2480);
nor U2798 (N_2798,N_2424,N_2554);
or U2799 (N_2799,N_2438,N_2527);
or U2800 (N_2800,N_2612,N_2750);
nand U2801 (N_2801,N_2754,N_2644);
nor U2802 (N_2802,N_2735,N_2647);
nand U2803 (N_2803,N_2734,N_2655);
xor U2804 (N_2804,N_2753,N_2628);
nor U2805 (N_2805,N_2712,N_2726);
xnor U2806 (N_2806,N_2605,N_2782);
xor U2807 (N_2807,N_2727,N_2739);
or U2808 (N_2808,N_2787,N_2718);
xnor U2809 (N_2809,N_2625,N_2758);
nand U2810 (N_2810,N_2618,N_2622);
xor U2811 (N_2811,N_2669,N_2645);
xnor U2812 (N_2812,N_2616,N_2763);
nor U2813 (N_2813,N_2662,N_2708);
and U2814 (N_2814,N_2690,N_2694);
or U2815 (N_2815,N_2770,N_2659);
nor U2816 (N_2816,N_2615,N_2676);
nor U2817 (N_2817,N_2776,N_2799);
nor U2818 (N_2818,N_2733,N_2725);
and U2819 (N_2819,N_2672,N_2643);
nor U2820 (N_2820,N_2654,N_2697);
nand U2821 (N_2821,N_2617,N_2639);
nand U2822 (N_2822,N_2757,N_2778);
nor U2823 (N_2823,N_2777,N_2620);
nand U2824 (N_2824,N_2685,N_2611);
nand U2825 (N_2825,N_2706,N_2723);
nor U2826 (N_2826,N_2765,N_2746);
xor U2827 (N_2827,N_2724,N_2684);
and U2828 (N_2828,N_2695,N_2696);
nand U2829 (N_2829,N_2744,N_2749);
or U2830 (N_2830,N_2607,N_2720);
xor U2831 (N_2831,N_2716,N_2798);
nand U2832 (N_2832,N_2774,N_2679);
and U2833 (N_2833,N_2624,N_2796);
xnor U2834 (N_2834,N_2630,N_2791);
xnor U2835 (N_2835,N_2674,N_2748);
nand U2836 (N_2836,N_2663,N_2772);
and U2837 (N_2837,N_2713,N_2736);
xor U2838 (N_2838,N_2670,N_2728);
nor U2839 (N_2839,N_2755,N_2722);
nor U2840 (N_2840,N_2707,N_2636);
nor U2841 (N_2841,N_2637,N_2691);
nand U2842 (N_2842,N_2661,N_2732);
and U2843 (N_2843,N_2714,N_2666);
and U2844 (N_2844,N_2703,N_2682);
or U2845 (N_2845,N_2677,N_2740);
nor U2846 (N_2846,N_2760,N_2797);
xnor U2847 (N_2847,N_2788,N_2786);
or U2848 (N_2848,N_2689,N_2642);
nand U2849 (N_2849,N_2784,N_2623);
nand U2850 (N_2850,N_2640,N_2742);
nand U2851 (N_2851,N_2619,N_2656);
or U2852 (N_2852,N_2650,N_2793);
nor U2853 (N_2853,N_2702,N_2638);
xor U2854 (N_2854,N_2609,N_2613);
and U2855 (N_2855,N_2602,N_2651);
nor U2856 (N_2856,N_2604,N_2704);
nand U2857 (N_2857,N_2603,N_2657);
and U2858 (N_2858,N_2715,N_2648);
nor U2859 (N_2859,N_2692,N_2610);
nor U2860 (N_2860,N_2693,N_2719);
nand U2861 (N_2861,N_2667,N_2653);
and U2862 (N_2862,N_2680,N_2792);
nand U2863 (N_2863,N_2683,N_2730);
or U2864 (N_2864,N_2766,N_2606);
xor U2865 (N_2865,N_2687,N_2737);
nand U2866 (N_2866,N_2633,N_2686);
and U2867 (N_2867,N_2794,N_2789);
nor U2868 (N_2868,N_2688,N_2705);
and U2869 (N_2869,N_2701,N_2635);
nor U2870 (N_2870,N_2731,N_2775);
and U2871 (N_2871,N_2721,N_2678);
and U2872 (N_2872,N_2785,N_2698);
nand U2873 (N_2873,N_2780,N_2658);
or U2874 (N_2874,N_2632,N_2756);
and U2875 (N_2875,N_2717,N_2627);
or U2876 (N_2876,N_2795,N_2665);
and U2877 (N_2877,N_2738,N_2768);
nor U2878 (N_2878,N_2629,N_2781);
and U2879 (N_2879,N_2626,N_2790);
nor U2880 (N_2880,N_2783,N_2769);
nand U2881 (N_2881,N_2646,N_2745);
nand U2882 (N_2882,N_2752,N_2711);
nand U2883 (N_2883,N_2700,N_2668);
nand U2884 (N_2884,N_2779,N_2741);
and U2885 (N_2885,N_2631,N_2751);
or U2886 (N_2886,N_2761,N_2641);
nor U2887 (N_2887,N_2671,N_2699);
nor U2888 (N_2888,N_2601,N_2764);
xnor U2889 (N_2889,N_2600,N_2759);
nor U2890 (N_2890,N_2614,N_2649);
or U2891 (N_2891,N_2660,N_2710);
or U2892 (N_2892,N_2762,N_2634);
xor U2893 (N_2893,N_2675,N_2729);
nor U2894 (N_2894,N_2709,N_2773);
and U2895 (N_2895,N_2664,N_2743);
or U2896 (N_2896,N_2608,N_2767);
and U2897 (N_2897,N_2747,N_2652);
and U2898 (N_2898,N_2681,N_2771);
and U2899 (N_2899,N_2621,N_2673);
nor U2900 (N_2900,N_2726,N_2671);
nor U2901 (N_2901,N_2707,N_2648);
xor U2902 (N_2902,N_2749,N_2719);
or U2903 (N_2903,N_2685,N_2763);
and U2904 (N_2904,N_2770,N_2752);
or U2905 (N_2905,N_2603,N_2608);
and U2906 (N_2906,N_2688,N_2714);
nor U2907 (N_2907,N_2635,N_2744);
and U2908 (N_2908,N_2744,N_2666);
xnor U2909 (N_2909,N_2797,N_2733);
xor U2910 (N_2910,N_2783,N_2670);
nand U2911 (N_2911,N_2704,N_2700);
xnor U2912 (N_2912,N_2740,N_2799);
nand U2913 (N_2913,N_2657,N_2706);
xnor U2914 (N_2914,N_2717,N_2784);
nand U2915 (N_2915,N_2709,N_2765);
or U2916 (N_2916,N_2661,N_2781);
nor U2917 (N_2917,N_2639,N_2783);
and U2918 (N_2918,N_2608,N_2712);
nor U2919 (N_2919,N_2785,N_2756);
or U2920 (N_2920,N_2759,N_2690);
or U2921 (N_2921,N_2614,N_2663);
xor U2922 (N_2922,N_2743,N_2634);
or U2923 (N_2923,N_2668,N_2760);
or U2924 (N_2924,N_2623,N_2715);
nor U2925 (N_2925,N_2711,N_2786);
and U2926 (N_2926,N_2608,N_2701);
nand U2927 (N_2927,N_2776,N_2729);
xnor U2928 (N_2928,N_2747,N_2738);
xor U2929 (N_2929,N_2615,N_2700);
and U2930 (N_2930,N_2709,N_2680);
or U2931 (N_2931,N_2612,N_2700);
xnor U2932 (N_2932,N_2621,N_2658);
and U2933 (N_2933,N_2694,N_2648);
xnor U2934 (N_2934,N_2797,N_2759);
nor U2935 (N_2935,N_2624,N_2674);
and U2936 (N_2936,N_2741,N_2660);
or U2937 (N_2937,N_2630,N_2674);
and U2938 (N_2938,N_2744,N_2710);
and U2939 (N_2939,N_2744,N_2687);
and U2940 (N_2940,N_2775,N_2664);
nand U2941 (N_2941,N_2700,N_2795);
xor U2942 (N_2942,N_2644,N_2628);
or U2943 (N_2943,N_2602,N_2726);
and U2944 (N_2944,N_2698,N_2606);
xor U2945 (N_2945,N_2697,N_2653);
nor U2946 (N_2946,N_2789,N_2630);
xnor U2947 (N_2947,N_2674,N_2784);
or U2948 (N_2948,N_2732,N_2635);
nor U2949 (N_2949,N_2713,N_2700);
nor U2950 (N_2950,N_2608,N_2659);
nor U2951 (N_2951,N_2738,N_2632);
xor U2952 (N_2952,N_2627,N_2647);
xnor U2953 (N_2953,N_2725,N_2710);
nor U2954 (N_2954,N_2665,N_2729);
or U2955 (N_2955,N_2668,N_2643);
nor U2956 (N_2956,N_2656,N_2796);
xor U2957 (N_2957,N_2689,N_2767);
xnor U2958 (N_2958,N_2624,N_2697);
nor U2959 (N_2959,N_2769,N_2633);
or U2960 (N_2960,N_2603,N_2719);
nor U2961 (N_2961,N_2681,N_2770);
nand U2962 (N_2962,N_2780,N_2714);
and U2963 (N_2963,N_2715,N_2790);
and U2964 (N_2964,N_2789,N_2626);
xor U2965 (N_2965,N_2704,N_2750);
and U2966 (N_2966,N_2731,N_2630);
xor U2967 (N_2967,N_2783,N_2778);
and U2968 (N_2968,N_2600,N_2659);
nand U2969 (N_2969,N_2753,N_2693);
nand U2970 (N_2970,N_2781,N_2695);
nor U2971 (N_2971,N_2708,N_2628);
or U2972 (N_2972,N_2669,N_2702);
and U2973 (N_2973,N_2713,N_2731);
and U2974 (N_2974,N_2779,N_2659);
and U2975 (N_2975,N_2609,N_2636);
xnor U2976 (N_2976,N_2793,N_2722);
nand U2977 (N_2977,N_2648,N_2794);
or U2978 (N_2978,N_2707,N_2627);
nand U2979 (N_2979,N_2684,N_2790);
and U2980 (N_2980,N_2635,N_2680);
nand U2981 (N_2981,N_2638,N_2671);
or U2982 (N_2982,N_2716,N_2654);
nand U2983 (N_2983,N_2691,N_2603);
nor U2984 (N_2984,N_2696,N_2777);
nand U2985 (N_2985,N_2645,N_2662);
xnor U2986 (N_2986,N_2788,N_2708);
xnor U2987 (N_2987,N_2612,N_2611);
or U2988 (N_2988,N_2711,N_2731);
or U2989 (N_2989,N_2677,N_2728);
nand U2990 (N_2990,N_2617,N_2613);
xor U2991 (N_2991,N_2753,N_2714);
and U2992 (N_2992,N_2601,N_2794);
nor U2993 (N_2993,N_2768,N_2765);
xnor U2994 (N_2994,N_2789,N_2763);
or U2995 (N_2995,N_2798,N_2632);
nand U2996 (N_2996,N_2748,N_2688);
nand U2997 (N_2997,N_2613,N_2623);
nand U2998 (N_2998,N_2661,N_2682);
xor U2999 (N_2999,N_2719,N_2717);
nor U3000 (N_3000,N_2896,N_2921);
xnor U3001 (N_3001,N_2866,N_2969);
and U3002 (N_3002,N_2957,N_2887);
nand U3003 (N_3003,N_2811,N_2905);
nand U3004 (N_3004,N_2936,N_2915);
nand U3005 (N_3005,N_2844,N_2837);
or U3006 (N_3006,N_2922,N_2865);
nand U3007 (N_3007,N_2986,N_2924);
nand U3008 (N_3008,N_2966,N_2952);
and U3009 (N_3009,N_2870,N_2963);
nor U3010 (N_3010,N_2933,N_2939);
nor U3011 (N_3011,N_2850,N_2805);
or U3012 (N_3012,N_2882,N_2889);
nor U3013 (N_3013,N_2959,N_2836);
xor U3014 (N_3014,N_2843,N_2877);
nor U3015 (N_3015,N_2995,N_2958);
and U3016 (N_3016,N_2853,N_2816);
and U3017 (N_3017,N_2947,N_2984);
xnor U3018 (N_3018,N_2810,N_2983);
or U3019 (N_3019,N_2817,N_2938);
nor U3020 (N_3020,N_2895,N_2916);
xor U3021 (N_3021,N_2824,N_2885);
or U3022 (N_3022,N_2934,N_2860);
nor U3023 (N_3023,N_2935,N_2872);
and U3024 (N_3024,N_2980,N_2847);
nor U3025 (N_3025,N_2826,N_2903);
and U3026 (N_3026,N_2912,N_2869);
or U3027 (N_3027,N_2875,N_2845);
or U3028 (N_3028,N_2953,N_2914);
or U3029 (N_3029,N_2876,N_2891);
nor U3030 (N_3030,N_2863,N_2800);
xnor U3031 (N_3031,N_2890,N_2991);
or U3032 (N_3032,N_2929,N_2808);
xor U3033 (N_3033,N_2910,N_2954);
xor U3034 (N_3034,N_2878,N_2928);
nand U3035 (N_3035,N_2967,N_2972);
xor U3036 (N_3036,N_2806,N_2812);
xnor U3037 (N_3037,N_2804,N_2940);
nor U3038 (N_3038,N_2907,N_2849);
and U3039 (N_3039,N_2923,N_2948);
xor U3040 (N_3040,N_2814,N_2900);
and U3041 (N_3041,N_2888,N_2978);
xnor U3042 (N_3042,N_2973,N_2994);
and U3043 (N_3043,N_2856,N_2813);
nand U3044 (N_3044,N_2820,N_2868);
and U3045 (N_3045,N_2827,N_2977);
nor U3046 (N_3046,N_2988,N_2899);
or U3047 (N_3047,N_2927,N_2828);
and U3048 (N_3048,N_2913,N_2852);
nand U3049 (N_3049,N_2803,N_2884);
and U3050 (N_3050,N_2943,N_2864);
xor U3051 (N_3051,N_2955,N_2989);
and U3052 (N_3052,N_2840,N_2846);
xnor U3053 (N_3053,N_2861,N_2975);
nand U3054 (N_3054,N_2883,N_2944);
or U3055 (N_3055,N_2981,N_2998);
xnor U3056 (N_3056,N_2990,N_2946);
nand U3057 (N_3057,N_2964,N_2961);
or U3058 (N_3058,N_2829,N_2880);
xnor U3059 (N_3059,N_2979,N_2819);
or U3060 (N_3060,N_2881,N_2902);
xor U3061 (N_3061,N_2841,N_2976);
or U3062 (N_3062,N_2833,N_2830);
nand U3063 (N_3063,N_2823,N_2997);
xnor U3064 (N_3064,N_2931,N_2821);
nand U3065 (N_3065,N_2909,N_2809);
nand U3066 (N_3066,N_2892,N_2897);
nor U3067 (N_3067,N_2965,N_2960);
nand U3068 (N_3068,N_2925,N_2838);
or U3069 (N_3069,N_2857,N_2992);
xnor U3070 (N_3070,N_2950,N_2908);
nand U3071 (N_3071,N_2996,N_2839);
or U3072 (N_3072,N_2918,N_2949);
xnor U3073 (N_3073,N_2858,N_2971);
xnor U3074 (N_3074,N_2815,N_2894);
nor U3075 (N_3075,N_2901,N_2801);
or U3076 (N_3076,N_2974,N_2835);
nor U3077 (N_3077,N_2985,N_2911);
or U3078 (N_3078,N_2930,N_2987);
nor U3079 (N_3079,N_2945,N_2906);
nand U3080 (N_3080,N_2873,N_2825);
and U3081 (N_3081,N_2926,N_2970);
xor U3082 (N_3082,N_2807,N_2879);
xnor U3083 (N_3083,N_2920,N_2951);
and U3084 (N_3084,N_2867,N_2993);
xor U3085 (N_3085,N_2898,N_2862);
and U3086 (N_3086,N_2848,N_2982);
nand U3087 (N_3087,N_2937,N_2941);
nand U3088 (N_3088,N_2842,N_2832);
or U3089 (N_3089,N_2831,N_2818);
nor U3090 (N_3090,N_2851,N_2942);
or U3091 (N_3091,N_2956,N_2874);
xnor U3092 (N_3092,N_2999,N_2962);
xnor U3093 (N_3093,N_2855,N_2904);
nand U3094 (N_3094,N_2893,N_2822);
nand U3095 (N_3095,N_2854,N_2834);
nor U3096 (N_3096,N_2917,N_2932);
nor U3097 (N_3097,N_2919,N_2871);
or U3098 (N_3098,N_2802,N_2859);
nor U3099 (N_3099,N_2886,N_2968);
nand U3100 (N_3100,N_2899,N_2934);
nor U3101 (N_3101,N_2824,N_2980);
nand U3102 (N_3102,N_2973,N_2854);
xor U3103 (N_3103,N_2959,N_2992);
or U3104 (N_3104,N_2873,N_2979);
nor U3105 (N_3105,N_2965,N_2808);
or U3106 (N_3106,N_2851,N_2825);
xnor U3107 (N_3107,N_2929,N_2893);
nor U3108 (N_3108,N_2905,N_2869);
xnor U3109 (N_3109,N_2926,N_2976);
nand U3110 (N_3110,N_2990,N_2960);
xor U3111 (N_3111,N_2841,N_2801);
and U3112 (N_3112,N_2813,N_2853);
nand U3113 (N_3113,N_2990,N_2805);
nand U3114 (N_3114,N_2945,N_2996);
and U3115 (N_3115,N_2862,N_2846);
and U3116 (N_3116,N_2804,N_2981);
and U3117 (N_3117,N_2938,N_2877);
nor U3118 (N_3118,N_2998,N_2961);
nor U3119 (N_3119,N_2807,N_2959);
or U3120 (N_3120,N_2825,N_2859);
nand U3121 (N_3121,N_2825,N_2812);
and U3122 (N_3122,N_2923,N_2970);
nor U3123 (N_3123,N_2850,N_2873);
nand U3124 (N_3124,N_2907,N_2829);
nand U3125 (N_3125,N_2929,N_2823);
xor U3126 (N_3126,N_2824,N_2848);
nand U3127 (N_3127,N_2972,N_2989);
nor U3128 (N_3128,N_2938,N_2906);
nand U3129 (N_3129,N_2855,N_2949);
nor U3130 (N_3130,N_2923,N_2914);
and U3131 (N_3131,N_2987,N_2836);
nor U3132 (N_3132,N_2903,N_2884);
xnor U3133 (N_3133,N_2944,N_2889);
nor U3134 (N_3134,N_2903,N_2898);
xor U3135 (N_3135,N_2993,N_2899);
nand U3136 (N_3136,N_2811,N_2822);
nand U3137 (N_3137,N_2879,N_2918);
or U3138 (N_3138,N_2833,N_2995);
nor U3139 (N_3139,N_2961,N_2955);
or U3140 (N_3140,N_2842,N_2910);
nor U3141 (N_3141,N_2855,N_2915);
nor U3142 (N_3142,N_2879,N_2883);
nor U3143 (N_3143,N_2945,N_2862);
nand U3144 (N_3144,N_2955,N_2994);
nor U3145 (N_3145,N_2909,N_2924);
nand U3146 (N_3146,N_2950,N_2958);
and U3147 (N_3147,N_2824,N_2915);
and U3148 (N_3148,N_2975,N_2816);
nand U3149 (N_3149,N_2975,N_2860);
and U3150 (N_3150,N_2914,N_2988);
and U3151 (N_3151,N_2928,N_2964);
nand U3152 (N_3152,N_2822,N_2972);
or U3153 (N_3153,N_2806,N_2819);
and U3154 (N_3154,N_2875,N_2963);
nor U3155 (N_3155,N_2823,N_2949);
nand U3156 (N_3156,N_2815,N_2832);
and U3157 (N_3157,N_2848,N_2888);
or U3158 (N_3158,N_2920,N_2937);
nand U3159 (N_3159,N_2857,N_2809);
nor U3160 (N_3160,N_2943,N_2985);
nand U3161 (N_3161,N_2832,N_2830);
xor U3162 (N_3162,N_2842,N_2837);
and U3163 (N_3163,N_2888,N_2906);
or U3164 (N_3164,N_2978,N_2933);
nand U3165 (N_3165,N_2992,N_2875);
or U3166 (N_3166,N_2978,N_2809);
or U3167 (N_3167,N_2837,N_2993);
nand U3168 (N_3168,N_2878,N_2977);
or U3169 (N_3169,N_2813,N_2942);
nor U3170 (N_3170,N_2953,N_2956);
or U3171 (N_3171,N_2905,N_2943);
or U3172 (N_3172,N_2981,N_2808);
and U3173 (N_3173,N_2985,N_2880);
nand U3174 (N_3174,N_2930,N_2849);
nand U3175 (N_3175,N_2847,N_2925);
and U3176 (N_3176,N_2864,N_2816);
xor U3177 (N_3177,N_2962,N_2928);
xnor U3178 (N_3178,N_2960,N_2981);
xnor U3179 (N_3179,N_2860,N_2971);
or U3180 (N_3180,N_2881,N_2921);
and U3181 (N_3181,N_2952,N_2994);
xnor U3182 (N_3182,N_2803,N_2962);
xnor U3183 (N_3183,N_2910,N_2820);
or U3184 (N_3184,N_2987,N_2928);
or U3185 (N_3185,N_2899,N_2802);
xnor U3186 (N_3186,N_2985,N_2865);
or U3187 (N_3187,N_2959,N_2921);
xor U3188 (N_3188,N_2814,N_2831);
xnor U3189 (N_3189,N_2865,N_2921);
nor U3190 (N_3190,N_2806,N_2845);
nor U3191 (N_3191,N_2966,N_2921);
or U3192 (N_3192,N_2951,N_2851);
nor U3193 (N_3193,N_2960,N_2956);
nand U3194 (N_3194,N_2940,N_2842);
xnor U3195 (N_3195,N_2989,N_2889);
nor U3196 (N_3196,N_2865,N_2926);
and U3197 (N_3197,N_2840,N_2833);
nand U3198 (N_3198,N_2964,N_2917);
nand U3199 (N_3199,N_2841,N_2862);
or U3200 (N_3200,N_3144,N_3147);
and U3201 (N_3201,N_3104,N_3077);
xnor U3202 (N_3202,N_3198,N_3155);
nand U3203 (N_3203,N_3195,N_3022);
nand U3204 (N_3204,N_3135,N_3036);
nand U3205 (N_3205,N_3093,N_3148);
and U3206 (N_3206,N_3040,N_3037);
or U3207 (N_3207,N_3019,N_3152);
or U3208 (N_3208,N_3119,N_3051);
xor U3209 (N_3209,N_3114,N_3165);
and U3210 (N_3210,N_3164,N_3023);
nor U3211 (N_3211,N_3065,N_3010);
xor U3212 (N_3212,N_3140,N_3158);
nand U3213 (N_3213,N_3009,N_3141);
nor U3214 (N_3214,N_3126,N_3060);
and U3215 (N_3215,N_3125,N_3074);
nor U3216 (N_3216,N_3149,N_3151);
nand U3217 (N_3217,N_3012,N_3015);
and U3218 (N_3218,N_3177,N_3002);
and U3219 (N_3219,N_3150,N_3039);
and U3220 (N_3220,N_3187,N_3079);
or U3221 (N_3221,N_3008,N_3053);
nor U3222 (N_3222,N_3184,N_3007);
and U3223 (N_3223,N_3196,N_3067);
xnor U3224 (N_3224,N_3115,N_3075);
xor U3225 (N_3225,N_3143,N_3068);
xnor U3226 (N_3226,N_3156,N_3084);
or U3227 (N_3227,N_3044,N_3167);
xor U3228 (N_3228,N_3056,N_3088);
and U3229 (N_3229,N_3081,N_3050);
nor U3230 (N_3230,N_3041,N_3063);
nor U3231 (N_3231,N_3070,N_3153);
or U3232 (N_3232,N_3188,N_3017);
and U3233 (N_3233,N_3059,N_3159);
nand U3234 (N_3234,N_3082,N_3111);
xor U3235 (N_3235,N_3013,N_3197);
and U3236 (N_3236,N_3049,N_3011);
or U3237 (N_3237,N_3107,N_3090);
xor U3238 (N_3238,N_3194,N_3179);
xnor U3239 (N_3239,N_3096,N_3110);
or U3240 (N_3240,N_3109,N_3100);
or U3241 (N_3241,N_3116,N_3089);
nor U3242 (N_3242,N_3024,N_3138);
or U3243 (N_3243,N_3083,N_3055);
xnor U3244 (N_3244,N_3026,N_3062);
xnor U3245 (N_3245,N_3146,N_3168);
and U3246 (N_3246,N_3029,N_3098);
nor U3247 (N_3247,N_3154,N_3004);
nor U3248 (N_3248,N_3170,N_3066);
and U3249 (N_3249,N_3129,N_3130);
nand U3250 (N_3250,N_3185,N_3020);
and U3251 (N_3251,N_3157,N_3192);
nor U3252 (N_3252,N_3193,N_3064);
nor U3253 (N_3253,N_3128,N_3103);
xnor U3254 (N_3254,N_3131,N_3134);
xnor U3255 (N_3255,N_3127,N_3080);
xor U3256 (N_3256,N_3145,N_3174);
and U3257 (N_3257,N_3061,N_3035);
and U3258 (N_3258,N_3120,N_3097);
nor U3259 (N_3259,N_3005,N_3101);
nand U3260 (N_3260,N_3175,N_3122);
xor U3261 (N_3261,N_3031,N_3118);
nor U3262 (N_3262,N_3112,N_3182);
xor U3263 (N_3263,N_3001,N_3014);
nand U3264 (N_3264,N_3087,N_3071);
or U3265 (N_3265,N_3190,N_3160);
and U3266 (N_3266,N_3176,N_3132);
and U3267 (N_3267,N_3072,N_3106);
and U3268 (N_3268,N_3048,N_3043);
and U3269 (N_3269,N_3034,N_3133);
or U3270 (N_3270,N_3028,N_3163);
nand U3271 (N_3271,N_3058,N_3136);
nor U3272 (N_3272,N_3046,N_3052);
and U3273 (N_3273,N_3045,N_3178);
and U3274 (N_3274,N_3092,N_3105);
and U3275 (N_3275,N_3000,N_3042);
xnor U3276 (N_3276,N_3123,N_3073);
and U3277 (N_3277,N_3057,N_3139);
nor U3278 (N_3278,N_3016,N_3095);
nor U3279 (N_3279,N_3085,N_3171);
xor U3280 (N_3280,N_3189,N_3181);
nor U3281 (N_3281,N_3142,N_3006);
nor U3282 (N_3282,N_3069,N_3047);
or U3283 (N_3283,N_3027,N_3099);
nand U3284 (N_3284,N_3003,N_3191);
xor U3285 (N_3285,N_3117,N_3054);
xor U3286 (N_3286,N_3032,N_3033);
nand U3287 (N_3287,N_3086,N_3172);
or U3288 (N_3288,N_3078,N_3180);
or U3289 (N_3289,N_3021,N_3199);
xor U3290 (N_3290,N_3102,N_3173);
nor U3291 (N_3291,N_3166,N_3025);
nor U3292 (N_3292,N_3108,N_3169);
xor U3293 (N_3293,N_3161,N_3186);
and U3294 (N_3294,N_3030,N_3124);
nor U3295 (N_3295,N_3121,N_3038);
or U3296 (N_3296,N_3091,N_3076);
and U3297 (N_3297,N_3018,N_3113);
or U3298 (N_3298,N_3183,N_3162);
or U3299 (N_3299,N_3137,N_3094);
xor U3300 (N_3300,N_3152,N_3023);
nor U3301 (N_3301,N_3001,N_3192);
or U3302 (N_3302,N_3194,N_3006);
xor U3303 (N_3303,N_3183,N_3015);
or U3304 (N_3304,N_3091,N_3159);
and U3305 (N_3305,N_3001,N_3050);
nor U3306 (N_3306,N_3013,N_3034);
and U3307 (N_3307,N_3029,N_3099);
xnor U3308 (N_3308,N_3100,N_3080);
nor U3309 (N_3309,N_3036,N_3094);
xnor U3310 (N_3310,N_3111,N_3105);
or U3311 (N_3311,N_3081,N_3147);
and U3312 (N_3312,N_3154,N_3084);
xor U3313 (N_3313,N_3194,N_3083);
or U3314 (N_3314,N_3165,N_3106);
or U3315 (N_3315,N_3019,N_3055);
nor U3316 (N_3316,N_3115,N_3147);
xor U3317 (N_3317,N_3047,N_3131);
nand U3318 (N_3318,N_3196,N_3009);
nand U3319 (N_3319,N_3009,N_3171);
or U3320 (N_3320,N_3110,N_3165);
and U3321 (N_3321,N_3105,N_3086);
or U3322 (N_3322,N_3028,N_3024);
xor U3323 (N_3323,N_3142,N_3029);
or U3324 (N_3324,N_3100,N_3182);
xor U3325 (N_3325,N_3076,N_3143);
nor U3326 (N_3326,N_3183,N_3009);
and U3327 (N_3327,N_3123,N_3083);
xor U3328 (N_3328,N_3147,N_3009);
nor U3329 (N_3329,N_3191,N_3127);
and U3330 (N_3330,N_3055,N_3081);
or U3331 (N_3331,N_3164,N_3038);
or U3332 (N_3332,N_3012,N_3070);
nand U3333 (N_3333,N_3007,N_3148);
and U3334 (N_3334,N_3085,N_3110);
xnor U3335 (N_3335,N_3084,N_3002);
nand U3336 (N_3336,N_3195,N_3043);
or U3337 (N_3337,N_3040,N_3160);
nor U3338 (N_3338,N_3018,N_3080);
xnor U3339 (N_3339,N_3166,N_3056);
or U3340 (N_3340,N_3074,N_3135);
or U3341 (N_3341,N_3151,N_3011);
and U3342 (N_3342,N_3113,N_3121);
nand U3343 (N_3343,N_3086,N_3024);
xor U3344 (N_3344,N_3025,N_3138);
nand U3345 (N_3345,N_3081,N_3193);
nand U3346 (N_3346,N_3194,N_3144);
or U3347 (N_3347,N_3153,N_3130);
xor U3348 (N_3348,N_3107,N_3106);
nor U3349 (N_3349,N_3033,N_3175);
or U3350 (N_3350,N_3167,N_3149);
or U3351 (N_3351,N_3139,N_3168);
xor U3352 (N_3352,N_3154,N_3043);
or U3353 (N_3353,N_3051,N_3086);
and U3354 (N_3354,N_3140,N_3075);
xor U3355 (N_3355,N_3065,N_3012);
or U3356 (N_3356,N_3003,N_3102);
and U3357 (N_3357,N_3181,N_3077);
nor U3358 (N_3358,N_3181,N_3074);
nor U3359 (N_3359,N_3105,N_3186);
and U3360 (N_3360,N_3156,N_3179);
nor U3361 (N_3361,N_3028,N_3081);
or U3362 (N_3362,N_3025,N_3180);
nor U3363 (N_3363,N_3152,N_3004);
nor U3364 (N_3364,N_3182,N_3029);
or U3365 (N_3365,N_3090,N_3050);
or U3366 (N_3366,N_3118,N_3161);
nor U3367 (N_3367,N_3025,N_3092);
nor U3368 (N_3368,N_3071,N_3154);
or U3369 (N_3369,N_3027,N_3086);
nand U3370 (N_3370,N_3106,N_3168);
or U3371 (N_3371,N_3182,N_3019);
nor U3372 (N_3372,N_3144,N_3091);
nand U3373 (N_3373,N_3045,N_3111);
and U3374 (N_3374,N_3024,N_3152);
and U3375 (N_3375,N_3131,N_3187);
or U3376 (N_3376,N_3143,N_3004);
nor U3377 (N_3377,N_3052,N_3141);
xor U3378 (N_3378,N_3030,N_3185);
nor U3379 (N_3379,N_3050,N_3148);
or U3380 (N_3380,N_3148,N_3026);
and U3381 (N_3381,N_3117,N_3043);
xnor U3382 (N_3382,N_3042,N_3065);
nand U3383 (N_3383,N_3054,N_3111);
xor U3384 (N_3384,N_3053,N_3016);
and U3385 (N_3385,N_3158,N_3024);
nand U3386 (N_3386,N_3170,N_3189);
or U3387 (N_3387,N_3195,N_3081);
and U3388 (N_3388,N_3181,N_3089);
nand U3389 (N_3389,N_3059,N_3189);
or U3390 (N_3390,N_3188,N_3040);
nor U3391 (N_3391,N_3061,N_3168);
nor U3392 (N_3392,N_3060,N_3143);
nand U3393 (N_3393,N_3096,N_3002);
nand U3394 (N_3394,N_3007,N_3062);
nand U3395 (N_3395,N_3199,N_3165);
or U3396 (N_3396,N_3090,N_3095);
and U3397 (N_3397,N_3172,N_3016);
or U3398 (N_3398,N_3036,N_3186);
nand U3399 (N_3399,N_3199,N_3028);
and U3400 (N_3400,N_3298,N_3350);
or U3401 (N_3401,N_3202,N_3391);
nor U3402 (N_3402,N_3356,N_3274);
nor U3403 (N_3403,N_3390,N_3313);
nand U3404 (N_3404,N_3263,N_3302);
xnor U3405 (N_3405,N_3281,N_3395);
nor U3406 (N_3406,N_3246,N_3222);
xnor U3407 (N_3407,N_3327,N_3223);
nand U3408 (N_3408,N_3292,N_3229);
xor U3409 (N_3409,N_3207,N_3251);
and U3410 (N_3410,N_3219,N_3373);
nand U3411 (N_3411,N_3394,N_3340);
or U3412 (N_3412,N_3325,N_3264);
nor U3413 (N_3413,N_3288,N_3291);
and U3414 (N_3414,N_3224,N_3268);
nand U3415 (N_3415,N_3284,N_3342);
nor U3416 (N_3416,N_3205,N_3399);
xor U3417 (N_3417,N_3280,N_3217);
nand U3418 (N_3418,N_3321,N_3343);
or U3419 (N_3419,N_3286,N_3267);
nand U3420 (N_3420,N_3308,N_3386);
or U3421 (N_3421,N_3220,N_3297);
nor U3422 (N_3422,N_3260,N_3293);
and U3423 (N_3423,N_3314,N_3369);
and U3424 (N_3424,N_3273,N_3261);
xnor U3425 (N_3425,N_3335,N_3221);
nand U3426 (N_3426,N_3269,N_3357);
or U3427 (N_3427,N_3243,N_3257);
nand U3428 (N_3428,N_3360,N_3320);
or U3429 (N_3429,N_3277,N_3240);
xnor U3430 (N_3430,N_3236,N_3275);
nor U3431 (N_3431,N_3228,N_3363);
or U3432 (N_3432,N_3227,N_3290);
and U3433 (N_3433,N_3309,N_3361);
or U3434 (N_3434,N_3215,N_3254);
and U3435 (N_3435,N_3244,N_3330);
and U3436 (N_3436,N_3364,N_3262);
nand U3437 (N_3437,N_3326,N_3295);
nand U3438 (N_3438,N_3365,N_3331);
xnor U3439 (N_3439,N_3241,N_3358);
or U3440 (N_3440,N_3255,N_3301);
nand U3441 (N_3441,N_3375,N_3209);
nand U3442 (N_3442,N_3249,N_3256);
or U3443 (N_3443,N_3247,N_3259);
xnor U3444 (N_3444,N_3283,N_3278);
or U3445 (N_3445,N_3370,N_3347);
nand U3446 (N_3446,N_3334,N_3387);
nand U3447 (N_3447,N_3248,N_3332);
or U3448 (N_3448,N_3374,N_3235);
nor U3449 (N_3449,N_3388,N_3352);
nor U3450 (N_3450,N_3378,N_3234);
xnor U3451 (N_3451,N_3204,N_3294);
nand U3452 (N_3452,N_3226,N_3316);
nand U3453 (N_3453,N_3203,N_3230);
nor U3454 (N_3454,N_3368,N_3385);
and U3455 (N_3455,N_3276,N_3303);
and U3456 (N_3456,N_3201,N_3318);
or U3457 (N_3457,N_3237,N_3362);
or U3458 (N_3458,N_3367,N_3306);
or U3459 (N_3459,N_3351,N_3384);
and U3460 (N_3460,N_3376,N_3353);
or U3461 (N_3461,N_3305,N_3285);
nor U3462 (N_3462,N_3250,N_3382);
and U3463 (N_3463,N_3231,N_3393);
nand U3464 (N_3464,N_3265,N_3397);
nand U3465 (N_3465,N_3296,N_3272);
nor U3466 (N_3466,N_3289,N_3300);
xor U3467 (N_3467,N_3315,N_3212);
nand U3468 (N_3468,N_3266,N_3396);
nor U3469 (N_3469,N_3398,N_3366);
or U3470 (N_3470,N_3339,N_3206);
xnor U3471 (N_3471,N_3372,N_3242);
xor U3472 (N_3472,N_3379,N_3349);
nand U3473 (N_3473,N_3355,N_3328);
nand U3474 (N_3474,N_3218,N_3329);
nand U3475 (N_3475,N_3322,N_3389);
nand U3476 (N_3476,N_3381,N_3311);
and U3477 (N_3477,N_3345,N_3344);
nand U3478 (N_3478,N_3348,N_3341);
nand U3479 (N_3479,N_3279,N_3211);
xor U3480 (N_3480,N_3323,N_3239);
xor U3481 (N_3481,N_3299,N_3216);
or U3482 (N_3482,N_3346,N_3312);
nor U3483 (N_3483,N_3253,N_3213);
nand U3484 (N_3484,N_3337,N_3333);
nor U3485 (N_3485,N_3336,N_3214);
nand U3486 (N_3486,N_3210,N_3270);
or U3487 (N_3487,N_3377,N_3383);
or U3488 (N_3488,N_3307,N_3287);
xor U3489 (N_3489,N_3310,N_3304);
xnor U3490 (N_3490,N_3319,N_3324);
and U3491 (N_3491,N_3354,N_3252);
nor U3492 (N_3492,N_3317,N_3359);
xnor U3493 (N_3493,N_3338,N_3258);
and U3494 (N_3494,N_3392,N_3371);
nand U3495 (N_3495,N_3271,N_3200);
and U3496 (N_3496,N_3232,N_3238);
xor U3497 (N_3497,N_3282,N_3233);
nand U3498 (N_3498,N_3225,N_3380);
nand U3499 (N_3499,N_3245,N_3208);
nor U3500 (N_3500,N_3216,N_3368);
nand U3501 (N_3501,N_3231,N_3336);
and U3502 (N_3502,N_3264,N_3330);
and U3503 (N_3503,N_3284,N_3259);
nand U3504 (N_3504,N_3371,N_3209);
and U3505 (N_3505,N_3339,N_3239);
nand U3506 (N_3506,N_3335,N_3367);
nor U3507 (N_3507,N_3318,N_3398);
nor U3508 (N_3508,N_3234,N_3272);
nand U3509 (N_3509,N_3267,N_3278);
nor U3510 (N_3510,N_3270,N_3388);
nor U3511 (N_3511,N_3264,N_3244);
nand U3512 (N_3512,N_3332,N_3329);
or U3513 (N_3513,N_3262,N_3206);
and U3514 (N_3514,N_3393,N_3332);
nor U3515 (N_3515,N_3278,N_3394);
nand U3516 (N_3516,N_3247,N_3392);
nor U3517 (N_3517,N_3231,N_3294);
xnor U3518 (N_3518,N_3220,N_3298);
nor U3519 (N_3519,N_3348,N_3364);
or U3520 (N_3520,N_3389,N_3293);
nor U3521 (N_3521,N_3337,N_3211);
nand U3522 (N_3522,N_3233,N_3224);
xnor U3523 (N_3523,N_3330,N_3363);
or U3524 (N_3524,N_3382,N_3221);
or U3525 (N_3525,N_3200,N_3348);
and U3526 (N_3526,N_3272,N_3389);
and U3527 (N_3527,N_3204,N_3326);
and U3528 (N_3528,N_3319,N_3335);
nand U3529 (N_3529,N_3384,N_3367);
or U3530 (N_3530,N_3372,N_3373);
nor U3531 (N_3531,N_3284,N_3367);
nor U3532 (N_3532,N_3263,N_3226);
and U3533 (N_3533,N_3232,N_3303);
nor U3534 (N_3534,N_3348,N_3310);
nor U3535 (N_3535,N_3242,N_3353);
xor U3536 (N_3536,N_3378,N_3380);
and U3537 (N_3537,N_3250,N_3335);
nor U3538 (N_3538,N_3211,N_3285);
and U3539 (N_3539,N_3380,N_3390);
or U3540 (N_3540,N_3325,N_3337);
xnor U3541 (N_3541,N_3262,N_3297);
or U3542 (N_3542,N_3251,N_3204);
or U3543 (N_3543,N_3213,N_3271);
nor U3544 (N_3544,N_3227,N_3353);
and U3545 (N_3545,N_3296,N_3343);
nor U3546 (N_3546,N_3257,N_3393);
or U3547 (N_3547,N_3233,N_3229);
nand U3548 (N_3548,N_3366,N_3225);
and U3549 (N_3549,N_3311,N_3280);
xor U3550 (N_3550,N_3359,N_3278);
nor U3551 (N_3551,N_3379,N_3326);
or U3552 (N_3552,N_3226,N_3215);
xnor U3553 (N_3553,N_3226,N_3309);
nand U3554 (N_3554,N_3263,N_3340);
or U3555 (N_3555,N_3233,N_3244);
or U3556 (N_3556,N_3232,N_3375);
and U3557 (N_3557,N_3284,N_3206);
nand U3558 (N_3558,N_3355,N_3291);
or U3559 (N_3559,N_3218,N_3343);
or U3560 (N_3560,N_3238,N_3306);
and U3561 (N_3561,N_3356,N_3265);
xnor U3562 (N_3562,N_3392,N_3275);
or U3563 (N_3563,N_3332,N_3264);
and U3564 (N_3564,N_3211,N_3388);
nand U3565 (N_3565,N_3284,N_3317);
or U3566 (N_3566,N_3205,N_3335);
or U3567 (N_3567,N_3211,N_3297);
nor U3568 (N_3568,N_3221,N_3255);
nor U3569 (N_3569,N_3282,N_3290);
and U3570 (N_3570,N_3254,N_3262);
nand U3571 (N_3571,N_3276,N_3367);
or U3572 (N_3572,N_3217,N_3376);
and U3573 (N_3573,N_3256,N_3215);
nand U3574 (N_3574,N_3361,N_3333);
nand U3575 (N_3575,N_3290,N_3277);
nor U3576 (N_3576,N_3256,N_3390);
and U3577 (N_3577,N_3369,N_3327);
nand U3578 (N_3578,N_3349,N_3346);
xnor U3579 (N_3579,N_3243,N_3209);
nand U3580 (N_3580,N_3364,N_3362);
or U3581 (N_3581,N_3216,N_3301);
or U3582 (N_3582,N_3330,N_3378);
nor U3583 (N_3583,N_3225,N_3262);
xor U3584 (N_3584,N_3224,N_3326);
xnor U3585 (N_3585,N_3211,N_3347);
and U3586 (N_3586,N_3263,N_3323);
nand U3587 (N_3587,N_3340,N_3309);
nor U3588 (N_3588,N_3296,N_3256);
xor U3589 (N_3589,N_3286,N_3204);
or U3590 (N_3590,N_3364,N_3267);
xnor U3591 (N_3591,N_3346,N_3332);
nand U3592 (N_3592,N_3248,N_3244);
nor U3593 (N_3593,N_3318,N_3388);
xor U3594 (N_3594,N_3299,N_3265);
and U3595 (N_3595,N_3395,N_3324);
nor U3596 (N_3596,N_3351,N_3385);
nand U3597 (N_3597,N_3375,N_3287);
and U3598 (N_3598,N_3313,N_3276);
xor U3599 (N_3599,N_3237,N_3224);
and U3600 (N_3600,N_3458,N_3480);
xnor U3601 (N_3601,N_3592,N_3438);
nor U3602 (N_3602,N_3474,N_3552);
nand U3603 (N_3603,N_3518,N_3578);
nand U3604 (N_3604,N_3506,N_3455);
nand U3605 (N_3605,N_3441,N_3416);
nor U3606 (N_3606,N_3580,N_3529);
or U3607 (N_3607,N_3428,N_3510);
and U3608 (N_3608,N_3443,N_3499);
nor U3609 (N_3609,N_3485,N_3589);
xor U3610 (N_3610,N_3465,N_3525);
nand U3611 (N_3611,N_3425,N_3456);
xnor U3612 (N_3612,N_3496,N_3426);
or U3613 (N_3613,N_3431,N_3437);
nand U3614 (N_3614,N_3545,N_3445);
or U3615 (N_3615,N_3538,N_3422);
nor U3616 (N_3616,N_3436,N_3514);
and U3617 (N_3617,N_3566,N_3432);
nand U3618 (N_3618,N_3528,N_3421);
nand U3619 (N_3619,N_3473,N_3537);
and U3620 (N_3620,N_3430,N_3556);
nand U3621 (N_3621,N_3502,N_3493);
or U3622 (N_3622,N_3540,N_3504);
xnor U3623 (N_3623,N_3517,N_3560);
and U3624 (N_3624,N_3530,N_3500);
or U3625 (N_3625,N_3501,N_3484);
nand U3626 (N_3626,N_3562,N_3417);
nor U3627 (N_3627,N_3531,N_3450);
nand U3628 (N_3628,N_3483,N_3435);
or U3629 (N_3629,N_3524,N_3404);
xnor U3630 (N_3630,N_3551,N_3403);
or U3631 (N_3631,N_3587,N_3564);
xor U3632 (N_3632,N_3419,N_3581);
xnor U3633 (N_3633,N_3521,N_3548);
nand U3634 (N_3634,N_3519,N_3522);
or U3635 (N_3635,N_3497,N_3513);
and U3636 (N_3636,N_3492,N_3516);
and U3637 (N_3637,N_3415,N_3457);
xnor U3638 (N_3638,N_3579,N_3414);
and U3639 (N_3639,N_3568,N_3448);
or U3640 (N_3640,N_3572,N_3424);
and U3641 (N_3641,N_3406,N_3459);
nor U3642 (N_3642,N_3418,N_3462);
xor U3643 (N_3643,N_3554,N_3544);
and U3644 (N_3644,N_3463,N_3582);
and U3645 (N_3645,N_3583,N_3569);
and U3646 (N_3646,N_3471,N_3488);
nand U3647 (N_3647,N_3405,N_3434);
nor U3648 (N_3648,N_3588,N_3547);
nor U3649 (N_3649,N_3489,N_3447);
nand U3650 (N_3650,N_3527,N_3549);
nor U3651 (N_3651,N_3487,N_3557);
or U3652 (N_3652,N_3539,N_3520);
nand U3653 (N_3653,N_3571,N_3585);
xor U3654 (N_3654,N_3509,N_3594);
nand U3655 (N_3655,N_3512,N_3439);
xor U3656 (N_3656,N_3523,N_3472);
or U3657 (N_3657,N_3532,N_3402);
xnor U3658 (N_3658,N_3526,N_3481);
or U3659 (N_3659,N_3593,N_3536);
or U3660 (N_3660,N_3543,N_3558);
xnor U3661 (N_3661,N_3442,N_3508);
nor U3662 (N_3662,N_3440,N_3598);
xor U3663 (N_3663,N_3559,N_3565);
and U3664 (N_3664,N_3475,N_3570);
or U3665 (N_3665,N_3444,N_3413);
xor U3666 (N_3666,N_3479,N_3561);
or U3667 (N_3667,N_3446,N_3533);
or U3668 (N_3668,N_3453,N_3574);
and U3669 (N_3669,N_3468,N_3553);
xnor U3670 (N_3670,N_3505,N_3460);
xnor U3671 (N_3671,N_3467,N_3476);
nor U3672 (N_3672,N_3427,N_3411);
nand U3673 (N_3673,N_3482,N_3408);
xor U3674 (N_3674,N_3550,N_3573);
nor U3675 (N_3675,N_3423,N_3555);
nor U3676 (N_3676,N_3542,N_3400);
or U3677 (N_3677,N_3466,N_3534);
and U3678 (N_3678,N_3491,N_3469);
nand U3679 (N_3679,N_3584,N_3596);
nor U3680 (N_3680,N_3576,N_3590);
nand U3681 (N_3681,N_3449,N_3515);
xnor U3682 (N_3682,N_3498,N_3490);
xor U3683 (N_3683,N_3546,N_3586);
nor U3684 (N_3684,N_3486,N_3599);
or U3685 (N_3685,N_3429,N_3507);
and U3686 (N_3686,N_3407,N_3563);
xnor U3687 (N_3687,N_3410,N_3597);
nand U3688 (N_3688,N_3541,N_3494);
and U3689 (N_3689,N_3575,N_3477);
nor U3690 (N_3690,N_3452,N_3503);
xor U3691 (N_3691,N_3511,N_3464);
nor U3692 (N_3692,N_3567,N_3595);
nor U3693 (N_3693,N_3433,N_3461);
xor U3694 (N_3694,N_3401,N_3470);
nor U3695 (N_3695,N_3409,N_3591);
or U3696 (N_3696,N_3412,N_3535);
and U3697 (N_3697,N_3478,N_3495);
or U3698 (N_3698,N_3420,N_3451);
xnor U3699 (N_3699,N_3577,N_3454);
nand U3700 (N_3700,N_3517,N_3510);
xor U3701 (N_3701,N_3523,N_3586);
nand U3702 (N_3702,N_3424,N_3483);
and U3703 (N_3703,N_3408,N_3598);
and U3704 (N_3704,N_3502,N_3407);
and U3705 (N_3705,N_3583,N_3568);
or U3706 (N_3706,N_3534,N_3432);
or U3707 (N_3707,N_3432,N_3441);
xor U3708 (N_3708,N_3557,N_3408);
nor U3709 (N_3709,N_3415,N_3534);
or U3710 (N_3710,N_3581,N_3517);
and U3711 (N_3711,N_3428,N_3575);
nor U3712 (N_3712,N_3441,N_3578);
nand U3713 (N_3713,N_3574,N_3588);
nand U3714 (N_3714,N_3539,N_3410);
or U3715 (N_3715,N_3460,N_3414);
nor U3716 (N_3716,N_3598,N_3540);
nor U3717 (N_3717,N_3589,N_3481);
or U3718 (N_3718,N_3423,N_3489);
xor U3719 (N_3719,N_3435,N_3469);
nor U3720 (N_3720,N_3534,N_3481);
xor U3721 (N_3721,N_3545,N_3490);
nor U3722 (N_3722,N_3528,N_3550);
nand U3723 (N_3723,N_3593,N_3522);
and U3724 (N_3724,N_3540,N_3593);
nand U3725 (N_3725,N_3487,N_3458);
nor U3726 (N_3726,N_3468,N_3434);
and U3727 (N_3727,N_3539,N_3529);
nor U3728 (N_3728,N_3562,N_3524);
nor U3729 (N_3729,N_3524,N_3451);
xnor U3730 (N_3730,N_3470,N_3473);
or U3731 (N_3731,N_3480,N_3403);
xor U3732 (N_3732,N_3578,N_3500);
nand U3733 (N_3733,N_3563,N_3529);
nand U3734 (N_3734,N_3503,N_3583);
xnor U3735 (N_3735,N_3576,N_3454);
xor U3736 (N_3736,N_3466,N_3524);
nand U3737 (N_3737,N_3463,N_3543);
nand U3738 (N_3738,N_3402,N_3501);
nand U3739 (N_3739,N_3451,N_3407);
nor U3740 (N_3740,N_3554,N_3510);
nor U3741 (N_3741,N_3531,N_3495);
xnor U3742 (N_3742,N_3515,N_3456);
and U3743 (N_3743,N_3520,N_3579);
nor U3744 (N_3744,N_3430,N_3442);
nand U3745 (N_3745,N_3500,N_3407);
nand U3746 (N_3746,N_3434,N_3447);
xnor U3747 (N_3747,N_3589,N_3415);
and U3748 (N_3748,N_3461,N_3430);
or U3749 (N_3749,N_3445,N_3514);
xor U3750 (N_3750,N_3473,N_3434);
nand U3751 (N_3751,N_3525,N_3511);
nor U3752 (N_3752,N_3582,N_3592);
or U3753 (N_3753,N_3430,N_3432);
or U3754 (N_3754,N_3489,N_3504);
and U3755 (N_3755,N_3423,N_3403);
or U3756 (N_3756,N_3550,N_3447);
nor U3757 (N_3757,N_3511,N_3519);
nor U3758 (N_3758,N_3437,N_3464);
or U3759 (N_3759,N_3407,N_3546);
nand U3760 (N_3760,N_3598,N_3426);
or U3761 (N_3761,N_3549,N_3441);
xnor U3762 (N_3762,N_3438,N_3521);
and U3763 (N_3763,N_3438,N_3559);
or U3764 (N_3764,N_3505,N_3444);
and U3765 (N_3765,N_3400,N_3592);
nand U3766 (N_3766,N_3501,N_3593);
or U3767 (N_3767,N_3433,N_3568);
or U3768 (N_3768,N_3539,N_3493);
nand U3769 (N_3769,N_3485,N_3409);
xor U3770 (N_3770,N_3427,N_3513);
nand U3771 (N_3771,N_3426,N_3423);
and U3772 (N_3772,N_3420,N_3452);
and U3773 (N_3773,N_3454,N_3549);
xnor U3774 (N_3774,N_3481,N_3551);
or U3775 (N_3775,N_3530,N_3557);
xnor U3776 (N_3776,N_3480,N_3457);
xor U3777 (N_3777,N_3567,N_3513);
nand U3778 (N_3778,N_3574,N_3425);
or U3779 (N_3779,N_3467,N_3452);
and U3780 (N_3780,N_3436,N_3469);
nor U3781 (N_3781,N_3455,N_3447);
nand U3782 (N_3782,N_3557,N_3413);
nor U3783 (N_3783,N_3502,N_3590);
nand U3784 (N_3784,N_3499,N_3418);
and U3785 (N_3785,N_3433,N_3486);
nor U3786 (N_3786,N_3499,N_3502);
nor U3787 (N_3787,N_3526,N_3513);
xor U3788 (N_3788,N_3470,N_3462);
nor U3789 (N_3789,N_3415,N_3506);
or U3790 (N_3790,N_3456,N_3529);
nor U3791 (N_3791,N_3467,N_3522);
nand U3792 (N_3792,N_3568,N_3554);
or U3793 (N_3793,N_3421,N_3536);
nor U3794 (N_3794,N_3438,N_3491);
nand U3795 (N_3795,N_3513,N_3535);
xor U3796 (N_3796,N_3414,N_3542);
nand U3797 (N_3797,N_3503,N_3498);
nor U3798 (N_3798,N_3562,N_3564);
xnor U3799 (N_3799,N_3486,N_3444);
nand U3800 (N_3800,N_3730,N_3660);
xnor U3801 (N_3801,N_3619,N_3671);
and U3802 (N_3802,N_3767,N_3645);
nand U3803 (N_3803,N_3750,N_3777);
nand U3804 (N_3804,N_3673,N_3625);
nor U3805 (N_3805,N_3784,N_3614);
and U3806 (N_3806,N_3733,N_3612);
nand U3807 (N_3807,N_3719,N_3718);
nand U3808 (N_3808,N_3787,N_3623);
or U3809 (N_3809,N_3616,N_3712);
and U3810 (N_3810,N_3654,N_3615);
nand U3811 (N_3811,N_3791,N_3697);
and U3812 (N_3812,N_3650,N_3748);
nor U3813 (N_3813,N_3702,N_3735);
and U3814 (N_3814,N_3769,N_3698);
nor U3815 (N_3815,N_3694,N_3655);
and U3816 (N_3816,N_3795,N_3648);
nor U3817 (N_3817,N_3796,N_3674);
xor U3818 (N_3818,N_3688,N_3610);
nand U3819 (N_3819,N_3708,N_3653);
or U3820 (N_3820,N_3740,N_3644);
or U3821 (N_3821,N_3741,N_3755);
nor U3822 (N_3822,N_3634,N_3753);
nor U3823 (N_3823,N_3700,N_3731);
and U3824 (N_3824,N_3754,N_3649);
xor U3825 (N_3825,N_3627,N_3626);
or U3826 (N_3826,N_3770,N_3679);
nand U3827 (N_3827,N_3659,N_3678);
xnor U3828 (N_3828,N_3724,N_3797);
and U3829 (N_3829,N_3773,N_3662);
and U3830 (N_3830,N_3651,N_3752);
xor U3831 (N_3831,N_3604,N_3603);
and U3832 (N_3832,N_3643,N_3788);
or U3833 (N_3833,N_3756,N_3707);
xor U3834 (N_3834,N_3620,N_3768);
or U3835 (N_3835,N_3696,N_3792);
xor U3836 (N_3836,N_3647,N_3605);
and U3837 (N_3837,N_3613,N_3779);
and U3838 (N_3838,N_3761,N_3669);
and U3839 (N_3839,N_3666,N_3636);
or U3840 (N_3840,N_3732,N_3691);
and U3841 (N_3841,N_3789,N_3680);
and U3842 (N_3842,N_3664,N_3723);
xor U3843 (N_3843,N_3606,N_3781);
and U3844 (N_3844,N_3630,N_3764);
nor U3845 (N_3845,N_3635,N_3621);
nor U3846 (N_3846,N_3640,N_3722);
or U3847 (N_3847,N_3624,N_3729);
nand U3848 (N_3848,N_3747,N_3658);
xnor U3849 (N_3849,N_3628,N_3738);
nor U3850 (N_3850,N_3629,N_3672);
xnor U3851 (N_3851,N_3631,N_3745);
or U3852 (N_3852,N_3701,N_3646);
or U3853 (N_3853,N_3641,N_3771);
or U3854 (N_3854,N_3783,N_3780);
nand U3855 (N_3855,N_3736,N_3675);
nand U3856 (N_3856,N_3763,N_3676);
nor U3857 (N_3857,N_3601,N_3652);
xnor U3858 (N_3858,N_3607,N_3693);
or U3859 (N_3859,N_3692,N_3706);
nor U3860 (N_3860,N_3746,N_3775);
or U3861 (N_3861,N_3728,N_3744);
xnor U3862 (N_3862,N_3786,N_3642);
or U3863 (N_3863,N_3682,N_3661);
nor U3864 (N_3864,N_3685,N_3600);
nor U3865 (N_3865,N_3766,N_3798);
and U3866 (N_3866,N_3668,N_3703);
nor U3867 (N_3867,N_3737,N_3602);
nor U3868 (N_3868,N_3751,N_3665);
nand U3869 (N_3869,N_3695,N_3622);
xnor U3870 (N_3870,N_3794,N_3759);
or U3871 (N_3871,N_3705,N_3726);
nor U3872 (N_3872,N_3717,N_3657);
xor U3873 (N_3873,N_3739,N_3758);
and U3874 (N_3874,N_3721,N_3713);
and U3875 (N_3875,N_3699,N_3677);
xnor U3876 (N_3876,N_3734,N_3742);
nor U3877 (N_3877,N_3632,N_3785);
and U3878 (N_3878,N_3663,N_3715);
xnor U3879 (N_3879,N_3633,N_3684);
nor U3880 (N_3880,N_3689,N_3725);
nand U3881 (N_3881,N_3778,N_3714);
and U3882 (N_3882,N_3790,N_3757);
nor U3883 (N_3883,N_3667,N_3716);
nor U3884 (N_3884,N_3608,N_3772);
nand U3885 (N_3885,N_3711,N_3656);
xnor U3886 (N_3886,N_3720,N_3687);
or U3887 (N_3887,N_3782,N_3681);
and U3888 (N_3888,N_3611,N_3793);
nor U3889 (N_3889,N_3709,N_3617);
nand U3890 (N_3890,N_3760,N_3776);
and U3891 (N_3891,N_3762,N_3704);
and U3892 (N_3892,N_3609,N_3686);
nand U3893 (N_3893,N_3710,N_3799);
xnor U3894 (N_3894,N_3690,N_3765);
nand U3895 (N_3895,N_3618,N_3749);
and U3896 (N_3896,N_3639,N_3670);
xnor U3897 (N_3897,N_3743,N_3638);
xnor U3898 (N_3898,N_3683,N_3774);
xnor U3899 (N_3899,N_3637,N_3727);
and U3900 (N_3900,N_3656,N_3610);
and U3901 (N_3901,N_3649,N_3650);
or U3902 (N_3902,N_3709,N_3729);
nand U3903 (N_3903,N_3667,N_3776);
or U3904 (N_3904,N_3679,N_3686);
or U3905 (N_3905,N_3713,N_3708);
xnor U3906 (N_3906,N_3717,N_3778);
nand U3907 (N_3907,N_3616,N_3798);
nor U3908 (N_3908,N_3688,N_3692);
nor U3909 (N_3909,N_3754,N_3774);
and U3910 (N_3910,N_3611,N_3617);
xor U3911 (N_3911,N_3661,N_3645);
nor U3912 (N_3912,N_3703,N_3765);
and U3913 (N_3913,N_3776,N_3698);
and U3914 (N_3914,N_3664,N_3702);
xor U3915 (N_3915,N_3685,N_3721);
or U3916 (N_3916,N_3788,N_3667);
nor U3917 (N_3917,N_3782,N_3715);
nor U3918 (N_3918,N_3645,N_3668);
and U3919 (N_3919,N_3787,N_3633);
xnor U3920 (N_3920,N_3785,N_3684);
xor U3921 (N_3921,N_3797,N_3684);
and U3922 (N_3922,N_3607,N_3601);
and U3923 (N_3923,N_3638,N_3623);
or U3924 (N_3924,N_3710,N_3706);
nand U3925 (N_3925,N_3777,N_3687);
xnor U3926 (N_3926,N_3639,N_3669);
nand U3927 (N_3927,N_3794,N_3715);
or U3928 (N_3928,N_3650,N_3793);
nor U3929 (N_3929,N_3738,N_3630);
or U3930 (N_3930,N_3682,N_3691);
nor U3931 (N_3931,N_3705,N_3738);
or U3932 (N_3932,N_3740,N_3767);
and U3933 (N_3933,N_3721,N_3611);
xnor U3934 (N_3934,N_3636,N_3764);
nand U3935 (N_3935,N_3660,N_3610);
or U3936 (N_3936,N_3757,N_3692);
nor U3937 (N_3937,N_3723,N_3778);
or U3938 (N_3938,N_3612,N_3661);
or U3939 (N_3939,N_3787,N_3605);
xnor U3940 (N_3940,N_3728,N_3643);
nor U3941 (N_3941,N_3757,N_3716);
nor U3942 (N_3942,N_3629,N_3695);
nand U3943 (N_3943,N_3721,N_3772);
or U3944 (N_3944,N_3670,N_3741);
xnor U3945 (N_3945,N_3758,N_3694);
or U3946 (N_3946,N_3776,N_3770);
nor U3947 (N_3947,N_3613,N_3763);
xor U3948 (N_3948,N_3616,N_3618);
and U3949 (N_3949,N_3668,N_3670);
nor U3950 (N_3950,N_3714,N_3624);
nand U3951 (N_3951,N_3769,N_3744);
nand U3952 (N_3952,N_3743,N_3752);
nand U3953 (N_3953,N_3735,N_3697);
and U3954 (N_3954,N_3644,N_3653);
xor U3955 (N_3955,N_3784,N_3743);
and U3956 (N_3956,N_3782,N_3640);
nand U3957 (N_3957,N_3753,N_3722);
nor U3958 (N_3958,N_3755,N_3769);
nor U3959 (N_3959,N_3706,N_3640);
and U3960 (N_3960,N_3736,N_3614);
nand U3961 (N_3961,N_3657,N_3667);
or U3962 (N_3962,N_3757,N_3719);
nor U3963 (N_3963,N_3663,N_3625);
nand U3964 (N_3964,N_3724,N_3600);
nand U3965 (N_3965,N_3677,N_3792);
nor U3966 (N_3966,N_3638,N_3759);
and U3967 (N_3967,N_3794,N_3791);
nand U3968 (N_3968,N_3672,N_3698);
or U3969 (N_3969,N_3730,N_3714);
nor U3970 (N_3970,N_3612,N_3793);
xor U3971 (N_3971,N_3719,N_3722);
xor U3972 (N_3972,N_3778,N_3765);
or U3973 (N_3973,N_3719,N_3651);
or U3974 (N_3974,N_3738,N_3788);
xnor U3975 (N_3975,N_3737,N_3616);
or U3976 (N_3976,N_3781,N_3779);
or U3977 (N_3977,N_3661,N_3738);
and U3978 (N_3978,N_3678,N_3773);
or U3979 (N_3979,N_3665,N_3650);
and U3980 (N_3980,N_3792,N_3706);
or U3981 (N_3981,N_3771,N_3731);
or U3982 (N_3982,N_3754,N_3783);
and U3983 (N_3983,N_3713,N_3632);
or U3984 (N_3984,N_3765,N_3628);
or U3985 (N_3985,N_3793,N_3604);
nand U3986 (N_3986,N_3729,N_3779);
nor U3987 (N_3987,N_3799,N_3666);
or U3988 (N_3988,N_3632,N_3767);
xor U3989 (N_3989,N_3788,N_3603);
and U3990 (N_3990,N_3600,N_3652);
xor U3991 (N_3991,N_3688,N_3638);
nand U3992 (N_3992,N_3672,N_3773);
or U3993 (N_3993,N_3680,N_3783);
xnor U3994 (N_3994,N_3614,N_3602);
nor U3995 (N_3995,N_3611,N_3675);
xor U3996 (N_3996,N_3772,N_3691);
nor U3997 (N_3997,N_3620,N_3764);
or U3998 (N_3998,N_3702,N_3665);
nor U3999 (N_3999,N_3709,N_3799);
xnor U4000 (N_4000,N_3860,N_3961);
nor U4001 (N_4001,N_3894,N_3879);
nor U4002 (N_4002,N_3976,N_3964);
or U4003 (N_4003,N_3923,N_3973);
and U4004 (N_4004,N_3890,N_3908);
nand U4005 (N_4005,N_3844,N_3820);
nor U4006 (N_4006,N_3987,N_3944);
and U4007 (N_4007,N_3869,N_3899);
and U4008 (N_4008,N_3870,N_3943);
or U4009 (N_4009,N_3849,N_3813);
or U4010 (N_4010,N_3905,N_3913);
or U4011 (N_4011,N_3836,N_3975);
or U4012 (N_4012,N_3941,N_3934);
and U4013 (N_4013,N_3839,N_3978);
nand U4014 (N_4014,N_3972,N_3911);
nand U4015 (N_4015,N_3887,N_3931);
nor U4016 (N_4016,N_3924,N_3974);
nor U4017 (N_4017,N_3886,N_3998);
nand U4018 (N_4018,N_3970,N_3932);
or U4019 (N_4019,N_3925,N_3891);
or U4020 (N_4020,N_3919,N_3935);
and U4021 (N_4021,N_3865,N_3895);
and U4022 (N_4022,N_3817,N_3822);
nand U4023 (N_4023,N_3901,N_3880);
nand U4024 (N_4024,N_3854,N_3996);
nor U4025 (N_4025,N_3846,N_3856);
or U4026 (N_4026,N_3804,N_3858);
or U4027 (N_4027,N_3889,N_3936);
or U4028 (N_4028,N_3861,N_3878);
nor U4029 (N_4029,N_3990,N_3949);
and U4030 (N_4030,N_3893,N_3853);
nand U4031 (N_4031,N_3828,N_3994);
nand U4032 (N_4032,N_3912,N_3948);
xor U4033 (N_4033,N_3995,N_3906);
and U4034 (N_4034,N_3967,N_3966);
or U4035 (N_4035,N_3831,N_3914);
xnor U4036 (N_4036,N_3953,N_3947);
nand U4037 (N_4037,N_3985,N_3819);
nor U4038 (N_4038,N_3897,N_3875);
or U4039 (N_4039,N_3945,N_3814);
and U4040 (N_4040,N_3900,N_3868);
nand U4041 (N_4041,N_3827,N_3808);
nand U4042 (N_4042,N_3882,N_3837);
nand U4043 (N_4043,N_3946,N_3968);
or U4044 (N_4044,N_3991,N_3825);
nand U4045 (N_4045,N_3933,N_3818);
nor U4046 (N_4046,N_3927,N_3993);
nand U4047 (N_4047,N_3942,N_3824);
and U4048 (N_4048,N_3848,N_3957);
xnor U4049 (N_4049,N_3977,N_3845);
nor U4050 (N_4050,N_3959,N_3835);
and U4051 (N_4051,N_3840,N_3963);
nand U4052 (N_4052,N_3940,N_3956);
xor U4053 (N_4053,N_3806,N_3898);
and U4054 (N_4054,N_3971,N_3852);
nor U4055 (N_4055,N_3833,N_3962);
or U4056 (N_4056,N_3917,N_3850);
or U4057 (N_4057,N_3955,N_3902);
nor U4058 (N_4058,N_3881,N_3910);
nand U4059 (N_4059,N_3939,N_3988);
xor U4060 (N_4060,N_3812,N_3952);
or U4061 (N_4061,N_3809,N_3892);
xnor U4062 (N_4062,N_3929,N_3984);
or U4063 (N_4063,N_3829,N_3802);
xnor U4064 (N_4064,N_3872,N_3979);
xor U4065 (N_4065,N_3969,N_3830);
nor U4066 (N_4066,N_3816,N_3847);
nor U4067 (N_4067,N_3915,N_3862);
and U4068 (N_4068,N_3938,N_3871);
nor U4069 (N_4069,N_3866,N_3834);
or U4070 (N_4070,N_3986,N_3876);
or U4071 (N_4071,N_3982,N_3877);
nand U4072 (N_4072,N_3983,N_3928);
or U4073 (N_4073,N_3867,N_3821);
or U4074 (N_4074,N_3904,N_3930);
or U4075 (N_4075,N_3920,N_3926);
and U4076 (N_4076,N_3992,N_3859);
nand U4077 (N_4077,N_3803,N_3838);
and U4078 (N_4078,N_3857,N_3918);
xnor U4079 (N_4079,N_3801,N_3884);
nand U4080 (N_4080,N_3874,N_3907);
and U4081 (N_4081,N_3826,N_3863);
nand U4082 (N_4082,N_3811,N_3981);
nor U4083 (N_4083,N_3805,N_3800);
or U4084 (N_4084,N_3951,N_3989);
or U4085 (N_4085,N_3807,N_3873);
and U4086 (N_4086,N_3888,N_3885);
xnor U4087 (N_4087,N_3965,N_3823);
and U4088 (N_4088,N_3832,N_3842);
xnor U4089 (N_4089,N_3997,N_3950);
xor U4090 (N_4090,N_3903,N_3841);
and U4091 (N_4091,N_3815,N_3980);
or U4092 (N_4092,N_3922,N_3883);
xnor U4093 (N_4093,N_3843,N_3999);
or U4094 (N_4094,N_3954,N_3896);
xor U4095 (N_4095,N_3958,N_3851);
xor U4096 (N_4096,N_3921,N_3916);
nor U4097 (N_4097,N_3864,N_3937);
and U4098 (N_4098,N_3855,N_3909);
nand U4099 (N_4099,N_3810,N_3960);
nand U4100 (N_4100,N_3891,N_3872);
nand U4101 (N_4101,N_3806,N_3901);
and U4102 (N_4102,N_3861,N_3945);
and U4103 (N_4103,N_3877,N_3932);
nand U4104 (N_4104,N_3942,N_3935);
nand U4105 (N_4105,N_3811,N_3883);
xnor U4106 (N_4106,N_3858,N_3869);
and U4107 (N_4107,N_3912,N_3878);
nand U4108 (N_4108,N_3842,N_3833);
xnor U4109 (N_4109,N_3974,N_3865);
nand U4110 (N_4110,N_3991,N_3958);
and U4111 (N_4111,N_3852,N_3830);
and U4112 (N_4112,N_3834,N_3959);
or U4113 (N_4113,N_3923,N_3805);
and U4114 (N_4114,N_3976,N_3812);
xor U4115 (N_4115,N_3877,N_3800);
and U4116 (N_4116,N_3817,N_3849);
and U4117 (N_4117,N_3952,N_3906);
nor U4118 (N_4118,N_3931,N_3948);
or U4119 (N_4119,N_3935,N_3948);
nor U4120 (N_4120,N_3958,N_3862);
xnor U4121 (N_4121,N_3908,N_3958);
and U4122 (N_4122,N_3833,N_3861);
or U4123 (N_4123,N_3885,N_3830);
xor U4124 (N_4124,N_3920,N_3856);
xnor U4125 (N_4125,N_3997,N_3881);
and U4126 (N_4126,N_3967,N_3949);
nand U4127 (N_4127,N_3887,N_3981);
and U4128 (N_4128,N_3828,N_3879);
nand U4129 (N_4129,N_3829,N_3869);
or U4130 (N_4130,N_3973,N_3867);
nor U4131 (N_4131,N_3851,N_3984);
xor U4132 (N_4132,N_3964,N_3816);
nor U4133 (N_4133,N_3918,N_3996);
nand U4134 (N_4134,N_3829,N_3932);
or U4135 (N_4135,N_3966,N_3944);
xor U4136 (N_4136,N_3942,N_3920);
and U4137 (N_4137,N_3882,N_3848);
nor U4138 (N_4138,N_3860,N_3939);
or U4139 (N_4139,N_3813,N_3987);
or U4140 (N_4140,N_3987,N_3977);
nand U4141 (N_4141,N_3828,N_3802);
xnor U4142 (N_4142,N_3947,N_3850);
and U4143 (N_4143,N_3926,N_3924);
nor U4144 (N_4144,N_3877,N_3907);
or U4145 (N_4145,N_3938,N_3864);
or U4146 (N_4146,N_3894,N_3935);
and U4147 (N_4147,N_3825,N_3819);
xor U4148 (N_4148,N_3964,N_3905);
and U4149 (N_4149,N_3991,N_3812);
or U4150 (N_4150,N_3946,N_3868);
nor U4151 (N_4151,N_3929,N_3977);
xor U4152 (N_4152,N_3812,N_3974);
and U4153 (N_4153,N_3938,N_3900);
or U4154 (N_4154,N_3864,N_3839);
nor U4155 (N_4155,N_3834,N_3914);
nor U4156 (N_4156,N_3887,N_3800);
nor U4157 (N_4157,N_3824,N_3945);
or U4158 (N_4158,N_3960,N_3973);
nor U4159 (N_4159,N_3927,N_3930);
nand U4160 (N_4160,N_3994,N_3833);
and U4161 (N_4161,N_3809,N_3885);
and U4162 (N_4162,N_3920,N_3902);
nor U4163 (N_4163,N_3961,N_3820);
xor U4164 (N_4164,N_3829,N_3879);
or U4165 (N_4165,N_3875,N_3950);
xor U4166 (N_4166,N_3993,N_3944);
or U4167 (N_4167,N_3991,N_3919);
or U4168 (N_4168,N_3815,N_3945);
or U4169 (N_4169,N_3897,N_3994);
or U4170 (N_4170,N_3967,N_3939);
and U4171 (N_4171,N_3824,N_3965);
xnor U4172 (N_4172,N_3897,N_3925);
and U4173 (N_4173,N_3937,N_3819);
nor U4174 (N_4174,N_3842,N_3988);
or U4175 (N_4175,N_3891,N_3924);
xor U4176 (N_4176,N_3966,N_3901);
or U4177 (N_4177,N_3961,N_3927);
and U4178 (N_4178,N_3986,N_3994);
or U4179 (N_4179,N_3812,N_3928);
nand U4180 (N_4180,N_3904,N_3863);
nor U4181 (N_4181,N_3917,N_3872);
or U4182 (N_4182,N_3905,N_3867);
or U4183 (N_4183,N_3833,N_3960);
or U4184 (N_4184,N_3837,N_3947);
nand U4185 (N_4185,N_3866,N_3998);
nand U4186 (N_4186,N_3908,N_3854);
and U4187 (N_4187,N_3941,N_3959);
nor U4188 (N_4188,N_3881,N_3927);
or U4189 (N_4189,N_3841,N_3891);
nor U4190 (N_4190,N_3918,N_3961);
nor U4191 (N_4191,N_3905,N_3945);
xnor U4192 (N_4192,N_3909,N_3956);
nand U4193 (N_4193,N_3810,N_3903);
and U4194 (N_4194,N_3960,N_3885);
or U4195 (N_4195,N_3920,N_3987);
xor U4196 (N_4196,N_3846,N_3876);
nand U4197 (N_4197,N_3829,N_3906);
or U4198 (N_4198,N_3893,N_3863);
nor U4199 (N_4199,N_3873,N_3884);
or U4200 (N_4200,N_4035,N_4127);
or U4201 (N_4201,N_4033,N_4052);
xnor U4202 (N_4202,N_4132,N_4122);
nor U4203 (N_4203,N_4078,N_4092);
nand U4204 (N_4204,N_4162,N_4096);
nand U4205 (N_4205,N_4170,N_4040);
and U4206 (N_4206,N_4126,N_4068);
nand U4207 (N_4207,N_4198,N_4071);
or U4208 (N_4208,N_4007,N_4155);
nor U4209 (N_4209,N_4090,N_4081);
nor U4210 (N_4210,N_4185,N_4114);
or U4211 (N_4211,N_4177,N_4029);
nor U4212 (N_4212,N_4001,N_4050);
xnor U4213 (N_4213,N_4134,N_4065);
nand U4214 (N_4214,N_4077,N_4191);
or U4215 (N_4215,N_4037,N_4086);
xnor U4216 (N_4216,N_4051,N_4196);
or U4217 (N_4217,N_4169,N_4095);
nand U4218 (N_4218,N_4004,N_4197);
nor U4219 (N_4219,N_4110,N_4027);
or U4220 (N_4220,N_4047,N_4128);
xor U4221 (N_4221,N_4178,N_4183);
and U4222 (N_4222,N_4010,N_4016);
nor U4223 (N_4223,N_4061,N_4076);
nand U4224 (N_4224,N_4053,N_4159);
xor U4225 (N_4225,N_4190,N_4116);
and U4226 (N_4226,N_4121,N_4113);
and U4227 (N_4227,N_4049,N_4069);
nand U4228 (N_4228,N_4066,N_4039);
nand U4229 (N_4229,N_4102,N_4142);
or U4230 (N_4230,N_4104,N_4024);
and U4231 (N_4231,N_4008,N_4146);
and U4232 (N_4232,N_4042,N_4139);
nand U4233 (N_4233,N_4151,N_4109);
and U4234 (N_4234,N_4025,N_4176);
nor U4235 (N_4235,N_4156,N_4002);
xnor U4236 (N_4236,N_4072,N_4144);
or U4237 (N_4237,N_4145,N_4009);
nand U4238 (N_4238,N_4075,N_4173);
nand U4239 (N_4239,N_4080,N_4137);
or U4240 (N_4240,N_4148,N_4175);
nand U4241 (N_4241,N_4036,N_4083);
nor U4242 (N_4242,N_4011,N_4045);
and U4243 (N_4243,N_4044,N_4098);
and U4244 (N_4244,N_4120,N_4174);
xor U4245 (N_4245,N_4154,N_4131);
or U4246 (N_4246,N_4180,N_4101);
and U4247 (N_4247,N_4149,N_4038);
or U4248 (N_4248,N_4164,N_4118);
nand U4249 (N_4249,N_4105,N_4167);
and U4250 (N_4250,N_4140,N_4070);
and U4251 (N_4251,N_4133,N_4054);
nor U4252 (N_4252,N_4097,N_4056);
nor U4253 (N_4253,N_4182,N_4073);
nand U4254 (N_4254,N_4048,N_4015);
and U4255 (N_4255,N_4089,N_4179);
nand U4256 (N_4256,N_4012,N_4111);
xnor U4257 (N_4257,N_4093,N_4067);
nor U4258 (N_4258,N_4062,N_4184);
nand U4259 (N_4259,N_4041,N_4000);
and U4260 (N_4260,N_4195,N_4057);
xor U4261 (N_4261,N_4030,N_4166);
nand U4262 (N_4262,N_4129,N_4100);
nand U4263 (N_4263,N_4064,N_4088);
and U4264 (N_4264,N_4031,N_4085);
xor U4265 (N_4265,N_4005,N_4194);
nand U4266 (N_4266,N_4094,N_4091);
nand U4267 (N_4267,N_4153,N_4063);
or U4268 (N_4268,N_4171,N_4188);
and U4269 (N_4269,N_4124,N_4108);
nor U4270 (N_4270,N_4163,N_4034);
nor U4271 (N_4271,N_4150,N_4013);
or U4272 (N_4272,N_4152,N_4106);
or U4273 (N_4273,N_4157,N_4193);
nor U4274 (N_4274,N_4115,N_4074);
nand U4275 (N_4275,N_4158,N_4084);
nor U4276 (N_4276,N_4123,N_4082);
xnor U4277 (N_4277,N_4143,N_4168);
xnor U4278 (N_4278,N_4058,N_4055);
nor U4279 (N_4279,N_4019,N_4125);
nor U4280 (N_4280,N_4046,N_4014);
xor U4281 (N_4281,N_4160,N_4020);
nor U4282 (N_4282,N_4192,N_4199);
and U4283 (N_4283,N_4018,N_4172);
nor U4284 (N_4284,N_4130,N_4017);
xor U4285 (N_4285,N_4103,N_4107);
and U4286 (N_4286,N_4136,N_4023);
nor U4287 (N_4287,N_4189,N_4187);
nand U4288 (N_4288,N_4021,N_4147);
nand U4289 (N_4289,N_4165,N_4099);
nor U4290 (N_4290,N_4141,N_4087);
xor U4291 (N_4291,N_4079,N_4112);
and U4292 (N_4292,N_4059,N_4138);
nor U4293 (N_4293,N_4043,N_4161);
xor U4294 (N_4294,N_4026,N_4060);
or U4295 (N_4295,N_4022,N_4186);
nor U4296 (N_4296,N_4032,N_4119);
nor U4297 (N_4297,N_4135,N_4181);
or U4298 (N_4298,N_4028,N_4003);
nand U4299 (N_4299,N_4117,N_4006);
nand U4300 (N_4300,N_4028,N_4194);
xor U4301 (N_4301,N_4026,N_4044);
xor U4302 (N_4302,N_4164,N_4096);
and U4303 (N_4303,N_4187,N_4184);
nor U4304 (N_4304,N_4068,N_4194);
or U4305 (N_4305,N_4045,N_4042);
and U4306 (N_4306,N_4130,N_4109);
nor U4307 (N_4307,N_4092,N_4115);
xor U4308 (N_4308,N_4169,N_4080);
or U4309 (N_4309,N_4078,N_4023);
and U4310 (N_4310,N_4186,N_4035);
xor U4311 (N_4311,N_4156,N_4100);
xnor U4312 (N_4312,N_4101,N_4169);
xor U4313 (N_4313,N_4152,N_4080);
or U4314 (N_4314,N_4088,N_4155);
and U4315 (N_4315,N_4007,N_4108);
nand U4316 (N_4316,N_4179,N_4081);
nand U4317 (N_4317,N_4106,N_4123);
nor U4318 (N_4318,N_4136,N_4087);
xnor U4319 (N_4319,N_4151,N_4118);
nand U4320 (N_4320,N_4178,N_4002);
nor U4321 (N_4321,N_4068,N_4062);
or U4322 (N_4322,N_4074,N_4095);
nor U4323 (N_4323,N_4137,N_4041);
nand U4324 (N_4324,N_4137,N_4079);
xnor U4325 (N_4325,N_4021,N_4087);
and U4326 (N_4326,N_4110,N_4186);
nand U4327 (N_4327,N_4114,N_4117);
xnor U4328 (N_4328,N_4024,N_4156);
nand U4329 (N_4329,N_4049,N_4077);
and U4330 (N_4330,N_4073,N_4058);
or U4331 (N_4331,N_4037,N_4028);
or U4332 (N_4332,N_4044,N_4196);
nor U4333 (N_4333,N_4027,N_4061);
and U4334 (N_4334,N_4123,N_4037);
or U4335 (N_4335,N_4022,N_4072);
xor U4336 (N_4336,N_4155,N_4174);
nand U4337 (N_4337,N_4082,N_4156);
nor U4338 (N_4338,N_4046,N_4168);
and U4339 (N_4339,N_4064,N_4166);
nand U4340 (N_4340,N_4113,N_4058);
nand U4341 (N_4341,N_4116,N_4094);
xor U4342 (N_4342,N_4173,N_4008);
or U4343 (N_4343,N_4046,N_4197);
xor U4344 (N_4344,N_4029,N_4013);
xnor U4345 (N_4345,N_4054,N_4094);
xnor U4346 (N_4346,N_4038,N_4095);
and U4347 (N_4347,N_4134,N_4016);
nand U4348 (N_4348,N_4007,N_4184);
and U4349 (N_4349,N_4082,N_4122);
or U4350 (N_4350,N_4100,N_4166);
or U4351 (N_4351,N_4176,N_4142);
or U4352 (N_4352,N_4198,N_4140);
xnor U4353 (N_4353,N_4139,N_4179);
nand U4354 (N_4354,N_4139,N_4155);
nand U4355 (N_4355,N_4077,N_4097);
or U4356 (N_4356,N_4036,N_4072);
and U4357 (N_4357,N_4169,N_4081);
nand U4358 (N_4358,N_4034,N_4093);
and U4359 (N_4359,N_4132,N_4108);
xnor U4360 (N_4360,N_4055,N_4018);
or U4361 (N_4361,N_4033,N_4116);
or U4362 (N_4362,N_4140,N_4134);
nand U4363 (N_4363,N_4016,N_4159);
and U4364 (N_4364,N_4029,N_4142);
nor U4365 (N_4365,N_4143,N_4017);
nor U4366 (N_4366,N_4169,N_4147);
nor U4367 (N_4367,N_4136,N_4108);
xor U4368 (N_4368,N_4068,N_4009);
xor U4369 (N_4369,N_4165,N_4077);
or U4370 (N_4370,N_4082,N_4086);
nor U4371 (N_4371,N_4011,N_4083);
nor U4372 (N_4372,N_4036,N_4046);
nor U4373 (N_4373,N_4049,N_4004);
nand U4374 (N_4374,N_4157,N_4032);
and U4375 (N_4375,N_4024,N_4164);
and U4376 (N_4376,N_4172,N_4159);
nor U4377 (N_4377,N_4024,N_4134);
or U4378 (N_4378,N_4014,N_4123);
and U4379 (N_4379,N_4198,N_4156);
xor U4380 (N_4380,N_4182,N_4099);
nand U4381 (N_4381,N_4047,N_4043);
xnor U4382 (N_4382,N_4124,N_4104);
or U4383 (N_4383,N_4156,N_4007);
nor U4384 (N_4384,N_4083,N_4035);
nand U4385 (N_4385,N_4083,N_4165);
xnor U4386 (N_4386,N_4004,N_4059);
and U4387 (N_4387,N_4064,N_4169);
nand U4388 (N_4388,N_4131,N_4035);
and U4389 (N_4389,N_4028,N_4022);
nor U4390 (N_4390,N_4150,N_4152);
or U4391 (N_4391,N_4139,N_4112);
xnor U4392 (N_4392,N_4157,N_4134);
or U4393 (N_4393,N_4095,N_4194);
and U4394 (N_4394,N_4179,N_4059);
xnor U4395 (N_4395,N_4099,N_4057);
or U4396 (N_4396,N_4011,N_4012);
xor U4397 (N_4397,N_4169,N_4046);
xnor U4398 (N_4398,N_4188,N_4155);
nor U4399 (N_4399,N_4101,N_4091);
or U4400 (N_4400,N_4313,N_4214);
or U4401 (N_4401,N_4340,N_4366);
nand U4402 (N_4402,N_4234,N_4297);
xnor U4403 (N_4403,N_4223,N_4247);
or U4404 (N_4404,N_4376,N_4242);
nand U4405 (N_4405,N_4211,N_4341);
nand U4406 (N_4406,N_4374,N_4215);
nand U4407 (N_4407,N_4267,N_4385);
or U4408 (N_4408,N_4381,N_4253);
xor U4409 (N_4409,N_4369,N_4265);
and U4410 (N_4410,N_4316,N_4318);
nor U4411 (N_4411,N_4353,N_4302);
and U4412 (N_4412,N_4218,N_4217);
nor U4413 (N_4413,N_4288,N_4207);
nor U4414 (N_4414,N_4382,N_4326);
or U4415 (N_4415,N_4263,N_4268);
and U4416 (N_4416,N_4256,N_4232);
nor U4417 (N_4417,N_4249,N_4311);
xnor U4418 (N_4418,N_4283,N_4222);
or U4419 (N_4419,N_4252,N_4202);
nor U4420 (N_4420,N_4208,N_4379);
and U4421 (N_4421,N_4260,N_4261);
xnor U4422 (N_4422,N_4329,N_4350);
xor U4423 (N_4423,N_4317,N_4287);
nor U4424 (N_4424,N_4301,N_4310);
nand U4425 (N_4425,N_4282,N_4266);
nand U4426 (N_4426,N_4354,N_4306);
xor U4427 (N_4427,N_4216,N_4355);
or U4428 (N_4428,N_4264,N_4240);
nand U4429 (N_4429,N_4276,N_4281);
nor U4430 (N_4430,N_4221,N_4321);
xor U4431 (N_4431,N_4298,N_4206);
or U4432 (N_4432,N_4325,N_4258);
nor U4433 (N_4433,N_4314,N_4320);
xor U4434 (N_4434,N_4323,N_4322);
nor U4435 (N_4435,N_4271,N_4277);
xor U4436 (N_4436,N_4229,N_4349);
and U4437 (N_4437,N_4358,N_4336);
and U4438 (N_4438,N_4251,N_4227);
xnor U4439 (N_4439,N_4332,N_4371);
xor U4440 (N_4440,N_4289,N_4299);
nor U4441 (N_4441,N_4231,N_4334);
or U4442 (N_4442,N_4384,N_4209);
xor U4443 (N_4443,N_4273,N_4233);
nand U4444 (N_4444,N_4248,N_4370);
and U4445 (N_4445,N_4361,N_4360);
xor U4446 (N_4446,N_4303,N_4312);
nor U4447 (N_4447,N_4324,N_4399);
and U4448 (N_4448,N_4393,N_4274);
nand U4449 (N_4449,N_4278,N_4285);
nand U4450 (N_4450,N_4356,N_4389);
and U4451 (N_4451,N_4383,N_4396);
nor U4452 (N_4452,N_4330,N_4308);
xnor U4453 (N_4453,N_4262,N_4337);
or U4454 (N_4454,N_4254,N_4394);
nand U4455 (N_4455,N_4204,N_4269);
or U4456 (N_4456,N_4275,N_4398);
nand U4457 (N_4457,N_4375,N_4225);
nor U4458 (N_4458,N_4357,N_4280);
or U4459 (N_4459,N_4345,N_4377);
and U4460 (N_4460,N_4362,N_4338);
xnor U4461 (N_4461,N_4388,N_4296);
nor U4462 (N_4462,N_4238,N_4328);
nor U4463 (N_4463,N_4241,N_4305);
or U4464 (N_4464,N_4351,N_4307);
nor U4465 (N_4465,N_4364,N_4331);
nor U4466 (N_4466,N_4294,N_4348);
and U4467 (N_4467,N_4201,N_4200);
nand U4468 (N_4468,N_4284,N_4342);
nand U4469 (N_4469,N_4397,N_4212);
or U4470 (N_4470,N_4228,N_4239);
or U4471 (N_4471,N_4290,N_4395);
or U4472 (N_4472,N_4220,N_4270);
or U4473 (N_4473,N_4368,N_4259);
and U4474 (N_4474,N_4327,N_4315);
or U4475 (N_4475,N_4343,N_4244);
or U4476 (N_4476,N_4255,N_4279);
nor U4477 (N_4477,N_4205,N_4235);
or U4478 (N_4478,N_4257,N_4210);
nor U4479 (N_4479,N_4292,N_4224);
nand U4480 (N_4480,N_4295,N_4390);
nand U4481 (N_4481,N_4237,N_4243);
nand U4482 (N_4482,N_4286,N_4391);
nand U4483 (N_4483,N_4319,N_4300);
xor U4484 (N_4484,N_4272,N_4250);
nor U4485 (N_4485,N_4245,N_4339);
or U4486 (N_4486,N_4363,N_4372);
or U4487 (N_4487,N_4373,N_4378);
nand U4488 (N_4488,N_4304,N_4226);
or U4489 (N_4489,N_4203,N_4386);
xor U4490 (N_4490,N_4346,N_4309);
xnor U4491 (N_4491,N_4219,N_4333);
nor U4492 (N_4492,N_4365,N_4347);
or U4493 (N_4493,N_4344,N_4291);
nor U4494 (N_4494,N_4352,N_4293);
nor U4495 (N_4495,N_4213,N_4335);
nand U4496 (N_4496,N_4236,N_4230);
or U4497 (N_4497,N_4387,N_4367);
xor U4498 (N_4498,N_4246,N_4359);
nor U4499 (N_4499,N_4392,N_4380);
or U4500 (N_4500,N_4366,N_4329);
or U4501 (N_4501,N_4240,N_4208);
nand U4502 (N_4502,N_4329,N_4298);
nor U4503 (N_4503,N_4240,N_4215);
nand U4504 (N_4504,N_4384,N_4255);
and U4505 (N_4505,N_4254,N_4398);
nand U4506 (N_4506,N_4324,N_4261);
nand U4507 (N_4507,N_4346,N_4254);
nor U4508 (N_4508,N_4325,N_4316);
nor U4509 (N_4509,N_4215,N_4276);
xnor U4510 (N_4510,N_4304,N_4360);
nand U4511 (N_4511,N_4263,N_4330);
xnor U4512 (N_4512,N_4394,N_4327);
nor U4513 (N_4513,N_4326,N_4243);
xor U4514 (N_4514,N_4343,N_4210);
or U4515 (N_4515,N_4236,N_4283);
and U4516 (N_4516,N_4330,N_4231);
nand U4517 (N_4517,N_4240,N_4377);
and U4518 (N_4518,N_4298,N_4217);
xor U4519 (N_4519,N_4314,N_4255);
nor U4520 (N_4520,N_4228,N_4357);
nor U4521 (N_4521,N_4277,N_4362);
or U4522 (N_4522,N_4334,N_4331);
xor U4523 (N_4523,N_4345,N_4340);
or U4524 (N_4524,N_4276,N_4342);
nand U4525 (N_4525,N_4215,N_4289);
xnor U4526 (N_4526,N_4387,N_4255);
nand U4527 (N_4527,N_4260,N_4379);
xor U4528 (N_4528,N_4204,N_4262);
nand U4529 (N_4529,N_4392,N_4292);
or U4530 (N_4530,N_4288,N_4267);
and U4531 (N_4531,N_4371,N_4314);
xor U4532 (N_4532,N_4267,N_4230);
or U4533 (N_4533,N_4232,N_4360);
and U4534 (N_4534,N_4263,N_4357);
and U4535 (N_4535,N_4342,N_4238);
and U4536 (N_4536,N_4240,N_4351);
xnor U4537 (N_4537,N_4218,N_4276);
nor U4538 (N_4538,N_4364,N_4257);
and U4539 (N_4539,N_4278,N_4204);
xor U4540 (N_4540,N_4371,N_4271);
and U4541 (N_4541,N_4356,N_4271);
or U4542 (N_4542,N_4258,N_4319);
and U4543 (N_4543,N_4394,N_4214);
nand U4544 (N_4544,N_4362,N_4270);
and U4545 (N_4545,N_4315,N_4388);
and U4546 (N_4546,N_4201,N_4230);
xor U4547 (N_4547,N_4364,N_4250);
and U4548 (N_4548,N_4241,N_4244);
nor U4549 (N_4549,N_4218,N_4307);
xnor U4550 (N_4550,N_4382,N_4297);
nor U4551 (N_4551,N_4260,N_4245);
nand U4552 (N_4552,N_4353,N_4377);
xor U4553 (N_4553,N_4248,N_4209);
xor U4554 (N_4554,N_4260,N_4227);
and U4555 (N_4555,N_4313,N_4241);
nor U4556 (N_4556,N_4203,N_4338);
nor U4557 (N_4557,N_4272,N_4338);
nor U4558 (N_4558,N_4335,N_4304);
nand U4559 (N_4559,N_4393,N_4275);
xor U4560 (N_4560,N_4353,N_4383);
and U4561 (N_4561,N_4252,N_4349);
nand U4562 (N_4562,N_4341,N_4253);
nand U4563 (N_4563,N_4316,N_4242);
and U4564 (N_4564,N_4296,N_4252);
xor U4565 (N_4565,N_4209,N_4217);
and U4566 (N_4566,N_4397,N_4332);
xor U4567 (N_4567,N_4310,N_4355);
or U4568 (N_4568,N_4274,N_4287);
nor U4569 (N_4569,N_4337,N_4255);
nor U4570 (N_4570,N_4316,N_4229);
and U4571 (N_4571,N_4238,N_4207);
or U4572 (N_4572,N_4217,N_4342);
or U4573 (N_4573,N_4357,N_4336);
or U4574 (N_4574,N_4226,N_4300);
nand U4575 (N_4575,N_4258,N_4306);
nor U4576 (N_4576,N_4327,N_4349);
nand U4577 (N_4577,N_4332,N_4328);
or U4578 (N_4578,N_4277,N_4258);
xnor U4579 (N_4579,N_4215,N_4383);
and U4580 (N_4580,N_4374,N_4203);
nand U4581 (N_4581,N_4330,N_4316);
or U4582 (N_4582,N_4351,N_4206);
xor U4583 (N_4583,N_4267,N_4374);
nor U4584 (N_4584,N_4252,N_4271);
nand U4585 (N_4585,N_4223,N_4206);
and U4586 (N_4586,N_4272,N_4379);
xor U4587 (N_4587,N_4299,N_4205);
or U4588 (N_4588,N_4339,N_4230);
nor U4589 (N_4589,N_4252,N_4393);
nand U4590 (N_4590,N_4298,N_4343);
and U4591 (N_4591,N_4353,N_4380);
nor U4592 (N_4592,N_4264,N_4222);
nand U4593 (N_4593,N_4260,N_4299);
nand U4594 (N_4594,N_4309,N_4382);
nand U4595 (N_4595,N_4243,N_4232);
and U4596 (N_4596,N_4373,N_4254);
nor U4597 (N_4597,N_4343,N_4325);
or U4598 (N_4598,N_4345,N_4223);
nand U4599 (N_4599,N_4398,N_4246);
xor U4600 (N_4600,N_4532,N_4422);
or U4601 (N_4601,N_4551,N_4491);
xor U4602 (N_4602,N_4563,N_4572);
nor U4603 (N_4603,N_4454,N_4521);
and U4604 (N_4604,N_4407,N_4449);
xor U4605 (N_4605,N_4588,N_4584);
or U4606 (N_4606,N_4536,N_4444);
nand U4607 (N_4607,N_4587,N_4419);
or U4608 (N_4608,N_4544,N_4425);
nand U4609 (N_4609,N_4540,N_4562);
nand U4610 (N_4610,N_4408,N_4429);
xor U4611 (N_4611,N_4501,N_4576);
nand U4612 (N_4612,N_4525,N_4534);
xor U4613 (N_4613,N_4508,N_4446);
or U4614 (N_4614,N_4568,N_4402);
or U4615 (N_4615,N_4537,N_4533);
xor U4616 (N_4616,N_4528,N_4546);
nand U4617 (N_4617,N_4595,N_4490);
nor U4618 (N_4618,N_4498,N_4535);
nor U4619 (N_4619,N_4549,N_4493);
xnor U4620 (N_4620,N_4413,N_4478);
nand U4621 (N_4621,N_4529,N_4497);
xor U4622 (N_4622,N_4488,N_4565);
or U4623 (N_4623,N_4416,N_4482);
or U4624 (N_4624,N_4561,N_4530);
nor U4625 (N_4625,N_4404,N_4558);
nand U4626 (N_4626,N_4445,N_4513);
xnor U4627 (N_4627,N_4462,N_4585);
nand U4628 (N_4628,N_4505,N_4567);
and U4629 (N_4629,N_4423,N_4410);
nor U4630 (N_4630,N_4455,N_4420);
nand U4631 (N_4631,N_4571,N_4476);
or U4632 (N_4632,N_4443,N_4448);
and U4633 (N_4633,N_4502,N_4479);
nand U4634 (N_4634,N_4578,N_4465);
or U4635 (N_4635,N_4450,N_4557);
nor U4636 (N_4636,N_4519,N_4543);
and U4637 (N_4637,N_4492,N_4453);
nor U4638 (N_4638,N_4415,N_4593);
nand U4639 (N_4639,N_4426,N_4460);
and U4640 (N_4640,N_4589,N_4506);
nand U4641 (N_4641,N_4542,N_4470);
nor U4642 (N_4642,N_4417,N_4555);
xnor U4643 (N_4643,N_4489,N_4494);
nor U4644 (N_4644,N_4548,N_4487);
nand U4645 (N_4645,N_4512,N_4523);
or U4646 (N_4646,N_4586,N_4428);
and U4647 (N_4647,N_4499,N_4597);
nand U4648 (N_4648,N_4475,N_4468);
nor U4649 (N_4649,N_4591,N_4435);
or U4650 (N_4650,N_4507,N_4522);
and U4651 (N_4651,N_4447,N_4431);
and U4652 (N_4652,N_4594,N_4466);
or U4653 (N_4653,N_4458,N_4421);
and U4654 (N_4654,N_4592,N_4436);
nand U4655 (N_4655,N_4559,N_4411);
or U4656 (N_4656,N_4485,N_4496);
nand U4657 (N_4657,N_4439,N_4517);
and U4658 (N_4658,N_4554,N_4583);
xor U4659 (N_4659,N_4527,N_4550);
xor U4660 (N_4660,N_4486,N_4471);
nor U4661 (N_4661,N_4577,N_4509);
nand U4662 (N_4662,N_4541,N_4472);
or U4663 (N_4663,N_4504,N_4469);
or U4664 (N_4664,N_4500,N_4432);
xnor U4665 (N_4665,N_4456,N_4599);
or U4666 (N_4666,N_4480,N_4539);
or U4667 (N_4667,N_4405,N_4545);
and U4668 (N_4668,N_4459,N_4463);
nor U4669 (N_4669,N_4427,N_4495);
or U4670 (N_4670,N_4598,N_4516);
nand U4671 (N_4671,N_4538,N_4574);
and U4672 (N_4672,N_4573,N_4414);
nand U4673 (N_4673,N_4452,N_4409);
or U4674 (N_4674,N_4434,N_4582);
nand U4675 (N_4675,N_4457,N_4483);
or U4676 (N_4676,N_4556,N_4590);
nor U4677 (N_4677,N_4560,N_4520);
nor U4678 (N_4678,N_4518,N_4467);
nand U4679 (N_4679,N_4514,N_4503);
nand U4680 (N_4680,N_4400,N_4481);
nand U4681 (N_4681,N_4403,N_4406);
xnor U4682 (N_4682,N_4437,N_4570);
and U4683 (N_4683,N_4510,N_4412);
nand U4684 (N_4684,N_4418,N_4579);
and U4685 (N_4685,N_4440,N_4581);
nand U4686 (N_4686,N_4424,N_4547);
or U4687 (N_4687,N_4596,N_4461);
or U4688 (N_4688,N_4430,N_4524);
or U4689 (N_4689,N_4552,N_4442);
nor U4690 (N_4690,N_4484,N_4553);
nand U4691 (N_4691,N_4511,N_4451);
xnor U4692 (N_4692,N_4438,N_4575);
or U4693 (N_4693,N_4473,N_4526);
and U4694 (N_4694,N_4433,N_4580);
nor U4695 (N_4695,N_4564,N_4441);
or U4696 (N_4696,N_4474,N_4515);
nand U4697 (N_4697,N_4569,N_4566);
xnor U4698 (N_4698,N_4401,N_4477);
nand U4699 (N_4699,N_4464,N_4531);
nand U4700 (N_4700,N_4479,N_4408);
and U4701 (N_4701,N_4445,N_4529);
nor U4702 (N_4702,N_4533,N_4528);
and U4703 (N_4703,N_4427,N_4454);
or U4704 (N_4704,N_4588,N_4519);
or U4705 (N_4705,N_4464,N_4513);
and U4706 (N_4706,N_4587,N_4500);
or U4707 (N_4707,N_4522,N_4510);
nand U4708 (N_4708,N_4517,N_4574);
xor U4709 (N_4709,N_4548,N_4489);
xor U4710 (N_4710,N_4543,N_4440);
nor U4711 (N_4711,N_4449,N_4442);
xnor U4712 (N_4712,N_4481,N_4588);
xor U4713 (N_4713,N_4568,N_4473);
and U4714 (N_4714,N_4463,N_4492);
nand U4715 (N_4715,N_4497,N_4586);
and U4716 (N_4716,N_4438,N_4557);
nor U4717 (N_4717,N_4562,N_4566);
and U4718 (N_4718,N_4521,N_4502);
and U4719 (N_4719,N_4473,N_4558);
nor U4720 (N_4720,N_4593,N_4511);
and U4721 (N_4721,N_4445,N_4476);
xnor U4722 (N_4722,N_4536,N_4437);
nand U4723 (N_4723,N_4409,N_4537);
nor U4724 (N_4724,N_4567,N_4486);
xnor U4725 (N_4725,N_4415,N_4559);
and U4726 (N_4726,N_4593,N_4499);
or U4727 (N_4727,N_4451,N_4476);
xor U4728 (N_4728,N_4532,N_4408);
nand U4729 (N_4729,N_4505,N_4443);
or U4730 (N_4730,N_4588,N_4528);
or U4731 (N_4731,N_4589,N_4463);
nand U4732 (N_4732,N_4559,N_4495);
xnor U4733 (N_4733,N_4485,N_4449);
nand U4734 (N_4734,N_4454,N_4411);
xnor U4735 (N_4735,N_4473,N_4458);
nor U4736 (N_4736,N_4440,N_4432);
xor U4737 (N_4737,N_4446,N_4509);
xnor U4738 (N_4738,N_4599,N_4479);
xnor U4739 (N_4739,N_4407,N_4436);
or U4740 (N_4740,N_4594,N_4438);
nand U4741 (N_4741,N_4464,N_4535);
nor U4742 (N_4742,N_4519,N_4488);
xnor U4743 (N_4743,N_4576,N_4442);
nor U4744 (N_4744,N_4562,N_4517);
nand U4745 (N_4745,N_4546,N_4420);
or U4746 (N_4746,N_4446,N_4497);
nor U4747 (N_4747,N_4590,N_4595);
nor U4748 (N_4748,N_4444,N_4453);
or U4749 (N_4749,N_4509,N_4526);
nand U4750 (N_4750,N_4511,N_4422);
or U4751 (N_4751,N_4583,N_4543);
or U4752 (N_4752,N_4473,N_4495);
or U4753 (N_4753,N_4585,N_4446);
nor U4754 (N_4754,N_4579,N_4472);
nand U4755 (N_4755,N_4531,N_4479);
nand U4756 (N_4756,N_4489,N_4519);
or U4757 (N_4757,N_4419,N_4593);
nor U4758 (N_4758,N_4496,N_4424);
nand U4759 (N_4759,N_4528,N_4477);
and U4760 (N_4760,N_4403,N_4447);
nand U4761 (N_4761,N_4577,N_4403);
nand U4762 (N_4762,N_4526,N_4488);
and U4763 (N_4763,N_4479,N_4462);
and U4764 (N_4764,N_4596,N_4464);
nor U4765 (N_4765,N_4502,N_4584);
and U4766 (N_4766,N_4578,N_4416);
and U4767 (N_4767,N_4480,N_4582);
nand U4768 (N_4768,N_4571,N_4544);
nor U4769 (N_4769,N_4561,N_4455);
and U4770 (N_4770,N_4441,N_4517);
and U4771 (N_4771,N_4531,N_4556);
nor U4772 (N_4772,N_4583,N_4432);
nor U4773 (N_4773,N_4587,N_4497);
or U4774 (N_4774,N_4441,N_4581);
nand U4775 (N_4775,N_4575,N_4555);
xnor U4776 (N_4776,N_4532,N_4403);
nor U4777 (N_4777,N_4413,N_4428);
xnor U4778 (N_4778,N_4415,N_4406);
nor U4779 (N_4779,N_4588,N_4429);
nand U4780 (N_4780,N_4587,N_4516);
and U4781 (N_4781,N_4496,N_4404);
nor U4782 (N_4782,N_4566,N_4456);
nor U4783 (N_4783,N_4559,N_4450);
xor U4784 (N_4784,N_4441,N_4499);
or U4785 (N_4785,N_4431,N_4444);
or U4786 (N_4786,N_4592,N_4509);
nand U4787 (N_4787,N_4437,N_4566);
and U4788 (N_4788,N_4466,N_4501);
or U4789 (N_4789,N_4503,N_4467);
or U4790 (N_4790,N_4557,N_4402);
xnor U4791 (N_4791,N_4559,N_4552);
nand U4792 (N_4792,N_4594,N_4450);
nor U4793 (N_4793,N_4481,N_4520);
and U4794 (N_4794,N_4429,N_4470);
or U4795 (N_4795,N_4477,N_4593);
or U4796 (N_4796,N_4432,N_4495);
nor U4797 (N_4797,N_4449,N_4551);
nand U4798 (N_4798,N_4481,N_4521);
xnor U4799 (N_4799,N_4496,N_4412);
and U4800 (N_4800,N_4696,N_4622);
or U4801 (N_4801,N_4749,N_4635);
nand U4802 (N_4802,N_4674,N_4743);
and U4803 (N_4803,N_4692,N_4615);
or U4804 (N_4804,N_4764,N_4779);
nor U4805 (N_4805,N_4755,N_4753);
or U4806 (N_4806,N_4799,N_4678);
or U4807 (N_4807,N_4687,N_4617);
nand U4808 (N_4808,N_4688,N_4611);
and U4809 (N_4809,N_4715,N_4760);
or U4810 (N_4810,N_4654,N_4709);
and U4811 (N_4811,N_4768,N_4708);
nor U4812 (N_4812,N_4681,N_4778);
nor U4813 (N_4813,N_4607,N_4682);
or U4814 (N_4814,N_4649,N_4792);
nand U4815 (N_4815,N_4741,N_4765);
xor U4816 (N_4816,N_4699,N_4746);
nand U4817 (N_4817,N_4603,N_4773);
and U4818 (N_4818,N_4656,N_4659);
nand U4819 (N_4819,N_4723,N_4724);
nor U4820 (N_4820,N_4610,N_4677);
nand U4821 (N_4821,N_4721,N_4780);
and U4822 (N_4822,N_4706,N_4672);
nor U4823 (N_4823,N_4662,N_4619);
xor U4824 (N_4824,N_4733,N_4796);
nand U4825 (N_4825,N_4614,N_4790);
and U4826 (N_4826,N_4655,N_4673);
or U4827 (N_4827,N_4663,N_4713);
xor U4828 (N_4828,N_4618,N_4664);
nor U4829 (N_4829,N_4728,N_4629);
or U4830 (N_4830,N_4684,N_4758);
xor U4831 (N_4831,N_4665,N_4798);
or U4832 (N_4832,N_4602,N_4627);
nor U4833 (N_4833,N_4704,N_4707);
nand U4834 (N_4834,N_4786,N_4769);
nor U4835 (N_4835,N_4797,N_4642);
nand U4836 (N_4836,N_4734,N_4772);
nand U4837 (N_4837,N_4717,N_4703);
nand U4838 (N_4838,N_4620,N_4625);
nor U4839 (N_4839,N_4752,N_4700);
or U4840 (N_4840,N_4727,N_4714);
nor U4841 (N_4841,N_4631,N_4770);
or U4842 (N_4842,N_4777,N_4757);
or U4843 (N_4843,N_4771,N_4609);
nand U4844 (N_4844,N_4716,N_4787);
and U4845 (N_4845,N_4647,N_4701);
or U4846 (N_4846,N_4686,N_4621);
and U4847 (N_4847,N_4628,N_4794);
xor U4848 (N_4848,N_4657,N_4766);
nand U4849 (N_4849,N_4637,N_4775);
xor U4850 (N_4850,N_4683,N_4652);
nor U4851 (N_4851,N_4605,N_4623);
and U4852 (N_4852,N_4633,N_4740);
nand U4853 (N_4853,N_4651,N_4630);
and U4854 (N_4854,N_4650,N_4616);
xnor U4855 (N_4855,N_4648,N_4784);
nand U4856 (N_4856,N_4751,N_4667);
nor U4857 (N_4857,N_4712,N_4626);
nor U4858 (N_4858,N_4735,N_4782);
and U4859 (N_4859,N_4785,N_4731);
and U4860 (N_4860,N_4710,N_4754);
nand U4861 (N_4861,N_4601,N_4644);
nand U4862 (N_4862,N_4689,N_4685);
xor U4863 (N_4863,N_4679,N_4675);
xor U4864 (N_4864,N_4747,N_4756);
and U4865 (N_4865,N_4776,N_4763);
xor U4866 (N_4866,N_4767,N_4634);
or U4867 (N_4867,N_4729,N_4632);
and U4868 (N_4868,N_4781,N_4697);
or U4869 (N_4869,N_4666,N_4739);
nand U4870 (N_4870,N_4789,N_4624);
nand U4871 (N_4871,N_4705,N_4608);
nand U4872 (N_4872,N_4744,N_4718);
xor U4873 (N_4873,N_4736,N_4730);
nand U4874 (N_4874,N_4661,N_4646);
and U4875 (N_4875,N_4711,N_4774);
xnor U4876 (N_4876,N_4761,N_4791);
nand U4877 (N_4877,N_4720,N_4676);
nand U4878 (N_4878,N_4606,N_4671);
or U4879 (N_4879,N_4750,N_4638);
and U4880 (N_4880,N_4640,N_4738);
nand U4881 (N_4881,N_4613,N_4795);
nor U4882 (N_4882,N_4722,N_4612);
or U4883 (N_4883,N_4742,N_4748);
nand U4884 (N_4884,N_4762,N_4732);
and U4885 (N_4885,N_4783,N_4793);
and U4886 (N_4886,N_4645,N_4737);
nor U4887 (N_4887,N_4643,N_4690);
xnor U4888 (N_4888,N_4725,N_4745);
and U4889 (N_4889,N_4694,N_4600);
nor U4890 (N_4890,N_4641,N_4658);
xor U4891 (N_4891,N_4668,N_4680);
nand U4892 (N_4892,N_4669,N_4702);
nand U4893 (N_4893,N_4698,N_4636);
xor U4894 (N_4894,N_4670,N_4695);
or U4895 (N_4895,N_4719,N_4660);
or U4896 (N_4896,N_4691,N_4759);
nand U4897 (N_4897,N_4693,N_4653);
xnor U4898 (N_4898,N_4604,N_4788);
or U4899 (N_4899,N_4639,N_4726);
or U4900 (N_4900,N_4669,N_4793);
or U4901 (N_4901,N_4731,N_4770);
nand U4902 (N_4902,N_4712,N_4600);
xnor U4903 (N_4903,N_4775,N_4780);
or U4904 (N_4904,N_4690,N_4788);
xnor U4905 (N_4905,N_4647,N_4646);
or U4906 (N_4906,N_4692,N_4764);
xnor U4907 (N_4907,N_4630,N_4608);
or U4908 (N_4908,N_4694,N_4609);
or U4909 (N_4909,N_4694,N_4715);
xnor U4910 (N_4910,N_4666,N_4690);
xor U4911 (N_4911,N_4730,N_4674);
xnor U4912 (N_4912,N_4738,N_4718);
nand U4913 (N_4913,N_4794,N_4735);
or U4914 (N_4914,N_4670,N_4630);
and U4915 (N_4915,N_4710,N_4690);
nor U4916 (N_4916,N_4634,N_4667);
nor U4917 (N_4917,N_4722,N_4716);
and U4918 (N_4918,N_4630,N_4758);
nand U4919 (N_4919,N_4795,N_4698);
nor U4920 (N_4920,N_4767,N_4644);
xor U4921 (N_4921,N_4781,N_4616);
or U4922 (N_4922,N_4739,N_4686);
nand U4923 (N_4923,N_4766,N_4635);
or U4924 (N_4924,N_4705,N_4707);
and U4925 (N_4925,N_4694,N_4645);
or U4926 (N_4926,N_4665,N_4720);
xor U4927 (N_4927,N_4609,N_4687);
nor U4928 (N_4928,N_4662,N_4782);
or U4929 (N_4929,N_4689,N_4682);
xor U4930 (N_4930,N_4771,N_4718);
nand U4931 (N_4931,N_4625,N_4611);
or U4932 (N_4932,N_4615,N_4746);
or U4933 (N_4933,N_4707,N_4611);
nor U4934 (N_4934,N_4771,N_4779);
xor U4935 (N_4935,N_4621,N_4787);
or U4936 (N_4936,N_4786,N_4725);
and U4937 (N_4937,N_4717,N_4653);
nand U4938 (N_4938,N_4748,N_4612);
nor U4939 (N_4939,N_4759,N_4639);
or U4940 (N_4940,N_4731,N_4789);
and U4941 (N_4941,N_4698,N_4616);
nand U4942 (N_4942,N_4756,N_4796);
and U4943 (N_4943,N_4721,N_4723);
xnor U4944 (N_4944,N_4666,N_4616);
and U4945 (N_4945,N_4676,N_4779);
or U4946 (N_4946,N_4720,N_4672);
or U4947 (N_4947,N_4669,N_4795);
nor U4948 (N_4948,N_4781,N_4696);
nand U4949 (N_4949,N_4789,N_4736);
nand U4950 (N_4950,N_4795,N_4688);
nand U4951 (N_4951,N_4686,N_4669);
xnor U4952 (N_4952,N_4756,N_4692);
nand U4953 (N_4953,N_4797,N_4774);
xor U4954 (N_4954,N_4638,N_4631);
xor U4955 (N_4955,N_4718,N_4751);
nor U4956 (N_4956,N_4735,N_4753);
or U4957 (N_4957,N_4649,N_4743);
and U4958 (N_4958,N_4706,N_4689);
nand U4959 (N_4959,N_4771,N_4701);
nor U4960 (N_4960,N_4799,N_4642);
or U4961 (N_4961,N_4731,N_4623);
and U4962 (N_4962,N_4732,N_4670);
and U4963 (N_4963,N_4738,N_4798);
or U4964 (N_4964,N_4667,N_4699);
nor U4965 (N_4965,N_4678,N_4732);
xnor U4966 (N_4966,N_4760,N_4730);
or U4967 (N_4967,N_4757,N_4659);
or U4968 (N_4968,N_4796,N_4616);
and U4969 (N_4969,N_4705,N_4655);
nor U4970 (N_4970,N_4756,N_4799);
nor U4971 (N_4971,N_4614,N_4782);
nand U4972 (N_4972,N_4629,N_4741);
and U4973 (N_4973,N_4716,N_4742);
nand U4974 (N_4974,N_4766,N_4612);
and U4975 (N_4975,N_4620,N_4600);
xor U4976 (N_4976,N_4630,N_4665);
or U4977 (N_4977,N_4721,N_4604);
or U4978 (N_4978,N_4622,N_4670);
nand U4979 (N_4979,N_4695,N_4653);
and U4980 (N_4980,N_4602,N_4664);
and U4981 (N_4981,N_4778,N_4688);
or U4982 (N_4982,N_4769,N_4717);
nor U4983 (N_4983,N_4724,N_4736);
xnor U4984 (N_4984,N_4769,N_4624);
nor U4985 (N_4985,N_4767,N_4655);
nor U4986 (N_4986,N_4710,N_4717);
nand U4987 (N_4987,N_4645,N_4643);
nand U4988 (N_4988,N_4673,N_4770);
nand U4989 (N_4989,N_4751,N_4796);
nand U4990 (N_4990,N_4720,N_4636);
nand U4991 (N_4991,N_4625,N_4663);
nor U4992 (N_4992,N_4722,N_4726);
nor U4993 (N_4993,N_4652,N_4779);
or U4994 (N_4994,N_4712,N_4759);
or U4995 (N_4995,N_4711,N_4603);
or U4996 (N_4996,N_4638,N_4711);
and U4997 (N_4997,N_4711,N_4789);
or U4998 (N_4998,N_4614,N_4729);
and U4999 (N_4999,N_4714,N_4609);
nand UO_0 (O_0,N_4885,N_4809);
and UO_1 (O_1,N_4906,N_4917);
nand UO_2 (O_2,N_4932,N_4836);
nor UO_3 (O_3,N_4936,N_4852);
nand UO_4 (O_4,N_4958,N_4978);
nor UO_5 (O_5,N_4990,N_4831);
xnor UO_6 (O_6,N_4901,N_4878);
or UO_7 (O_7,N_4924,N_4876);
nand UO_8 (O_8,N_4972,N_4827);
or UO_9 (O_9,N_4947,N_4949);
nand UO_10 (O_10,N_4823,N_4940);
and UO_11 (O_11,N_4837,N_4986);
and UO_12 (O_12,N_4829,N_4839);
or UO_13 (O_13,N_4869,N_4900);
or UO_14 (O_14,N_4872,N_4842);
and UO_15 (O_15,N_4942,N_4925);
nand UO_16 (O_16,N_4930,N_4946);
nor UO_17 (O_17,N_4963,N_4887);
nor UO_18 (O_18,N_4902,N_4895);
nor UO_19 (O_19,N_4910,N_4985);
nor UO_20 (O_20,N_4992,N_4870);
nor UO_21 (O_21,N_4863,N_4886);
nand UO_22 (O_22,N_4998,N_4882);
xor UO_23 (O_23,N_4822,N_4899);
xor UO_24 (O_24,N_4953,N_4889);
nand UO_25 (O_25,N_4806,N_4974);
xnor UO_26 (O_26,N_4995,N_4982);
nand UO_27 (O_27,N_4832,N_4920);
and UO_28 (O_28,N_4989,N_4883);
nand UO_29 (O_29,N_4979,N_4981);
nand UO_30 (O_30,N_4977,N_4952);
nand UO_31 (O_31,N_4962,N_4879);
and UO_32 (O_32,N_4802,N_4996);
and UO_33 (O_33,N_4945,N_4987);
nand UO_34 (O_34,N_4815,N_4909);
nor UO_35 (O_35,N_4964,N_4824);
nor UO_36 (O_36,N_4817,N_4923);
or UO_37 (O_37,N_4954,N_4881);
or UO_38 (O_38,N_4904,N_4844);
or UO_39 (O_39,N_4926,N_4880);
nor UO_40 (O_40,N_4850,N_4834);
nor UO_41 (O_41,N_4847,N_4825);
and UO_42 (O_42,N_4907,N_4803);
or UO_43 (O_43,N_4905,N_4893);
or UO_44 (O_44,N_4833,N_4959);
nand UO_45 (O_45,N_4994,N_4931);
nand UO_46 (O_46,N_4939,N_4820);
nand UO_47 (O_47,N_4980,N_4911);
nor UO_48 (O_48,N_4968,N_4976);
or UO_49 (O_49,N_4805,N_4862);
xnor UO_50 (O_50,N_4961,N_4865);
or UO_51 (O_51,N_4848,N_4853);
nor UO_52 (O_52,N_4840,N_4816);
xor UO_53 (O_53,N_4922,N_4983);
xnor UO_54 (O_54,N_4935,N_4877);
or UO_55 (O_55,N_4871,N_4875);
nand UO_56 (O_56,N_4851,N_4971);
nor UO_57 (O_57,N_4898,N_4873);
or UO_58 (O_58,N_4908,N_4892);
or UO_59 (O_59,N_4858,N_4955);
or UO_60 (O_60,N_4903,N_4860);
or UO_61 (O_61,N_4843,N_4933);
nor UO_62 (O_62,N_4835,N_4966);
nand UO_63 (O_63,N_4800,N_4866);
nor UO_64 (O_64,N_4957,N_4944);
xnor UO_65 (O_65,N_4913,N_4801);
nand UO_66 (O_66,N_4819,N_4874);
and UO_67 (O_67,N_4894,N_4912);
xnor UO_68 (O_68,N_4970,N_4868);
nor UO_69 (O_69,N_4859,N_4967);
nor UO_70 (O_70,N_4896,N_4857);
or UO_71 (O_71,N_4956,N_4884);
and UO_72 (O_72,N_4846,N_4914);
nand UO_73 (O_73,N_4830,N_4804);
and UO_74 (O_74,N_4897,N_4973);
nand UO_75 (O_75,N_4861,N_4826);
or UO_76 (O_76,N_4807,N_4888);
and UO_77 (O_77,N_4960,N_4849);
xor UO_78 (O_78,N_4845,N_4934);
or UO_79 (O_79,N_4941,N_4821);
nor UO_80 (O_80,N_4915,N_4921);
or UO_81 (O_81,N_4818,N_4841);
xnor UO_82 (O_82,N_4991,N_4919);
or UO_83 (O_83,N_4812,N_4828);
and UO_84 (O_84,N_4891,N_4965);
nor UO_85 (O_85,N_4937,N_4808);
and UO_86 (O_86,N_4814,N_4948);
nor UO_87 (O_87,N_4854,N_4916);
xor UO_88 (O_88,N_4890,N_4855);
and UO_89 (O_89,N_4969,N_4811);
or UO_90 (O_90,N_4999,N_4943);
nand UO_91 (O_91,N_4938,N_4867);
or UO_92 (O_92,N_4984,N_4864);
or UO_93 (O_93,N_4838,N_4856);
nand UO_94 (O_94,N_4975,N_4929);
nand UO_95 (O_95,N_4928,N_4810);
or UO_96 (O_96,N_4988,N_4993);
or UO_97 (O_97,N_4918,N_4813);
nand UO_98 (O_98,N_4950,N_4997);
nor UO_99 (O_99,N_4927,N_4951);
nand UO_100 (O_100,N_4942,N_4872);
or UO_101 (O_101,N_4956,N_4856);
nor UO_102 (O_102,N_4882,N_4899);
and UO_103 (O_103,N_4995,N_4983);
or UO_104 (O_104,N_4838,N_4926);
xnor UO_105 (O_105,N_4896,N_4922);
or UO_106 (O_106,N_4858,N_4888);
nor UO_107 (O_107,N_4893,N_4958);
nand UO_108 (O_108,N_4889,N_4935);
and UO_109 (O_109,N_4869,N_4990);
nor UO_110 (O_110,N_4954,N_4885);
or UO_111 (O_111,N_4825,N_4916);
xor UO_112 (O_112,N_4853,N_4817);
or UO_113 (O_113,N_4818,N_4978);
and UO_114 (O_114,N_4866,N_4917);
xor UO_115 (O_115,N_4978,N_4905);
and UO_116 (O_116,N_4948,N_4908);
or UO_117 (O_117,N_4930,N_4876);
nor UO_118 (O_118,N_4961,N_4877);
xor UO_119 (O_119,N_4924,N_4913);
and UO_120 (O_120,N_4854,N_4805);
nand UO_121 (O_121,N_4919,N_4911);
nor UO_122 (O_122,N_4991,N_4993);
or UO_123 (O_123,N_4990,N_4899);
xnor UO_124 (O_124,N_4973,N_4979);
or UO_125 (O_125,N_4958,N_4982);
or UO_126 (O_126,N_4857,N_4838);
nand UO_127 (O_127,N_4998,N_4804);
and UO_128 (O_128,N_4905,N_4805);
nor UO_129 (O_129,N_4934,N_4889);
nand UO_130 (O_130,N_4902,N_4934);
and UO_131 (O_131,N_4978,N_4962);
nor UO_132 (O_132,N_4977,N_4908);
or UO_133 (O_133,N_4809,N_4972);
xor UO_134 (O_134,N_4818,N_4987);
nor UO_135 (O_135,N_4811,N_4866);
xor UO_136 (O_136,N_4850,N_4986);
xnor UO_137 (O_137,N_4962,N_4912);
and UO_138 (O_138,N_4963,N_4943);
and UO_139 (O_139,N_4992,N_4906);
nand UO_140 (O_140,N_4895,N_4976);
xnor UO_141 (O_141,N_4833,N_4937);
or UO_142 (O_142,N_4914,N_4994);
xor UO_143 (O_143,N_4900,N_4997);
nor UO_144 (O_144,N_4952,N_4925);
nand UO_145 (O_145,N_4814,N_4821);
nor UO_146 (O_146,N_4831,N_4842);
and UO_147 (O_147,N_4975,N_4879);
and UO_148 (O_148,N_4972,N_4860);
and UO_149 (O_149,N_4958,N_4962);
nand UO_150 (O_150,N_4982,N_4938);
nand UO_151 (O_151,N_4941,N_4829);
nor UO_152 (O_152,N_4957,N_4954);
xor UO_153 (O_153,N_4880,N_4854);
and UO_154 (O_154,N_4811,N_4858);
nand UO_155 (O_155,N_4880,N_4870);
nor UO_156 (O_156,N_4887,N_4908);
or UO_157 (O_157,N_4880,N_4839);
or UO_158 (O_158,N_4873,N_4817);
and UO_159 (O_159,N_4810,N_4938);
nor UO_160 (O_160,N_4805,N_4896);
or UO_161 (O_161,N_4840,N_4861);
xnor UO_162 (O_162,N_4829,N_4893);
nor UO_163 (O_163,N_4809,N_4961);
nand UO_164 (O_164,N_4802,N_4969);
or UO_165 (O_165,N_4989,N_4996);
xnor UO_166 (O_166,N_4938,N_4988);
nand UO_167 (O_167,N_4871,N_4836);
and UO_168 (O_168,N_4830,N_4864);
nand UO_169 (O_169,N_4835,N_4998);
and UO_170 (O_170,N_4874,N_4877);
xnor UO_171 (O_171,N_4994,N_4863);
nand UO_172 (O_172,N_4949,N_4922);
or UO_173 (O_173,N_4937,N_4849);
xnor UO_174 (O_174,N_4862,N_4843);
nand UO_175 (O_175,N_4969,N_4905);
nand UO_176 (O_176,N_4892,N_4841);
nor UO_177 (O_177,N_4916,N_4989);
nor UO_178 (O_178,N_4928,N_4847);
xnor UO_179 (O_179,N_4905,N_4890);
xnor UO_180 (O_180,N_4845,N_4977);
nor UO_181 (O_181,N_4924,N_4835);
and UO_182 (O_182,N_4888,N_4809);
nand UO_183 (O_183,N_4961,N_4895);
and UO_184 (O_184,N_4820,N_4862);
nor UO_185 (O_185,N_4907,N_4875);
and UO_186 (O_186,N_4909,N_4924);
and UO_187 (O_187,N_4936,N_4959);
nor UO_188 (O_188,N_4836,N_4915);
nor UO_189 (O_189,N_4881,N_4898);
nand UO_190 (O_190,N_4923,N_4836);
xnor UO_191 (O_191,N_4904,N_4815);
xnor UO_192 (O_192,N_4861,N_4972);
nor UO_193 (O_193,N_4944,N_4898);
or UO_194 (O_194,N_4841,N_4855);
nand UO_195 (O_195,N_4940,N_4816);
nand UO_196 (O_196,N_4821,N_4978);
or UO_197 (O_197,N_4914,N_4830);
and UO_198 (O_198,N_4878,N_4957);
nand UO_199 (O_199,N_4946,N_4815);
and UO_200 (O_200,N_4908,N_4989);
xnor UO_201 (O_201,N_4925,N_4809);
nor UO_202 (O_202,N_4846,N_4949);
or UO_203 (O_203,N_4842,N_4969);
nand UO_204 (O_204,N_4999,N_4969);
xor UO_205 (O_205,N_4961,N_4979);
nand UO_206 (O_206,N_4865,N_4949);
and UO_207 (O_207,N_4949,N_4837);
xnor UO_208 (O_208,N_4854,N_4852);
xor UO_209 (O_209,N_4999,N_4967);
and UO_210 (O_210,N_4879,N_4882);
nand UO_211 (O_211,N_4820,N_4998);
and UO_212 (O_212,N_4827,N_4849);
and UO_213 (O_213,N_4948,N_4834);
nand UO_214 (O_214,N_4833,N_4900);
xnor UO_215 (O_215,N_4863,N_4880);
and UO_216 (O_216,N_4883,N_4957);
and UO_217 (O_217,N_4927,N_4981);
and UO_218 (O_218,N_4871,N_4857);
and UO_219 (O_219,N_4923,N_4947);
nor UO_220 (O_220,N_4937,N_4938);
and UO_221 (O_221,N_4898,N_4952);
and UO_222 (O_222,N_4866,N_4830);
and UO_223 (O_223,N_4960,N_4844);
and UO_224 (O_224,N_4857,N_4800);
nand UO_225 (O_225,N_4825,N_4925);
xnor UO_226 (O_226,N_4886,N_4851);
nor UO_227 (O_227,N_4930,N_4962);
nand UO_228 (O_228,N_4808,N_4862);
nand UO_229 (O_229,N_4801,N_4831);
nand UO_230 (O_230,N_4965,N_4916);
nor UO_231 (O_231,N_4984,N_4835);
and UO_232 (O_232,N_4961,N_4843);
nand UO_233 (O_233,N_4917,N_4985);
nor UO_234 (O_234,N_4864,N_4832);
nor UO_235 (O_235,N_4991,N_4889);
xnor UO_236 (O_236,N_4909,N_4807);
nand UO_237 (O_237,N_4850,N_4898);
nor UO_238 (O_238,N_4972,N_4849);
and UO_239 (O_239,N_4883,N_4831);
or UO_240 (O_240,N_4955,N_4828);
xnor UO_241 (O_241,N_4815,N_4945);
nor UO_242 (O_242,N_4854,N_4807);
and UO_243 (O_243,N_4833,N_4899);
or UO_244 (O_244,N_4874,N_4902);
and UO_245 (O_245,N_4863,N_4856);
xor UO_246 (O_246,N_4830,N_4993);
nand UO_247 (O_247,N_4991,N_4910);
or UO_248 (O_248,N_4828,N_4977);
xor UO_249 (O_249,N_4854,N_4846);
nor UO_250 (O_250,N_4910,N_4900);
nor UO_251 (O_251,N_4901,N_4917);
nand UO_252 (O_252,N_4899,N_4823);
nor UO_253 (O_253,N_4937,N_4816);
nor UO_254 (O_254,N_4996,N_4935);
and UO_255 (O_255,N_4989,N_4925);
and UO_256 (O_256,N_4876,N_4801);
xor UO_257 (O_257,N_4995,N_4997);
and UO_258 (O_258,N_4996,N_4868);
or UO_259 (O_259,N_4930,N_4830);
and UO_260 (O_260,N_4956,N_4899);
xnor UO_261 (O_261,N_4819,N_4988);
and UO_262 (O_262,N_4859,N_4826);
and UO_263 (O_263,N_4845,N_4867);
or UO_264 (O_264,N_4959,N_4911);
nand UO_265 (O_265,N_4823,N_4951);
and UO_266 (O_266,N_4955,N_4872);
nor UO_267 (O_267,N_4946,N_4839);
or UO_268 (O_268,N_4979,N_4935);
nor UO_269 (O_269,N_4810,N_4920);
and UO_270 (O_270,N_4828,N_4951);
nor UO_271 (O_271,N_4997,N_4983);
xnor UO_272 (O_272,N_4896,N_4825);
nor UO_273 (O_273,N_4955,N_4878);
nand UO_274 (O_274,N_4841,N_4988);
or UO_275 (O_275,N_4826,N_4972);
and UO_276 (O_276,N_4998,N_4938);
nor UO_277 (O_277,N_4855,N_4935);
or UO_278 (O_278,N_4973,N_4826);
and UO_279 (O_279,N_4962,N_4800);
nor UO_280 (O_280,N_4828,N_4988);
and UO_281 (O_281,N_4964,N_4801);
nand UO_282 (O_282,N_4938,N_4913);
nor UO_283 (O_283,N_4963,N_4922);
or UO_284 (O_284,N_4965,N_4961);
xnor UO_285 (O_285,N_4875,N_4932);
xnor UO_286 (O_286,N_4973,N_4825);
xnor UO_287 (O_287,N_4829,N_4981);
or UO_288 (O_288,N_4911,N_4907);
nand UO_289 (O_289,N_4886,N_4921);
nand UO_290 (O_290,N_4943,N_4899);
nor UO_291 (O_291,N_4831,N_4910);
and UO_292 (O_292,N_4847,N_4802);
xor UO_293 (O_293,N_4873,N_4917);
and UO_294 (O_294,N_4889,N_4997);
nor UO_295 (O_295,N_4905,N_4870);
xor UO_296 (O_296,N_4950,N_4924);
nand UO_297 (O_297,N_4903,N_4951);
nand UO_298 (O_298,N_4925,N_4931);
nand UO_299 (O_299,N_4885,N_4909);
and UO_300 (O_300,N_4941,N_4855);
and UO_301 (O_301,N_4831,N_4911);
nor UO_302 (O_302,N_4829,N_4955);
xnor UO_303 (O_303,N_4903,N_4863);
xor UO_304 (O_304,N_4912,N_4917);
or UO_305 (O_305,N_4886,N_4996);
nor UO_306 (O_306,N_4917,N_4891);
or UO_307 (O_307,N_4980,N_4954);
or UO_308 (O_308,N_4910,N_4898);
or UO_309 (O_309,N_4982,N_4891);
nor UO_310 (O_310,N_4813,N_4949);
xor UO_311 (O_311,N_4872,N_4989);
nand UO_312 (O_312,N_4997,N_4886);
xor UO_313 (O_313,N_4815,N_4932);
nor UO_314 (O_314,N_4973,N_4951);
nand UO_315 (O_315,N_4949,N_4974);
and UO_316 (O_316,N_4889,N_4963);
nand UO_317 (O_317,N_4943,N_4888);
or UO_318 (O_318,N_4862,N_4884);
xnor UO_319 (O_319,N_4839,N_4975);
xnor UO_320 (O_320,N_4837,N_4969);
xnor UO_321 (O_321,N_4923,N_4934);
or UO_322 (O_322,N_4854,N_4850);
xor UO_323 (O_323,N_4865,N_4892);
or UO_324 (O_324,N_4952,N_4829);
or UO_325 (O_325,N_4896,N_4804);
xor UO_326 (O_326,N_4815,N_4846);
and UO_327 (O_327,N_4926,N_4967);
nor UO_328 (O_328,N_4835,N_4969);
or UO_329 (O_329,N_4886,N_4986);
and UO_330 (O_330,N_4849,N_4918);
nor UO_331 (O_331,N_4948,N_4963);
nor UO_332 (O_332,N_4894,N_4982);
nor UO_333 (O_333,N_4918,N_4854);
nand UO_334 (O_334,N_4990,N_4936);
and UO_335 (O_335,N_4928,N_4940);
nand UO_336 (O_336,N_4994,N_4944);
nor UO_337 (O_337,N_4883,N_4893);
nor UO_338 (O_338,N_4870,N_4817);
nor UO_339 (O_339,N_4804,N_4870);
nand UO_340 (O_340,N_4867,N_4969);
xnor UO_341 (O_341,N_4826,N_4820);
nor UO_342 (O_342,N_4892,N_4853);
or UO_343 (O_343,N_4889,N_4968);
or UO_344 (O_344,N_4882,N_4834);
and UO_345 (O_345,N_4894,N_4893);
and UO_346 (O_346,N_4985,N_4908);
and UO_347 (O_347,N_4862,N_4908);
nor UO_348 (O_348,N_4849,N_4840);
and UO_349 (O_349,N_4948,N_4940);
nand UO_350 (O_350,N_4837,N_4884);
xnor UO_351 (O_351,N_4874,N_4922);
nand UO_352 (O_352,N_4940,N_4835);
and UO_353 (O_353,N_4912,N_4828);
nand UO_354 (O_354,N_4820,N_4833);
and UO_355 (O_355,N_4846,N_4907);
or UO_356 (O_356,N_4874,N_4827);
xor UO_357 (O_357,N_4841,N_4806);
nor UO_358 (O_358,N_4875,N_4888);
nand UO_359 (O_359,N_4939,N_4940);
or UO_360 (O_360,N_4986,N_4883);
or UO_361 (O_361,N_4802,N_4815);
and UO_362 (O_362,N_4884,N_4902);
nand UO_363 (O_363,N_4904,N_4956);
nor UO_364 (O_364,N_4924,N_4947);
or UO_365 (O_365,N_4848,N_4852);
xnor UO_366 (O_366,N_4843,N_4996);
xnor UO_367 (O_367,N_4987,N_4879);
nand UO_368 (O_368,N_4830,N_4999);
or UO_369 (O_369,N_4936,N_4943);
or UO_370 (O_370,N_4939,N_4972);
xnor UO_371 (O_371,N_4866,N_4906);
and UO_372 (O_372,N_4981,N_4956);
xor UO_373 (O_373,N_4942,N_4860);
and UO_374 (O_374,N_4961,N_4836);
nor UO_375 (O_375,N_4940,N_4890);
and UO_376 (O_376,N_4851,N_4803);
xor UO_377 (O_377,N_4982,N_4997);
nand UO_378 (O_378,N_4995,N_4966);
nand UO_379 (O_379,N_4832,N_4940);
and UO_380 (O_380,N_4969,N_4968);
nor UO_381 (O_381,N_4847,N_4835);
nor UO_382 (O_382,N_4954,N_4877);
nand UO_383 (O_383,N_4849,N_4936);
or UO_384 (O_384,N_4856,N_4832);
and UO_385 (O_385,N_4887,N_4873);
xor UO_386 (O_386,N_4968,N_4982);
nor UO_387 (O_387,N_4997,N_4964);
nor UO_388 (O_388,N_4981,N_4851);
or UO_389 (O_389,N_4855,N_4834);
and UO_390 (O_390,N_4975,N_4832);
and UO_391 (O_391,N_4952,N_4813);
nor UO_392 (O_392,N_4984,N_4968);
xnor UO_393 (O_393,N_4962,N_4933);
and UO_394 (O_394,N_4839,N_4942);
nand UO_395 (O_395,N_4840,N_4969);
xnor UO_396 (O_396,N_4923,N_4801);
nor UO_397 (O_397,N_4933,N_4992);
nor UO_398 (O_398,N_4814,N_4999);
and UO_399 (O_399,N_4904,N_4906);
and UO_400 (O_400,N_4926,N_4929);
nor UO_401 (O_401,N_4804,N_4862);
nand UO_402 (O_402,N_4855,N_4962);
nor UO_403 (O_403,N_4892,N_4880);
or UO_404 (O_404,N_4993,N_4936);
nand UO_405 (O_405,N_4964,N_4841);
or UO_406 (O_406,N_4968,N_4869);
and UO_407 (O_407,N_4925,N_4921);
or UO_408 (O_408,N_4885,N_4998);
xor UO_409 (O_409,N_4814,N_4938);
nor UO_410 (O_410,N_4916,N_4945);
nand UO_411 (O_411,N_4849,N_4892);
nand UO_412 (O_412,N_4878,N_4978);
nor UO_413 (O_413,N_4853,N_4812);
nand UO_414 (O_414,N_4857,N_4962);
and UO_415 (O_415,N_4910,N_4826);
nor UO_416 (O_416,N_4830,N_4994);
or UO_417 (O_417,N_4896,N_4841);
and UO_418 (O_418,N_4843,N_4805);
xnor UO_419 (O_419,N_4872,N_4840);
nor UO_420 (O_420,N_4868,N_4921);
or UO_421 (O_421,N_4906,N_4905);
xor UO_422 (O_422,N_4831,N_4900);
or UO_423 (O_423,N_4961,N_4806);
nand UO_424 (O_424,N_4860,N_4950);
xnor UO_425 (O_425,N_4907,N_4848);
or UO_426 (O_426,N_4867,N_4812);
nor UO_427 (O_427,N_4864,N_4979);
xnor UO_428 (O_428,N_4833,N_4969);
or UO_429 (O_429,N_4863,N_4862);
nand UO_430 (O_430,N_4808,N_4972);
nand UO_431 (O_431,N_4833,N_4803);
or UO_432 (O_432,N_4901,N_4986);
or UO_433 (O_433,N_4928,N_4854);
nor UO_434 (O_434,N_4873,N_4901);
xnor UO_435 (O_435,N_4914,N_4967);
or UO_436 (O_436,N_4932,N_4856);
xor UO_437 (O_437,N_4973,N_4901);
or UO_438 (O_438,N_4846,N_4900);
nand UO_439 (O_439,N_4955,N_4850);
nand UO_440 (O_440,N_4937,N_4872);
and UO_441 (O_441,N_4938,N_4900);
xor UO_442 (O_442,N_4909,N_4952);
or UO_443 (O_443,N_4991,N_4837);
xnor UO_444 (O_444,N_4962,N_4953);
nand UO_445 (O_445,N_4896,N_4827);
nand UO_446 (O_446,N_4908,N_4939);
or UO_447 (O_447,N_4809,N_4862);
nor UO_448 (O_448,N_4991,N_4897);
xor UO_449 (O_449,N_4884,N_4887);
xor UO_450 (O_450,N_4935,N_4908);
and UO_451 (O_451,N_4958,N_4938);
and UO_452 (O_452,N_4871,N_4845);
nor UO_453 (O_453,N_4809,N_4852);
nor UO_454 (O_454,N_4938,N_4862);
and UO_455 (O_455,N_4834,N_4999);
and UO_456 (O_456,N_4825,N_4889);
and UO_457 (O_457,N_4820,N_4806);
or UO_458 (O_458,N_4804,N_4973);
nand UO_459 (O_459,N_4922,N_4826);
and UO_460 (O_460,N_4871,N_4907);
and UO_461 (O_461,N_4920,N_4892);
nor UO_462 (O_462,N_4975,N_4865);
nor UO_463 (O_463,N_4982,N_4833);
nor UO_464 (O_464,N_4973,N_4912);
or UO_465 (O_465,N_4972,N_4966);
and UO_466 (O_466,N_4970,N_4858);
nor UO_467 (O_467,N_4831,N_4835);
nor UO_468 (O_468,N_4992,N_4984);
and UO_469 (O_469,N_4874,N_4968);
and UO_470 (O_470,N_4865,N_4899);
nor UO_471 (O_471,N_4842,N_4829);
nand UO_472 (O_472,N_4810,N_4854);
and UO_473 (O_473,N_4894,N_4959);
nor UO_474 (O_474,N_4953,N_4915);
nand UO_475 (O_475,N_4905,N_4981);
nor UO_476 (O_476,N_4938,N_4918);
nor UO_477 (O_477,N_4800,N_4810);
nor UO_478 (O_478,N_4817,N_4859);
or UO_479 (O_479,N_4806,N_4977);
and UO_480 (O_480,N_4961,N_4838);
xnor UO_481 (O_481,N_4928,N_4980);
and UO_482 (O_482,N_4822,N_4948);
or UO_483 (O_483,N_4825,N_4812);
and UO_484 (O_484,N_4972,N_4990);
or UO_485 (O_485,N_4819,N_4953);
nor UO_486 (O_486,N_4971,N_4843);
and UO_487 (O_487,N_4952,N_4976);
nand UO_488 (O_488,N_4840,N_4995);
and UO_489 (O_489,N_4881,N_4828);
and UO_490 (O_490,N_4968,N_4922);
or UO_491 (O_491,N_4893,N_4813);
nand UO_492 (O_492,N_4992,N_4880);
nand UO_493 (O_493,N_4896,N_4883);
nor UO_494 (O_494,N_4872,N_4871);
nand UO_495 (O_495,N_4821,N_4801);
or UO_496 (O_496,N_4827,N_4933);
and UO_497 (O_497,N_4876,N_4915);
nand UO_498 (O_498,N_4830,N_4888);
nor UO_499 (O_499,N_4955,N_4824);
nor UO_500 (O_500,N_4953,N_4813);
nand UO_501 (O_501,N_4979,N_4948);
nor UO_502 (O_502,N_4809,N_4912);
and UO_503 (O_503,N_4827,N_4920);
nor UO_504 (O_504,N_4976,N_4979);
or UO_505 (O_505,N_4846,N_4919);
or UO_506 (O_506,N_4946,N_4952);
xnor UO_507 (O_507,N_4963,N_4817);
and UO_508 (O_508,N_4854,N_4888);
nand UO_509 (O_509,N_4970,N_4852);
and UO_510 (O_510,N_4912,N_4825);
nand UO_511 (O_511,N_4884,N_4879);
or UO_512 (O_512,N_4827,N_4939);
or UO_513 (O_513,N_4868,N_4836);
or UO_514 (O_514,N_4830,N_4983);
nor UO_515 (O_515,N_4926,N_4996);
xnor UO_516 (O_516,N_4828,N_4956);
xnor UO_517 (O_517,N_4942,N_4989);
nor UO_518 (O_518,N_4889,N_4816);
nand UO_519 (O_519,N_4882,N_4901);
or UO_520 (O_520,N_4904,N_4871);
or UO_521 (O_521,N_4950,N_4850);
nor UO_522 (O_522,N_4853,N_4865);
nor UO_523 (O_523,N_4822,N_4846);
or UO_524 (O_524,N_4895,N_4823);
and UO_525 (O_525,N_4837,N_4814);
and UO_526 (O_526,N_4913,N_4930);
and UO_527 (O_527,N_4979,N_4808);
and UO_528 (O_528,N_4806,N_4823);
xor UO_529 (O_529,N_4882,N_4822);
nand UO_530 (O_530,N_4979,N_4811);
xnor UO_531 (O_531,N_4932,N_4809);
nand UO_532 (O_532,N_4862,N_4824);
or UO_533 (O_533,N_4820,N_4838);
nand UO_534 (O_534,N_4976,N_4975);
xor UO_535 (O_535,N_4963,N_4843);
nand UO_536 (O_536,N_4939,N_4981);
and UO_537 (O_537,N_4844,N_4819);
xnor UO_538 (O_538,N_4943,N_4964);
or UO_539 (O_539,N_4924,N_4815);
or UO_540 (O_540,N_4886,N_4935);
nand UO_541 (O_541,N_4825,N_4900);
nor UO_542 (O_542,N_4871,N_4990);
nand UO_543 (O_543,N_4941,N_4859);
or UO_544 (O_544,N_4829,N_4865);
xor UO_545 (O_545,N_4828,N_4909);
and UO_546 (O_546,N_4958,N_4879);
nor UO_547 (O_547,N_4943,N_4993);
and UO_548 (O_548,N_4945,N_4824);
nand UO_549 (O_549,N_4835,N_4817);
nand UO_550 (O_550,N_4876,N_4986);
or UO_551 (O_551,N_4801,N_4961);
xor UO_552 (O_552,N_4949,N_4904);
nor UO_553 (O_553,N_4988,N_4911);
nor UO_554 (O_554,N_4899,N_4887);
nand UO_555 (O_555,N_4894,N_4857);
nand UO_556 (O_556,N_4919,N_4801);
xnor UO_557 (O_557,N_4898,N_4854);
nor UO_558 (O_558,N_4875,N_4817);
nand UO_559 (O_559,N_4905,N_4935);
and UO_560 (O_560,N_4908,N_4851);
and UO_561 (O_561,N_4804,N_4813);
xnor UO_562 (O_562,N_4909,N_4994);
nand UO_563 (O_563,N_4905,N_4887);
or UO_564 (O_564,N_4832,N_4812);
xor UO_565 (O_565,N_4973,N_4849);
or UO_566 (O_566,N_4950,N_4853);
or UO_567 (O_567,N_4857,N_4805);
nor UO_568 (O_568,N_4971,N_4865);
xnor UO_569 (O_569,N_4934,N_4857);
and UO_570 (O_570,N_4818,N_4839);
nor UO_571 (O_571,N_4858,N_4801);
and UO_572 (O_572,N_4865,N_4974);
and UO_573 (O_573,N_4946,N_4885);
xnor UO_574 (O_574,N_4830,N_4948);
and UO_575 (O_575,N_4840,N_4918);
and UO_576 (O_576,N_4930,N_4920);
xnor UO_577 (O_577,N_4924,N_4823);
and UO_578 (O_578,N_4856,N_4871);
nand UO_579 (O_579,N_4826,N_4810);
nand UO_580 (O_580,N_4945,N_4875);
xnor UO_581 (O_581,N_4984,N_4969);
xor UO_582 (O_582,N_4897,N_4965);
nand UO_583 (O_583,N_4971,N_4836);
or UO_584 (O_584,N_4803,N_4828);
nand UO_585 (O_585,N_4878,N_4908);
or UO_586 (O_586,N_4846,N_4837);
and UO_587 (O_587,N_4876,N_4866);
and UO_588 (O_588,N_4892,N_4879);
xor UO_589 (O_589,N_4906,N_4953);
nor UO_590 (O_590,N_4933,N_4862);
xnor UO_591 (O_591,N_4932,N_4937);
nor UO_592 (O_592,N_4923,N_4927);
and UO_593 (O_593,N_4989,N_4959);
and UO_594 (O_594,N_4992,N_4981);
nor UO_595 (O_595,N_4940,N_4828);
xnor UO_596 (O_596,N_4978,N_4969);
or UO_597 (O_597,N_4883,N_4971);
or UO_598 (O_598,N_4957,N_4937);
and UO_599 (O_599,N_4992,N_4803);
and UO_600 (O_600,N_4864,N_4856);
nor UO_601 (O_601,N_4921,N_4943);
nor UO_602 (O_602,N_4892,N_4977);
and UO_603 (O_603,N_4978,N_4935);
or UO_604 (O_604,N_4870,N_4987);
nand UO_605 (O_605,N_4882,N_4824);
xor UO_606 (O_606,N_4888,N_4939);
and UO_607 (O_607,N_4976,N_4969);
and UO_608 (O_608,N_4886,N_4936);
nor UO_609 (O_609,N_4870,N_4947);
or UO_610 (O_610,N_4808,N_4920);
or UO_611 (O_611,N_4823,N_4821);
or UO_612 (O_612,N_4956,N_4831);
or UO_613 (O_613,N_4808,N_4956);
or UO_614 (O_614,N_4999,N_4961);
and UO_615 (O_615,N_4952,N_4991);
xor UO_616 (O_616,N_4814,N_4918);
nor UO_617 (O_617,N_4817,N_4915);
or UO_618 (O_618,N_4873,N_4835);
xor UO_619 (O_619,N_4928,N_4927);
nand UO_620 (O_620,N_4931,N_4948);
and UO_621 (O_621,N_4945,N_4960);
nor UO_622 (O_622,N_4944,N_4863);
nor UO_623 (O_623,N_4924,N_4952);
nor UO_624 (O_624,N_4826,N_4834);
nand UO_625 (O_625,N_4930,N_4845);
or UO_626 (O_626,N_4825,N_4949);
xor UO_627 (O_627,N_4951,N_4933);
nor UO_628 (O_628,N_4971,N_4976);
and UO_629 (O_629,N_4971,N_4871);
or UO_630 (O_630,N_4836,N_4962);
xor UO_631 (O_631,N_4800,N_4851);
nor UO_632 (O_632,N_4937,N_4971);
nor UO_633 (O_633,N_4950,N_4843);
xnor UO_634 (O_634,N_4979,N_4933);
xnor UO_635 (O_635,N_4993,N_4954);
nand UO_636 (O_636,N_4823,N_4998);
nor UO_637 (O_637,N_4929,N_4974);
or UO_638 (O_638,N_4962,N_4942);
nand UO_639 (O_639,N_4991,N_4830);
and UO_640 (O_640,N_4869,N_4949);
or UO_641 (O_641,N_4806,N_4862);
xor UO_642 (O_642,N_4871,N_4963);
and UO_643 (O_643,N_4864,N_4801);
or UO_644 (O_644,N_4904,N_4986);
nand UO_645 (O_645,N_4805,N_4875);
and UO_646 (O_646,N_4899,N_4835);
and UO_647 (O_647,N_4887,N_4828);
nor UO_648 (O_648,N_4943,N_4989);
xor UO_649 (O_649,N_4821,N_4927);
and UO_650 (O_650,N_4894,N_4969);
and UO_651 (O_651,N_4911,N_4982);
nor UO_652 (O_652,N_4817,N_4809);
nand UO_653 (O_653,N_4880,N_4831);
nor UO_654 (O_654,N_4914,N_4861);
and UO_655 (O_655,N_4857,N_4935);
nand UO_656 (O_656,N_4876,N_4931);
xor UO_657 (O_657,N_4831,N_4813);
nand UO_658 (O_658,N_4886,N_4919);
nor UO_659 (O_659,N_4907,N_4807);
or UO_660 (O_660,N_4938,N_4824);
nand UO_661 (O_661,N_4904,N_4819);
nor UO_662 (O_662,N_4868,N_4838);
or UO_663 (O_663,N_4817,N_4897);
and UO_664 (O_664,N_4961,N_4908);
nand UO_665 (O_665,N_4832,N_4935);
xnor UO_666 (O_666,N_4834,N_4884);
xnor UO_667 (O_667,N_4866,N_4930);
and UO_668 (O_668,N_4932,N_4877);
and UO_669 (O_669,N_4914,N_4817);
nand UO_670 (O_670,N_4895,N_4905);
nor UO_671 (O_671,N_4909,N_4981);
nand UO_672 (O_672,N_4963,N_4960);
xor UO_673 (O_673,N_4827,N_4943);
and UO_674 (O_674,N_4840,N_4951);
and UO_675 (O_675,N_4831,N_4817);
nor UO_676 (O_676,N_4959,N_4934);
and UO_677 (O_677,N_4943,N_4816);
and UO_678 (O_678,N_4948,N_4866);
xnor UO_679 (O_679,N_4858,N_4922);
nor UO_680 (O_680,N_4834,N_4815);
xnor UO_681 (O_681,N_4869,N_4977);
xnor UO_682 (O_682,N_4938,N_4819);
nand UO_683 (O_683,N_4827,N_4969);
or UO_684 (O_684,N_4868,N_4881);
xor UO_685 (O_685,N_4850,N_4983);
or UO_686 (O_686,N_4859,N_4898);
nand UO_687 (O_687,N_4922,N_4905);
or UO_688 (O_688,N_4962,N_4893);
and UO_689 (O_689,N_4976,N_4851);
xnor UO_690 (O_690,N_4955,N_4869);
nor UO_691 (O_691,N_4822,N_4921);
and UO_692 (O_692,N_4943,N_4976);
xnor UO_693 (O_693,N_4995,N_4934);
or UO_694 (O_694,N_4820,N_4976);
and UO_695 (O_695,N_4858,N_4812);
and UO_696 (O_696,N_4882,N_4816);
or UO_697 (O_697,N_4841,N_4900);
or UO_698 (O_698,N_4880,N_4920);
nor UO_699 (O_699,N_4858,N_4994);
nor UO_700 (O_700,N_4861,N_4805);
xor UO_701 (O_701,N_4860,N_4999);
xor UO_702 (O_702,N_4811,N_4906);
xor UO_703 (O_703,N_4915,N_4875);
nor UO_704 (O_704,N_4880,N_4976);
or UO_705 (O_705,N_4827,N_4922);
nor UO_706 (O_706,N_4853,N_4866);
nand UO_707 (O_707,N_4972,N_4995);
or UO_708 (O_708,N_4975,N_4840);
xor UO_709 (O_709,N_4985,N_4855);
xor UO_710 (O_710,N_4994,N_4976);
and UO_711 (O_711,N_4882,N_4877);
and UO_712 (O_712,N_4959,N_4867);
nand UO_713 (O_713,N_4867,N_4989);
or UO_714 (O_714,N_4990,N_4964);
nor UO_715 (O_715,N_4901,N_4893);
nand UO_716 (O_716,N_4820,N_4887);
nand UO_717 (O_717,N_4860,N_4877);
nand UO_718 (O_718,N_4817,N_4903);
xnor UO_719 (O_719,N_4850,N_4873);
and UO_720 (O_720,N_4940,N_4983);
nor UO_721 (O_721,N_4959,N_4841);
or UO_722 (O_722,N_4880,N_4821);
or UO_723 (O_723,N_4963,N_4857);
nand UO_724 (O_724,N_4820,N_4971);
xor UO_725 (O_725,N_4951,N_4894);
nor UO_726 (O_726,N_4886,N_4847);
nor UO_727 (O_727,N_4918,N_4952);
and UO_728 (O_728,N_4928,N_4954);
and UO_729 (O_729,N_4941,N_4808);
nor UO_730 (O_730,N_4827,N_4803);
nor UO_731 (O_731,N_4955,N_4924);
xnor UO_732 (O_732,N_4957,N_4976);
nor UO_733 (O_733,N_4819,N_4864);
and UO_734 (O_734,N_4987,N_4935);
or UO_735 (O_735,N_4849,N_4884);
nor UO_736 (O_736,N_4892,N_4844);
xor UO_737 (O_737,N_4879,N_4914);
nand UO_738 (O_738,N_4952,N_4814);
nand UO_739 (O_739,N_4882,N_4991);
nand UO_740 (O_740,N_4808,N_4801);
nand UO_741 (O_741,N_4824,N_4899);
nor UO_742 (O_742,N_4902,N_4939);
or UO_743 (O_743,N_4972,N_4969);
nand UO_744 (O_744,N_4987,N_4838);
xnor UO_745 (O_745,N_4832,N_4844);
nor UO_746 (O_746,N_4801,N_4832);
and UO_747 (O_747,N_4829,N_4954);
or UO_748 (O_748,N_4912,N_4836);
and UO_749 (O_749,N_4872,N_4909);
or UO_750 (O_750,N_4836,N_4954);
or UO_751 (O_751,N_4930,N_4902);
nand UO_752 (O_752,N_4951,N_4994);
or UO_753 (O_753,N_4942,N_4863);
and UO_754 (O_754,N_4825,N_4919);
xnor UO_755 (O_755,N_4950,N_4975);
and UO_756 (O_756,N_4824,N_4948);
nand UO_757 (O_757,N_4948,N_4839);
nand UO_758 (O_758,N_4851,N_4813);
nor UO_759 (O_759,N_4802,N_4975);
nand UO_760 (O_760,N_4824,N_4952);
and UO_761 (O_761,N_4958,N_4930);
or UO_762 (O_762,N_4836,N_4870);
and UO_763 (O_763,N_4821,N_4881);
or UO_764 (O_764,N_4920,N_4914);
or UO_765 (O_765,N_4959,N_4901);
xor UO_766 (O_766,N_4957,N_4835);
or UO_767 (O_767,N_4836,N_4857);
xnor UO_768 (O_768,N_4952,N_4934);
xor UO_769 (O_769,N_4828,N_4950);
or UO_770 (O_770,N_4916,N_4861);
nand UO_771 (O_771,N_4840,N_4900);
or UO_772 (O_772,N_4837,N_4908);
and UO_773 (O_773,N_4852,N_4841);
nor UO_774 (O_774,N_4871,N_4936);
and UO_775 (O_775,N_4887,N_4970);
nand UO_776 (O_776,N_4904,N_4942);
or UO_777 (O_777,N_4978,N_4901);
and UO_778 (O_778,N_4965,N_4902);
nor UO_779 (O_779,N_4898,N_4926);
nand UO_780 (O_780,N_4927,N_4962);
or UO_781 (O_781,N_4851,N_4956);
and UO_782 (O_782,N_4996,N_4924);
and UO_783 (O_783,N_4843,N_4844);
xnor UO_784 (O_784,N_4979,N_4969);
nand UO_785 (O_785,N_4873,N_4926);
or UO_786 (O_786,N_4892,N_4893);
or UO_787 (O_787,N_4837,N_4957);
xor UO_788 (O_788,N_4882,N_4944);
nand UO_789 (O_789,N_4919,N_4883);
nor UO_790 (O_790,N_4941,N_4909);
nor UO_791 (O_791,N_4959,N_4803);
xor UO_792 (O_792,N_4976,N_4885);
nor UO_793 (O_793,N_4935,N_4902);
nand UO_794 (O_794,N_4912,N_4950);
nand UO_795 (O_795,N_4999,N_4977);
nand UO_796 (O_796,N_4999,N_4817);
or UO_797 (O_797,N_4920,N_4945);
nor UO_798 (O_798,N_4869,N_4896);
nand UO_799 (O_799,N_4941,N_4985);
nand UO_800 (O_800,N_4889,N_4817);
nor UO_801 (O_801,N_4899,N_4957);
or UO_802 (O_802,N_4932,N_4941);
and UO_803 (O_803,N_4846,N_4995);
nand UO_804 (O_804,N_4902,N_4982);
or UO_805 (O_805,N_4915,N_4974);
nor UO_806 (O_806,N_4901,N_4962);
or UO_807 (O_807,N_4990,N_4884);
or UO_808 (O_808,N_4960,N_4813);
or UO_809 (O_809,N_4823,N_4853);
or UO_810 (O_810,N_4823,N_4969);
or UO_811 (O_811,N_4897,N_4981);
xnor UO_812 (O_812,N_4894,N_4814);
or UO_813 (O_813,N_4906,N_4973);
or UO_814 (O_814,N_4806,N_4972);
and UO_815 (O_815,N_4886,N_4810);
and UO_816 (O_816,N_4971,N_4926);
nand UO_817 (O_817,N_4941,N_4805);
nand UO_818 (O_818,N_4995,N_4875);
or UO_819 (O_819,N_4988,N_4816);
or UO_820 (O_820,N_4945,N_4917);
nor UO_821 (O_821,N_4938,N_4879);
or UO_822 (O_822,N_4812,N_4965);
nor UO_823 (O_823,N_4825,N_4882);
and UO_824 (O_824,N_4967,N_4800);
xor UO_825 (O_825,N_4889,N_4862);
nand UO_826 (O_826,N_4869,N_4944);
nand UO_827 (O_827,N_4963,N_4885);
nor UO_828 (O_828,N_4811,N_4985);
or UO_829 (O_829,N_4897,N_4803);
nand UO_830 (O_830,N_4895,N_4990);
and UO_831 (O_831,N_4990,N_4977);
and UO_832 (O_832,N_4871,N_4909);
nor UO_833 (O_833,N_4814,N_4914);
nor UO_834 (O_834,N_4806,N_4998);
nand UO_835 (O_835,N_4830,N_4924);
nor UO_836 (O_836,N_4984,N_4854);
nand UO_837 (O_837,N_4829,N_4965);
and UO_838 (O_838,N_4825,N_4970);
and UO_839 (O_839,N_4884,N_4909);
xor UO_840 (O_840,N_4815,N_4997);
nor UO_841 (O_841,N_4827,N_4861);
nor UO_842 (O_842,N_4982,N_4866);
xor UO_843 (O_843,N_4849,N_4863);
xor UO_844 (O_844,N_4956,N_4858);
nand UO_845 (O_845,N_4821,N_4984);
nor UO_846 (O_846,N_4828,N_4922);
and UO_847 (O_847,N_4826,N_4850);
or UO_848 (O_848,N_4827,N_4995);
nor UO_849 (O_849,N_4952,N_4912);
or UO_850 (O_850,N_4913,N_4986);
nand UO_851 (O_851,N_4803,N_4868);
nand UO_852 (O_852,N_4869,N_4847);
or UO_853 (O_853,N_4968,N_4827);
xnor UO_854 (O_854,N_4922,N_4901);
xor UO_855 (O_855,N_4989,N_4802);
nor UO_856 (O_856,N_4976,N_4816);
nor UO_857 (O_857,N_4908,N_4864);
nand UO_858 (O_858,N_4803,N_4974);
or UO_859 (O_859,N_4833,N_4843);
or UO_860 (O_860,N_4893,N_4997);
nand UO_861 (O_861,N_4939,N_4836);
xnor UO_862 (O_862,N_4851,N_4861);
and UO_863 (O_863,N_4886,N_4991);
nor UO_864 (O_864,N_4847,N_4824);
nand UO_865 (O_865,N_4880,N_4893);
xnor UO_866 (O_866,N_4941,N_4815);
and UO_867 (O_867,N_4951,N_4901);
nand UO_868 (O_868,N_4987,N_4970);
xnor UO_869 (O_869,N_4866,N_4998);
and UO_870 (O_870,N_4998,N_4921);
xor UO_871 (O_871,N_4912,N_4878);
nor UO_872 (O_872,N_4800,N_4903);
or UO_873 (O_873,N_4873,N_4894);
and UO_874 (O_874,N_4923,N_4946);
xor UO_875 (O_875,N_4801,N_4845);
nor UO_876 (O_876,N_4949,N_4864);
or UO_877 (O_877,N_4853,N_4957);
nand UO_878 (O_878,N_4951,N_4864);
nand UO_879 (O_879,N_4864,N_4904);
and UO_880 (O_880,N_4833,N_4850);
nor UO_881 (O_881,N_4912,N_4991);
nand UO_882 (O_882,N_4837,N_4821);
nor UO_883 (O_883,N_4830,N_4853);
nand UO_884 (O_884,N_4893,N_4993);
or UO_885 (O_885,N_4856,N_4844);
nor UO_886 (O_886,N_4936,N_4814);
nor UO_887 (O_887,N_4954,N_4948);
xor UO_888 (O_888,N_4921,N_4963);
and UO_889 (O_889,N_4917,N_4833);
nand UO_890 (O_890,N_4880,N_4866);
or UO_891 (O_891,N_4948,N_4987);
nand UO_892 (O_892,N_4838,N_4970);
xor UO_893 (O_893,N_4843,N_4909);
and UO_894 (O_894,N_4957,N_4983);
nand UO_895 (O_895,N_4882,N_4900);
nor UO_896 (O_896,N_4926,N_4805);
or UO_897 (O_897,N_4952,N_4811);
and UO_898 (O_898,N_4880,N_4942);
nand UO_899 (O_899,N_4889,N_4995);
and UO_900 (O_900,N_4960,N_4919);
xor UO_901 (O_901,N_4931,N_4912);
or UO_902 (O_902,N_4993,N_4888);
and UO_903 (O_903,N_4881,N_4872);
nor UO_904 (O_904,N_4956,N_4885);
and UO_905 (O_905,N_4974,N_4914);
nor UO_906 (O_906,N_4925,N_4838);
nor UO_907 (O_907,N_4913,N_4832);
nand UO_908 (O_908,N_4997,N_4818);
xnor UO_909 (O_909,N_4951,N_4862);
or UO_910 (O_910,N_4862,N_4967);
nor UO_911 (O_911,N_4833,N_4972);
xnor UO_912 (O_912,N_4826,N_4961);
nor UO_913 (O_913,N_4919,N_4815);
xor UO_914 (O_914,N_4890,N_4974);
xnor UO_915 (O_915,N_4866,N_4819);
xor UO_916 (O_916,N_4972,N_4892);
and UO_917 (O_917,N_4883,N_4946);
xor UO_918 (O_918,N_4864,N_4980);
nor UO_919 (O_919,N_4944,N_4918);
nand UO_920 (O_920,N_4893,N_4875);
and UO_921 (O_921,N_4948,N_4996);
nor UO_922 (O_922,N_4856,N_4918);
nor UO_923 (O_923,N_4954,N_4851);
or UO_924 (O_924,N_4806,N_4907);
nand UO_925 (O_925,N_4833,N_4907);
nor UO_926 (O_926,N_4855,N_4902);
nand UO_927 (O_927,N_4978,N_4834);
xnor UO_928 (O_928,N_4806,N_4925);
xnor UO_929 (O_929,N_4969,N_4911);
xnor UO_930 (O_930,N_4803,N_4819);
and UO_931 (O_931,N_4997,N_4980);
xnor UO_932 (O_932,N_4871,N_4826);
nand UO_933 (O_933,N_4895,N_4963);
xor UO_934 (O_934,N_4975,N_4884);
nand UO_935 (O_935,N_4837,N_4916);
nor UO_936 (O_936,N_4811,N_4962);
xnor UO_937 (O_937,N_4929,N_4910);
nor UO_938 (O_938,N_4990,N_4942);
nor UO_939 (O_939,N_4838,N_4817);
and UO_940 (O_940,N_4908,N_4960);
or UO_941 (O_941,N_4823,N_4977);
and UO_942 (O_942,N_4990,N_4981);
nor UO_943 (O_943,N_4929,N_4887);
xnor UO_944 (O_944,N_4944,N_4926);
nor UO_945 (O_945,N_4970,N_4940);
nand UO_946 (O_946,N_4852,N_4956);
xnor UO_947 (O_947,N_4896,N_4816);
and UO_948 (O_948,N_4911,N_4960);
or UO_949 (O_949,N_4841,N_4878);
and UO_950 (O_950,N_4987,N_4958);
nor UO_951 (O_951,N_4988,N_4960);
xor UO_952 (O_952,N_4849,N_4925);
nor UO_953 (O_953,N_4914,N_4818);
nor UO_954 (O_954,N_4898,N_4805);
nor UO_955 (O_955,N_4917,N_4882);
nor UO_956 (O_956,N_4810,N_4994);
and UO_957 (O_957,N_4932,N_4806);
and UO_958 (O_958,N_4893,N_4924);
nor UO_959 (O_959,N_4821,N_4951);
xnor UO_960 (O_960,N_4807,N_4857);
nor UO_961 (O_961,N_4929,N_4846);
and UO_962 (O_962,N_4919,N_4956);
and UO_963 (O_963,N_4886,N_4877);
nor UO_964 (O_964,N_4986,N_4872);
and UO_965 (O_965,N_4881,N_4930);
nor UO_966 (O_966,N_4993,N_4995);
xor UO_967 (O_967,N_4853,N_4930);
and UO_968 (O_968,N_4816,N_4873);
xnor UO_969 (O_969,N_4820,N_4884);
nand UO_970 (O_970,N_4842,N_4854);
and UO_971 (O_971,N_4851,N_4841);
xor UO_972 (O_972,N_4951,N_4805);
xnor UO_973 (O_973,N_4842,N_4866);
nand UO_974 (O_974,N_4825,N_4923);
nand UO_975 (O_975,N_4898,N_4997);
and UO_976 (O_976,N_4939,N_4867);
nand UO_977 (O_977,N_4843,N_4827);
nand UO_978 (O_978,N_4881,N_4829);
xnor UO_979 (O_979,N_4853,N_4916);
nand UO_980 (O_980,N_4826,N_4931);
xor UO_981 (O_981,N_4926,N_4955);
or UO_982 (O_982,N_4937,N_4865);
nor UO_983 (O_983,N_4925,N_4965);
and UO_984 (O_984,N_4932,N_4926);
and UO_985 (O_985,N_4937,N_4967);
and UO_986 (O_986,N_4863,N_4974);
and UO_987 (O_987,N_4967,N_4955);
and UO_988 (O_988,N_4951,N_4967);
and UO_989 (O_989,N_4805,N_4816);
xor UO_990 (O_990,N_4997,N_4905);
or UO_991 (O_991,N_4985,N_4903);
nor UO_992 (O_992,N_4870,N_4959);
or UO_993 (O_993,N_4806,N_4816);
nand UO_994 (O_994,N_4944,N_4897);
or UO_995 (O_995,N_4945,N_4892);
nand UO_996 (O_996,N_4970,N_4999);
and UO_997 (O_997,N_4940,N_4912);
nand UO_998 (O_998,N_4968,N_4938);
nand UO_999 (O_999,N_4911,N_4866);
endmodule