module basic_3000_30000_3500_30_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1481,In_264);
nand U1 (N_1,In_1993,In_2428);
nor U2 (N_2,In_498,In_2073);
nor U3 (N_3,In_2356,In_2062);
nor U4 (N_4,In_2063,In_531);
xnor U5 (N_5,In_1748,In_2900);
xnor U6 (N_6,In_1423,In_823);
nand U7 (N_7,In_817,In_2658);
nor U8 (N_8,In_1773,In_494);
nand U9 (N_9,In_1323,In_759);
nor U10 (N_10,In_622,In_1177);
nor U11 (N_11,In_1170,In_2313);
xor U12 (N_12,In_2746,In_939);
and U13 (N_13,In_411,In_1353);
nand U14 (N_14,In_268,In_1247);
nand U15 (N_15,In_1977,In_2638);
or U16 (N_16,In_2924,In_1191);
nand U17 (N_17,In_2701,In_2446);
xor U18 (N_18,In_1223,In_2174);
and U19 (N_19,In_157,In_1349);
and U20 (N_20,In_2140,In_550);
xor U21 (N_21,In_1290,In_1689);
xor U22 (N_22,In_2159,In_2411);
xor U23 (N_23,In_953,In_1712);
nand U24 (N_24,In_1233,In_260);
and U25 (N_25,In_994,In_2917);
nand U26 (N_26,In_565,In_2022);
nor U27 (N_27,In_1669,In_974);
nand U28 (N_28,In_1457,In_1617);
nand U29 (N_29,In_446,In_1976);
nor U30 (N_30,In_927,In_168);
xnor U31 (N_31,In_1996,In_1698);
or U32 (N_32,In_1044,In_1259);
and U33 (N_33,In_2755,In_1809);
and U34 (N_34,In_102,In_1483);
or U35 (N_35,In_595,In_77);
nor U36 (N_36,In_2271,In_990);
nor U37 (N_37,In_434,In_2191);
and U38 (N_38,In_2883,In_2728);
or U39 (N_39,In_1274,In_1393);
nor U40 (N_40,In_2896,In_2686);
xor U41 (N_41,In_2552,In_75);
and U42 (N_42,In_1872,In_1547);
xor U43 (N_43,In_1798,In_147);
or U44 (N_44,In_697,In_204);
xor U45 (N_45,In_2311,In_1186);
nand U46 (N_46,In_860,In_2644);
nand U47 (N_47,In_1578,In_2669);
xor U48 (N_48,In_2793,In_786);
and U49 (N_49,In_2057,In_2088);
nor U50 (N_50,In_1100,In_1509);
or U51 (N_51,In_1720,In_2152);
xor U52 (N_52,In_611,In_1376);
xor U53 (N_53,In_2745,In_1168);
nor U54 (N_54,In_2231,In_2808);
and U55 (N_55,In_629,In_1126);
nand U56 (N_56,In_92,In_2371);
or U57 (N_57,In_1466,In_153);
and U58 (N_58,In_2656,In_1709);
nand U59 (N_59,In_230,In_19);
or U60 (N_60,In_2027,In_547);
nor U61 (N_61,In_2420,In_671);
xnor U62 (N_62,In_49,In_2744);
nor U63 (N_63,In_1018,In_1447);
nor U64 (N_64,In_435,In_617);
and U65 (N_65,In_1943,In_445);
nor U66 (N_66,In_1987,In_978);
nand U67 (N_67,In_1127,In_185);
nand U68 (N_68,In_1485,In_1317);
and U69 (N_69,In_2981,In_2256);
or U70 (N_70,In_1704,In_453);
and U71 (N_71,In_2662,In_1360);
or U72 (N_72,In_1192,In_1900);
nor U73 (N_73,In_683,In_2984);
nand U74 (N_74,In_1634,In_2943);
xor U75 (N_75,In_1021,In_2992);
nor U76 (N_76,In_2399,In_416);
nand U77 (N_77,In_2978,In_288);
or U78 (N_78,In_1421,In_1874);
xor U79 (N_79,In_1143,In_1591);
xnor U80 (N_80,In_55,In_1020);
and U81 (N_81,In_928,In_1877);
and U82 (N_82,In_1907,In_1867);
xnor U83 (N_83,In_2930,In_703);
and U84 (N_84,In_1273,In_359);
and U85 (N_85,In_1929,In_947);
nor U86 (N_86,In_428,In_81);
xnor U87 (N_87,In_2634,In_1472);
and U88 (N_88,In_930,In_2763);
xor U89 (N_89,In_919,In_2532);
and U90 (N_90,In_2330,In_2121);
and U91 (N_91,In_2483,In_2011);
or U92 (N_92,In_734,In_1388);
and U93 (N_93,In_2690,In_1230);
nand U94 (N_94,In_2869,In_174);
nand U95 (N_95,In_2214,In_2989);
nor U96 (N_96,In_457,In_2895);
nand U97 (N_97,In_1546,In_122);
xor U98 (N_98,In_871,In_2245);
nand U99 (N_99,In_320,In_2509);
or U100 (N_100,In_551,In_235);
or U101 (N_101,In_339,In_1201);
nor U102 (N_102,In_383,In_32);
nand U103 (N_103,In_1014,In_117);
xor U104 (N_104,In_2787,In_2444);
nor U105 (N_105,In_1846,In_738);
or U106 (N_106,In_1831,In_2406);
nand U107 (N_107,In_1415,In_948);
or U108 (N_108,In_1735,In_2849);
and U109 (N_109,In_845,In_1304);
xor U110 (N_110,In_2613,In_1626);
xor U111 (N_111,In_1113,In_1582);
or U112 (N_112,In_1162,In_266);
or U113 (N_113,In_2370,In_2248);
nand U114 (N_114,In_1428,In_2844);
or U115 (N_115,In_941,In_2113);
nor U116 (N_116,In_1569,In_818);
or U117 (N_117,In_1622,In_2529);
xnor U118 (N_118,In_376,In_1010);
and U119 (N_119,In_917,In_1275);
or U120 (N_120,In_283,In_1329);
xnor U121 (N_121,In_1053,In_1718);
nand U122 (N_122,In_90,In_2516);
nor U123 (N_123,In_2819,In_783);
nor U124 (N_124,In_1465,In_2608);
nor U125 (N_125,In_1612,In_1486);
nor U126 (N_126,In_760,In_1656);
and U127 (N_127,In_1158,In_1737);
nand U128 (N_128,In_854,In_1971);
or U129 (N_129,In_2855,In_280);
and U130 (N_130,In_72,In_542);
xnor U131 (N_131,In_2203,In_605);
xor U132 (N_132,In_1086,In_2751);
nand U133 (N_133,In_1570,In_1592);
nor U134 (N_134,In_1864,In_2747);
xor U135 (N_135,In_1330,In_2202);
nand U136 (N_136,In_1912,In_321);
xor U137 (N_137,In_2782,In_1901);
and U138 (N_138,In_1286,In_2725);
nand U139 (N_139,In_2825,In_2103);
or U140 (N_140,In_1318,In_2069);
nor U141 (N_141,In_596,In_532);
nor U142 (N_142,In_1299,In_1052);
and U143 (N_143,In_2035,In_1713);
or U144 (N_144,In_368,In_2920);
nor U145 (N_145,In_223,In_731);
nand U146 (N_146,In_2902,In_1117);
xor U147 (N_147,In_2734,In_1830);
or U148 (N_148,In_1670,In_1104);
nand U149 (N_149,In_2230,In_313);
nor U150 (N_150,In_1433,In_552);
xnor U151 (N_151,In_166,In_2589);
and U152 (N_152,In_281,In_2340);
nand U153 (N_153,In_2070,In_2165);
xnor U154 (N_154,In_2997,In_556);
or U155 (N_155,In_2864,In_1611);
and U156 (N_156,In_2814,In_897);
xor U157 (N_157,In_342,In_2228);
nand U158 (N_158,In_152,In_2031);
xor U159 (N_159,In_2386,In_2729);
nor U160 (N_160,In_332,In_802);
and U161 (N_161,In_1309,In_1429);
or U162 (N_162,In_2923,In_298);
nand U163 (N_163,In_2307,In_1639);
nand U164 (N_164,In_1489,In_1512);
or U165 (N_165,In_2440,In_619);
or U166 (N_166,In_140,In_1694);
nand U167 (N_167,In_796,In_2049);
nor U168 (N_168,In_30,In_1125);
nand U169 (N_169,In_2253,In_849);
xnor U170 (N_170,In_2522,In_2128);
xnor U171 (N_171,In_1710,In_2741);
nand U172 (N_172,In_2267,In_2938);
xnor U173 (N_173,In_2560,In_2919);
or U174 (N_174,In_1974,In_123);
nand U175 (N_175,In_1576,In_2710);
nand U176 (N_176,In_1716,In_1940);
xnor U177 (N_177,In_139,In_704);
xnor U178 (N_178,In_2309,In_1862);
nand U179 (N_179,In_1244,In_643);
nor U180 (N_180,In_634,In_2602);
and U181 (N_181,In_1387,In_1848);
or U182 (N_182,In_415,In_2162);
nand U183 (N_183,In_1280,In_2562);
or U184 (N_184,In_878,In_1377);
xor U185 (N_185,In_2637,In_2357);
or U186 (N_186,In_913,In_1695);
nand U187 (N_187,In_1559,In_966);
or U188 (N_188,In_2952,In_150);
xor U189 (N_189,In_1400,In_2795);
nor U190 (N_190,In_1654,In_2722);
or U191 (N_191,In_540,In_142);
nor U192 (N_192,In_1498,In_912);
nand U193 (N_193,In_2675,In_2236);
or U194 (N_194,In_1785,In_156);
and U195 (N_195,In_2880,In_2287);
or U196 (N_196,In_748,In_2369);
or U197 (N_197,In_1897,In_1727);
or U198 (N_198,In_1346,In_539);
xnor U199 (N_199,In_1607,In_1517);
or U200 (N_200,In_2665,In_581);
or U201 (N_201,In_1205,In_2769);
xor U202 (N_202,In_792,In_664);
nor U203 (N_203,In_2495,In_1787);
xnor U204 (N_204,In_421,In_1527);
nand U205 (N_205,In_2834,In_1101);
or U206 (N_206,In_1175,In_2947);
or U207 (N_207,In_2812,In_2192);
or U208 (N_208,In_85,In_1240);
xor U209 (N_209,In_2342,In_2991);
nor U210 (N_210,In_2204,In_2946);
nor U211 (N_211,In_1955,In_2142);
xnor U212 (N_212,In_2577,In_1478);
nor U213 (N_213,In_2008,In_2545);
or U214 (N_214,In_839,In_371);
nor U215 (N_215,In_1746,In_2845);
xor U216 (N_216,In_1542,In_1772);
xnor U217 (N_217,In_2618,In_1045);
and U218 (N_218,In_2242,In_2884);
xnor U219 (N_219,In_2506,In_1573);
and U220 (N_220,In_128,In_1790);
or U221 (N_221,In_2765,In_699);
or U222 (N_222,In_2828,In_2655);
xor U223 (N_223,In_1236,In_754);
and U224 (N_224,In_663,In_2372);
or U225 (N_225,In_1535,In_1167);
and U226 (N_226,In_379,In_1159);
nor U227 (N_227,In_2972,In_613);
or U228 (N_228,In_2350,In_2133);
and U229 (N_229,In_2630,In_847);
xor U230 (N_230,In_1339,In_2859);
nand U231 (N_231,In_625,In_536);
nor U232 (N_232,In_258,In_2810);
nor U233 (N_233,In_1118,In_237);
nor U234 (N_234,In_2705,In_1320);
or U235 (N_235,In_1895,In_1190);
nand U236 (N_236,In_440,In_2161);
nand U237 (N_237,In_2857,In_56);
nor U238 (N_238,In_1111,In_2543);
xor U239 (N_239,In_2061,In_1051);
nand U240 (N_240,In_1555,In_2820);
or U241 (N_241,In_696,In_68);
and U242 (N_242,In_2328,In_915);
nor U243 (N_243,In_1928,In_2282);
nor U244 (N_244,In_2612,In_1814);
nand U245 (N_245,In_389,In_631);
nor U246 (N_246,In_2974,In_820);
nor U247 (N_247,In_1313,In_2831);
nand U248 (N_248,In_574,In_480);
nor U249 (N_249,In_1794,In_831);
nand U250 (N_250,In_702,In_322);
or U251 (N_251,In_187,In_658);
or U252 (N_252,In_2870,In_183);
nand U253 (N_253,In_2575,In_2911);
or U254 (N_254,In_370,In_609);
or U255 (N_255,In_1887,In_1919);
nor U256 (N_256,In_296,In_220);
nor U257 (N_257,In_1635,In_2051);
nand U258 (N_258,In_2776,In_1705);
xor U259 (N_259,In_1147,In_2479);
nor U260 (N_260,In_1030,In_1650);
or U261 (N_261,In_357,In_2540);
or U262 (N_262,In_1595,In_1381);
or U263 (N_263,In_483,In_1185);
nor U264 (N_264,In_2866,In_893);
nand U265 (N_265,In_148,In_1491);
xor U266 (N_266,In_1050,In_2709);
xor U267 (N_267,In_2183,In_2316);
or U268 (N_268,In_2156,In_2100);
and U269 (N_269,In_753,In_2858);
xnor U270 (N_270,In_872,In_891);
xnor U271 (N_271,In_84,In_2962);
or U272 (N_272,In_2447,In_1131);
nand U273 (N_273,In_291,In_1495);
and U274 (N_274,In_2032,In_1193);
or U275 (N_275,In_2374,In_1751);
nor U276 (N_276,In_2742,In_1648);
or U277 (N_277,In_196,In_51);
xnor U278 (N_278,In_916,In_2778);
xor U279 (N_279,In_1740,In_1629);
xnor U280 (N_280,In_1777,In_215);
nor U281 (N_281,In_2549,In_361);
nor U282 (N_282,In_2368,In_182);
or U283 (N_283,In_401,In_894);
nor U284 (N_284,In_1386,In_1276);
nand U285 (N_285,In_95,In_713);
and U286 (N_286,In_1107,In_1249);
or U287 (N_287,In_1951,In_1769);
nand U288 (N_288,In_2721,In_2237);
xor U289 (N_289,In_2412,In_97);
nor U290 (N_290,In_986,In_508);
or U291 (N_291,In_501,In_2891);
or U292 (N_292,In_1451,In_1029);
and U293 (N_293,In_518,In_1646);
and U294 (N_294,In_2762,In_1587);
and U295 (N_295,In_2581,In_460);
nor U296 (N_296,In_1343,In_2714);
nor U297 (N_297,In_420,In_1268);
nor U298 (N_298,In_1950,In_2334);
nor U299 (N_299,In_2757,In_2800);
nand U300 (N_300,In_770,In_1416);
xor U301 (N_301,In_492,In_206);
and U302 (N_302,In_26,In_2535);
or U303 (N_303,In_1925,In_1293);
nor U304 (N_304,In_2736,In_945);
xor U305 (N_305,In_2918,In_724);
xor U306 (N_306,In_2942,In_1970);
nor U307 (N_307,In_251,In_209);
and U308 (N_308,In_1090,In_57);
and U309 (N_309,In_373,In_1953);
nor U310 (N_310,In_650,In_2590);
and U311 (N_311,In_618,In_2789);
or U312 (N_312,In_2862,In_289);
nor U313 (N_313,In_2053,In_1399);
xor U314 (N_314,In_835,In_2885);
xnor U315 (N_315,In_2886,In_1812);
and U316 (N_316,In_245,In_2117);
and U317 (N_317,In_331,In_982);
or U318 (N_318,In_2670,In_274);
nor U319 (N_319,In_2401,In_319);
or U320 (N_320,In_398,In_1992);
nor U321 (N_321,In_240,In_2302);
and U322 (N_322,In_2487,In_1544);
nor U323 (N_323,In_2127,In_348);
nand U324 (N_324,In_126,In_2004);
nor U325 (N_325,In_995,In_846);
or U326 (N_326,In_1039,In_239);
xnor U327 (N_327,In_2044,In_1915);
and U328 (N_328,In_422,In_2515);
and U329 (N_329,In_1606,In_2771);
xor U330 (N_330,In_2317,In_2259);
xor U331 (N_331,In_692,In_2012);
xor U332 (N_332,In_2286,In_448);
nand U333 (N_333,In_832,In_44);
and U334 (N_334,In_795,In_1696);
or U335 (N_335,In_1528,In_2818);
nor U336 (N_336,In_1514,In_2905);
xnor U337 (N_337,In_2272,In_232);
nor U338 (N_338,In_1764,In_1964);
or U339 (N_339,In_2505,In_2116);
nand U340 (N_340,In_1181,In_1176);
nand U341 (N_341,In_1148,In_808);
nand U342 (N_342,In_450,In_730);
xor U343 (N_343,In_1803,In_1620);
xor U344 (N_344,In_218,In_1009);
or U345 (N_345,In_1644,In_2284);
and U346 (N_346,In_1609,In_113);
nand U347 (N_347,In_1657,In_2914);
xor U348 (N_348,In_1923,In_890);
nand U349 (N_349,In_1766,In_1963);
and U350 (N_350,In_1728,In_1816);
nand U351 (N_351,In_541,In_700);
nand U352 (N_352,In_2455,In_2957);
xor U353 (N_353,In_2743,In_1526);
and U354 (N_354,In_1337,In_249);
nand U355 (N_355,In_2898,In_1700);
and U356 (N_356,In_2007,In_165);
or U357 (N_357,In_2243,In_59);
and U358 (N_358,In_1425,In_1824);
xnor U359 (N_359,In_1732,In_1999);
or U360 (N_360,In_2325,In_366);
nand U361 (N_361,In_2454,In_709);
nor U362 (N_362,In_2564,In_2783);
and U363 (N_363,In_1212,In_391);
or U364 (N_364,In_2018,In_2093);
nand U365 (N_365,In_1532,In_1757);
or U366 (N_366,In_638,In_146);
and U367 (N_367,In_644,In_311);
or U368 (N_368,In_306,In_728);
xnor U369 (N_369,In_1667,In_295);
xor U370 (N_370,In_353,In_1308);
xor U371 (N_371,In_2339,In_2636);
nand U372 (N_372,In_1693,In_277);
nand U373 (N_373,In_1924,In_2711);
and U374 (N_374,In_1361,In_1397);
xnor U375 (N_375,In_10,In_884);
nor U376 (N_376,In_1701,In_549);
nor U377 (N_377,In_645,In_314);
and U378 (N_378,In_468,In_954);
nand U379 (N_379,In_2265,In_1366);
nand U380 (N_380,In_842,In_2352);
xor U381 (N_381,In_1982,In_2042);
and U382 (N_382,In_1434,In_1340);
nor U383 (N_383,In_962,In_1444);
xnor U384 (N_384,In_1161,In_2582);
xnor U385 (N_385,In_1843,In_2065);
nand U386 (N_386,In_431,In_1703);
nor U387 (N_387,In_1155,In_2358);
nand U388 (N_388,In_37,In_855);
or U389 (N_389,In_1019,In_1768);
xor U390 (N_390,In_1197,In_336);
xnor U391 (N_391,In_127,In_2470);
xnor U392 (N_392,In_1204,In_1692);
xnor U393 (N_393,In_74,In_2171);
nor U394 (N_394,In_1891,In_270);
or U395 (N_395,In_1404,In_144);
nand U396 (N_396,In_1658,In_648);
and U397 (N_397,In_488,In_2348);
nand U398 (N_398,In_725,In_2347);
and U399 (N_399,In_1754,In_2468);
xnor U400 (N_400,In_224,In_761);
xnor U401 (N_401,In_2474,In_2803);
nor U402 (N_402,In_621,In_1112);
nor U403 (N_403,In_307,In_2132);
or U404 (N_404,In_2547,In_63);
or U405 (N_405,In_259,In_2226);
xor U406 (N_406,In_0,In_749);
and U407 (N_407,In_506,In_426);
or U408 (N_408,In_620,In_17);
xnor U409 (N_409,In_364,In_2615);
nor U410 (N_410,In_2092,In_1157);
nand U411 (N_411,In_2623,In_1407);
xor U412 (N_412,In_1847,In_2212);
nand U413 (N_413,In_1518,In_2723);
nand U414 (N_414,In_1672,In_1771);
and U415 (N_415,In_2335,In_1707);
xor U416 (N_416,In_1149,In_413);
nand U417 (N_417,In_1123,In_1080);
xor U418 (N_418,In_1091,In_2198);
nand U419 (N_419,In_2996,In_1257);
nor U420 (N_420,In_184,In_2625);
xnor U421 (N_421,In_2944,In_1972);
or U422 (N_422,In_456,In_124);
nor U423 (N_423,In_1326,In_2512);
or U424 (N_424,In_1110,In_2046);
nor U425 (N_425,In_1464,In_1202);
xor U426 (N_426,In_2036,In_2843);
and U427 (N_427,In_1427,In_938);
xnor U428 (N_428,In_993,In_815);
nand U429 (N_429,In_2852,In_2966);
xnor U430 (N_430,In_2708,In_1579);
nor U431 (N_431,In_2960,In_372);
xor U432 (N_432,In_1808,In_2402);
and U433 (N_433,In_112,In_2407);
xor U434 (N_434,In_825,In_2616);
xor U435 (N_435,In_1668,In_1165);
xor U436 (N_436,In_137,In_992);
or U437 (N_437,In_1437,In_61);
xnor U438 (N_438,In_104,In_951);
xnor U439 (N_439,In_757,In_1796);
nand U440 (N_440,In_880,In_2520);
xor U441 (N_441,In_1375,In_1122);
xnor U442 (N_442,In_665,In_2856);
nand U443 (N_443,In_2089,In_2097);
xor U444 (N_444,In_1163,In_2481);
and U445 (N_445,In_1742,In_1885);
xnor U446 (N_446,In_686,In_191);
or U447 (N_447,In_1279,In_1580);
xor U448 (N_448,In_86,In_2014);
nand U449 (N_449,In_1784,In_2200);
xnor U450 (N_450,In_1730,In_46);
and U451 (N_451,In_1917,In_2893);
and U452 (N_452,In_533,In_933);
xnor U453 (N_453,In_1139,In_1908);
xor U454 (N_454,In_582,In_538);
nor U455 (N_455,In_1477,In_1586);
nor U456 (N_456,In_1537,In_2244);
and U457 (N_457,In_2377,In_50);
or U458 (N_458,In_308,In_1775);
nor U459 (N_459,In_2109,In_315);
nand U460 (N_460,In_449,In_2169);
nand U461 (N_461,In_2383,In_1027);
xnor U462 (N_462,In_226,In_1032);
nand U463 (N_463,In_1820,In_1246);
xnor U464 (N_464,In_2426,In_2164);
or U465 (N_465,In_1140,In_466);
nand U466 (N_466,In_1173,In_2082);
and U467 (N_467,In_1833,In_1556);
nor U468 (N_468,In_745,In_1844);
nand U469 (N_469,In_1443,In_2262);
nor U470 (N_470,In_769,In_1322);
and U471 (N_471,In_1837,In_2851);
or U472 (N_472,In_1467,In_1819);
nand U473 (N_473,In_1235,In_2683);
nand U474 (N_474,In_405,In_2737);
nor U475 (N_475,In_553,In_544);
or U476 (N_476,In_2542,In_423);
nand U477 (N_477,In_15,In_682);
nor U478 (N_478,In_175,In_2201);
or U479 (N_479,In_908,In_1958);
nor U480 (N_480,In_1084,In_830);
or U481 (N_481,In_2318,In_2621);
or U482 (N_482,In_2712,In_2748);
or U483 (N_483,In_1055,In_859);
nor U484 (N_484,In_1673,In_558);
nor U485 (N_485,In_2176,In_1327);
xnor U486 (N_486,In_2892,In_1179);
or U487 (N_487,In_2830,In_469);
nor U488 (N_488,In_1463,In_1662);
and U489 (N_489,In_586,In_2592);
and U490 (N_490,In_1767,In_1380);
or U491 (N_491,In_130,In_784);
nor U492 (N_492,In_726,In_2847);
nor U493 (N_493,In_2939,In_657);
and U494 (N_494,In_1926,In_2416);
nor U495 (N_495,In_684,In_2601);
xnor U496 (N_496,In_1553,In_2873);
nand U497 (N_497,In_2780,In_1141);
and U498 (N_498,In_2538,In_1681);
xor U499 (N_499,In_2593,In_2055);
and U500 (N_500,In_1288,In_2405);
nor U501 (N_501,In_656,In_2530);
or U502 (N_502,In_427,In_1749);
nor U503 (N_503,In_1406,In_2039);
nand U504 (N_504,In_2308,In_996);
xnor U505 (N_505,In_2700,In_2788);
xnor U506 (N_506,In_1097,In_2563);
xnor U507 (N_507,In_895,In_1362);
nor U508 (N_508,In_868,In_2422);
xor U509 (N_509,In_47,In_2707);
nor U510 (N_510,In_62,In_2689);
nor U511 (N_511,In_212,In_1541);
nor U512 (N_512,In_2457,In_1956);
or U513 (N_513,In_2072,In_2460);
xor U514 (N_514,In_1153,In_2807);
nor U515 (N_515,In_837,In_2727);
xor U516 (N_516,In_1813,In_766);
nand U517 (N_517,In_1741,In_484);
and U518 (N_518,In_1253,In_1596);
nand U519 (N_519,In_465,In_2731);
nor U520 (N_520,In_1390,In_563);
nor U521 (N_521,In_1410,In_1988);
and U522 (N_522,In_2754,In_247);
and U523 (N_523,In_101,In_2827);
or U524 (N_524,In_358,In_151);
nand U525 (N_525,In_666,In_341);
nand U526 (N_526,In_1085,In_1726);
or U527 (N_527,In_639,In_675);
nor U528 (N_528,In_513,In_1488);
nand U529 (N_529,In_1272,In_70);
nor U530 (N_530,In_1060,In_2289);
nand U531 (N_531,In_500,In_143);
or U532 (N_532,In_351,In_1401);
nand U533 (N_533,In_2429,In_2817);
and U534 (N_534,In_1385,In_2343);
or U535 (N_535,In_1238,In_177);
nand U536 (N_536,In_1405,In_1560);
and U537 (N_537,In_7,In_385);
nand U538 (N_538,In_2054,In_111);
or U539 (N_539,In_2551,In_2336);
xor U540 (N_540,In_1025,In_2270);
nand U541 (N_541,In_2587,In_2585);
xnor U542 (N_542,In_2663,In_2597);
or U543 (N_543,In_821,In_2076);
xor U544 (N_544,In_2341,In_1931);
or U545 (N_545,In_2629,In_487);
nand U546 (N_546,In_2450,In_2977);
nor U547 (N_547,In_2079,In_922);
xnor U548 (N_548,In_2492,In_780);
nor U549 (N_549,In_2798,In_1878);
nor U550 (N_550,In_1154,In_408);
nand U551 (N_551,In_33,In_1187);
or U552 (N_552,In_876,In_2019);
or U553 (N_553,In_2280,In_2059);
nand U554 (N_554,In_131,In_592);
and U555 (N_555,In_1336,In_2149);
xor U556 (N_556,In_1699,In_316);
nor U557 (N_557,In_2151,In_567);
or U558 (N_558,In_1838,In_2364);
xnor U559 (N_559,In_2120,In_2091);
or U560 (N_560,In_2124,In_355);
and U561 (N_561,In_2222,In_2801);
nand U562 (N_562,In_750,In_1383);
nor U563 (N_563,In_115,In_442);
and U564 (N_564,In_1420,In_1575);
or U565 (N_565,In_1879,In_2002);
and U566 (N_566,In_2217,In_1920);
and U567 (N_567,In_2170,In_673);
nor U568 (N_568,In_526,In_999);
xnor U569 (N_569,In_2137,In_1074);
nor U570 (N_570,In_1857,In_924);
xor U571 (N_571,In_2102,In_198);
or U572 (N_572,In_2067,In_2344);
and U573 (N_573,In_2080,In_346);
nor U574 (N_574,In_1945,In_560);
or U575 (N_575,In_869,In_2840);
nand U576 (N_576,In_1134,In_2986);
nor U577 (N_577,In_546,In_129);
xor U578 (N_578,In_39,In_2375);
and U579 (N_579,In_231,In_944);
and U580 (N_580,In_2408,In_594);
or U581 (N_581,In_1733,In_2600);
nand U582 (N_582,In_463,In_1108);
xnor U583 (N_583,In_1225,In_1598);
xnor U584 (N_584,In_40,In_1414);
and U585 (N_585,In_2699,In_2519);
nand U586 (N_586,In_2373,In_2392);
xor U587 (N_587,In_2674,In_1828);
nor U588 (N_588,In_900,In_1363);
and U589 (N_589,In_1690,In_2464);
xnor U590 (N_590,In_2688,In_1260);
or U591 (N_591,In_257,In_1765);
and U592 (N_592,In_1600,In_2257);
and U593 (N_593,In_2441,In_1218);
xnor U594 (N_594,In_1208,In_414);
nand U595 (N_595,In_2871,In_2667);
or U596 (N_596,In_2013,In_1524);
nand U597 (N_597,In_1358,In_740);
or U598 (N_598,In_199,In_2482);
xnor U599 (N_599,In_1145,In_777);
nor U600 (N_600,In_1169,In_1494);
or U601 (N_601,In_1960,In_425);
or U602 (N_602,In_668,In_1529);
xnor U603 (N_603,In_569,In_1351);
nor U604 (N_604,In_873,In_1446);
xor U605 (N_605,In_503,In_2907);
nor U606 (N_606,In_2521,In_350);
nand U607 (N_607,In_1630,In_829);
nand U608 (N_608,In_719,In_244);
nand U609 (N_609,In_615,In_1378);
and U610 (N_610,In_1655,In_1389);
or U611 (N_611,In_2523,In_2779);
and U612 (N_612,In_222,In_801);
nor U613 (N_613,In_2687,In_2250);
and U614 (N_614,In_2233,In_2649);
xnor U615 (N_615,In_989,In_1432);
nor U616 (N_616,In_1763,In_998);
or U617 (N_617,In_2135,In_470);
nand U618 (N_618,In_2985,In_499);
nand U619 (N_619,In_109,In_952);
nand U620 (N_620,In_2878,In_1935);
xor U621 (N_621,In_2258,In_2901);
nand U622 (N_622,In_2921,In_360);
and U623 (N_623,In_1708,In_1674);
and U624 (N_624,In_1585,In_1312);
nand U625 (N_625,In_2025,In_1990);
xnor U626 (N_626,In_1136,In_301);
nand U627 (N_627,In_767,In_712);
or U628 (N_628,In_141,In_1368);
nand U629 (N_629,In_2887,In_1557);
nand U630 (N_630,In_386,In_852);
xnor U631 (N_631,In_490,In_2430);
nor U632 (N_632,In_1316,In_827);
nand U633 (N_633,In_747,In_20);
xnor U634 (N_634,In_680,In_811);
or U635 (N_635,In_2136,In_2584);
nand U636 (N_636,In_18,In_1936);
or U637 (N_637,In_2567,In_2016);
and U638 (N_638,In_814,In_1997);
nand U639 (N_639,In_1978,In_773);
or U640 (N_640,In_1228,In_263);
xor U641 (N_641,In_297,In_937);
and U642 (N_642,In_2556,In_1590);
nor U643 (N_643,In_179,In_2195);
xnor U644 (N_644,In_545,In_1254);
nor U645 (N_645,In_1264,In_80);
nand U646 (N_646,In_1503,In_2982);
nor U647 (N_647,In_2832,In_2620);
nor U648 (N_648,In_936,In_2648);
and U649 (N_649,In_2614,In_2398);
and U650 (N_650,In_762,In_2153);
and U651 (N_651,In_520,In_2635);
nor U652 (N_652,In_1120,In_534);
and U653 (N_653,In_1015,In_1632);
xnor U654 (N_654,In_1115,In_1295);
nand U655 (N_655,In_1893,In_653);
nand U656 (N_656,In_340,In_2726);
and U657 (N_657,In_197,In_660);
and U658 (N_658,In_1636,In_1067);
xor U659 (N_659,In_2837,In_1851);
or U660 (N_660,In_1865,In_1142);
nand U661 (N_661,In_926,In_1680);
nor U662 (N_662,In_509,In_778);
nor U663 (N_663,In_2172,In_746);
nand U664 (N_664,In_2525,In_94);
xnor U665 (N_665,In_688,In_1203);
or U666 (N_666,In_1475,In_790);
xnor U667 (N_667,In_2899,In_1782);
or U668 (N_668,In_987,In_2945);
xnor U669 (N_669,In_337,In_1178);
nand U670 (N_670,In_424,In_403);
or U671 (N_671,In_1666,In_238);
and U672 (N_672,In_2653,In_1220);
or U673 (N_673,In_2881,In_12);
or U674 (N_674,In_333,In_2197);
or U675 (N_675,In_2720,In_554);
or U676 (N_676,In_2703,In_1627);
nand U677 (N_677,In_1370,In_1603);
and U678 (N_678,In_883,In_561);
nand U679 (N_679,In_2305,In_2933);
and U680 (N_680,In_1476,In_2131);
or U681 (N_681,In_384,In_1371);
nand U682 (N_682,In_447,In_812);
nor U683 (N_683,In_2794,In_755);
nand U684 (N_684,In_1297,In_2000);
xor U685 (N_685,In_2749,In_1037);
and U686 (N_686,In_481,In_706);
and U687 (N_687,In_1817,In_159);
and U688 (N_688,In_1981,In_628);
or U689 (N_689,In_2215,In_1979);
or U690 (N_690,In_1540,In_1449);
and U691 (N_691,In_1300,In_1671);
nor U692 (N_692,In_2579,In_362);
xnor U693 (N_693,In_2112,In_1171);
and U694 (N_694,In_929,In_816);
and U695 (N_695,In_2973,In_1196);
or U696 (N_696,In_282,In_1861);
nand U697 (N_697,In_1653,In_2475);
or U698 (N_698,In_2976,In_882);
nor U699 (N_699,In_106,In_741);
or U700 (N_700,In_2713,In_2148);
or U701 (N_701,In_718,In_1007);
nand U702 (N_702,In_1001,In_1687);
nand U703 (N_703,In_1207,In_2595);
nor U704 (N_704,In_972,In_234);
xor U705 (N_705,In_318,In_557);
nor U706 (N_706,In_269,In_983);
and U707 (N_707,In_2485,In_1903);
xor U708 (N_708,In_1664,In_2376);
nor U709 (N_709,In_2326,In_1035);
and U710 (N_710,In_981,In_1789);
xor U711 (N_711,In_96,In_2403);
or U712 (N_712,In_1121,In_2647);
nor U713 (N_713,In_1077,In_902);
nor U714 (N_714,In_1038,In_2719);
xnor U715 (N_715,In_2497,In_1000);
nand U716 (N_716,In_2138,In_1087);
nor U717 (N_717,In_2077,In_742);
or U718 (N_718,In_2210,In_2266);
or U719 (N_719,In_1103,In_841);
nand U720 (N_720,In_2805,In_286);
or U721 (N_721,In_2548,In_1119);
and U722 (N_722,In_1195,In_2469);
and U723 (N_723,In_252,In_1952);
and U724 (N_724,In_1581,In_293);
nor U725 (N_725,In_1850,In_2486);
nand U726 (N_726,In_284,In_1382);
nand U727 (N_727,In_2833,In_573);
or U728 (N_728,In_2975,In_2682);
and U729 (N_729,In_169,In_419);
and U730 (N_730,In_775,In_2958);
nand U731 (N_731,In_2861,In_1792);
nand U732 (N_732,In_2550,In_875);
nor U733 (N_733,In_262,In_2961);
nor U734 (N_734,In_721,In_400);
or U735 (N_735,In_2951,In_1810);
or U736 (N_736,In_2115,In_2268);
nand U737 (N_737,In_2365,In_2659);
or U738 (N_738,In_1932,In_659);
or U739 (N_739,In_973,In_496);
nor U740 (N_740,In_9,In_1088);
nor U741 (N_741,In_1934,In_959);
nand U742 (N_742,In_367,In_2606);
nor U743 (N_743,In_1135,In_2363);
nand U744 (N_744,In_324,In_2379);
nand U745 (N_745,In_1270,In_64);
or U746 (N_746,In_2388,In_507);
nor U747 (N_747,In_2427,In_2393);
or U748 (N_748,In_1271,In_171);
nand U749 (N_749,In_909,In_717);
nor U750 (N_750,In_1474,In_1468);
nand U751 (N_751,In_119,In_2641);
and U752 (N_752,In_1028,In_2194);
and U753 (N_753,In_708,In_633);
and U754 (N_754,In_2297,In_2196);
nand U755 (N_755,In_2304,In_2792);
nor U756 (N_756,In_2123,In_1328);
nand U757 (N_757,In_2611,In_91);
xnor U758 (N_758,In_2987,In_2261);
and U759 (N_759,In_66,In_1930);
or U760 (N_760,In_2472,In_2696);
xnor U761 (N_761,In_510,In_980);
nand U762 (N_762,In_255,In_836);
xnor U763 (N_763,In_1031,In_2385);
nand U764 (N_764,In_393,In_570);
and U765 (N_765,In_2083,In_1255);
or U766 (N_766,In_381,In_906);
xor U767 (N_767,In_13,In_54);
or U768 (N_768,In_2434,In_2490);
xnor U769 (N_769,In_1536,In_1706);
or U770 (N_770,In_2740,In_1543);
and U771 (N_771,In_1916,In_1859);
nand U772 (N_772,In_356,In_261);
nand U773 (N_773,In_493,In_310);
and U774 (N_774,In_1229,In_1493);
nand U775 (N_775,In_439,In_1899);
or U776 (N_776,In_1853,In_1624);
xnor U777 (N_777,In_963,In_866);
and U778 (N_778,In_2533,In_1241);
and U779 (N_779,In_942,In_217);
and U780 (N_780,In_211,In_2264);
and U781 (N_781,In_1539,In_1473);
nor U782 (N_782,In_2096,In_1855);
and U783 (N_783,In_1722,In_2206);
xor U784 (N_784,In_2681,In_967);
nand U785 (N_785,In_387,In_1256);
or U786 (N_786,In_369,In_528);
or U787 (N_787,In_181,In_1023);
nand U788 (N_788,In_1989,In_418);
and U789 (N_789,In_1752,In_118);
nor U790 (N_790,In_2994,In_205);
nand U791 (N_791,In_1608,In_1738);
and U792 (N_792,In_2598,In_1319);
xnor U793 (N_793,In_804,In_2574);
nand U794 (N_794,In_597,In_1354);
and U795 (N_795,In_707,In_1948);
xor U796 (N_796,In_2501,In_82);
xnor U797 (N_797,In_2387,In_2225);
and U798 (N_798,In_756,In_591);
and U799 (N_799,In_2098,In_436);
nor U800 (N_800,In_265,In_1439);
xor U801 (N_801,In_2232,In_2842);
or U802 (N_802,In_543,In_233);
or U803 (N_803,In_2565,In_693);
or U804 (N_804,In_958,In_29);
xor U805 (N_805,In_248,In_2531);
and U806 (N_806,In_2569,In_375);
and U807 (N_807,In_325,In_451);
nor U808 (N_808,In_71,In_1643);
and U809 (N_809,In_406,In_2185);
and U810 (N_810,In_1454,In_2846);
or U811 (N_811,In_1909,In_392);
nand U812 (N_812,In_840,In_2048);
nand U813 (N_813,In_110,In_1394);
and U814 (N_814,In_935,In_857);
and U815 (N_815,In_1221,In_1827);
nor U816 (N_816,In_1243,In_272);
nor U817 (N_817,In_2400,In_202);
or U818 (N_818,In_587,In_23);
nand U819 (N_819,In_2126,In_806);
xor U820 (N_820,In_2,In_1593);
nand U821 (N_821,In_1558,In_564);
nor U822 (N_822,In_2106,In_2213);
or U823 (N_823,In_2425,In_2785);
nor U824 (N_824,In_276,In_2037);
and U825 (N_825,In_1683,In_2458);
nor U826 (N_826,In_630,In_2249);
nor U827 (N_827,In_2836,In_2315);
xor U828 (N_828,In_1884,In_1869);
and U829 (N_829,In_997,In_2626);
nor U830 (N_830,In_968,In_523);
xor U831 (N_831,In_2229,In_2017);
nand U832 (N_832,In_525,In_2397);
nand U833 (N_833,In_646,In_517);
and U834 (N_834,In_1715,In_1502);
nand U835 (N_835,In_1095,In_2331);
and U836 (N_836,In_1284,In_48);
xor U837 (N_837,In_1496,In_482);
nand U838 (N_838,In_2150,In_865);
and U839 (N_839,In_2580,In_2759);
nor U840 (N_840,In_1615,In_1231);
and U841 (N_841,In_1525,In_377);
nor U842 (N_842,In_904,In_1825);
nor U843 (N_843,In_2360,In_43);
xor U844 (N_844,In_2998,In_2654);
nand U845 (N_845,In_1436,In_2218);
xor U846 (N_846,In_2338,In_2594);
xnor U847 (N_847,In_65,In_2566);
or U848 (N_848,In_2030,In_1719);
and U849 (N_849,In_1610,In_2224);
or U850 (N_850,In_136,In_2129);
xor U851 (N_851,In_735,In_1094);
xnor U852 (N_852,In_1324,In_2640);
nor U853 (N_853,In_1745,In_2345);
and U854 (N_854,In_694,In_1184);
nand U855 (N_855,In_1640,In_228);
xnor U856 (N_856,In_2160,In_1492);
xnor U857 (N_857,In_1079,In_1734);
xnor U858 (N_858,In_681,In_2718);
xnor U859 (N_859,In_343,In_2959);
xor U860 (N_860,In_363,In_1910);
nor U861 (N_861,In_2677,In_2835);
xnor U862 (N_862,In_2500,In_2784);
and U863 (N_863,In_2353,In_2791);
and U864 (N_864,In_701,In_1962);
nand U865 (N_865,In_2180,In_1047);
or U866 (N_866,In_2134,In_2555);
xor U867 (N_867,In_1918,In_1332);
nor U868 (N_868,In_246,In_1338);
nor U869 (N_869,In_2863,In_1842);
or U870 (N_870,In_647,In_2275);
and U871 (N_871,In_642,In_1359);
or U872 (N_872,In_2724,In_2889);
and U873 (N_873,In_1156,In_214);
and U874 (N_874,In_1697,In_1938);
or U875 (N_875,In_98,In_1995);
nand U876 (N_876,In_1954,In_2139);
nor U877 (N_877,In_1310,In_1482);
nor U878 (N_878,In_1702,In_661);
nand U879 (N_879,In_809,In_2983);
or U880 (N_880,In_763,In_116);
xor U881 (N_881,In_417,In_1216);
nor U882 (N_882,In_2668,In_1083);
xor U883 (N_883,In_2816,In_2312);
xnor U884 (N_884,In_1285,In_409);
xnor U885 (N_885,In_273,In_2449);
nor U886 (N_886,In_2118,In_271);
and U887 (N_887,In_2617,In_2381);
xor U888 (N_888,In_1572,In_1870);
and U889 (N_889,In_1513,In_2303);
nand U890 (N_890,In_1500,In_1403);
and U891 (N_891,In_521,In_2323);
nand U892 (N_892,In_2882,In_1835);
nand U893 (N_893,In_412,In_338);
or U894 (N_894,In_1081,In_2796);
or U895 (N_895,In_2337,In_2511);
and U896 (N_896,In_1793,In_1043);
nor U897 (N_897,In_2060,In_1089);
xor U898 (N_898,In_2473,In_1969);
and U899 (N_899,In_1398,In_2839);
xor U900 (N_900,In_2247,In_584);
and U901 (N_901,In_1642,In_2001);
or U902 (N_902,In_221,In_31);
nand U903 (N_903,In_2693,In_1804);
nor U904 (N_904,In_1588,In_758);
or U905 (N_905,In_2090,In_2329);
and U906 (N_906,In_1068,In_527);
xnor U907 (N_907,In_267,In_22);
xor U908 (N_908,In_2314,In_2404);
nand U909 (N_909,In_1811,In_2926);
nand U910 (N_910,In_940,In_36);
nand U911 (N_911,In_2058,In_1278);
nor U912 (N_912,In_1426,In_1788);
xnor U913 (N_913,In_985,In_2806);
xor U914 (N_914,In_2189,In_1921);
and U915 (N_915,In_1011,In_2774);
nor U916 (N_916,In_2047,In_1876);
xnor U917 (N_917,In_2823,In_2166);
and U918 (N_918,In_1786,In_1305);
nor U919 (N_919,In_2518,In_1933);
xor U920 (N_920,In_2066,In_253);
xor U921 (N_921,In_1102,In_956);
nor U922 (N_922,In_2822,In_219);
or U923 (N_923,In_722,In_1967);
nor U924 (N_924,In_2114,In_1471);
or U925 (N_925,In_2684,In_2221);
and U926 (N_926,In_2319,In_1072);
nand U927 (N_927,In_583,In_685);
xnor U928 (N_928,In_2967,In_2537);
xnor U929 (N_929,In_100,In_1645);
xnor U930 (N_930,In_1589,In_2251);
xnor U931 (N_931,In_2619,In_1182);
or U932 (N_932,In_1041,In_2979);
or U933 (N_933,In_2572,In_921);
xor U934 (N_934,In_1621,In_2389);
xor U935 (N_935,In_920,In_2698);
and U936 (N_936,In_602,In_2671);
xnor U937 (N_937,In_1075,In_79);
nor U938 (N_938,In_1551,In_885);
and U939 (N_939,In_2038,In_610);
nor U940 (N_940,In_69,In_250);
nand U941 (N_941,In_651,In_1269);
nor U942 (N_942,In_461,In_874);
xor U943 (N_943,In_677,In_299);
nor U944 (N_944,In_14,In_861);
nand U945 (N_945,In_154,In_969);
xor U946 (N_946,In_162,In_73);
and U947 (N_947,In_2499,In_1998);
or U948 (N_948,In_1685,In_430);
nand U949 (N_949,In_2293,In_304);
nand U950 (N_950,In_1061,In_2664);
or U951 (N_951,In_723,In_1684);
or U952 (N_952,In_2298,In_2321);
nor U953 (N_953,In_479,In_1723);
nand U954 (N_954,In_632,In_241);
nor U955 (N_955,In_1296,In_1574);
or U956 (N_956,In_2678,In_1686);
nor U957 (N_957,In_1947,In_1957);
and U958 (N_958,In_2484,In_1839);
and U959 (N_959,In_711,In_200);
and U960 (N_960,In_1188,In_2005);
nor U961 (N_961,In_907,In_805);
and U962 (N_962,In_2706,In_678);
nand U963 (N_963,In_2950,In_2527);
nor U964 (N_964,In_2466,In_1652);
nor U965 (N_965,In_2260,In_1294);
xnor U966 (N_966,In_2903,In_716);
nand U967 (N_967,In_1871,In_2177);
or U968 (N_968,In_2471,In_108);
nand U969 (N_969,In_2291,In_578);
xor U970 (N_970,In_2366,In_1448);
nor U971 (N_971,In_1130,In_2193);
or U972 (N_972,In_1277,In_2477);
xnor U973 (N_973,In_672,In_1906);
and U974 (N_974,In_1321,In_1937);
nand U975 (N_975,In_1770,In_242);
and U976 (N_976,In_2559,In_903);
xor U977 (N_977,In_1265,In_164);
or U978 (N_978,In_1563,In_2241);
xor U979 (N_979,In_2300,In_1440);
and U980 (N_980,In_2084,In_950);
nand U981 (N_981,In_1198,In_2909);
nor U982 (N_982,In_1129,In_752);
and U983 (N_983,In_2588,In_867);
xor U984 (N_984,In_1209,In_1807);
and U985 (N_985,In_76,In_1263);
nand U986 (N_986,In_2968,In_2928);
and U987 (N_987,In_429,In_2990);
or U988 (N_988,In_1261,In_1679);
xor U989 (N_989,In_2453,In_2773);
and U990 (N_990,In_2391,In_1453);
and U991 (N_991,In_791,In_1756);
nand U992 (N_992,In_627,In_1845);
xnor U993 (N_993,In_2809,In_2932);
nand U994 (N_994,In_1986,In_2301);
nand U995 (N_995,In_1818,In_2571);
nor U996 (N_996,In_1949,In_2876);
nor U997 (N_997,In_1344,In_1266);
nand U998 (N_998,In_2292,In_1082);
or U999 (N_999,In_1356,In_794);
or U1000 (N_1000,In_349,N_327);
nand U1001 (N_1001,N_63,In_132);
or U1002 (N_1002,In_88,N_584);
xor U1003 (N_1003,In_1898,In_21);
nand U1004 (N_1004,In_2219,In_772);
xor U1005 (N_1005,In_2730,In_1744);
nand U1006 (N_1006,N_764,In_537);
or U1007 (N_1007,In_2906,N_611);
nand U1008 (N_1008,N_779,In_176);
or U1009 (N_1009,N_305,In_2125);
nor U1010 (N_1010,In_943,N_150);
nor U1011 (N_1011,N_83,N_130);
nand U1012 (N_1012,In_471,N_988);
and U1013 (N_1013,In_388,In_511);
or U1014 (N_1014,In_2622,N_682);
nand U1015 (N_1015,N_939,N_484);
nor U1016 (N_1016,In_2524,In_1985);
nor U1017 (N_1017,In_1523,In_2496);
nor U1018 (N_1018,In_2607,N_959);
nand U1019 (N_1019,N_981,N_30);
xor U1020 (N_1020,In_444,In_1888);
and U1021 (N_1021,In_1802,N_900);
nand U1022 (N_1022,In_45,N_567);
nor U1023 (N_1023,In_475,N_366);
xor U1024 (N_1024,N_753,N_465);
xor U1025 (N_1025,In_1046,In_2020);
nand U1026 (N_1026,N_646,N_756);
or U1027 (N_1027,In_1533,In_1250);
xor U1028 (N_1028,In_2980,In_103);
nor U1029 (N_1029,In_1217,N_417);
or U1030 (N_1030,N_24,In_2739);
or U1031 (N_1031,In_2006,In_2026);
nand U1032 (N_1032,In_459,N_521);
nor U1033 (N_1033,N_241,In_2435);
or U1034 (N_1034,In_2915,N_291);
and U1035 (N_1035,N_159,N_823);
or U1036 (N_1036,In_1959,N_675);
nor U1037 (N_1037,N_459,N_18);
and U1038 (N_1038,N_258,N_555);
and U1039 (N_1039,N_0,N_341);
or U1040 (N_1040,N_609,N_236);
nand U1041 (N_1041,In_5,N_841);
and U1042 (N_1042,In_1747,In_1760);
nand U1043 (N_1043,N_588,In_1215);
and U1044 (N_1044,N_397,N_804);
xor U1045 (N_1045,N_902,N_836);
or U1046 (N_1046,In_2732,N_479);
xnor U1047 (N_1047,In_555,In_1675);
and U1048 (N_1048,In_1092,In_2355);
xnor U1049 (N_1049,N_961,N_919);
and U1050 (N_1050,N_784,N_73);
and U1051 (N_1051,N_577,N_32);
nor U1052 (N_1052,In_1460,In_1469);
or U1053 (N_1053,N_363,N_903);
nand U1054 (N_1054,N_447,In_1292);
nor U1055 (N_1055,In_502,In_410);
and U1056 (N_1056,In_715,N_904);
nor U1057 (N_1057,In_803,In_2147);
nand U1058 (N_1058,N_590,N_40);
nor U1059 (N_1059,In_2021,In_3);
nor U1060 (N_1060,N_37,N_109);
and U1061 (N_1061,N_944,In_1334);
and U1062 (N_1062,In_732,In_1350);
and U1063 (N_1063,In_1058,In_824);
and U1064 (N_1064,N_532,N_982);
xor U1065 (N_1065,In_41,N_145);
xnor U1066 (N_1066,N_834,In_1239);
or U1067 (N_1067,In_134,N_998);
and U1068 (N_1068,In_787,In_2445);
nand U1069 (N_1069,In_1412,N_286);
and U1070 (N_1070,N_255,In_1237);
nand U1071 (N_1071,N_14,N_833);
nor U1072 (N_1072,In_1174,N_249);
or U1073 (N_1073,N_411,In_2692);
and U1074 (N_1074,In_1823,N_580);
nor U1075 (N_1075,N_519,In_2642);
or U1076 (N_1076,N_106,In_2234);
and U1077 (N_1077,N_837,In_2488);
and U1078 (N_1078,In_2931,In_1289);
xnor U1079 (N_1079,In_1599,N_811);
nand U1080 (N_1080,N_140,N_882);
xnor U1081 (N_1081,In_1805,In_515);
and U1082 (N_1082,N_325,N_138);
nand U1083 (N_1083,N_490,In_2821);
xnor U1084 (N_1084,In_1554,In_2010);
or U1085 (N_1085,N_516,In_2451);
nor U1086 (N_1086,N_414,In_2639);
xnor U1087 (N_1087,N_781,N_520);
xor U1088 (N_1088,In_2437,In_2995);
and U1089 (N_1089,N_283,In_443);
or U1090 (N_1090,N_825,N_463);
nor U1091 (N_1091,In_53,In_888);
nor U1092 (N_1092,N_443,N_565);
and U1093 (N_1093,In_25,In_910);
nor U1094 (N_1094,N_574,N_579);
nor U1095 (N_1095,N_649,N_347);
xor U1096 (N_1096,In_1116,N_776);
or U1097 (N_1097,In_1795,In_1531);
or U1098 (N_1098,In_309,N_774);
nand U1099 (N_1099,In_813,N_300);
nor U1100 (N_1100,N_754,N_458);
or U1101 (N_1101,N_438,N_543);
nand U1102 (N_1102,In_1562,In_689);
and U1103 (N_1103,N_2,In_1234);
and U1104 (N_1104,In_834,N_313);
xnor U1105 (N_1105,In_2680,In_458);
and U1106 (N_1106,N_388,In_2144);
nand U1107 (N_1107,N_268,In_1096);
nand U1108 (N_1108,N_566,In_1755);
nand U1109 (N_1109,In_828,In_1109);
nor U1110 (N_1110,N_620,N_715);
and U1111 (N_1111,N_663,In_2627);
nor U1112 (N_1112,N_743,N_999);
or U1113 (N_1113,In_2999,N_108);
xor U1114 (N_1114,In_2940,In_635);
and U1115 (N_1115,N_600,N_434);
nor U1116 (N_1116,In_1750,In_1409);
and U1117 (N_1117,N_420,In_4);
and U1118 (N_1118,N_133,N_911);
nor U1119 (N_1119,N_701,N_142);
and U1120 (N_1120,In_2631,N_801);
and U1121 (N_1121,In_278,In_210);
and U1122 (N_1122,In_2877,N_147);
or U1123 (N_1123,N_707,N_129);
or U1124 (N_1124,In_133,N_750);
and U1125 (N_1125,In_173,N_19);
and U1126 (N_1126,In_1628,N_167);
nand U1127 (N_1127,In_2553,N_713);
xnor U1128 (N_1128,N_791,N_309);
and U1129 (N_1129,N_28,N_968);
xnor U1130 (N_1130,N_780,In_1834);
xor U1131 (N_1131,In_1022,In_1661);
xor U1132 (N_1132,N_627,In_1301);
xnor U1133 (N_1133,In_1883,In_207);
or U1134 (N_1134,In_1307,N_31);
nor U1135 (N_1135,N_830,In_2695);
nor U1136 (N_1136,In_1881,N_412);
nand U1137 (N_1137,N_410,In_1922);
nand U1138 (N_1138,N_86,In_1419);
or U1139 (N_1139,In_2599,N_739);
xor U1140 (N_1140,N_728,In_2252);
nor U1141 (N_1141,N_936,In_1124);
nand U1142 (N_1142,In_2702,In_1431);
or U1143 (N_1143,In_1549,N_890);
or U1144 (N_1144,N_351,In_2767);
nor U1145 (N_1145,In_1441,In_2432);
and U1146 (N_1146,N_812,N_908);
nor U1147 (N_1147,In_898,N_918);
nand U1148 (N_1148,In_979,In_2941);
nand U1149 (N_1149,In_714,N_460);
nand U1150 (N_1150,N_42,In_575);
and U1151 (N_1151,In_886,N_334);
nand U1152 (N_1152,In_640,N_170);
nor U1153 (N_1153,N_500,In_2715);
or U1154 (N_1154,In_975,N_552);
nor U1155 (N_1155,In_1224,N_321);
or U1156 (N_1156,In_529,N_72);
or U1157 (N_1157,N_554,In_2436);
nand U1158 (N_1158,N_891,In_1753);
nor U1159 (N_1159,In_2507,N_881);
nor U1160 (N_1160,N_861,N_183);
nor U1161 (N_1161,N_669,In_216);
nand U1162 (N_1162,In_1506,N_551);
nand U1163 (N_1163,N_466,In_1470);
nand U1164 (N_1164,In_305,N_820);
nand U1165 (N_1165,N_700,In_522);
nand U1166 (N_1166,In_1364,In_1418);
and U1167 (N_1167,In_2879,In_2045);
xnor U1168 (N_1168,N_79,In_120);
xor U1169 (N_1169,N_690,N_474);
nand U1170 (N_1170,N_243,In_2154);
and U1171 (N_1171,N_204,In_1649);
xnor U1172 (N_1172,N_477,In_2491);
xor U1173 (N_1173,N_905,N_909);
and U1174 (N_1174,In_1042,In_1281);
or U1175 (N_1175,In_378,In_2539);
nand U1176 (N_1176,In_1619,N_851);
xnor U1177 (N_1177,In_160,N_467);
xnor U1178 (N_1178,N_835,In_624);
nand U1179 (N_1179,In_1641,N_61);
nor U1180 (N_1180,In_652,In_2583);
and U1181 (N_1181,N_828,N_696);
nand U1182 (N_1182,In_89,In_1965);
nand U1183 (N_1183,N_238,In_580);
xnor U1184 (N_1184,In_2561,N_992);
or U1185 (N_1185,N_95,In_1875);
xor U1186 (N_1186,In_2087,N_342);
and U1187 (N_1187,N_966,N_857);
and U1188 (N_1188,In_2417,N_180);
or U1189 (N_1189,In_1490,In_1189);
nor U1190 (N_1190,In_2897,N_893);
nand U1191 (N_1191,N_288,In_1333);
and U1192 (N_1192,In_881,N_608);
and U1193 (N_1193,In_1445,N_15);
or U1194 (N_1194,In_2853,N_263);
and U1195 (N_1195,In_2056,N_668);
xnor U1196 (N_1196,N_480,In_1616);
xnor U1197 (N_1197,In_2277,In_514);
xnor U1198 (N_1198,In_1841,N_271);
and U1199 (N_1199,In_1098,In_2573);
xnor U1200 (N_1200,N_261,N_124);
and U1201 (N_1201,In_1210,N_11);
nor U1202 (N_1202,N_483,In_807);
and U1203 (N_1203,In_2576,N_974);
nor U1204 (N_1204,In_330,In_1365);
or U1205 (N_1205,N_657,N_508);
nor U1206 (N_1206,N_302,In_203);
xnor U1207 (N_1207,N_278,N_494);
nand U1208 (N_1208,In_1660,N_749);
nor U1209 (N_1209,In_604,N_260);
nand U1210 (N_1210,N_176,In_1530);
and U1211 (N_1211,In_2534,In_923);
nand U1212 (N_1212,In_1863,N_113);
nor U1213 (N_1213,In_2875,N_610);
or U1214 (N_1214,In_1219,In_2643);
nor U1215 (N_1215,N_237,N_925);
and U1216 (N_1216,N_762,In_1367);
nand U1217 (N_1217,N_832,N_253);
nand U1218 (N_1218,N_132,In_402);
nor U1219 (N_1219,In_2766,In_1538);
xnor U1220 (N_1220,N_643,In_2122);
xor U1221 (N_1221,N_57,N_77);
nand U1222 (N_1222,N_115,N_658);
nand U1223 (N_1223,In_1889,N_615);
or U1224 (N_1224,In_2029,N_373);
nand U1225 (N_1225,In_2503,In_1880);
nor U1226 (N_1226,In_334,N_210);
and U1227 (N_1227,In_1245,N_429);
nor U1228 (N_1228,N_67,In_190);
nand U1229 (N_1229,In_1314,N_693);
nand U1230 (N_1230,In_2772,In_674);
and U1231 (N_1231,N_938,N_993);
xnor U1232 (N_1232,In_2672,In_2367);
nand U1233 (N_1233,N_990,In_1896);
nor U1234 (N_1234,In_317,In_1099);
xnor U1235 (N_1235,N_116,In_1980);
nor U1236 (N_1236,In_793,N_287);
or U1237 (N_1237,N_654,N_957);
and U1238 (N_1238,In_1577,In_1002);
xnor U1239 (N_1239,N_547,In_1070);
and U1240 (N_1240,N_499,N_738);
nor U1241 (N_1241,In_1150,In_478);
and U1242 (N_1242,In_328,In_2824);
nand U1243 (N_1243,N_296,In_438);
nor U1244 (N_1244,In_2633,N_378);
nor U1245 (N_1245,In_2068,In_6);
and U1246 (N_1246,N_767,In_344);
nor U1247 (N_1247,In_24,N_534);
nand U1248 (N_1248,In_432,N_361);
nand U1249 (N_1249,In_889,N_9);
xnor U1250 (N_1250,N_34,N_187);
nand U1251 (N_1251,N_783,N_651);
nor U1252 (N_1252,N_793,N_175);
nor U1253 (N_1253,N_105,N_585);
xor U1254 (N_1254,N_156,In_1882);
and U1255 (N_1255,In_201,N_403);
xnor U1256 (N_1256,N_62,In_626);
nor U1257 (N_1257,In_93,N_813);
xnor U1258 (N_1258,In_590,N_433);
nor U1259 (N_1259,In_2544,N_949);
and U1260 (N_1260,N_848,In_850);
nand U1261 (N_1261,In_189,In_2476);
nor U1262 (N_1262,N_879,N_171);
xor U1263 (N_1263,In_655,N_724);
or U1264 (N_1264,N_69,N_583);
nor U1265 (N_1265,In_194,In_877);
nand U1266 (N_1266,In_931,In_2299);
nor U1267 (N_1267,N_324,In_949);
and U1268 (N_1268,In_1114,In_394);
nor U1269 (N_1269,In_1013,In_1341);
xnor U1270 (N_1270,In_2478,In_1408);
nor U1271 (N_1271,In_2508,In_2536);
xnor U1272 (N_1272,N_575,In_302);
xor U1273 (N_1273,N_284,N_144);
or U1274 (N_1274,In_810,N_768);
xnor U1275 (N_1275,N_969,N_729);
xnor U1276 (N_1276,In_1866,In_495);
nor U1277 (N_1277,N_561,N_310);
and U1278 (N_1278,N_978,In_2351);
and U1279 (N_1279,In_670,In_568);
and U1280 (N_1280,N_201,N_640);
nand U1281 (N_1281,In_2510,In_2768);
and U1282 (N_1282,In_1973,N_336);
nand U1283 (N_1283,N_872,N_942);
xnor U1284 (N_1284,In_2691,N_424);
and U1285 (N_1285,N_164,N_346);
nor U1286 (N_1286,N_89,N_205);
nand U1287 (N_1287,N_368,In_1049);
and U1288 (N_1288,In_236,In_1026);
or U1289 (N_1289,N_442,In_1499);
nand U1290 (N_1290,N_307,N_216);
nand U1291 (N_1291,N_413,N_504);
nand U1292 (N_1292,N_141,In_679);
and U1293 (N_1293,N_267,In_858);
or U1294 (N_1294,N_456,N_110);
xor U1295 (N_1295,N_228,In_1944);
nor U1296 (N_1296,In_2294,N_556);
nand U1297 (N_1297,In_1780,In_2327);
xnor U1298 (N_1298,In_676,In_208);
nor U1299 (N_1299,In_1868,N_899);
or U1300 (N_1300,In_2955,N_592);
and U1301 (N_1301,N_497,In_2254);
xor U1302 (N_1302,N_349,N_597);
nor U1303 (N_1303,N_695,In_1066);
nor U1304 (N_1304,In_1739,N_319);
nand U1305 (N_1305,N_408,N_104);
and U1306 (N_1306,In_472,N_970);
xnor U1307 (N_1307,N_119,In_2346);
nor U1308 (N_1308,In_649,N_248);
or U1309 (N_1309,N_572,N_818);
xor U1310 (N_1310,N_482,N_867);
or U1311 (N_1311,N_430,In_497);
nor U1312 (N_1312,In_2971,N_436);
or U1313 (N_1313,N_873,N_810);
nand U1314 (N_1314,In_2110,N_274);
nor U1315 (N_1315,In_2964,In_2456);
nand U1316 (N_1316,N_887,In_1347);
or U1317 (N_1317,N_163,N_404);
nand U1318 (N_1318,In_1516,In_1721);
and U1319 (N_1319,In_1402,N_343);
xor U1320 (N_1320,In_2168,In_2929);
nand U1321 (N_1321,N_796,N_514);
nand U1322 (N_1322,In_2802,N_963);
xnor U1323 (N_1323,N_672,In_2494);
nand U1324 (N_1324,In_1395,In_1725);
and U1325 (N_1325,N_470,In_2908);
nor U1326 (N_1326,In_1226,N_621);
or U1327 (N_1327,N_568,N_265);
or U1328 (N_1328,In_149,In_2015);
nand U1329 (N_1329,In_2890,N_849);
xor U1330 (N_1330,N_365,In_2099);
and U1331 (N_1331,In_2666,In_1056);
and U1332 (N_1332,N_234,N_364);
or U1333 (N_1333,In_1004,In_1413);
xnor U1334 (N_1334,In_687,In_2433);
xnor U1335 (N_1335,N_950,In_1983);
nor U1336 (N_1336,In_505,In_11);
and U1337 (N_1337,N_956,N_282);
or U1338 (N_1338,N_359,In_2965);
or U1339 (N_1339,In_476,N_855);
nand U1340 (N_1340,In_2554,N_207);
nand U1341 (N_1341,N_569,In_1663);
nand U1342 (N_1342,In_2716,N_977);
or U1343 (N_1343,N_44,In_1665);
xnor U1344 (N_1344,In_1724,N_94);
or U1345 (N_1345,N_16,N_85);
nor U1346 (N_1346,In_1515,In_1691);
nor U1347 (N_1347,N_752,N_421);
nand U1348 (N_1348,N_613,In_1781);
xnor U1349 (N_1349,N_578,N_212);
nor U1350 (N_1350,In_474,In_477);
and U1351 (N_1351,In_2850,In_2078);
nand U1352 (N_1352,N_154,N_888);
xor U1353 (N_1353,N_233,In_736);
or U1354 (N_1354,In_1480,N_318);
nor U1355 (N_1355,N_614,In_1484);
nand U1356 (N_1356,N_392,In_121);
and U1357 (N_1357,In_473,In_566);
nand U1358 (N_1358,N_20,In_1604);
xnor U1359 (N_1359,In_1057,In_99);
and U1360 (N_1360,N_496,N_435);
and U1361 (N_1361,N_495,In_2382);
xor U1362 (N_1362,In_243,In_1093);
and U1363 (N_1363,N_515,N_557);
nor U1364 (N_1364,N_462,N_702);
nand U1365 (N_1365,In_2269,N_639);
or U1366 (N_1366,N_68,In_1064);
nand U1367 (N_1367,In_2074,In_1164);
nand U1368 (N_1368,N_708,N_379);
and U1369 (N_1369,In_8,In_918);
xor U1370 (N_1370,N_720,In_2283);
nor U1371 (N_1371,N_375,N_522);
or U1372 (N_1372,In_1994,N_634);
nor U1373 (N_1373,In_535,N_127);
nor U1374 (N_1374,N_790,In_2246);
nand U1375 (N_1375,N_576,In_1040);
nand U1376 (N_1376,N_647,N_795);
nor U1377 (N_1377,N_316,N_224);
or U1378 (N_1378,N_437,N_446);
nand U1379 (N_1379,In_300,N_755);
or U1380 (N_1380,N_314,N_965);
or U1381 (N_1381,N_935,In_1860);
and U1382 (N_1382,In_1758,In_2288);
nand U1383 (N_1383,In_1194,In_2557);
and U1384 (N_1384,In_1213,In_42);
nand U1385 (N_1385,In_178,In_2255);
xor U1386 (N_1386,In_2281,In_1369);
nor U1387 (N_1387,In_870,In_2086);
nor U1388 (N_1388,N_883,In_2752);
xnor U1389 (N_1389,N_719,N_488);
xnor U1390 (N_1390,N_54,In_254);
nand U1391 (N_1391,In_2033,In_2188);
nand U1392 (N_1392,N_440,N_799);
or U1393 (N_1393,In_2395,In_2380);
nor U1394 (N_1394,In_887,In_2378);
xor U1395 (N_1395,N_425,N_531);
nand U1396 (N_1396,N_122,In_879);
and U1397 (N_1397,In_1430,N_226);
nor U1398 (N_1398,In_2418,In_599);
xnor U1399 (N_1399,N_741,N_537);
xor U1400 (N_1400,In_691,N_209);
nor U1401 (N_1401,N_197,N_709);
nand U1402 (N_1402,In_2777,N_51);
nand U1403 (N_1403,In_2274,N_203);
and U1404 (N_1404,N_808,In_16);
xnor U1405 (N_1405,N_118,In_1711);
and U1406 (N_1406,N_636,N_173);
or U1407 (N_1407,In_2104,In_1016);
and U1408 (N_1408,N_391,N_338);
and U1409 (N_1409,N_865,N_571);
nor U1410 (N_1410,N_454,In_1166);
or U1411 (N_1411,N_792,In_1062);
xnor U1412 (N_1412,N_427,In_2186);
nor U1413 (N_1413,In_27,N_80);
xor U1414 (N_1414,In_1651,In_2322);
nand U1415 (N_1415,In_2263,N_798);
xnor U1416 (N_1416,In_1355,N_549);
or U1417 (N_1417,N_983,In_1242);
and U1418 (N_1418,N_725,In_1968);
or U1419 (N_1419,N_387,In_380);
nor U1420 (N_1420,In_1731,N_985);
or U1421 (N_1421,In_1459,In_1873);
or U1422 (N_1422,N_50,In_1211);
or U1423 (N_1423,N_280,N_181);
nand U1424 (N_1424,In_984,In_155);
nand U1425 (N_1425,In_1012,In_2413);
nor U1426 (N_1426,N_335,N_751);
xor U1427 (N_1427,In_2075,In_2829);
or U1428 (N_1428,N_148,N_877);
xor U1429 (N_1429,In_1422,N_328);
or U1430 (N_1430,In_988,N_97);
xor U1431 (N_1431,In_1779,In_454);
xor U1432 (N_1432,In_1345,N_923);
or U1433 (N_1433,In_851,N_892);
and U1434 (N_1434,In_87,N_689);
nand U1435 (N_1435,N_107,N_678);
nor U1436 (N_1436,N_117,In_1597);
nor U1437 (N_1437,N_996,N_475);
and U1438 (N_1438,In_901,In_695);
or U1439 (N_1439,In_462,N_995);
and U1440 (N_1440,In_1144,N_619);
nor U1441 (N_1441,N_158,In_1911);
nor U1442 (N_1442,N_311,N_652);
nor U1443 (N_1443,In_1507,N_194);
nand U1444 (N_1444,N_53,In_1214);
xnor U1445 (N_1445,N_367,N_453);
nor U1446 (N_1446,In_195,In_2661);
xor U1447 (N_1447,In_2278,In_1800);
nand U1448 (N_1448,In_2071,N_322);
and U1449 (N_1449,N_22,N_660);
xor U1450 (N_1450,N_612,In_1331);
nand U1451 (N_1451,In_2384,In_1567);
nor U1452 (N_1452,N_945,N_816);
and U1453 (N_1453,In_776,In_729);
or U1454 (N_1454,In_1806,In_1761);
or U1455 (N_1455,N_227,N_775);
nand U1456 (N_1456,In_2761,In_965);
and U1457 (N_1457,N_206,In_60);
nand U1458 (N_1458,In_158,In_2514);
nand U1459 (N_1459,N_168,In_1071);
xnor U1460 (N_1460,In_1105,N_530);
nand U1461 (N_1461,In_2628,In_2310);
xor U1462 (N_1462,In_303,In_1797);
nand U1463 (N_1463,N_222,In_1504);
and U1464 (N_1464,N_350,N_45);
nand U1465 (N_1465,In_751,N_377);
nor U1466 (N_1466,In_2624,N_174);
or U1467 (N_1467,In_2517,N_123);
or U1468 (N_1468,N_393,In_1890);
or U1469 (N_1469,In_2143,In_2285);
nand U1470 (N_1470,In_572,N_5);
nor U1471 (N_1471,N_36,N_178);
nand U1472 (N_1472,In_2439,In_365);
or U1473 (N_1473,In_1659,In_2362);
nor U1474 (N_1474,In_2227,N_135);
or U1475 (N_1475,In_1152,N_599);
and U1476 (N_1476,N_853,N_431);
and U1477 (N_1477,In_2324,In_2333);
or U1478 (N_1478,N_394,N_82);
and U1479 (N_1479,In_2003,In_1151);
nand U1480 (N_1480,In_641,In_1520);
xnor U1481 (N_1481,N_606,N_676);
or U1482 (N_1482,In_2111,N_213);
or U1483 (N_1483,N_760,In_603);
nand U1484 (N_1484,N_457,N_625);
or U1485 (N_1485,N_826,N_710);
or U1486 (N_1486,N_558,N_46);
nand U1487 (N_1487,N_716,N_921);
nor U1488 (N_1488,N_445,N_423);
and U1489 (N_1489,N_422,In_2528);
or U1490 (N_1490,N_758,N_360);
nand U1491 (N_1491,N_717,N_723);
and U1492 (N_1492,N_517,N_264);
and U1493 (N_1493,In_1565,In_2632);
or U1494 (N_1494,N_279,In_404);
nand U1495 (N_1495,N_126,N_452);
nand U1496 (N_1496,N_242,N_476);
xor U1497 (N_1497,N_485,N_598);
nand U1498 (N_1498,N_455,In_2493);
nor U1499 (N_1499,In_1291,N_971);
nand U1500 (N_1500,In_1357,In_2912);
xor U1501 (N_1501,In_524,N_850);
nor U1502 (N_1502,N_635,N_449);
nor U1503 (N_1503,N_240,N_523);
or U1504 (N_1504,In_2948,N_674);
xor U1505 (N_1505,In_2694,In_577);
nand U1506 (N_1506,N_868,In_1303);
nor U1507 (N_1507,N_103,In_1435);
xnor U1508 (N_1508,N_87,In_1647);
xor U1509 (N_1509,In_1,N_533);
and U1510 (N_1510,In_548,N_332);
and U1511 (N_1511,N_162,In_464);
nor U1512 (N_1512,In_2513,In_826);
and U1513 (N_1513,N_230,In_1008);
xor U1514 (N_1514,In_1550,In_2273);
xor U1515 (N_1515,In_1222,N_972);
nor U1516 (N_1516,N_400,N_513);
or U1517 (N_1517,In_1442,N_289);
xnor U1518 (N_1518,N_471,In_2410);
or U1519 (N_1519,N_786,N_822);
nor U1520 (N_1520,In_2756,In_1682);
xor U1521 (N_1521,N_439,In_396);
or U1522 (N_1522,N_898,N_677);
or U1523 (N_1523,N_330,N_3);
and U1524 (N_1524,In_844,In_163);
xnor U1525 (N_1525,N_769,In_161);
xnor U1526 (N_1526,In_34,N_215);
nor U1527 (N_1527,N_542,In_2489);
and U1528 (N_1528,N_402,N_979);
xnor U1529 (N_1529,In_1078,In_2815);
nor U1530 (N_1530,In_2660,In_1991);
nor U1531 (N_1531,In_390,In_2459);
and U1532 (N_1532,N_290,In_2108);
nand U1533 (N_1533,In_2753,N_90);
and U1534 (N_1534,N_641,In_1497);
xnor U1535 (N_1535,N_623,In_38);
or U1536 (N_1536,N_711,In_213);
or U1537 (N_1537,N_856,In_1623);
nand U1538 (N_1538,N_631,In_2760);
nor U1539 (N_1539,N_896,N_540);
and U1540 (N_1540,In_2790,N_492);
xor U1541 (N_1541,N_559,In_1396);
xnor U1542 (N_1542,In_960,N_687);
xnor U1543 (N_1543,In_28,N_74);
or U1544 (N_1544,N_401,In_1602);
or U1545 (N_1545,N_847,In_1005);
or U1546 (N_1546,N_759,In_1342);
nor U1547 (N_1547,In_516,In_1939);
nand U1548 (N_1548,In_399,In_1132);
nor U1549 (N_1549,In_934,In_2452);
nor U1550 (N_1550,In_2040,In_788);
or U1551 (N_1551,In_2894,In_970);
xnor U1552 (N_1552,In_485,N_917);
or U1553 (N_1553,N_64,N_875);
xnor U1554 (N_1554,N_270,In_1678);
and U1555 (N_1555,In_1183,In_290);
nor U1556 (N_1556,N_75,In_1298);
nor U1557 (N_1557,N_880,In_2424);
and U1558 (N_1558,In_2179,N_161);
nand U1559 (N_1559,In_2697,N_186);
and U1560 (N_1560,N_510,N_871);
nor U1561 (N_1561,In_2359,In_1927);
nor U1562 (N_1562,In_227,In_843);
or U1563 (N_1563,N_656,In_2797);
xor U1564 (N_1564,N_952,In_1676);
xnor U1565 (N_1565,N_137,In_853);
nor U1566 (N_1566,In_1372,In_489);
or U1567 (N_1567,In_1583,In_899);
or U1568 (N_1568,In_1487,In_2290);
nand U1569 (N_1569,N_637,N_607);
or U1570 (N_1570,N_937,N_670);
nor U1571 (N_1571,N_831,N_560);
or U1572 (N_1572,In_2956,In_1832);
and U1573 (N_1573,In_2750,In_1942);
xnor U1574 (N_1574,In_744,In_1829);
nor U1575 (N_1575,In_312,N_844);
nor U1576 (N_1576,In_2220,In_1258);
or U1577 (N_1577,In_1335,N_329);
or U1578 (N_1578,In_559,N_539);
nand U1579 (N_1579,N_681,In_1392);
xor U1580 (N_1580,In_1736,N_415);
and U1581 (N_1581,N_337,In_1373);
nand U1582 (N_1582,In_2306,N_889);
nand U1583 (N_1583,In_2462,N_251);
and U1584 (N_1584,N_928,N_312);
nor U1585 (N_1585,In_1552,N_441);
or U1586 (N_1586,In_2717,N_787);
nand U1587 (N_1587,N_12,N_846);
xnor U1588 (N_1588,N_93,N_772);
or U1589 (N_1589,In_1961,In_779);
nand U1590 (N_1590,N_683,In_1743);
and U1591 (N_1591,N_732,In_1461);
xor U1592 (N_1592,N_933,In_1424);
nand U1593 (N_1593,N_740,N_946);
nor U1594 (N_1594,N_189,N_763);
nand U1595 (N_1595,N_102,N_217);
or U1596 (N_1596,In_2438,In_395);
and U1597 (N_1597,In_2173,In_593);
and U1598 (N_1598,N_406,N_21);
nand U1599 (N_1599,In_1348,In_2332);
or U1600 (N_1600,In_2094,N_208);
xor U1601 (N_1601,In_256,N_688);
nand U1602 (N_1602,N_317,In_1065);
nor U1603 (N_1603,N_23,In_2949);
xnor U1604 (N_1604,N_924,N_254);
xor U1605 (N_1605,N_926,N_862);
xor U1606 (N_1606,In_467,In_279);
nor U1607 (N_1607,N_852,N_941);
or U1608 (N_1608,In_192,In_2652);
xor U1609 (N_1609,N_770,In_1984);
xnor U1610 (N_1610,In_2910,In_2993);
and U1611 (N_1611,N_745,In_1501);
or U1612 (N_1612,N_536,In_608);
nor U1613 (N_1613,In_789,N_179);
xor U1614 (N_1614,N_225,N_870);
nor U1615 (N_1615,N_843,N_948);
xnor U1616 (N_1616,In_1452,N_88);
or U1617 (N_1617,In_1548,N_765);
and U1618 (N_1618,N_8,In_1252);
xnor U1619 (N_1619,N_650,In_2181);
xor U1620 (N_1620,N_38,In_925);
nor U1621 (N_1621,In_1059,In_135);
nor U1622 (N_1622,In_1455,In_1571);
xnor U1623 (N_1623,N_906,N_121);
nor U1624 (N_1624,N_778,N_33);
or U1625 (N_1625,N_252,In_607);
nand U1626 (N_1626,In_1034,N_512);
and U1627 (N_1627,In_2685,N_605);
and U1628 (N_1628,In_1822,N_815);
nand U1629 (N_1629,N_199,N_800);
xnor U1630 (N_1630,In_2396,In_1519);
nand U1631 (N_1631,N_975,N_686);
and U1632 (N_1632,In_2811,In_1232);
or U1633 (N_1633,In_896,In_2130);
or U1634 (N_1634,N_277,In_170);
and U1635 (N_1635,N_785,In_78);
nand U1636 (N_1636,N_259,N_188);
or U1637 (N_1637,N_821,N_962);
nand U1638 (N_1638,N_323,N_645);
and U1639 (N_1639,N_35,N_376);
nor U1640 (N_1640,In_186,In_798);
nor U1641 (N_1641,N_390,In_2240);
or U1642 (N_1642,In_1613,N_819);
nand U1643 (N_1643,In_2167,N_589);
or U1644 (N_1644,In_964,In_2409);
xnor U1645 (N_1645,In_1417,In_2085);
and U1646 (N_1646,In_285,In_1783);
and U1647 (N_1647,In_1601,In_833);
xor U1648 (N_1648,N_929,N_49);
xnor U1649 (N_1649,In_606,In_2034);
nor U1650 (N_1650,N_691,In_2679);
or U1651 (N_1651,In_1913,N_395);
xor U1652 (N_1652,In_2651,In_598);
xor U1653 (N_1653,N_389,In_2860);
nor U1654 (N_1654,N_71,In_1856);
xnor U1655 (N_1655,N_544,In_2922);
and U1656 (N_1656,In_374,In_2081);
nand U1657 (N_1657,In_1840,N_428);
nand U1658 (N_1658,N_794,In_452);
nor U1659 (N_1659,N_157,In_905);
nor U1660 (N_1660,In_2184,In_932);
nand U1661 (N_1661,N_727,N_464);
and U1662 (N_1662,N_742,N_444);
nor U1663 (N_1663,In_2841,N_951);
nand U1664 (N_1664,In_1975,N_845);
nand U1665 (N_1665,N_761,In_2936);
nand U1666 (N_1666,In_1374,N_60);
nor U1667 (N_1667,In_2646,In_1508);
nand U1668 (N_1668,In_2526,In_2239);
and U1669 (N_1669,N_722,In_2178);
nor U1670 (N_1670,N_806,N_503);
and U1671 (N_1671,N_782,N_838);
xnor U1672 (N_1672,N_221,In_588);
nand U1673 (N_1673,In_2913,N_6);
nor U1674 (N_1674,N_65,In_335);
and U1675 (N_1675,N_653,N_372);
nand U1676 (N_1676,In_1762,N_582);
or U1677 (N_1677,In_976,N_550);
and U1678 (N_1678,In_589,In_2865);
nand U1679 (N_1679,N_502,N_281);
xnor U1680 (N_1680,N_128,N_525);
nand U1681 (N_1681,In_2052,In_329);
or U1682 (N_1682,N_869,N_616);
nor U1683 (N_1683,N_269,N_726);
nand U1684 (N_1684,In_2442,N_374);
or U1685 (N_1685,N_184,N_468);
and U1686 (N_1686,N_354,In_35);
nand U1687 (N_1687,In_2904,N_524);
nor U1688 (N_1688,In_2461,N_736);
xnor U1689 (N_1689,N_528,N_581);
and U1690 (N_1690,N_125,In_1172);
or U1691 (N_1691,N_245,In_1688);
or U1692 (N_1692,In_1248,N_596);
or U1693 (N_1693,In_2867,N_98);
xor U1694 (N_1694,N_994,N_771);
and U1695 (N_1695,In_83,In_2414);
nand U1696 (N_1696,N_507,N_986);
nand U1697 (N_1697,In_1283,In_1894);
xor U1698 (N_1698,N_195,In_1048);
xor U1699 (N_1699,In_838,N_348);
and U1700 (N_1700,N_262,In_2101);
xnor U1701 (N_1701,N_860,In_1618);
and U1702 (N_1702,N_26,N_182);
and U1703 (N_1703,N_405,In_743);
or U1704 (N_1704,In_327,N_927);
xor U1705 (N_1705,N_59,N_735);
or U1706 (N_1706,N_353,N_247);
and U1707 (N_1707,In_1941,N_292);
or U1708 (N_1708,N_214,In_2733);
xnor U1709 (N_1709,In_616,N_564);
nand U1710 (N_1710,N_603,In_1063);
and U1711 (N_1711,N_96,In_2838);
nand U1712 (N_1712,In_2141,N_916);
nand U1713 (N_1713,N_618,In_2591);
and U1714 (N_1714,N_177,N_301);
nand U1715 (N_1715,In_1505,N_538);
nand U1716 (N_1716,In_1054,N_629);
xnor U1717 (N_1717,In_2296,N_730);
xnor U1718 (N_1718,N_25,In_822);
nand U1719 (N_1719,In_961,In_771);
or U1720 (N_1720,N_398,In_2546);
nor U1721 (N_1721,N_997,In_1966);
or U1722 (N_1722,N_381,In_1904);
nand U1723 (N_1723,In_576,In_1006);
or U1724 (N_1724,N_858,In_614);
or U1725 (N_1725,In_2295,In_2786);
or U1726 (N_1726,In_188,In_2349);
or U1727 (N_1727,In_2954,N_139);
xnor U1728 (N_1728,In_1568,N_884);
or U1729 (N_1729,In_2465,In_2764);
and U1730 (N_1730,In_326,In_585);
xnor U1731 (N_1731,In_1564,N_626);
nand U1732 (N_1732,In_2209,In_667);
xnor U1733 (N_1733,In_2969,N_897);
nor U1734 (N_1734,N_747,In_764);
nor U1735 (N_1735,N_601,N_748);
and U1736 (N_1736,In_690,In_2586);
nor U1737 (N_1737,In_2064,N_92);
nor U1738 (N_1738,In_172,In_856);
nand U1739 (N_1739,In_193,N_914);
xor U1740 (N_1740,N_671,In_911);
nor U1741 (N_1741,In_977,N_1);
or U1742 (N_1742,N_111,In_1458);
nor U1743 (N_1743,N_943,In_2463);
nor U1744 (N_1744,N_275,N_190);
nand U1745 (N_1745,N_489,In_1033);
nor U1746 (N_1746,In_512,In_2223);
and U1747 (N_1747,N_81,In_768);
xnor U1748 (N_1748,In_1729,In_2609);
and U1749 (N_1749,N_662,In_2431);
nand U1750 (N_1750,In_287,In_1282);
xor U1751 (N_1751,In_2676,In_1854);
or U1752 (N_1752,In_892,In_52);
nand U1753 (N_1753,N_134,N_684);
nand U1754 (N_1754,N_665,In_455);
and U1755 (N_1755,N_586,In_292);
nor U1756 (N_1756,N_685,In_1200);
or U1757 (N_1757,In_612,In_864);
and U1758 (N_1758,In_433,In_2107);
and U1759 (N_1759,N_633,N_718);
nor U1760 (N_1760,In_1073,In_229);
and U1761 (N_1761,In_2105,In_797);
or U1762 (N_1762,In_2657,In_2799);
nor U1763 (N_1763,N_744,In_705);
nor U1764 (N_1764,N_953,N_706);
nor U1765 (N_1765,In_1584,N_648);
xor U1766 (N_1766,N_112,In_2735);
and U1767 (N_1767,In_727,N_491);
xor U1768 (N_1768,In_1677,N_714);
and U1769 (N_1769,In_1106,In_971);
nand U1770 (N_1770,N_661,In_1138);
xor U1771 (N_1771,N_664,N_989);
nor U1772 (N_1772,N_344,N_285);
or U1773 (N_1773,N_153,N_273);
nand U1774 (N_1774,In_2175,In_1076);
nand U1775 (N_1775,N_591,N_136);
and U1776 (N_1776,N_220,N_984);
nor U1777 (N_1777,N_562,In_1852);
nor U1778 (N_1778,N_694,N_448);
nand U1779 (N_1779,In_1815,N_101);
and U1780 (N_1780,In_2023,N_48);
nand U1781 (N_1781,In_2354,In_2874);
nor U1782 (N_1782,In_957,In_785);
xor U1783 (N_1783,In_1633,N_166);
nand U1784 (N_1784,N_757,In_2448);
and U1785 (N_1785,N_814,N_737);
nand U1786 (N_1786,N_315,In_486);
xnor U1787 (N_1787,N_160,In_1946);
xnor U1788 (N_1788,N_788,N_940);
nor U1789 (N_1789,In_1003,N_293);
and U1790 (N_1790,N_655,N_481);
nor U1791 (N_1791,In_2024,In_1069);
nand U1792 (N_1792,In_1511,In_1776);
xnor U1793 (N_1793,N_396,In_1821);
or U1794 (N_1794,In_1594,N_29);
nand U1795 (N_1795,In_1778,In_180);
or U1796 (N_1796,N_802,N_461);
nor U1797 (N_1797,N_667,In_1799);
and U1798 (N_1798,In_1411,In_2925);
or U1799 (N_1799,In_1858,N_399);
or U1800 (N_1800,N_518,In_2415);
nor U1801 (N_1801,In_2041,In_2848);
xnor U1802 (N_1802,N_91,N_146);
and U1803 (N_1803,N_306,In_2211);
nor U1804 (N_1804,N_704,N_78);
nand U1805 (N_1805,In_125,In_519);
nand U1806 (N_1806,In_437,N_545);
or U1807 (N_1807,In_1325,N_155);
and U1808 (N_1808,N_932,In_1462);
nor U1809 (N_1809,In_2826,N_680);
and U1810 (N_1810,N_384,In_1450);
nor U1811 (N_1811,N_358,N_486);
nand U1812 (N_1812,In_2157,N_131);
nand U1813 (N_1813,N_304,In_1905);
xor U1814 (N_1814,N_915,N_223);
nand U1815 (N_1815,In_138,N_55);
xor U1816 (N_1816,N_498,N_712);
and U1817 (N_1817,In_2541,In_2208);
xnor U1818 (N_1818,In_2645,In_1566);
or U1819 (N_1819,In_2421,In_710);
xor U1820 (N_1820,In_354,In_2190);
and U1821 (N_1821,In_1605,N_371);
xnor U1822 (N_1822,N_546,N_630);
nor U1823 (N_1823,In_1638,In_781);
nor U1824 (N_1824,In_2158,In_2916);
or U1825 (N_1825,In_1534,N_257);
nand U1826 (N_1826,In_862,In_1631);
or U1827 (N_1827,In_2781,N_76);
or U1828 (N_1828,N_842,N_807);
xor U1829 (N_1829,In_720,N_84);
and U1830 (N_1830,In_1849,N_548);
and U1831 (N_1831,N_246,In_2443);
nand U1832 (N_1832,In_2419,N_697);
and U1833 (N_1833,In_1902,N_419);
xnor U1834 (N_1834,In_1017,In_739);
xor U1835 (N_1835,In_2467,N_380);
xnor U1836 (N_1836,N_219,N_10);
nand U1837 (N_1837,N_256,N_356);
and U1838 (N_1838,In_2279,N_526);
and U1839 (N_1839,N_570,In_799);
nor U1840 (N_1840,N_827,In_58);
or U1841 (N_1841,N_973,N_960);
xor U1842 (N_1842,In_848,In_623);
or U1843 (N_1843,In_2238,In_2854);
or U1844 (N_1844,N_930,In_1826);
nand U1845 (N_1845,In_2578,N_803);
nor U1846 (N_1846,In_571,N_432);
nor U1847 (N_1847,N_487,In_504);
xnor U1848 (N_1848,In_1306,In_1521);
nor U1849 (N_1849,In_2498,In_2502);
nor U1850 (N_1850,In_1146,N_409);
or U1851 (N_1851,N_703,N_27);
nand U1852 (N_1852,N_931,N_407);
nor U1853 (N_1853,In_294,In_167);
or U1854 (N_1854,N_370,N_817);
nor U1855 (N_1855,N_644,N_692);
or U1856 (N_1856,In_2868,N_976);
or U1857 (N_1857,In_530,In_2934);
nor U1858 (N_1858,In_2187,In_1180);
or U1859 (N_1859,In_991,N_469);
or U1860 (N_1860,In_2009,In_2182);
xnor U1861 (N_1861,N_824,N_922);
nor U1862 (N_1862,N_805,In_1625);
or U1863 (N_1863,N_56,N_628);
xnor U1864 (N_1864,N_120,N_451);
nor U1865 (N_1865,In_1801,N_211);
and U1866 (N_1866,N_563,In_2568);
and U1867 (N_1867,N_746,N_192);
and U1868 (N_1868,N_239,N_733);
nand U1869 (N_1869,In_1637,N_987);
or U1870 (N_1870,In_1384,N_416);
or U1871 (N_1871,In_782,In_1302);
and U1872 (N_1872,In_2937,N_617);
xor U1873 (N_1873,N_840,In_1262);
and U1874 (N_1874,In_352,In_145);
nor U1875 (N_1875,N_345,In_654);
nor U1876 (N_1876,N_602,N_511);
and U1877 (N_1877,N_185,In_2953);
nor U1878 (N_1878,In_733,In_2963);
xor U1879 (N_1879,N_339,In_1510);
xor U1880 (N_1880,In_1438,N_52);
or U1881 (N_1881,N_229,N_58);
or U1882 (N_1882,N_143,N_624);
nand U1883 (N_1883,N_901,N_333);
nand U1884 (N_1884,N_232,N_196);
nor U1885 (N_1885,N_642,In_1315);
xnor U1886 (N_1886,In_2205,N_839);
xor U1887 (N_1887,N_731,N_535);
or U1888 (N_1888,N_876,N_172);
nand U1889 (N_1889,In_2390,In_2146);
nor U1890 (N_1890,N_866,N_553);
xor U1891 (N_1891,N_7,In_1206);
or U1892 (N_1892,N_426,In_2320);
nor U1893 (N_1893,In_1614,In_662);
nand U1894 (N_1894,In_2738,N_13);
and U1895 (N_1895,In_2155,N_385);
nand U1896 (N_1896,In_1160,In_1137);
and U1897 (N_1897,N_17,N_913);
and U1898 (N_1898,In_2235,N_766);
nand U1899 (N_1899,N_478,In_2673);
nor U1900 (N_1900,In_2276,In_1311);
nand U1901 (N_1901,In_1522,N_99);
nor U1902 (N_1902,In_2199,In_2872);
or U1903 (N_1903,N_679,N_964);
nand U1904 (N_1904,In_698,N_699);
and U1905 (N_1905,N_501,N_357);
or U1906 (N_1906,N_864,N_632);
nand U1907 (N_1907,N_659,In_2888);
nor U1908 (N_1908,N_369,In_955);
nand U1909 (N_1909,N_698,In_1892);
nor U1910 (N_1910,N_299,N_886);
nor U1911 (N_1911,In_2480,In_946);
or U1912 (N_1912,N_198,In_2163);
nand U1913 (N_1913,N_854,N_595);
and U1914 (N_1914,N_244,In_2504);
and U1915 (N_1915,N_874,In_2970);
and U1916 (N_1916,In_1479,N_326);
and U1917 (N_1917,N_41,In_107);
nand U1918 (N_1918,N_721,In_562);
or U1919 (N_1919,In_114,In_441);
or U1920 (N_1920,In_669,In_2145);
or U1921 (N_1921,N_912,In_774);
xor U1922 (N_1922,In_914,N_169);
nor U1923 (N_1923,N_4,In_2804);
or U1924 (N_1924,N_303,In_407);
and U1925 (N_1925,In_67,In_1886);
xor U1926 (N_1926,In_2119,N_250);
or U1927 (N_1927,N_666,N_829);
xor U1928 (N_1928,N_298,N_773);
or U1929 (N_1929,In_323,N_382);
xnor U1930 (N_1930,N_527,In_2596);
and U1931 (N_1931,In_225,In_2050);
xnor U1932 (N_1932,N_604,In_637);
xnor U1933 (N_1933,N_418,In_1717);
nor U1934 (N_1934,N_235,In_800);
nor U1935 (N_1935,N_165,N_352);
or U1936 (N_1936,N_958,In_2770);
and U1937 (N_1937,N_529,N_885);
and U1938 (N_1938,N_202,N_638);
nor U1939 (N_1939,N_276,N_947);
nor U1940 (N_1940,N_218,N_295);
nor U1941 (N_1941,N_340,In_1267);
nor U1942 (N_1942,N_894,N_331);
and U1943 (N_1943,In_863,N_863);
nor U1944 (N_1944,N_472,In_2558);
xor U1945 (N_1945,N_151,N_920);
and U1946 (N_1946,In_1759,In_2605);
nand U1947 (N_1947,In_1456,N_493);
or U1948 (N_1948,In_1227,In_2028);
xnor U1949 (N_1949,In_345,In_275);
nand U1950 (N_1950,In_105,N_70);
nor U1951 (N_1951,N_991,N_355);
nor U1952 (N_1952,N_66,In_397);
nand U1953 (N_1953,N_191,In_2603);
nor U1954 (N_1954,In_579,In_1774);
or U1955 (N_1955,In_819,N_473);
nand U1956 (N_1956,N_193,N_231);
xor U1957 (N_1957,N_149,In_1352);
xor U1958 (N_1958,N_266,N_386);
nor U1959 (N_1959,N_859,In_1391);
xnor U1960 (N_1960,In_2043,N_777);
and U1961 (N_1961,In_2570,N_895);
or U1962 (N_1962,N_934,N_200);
and U1963 (N_1963,N_907,In_2216);
and U1964 (N_1964,In_2361,N_297);
nor U1965 (N_1965,In_347,In_2927);
xnor U1966 (N_1966,N_789,In_2758);
nand U1967 (N_1967,In_2935,In_2423);
nor U1968 (N_1968,N_541,In_1791);
or U1969 (N_1969,N_308,N_622);
nor U1970 (N_1970,N_114,In_2775);
xor U1971 (N_1971,In_2610,N_383);
xor U1972 (N_1972,N_809,N_152);
and U1973 (N_1973,In_737,In_765);
and U1974 (N_1974,N_734,N_593);
or U1975 (N_1975,N_955,In_2207);
or U1976 (N_1976,In_636,In_1561);
nor U1977 (N_1977,In_1545,In_2394);
nand U1978 (N_1978,In_1914,In_2095);
or U1979 (N_1979,In_2988,N_594);
and U1980 (N_1980,In_382,In_1287);
and U1981 (N_1981,In_2604,In_601);
nand U1982 (N_1982,N_362,In_1128);
nor U1983 (N_1983,N_272,N_910);
or U1984 (N_1984,N_587,In_2704);
xnor U1985 (N_1985,N_797,N_100);
and U1986 (N_1986,N_954,N_967);
or U1987 (N_1987,In_491,N_294);
nor U1988 (N_1988,N_509,N_505);
and U1989 (N_1989,N_506,N_878);
nand U1990 (N_1990,In_1714,In_1036);
and U1991 (N_1991,In_2650,N_47);
and U1992 (N_1992,N_320,In_1024);
nand U1993 (N_1993,In_1251,N_673);
nor U1994 (N_1994,N_980,N_573);
nand U1995 (N_1995,In_1133,In_1199);
nand U1996 (N_1996,In_1836,N_39);
nand U1997 (N_1997,In_2813,N_450);
and U1998 (N_1998,N_705,N_43);
xor U1999 (N_1999,In_600,In_1379);
nand U2000 (N_2000,N_1829,N_1533);
and U2001 (N_2001,N_1292,N_1118);
nand U2002 (N_2002,N_1468,N_1095);
nor U2003 (N_2003,N_1338,N_1859);
nand U2004 (N_2004,N_1394,N_1728);
xnor U2005 (N_2005,N_1400,N_1293);
or U2006 (N_2006,N_1390,N_1249);
or U2007 (N_2007,N_1510,N_1992);
and U2008 (N_2008,N_1818,N_1705);
nand U2009 (N_2009,N_1697,N_1792);
xnor U2010 (N_2010,N_1704,N_1326);
xnor U2011 (N_2011,N_1513,N_1968);
xnor U2012 (N_2012,N_1226,N_1843);
and U2013 (N_2013,N_1813,N_1879);
nand U2014 (N_2014,N_1469,N_1880);
or U2015 (N_2015,N_1679,N_1972);
nor U2016 (N_2016,N_1442,N_1606);
xor U2017 (N_2017,N_1447,N_1602);
nor U2018 (N_2018,N_1096,N_1785);
nor U2019 (N_2019,N_1842,N_1558);
xor U2020 (N_2020,N_1406,N_1170);
xnor U2021 (N_2021,N_1472,N_1335);
or U2022 (N_2022,N_1799,N_1932);
or U2023 (N_2023,N_1074,N_1159);
xor U2024 (N_2024,N_1482,N_1666);
nor U2025 (N_2025,N_1862,N_1171);
or U2026 (N_2026,N_1929,N_1795);
nand U2027 (N_2027,N_1612,N_1939);
or U2028 (N_2028,N_1512,N_1619);
and U2029 (N_2029,N_1828,N_1933);
nor U2030 (N_2030,N_1415,N_1242);
nand U2031 (N_2031,N_1057,N_1032);
nand U2032 (N_2032,N_1494,N_1375);
xnor U2033 (N_2033,N_1451,N_1459);
nand U2034 (N_2034,N_1322,N_1524);
nand U2035 (N_2035,N_1886,N_1092);
or U2036 (N_2036,N_1868,N_1700);
nand U2037 (N_2037,N_1580,N_1274);
and U2038 (N_2038,N_1324,N_1884);
nand U2039 (N_2039,N_1617,N_1013);
nand U2040 (N_2040,N_1568,N_1804);
xnor U2041 (N_2041,N_1291,N_1232);
nand U2042 (N_2042,N_1867,N_1976);
xnor U2043 (N_2043,N_1890,N_1934);
or U2044 (N_2044,N_1045,N_1178);
nor U2045 (N_2045,N_1647,N_1626);
or U2046 (N_2046,N_1332,N_1997);
nor U2047 (N_2047,N_1334,N_1812);
nand U2048 (N_2048,N_1416,N_1098);
and U2049 (N_2049,N_1002,N_1120);
and U2050 (N_2050,N_1686,N_1424);
xor U2051 (N_2051,N_1085,N_1805);
xnor U2052 (N_2052,N_1033,N_1019);
xnor U2053 (N_2053,N_1764,N_1486);
or U2054 (N_2054,N_1729,N_1191);
nor U2055 (N_2055,N_1581,N_1759);
nor U2056 (N_2056,N_1803,N_1056);
and U2057 (N_2057,N_1866,N_1417);
xor U2058 (N_2058,N_1778,N_1353);
or U2059 (N_2059,N_1201,N_1632);
nor U2060 (N_2060,N_1681,N_1461);
and U2061 (N_2061,N_1789,N_1498);
or U2062 (N_2062,N_1597,N_1410);
or U2063 (N_2063,N_1656,N_1991);
or U2064 (N_2064,N_1959,N_1102);
nand U2065 (N_2065,N_1490,N_1044);
nor U2066 (N_2066,N_1702,N_1426);
nand U2067 (N_2067,N_1064,N_1714);
nand U2068 (N_2068,N_1907,N_1673);
xnor U2069 (N_2069,N_1450,N_1217);
nor U2070 (N_2070,N_1346,N_1207);
or U2071 (N_2071,N_1475,N_1430);
nand U2072 (N_2072,N_1245,N_1589);
or U2073 (N_2073,N_1137,N_1248);
nor U2074 (N_2074,N_1832,N_1642);
and U2075 (N_2075,N_1822,N_1199);
nand U2076 (N_2076,N_1631,N_1331);
or U2077 (N_2077,N_1108,N_1132);
and U2078 (N_2078,N_1979,N_1358);
nand U2079 (N_2079,N_1749,N_1628);
nand U2080 (N_2080,N_1618,N_1550);
xnor U2081 (N_2081,N_1620,N_1029);
nor U2082 (N_2082,N_1635,N_1360);
xor U2083 (N_2083,N_1005,N_1600);
and U2084 (N_2084,N_1241,N_1624);
xor U2085 (N_2085,N_1196,N_1927);
nand U2086 (N_2086,N_1103,N_1831);
nor U2087 (N_2087,N_1562,N_1398);
xor U2088 (N_2088,N_1149,N_1348);
and U2089 (N_2089,N_1182,N_1753);
or U2090 (N_2090,N_1369,N_1680);
xor U2091 (N_2091,N_1297,N_1088);
nand U2092 (N_2092,N_1903,N_1347);
nor U2093 (N_2093,N_1918,N_1720);
nand U2094 (N_2094,N_1777,N_1576);
and U2095 (N_2095,N_1961,N_1039);
nor U2096 (N_2096,N_1001,N_1971);
or U2097 (N_2097,N_1990,N_1474);
xnor U2098 (N_2098,N_1925,N_1615);
nor U2099 (N_2099,N_1891,N_1769);
nor U2100 (N_2100,N_1657,N_1139);
and U2101 (N_2101,N_1214,N_1622);
nor U2102 (N_2102,N_1167,N_1821);
and U2103 (N_2103,N_1689,N_1330);
and U2104 (N_2104,N_1372,N_1945);
xor U2105 (N_2105,N_1501,N_1713);
nand U2106 (N_2106,N_1252,N_1380);
and U2107 (N_2107,N_1844,N_1011);
or U2108 (N_2108,N_1819,N_1758);
nand U2109 (N_2109,N_1141,N_1955);
xor U2110 (N_2110,N_1770,N_1889);
or U2111 (N_2111,N_1411,N_1559);
nor U2112 (N_2112,N_1185,N_1190);
xnor U2113 (N_2113,N_1838,N_1731);
nand U2114 (N_2114,N_1847,N_1757);
or U2115 (N_2115,N_1532,N_1640);
nand U2116 (N_2116,N_1594,N_1601);
or U2117 (N_2117,N_1458,N_1113);
nand U2118 (N_2118,N_1549,N_1671);
and U2119 (N_2119,N_1609,N_1476);
xor U2120 (N_2120,N_1554,N_1244);
nor U2121 (N_2121,N_1412,N_1523);
xor U2122 (N_2122,N_1385,N_1957);
and U2123 (N_2123,N_1370,N_1392);
xor U2124 (N_2124,N_1089,N_1026);
xor U2125 (N_2125,N_1556,N_1439);
nand U2126 (N_2126,N_1783,N_1179);
and U2127 (N_2127,N_1897,N_1161);
nor U2128 (N_2128,N_1920,N_1023);
and U2129 (N_2129,N_1900,N_1634);
nor U2130 (N_2130,N_1467,N_1522);
or U2131 (N_2131,N_1854,N_1973);
or U2132 (N_2132,N_1999,N_1623);
and U2133 (N_2133,N_1489,N_1809);
nand U2134 (N_2134,N_1151,N_1455);
or U2135 (N_2135,N_1893,N_1371);
xor U2136 (N_2136,N_1786,N_1200);
nor U2137 (N_2137,N_1464,N_1740);
and U2138 (N_2138,N_1124,N_1446);
and U2139 (N_2139,N_1708,N_1100);
xor U2140 (N_2140,N_1440,N_1717);
or U2141 (N_2141,N_1130,N_1760);
and U2142 (N_2142,N_1342,N_1691);
nor U2143 (N_2143,N_1156,N_1833);
nor U2144 (N_2144,N_1284,N_1329);
and U2145 (N_2145,N_1846,N_1008);
nand U2146 (N_2146,N_1655,N_1716);
nor U2147 (N_2147,N_1443,N_1354);
xor U2148 (N_2148,N_1077,N_1881);
nand U2149 (N_2149,N_1418,N_1213);
xor U2150 (N_2150,N_1505,N_1734);
nor U2151 (N_2151,N_1935,N_1824);
or U2152 (N_2152,N_1566,N_1452);
and U2153 (N_2153,N_1107,N_1014);
and U2154 (N_2154,N_1176,N_1998);
or U2155 (N_2155,N_1035,N_1208);
nor U2156 (N_2156,N_1825,N_1855);
and U2157 (N_2157,N_1240,N_1802);
nor U2158 (N_2158,N_1873,N_1362);
or U2159 (N_2159,N_1021,N_1896);
nand U2160 (N_2160,N_1851,N_1793);
or U2161 (N_2161,N_1962,N_1563);
or U2162 (N_2162,N_1738,N_1682);
or U2163 (N_2163,N_1956,N_1826);
and U2164 (N_2164,N_1377,N_1283);
xor U2165 (N_2165,N_1944,N_1947);
nand U2166 (N_2166,N_1718,N_1471);
nand U2167 (N_2167,N_1491,N_1794);
or U2168 (N_2168,N_1857,N_1441);
nand U2169 (N_2169,N_1904,N_1987);
or U2170 (N_2170,N_1257,N_1036);
nand U2171 (N_2171,N_1169,N_1106);
nand U2172 (N_2172,N_1662,N_1517);
xnor U2173 (N_2173,N_1020,N_1365);
and U2174 (N_2174,N_1871,N_1314);
and U2175 (N_2175,N_1911,N_1894);
nand U2176 (N_2176,N_1616,N_1025);
and U2177 (N_2177,N_1389,N_1808);
or U2178 (N_2178,N_1310,N_1285);
and U2179 (N_2179,N_1397,N_1496);
nand U2180 (N_2180,N_1269,N_1004);
or U2181 (N_2181,N_1433,N_1906);
nand U2182 (N_2182,N_1395,N_1122);
and U2183 (N_2183,N_1943,N_1967);
and U2184 (N_2184,N_1684,N_1305);
nand U2185 (N_2185,N_1951,N_1311);
nand U2186 (N_2186,N_1247,N_1255);
or U2187 (N_2187,N_1018,N_1267);
or U2188 (N_2188,N_1937,N_1277);
nor U2189 (N_2189,N_1983,N_1688);
xnor U2190 (N_2190,N_1773,N_1931);
or U2191 (N_2191,N_1270,N_1084);
nand U2192 (N_2192,N_1963,N_1827);
nor U2193 (N_2193,N_1781,N_1080);
and U2194 (N_2194,N_1123,N_1586);
nor U2195 (N_2195,N_1670,N_1638);
and U2196 (N_2196,N_1858,N_1076);
or U2197 (N_2197,N_1922,N_1564);
and U2198 (N_2198,N_1253,N_1614);
or U2199 (N_2199,N_1633,N_1230);
nor U2200 (N_2200,N_1519,N_1239);
nor U2201 (N_2201,N_1340,N_1970);
or U2202 (N_2202,N_1384,N_1940);
nor U2203 (N_2203,N_1645,N_1093);
and U2204 (N_2204,N_1062,N_1402);
xor U2205 (N_2205,N_1470,N_1869);
nor U2206 (N_2206,N_1352,N_1981);
or U2207 (N_2207,N_1229,N_1912);
xnor U2208 (N_2208,N_1184,N_1328);
or U2209 (N_2209,N_1861,N_1082);
nand U2210 (N_2210,N_1478,N_1115);
nand U2211 (N_2211,N_1155,N_1220);
or U2212 (N_2212,N_1423,N_1078);
nand U2213 (N_2213,N_1675,N_1150);
or U2214 (N_2214,N_1099,N_1480);
or U2215 (N_2215,N_1094,N_1752);
xor U2216 (N_2216,N_1946,N_1425);
or U2217 (N_2217,N_1473,N_1058);
or U2218 (N_2218,N_1853,N_1488);
and U2219 (N_2219,N_1665,N_1776);
and U2220 (N_2220,N_1678,N_1706);
xnor U2221 (N_2221,N_1457,N_1361);
nor U2222 (N_2222,N_1047,N_1690);
and U2223 (N_2223,N_1500,N_1485);
xor U2224 (N_2224,N_1661,N_1952);
nor U2225 (N_2225,N_1901,N_1303);
nand U2226 (N_2226,N_1404,N_1327);
or U2227 (N_2227,N_1263,N_1028);
and U2228 (N_2228,N_1349,N_1031);
nor U2229 (N_2229,N_1111,N_1766);
and U2230 (N_2230,N_1836,N_1131);
nor U2231 (N_2231,N_1069,N_1212);
and U2232 (N_2232,N_1754,N_1243);
nor U2233 (N_2233,N_1965,N_1216);
or U2234 (N_2234,N_1436,N_1745);
xor U2235 (N_2235,N_1579,N_1477);
nor U2236 (N_2236,N_1646,N_1453);
xnor U2237 (N_2237,N_1739,N_1350);
and U2238 (N_2238,N_1189,N_1038);
nand U2239 (N_2239,N_1712,N_1321);
and U2240 (N_2240,N_1636,N_1978);
nand U2241 (N_2241,N_1109,N_1726);
nor U2242 (N_2242,N_1767,N_1166);
nor U2243 (N_2243,N_1839,N_1165);
nand U2244 (N_2244,N_1403,N_1698);
nand U2245 (N_2245,N_1641,N_1723);
xnor U2246 (N_2246,N_1386,N_1654);
nor U2247 (N_2247,N_1629,N_1810);
nand U2248 (N_2248,N_1279,N_1336);
nand U2249 (N_2249,N_1333,N_1231);
and U2250 (N_2250,N_1408,N_1246);
nand U2251 (N_2251,N_1650,N_1787);
or U2252 (N_2252,N_1233,N_1570);
nor U2253 (N_2253,N_1543,N_1393);
and U2254 (N_2254,N_1068,N_1692);
xnor U2255 (N_2255,N_1652,N_1071);
or U2256 (N_2256,N_1223,N_1125);
nor U2257 (N_2257,N_1954,N_1902);
nand U2258 (N_2258,N_1016,N_1514);
or U2259 (N_2259,N_1308,N_1133);
and U2260 (N_2260,N_1449,N_1663);
and U2261 (N_2261,N_1721,N_1814);
nand U2262 (N_2262,N_1750,N_1966);
nor U2263 (N_2263,N_1495,N_1275);
or U2264 (N_2264,N_1256,N_1224);
or U2265 (N_2265,N_1409,N_1807);
nand U2266 (N_2266,N_1806,N_1788);
xor U2267 (N_2267,N_1237,N_1582);
or U2268 (N_2268,N_1126,N_1320);
or U2269 (N_2269,N_1528,N_1590);
xor U2270 (N_2270,N_1290,N_1266);
nand U2271 (N_2271,N_1864,N_1537);
or U2272 (N_2272,N_1709,N_1438);
xor U2273 (N_2273,N_1083,N_1059);
and U2274 (N_2274,N_1525,N_1572);
and U2275 (N_2275,N_1079,N_1427);
and U2276 (N_2276,N_1748,N_1565);
and U2277 (N_2277,N_1577,N_1435);
nor U2278 (N_2278,N_1157,N_1129);
xnor U2279 (N_2279,N_1984,N_1262);
nand U2280 (N_2280,N_1209,N_1168);
xor U2281 (N_2281,N_1306,N_1027);
and U2282 (N_2282,N_1276,N_1669);
nand U2283 (N_2283,N_1228,N_1382);
and U2284 (N_2284,N_1660,N_1264);
and U2285 (N_2285,N_1504,N_1527);
or U2286 (N_2286,N_1067,N_1363);
nand U2287 (N_2287,N_1101,N_1701);
xor U2288 (N_2288,N_1289,N_1399);
xor U2289 (N_2289,N_1696,N_1298);
nand U2290 (N_2290,N_1188,N_1312);
nand U2291 (N_2291,N_1598,N_1508);
nor U2292 (N_2292,N_1388,N_1996);
or U2293 (N_2293,N_1466,N_1172);
nor U2294 (N_2294,N_1849,N_1053);
nor U2295 (N_2295,N_1711,N_1227);
or U2296 (N_2296,N_1075,N_1300);
and U2297 (N_2297,N_1260,N_1599);
and U2298 (N_2298,N_1569,N_1722);
nor U2299 (N_2299,N_1315,N_1936);
or U2300 (N_2300,N_1542,N_1186);
xnor U2301 (N_2301,N_1539,N_1000);
nor U2302 (N_2302,N_1921,N_1593);
xor U2303 (N_2303,N_1481,N_1552);
nand U2304 (N_2304,N_1516,N_1359);
and U2305 (N_2305,N_1462,N_1982);
nand U2306 (N_2306,N_1281,N_1204);
nand U2307 (N_2307,N_1800,N_1090);
xor U2308 (N_2308,N_1658,N_1719);
and U2309 (N_2309,N_1117,N_1948);
nand U2310 (N_2310,N_1041,N_1378);
or U2311 (N_2311,N_1148,N_1070);
xnor U2312 (N_2312,N_1175,N_1487);
and U2313 (N_2313,N_1977,N_1782);
and U2314 (N_2314,N_1885,N_1715);
nor U2315 (N_2315,N_1737,N_1643);
and U2316 (N_2316,N_1309,N_1603);
nand U2317 (N_2317,N_1648,N_1621);
xnor U2318 (N_2318,N_1725,N_1339);
and U2319 (N_2319,N_1584,N_1206);
nand U2320 (N_2320,N_1009,N_1520);
and U2321 (N_2321,N_1351,N_1762);
nand U2322 (N_2322,N_1790,N_1448);
nor U2323 (N_2323,N_1273,N_1343);
and U2324 (N_2324,N_1138,N_1499);
and U2325 (N_2325,N_1429,N_1664);
or U2326 (N_2326,N_1373,N_1742);
nor U2327 (N_2327,N_1541,N_1153);
xor U2328 (N_2328,N_1693,N_1659);
xor U2329 (N_2329,N_1205,N_1234);
nor U2330 (N_2330,N_1540,N_1272);
nor U2331 (N_2331,N_1366,N_1526);
and U2332 (N_2332,N_1548,N_1639);
and U2333 (N_2333,N_1432,N_1140);
and U2334 (N_2334,N_1765,N_1147);
nand U2335 (N_2335,N_1192,N_1143);
nand U2336 (N_2336,N_1695,N_1958);
xor U2337 (N_2337,N_1780,N_1667);
nand U2338 (N_2338,N_1048,N_1942);
xor U2339 (N_2339,N_1325,N_1699);
and U2340 (N_2340,N_1022,N_1483);
nand U2341 (N_2341,N_1465,N_1054);
nand U2342 (N_2342,N_1183,N_1401);
nor U2343 (N_2343,N_1534,N_1225);
and U2344 (N_2344,N_1114,N_1086);
nand U2345 (N_2345,N_1924,N_1596);
or U2346 (N_2346,N_1674,N_1863);
nor U2347 (N_2347,N_1050,N_1685);
nor U2348 (N_2348,N_1817,N_1898);
xor U2349 (N_2349,N_1034,N_1374);
and U2350 (N_2350,N_1105,N_1007);
nand U2351 (N_2351,N_1875,N_1964);
xnor U2352 (N_2352,N_1091,N_1278);
nand U2353 (N_2353,N_1730,N_1953);
nand U2354 (N_2354,N_1870,N_1164);
xor U2355 (N_2355,N_1974,N_1052);
xor U2356 (N_2356,N_1538,N_1733);
and U2357 (N_2357,N_1222,N_1040);
nor U2358 (N_2358,N_1060,N_1683);
and U2359 (N_2359,N_1259,N_1042);
nor U2360 (N_2360,N_1081,N_1914);
and U2361 (N_2361,N_1142,N_1518);
xor U2362 (N_2362,N_1756,N_1915);
and U2363 (N_2363,N_1506,N_1061);
or U2364 (N_2364,N_1128,N_1774);
or U2365 (N_2365,N_1637,N_1319);
nor U2366 (N_2366,N_1145,N_1567);
and U2367 (N_2367,N_1801,N_1649);
xor U2368 (N_2368,N_1364,N_1055);
xor U2369 (N_2369,N_1895,N_1152);
or U2370 (N_2370,N_1823,N_1530);
nand U2371 (N_2371,N_1271,N_1816);
or U2372 (N_2372,N_1743,N_1553);
nand U2373 (N_2373,N_1775,N_1280);
nand U2374 (N_2374,N_1454,N_1980);
and U2375 (N_2375,N_1006,N_1509);
and U2376 (N_2376,N_1841,N_1511);
and U2377 (N_2377,N_1046,N_1174);
nor U2378 (N_2378,N_1317,N_1419);
nor U2379 (N_2379,N_1295,N_1507);
nor U2380 (N_2380,N_1771,N_1941);
nand U2381 (N_2381,N_1445,N_1356);
nand U2382 (N_2382,N_1261,N_1888);
nand U2383 (N_2383,N_1268,N_1710);
xor U2384 (N_2384,N_1994,N_1547);
or U2385 (N_2385,N_1557,N_1063);
nand U2386 (N_2386,N_1238,N_1988);
nor U2387 (N_2387,N_1677,N_1065);
nor U2388 (N_2388,N_1848,N_1917);
nand U2389 (N_2389,N_1573,N_1908);
nand U2390 (N_2390,N_1136,N_1405);
nor U2391 (N_2391,N_1950,N_1479);
nor U2392 (N_2392,N_1187,N_1421);
xnor U2393 (N_2393,N_1845,N_1529);
xnor U2394 (N_2394,N_1049,N_1724);
xor U2395 (N_2395,N_1177,N_1413);
or U2396 (N_2396,N_1236,N_1625);
nor U2397 (N_2397,N_1344,N_1521);
nor U2398 (N_2398,N_1012,N_1544);
nand U2399 (N_2399,N_1611,N_1254);
or U2400 (N_2400,N_1337,N_1747);
nor U2401 (N_2401,N_1892,N_1073);
and U2402 (N_2402,N_1872,N_1928);
or U2403 (N_2403,N_1850,N_1592);
and U2404 (N_2404,N_1546,N_1923);
or U2405 (N_2405,N_1751,N_1840);
and U2406 (N_2406,N_1995,N_1503);
and U2407 (N_2407,N_1672,N_1288);
and U2408 (N_2408,N_1037,N_1555);
nand U2409 (N_2409,N_1112,N_1736);
or U2410 (N_2410,N_1811,N_1969);
or U2411 (N_2411,N_1135,N_1194);
nor U2412 (N_2412,N_1856,N_1318);
or U2413 (N_2413,N_1024,N_1163);
or U2414 (N_2414,N_1820,N_1497);
xor U2415 (N_2415,N_1414,N_1574);
nor U2416 (N_2416,N_1938,N_1197);
and U2417 (N_2417,N_1345,N_1583);
or U2418 (N_2418,N_1119,N_1087);
nand U2419 (N_2419,N_1407,N_1707);
and U2420 (N_2420,N_1154,N_1926);
nor U2421 (N_2421,N_1313,N_1798);
xor U2422 (N_2422,N_1993,N_1909);
or U2423 (N_2423,N_1561,N_1250);
nand U2424 (N_2424,N_1422,N_1651);
xnor U2425 (N_2425,N_1545,N_1746);
nand U2426 (N_2426,N_1551,N_1431);
nand U2427 (N_2427,N_1930,N_1387);
nand U2428 (N_2428,N_1381,N_1755);
nor U2429 (N_2429,N_1668,N_1986);
and U2430 (N_2430,N_1210,N_1376);
and U2431 (N_2431,N_1379,N_1605);
and U2432 (N_2432,N_1905,N_1134);
nor U2433 (N_2433,N_1301,N_1607);
nand U2434 (N_2434,N_1072,N_1535);
nor U2435 (N_2435,N_1910,N_1296);
and U2436 (N_2436,N_1304,N_1251);
or U2437 (N_2437,N_1097,N_1396);
nand U2438 (N_2438,N_1127,N_1727);
xor U2439 (N_2439,N_1146,N_1578);
or U2440 (N_2440,N_1536,N_1830);
xnor U2441 (N_2441,N_1193,N_1768);
nor U2442 (N_2442,N_1796,N_1608);
nor U2443 (N_2443,N_1591,N_1181);
and U2444 (N_2444,N_1420,N_1815);
xnor U2445 (N_2445,N_1158,N_1919);
nand U2446 (N_2446,N_1218,N_1694);
nand U2447 (N_2447,N_1687,N_1860);
or U2448 (N_2448,N_1460,N_1610);
and U2449 (N_2449,N_1916,N_1355);
and U2450 (N_2450,N_1066,N_1307);
nand U2451 (N_2451,N_1030,N_1463);
or U2452 (N_2452,N_1874,N_1434);
nor U2453 (N_2453,N_1852,N_1835);
or U2454 (N_2454,N_1630,N_1258);
and U2455 (N_2455,N_1732,N_1913);
or U2456 (N_2456,N_1121,N_1949);
xor U2457 (N_2457,N_1878,N_1221);
nand U2458 (N_2458,N_1585,N_1287);
xnor U2459 (N_2459,N_1160,N_1613);
or U2460 (N_2460,N_1735,N_1575);
or U2461 (N_2461,N_1791,N_1883);
and U2462 (N_2462,N_1162,N_1865);
or U2463 (N_2463,N_1316,N_1195);
and U2464 (N_2464,N_1010,N_1899);
nand U2465 (N_2465,N_1456,N_1104);
or U2466 (N_2466,N_1975,N_1703);
and U2467 (N_2467,N_1173,N_1235);
nand U2468 (N_2468,N_1587,N_1302);
or U2469 (N_2469,N_1588,N_1772);
nand U2470 (N_2470,N_1110,N_1779);
and U2471 (N_2471,N_1391,N_1211);
or U2472 (N_2472,N_1887,N_1219);
and U2473 (N_2473,N_1595,N_1203);
or U2474 (N_2474,N_1367,N_1017);
or U2475 (N_2475,N_1627,N_1323);
or U2476 (N_2476,N_1877,N_1202);
nand U2477 (N_2477,N_1653,N_1571);
nand U2478 (N_2478,N_1560,N_1744);
and U2479 (N_2479,N_1341,N_1444);
or U2480 (N_2480,N_1357,N_1198);
nor U2481 (N_2481,N_1144,N_1985);
xnor U2482 (N_2482,N_1299,N_1882);
nor U2483 (N_2483,N_1180,N_1876);
xor U2484 (N_2484,N_1437,N_1834);
nand U2485 (N_2485,N_1741,N_1837);
or U2486 (N_2486,N_1531,N_1294);
or U2487 (N_2487,N_1116,N_1784);
nand U2488 (N_2488,N_1797,N_1644);
nor U2489 (N_2489,N_1502,N_1763);
and U2490 (N_2490,N_1282,N_1484);
or U2491 (N_2491,N_1383,N_1989);
nor U2492 (N_2492,N_1043,N_1515);
nor U2493 (N_2493,N_1493,N_1604);
xnor U2494 (N_2494,N_1960,N_1286);
or U2495 (N_2495,N_1265,N_1676);
or U2496 (N_2496,N_1492,N_1015);
nand U2497 (N_2497,N_1215,N_1368);
nor U2498 (N_2498,N_1761,N_1003);
and U2499 (N_2499,N_1428,N_1051);
nor U2500 (N_2500,N_1288,N_1528);
nor U2501 (N_2501,N_1613,N_1044);
nand U2502 (N_2502,N_1722,N_1392);
nand U2503 (N_2503,N_1455,N_1233);
nor U2504 (N_2504,N_1989,N_1156);
nand U2505 (N_2505,N_1726,N_1207);
and U2506 (N_2506,N_1907,N_1919);
nor U2507 (N_2507,N_1120,N_1477);
nand U2508 (N_2508,N_1510,N_1840);
nor U2509 (N_2509,N_1307,N_1773);
and U2510 (N_2510,N_1635,N_1717);
or U2511 (N_2511,N_1083,N_1555);
nand U2512 (N_2512,N_1186,N_1260);
nand U2513 (N_2513,N_1670,N_1888);
or U2514 (N_2514,N_1897,N_1267);
nand U2515 (N_2515,N_1267,N_1785);
and U2516 (N_2516,N_1907,N_1741);
nor U2517 (N_2517,N_1407,N_1035);
or U2518 (N_2518,N_1631,N_1367);
nand U2519 (N_2519,N_1293,N_1470);
xor U2520 (N_2520,N_1797,N_1286);
or U2521 (N_2521,N_1037,N_1532);
nand U2522 (N_2522,N_1498,N_1602);
and U2523 (N_2523,N_1302,N_1498);
nor U2524 (N_2524,N_1720,N_1517);
and U2525 (N_2525,N_1306,N_1924);
nand U2526 (N_2526,N_1980,N_1399);
nor U2527 (N_2527,N_1451,N_1525);
and U2528 (N_2528,N_1103,N_1947);
nand U2529 (N_2529,N_1708,N_1995);
nand U2530 (N_2530,N_1786,N_1783);
nor U2531 (N_2531,N_1490,N_1061);
xnor U2532 (N_2532,N_1810,N_1635);
nor U2533 (N_2533,N_1153,N_1155);
or U2534 (N_2534,N_1725,N_1675);
and U2535 (N_2535,N_1536,N_1434);
xnor U2536 (N_2536,N_1743,N_1834);
and U2537 (N_2537,N_1811,N_1292);
xnor U2538 (N_2538,N_1789,N_1640);
or U2539 (N_2539,N_1856,N_1099);
or U2540 (N_2540,N_1302,N_1992);
nand U2541 (N_2541,N_1232,N_1260);
nor U2542 (N_2542,N_1233,N_1978);
nand U2543 (N_2543,N_1726,N_1561);
xor U2544 (N_2544,N_1249,N_1403);
nor U2545 (N_2545,N_1146,N_1520);
xor U2546 (N_2546,N_1856,N_1800);
nor U2547 (N_2547,N_1436,N_1947);
xnor U2548 (N_2548,N_1139,N_1983);
and U2549 (N_2549,N_1841,N_1455);
or U2550 (N_2550,N_1043,N_1008);
xor U2551 (N_2551,N_1705,N_1070);
nand U2552 (N_2552,N_1705,N_1123);
nand U2553 (N_2553,N_1722,N_1439);
nand U2554 (N_2554,N_1112,N_1673);
xor U2555 (N_2555,N_1624,N_1306);
and U2556 (N_2556,N_1025,N_1950);
xnor U2557 (N_2557,N_1648,N_1614);
and U2558 (N_2558,N_1813,N_1051);
xnor U2559 (N_2559,N_1406,N_1619);
or U2560 (N_2560,N_1470,N_1691);
nand U2561 (N_2561,N_1582,N_1786);
xor U2562 (N_2562,N_1026,N_1857);
and U2563 (N_2563,N_1562,N_1809);
nor U2564 (N_2564,N_1134,N_1061);
nor U2565 (N_2565,N_1794,N_1571);
and U2566 (N_2566,N_1732,N_1048);
and U2567 (N_2567,N_1797,N_1854);
xor U2568 (N_2568,N_1538,N_1179);
nand U2569 (N_2569,N_1220,N_1647);
xnor U2570 (N_2570,N_1201,N_1457);
nand U2571 (N_2571,N_1551,N_1416);
and U2572 (N_2572,N_1231,N_1644);
xnor U2573 (N_2573,N_1927,N_1276);
xor U2574 (N_2574,N_1059,N_1249);
and U2575 (N_2575,N_1984,N_1162);
nor U2576 (N_2576,N_1097,N_1432);
nand U2577 (N_2577,N_1023,N_1058);
and U2578 (N_2578,N_1690,N_1651);
xnor U2579 (N_2579,N_1836,N_1700);
and U2580 (N_2580,N_1275,N_1795);
xnor U2581 (N_2581,N_1314,N_1055);
nand U2582 (N_2582,N_1645,N_1859);
nor U2583 (N_2583,N_1123,N_1089);
nand U2584 (N_2584,N_1753,N_1180);
nand U2585 (N_2585,N_1920,N_1758);
or U2586 (N_2586,N_1357,N_1916);
nor U2587 (N_2587,N_1720,N_1705);
nand U2588 (N_2588,N_1545,N_1990);
or U2589 (N_2589,N_1775,N_1842);
nand U2590 (N_2590,N_1112,N_1511);
nor U2591 (N_2591,N_1400,N_1746);
nand U2592 (N_2592,N_1856,N_1730);
xnor U2593 (N_2593,N_1731,N_1069);
nand U2594 (N_2594,N_1770,N_1048);
nand U2595 (N_2595,N_1927,N_1751);
and U2596 (N_2596,N_1590,N_1599);
nor U2597 (N_2597,N_1568,N_1093);
nor U2598 (N_2598,N_1710,N_1488);
or U2599 (N_2599,N_1772,N_1009);
or U2600 (N_2600,N_1692,N_1425);
nor U2601 (N_2601,N_1021,N_1479);
xnor U2602 (N_2602,N_1783,N_1437);
and U2603 (N_2603,N_1421,N_1837);
or U2604 (N_2604,N_1972,N_1186);
or U2605 (N_2605,N_1778,N_1774);
xor U2606 (N_2606,N_1240,N_1612);
or U2607 (N_2607,N_1168,N_1592);
nand U2608 (N_2608,N_1439,N_1451);
xor U2609 (N_2609,N_1662,N_1478);
nor U2610 (N_2610,N_1488,N_1991);
and U2611 (N_2611,N_1986,N_1372);
nand U2612 (N_2612,N_1536,N_1543);
nor U2613 (N_2613,N_1789,N_1991);
xor U2614 (N_2614,N_1679,N_1492);
nor U2615 (N_2615,N_1780,N_1611);
nor U2616 (N_2616,N_1542,N_1316);
and U2617 (N_2617,N_1269,N_1106);
or U2618 (N_2618,N_1397,N_1061);
and U2619 (N_2619,N_1448,N_1742);
and U2620 (N_2620,N_1349,N_1821);
and U2621 (N_2621,N_1721,N_1786);
or U2622 (N_2622,N_1380,N_1619);
or U2623 (N_2623,N_1621,N_1855);
and U2624 (N_2624,N_1924,N_1920);
and U2625 (N_2625,N_1344,N_1704);
xnor U2626 (N_2626,N_1199,N_1338);
and U2627 (N_2627,N_1907,N_1019);
and U2628 (N_2628,N_1318,N_1257);
xnor U2629 (N_2629,N_1793,N_1231);
nand U2630 (N_2630,N_1692,N_1820);
nand U2631 (N_2631,N_1372,N_1310);
or U2632 (N_2632,N_1858,N_1303);
xnor U2633 (N_2633,N_1551,N_1390);
nor U2634 (N_2634,N_1050,N_1833);
and U2635 (N_2635,N_1134,N_1426);
and U2636 (N_2636,N_1020,N_1525);
and U2637 (N_2637,N_1235,N_1587);
xnor U2638 (N_2638,N_1788,N_1231);
nand U2639 (N_2639,N_1354,N_1636);
nor U2640 (N_2640,N_1676,N_1130);
nand U2641 (N_2641,N_1423,N_1333);
nor U2642 (N_2642,N_1002,N_1967);
nor U2643 (N_2643,N_1397,N_1734);
or U2644 (N_2644,N_1536,N_1442);
nand U2645 (N_2645,N_1050,N_1080);
or U2646 (N_2646,N_1736,N_1061);
xnor U2647 (N_2647,N_1248,N_1256);
and U2648 (N_2648,N_1113,N_1641);
xor U2649 (N_2649,N_1466,N_1631);
xor U2650 (N_2650,N_1938,N_1634);
or U2651 (N_2651,N_1442,N_1896);
xnor U2652 (N_2652,N_1212,N_1116);
xnor U2653 (N_2653,N_1194,N_1656);
or U2654 (N_2654,N_1198,N_1939);
or U2655 (N_2655,N_1598,N_1086);
and U2656 (N_2656,N_1494,N_1912);
and U2657 (N_2657,N_1095,N_1138);
xor U2658 (N_2658,N_1557,N_1437);
or U2659 (N_2659,N_1119,N_1253);
and U2660 (N_2660,N_1799,N_1675);
and U2661 (N_2661,N_1122,N_1037);
and U2662 (N_2662,N_1569,N_1801);
and U2663 (N_2663,N_1980,N_1453);
nand U2664 (N_2664,N_1319,N_1962);
xnor U2665 (N_2665,N_1271,N_1934);
nand U2666 (N_2666,N_1740,N_1809);
or U2667 (N_2667,N_1199,N_1773);
nor U2668 (N_2668,N_1000,N_1022);
xor U2669 (N_2669,N_1522,N_1449);
and U2670 (N_2670,N_1632,N_1321);
nand U2671 (N_2671,N_1965,N_1968);
and U2672 (N_2672,N_1791,N_1321);
nor U2673 (N_2673,N_1741,N_1800);
nor U2674 (N_2674,N_1444,N_1070);
xnor U2675 (N_2675,N_1661,N_1301);
and U2676 (N_2676,N_1120,N_1623);
nand U2677 (N_2677,N_1036,N_1522);
nor U2678 (N_2678,N_1177,N_1412);
nor U2679 (N_2679,N_1728,N_1528);
or U2680 (N_2680,N_1128,N_1219);
or U2681 (N_2681,N_1946,N_1749);
nor U2682 (N_2682,N_1226,N_1196);
or U2683 (N_2683,N_1808,N_1983);
nor U2684 (N_2684,N_1912,N_1353);
xnor U2685 (N_2685,N_1194,N_1677);
and U2686 (N_2686,N_1870,N_1007);
xnor U2687 (N_2687,N_1940,N_1392);
nand U2688 (N_2688,N_1240,N_1598);
and U2689 (N_2689,N_1717,N_1225);
xnor U2690 (N_2690,N_1353,N_1337);
or U2691 (N_2691,N_1293,N_1002);
xnor U2692 (N_2692,N_1775,N_1441);
nor U2693 (N_2693,N_1370,N_1147);
and U2694 (N_2694,N_1579,N_1767);
nand U2695 (N_2695,N_1412,N_1266);
or U2696 (N_2696,N_1136,N_1760);
and U2697 (N_2697,N_1608,N_1685);
and U2698 (N_2698,N_1577,N_1178);
nand U2699 (N_2699,N_1011,N_1510);
and U2700 (N_2700,N_1222,N_1481);
xor U2701 (N_2701,N_1876,N_1575);
and U2702 (N_2702,N_1736,N_1339);
and U2703 (N_2703,N_1178,N_1612);
and U2704 (N_2704,N_1887,N_1943);
and U2705 (N_2705,N_1665,N_1299);
or U2706 (N_2706,N_1866,N_1754);
nor U2707 (N_2707,N_1667,N_1945);
nand U2708 (N_2708,N_1116,N_1687);
xor U2709 (N_2709,N_1290,N_1784);
and U2710 (N_2710,N_1588,N_1864);
nand U2711 (N_2711,N_1940,N_1673);
or U2712 (N_2712,N_1866,N_1241);
xor U2713 (N_2713,N_1784,N_1677);
and U2714 (N_2714,N_1592,N_1519);
and U2715 (N_2715,N_1966,N_1352);
xnor U2716 (N_2716,N_1081,N_1370);
nor U2717 (N_2717,N_1591,N_1480);
and U2718 (N_2718,N_1400,N_1902);
or U2719 (N_2719,N_1181,N_1623);
nor U2720 (N_2720,N_1604,N_1474);
nand U2721 (N_2721,N_1621,N_1013);
nand U2722 (N_2722,N_1481,N_1354);
or U2723 (N_2723,N_1838,N_1543);
and U2724 (N_2724,N_1584,N_1658);
xor U2725 (N_2725,N_1471,N_1433);
nor U2726 (N_2726,N_1134,N_1852);
and U2727 (N_2727,N_1680,N_1755);
xor U2728 (N_2728,N_1110,N_1626);
nand U2729 (N_2729,N_1631,N_1609);
or U2730 (N_2730,N_1330,N_1385);
and U2731 (N_2731,N_1441,N_1853);
xor U2732 (N_2732,N_1389,N_1149);
or U2733 (N_2733,N_1872,N_1561);
nand U2734 (N_2734,N_1023,N_1145);
or U2735 (N_2735,N_1114,N_1834);
nand U2736 (N_2736,N_1259,N_1142);
nor U2737 (N_2737,N_1505,N_1594);
xor U2738 (N_2738,N_1482,N_1476);
xnor U2739 (N_2739,N_1662,N_1066);
xnor U2740 (N_2740,N_1649,N_1358);
or U2741 (N_2741,N_1453,N_1527);
nor U2742 (N_2742,N_1576,N_1592);
and U2743 (N_2743,N_1300,N_1086);
nor U2744 (N_2744,N_1878,N_1666);
nor U2745 (N_2745,N_1568,N_1298);
and U2746 (N_2746,N_1244,N_1774);
nor U2747 (N_2747,N_1505,N_1421);
and U2748 (N_2748,N_1817,N_1071);
or U2749 (N_2749,N_1083,N_1598);
nand U2750 (N_2750,N_1054,N_1815);
nand U2751 (N_2751,N_1053,N_1257);
xor U2752 (N_2752,N_1234,N_1715);
xnor U2753 (N_2753,N_1175,N_1401);
nand U2754 (N_2754,N_1351,N_1675);
nor U2755 (N_2755,N_1893,N_1325);
xnor U2756 (N_2756,N_1081,N_1175);
nand U2757 (N_2757,N_1807,N_1082);
and U2758 (N_2758,N_1146,N_1756);
xnor U2759 (N_2759,N_1058,N_1576);
xnor U2760 (N_2760,N_1360,N_1128);
xnor U2761 (N_2761,N_1060,N_1777);
nor U2762 (N_2762,N_1361,N_1584);
nand U2763 (N_2763,N_1811,N_1681);
xnor U2764 (N_2764,N_1540,N_1820);
and U2765 (N_2765,N_1851,N_1862);
and U2766 (N_2766,N_1695,N_1620);
or U2767 (N_2767,N_1469,N_1856);
nand U2768 (N_2768,N_1101,N_1017);
nand U2769 (N_2769,N_1400,N_1604);
xor U2770 (N_2770,N_1579,N_1791);
xor U2771 (N_2771,N_1578,N_1144);
or U2772 (N_2772,N_1133,N_1556);
xnor U2773 (N_2773,N_1675,N_1616);
nand U2774 (N_2774,N_1196,N_1372);
and U2775 (N_2775,N_1616,N_1572);
nand U2776 (N_2776,N_1675,N_1280);
or U2777 (N_2777,N_1204,N_1695);
or U2778 (N_2778,N_1753,N_1784);
and U2779 (N_2779,N_1483,N_1642);
nor U2780 (N_2780,N_1996,N_1556);
and U2781 (N_2781,N_1272,N_1145);
and U2782 (N_2782,N_1324,N_1529);
nand U2783 (N_2783,N_1632,N_1974);
or U2784 (N_2784,N_1436,N_1377);
nand U2785 (N_2785,N_1414,N_1730);
xnor U2786 (N_2786,N_1538,N_1099);
nor U2787 (N_2787,N_1262,N_1846);
xnor U2788 (N_2788,N_1581,N_1956);
nor U2789 (N_2789,N_1338,N_1335);
nand U2790 (N_2790,N_1945,N_1063);
xor U2791 (N_2791,N_1287,N_1957);
nor U2792 (N_2792,N_1594,N_1514);
xor U2793 (N_2793,N_1560,N_1176);
nand U2794 (N_2794,N_1925,N_1915);
nor U2795 (N_2795,N_1456,N_1018);
nand U2796 (N_2796,N_1133,N_1159);
and U2797 (N_2797,N_1007,N_1207);
nor U2798 (N_2798,N_1884,N_1203);
nand U2799 (N_2799,N_1172,N_1428);
xor U2800 (N_2800,N_1365,N_1042);
or U2801 (N_2801,N_1297,N_1566);
nor U2802 (N_2802,N_1304,N_1413);
xnor U2803 (N_2803,N_1002,N_1681);
and U2804 (N_2804,N_1006,N_1159);
xor U2805 (N_2805,N_1628,N_1764);
nand U2806 (N_2806,N_1855,N_1430);
and U2807 (N_2807,N_1918,N_1707);
xor U2808 (N_2808,N_1643,N_1541);
and U2809 (N_2809,N_1482,N_1216);
and U2810 (N_2810,N_1365,N_1328);
xor U2811 (N_2811,N_1675,N_1752);
xor U2812 (N_2812,N_1358,N_1494);
xor U2813 (N_2813,N_1853,N_1344);
nor U2814 (N_2814,N_1236,N_1639);
nand U2815 (N_2815,N_1647,N_1252);
nor U2816 (N_2816,N_1886,N_1227);
xnor U2817 (N_2817,N_1977,N_1406);
nor U2818 (N_2818,N_1346,N_1671);
and U2819 (N_2819,N_1867,N_1634);
and U2820 (N_2820,N_1417,N_1796);
nor U2821 (N_2821,N_1290,N_1004);
or U2822 (N_2822,N_1727,N_1954);
nand U2823 (N_2823,N_1625,N_1538);
xor U2824 (N_2824,N_1454,N_1645);
nand U2825 (N_2825,N_1515,N_1063);
nor U2826 (N_2826,N_1141,N_1534);
nand U2827 (N_2827,N_1938,N_1581);
nand U2828 (N_2828,N_1680,N_1740);
xor U2829 (N_2829,N_1616,N_1678);
xnor U2830 (N_2830,N_1231,N_1554);
and U2831 (N_2831,N_1566,N_1900);
or U2832 (N_2832,N_1332,N_1629);
or U2833 (N_2833,N_1082,N_1503);
or U2834 (N_2834,N_1800,N_1573);
or U2835 (N_2835,N_1998,N_1806);
xor U2836 (N_2836,N_1328,N_1353);
and U2837 (N_2837,N_1289,N_1235);
nand U2838 (N_2838,N_1481,N_1850);
and U2839 (N_2839,N_1665,N_1012);
xor U2840 (N_2840,N_1667,N_1002);
or U2841 (N_2841,N_1945,N_1919);
nor U2842 (N_2842,N_1026,N_1319);
or U2843 (N_2843,N_1633,N_1348);
and U2844 (N_2844,N_1932,N_1325);
nor U2845 (N_2845,N_1190,N_1758);
xnor U2846 (N_2846,N_1011,N_1125);
or U2847 (N_2847,N_1153,N_1441);
xnor U2848 (N_2848,N_1110,N_1596);
or U2849 (N_2849,N_1610,N_1931);
and U2850 (N_2850,N_1934,N_1941);
nand U2851 (N_2851,N_1638,N_1594);
xor U2852 (N_2852,N_1472,N_1560);
xnor U2853 (N_2853,N_1071,N_1302);
or U2854 (N_2854,N_1691,N_1674);
nand U2855 (N_2855,N_1645,N_1335);
xnor U2856 (N_2856,N_1497,N_1486);
nand U2857 (N_2857,N_1575,N_1825);
or U2858 (N_2858,N_1801,N_1003);
nand U2859 (N_2859,N_1299,N_1134);
nor U2860 (N_2860,N_1097,N_1480);
or U2861 (N_2861,N_1842,N_1801);
and U2862 (N_2862,N_1344,N_1641);
xnor U2863 (N_2863,N_1400,N_1021);
or U2864 (N_2864,N_1871,N_1875);
xnor U2865 (N_2865,N_1784,N_1355);
or U2866 (N_2866,N_1336,N_1564);
nor U2867 (N_2867,N_1760,N_1671);
xnor U2868 (N_2868,N_1448,N_1598);
or U2869 (N_2869,N_1816,N_1640);
and U2870 (N_2870,N_1917,N_1858);
xnor U2871 (N_2871,N_1218,N_1697);
nand U2872 (N_2872,N_1711,N_1483);
nand U2873 (N_2873,N_1567,N_1959);
and U2874 (N_2874,N_1685,N_1070);
and U2875 (N_2875,N_1599,N_1348);
xor U2876 (N_2876,N_1150,N_1375);
nand U2877 (N_2877,N_1349,N_1502);
xnor U2878 (N_2878,N_1384,N_1072);
and U2879 (N_2879,N_1719,N_1763);
nor U2880 (N_2880,N_1435,N_1555);
nor U2881 (N_2881,N_1838,N_1604);
nand U2882 (N_2882,N_1639,N_1387);
or U2883 (N_2883,N_1375,N_1991);
nand U2884 (N_2884,N_1785,N_1544);
and U2885 (N_2885,N_1117,N_1425);
or U2886 (N_2886,N_1450,N_1555);
xnor U2887 (N_2887,N_1480,N_1182);
and U2888 (N_2888,N_1292,N_1158);
xnor U2889 (N_2889,N_1194,N_1386);
nand U2890 (N_2890,N_1254,N_1733);
nor U2891 (N_2891,N_1835,N_1634);
xnor U2892 (N_2892,N_1827,N_1701);
xor U2893 (N_2893,N_1889,N_1082);
xor U2894 (N_2894,N_1272,N_1013);
nand U2895 (N_2895,N_1494,N_1475);
nand U2896 (N_2896,N_1214,N_1352);
nor U2897 (N_2897,N_1703,N_1261);
xnor U2898 (N_2898,N_1752,N_1864);
xor U2899 (N_2899,N_1942,N_1972);
and U2900 (N_2900,N_1419,N_1981);
and U2901 (N_2901,N_1973,N_1181);
nand U2902 (N_2902,N_1688,N_1361);
and U2903 (N_2903,N_1652,N_1757);
nor U2904 (N_2904,N_1843,N_1423);
and U2905 (N_2905,N_1937,N_1410);
xnor U2906 (N_2906,N_1897,N_1162);
nor U2907 (N_2907,N_1883,N_1547);
nor U2908 (N_2908,N_1268,N_1646);
nand U2909 (N_2909,N_1277,N_1550);
nor U2910 (N_2910,N_1310,N_1094);
nor U2911 (N_2911,N_1125,N_1134);
xor U2912 (N_2912,N_1616,N_1329);
and U2913 (N_2913,N_1054,N_1527);
or U2914 (N_2914,N_1090,N_1592);
nand U2915 (N_2915,N_1636,N_1980);
xnor U2916 (N_2916,N_1959,N_1405);
nor U2917 (N_2917,N_1729,N_1782);
nand U2918 (N_2918,N_1517,N_1473);
xor U2919 (N_2919,N_1459,N_1820);
or U2920 (N_2920,N_1604,N_1362);
and U2921 (N_2921,N_1893,N_1382);
nand U2922 (N_2922,N_1495,N_1760);
xor U2923 (N_2923,N_1152,N_1897);
nand U2924 (N_2924,N_1383,N_1130);
nand U2925 (N_2925,N_1615,N_1597);
and U2926 (N_2926,N_1550,N_1944);
xor U2927 (N_2927,N_1658,N_1043);
nor U2928 (N_2928,N_1064,N_1072);
and U2929 (N_2929,N_1634,N_1732);
nor U2930 (N_2930,N_1560,N_1251);
xnor U2931 (N_2931,N_1937,N_1348);
nor U2932 (N_2932,N_1079,N_1159);
nor U2933 (N_2933,N_1683,N_1016);
nor U2934 (N_2934,N_1561,N_1105);
nor U2935 (N_2935,N_1427,N_1411);
and U2936 (N_2936,N_1700,N_1146);
and U2937 (N_2937,N_1827,N_1649);
xor U2938 (N_2938,N_1870,N_1133);
and U2939 (N_2939,N_1221,N_1592);
nand U2940 (N_2940,N_1206,N_1488);
nand U2941 (N_2941,N_1841,N_1975);
and U2942 (N_2942,N_1521,N_1768);
xor U2943 (N_2943,N_1256,N_1318);
nor U2944 (N_2944,N_1673,N_1918);
or U2945 (N_2945,N_1239,N_1401);
and U2946 (N_2946,N_1793,N_1444);
nor U2947 (N_2947,N_1988,N_1032);
xor U2948 (N_2948,N_1983,N_1932);
nand U2949 (N_2949,N_1780,N_1956);
or U2950 (N_2950,N_1897,N_1992);
nor U2951 (N_2951,N_1081,N_1496);
xor U2952 (N_2952,N_1323,N_1012);
xor U2953 (N_2953,N_1822,N_1097);
or U2954 (N_2954,N_1988,N_1751);
xnor U2955 (N_2955,N_1065,N_1229);
or U2956 (N_2956,N_1755,N_1737);
nand U2957 (N_2957,N_1993,N_1304);
nor U2958 (N_2958,N_1363,N_1820);
xnor U2959 (N_2959,N_1598,N_1344);
nand U2960 (N_2960,N_1394,N_1388);
and U2961 (N_2961,N_1069,N_1486);
xor U2962 (N_2962,N_1791,N_1625);
xnor U2963 (N_2963,N_1625,N_1562);
and U2964 (N_2964,N_1233,N_1784);
nor U2965 (N_2965,N_1875,N_1560);
nand U2966 (N_2966,N_1457,N_1143);
xor U2967 (N_2967,N_1313,N_1647);
xnor U2968 (N_2968,N_1926,N_1814);
nor U2969 (N_2969,N_1161,N_1821);
nor U2970 (N_2970,N_1638,N_1343);
xor U2971 (N_2971,N_1718,N_1656);
and U2972 (N_2972,N_1697,N_1965);
or U2973 (N_2973,N_1670,N_1405);
xor U2974 (N_2974,N_1201,N_1451);
xnor U2975 (N_2975,N_1903,N_1869);
nor U2976 (N_2976,N_1808,N_1615);
nor U2977 (N_2977,N_1947,N_1633);
xor U2978 (N_2978,N_1952,N_1227);
nor U2979 (N_2979,N_1533,N_1613);
xnor U2980 (N_2980,N_1551,N_1923);
nor U2981 (N_2981,N_1169,N_1896);
or U2982 (N_2982,N_1496,N_1851);
nor U2983 (N_2983,N_1611,N_1139);
nand U2984 (N_2984,N_1749,N_1993);
nand U2985 (N_2985,N_1690,N_1700);
nor U2986 (N_2986,N_1602,N_1041);
nand U2987 (N_2987,N_1576,N_1294);
xnor U2988 (N_2988,N_1280,N_1214);
nand U2989 (N_2989,N_1507,N_1024);
and U2990 (N_2990,N_1945,N_1786);
or U2991 (N_2991,N_1017,N_1438);
nand U2992 (N_2992,N_1917,N_1901);
xor U2993 (N_2993,N_1527,N_1953);
xor U2994 (N_2994,N_1726,N_1598);
xnor U2995 (N_2995,N_1226,N_1594);
or U2996 (N_2996,N_1993,N_1771);
nand U2997 (N_2997,N_1732,N_1594);
or U2998 (N_2998,N_1961,N_1547);
xor U2999 (N_2999,N_1871,N_1621);
or U3000 (N_3000,N_2245,N_2323);
nand U3001 (N_3001,N_2355,N_2979);
or U3002 (N_3002,N_2678,N_2110);
nor U3003 (N_3003,N_2268,N_2390);
xor U3004 (N_3004,N_2457,N_2755);
nand U3005 (N_3005,N_2008,N_2003);
nor U3006 (N_3006,N_2058,N_2122);
xnor U3007 (N_3007,N_2121,N_2502);
xor U3008 (N_3008,N_2252,N_2057);
or U3009 (N_3009,N_2509,N_2223);
xnor U3010 (N_3010,N_2129,N_2653);
and U3011 (N_3011,N_2210,N_2422);
and U3012 (N_3012,N_2490,N_2750);
or U3013 (N_3013,N_2764,N_2956);
or U3014 (N_3014,N_2507,N_2049);
nor U3015 (N_3015,N_2256,N_2214);
or U3016 (N_3016,N_2917,N_2135);
nor U3017 (N_3017,N_2155,N_2530);
xnor U3018 (N_3018,N_2083,N_2013);
or U3019 (N_3019,N_2221,N_2233);
nand U3020 (N_3020,N_2952,N_2145);
nand U3021 (N_3021,N_2515,N_2191);
and U3022 (N_3022,N_2877,N_2452);
or U3023 (N_3023,N_2026,N_2649);
nand U3024 (N_3024,N_2718,N_2685);
nand U3025 (N_3025,N_2944,N_2435);
xnor U3026 (N_3026,N_2666,N_2411);
nand U3027 (N_3027,N_2265,N_2237);
nor U3028 (N_3028,N_2019,N_2137);
or U3029 (N_3029,N_2698,N_2269);
and U3030 (N_3030,N_2364,N_2492);
nor U3031 (N_3031,N_2747,N_2097);
nor U3032 (N_3032,N_2186,N_2152);
nor U3033 (N_3033,N_2427,N_2392);
nand U3034 (N_3034,N_2339,N_2220);
nand U3035 (N_3035,N_2286,N_2035);
or U3036 (N_3036,N_2527,N_2591);
nand U3037 (N_3037,N_2535,N_2384);
nor U3038 (N_3038,N_2838,N_2119);
or U3039 (N_3039,N_2825,N_2880);
and U3040 (N_3040,N_2402,N_2549);
or U3041 (N_3041,N_2925,N_2757);
nand U3042 (N_3042,N_2520,N_2229);
or U3043 (N_3043,N_2327,N_2499);
or U3044 (N_3044,N_2789,N_2031);
xor U3045 (N_3045,N_2556,N_2710);
or U3046 (N_3046,N_2408,N_2335);
nand U3047 (N_3047,N_2354,N_2234);
nand U3048 (N_3048,N_2612,N_2028);
and U3049 (N_3049,N_2105,N_2892);
nor U3050 (N_3050,N_2174,N_2781);
nor U3051 (N_3051,N_2547,N_2136);
and U3052 (N_3052,N_2118,N_2450);
and U3053 (N_3053,N_2166,N_2333);
xor U3054 (N_3054,N_2273,N_2846);
and U3055 (N_3055,N_2874,N_2644);
and U3056 (N_3056,N_2768,N_2312);
or U3057 (N_3057,N_2990,N_2040);
and U3058 (N_3058,N_2720,N_2397);
and U3059 (N_3059,N_2976,N_2093);
xnor U3060 (N_3060,N_2444,N_2203);
and U3061 (N_3061,N_2580,N_2984);
or U3062 (N_3062,N_2317,N_2211);
or U3063 (N_3063,N_2033,N_2544);
and U3064 (N_3064,N_2721,N_2421);
nor U3065 (N_3065,N_2415,N_2651);
or U3066 (N_3066,N_2348,N_2792);
or U3067 (N_3067,N_2997,N_2039);
nand U3068 (N_3068,N_2887,N_2868);
nand U3069 (N_3069,N_2261,N_2297);
nand U3070 (N_3070,N_2821,N_2271);
xor U3071 (N_3071,N_2740,N_2241);
or U3072 (N_3072,N_2852,N_2529);
and U3073 (N_3073,N_2132,N_2611);
nor U3074 (N_3074,N_2733,N_2454);
and U3075 (N_3075,N_2985,N_2262);
nor U3076 (N_3076,N_2077,N_2120);
or U3077 (N_3077,N_2487,N_2730);
xor U3078 (N_3078,N_2400,N_2212);
nor U3079 (N_3079,N_2907,N_2690);
nand U3080 (N_3080,N_2282,N_2441);
nor U3081 (N_3081,N_2064,N_2330);
nand U3082 (N_3082,N_2622,N_2053);
xnor U3083 (N_3083,N_2518,N_2165);
nor U3084 (N_3084,N_2066,N_2618);
xnor U3085 (N_3085,N_2715,N_2981);
xor U3086 (N_3086,N_2108,N_2695);
and U3087 (N_3087,N_2560,N_2894);
or U3088 (N_3088,N_2876,N_2939);
nand U3089 (N_3089,N_2117,N_2586);
xnor U3090 (N_3090,N_2433,N_2180);
nor U3091 (N_3091,N_2404,N_2055);
xnor U3092 (N_3092,N_2929,N_2193);
and U3093 (N_3093,N_2731,N_2970);
nand U3094 (N_3094,N_2687,N_2293);
and U3095 (N_3095,N_2773,N_2665);
nor U3096 (N_3096,N_2722,N_2187);
nand U3097 (N_3097,N_2541,N_2555);
xor U3098 (N_3098,N_2379,N_2760);
and U3099 (N_3099,N_2729,N_2709);
or U3100 (N_3100,N_2700,N_2216);
and U3101 (N_3101,N_2482,N_2603);
or U3102 (N_3102,N_2368,N_2928);
nand U3103 (N_3103,N_2414,N_2664);
or U3104 (N_3104,N_2817,N_2696);
nand U3105 (N_3105,N_2858,N_2699);
xor U3106 (N_3106,N_2385,N_2124);
or U3107 (N_3107,N_2519,N_2113);
nand U3108 (N_3108,N_2139,N_2326);
nor U3109 (N_3109,N_2481,N_2258);
and U3110 (N_3110,N_2996,N_2311);
or U3111 (N_3111,N_2409,N_2636);
or U3112 (N_3112,N_2426,N_2992);
and U3113 (N_3113,N_2360,N_2631);
and U3114 (N_3114,N_2926,N_2418);
or U3115 (N_3115,N_2043,N_2584);
or U3116 (N_3116,N_2913,N_2465);
or U3117 (N_3117,N_2671,N_2375);
nor U3118 (N_3118,N_2936,N_2147);
and U3119 (N_3119,N_2488,N_2613);
xnor U3120 (N_3120,N_2153,N_2771);
or U3121 (N_3121,N_2227,N_2986);
and U3122 (N_3122,N_2845,N_2102);
nand U3123 (N_3123,N_2403,N_2785);
nand U3124 (N_3124,N_2957,N_2483);
xor U3125 (N_3125,N_2107,N_2809);
and U3126 (N_3126,N_2272,N_2472);
xnor U3127 (N_3127,N_2562,N_2445);
nor U3128 (N_3128,N_2862,N_2370);
or U3129 (N_3129,N_2471,N_2900);
nand U3130 (N_3130,N_2103,N_2559);
or U3131 (N_3131,N_2299,N_2030);
and U3132 (N_3132,N_2170,N_2181);
and U3133 (N_3133,N_2577,N_2667);
and U3134 (N_3134,N_2126,N_2082);
xor U3135 (N_3135,N_2842,N_2176);
nor U3136 (N_3136,N_2313,N_2151);
nand U3137 (N_3137,N_2154,N_2701);
nand U3138 (N_3138,N_2167,N_2937);
xor U3139 (N_3139,N_2728,N_2278);
and U3140 (N_3140,N_2410,N_2006);
nand U3141 (N_3141,N_2919,N_2989);
and U3142 (N_3142,N_2448,N_2079);
and U3143 (N_3143,N_2524,N_2340);
xnor U3144 (N_3144,N_2206,N_2620);
or U3145 (N_3145,N_2169,N_2829);
nand U3146 (N_3146,N_2726,N_2969);
and U3147 (N_3147,N_2534,N_2351);
or U3148 (N_3148,N_2114,N_2383);
xnor U3149 (N_3149,N_2776,N_2194);
and U3150 (N_3150,N_2587,N_2548);
and U3151 (N_3151,N_2904,N_2641);
xor U3152 (N_3152,N_2546,N_2761);
nand U3153 (N_3153,N_2861,N_2982);
nor U3154 (N_3154,N_2707,N_2660);
and U3155 (N_3155,N_2735,N_2935);
xnor U3156 (N_3156,N_2020,N_2627);
xor U3157 (N_3157,N_2998,N_2634);
xor U3158 (N_3158,N_2069,N_2865);
nor U3159 (N_3159,N_2600,N_2443);
nand U3160 (N_3160,N_2253,N_2532);
xnor U3161 (N_3161,N_2281,N_2012);
or U3162 (N_3162,N_2350,N_2288);
or U3163 (N_3163,N_2086,N_2867);
or U3164 (N_3164,N_2745,N_2372);
xor U3165 (N_3165,N_2361,N_2793);
nand U3166 (N_3166,N_2898,N_2849);
nand U3167 (N_3167,N_2130,N_2319);
xnor U3168 (N_3168,N_2300,N_2816);
xnor U3169 (N_3169,N_2830,N_2772);
and U3170 (N_3170,N_2276,N_2801);
nor U3171 (N_3171,N_2094,N_2207);
and U3172 (N_3172,N_2381,N_2419);
nor U3173 (N_3173,N_2920,N_2891);
xor U3174 (N_3174,N_2914,N_2938);
and U3175 (N_3175,N_2249,N_2398);
and U3176 (N_3176,N_2828,N_2479);
nor U3177 (N_3177,N_2609,N_2374);
xnor U3178 (N_3178,N_2041,N_2934);
and U3179 (N_3179,N_2759,N_2820);
or U3180 (N_3180,N_2886,N_2557);
nor U3181 (N_3181,N_2623,N_2686);
and U3182 (N_3182,N_2150,N_2042);
xnor U3183 (N_3183,N_2598,N_2065);
xor U3184 (N_3184,N_2633,N_2460);
nand U3185 (N_3185,N_2185,N_2201);
nor U3186 (N_3186,N_2133,N_2542);
nand U3187 (N_3187,N_2236,N_2942);
xnor U3188 (N_3188,N_2022,N_2257);
nor U3189 (N_3189,N_2883,N_2684);
and U3190 (N_3190,N_2682,N_2960);
or U3191 (N_3191,N_2209,N_2583);
and U3192 (N_3192,N_2662,N_2554);
or U3193 (N_3193,N_2439,N_2654);
nand U3194 (N_3194,N_2142,N_2163);
nand U3195 (N_3195,N_2356,N_2841);
or U3196 (N_3196,N_2589,N_2178);
and U3197 (N_3197,N_2357,N_2279);
xnor U3198 (N_3198,N_2882,N_2916);
xnor U3199 (N_3199,N_2850,N_2432);
or U3200 (N_3200,N_2184,N_2791);
nor U3201 (N_3201,N_2966,N_2582);
and U3202 (N_3202,N_2819,N_2736);
nand U3203 (N_3203,N_2870,N_2744);
nand U3204 (N_3204,N_2329,N_2506);
and U3205 (N_3205,N_2576,N_2787);
xor U3206 (N_3206,N_2769,N_2840);
or U3207 (N_3207,N_2538,N_2005);
xnor U3208 (N_3208,N_2616,N_2804);
and U3209 (N_3209,N_2436,N_2200);
or U3210 (N_3210,N_2672,N_2522);
nand U3211 (N_3211,N_2024,N_2243);
and U3212 (N_3212,N_2988,N_2303);
nand U3213 (N_3213,N_2172,N_2663);
and U3214 (N_3214,N_2797,N_2014);
xor U3215 (N_3215,N_2235,N_2247);
nor U3216 (N_3216,N_2061,N_2503);
nand U3217 (N_3217,N_2608,N_2645);
xnor U3218 (N_3218,N_2343,N_2358);
xor U3219 (N_3219,N_2377,N_2910);
or U3220 (N_3220,N_2959,N_2972);
xor U3221 (N_3221,N_2625,N_2902);
and U3222 (N_3222,N_2440,N_2141);
or U3223 (N_3223,N_2011,N_2521);
nor U3224 (N_3224,N_2060,N_2630);
nor U3225 (N_3225,N_2318,N_2067);
nor U3226 (N_3226,N_2007,N_2470);
and U3227 (N_3227,N_2885,N_2078);
nand U3228 (N_3228,N_2869,N_2903);
or U3229 (N_3229,N_2248,N_2459);
xor U3230 (N_3230,N_2328,N_2376);
or U3231 (N_3231,N_2073,N_2018);
and U3232 (N_3232,N_2795,N_2691);
nand U3233 (N_3233,N_2179,N_2978);
or U3234 (N_3234,N_2893,N_2637);
nand U3235 (N_3235,N_2911,N_2713);
nor U3236 (N_3236,N_2341,N_2805);
and U3237 (N_3237,N_2337,N_2578);
nand U3238 (N_3238,N_2688,N_2983);
xor U3239 (N_3239,N_2566,N_2486);
nor U3240 (N_3240,N_2629,N_2594);
and U3241 (N_3241,N_2752,N_2332);
xor U3242 (N_3242,N_2453,N_2474);
and U3243 (N_3243,N_2489,N_2756);
xnor U3244 (N_3244,N_2263,N_2463);
nor U3245 (N_3245,N_2270,N_2412);
and U3246 (N_3246,N_2941,N_2674);
or U3247 (N_3247,N_2727,N_2071);
or U3248 (N_3248,N_2912,N_2267);
xnor U3249 (N_3249,N_2588,N_2540);
and U3250 (N_3250,N_2128,N_2423);
nor U3251 (N_3251,N_2951,N_2669);
nand U3252 (N_3252,N_2425,N_2283);
xor U3253 (N_3253,N_2628,N_2306);
and U3254 (N_3254,N_2724,N_2708);
nand U3255 (N_3255,N_2601,N_2860);
and U3256 (N_3256,N_2950,N_2188);
and U3257 (N_3257,N_2505,N_2794);
nand U3258 (N_3258,N_2689,N_2626);
nand U3259 (N_3259,N_2373,N_2813);
xor U3260 (N_3260,N_2469,N_2417);
and U3261 (N_3261,N_2146,N_2182);
xor U3262 (N_3262,N_2851,N_2796);
and U3263 (N_3263,N_2751,N_2536);
nand U3264 (N_3264,N_2703,N_2516);
nand U3265 (N_3265,N_2899,N_2431);
xor U3266 (N_3266,N_2034,N_2072);
and U3267 (N_3267,N_2823,N_2037);
and U3268 (N_3268,N_2219,N_2572);
nand U3269 (N_3269,N_2717,N_2856);
nor U3270 (N_3270,N_2552,N_2734);
and U3271 (N_3271,N_2054,N_2602);
or U3272 (N_3272,N_2059,N_2918);
nand U3273 (N_3273,N_2029,N_2810);
and U3274 (N_3274,N_2430,N_2676);
xor U3275 (N_3275,N_2619,N_2106);
or U3276 (N_3276,N_2994,N_2812);
nor U3277 (N_3277,N_2705,N_2712);
and U3278 (N_3278,N_2822,N_2692);
nor U3279 (N_3279,N_2826,N_2510);
and U3280 (N_3280,N_2224,N_2254);
nor U3281 (N_3281,N_2954,N_2240);
and U3282 (N_3282,N_2526,N_2777);
xor U3283 (N_3283,N_2251,N_2101);
or U3284 (N_3284,N_2009,N_2407);
or U3285 (N_3285,N_2016,N_2818);
and U3286 (N_3286,N_2884,N_2084);
or U3287 (N_3287,N_2001,N_2015);
xnor U3288 (N_3288,N_2790,N_2087);
nand U3289 (N_3289,N_2378,N_2275);
or U3290 (N_3290,N_2295,N_2774);
or U3291 (N_3291,N_2324,N_2814);
or U3292 (N_3292,N_2561,N_2824);
or U3293 (N_3293,N_2640,N_2632);
xnor U3294 (N_3294,N_2239,N_2746);
or U3295 (N_3295,N_2112,N_2274);
nand U3296 (N_3296,N_2606,N_2881);
nor U3297 (N_3297,N_2593,N_2585);
nor U3298 (N_3298,N_2833,N_2635);
nor U3299 (N_3299,N_2565,N_2766);
xor U3300 (N_3300,N_2010,N_2109);
nand U3301 (N_3301,N_2788,N_2215);
nand U3302 (N_3302,N_2831,N_2366);
nand U3303 (N_3303,N_2322,N_2943);
and U3304 (N_3304,N_2171,N_2706);
and U3305 (N_3305,N_2661,N_2802);
or U3306 (N_3306,N_2347,N_2222);
or U3307 (N_3307,N_2617,N_2429);
and U3308 (N_3308,N_2396,N_2310);
nand U3309 (N_3309,N_2111,N_2308);
or U3310 (N_3310,N_2099,N_2023);
xnor U3311 (N_3311,N_2570,N_2052);
nand U3312 (N_3312,N_2621,N_2140);
or U3313 (N_3313,N_2779,N_2843);
or U3314 (N_3314,N_2697,N_2681);
nand U3315 (N_3315,N_2504,N_2859);
and U3316 (N_3316,N_2314,N_2517);
or U3317 (N_3317,N_2763,N_2497);
nand U3318 (N_3318,N_2284,N_2144);
nand U3319 (N_3319,N_2704,N_2915);
xnor U3320 (N_3320,N_2424,N_2362);
xnor U3321 (N_3321,N_2924,N_2056);
nor U3322 (N_3322,N_2879,N_2342);
and U3323 (N_3323,N_2890,N_2449);
and U3324 (N_3324,N_2947,N_2080);
and U3325 (N_3325,N_2615,N_2693);
nor U3326 (N_3326,N_2420,N_2778);
or U3327 (N_3327,N_2204,N_2352);
nor U3328 (N_3328,N_2655,N_2017);
or U3329 (N_3329,N_2437,N_2955);
xnor U3330 (N_3330,N_2298,N_2550);
nor U3331 (N_3331,N_2783,N_2296);
nand U3332 (N_3332,N_2451,N_2940);
or U3333 (N_3333,N_2558,N_2406);
xnor U3334 (N_3334,N_2605,N_2723);
nand U3335 (N_3335,N_2250,N_2091);
nand U3336 (N_3336,N_2889,N_2305);
xor U3337 (N_3337,N_2725,N_2977);
nor U3338 (N_3338,N_2604,N_2315);
xor U3339 (N_3339,N_2599,N_2088);
nor U3340 (N_3340,N_2480,N_2199);
nor U3341 (N_3341,N_2905,N_2921);
nand U3342 (N_3342,N_2157,N_2349);
xor U3343 (N_3343,N_2738,N_2658);
and U3344 (N_3344,N_2213,N_2189);
nor U3345 (N_3345,N_2786,N_2508);
and U3346 (N_3346,N_2906,N_2075);
or U3347 (N_3347,N_2719,N_2543);
and U3348 (N_3348,N_2711,N_2878);
and U3349 (N_3349,N_2923,N_2447);
and U3350 (N_3350,N_2739,N_2477);
xor U3351 (N_3351,N_2922,N_2456);
nand U3352 (N_3352,N_2592,N_2948);
or U3353 (N_3353,N_2573,N_2473);
xnor U3354 (N_3354,N_2002,N_2334);
nor U3355 (N_3355,N_2149,N_2607);
nor U3356 (N_3356,N_2945,N_2036);
xnor U3357 (N_3357,N_2673,N_2993);
or U3358 (N_3358,N_2044,N_2564);
nor U3359 (N_3359,N_2624,N_2595);
or U3360 (N_3360,N_2501,N_2382);
and U3361 (N_3361,N_2962,N_2369);
and U3362 (N_3362,N_2827,N_2742);
nor U3363 (N_3363,N_2597,N_2895);
nand U3364 (N_3364,N_2127,N_2173);
or U3365 (N_3365,N_2967,N_2748);
nor U3366 (N_3366,N_2571,N_2123);
xor U3367 (N_3367,N_2961,N_2949);
and U3368 (N_3368,N_2873,N_2574);
nor U3369 (N_3369,N_2965,N_2980);
and U3370 (N_3370,N_2537,N_2875);
xnor U3371 (N_3371,N_2659,N_2964);
xnor U3372 (N_3372,N_2231,N_2089);
nand U3373 (N_3373,N_2391,N_2438);
nand U3374 (N_3374,N_2468,N_2754);
nand U3375 (N_3375,N_2836,N_2834);
nand U3376 (N_3376,N_2289,N_2901);
nor U3377 (N_3377,N_2192,N_2590);
nand U3378 (N_3378,N_2762,N_2177);
and U3379 (N_3379,N_2025,N_2539);
xnor U3380 (N_3380,N_2496,N_2394);
xor U3381 (N_3381,N_2897,N_2975);
and U3382 (N_3382,N_2244,N_2927);
nand U3383 (N_3383,N_2027,N_2161);
or U3384 (N_3384,N_2255,N_2325);
nor U3385 (N_3385,N_2683,N_2260);
or U3386 (N_3386,N_2680,N_2800);
nand U3387 (N_3387,N_2386,N_2467);
xnor U3388 (N_3388,N_2525,N_2413);
and U3389 (N_3389,N_2485,N_2478);
nor U3390 (N_3390,N_2032,N_2047);
nand U3391 (N_3391,N_2183,N_2092);
and U3392 (N_3392,N_2643,N_2000);
or U3393 (N_3393,N_2365,N_2958);
xnor U3394 (N_3394,N_2125,N_2464);
or U3395 (N_3395,N_2076,N_2553);
or U3396 (N_3396,N_2280,N_2259);
nor U3397 (N_3397,N_2090,N_2301);
nor U3398 (N_3398,N_2070,N_2749);
and U3399 (N_3399,N_2732,N_2021);
nand U3400 (N_3400,N_2514,N_2931);
nand U3401 (N_3401,N_2835,N_2971);
nor U3402 (N_3402,N_2782,N_2551);
nor U3403 (N_3403,N_2395,N_2484);
or U3404 (N_3404,N_2495,N_2238);
xor U3405 (N_3405,N_2932,N_2353);
nor U3406 (N_3406,N_2675,N_2371);
and U3407 (N_3407,N_2491,N_2610);
nor U3408 (N_3408,N_2714,N_2896);
and U3409 (N_3409,N_2987,N_2045);
or U3410 (N_3410,N_2434,N_2500);
xnor U3411 (N_3411,N_2798,N_2513);
and U3412 (N_3412,N_2848,N_2815);
xor U3413 (N_3413,N_2226,N_2716);
nand U3414 (N_3414,N_2569,N_2933);
or U3415 (N_3415,N_2694,N_2854);
or U3416 (N_3416,N_2098,N_2331);
or U3417 (N_3417,N_2399,N_2156);
nor U3418 (N_3418,N_2668,N_2498);
nor U3419 (N_3419,N_2533,N_2100);
or U3420 (N_3420,N_2837,N_2266);
nor U3421 (N_3421,N_2999,N_2346);
nor U3422 (N_3422,N_2148,N_2232);
xnor U3423 (N_3423,N_2531,N_2446);
nand U3424 (N_3424,N_2051,N_2758);
nor U3425 (N_3425,N_2175,N_2642);
nor U3426 (N_3426,N_2866,N_2345);
or U3427 (N_3427,N_2839,N_2038);
and U3428 (N_3428,N_2770,N_2442);
and U3429 (N_3429,N_2162,N_2466);
xnor U3430 (N_3430,N_2277,N_2799);
nor U3431 (N_3431,N_2784,N_2294);
and U3432 (N_3432,N_2225,N_2545);
nor U3433 (N_3433,N_2462,N_2202);
nor U3434 (N_3434,N_2387,N_2285);
and U3435 (N_3435,N_2316,N_2638);
and U3436 (N_3436,N_2648,N_2190);
nor U3437 (N_3437,N_2405,N_2344);
xor U3438 (N_3438,N_2872,N_2198);
or U3439 (N_3439,N_2458,N_2995);
nand U3440 (N_3440,N_2806,N_2767);
nor U3441 (N_3441,N_2416,N_2096);
nor U3442 (N_3442,N_2568,N_2085);
and U3443 (N_3443,N_2832,N_2290);
nand U3444 (N_3444,N_2614,N_2775);
nor U3445 (N_3445,N_2380,N_2476);
and U3446 (N_3446,N_2575,N_2855);
or U3447 (N_3447,N_2197,N_2228);
nor U3448 (N_3448,N_2888,N_2808);
or U3449 (N_3449,N_2104,N_2304);
xor U3450 (N_3450,N_2677,N_2242);
xor U3451 (N_3451,N_2218,N_2230);
or U3452 (N_3452,N_2702,N_2196);
or U3453 (N_3453,N_2946,N_2063);
or U3454 (N_3454,N_2953,N_2307);
and U3455 (N_3455,N_2567,N_2074);
or U3456 (N_3456,N_2670,N_2363);
nor U3457 (N_3457,N_2579,N_2336);
nand U3458 (N_3458,N_2963,N_2753);
nand U3459 (N_3459,N_2168,N_2863);
nor U3460 (N_3460,N_2646,N_2974);
nor U3461 (N_3461,N_2679,N_2657);
or U3462 (N_3462,N_2743,N_2068);
nand U3463 (N_3463,N_2050,N_2143);
nor U3464 (N_3464,N_2393,N_2401);
and U3465 (N_3465,N_2475,N_2116);
nand U3466 (N_3466,N_2737,N_2493);
nand U3467 (N_3467,N_2246,N_2428);
xnor U3468 (N_3468,N_2844,N_2494);
xor U3469 (N_3469,N_2205,N_2511);
nor U3470 (N_3470,N_2596,N_2048);
nand U3471 (N_3471,N_2302,N_2388);
or U3472 (N_3472,N_2803,N_2159);
or U3473 (N_3473,N_2652,N_2164);
and U3474 (N_3474,N_2338,N_2847);
nor U3475 (N_3475,N_2639,N_2864);
or U3476 (N_3476,N_2004,N_2309);
or U3477 (N_3477,N_2853,N_2930);
and U3478 (N_3478,N_2647,N_2563);
nand U3479 (N_3479,N_2291,N_2807);
xor U3480 (N_3480,N_2160,N_2367);
nor U3481 (N_3481,N_2765,N_2991);
and U3482 (N_3482,N_2264,N_2741);
and U3483 (N_3483,N_2131,N_2389);
xnor U3484 (N_3484,N_2871,N_2968);
or U3485 (N_3485,N_2461,N_2528);
nor U3486 (N_3486,N_2062,N_2359);
nor U3487 (N_3487,N_2115,N_2857);
nor U3488 (N_3488,N_2973,N_2287);
or U3489 (N_3489,N_2134,N_2656);
nand U3490 (N_3490,N_2908,N_2650);
nor U3491 (N_3491,N_2046,N_2581);
nand U3492 (N_3492,N_2320,N_2455);
and U3493 (N_3493,N_2195,N_2292);
and U3494 (N_3494,N_2523,N_2138);
or U3495 (N_3495,N_2095,N_2909);
or U3496 (N_3496,N_2158,N_2081);
and U3497 (N_3497,N_2321,N_2512);
nor U3498 (N_3498,N_2217,N_2780);
xor U3499 (N_3499,N_2811,N_2208);
nor U3500 (N_3500,N_2530,N_2061);
or U3501 (N_3501,N_2929,N_2226);
nor U3502 (N_3502,N_2320,N_2714);
and U3503 (N_3503,N_2482,N_2339);
or U3504 (N_3504,N_2501,N_2627);
nor U3505 (N_3505,N_2122,N_2160);
nor U3506 (N_3506,N_2782,N_2291);
or U3507 (N_3507,N_2974,N_2585);
nor U3508 (N_3508,N_2519,N_2071);
nor U3509 (N_3509,N_2285,N_2404);
nor U3510 (N_3510,N_2818,N_2546);
and U3511 (N_3511,N_2411,N_2972);
or U3512 (N_3512,N_2064,N_2022);
or U3513 (N_3513,N_2310,N_2088);
or U3514 (N_3514,N_2038,N_2869);
nand U3515 (N_3515,N_2789,N_2089);
xor U3516 (N_3516,N_2531,N_2355);
or U3517 (N_3517,N_2525,N_2343);
and U3518 (N_3518,N_2733,N_2402);
or U3519 (N_3519,N_2006,N_2374);
or U3520 (N_3520,N_2550,N_2121);
or U3521 (N_3521,N_2524,N_2558);
and U3522 (N_3522,N_2619,N_2366);
nand U3523 (N_3523,N_2549,N_2858);
or U3524 (N_3524,N_2100,N_2416);
xnor U3525 (N_3525,N_2810,N_2596);
or U3526 (N_3526,N_2991,N_2870);
xnor U3527 (N_3527,N_2267,N_2675);
nand U3528 (N_3528,N_2856,N_2030);
xor U3529 (N_3529,N_2707,N_2992);
or U3530 (N_3530,N_2341,N_2200);
or U3531 (N_3531,N_2102,N_2516);
nor U3532 (N_3532,N_2885,N_2119);
nand U3533 (N_3533,N_2684,N_2141);
nand U3534 (N_3534,N_2937,N_2258);
nor U3535 (N_3535,N_2313,N_2898);
xor U3536 (N_3536,N_2027,N_2117);
nand U3537 (N_3537,N_2728,N_2613);
xnor U3538 (N_3538,N_2909,N_2637);
nand U3539 (N_3539,N_2082,N_2758);
or U3540 (N_3540,N_2390,N_2601);
nor U3541 (N_3541,N_2711,N_2458);
nor U3542 (N_3542,N_2496,N_2472);
or U3543 (N_3543,N_2515,N_2619);
or U3544 (N_3544,N_2115,N_2169);
and U3545 (N_3545,N_2246,N_2696);
nand U3546 (N_3546,N_2683,N_2209);
nand U3547 (N_3547,N_2875,N_2250);
nand U3548 (N_3548,N_2422,N_2167);
or U3549 (N_3549,N_2806,N_2850);
or U3550 (N_3550,N_2933,N_2735);
nand U3551 (N_3551,N_2193,N_2149);
or U3552 (N_3552,N_2879,N_2624);
or U3553 (N_3553,N_2997,N_2379);
xnor U3554 (N_3554,N_2592,N_2173);
nor U3555 (N_3555,N_2520,N_2069);
or U3556 (N_3556,N_2654,N_2112);
xor U3557 (N_3557,N_2799,N_2725);
nor U3558 (N_3558,N_2017,N_2208);
nand U3559 (N_3559,N_2679,N_2133);
nor U3560 (N_3560,N_2598,N_2257);
nand U3561 (N_3561,N_2240,N_2241);
nand U3562 (N_3562,N_2715,N_2428);
nand U3563 (N_3563,N_2745,N_2273);
or U3564 (N_3564,N_2091,N_2766);
nor U3565 (N_3565,N_2033,N_2907);
and U3566 (N_3566,N_2739,N_2908);
or U3567 (N_3567,N_2936,N_2121);
nand U3568 (N_3568,N_2970,N_2619);
and U3569 (N_3569,N_2962,N_2496);
or U3570 (N_3570,N_2441,N_2011);
nand U3571 (N_3571,N_2309,N_2622);
nor U3572 (N_3572,N_2511,N_2387);
and U3573 (N_3573,N_2178,N_2332);
xnor U3574 (N_3574,N_2315,N_2290);
or U3575 (N_3575,N_2329,N_2519);
nor U3576 (N_3576,N_2438,N_2260);
nor U3577 (N_3577,N_2215,N_2492);
xor U3578 (N_3578,N_2368,N_2162);
nand U3579 (N_3579,N_2889,N_2795);
and U3580 (N_3580,N_2447,N_2721);
xnor U3581 (N_3581,N_2613,N_2468);
nor U3582 (N_3582,N_2989,N_2710);
nand U3583 (N_3583,N_2068,N_2456);
nor U3584 (N_3584,N_2757,N_2710);
or U3585 (N_3585,N_2678,N_2395);
nor U3586 (N_3586,N_2588,N_2526);
xnor U3587 (N_3587,N_2724,N_2328);
nand U3588 (N_3588,N_2153,N_2290);
nand U3589 (N_3589,N_2463,N_2765);
or U3590 (N_3590,N_2086,N_2918);
and U3591 (N_3591,N_2483,N_2407);
or U3592 (N_3592,N_2951,N_2538);
nor U3593 (N_3593,N_2943,N_2965);
or U3594 (N_3594,N_2431,N_2651);
xor U3595 (N_3595,N_2672,N_2012);
or U3596 (N_3596,N_2202,N_2777);
or U3597 (N_3597,N_2250,N_2628);
nand U3598 (N_3598,N_2481,N_2222);
or U3599 (N_3599,N_2942,N_2240);
nor U3600 (N_3600,N_2816,N_2593);
nand U3601 (N_3601,N_2977,N_2868);
nor U3602 (N_3602,N_2321,N_2547);
xnor U3603 (N_3603,N_2486,N_2383);
and U3604 (N_3604,N_2466,N_2214);
xor U3605 (N_3605,N_2166,N_2328);
nor U3606 (N_3606,N_2277,N_2921);
nand U3607 (N_3607,N_2467,N_2619);
nand U3608 (N_3608,N_2487,N_2312);
or U3609 (N_3609,N_2621,N_2457);
or U3610 (N_3610,N_2402,N_2671);
nor U3611 (N_3611,N_2690,N_2248);
xor U3612 (N_3612,N_2690,N_2458);
or U3613 (N_3613,N_2757,N_2376);
nand U3614 (N_3614,N_2580,N_2543);
and U3615 (N_3615,N_2920,N_2927);
nor U3616 (N_3616,N_2849,N_2572);
xnor U3617 (N_3617,N_2736,N_2003);
xor U3618 (N_3618,N_2250,N_2074);
and U3619 (N_3619,N_2514,N_2326);
nor U3620 (N_3620,N_2670,N_2014);
xor U3621 (N_3621,N_2492,N_2163);
nand U3622 (N_3622,N_2666,N_2869);
and U3623 (N_3623,N_2927,N_2677);
xor U3624 (N_3624,N_2165,N_2910);
nand U3625 (N_3625,N_2420,N_2504);
or U3626 (N_3626,N_2220,N_2699);
nand U3627 (N_3627,N_2182,N_2678);
nand U3628 (N_3628,N_2614,N_2337);
or U3629 (N_3629,N_2279,N_2804);
nand U3630 (N_3630,N_2238,N_2659);
or U3631 (N_3631,N_2838,N_2891);
nor U3632 (N_3632,N_2341,N_2357);
xor U3633 (N_3633,N_2248,N_2356);
nor U3634 (N_3634,N_2449,N_2223);
xor U3635 (N_3635,N_2471,N_2174);
and U3636 (N_3636,N_2089,N_2489);
and U3637 (N_3637,N_2495,N_2955);
nand U3638 (N_3638,N_2886,N_2479);
nor U3639 (N_3639,N_2838,N_2500);
xor U3640 (N_3640,N_2323,N_2886);
nor U3641 (N_3641,N_2268,N_2020);
xnor U3642 (N_3642,N_2121,N_2939);
nor U3643 (N_3643,N_2596,N_2339);
xnor U3644 (N_3644,N_2949,N_2826);
xor U3645 (N_3645,N_2980,N_2620);
or U3646 (N_3646,N_2921,N_2368);
and U3647 (N_3647,N_2735,N_2170);
nand U3648 (N_3648,N_2371,N_2426);
nor U3649 (N_3649,N_2017,N_2670);
or U3650 (N_3650,N_2950,N_2652);
nor U3651 (N_3651,N_2944,N_2558);
xnor U3652 (N_3652,N_2328,N_2180);
nand U3653 (N_3653,N_2109,N_2436);
nor U3654 (N_3654,N_2380,N_2832);
nand U3655 (N_3655,N_2905,N_2022);
nand U3656 (N_3656,N_2989,N_2633);
or U3657 (N_3657,N_2906,N_2478);
nor U3658 (N_3658,N_2457,N_2056);
xnor U3659 (N_3659,N_2629,N_2802);
nand U3660 (N_3660,N_2729,N_2804);
xnor U3661 (N_3661,N_2727,N_2765);
or U3662 (N_3662,N_2014,N_2224);
xor U3663 (N_3663,N_2888,N_2308);
xor U3664 (N_3664,N_2718,N_2414);
and U3665 (N_3665,N_2115,N_2409);
or U3666 (N_3666,N_2562,N_2602);
nand U3667 (N_3667,N_2292,N_2360);
nor U3668 (N_3668,N_2587,N_2934);
nand U3669 (N_3669,N_2715,N_2246);
nor U3670 (N_3670,N_2128,N_2407);
and U3671 (N_3671,N_2231,N_2946);
xnor U3672 (N_3672,N_2645,N_2586);
and U3673 (N_3673,N_2429,N_2703);
or U3674 (N_3674,N_2629,N_2336);
nor U3675 (N_3675,N_2538,N_2549);
nand U3676 (N_3676,N_2516,N_2849);
nor U3677 (N_3677,N_2458,N_2759);
and U3678 (N_3678,N_2181,N_2596);
nand U3679 (N_3679,N_2317,N_2745);
nor U3680 (N_3680,N_2497,N_2416);
and U3681 (N_3681,N_2436,N_2176);
and U3682 (N_3682,N_2136,N_2304);
nand U3683 (N_3683,N_2571,N_2283);
or U3684 (N_3684,N_2928,N_2798);
and U3685 (N_3685,N_2744,N_2525);
nor U3686 (N_3686,N_2919,N_2680);
nand U3687 (N_3687,N_2066,N_2481);
xnor U3688 (N_3688,N_2129,N_2520);
nor U3689 (N_3689,N_2568,N_2214);
or U3690 (N_3690,N_2225,N_2239);
xor U3691 (N_3691,N_2633,N_2732);
xnor U3692 (N_3692,N_2522,N_2067);
xor U3693 (N_3693,N_2975,N_2486);
nand U3694 (N_3694,N_2023,N_2216);
nor U3695 (N_3695,N_2301,N_2581);
or U3696 (N_3696,N_2577,N_2230);
nor U3697 (N_3697,N_2648,N_2218);
nor U3698 (N_3698,N_2428,N_2217);
and U3699 (N_3699,N_2111,N_2459);
nor U3700 (N_3700,N_2568,N_2054);
and U3701 (N_3701,N_2467,N_2526);
xnor U3702 (N_3702,N_2887,N_2633);
xor U3703 (N_3703,N_2569,N_2083);
and U3704 (N_3704,N_2648,N_2090);
or U3705 (N_3705,N_2927,N_2055);
nand U3706 (N_3706,N_2373,N_2517);
or U3707 (N_3707,N_2153,N_2184);
nand U3708 (N_3708,N_2424,N_2306);
xor U3709 (N_3709,N_2594,N_2550);
xor U3710 (N_3710,N_2126,N_2985);
nor U3711 (N_3711,N_2332,N_2593);
and U3712 (N_3712,N_2479,N_2921);
or U3713 (N_3713,N_2889,N_2206);
and U3714 (N_3714,N_2800,N_2684);
or U3715 (N_3715,N_2288,N_2233);
nor U3716 (N_3716,N_2165,N_2515);
and U3717 (N_3717,N_2234,N_2827);
nand U3718 (N_3718,N_2663,N_2132);
and U3719 (N_3719,N_2039,N_2279);
nand U3720 (N_3720,N_2160,N_2206);
nor U3721 (N_3721,N_2732,N_2367);
nand U3722 (N_3722,N_2075,N_2773);
xnor U3723 (N_3723,N_2605,N_2219);
nand U3724 (N_3724,N_2472,N_2124);
and U3725 (N_3725,N_2899,N_2077);
or U3726 (N_3726,N_2082,N_2408);
nand U3727 (N_3727,N_2485,N_2656);
or U3728 (N_3728,N_2608,N_2497);
nand U3729 (N_3729,N_2327,N_2439);
or U3730 (N_3730,N_2042,N_2890);
nand U3731 (N_3731,N_2934,N_2027);
xor U3732 (N_3732,N_2799,N_2756);
and U3733 (N_3733,N_2730,N_2603);
nor U3734 (N_3734,N_2633,N_2267);
xnor U3735 (N_3735,N_2998,N_2493);
and U3736 (N_3736,N_2101,N_2955);
nand U3737 (N_3737,N_2837,N_2117);
xor U3738 (N_3738,N_2890,N_2903);
nor U3739 (N_3739,N_2988,N_2485);
nand U3740 (N_3740,N_2448,N_2660);
nand U3741 (N_3741,N_2677,N_2164);
nand U3742 (N_3742,N_2180,N_2476);
or U3743 (N_3743,N_2104,N_2506);
nand U3744 (N_3744,N_2767,N_2644);
or U3745 (N_3745,N_2818,N_2699);
nand U3746 (N_3746,N_2716,N_2027);
xor U3747 (N_3747,N_2040,N_2736);
and U3748 (N_3748,N_2238,N_2072);
nand U3749 (N_3749,N_2671,N_2909);
nand U3750 (N_3750,N_2700,N_2063);
nor U3751 (N_3751,N_2109,N_2860);
nand U3752 (N_3752,N_2911,N_2317);
and U3753 (N_3753,N_2740,N_2270);
nor U3754 (N_3754,N_2550,N_2171);
or U3755 (N_3755,N_2705,N_2066);
or U3756 (N_3756,N_2946,N_2698);
nand U3757 (N_3757,N_2265,N_2694);
xor U3758 (N_3758,N_2205,N_2579);
and U3759 (N_3759,N_2573,N_2885);
nand U3760 (N_3760,N_2209,N_2325);
and U3761 (N_3761,N_2489,N_2805);
or U3762 (N_3762,N_2896,N_2620);
nand U3763 (N_3763,N_2394,N_2904);
nor U3764 (N_3764,N_2203,N_2701);
nand U3765 (N_3765,N_2539,N_2648);
nor U3766 (N_3766,N_2840,N_2002);
nor U3767 (N_3767,N_2943,N_2515);
or U3768 (N_3768,N_2701,N_2369);
or U3769 (N_3769,N_2483,N_2910);
nor U3770 (N_3770,N_2523,N_2365);
or U3771 (N_3771,N_2798,N_2602);
and U3772 (N_3772,N_2435,N_2623);
and U3773 (N_3773,N_2704,N_2234);
nand U3774 (N_3774,N_2542,N_2973);
and U3775 (N_3775,N_2054,N_2556);
nor U3776 (N_3776,N_2063,N_2777);
xor U3777 (N_3777,N_2476,N_2731);
nor U3778 (N_3778,N_2291,N_2371);
nand U3779 (N_3779,N_2246,N_2802);
and U3780 (N_3780,N_2424,N_2413);
nor U3781 (N_3781,N_2818,N_2081);
or U3782 (N_3782,N_2776,N_2834);
nand U3783 (N_3783,N_2237,N_2133);
xnor U3784 (N_3784,N_2302,N_2120);
xnor U3785 (N_3785,N_2108,N_2593);
xnor U3786 (N_3786,N_2590,N_2568);
nand U3787 (N_3787,N_2732,N_2728);
nor U3788 (N_3788,N_2806,N_2759);
nor U3789 (N_3789,N_2199,N_2451);
xor U3790 (N_3790,N_2735,N_2995);
nor U3791 (N_3791,N_2038,N_2540);
xor U3792 (N_3792,N_2653,N_2309);
and U3793 (N_3793,N_2779,N_2427);
nand U3794 (N_3794,N_2865,N_2100);
xnor U3795 (N_3795,N_2932,N_2710);
or U3796 (N_3796,N_2180,N_2452);
xnor U3797 (N_3797,N_2262,N_2604);
nor U3798 (N_3798,N_2223,N_2258);
xnor U3799 (N_3799,N_2828,N_2151);
or U3800 (N_3800,N_2450,N_2954);
and U3801 (N_3801,N_2975,N_2535);
nand U3802 (N_3802,N_2114,N_2106);
or U3803 (N_3803,N_2221,N_2230);
xor U3804 (N_3804,N_2246,N_2296);
nor U3805 (N_3805,N_2936,N_2375);
xor U3806 (N_3806,N_2528,N_2931);
nand U3807 (N_3807,N_2879,N_2912);
nor U3808 (N_3808,N_2080,N_2283);
nand U3809 (N_3809,N_2309,N_2183);
and U3810 (N_3810,N_2405,N_2946);
or U3811 (N_3811,N_2358,N_2325);
xor U3812 (N_3812,N_2263,N_2760);
nand U3813 (N_3813,N_2746,N_2351);
nor U3814 (N_3814,N_2089,N_2342);
xor U3815 (N_3815,N_2461,N_2651);
and U3816 (N_3816,N_2123,N_2736);
nand U3817 (N_3817,N_2720,N_2110);
nor U3818 (N_3818,N_2824,N_2434);
and U3819 (N_3819,N_2624,N_2787);
nand U3820 (N_3820,N_2437,N_2191);
nor U3821 (N_3821,N_2744,N_2696);
xor U3822 (N_3822,N_2057,N_2441);
and U3823 (N_3823,N_2894,N_2157);
and U3824 (N_3824,N_2988,N_2566);
nor U3825 (N_3825,N_2385,N_2174);
nand U3826 (N_3826,N_2216,N_2068);
nor U3827 (N_3827,N_2128,N_2154);
nor U3828 (N_3828,N_2919,N_2735);
nand U3829 (N_3829,N_2910,N_2310);
xnor U3830 (N_3830,N_2351,N_2499);
and U3831 (N_3831,N_2175,N_2359);
nor U3832 (N_3832,N_2740,N_2906);
and U3833 (N_3833,N_2597,N_2968);
xor U3834 (N_3834,N_2646,N_2127);
xnor U3835 (N_3835,N_2586,N_2738);
xnor U3836 (N_3836,N_2031,N_2249);
or U3837 (N_3837,N_2901,N_2530);
and U3838 (N_3838,N_2008,N_2811);
xnor U3839 (N_3839,N_2934,N_2318);
or U3840 (N_3840,N_2127,N_2361);
nor U3841 (N_3841,N_2010,N_2785);
and U3842 (N_3842,N_2678,N_2544);
or U3843 (N_3843,N_2607,N_2895);
nor U3844 (N_3844,N_2526,N_2927);
nor U3845 (N_3845,N_2904,N_2721);
and U3846 (N_3846,N_2513,N_2807);
xnor U3847 (N_3847,N_2231,N_2262);
and U3848 (N_3848,N_2618,N_2193);
or U3849 (N_3849,N_2811,N_2321);
and U3850 (N_3850,N_2163,N_2104);
nor U3851 (N_3851,N_2722,N_2261);
or U3852 (N_3852,N_2221,N_2257);
xor U3853 (N_3853,N_2393,N_2141);
or U3854 (N_3854,N_2294,N_2198);
xnor U3855 (N_3855,N_2387,N_2071);
or U3856 (N_3856,N_2498,N_2767);
nand U3857 (N_3857,N_2712,N_2830);
or U3858 (N_3858,N_2427,N_2739);
or U3859 (N_3859,N_2009,N_2004);
nand U3860 (N_3860,N_2984,N_2010);
xor U3861 (N_3861,N_2309,N_2588);
nand U3862 (N_3862,N_2476,N_2346);
or U3863 (N_3863,N_2237,N_2463);
nand U3864 (N_3864,N_2990,N_2018);
and U3865 (N_3865,N_2284,N_2386);
xnor U3866 (N_3866,N_2696,N_2535);
or U3867 (N_3867,N_2550,N_2201);
and U3868 (N_3868,N_2549,N_2811);
nand U3869 (N_3869,N_2975,N_2692);
and U3870 (N_3870,N_2478,N_2640);
or U3871 (N_3871,N_2766,N_2651);
nor U3872 (N_3872,N_2449,N_2166);
nand U3873 (N_3873,N_2587,N_2278);
nand U3874 (N_3874,N_2698,N_2814);
xor U3875 (N_3875,N_2765,N_2513);
xor U3876 (N_3876,N_2956,N_2863);
xnor U3877 (N_3877,N_2548,N_2777);
or U3878 (N_3878,N_2259,N_2610);
and U3879 (N_3879,N_2833,N_2153);
or U3880 (N_3880,N_2914,N_2183);
xor U3881 (N_3881,N_2213,N_2775);
and U3882 (N_3882,N_2949,N_2173);
xor U3883 (N_3883,N_2153,N_2818);
and U3884 (N_3884,N_2693,N_2977);
or U3885 (N_3885,N_2498,N_2074);
xnor U3886 (N_3886,N_2672,N_2290);
nand U3887 (N_3887,N_2218,N_2798);
xor U3888 (N_3888,N_2961,N_2060);
nand U3889 (N_3889,N_2737,N_2002);
or U3890 (N_3890,N_2939,N_2976);
xnor U3891 (N_3891,N_2626,N_2001);
and U3892 (N_3892,N_2432,N_2308);
and U3893 (N_3893,N_2084,N_2902);
or U3894 (N_3894,N_2012,N_2600);
and U3895 (N_3895,N_2106,N_2025);
xnor U3896 (N_3896,N_2153,N_2530);
nand U3897 (N_3897,N_2304,N_2035);
nand U3898 (N_3898,N_2690,N_2792);
or U3899 (N_3899,N_2633,N_2339);
xor U3900 (N_3900,N_2374,N_2884);
and U3901 (N_3901,N_2315,N_2580);
and U3902 (N_3902,N_2876,N_2185);
nand U3903 (N_3903,N_2784,N_2112);
or U3904 (N_3904,N_2258,N_2593);
nand U3905 (N_3905,N_2198,N_2325);
and U3906 (N_3906,N_2309,N_2580);
nor U3907 (N_3907,N_2284,N_2375);
or U3908 (N_3908,N_2944,N_2374);
and U3909 (N_3909,N_2519,N_2875);
xor U3910 (N_3910,N_2139,N_2313);
or U3911 (N_3911,N_2174,N_2053);
nand U3912 (N_3912,N_2754,N_2221);
and U3913 (N_3913,N_2353,N_2476);
or U3914 (N_3914,N_2073,N_2068);
nand U3915 (N_3915,N_2263,N_2866);
xnor U3916 (N_3916,N_2100,N_2601);
or U3917 (N_3917,N_2177,N_2467);
and U3918 (N_3918,N_2880,N_2455);
xor U3919 (N_3919,N_2390,N_2585);
xnor U3920 (N_3920,N_2254,N_2152);
xor U3921 (N_3921,N_2853,N_2384);
and U3922 (N_3922,N_2579,N_2581);
nand U3923 (N_3923,N_2013,N_2107);
xnor U3924 (N_3924,N_2823,N_2318);
nand U3925 (N_3925,N_2682,N_2156);
xnor U3926 (N_3926,N_2719,N_2720);
xor U3927 (N_3927,N_2776,N_2933);
xnor U3928 (N_3928,N_2157,N_2863);
nand U3929 (N_3929,N_2122,N_2825);
and U3930 (N_3930,N_2971,N_2538);
and U3931 (N_3931,N_2393,N_2566);
nand U3932 (N_3932,N_2612,N_2913);
xor U3933 (N_3933,N_2463,N_2328);
nand U3934 (N_3934,N_2918,N_2808);
nand U3935 (N_3935,N_2560,N_2528);
and U3936 (N_3936,N_2885,N_2125);
nor U3937 (N_3937,N_2592,N_2413);
or U3938 (N_3938,N_2254,N_2033);
nand U3939 (N_3939,N_2166,N_2935);
nand U3940 (N_3940,N_2165,N_2946);
nor U3941 (N_3941,N_2665,N_2777);
nand U3942 (N_3942,N_2862,N_2788);
nor U3943 (N_3943,N_2294,N_2836);
and U3944 (N_3944,N_2420,N_2347);
or U3945 (N_3945,N_2726,N_2750);
or U3946 (N_3946,N_2048,N_2414);
or U3947 (N_3947,N_2643,N_2826);
or U3948 (N_3948,N_2116,N_2834);
and U3949 (N_3949,N_2268,N_2550);
xor U3950 (N_3950,N_2751,N_2456);
and U3951 (N_3951,N_2404,N_2230);
nand U3952 (N_3952,N_2931,N_2148);
nor U3953 (N_3953,N_2173,N_2296);
nor U3954 (N_3954,N_2313,N_2770);
or U3955 (N_3955,N_2404,N_2985);
or U3956 (N_3956,N_2426,N_2885);
and U3957 (N_3957,N_2742,N_2015);
and U3958 (N_3958,N_2666,N_2279);
xnor U3959 (N_3959,N_2605,N_2497);
xnor U3960 (N_3960,N_2619,N_2351);
nand U3961 (N_3961,N_2249,N_2891);
or U3962 (N_3962,N_2349,N_2791);
xnor U3963 (N_3963,N_2331,N_2268);
and U3964 (N_3964,N_2321,N_2471);
or U3965 (N_3965,N_2088,N_2704);
or U3966 (N_3966,N_2067,N_2813);
nand U3967 (N_3967,N_2621,N_2085);
xnor U3968 (N_3968,N_2999,N_2232);
nor U3969 (N_3969,N_2832,N_2237);
and U3970 (N_3970,N_2837,N_2724);
or U3971 (N_3971,N_2000,N_2235);
nor U3972 (N_3972,N_2498,N_2568);
nand U3973 (N_3973,N_2838,N_2835);
xnor U3974 (N_3974,N_2623,N_2912);
xnor U3975 (N_3975,N_2444,N_2818);
or U3976 (N_3976,N_2131,N_2168);
nor U3977 (N_3977,N_2621,N_2536);
nor U3978 (N_3978,N_2931,N_2716);
and U3979 (N_3979,N_2830,N_2858);
and U3980 (N_3980,N_2986,N_2969);
nand U3981 (N_3981,N_2291,N_2343);
nand U3982 (N_3982,N_2797,N_2305);
or U3983 (N_3983,N_2650,N_2219);
nor U3984 (N_3984,N_2032,N_2856);
or U3985 (N_3985,N_2238,N_2695);
nor U3986 (N_3986,N_2103,N_2024);
nand U3987 (N_3987,N_2623,N_2184);
nor U3988 (N_3988,N_2299,N_2335);
and U3989 (N_3989,N_2736,N_2022);
nor U3990 (N_3990,N_2574,N_2547);
xnor U3991 (N_3991,N_2799,N_2360);
xor U3992 (N_3992,N_2732,N_2468);
nand U3993 (N_3993,N_2789,N_2924);
nor U3994 (N_3994,N_2108,N_2905);
nor U3995 (N_3995,N_2148,N_2425);
nand U3996 (N_3996,N_2342,N_2331);
and U3997 (N_3997,N_2291,N_2363);
xnor U3998 (N_3998,N_2893,N_2379);
nor U3999 (N_3999,N_2530,N_2171);
or U4000 (N_4000,N_3192,N_3281);
or U4001 (N_4001,N_3596,N_3983);
and U4002 (N_4002,N_3798,N_3120);
xnor U4003 (N_4003,N_3276,N_3986);
nand U4004 (N_4004,N_3115,N_3288);
and U4005 (N_4005,N_3413,N_3989);
nor U4006 (N_4006,N_3971,N_3965);
or U4007 (N_4007,N_3100,N_3722);
nor U4008 (N_4008,N_3287,N_3956);
or U4009 (N_4009,N_3300,N_3271);
nor U4010 (N_4010,N_3210,N_3675);
xnor U4011 (N_4011,N_3311,N_3072);
or U4012 (N_4012,N_3392,N_3724);
xor U4013 (N_4013,N_3107,N_3214);
or U4014 (N_4014,N_3329,N_3712);
and U4015 (N_4015,N_3158,N_3903);
nand U4016 (N_4016,N_3479,N_3929);
nand U4017 (N_4017,N_3713,N_3633);
nand U4018 (N_4018,N_3444,N_3146);
xor U4019 (N_4019,N_3901,N_3773);
and U4020 (N_4020,N_3246,N_3978);
nand U4021 (N_4021,N_3787,N_3314);
nand U4022 (N_4022,N_3186,N_3318);
xnor U4023 (N_4023,N_3942,N_3203);
nand U4024 (N_4024,N_3257,N_3124);
xor U4025 (N_4025,N_3395,N_3762);
xor U4026 (N_4026,N_3509,N_3967);
or U4027 (N_4027,N_3940,N_3735);
nor U4028 (N_4028,N_3524,N_3269);
nand U4029 (N_4029,N_3844,N_3270);
or U4030 (N_4030,N_3690,N_3157);
xor U4031 (N_4031,N_3170,N_3824);
nand U4032 (N_4032,N_3686,N_3662);
nor U4033 (N_4033,N_3795,N_3458);
nor U4034 (N_4034,N_3451,N_3799);
or U4035 (N_4035,N_3359,N_3499);
and U4036 (N_4036,N_3061,N_3969);
and U4037 (N_4037,N_3205,N_3467);
or U4038 (N_4038,N_3247,N_3278);
xor U4039 (N_4039,N_3382,N_3498);
nand U4040 (N_4040,N_3282,N_3054);
or U4041 (N_4041,N_3880,N_3347);
nand U4042 (N_4042,N_3216,N_3923);
xor U4043 (N_4043,N_3025,N_3489);
and U4044 (N_4044,N_3779,N_3400);
nand U4045 (N_4045,N_3226,N_3196);
or U4046 (N_4046,N_3574,N_3449);
nor U4047 (N_4047,N_3708,N_3757);
xor U4048 (N_4048,N_3551,N_3432);
or U4049 (N_4049,N_3599,N_3737);
and U4050 (N_4050,N_3114,N_3109);
xnor U4051 (N_4051,N_3731,N_3530);
or U4052 (N_4052,N_3304,N_3076);
nor U4053 (N_4053,N_3985,N_3587);
nor U4054 (N_4054,N_3041,N_3674);
and U4055 (N_4055,N_3485,N_3628);
nand U4056 (N_4056,N_3045,N_3249);
and U4057 (N_4057,N_3768,N_3084);
or U4058 (N_4058,N_3441,N_3884);
nor U4059 (N_4059,N_3429,N_3029);
nor U4060 (N_4060,N_3391,N_3906);
nor U4061 (N_4061,N_3236,N_3369);
and U4062 (N_4062,N_3122,N_3071);
nand U4063 (N_4063,N_3896,N_3046);
or U4064 (N_4064,N_3207,N_3062);
nand U4065 (N_4065,N_3361,N_3384);
xor U4066 (N_4066,N_3398,N_3232);
nor U4067 (N_4067,N_3776,N_3440);
and U4068 (N_4068,N_3190,N_3058);
or U4069 (N_4069,N_3865,N_3316);
or U4070 (N_4070,N_3958,N_3845);
or U4071 (N_4071,N_3945,N_3155);
xor U4072 (N_4072,N_3090,N_3411);
nand U4073 (N_4073,N_3693,N_3153);
and U4074 (N_4074,N_3434,N_3218);
nor U4075 (N_4075,N_3303,N_3982);
or U4076 (N_4076,N_3952,N_3372);
xnor U4077 (N_4077,N_3745,N_3809);
nor U4078 (N_4078,N_3459,N_3317);
or U4079 (N_4079,N_3033,N_3163);
nor U4080 (N_4080,N_3366,N_3728);
nand U4081 (N_4081,N_3723,N_3131);
nand U4082 (N_4082,N_3555,N_3789);
nand U4083 (N_4083,N_3658,N_3997);
and U4084 (N_4084,N_3556,N_3103);
nor U4085 (N_4085,N_3572,N_3618);
xor U4086 (N_4086,N_3553,N_3219);
and U4087 (N_4087,N_3493,N_3177);
nor U4088 (N_4088,N_3848,N_3537);
nand U4089 (N_4089,N_3515,N_3322);
and U4090 (N_4090,N_3563,N_3950);
or U4091 (N_4091,N_3520,N_3560);
and U4092 (N_4092,N_3354,N_3112);
and U4093 (N_4093,N_3665,N_3935);
and U4094 (N_4094,N_3301,N_3160);
or U4095 (N_4095,N_3453,N_3279);
or U4096 (N_4096,N_3682,N_3919);
or U4097 (N_4097,N_3603,N_3885);
xor U4098 (N_4098,N_3639,N_3904);
or U4099 (N_4099,N_3769,N_3073);
nand U4100 (N_4100,N_3777,N_3179);
nand U4101 (N_4101,N_3830,N_3250);
and U4102 (N_4102,N_3383,N_3476);
xor U4103 (N_4103,N_3835,N_3334);
nand U4104 (N_4104,N_3245,N_3889);
xor U4105 (N_4105,N_3370,N_3486);
xnor U4106 (N_4106,N_3636,N_3823);
nor U4107 (N_4107,N_3235,N_3379);
nor U4108 (N_4108,N_3828,N_3345);
and U4109 (N_4109,N_3943,N_3529);
nor U4110 (N_4110,N_3924,N_3204);
xor U4111 (N_4111,N_3150,N_3755);
xor U4112 (N_4112,N_3502,N_3512);
nor U4113 (N_4113,N_3957,N_3862);
xnor U4114 (N_4114,N_3389,N_3748);
or U4115 (N_4115,N_3129,N_3536);
or U4116 (N_4116,N_3454,N_3785);
xor U4117 (N_4117,N_3975,N_3653);
nand U4118 (N_4118,N_3183,N_3299);
or U4119 (N_4119,N_3496,N_3854);
nor U4120 (N_4120,N_3034,N_3240);
xnor U4121 (N_4121,N_3918,N_3101);
xnor U4122 (N_4122,N_3871,N_3656);
nand U4123 (N_4123,N_3173,N_3792);
xor U4124 (N_4124,N_3456,N_3030);
nor U4125 (N_4125,N_3710,N_3364);
nor U4126 (N_4126,N_3998,N_3925);
xnor U4127 (N_4127,N_3315,N_3199);
nand U4128 (N_4128,N_3894,N_3293);
nand U4129 (N_4129,N_3996,N_3546);
nor U4130 (N_4130,N_3966,N_3338);
and U4131 (N_4131,N_3035,N_3691);
xnor U4132 (N_4132,N_3137,N_3254);
or U4133 (N_4133,N_3740,N_3552);
nor U4134 (N_4134,N_3143,N_3988);
nor U4135 (N_4135,N_3651,N_3002);
or U4136 (N_4136,N_3351,N_3853);
xor U4137 (N_4137,N_3744,N_3201);
and U4138 (N_4138,N_3911,N_3081);
and U4139 (N_4139,N_3800,N_3914);
or U4140 (N_4140,N_3284,N_3168);
and U4141 (N_4141,N_3027,N_3718);
nor U4142 (N_4142,N_3102,N_3857);
xor U4143 (N_4143,N_3538,N_3811);
or U4144 (N_4144,N_3253,N_3557);
or U4145 (N_4145,N_3415,N_3283);
or U4146 (N_4146,N_3421,N_3344);
nor U4147 (N_4147,N_3565,N_3772);
nand U4148 (N_4148,N_3267,N_3539);
xor U4149 (N_4149,N_3044,N_3012);
and U4150 (N_4150,N_3584,N_3607);
or U4151 (N_4151,N_3427,N_3770);
xnor U4152 (N_4152,N_3937,N_3938);
or U4153 (N_4153,N_3622,N_3910);
nand U4154 (N_4154,N_3841,N_3133);
or U4155 (N_4155,N_3482,N_3362);
nand U4156 (N_4156,N_3118,N_3891);
or U4157 (N_4157,N_3028,N_3660);
or U4158 (N_4158,N_3144,N_3328);
nand U4159 (N_4159,N_3360,N_3187);
xor U4160 (N_4160,N_3241,N_3796);
nand U4161 (N_4161,N_3700,N_3688);
xnor U4162 (N_4162,N_3393,N_3510);
nor U4163 (N_4163,N_3588,N_3961);
xnor U4164 (N_4164,N_3464,N_3922);
and U4165 (N_4165,N_3864,N_3088);
nand U4166 (N_4166,N_3503,N_3726);
and U4167 (N_4167,N_3403,N_3481);
nor U4168 (N_4168,N_3739,N_3264);
and U4169 (N_4169,N_3839,N_3976);
nor U4170 (N_4170,N_3319,N_3741);
xnor U4171 (N_4171,N_3290,N_3428);
nand U4172 (N_4172,N_3561,N_3015);
nor U4173 (N_4173,N_3963,N_3559);
xor U4174 (N_4174,N_3962,N_3332);
or U4175 (N_4175,N_3843,N_3649);
nand U4176 (N_4176,N_3635,N_3374);
xnor U4177 (N_4177,N_3514,N_3490);
or U4178 (N_4178,N_3475,N_3586);
or U4179 (N_4179,N_3380,N_3410);
nand U4180 (N_4180,N_3671,N_3385);
xnor U4181 (N_4181,N_3087,N_3888);
or U4182 (N_4182,N_3766,N_3794);
nand U4183 (N_4183,N_3927,N_3964);
nor U4184 (N_4184,N_3184,N_3926);
xor U4185 (N_4185,N_3518,N_3709);
nor U4186 (N_4186,N_3677,N_3343);
xor U4187 (N_4187,N_3544,N_3790);
and U4188 (N_4188,N_3019,N_3615);
or U4189 (N_4189,N_3363,N_3591);
xnor U4190 (N_4190,N_3683,N_3604);
nand U4191 (N_4191,N_3443,N_3791);
nor U4192 (N_4192,N_3111,N_3139);
xor U4193 (N_4193,N_3980,N_3172);
or U4194 (N_4194,N_3011,N_3861);
or U4195 (N_4195,N_3176,N_3039);
and U4196 (N_4196,N_3409,N_3225);
xor U4197 (N_4197,N_3274,N_3513);
xnor U4198 (N_4198,N_3681,N_3913);
or U4199 (N_4199,N_3221,N_3840);
xor U4200 (N_4200,N_3720,N_3350);
xor U4201 (N_4201,N_3113,N_3532);
nor U4202 (N_4202,N_3142,N_3230);
nand U4203 (N_4203,N_3178,N_3180);
nand U4204 (N_4204,N_3043,N_3883);
or U4205 (N_4205,N_3542,N_3188);
nor U4206 (N_4206,N_3620,N_3960);
nor U4207 (N_4207,N_3685,N_3702);
xor U4208 (N_4208,N_3916,N_3431);
and U4209 (N_4209,N_3223,N_3305);
nand U4210 (N_4210,N_3148,N_3959);
or U4211 (N_4211,N_3528,N_3801);
or U4212 (N_4212,N_3189,N_3121);
nor U4213 (N_4213,N_3605,N_3667);
xor U4214 (N_4214,N_3611,N_3175);
or U4215 (N_4215,N_3474,N_3075);
xor U4216 (N_4216,N_3418,N_3699);
xor U4217 (N_4217,N_3016,N_3472);
nor U4218 (N_4218,N_3097,N_3580);
or U4219 (N_4219,N_3302,N_3094);
nand U4220 (N_4220,N_3793,N_3010);
nand U4221 (N_4221,N_3069,N_3083);
and U4222 (N_4222,N_3086,N_3602);
xor U4223 (N_4223,N_3308,N_3838);
xor U4224 (N_4224,N_3953,N_3680);
and U4225 (N_4225,N_3535,N_3994);
or U4226 (N_4226,N_3321,N_3543);
nor U4227 (N_4227,N_3826,N_3078);
nor U4228 (N_4228,N_3941,N_3265);
or U4229 (N_4229,N_3469,N_3323);
and U4230 (N_4230,N_3417,N_3217);
or U4231 (N_4231,N_3774,N_3706);
nor U4232 (N_4232,N_3614,N_3208);
or U4233 (N_4233,N_3388,N_3096);
xnor U4234 (N_4234,N_3080,N_3928);
xnor U4235 (N_4235,N_3297,N_3753);
xnor U4236 (N_4236,N_3294,N_3036);
nand U4237 (N_4237,N_3024,N_3650);
or U4238 (N_4238,N_3820,N_3352);
nand U4239 (N_4239,N_3042,N_3438);
nand U4240 (N_4240,N_3729,N_3198);
and U4241 (N_4241,N_3435,N_3661);
nor U4242 (N_4242,N_3008,N_3306);
and U4243 (N_4243,N_3562,N_3815);
xnor U4244 (N_4244,N_3378,N_3972);
and U4245 (N_4245,N_3408,N_3664);
and U4246 (N_4246,N_3715,N_3298);
xor U4247 (N_4247,N_3295,N_3377);
or U4248 (N_4248,N_3095,N_3589);
nor U4249 (N_4249,N_3895,N_3642);
nor U4250 (N_4250,N_3161,N_3505);
nor U4251 (N_4251,N_3516,N_3836);
nor U4252 (N_4252,N_3445,N_3309);
and U4253 (N_4253,N_3743,N_3074);
or U4254 (N_4254,N_3348,N_3993);
xor U4255 (N_4255,N_3749,N_3920);
xor U4256 (N_4256,N_3292,N_3128);
and U4257 (N_4257,N_3990,N_3874);
nor U4258 (N_4258,N_3765,N_3386);
and U4259 (N_4259,N_3872,N_3873);
nor U4260 (N_4260,N_3406,N_3404);
and U4261 (N_4261,N_3324,N_3788);
and U4262 (N_4262,N_3231,N_3999);
and U4263 (N_4263,N_3627,N_3761);
nor U4264 (N_4264,N_3878,N_3654);
or U4265 (N_4265,N_3104,N_3979);
and U4266 (N_4266,N_3123,N_3613);
nor U4267 (N_4267,N_3169,N_3151);
nor U4268 (N_4268,N_3166,N_3721);
or U4269 (N_4269,N_3968,N_3519);
and U4270 (N_4270,N_3127,N_3575);
or U4271 (N_4271,N_3759,N_3638);
or U4272 (N_4272,N_3508,N_3932);
or U4273 (N_4273,N_3549,N_3786);
nand U4274 (N_4274,N_3419,N_3719);
xor U4275 (N_4275,N_3717,N_3598);
or U4276 (N_4276,N_3422,N_3814);
and U4277 (N_4277,N_3846,N_3063);
xnor U4278 (N_4278,N_3523,N_3213);
or U4279 (N_4279,N_3752,N_3984);
and U4280 (N_4280,N_3668,N_3870);
xor U4281 (N_4281,N_3758,N_3849);
nand U4282 (N_4282,N_3229,N_3407);
and U4283 (N_4283,N_3145,N_3056);
or U4284 (N_4284,N_3387,N_3255);
or U4285 (N_4285,N_3727,N_3152);
or U4286 (N_4286,N_3504,N_3349);
xnor U4287 (N_4287,N_3738,N_3626);
and U4288 (N_4288,N_3468,N_3646);
nor U4289 (N_4289,N_3066,N_3805);
xor U4290 (N_4290,N_3399,N_3534);
or U4291 (N_4291,N_3858,N_3623);
nor U4292 (N_4292,N_3825,N_3763);
xor U4293 (N_4293,N_3897,N_3209);
nor U4294 (N_4294,N_3296,N_3936);
nand U4295 (N_4295,N_3608,N_3951);
nand U4296 (N_4296,N_3325,N_3197);
or U4297 (N_4297,N_3659,N_3736);
or U4298 (N_4298,N_3526,N_3954);
nand U4299 (N_4299,N_3003,N_3780);
nand U4300 (N_4300,N_3473,N_3578);
nor U4301 (N_4301,N_3564,N_3746);
and U4302 (N_4302,N_3110,N_3947);
or U4303 (N_4303,N_3371,N_3666);
nor U4304 (N_4304,N_3463,N_3547);
xnor U4305 (N_4305,N_3695,N_3856);
nand U4306 (N_4306,N_3126,N_3307);
or U4307 (N_4307,N_3816,N_3140);
nand U4308 (N_4308,N_3079,N_3009);
or U4309 (N_4309,N_3068,N_3093);
xor U4310 (N_4310,N_3669,N_3141);
or U4311 (N_4311,N_3414,N_3750);
or U4312 (N_4312,N_3067,N_3452);
or U4313 (N_4313,N_3433,N_3089);
nand U4314 (N_4314,N_3521,N_3732);
nor U4315 (N_4315,N_3698,N_3579);
xor U4316 (N_4316,N_3827,N_3898);
nand U4317 (N_4317,N_3420,N_3259);
or U4318 (N_4318,N_3340,N_3138);
xnor U4319 (N_4319,N_3132,N_3423);
nor U4320 (N_4320,N_3052,N_3014);
xor U4321 (N_4321,N_3531,N_3212);
xor U4322 (N_4322,N_3527,N_3655);
xnor U4323 (N_4323,N_3829,N_3200);
xnor U4324 (N_4324,N_3194,N_3931);
or U4325 (N_4325,N_3593,N_3697);
nor U4326 (N_4326,N_3248,N_3821);
and U4327 (N_4327,N_3040,N_3206);
and U4328 (N_4328,N_3396,N_3866);
or U4329 (N_4329,N_3480,N_3970);
or U4330 (N_4330,N_3760,N_3991);
xnor U4331 (N_4331,N_3202,N_3879);
xnor U4332 (N_4332,N_3171,N_3944);
nor U4333 (N_4333,N_3902,N_3850);
and U4334 (N_4334,N_3026,N_3291);
and U4335 (N_4335,N_3237,N_3834);
and U4336 (N_4336,N_3939,N_3487);
nand U4337 (N_4337,N_3915,N_3657);
and U4338 (N_4338,N_3313,N_3381);
nor U4339 (N_4339,N_3442,N_3065);
xor U4340 (N_4340,N_3368,N_3673);
nor U4341 (N_4341,N_3995,N_3149);
nor U4342 (N_4342,N_3581,N_3446);
and U4343 (N_4343,N_3285,N_3082);
nand U4344 (N_4344,N_3105,N_3554);
and U4345 (N_4345,N_3624,N_3260);
nand U4346 (N_4346,N_3908,N_3670);
or U4347 (N_4347,N_3327,N_3600);
and U4348 (N_4348,N_3573,N_3426);
or U4349 (N_4349,N_3807,N_3852);
and U4350 (N_4350,N_3684,N_3416);
nor U4351 (N_4351,N_3147,N_3436);
nand U4352 (N_4352,N_3167,N_3784);
xor U4353 (N_4353,N_3022,N_3222);
nor U4354 (N_4354,N_3507,N_3921);
nand U4355 (N_4355,N_3397,N_3320);
and U4356 (N_4356,N_3637,N_3460);
xor U4357 (N_4357,N_3876,N_3569);
or U4358 (N_4358,N_3483,N_3813);
xnor U4359 (N_4359,N_3211,N_3017);
and U4360 (N_4360,N_3863,N_3091);
or U4361 (N_4361,N_3571,N_3612);
and U4362 (N_4362,N_3867,N_3892);
and U4363 (N_4363,N_3730,N_3687);
nor U4364 (N_4364,N_3405,N_3135);
or U4365 (N_4365,N_3032,N_3905);
xnor U4366 (N_4366,N_3020,N_3601);
and U4367 (N_4367,N_3466,N_3868);
or U4368 (N_4368,N_3747,N_3855);
and U4369 (N_4369,N_3893,N_3881);
nand U4370 (N_4370,N_3280,N_3023);
or U4371 (N_4371,N_3117,N_3679);
and U4372 (N_4372,N_3031,N_3678);
nand U4373 (N_4373,N_3261,N_3716);
or U4374 (N_4374,N_3098,N_3000);
and U4375 (N_4375,N_3592,N_3239);
xor U4376 (N_4376,N_3648,N_3540);
nor U4377 (N_4377,N_3227,N_3193);
xor U4378 (N_4378,N_3286,N_3517);
and U4379 (N_4379,N_3842,N_3819);
xnor U4380 (N_4380,N_3640,N_3242);
nor U4381 (N_4381,N_3810,N_3558);
nand U4382 (N_4382,N_3771,N_3860);
or U4383 (N_4383,N_3491,N_3220);
nor U4384 (N_4384,N_3244,N_3631);
nand U4385 (N_4385,N_3930,N_3048);
xnor U4386 (N_4386,N_3689,N_3013);
or U4387 (N_4387,N_3018,N_3390);
or U4388 (N_4388,N_3625,N_3162);
nor U4389 (N_4389,N_3001,N_3567);
and U4390 (N_4390,N_3887,N_3714);
nor U4391 (N_4391,N_3570,N_3099);
and U4392 (N_4392,N_3165,N_3488);
nor U4393 (N_4393,N_3262,N_3005);
nor U4394 (N_4394,N_3783,N_3055);
and U4395 (N_4395,N_3341,N_3376);
nor U4396 (N_4396,N_3645,N_3974);
nor U4397 (N_4397,N_3831,N_3533);
xnor U4398 (N_4398,N_3224,N_3775);
or U4399 (N_4399,N_3595,N_3987);
nor U4400 (N_4400,N_3275,N_3154);
or U4401 (N_4401,N_3899,N_3694);
and U4402 (N_4402,N_3330,N_3859);
and U4403 (N_4403,N_3797,N_3060);
and U4404 (N_4404,N_3676,N_3701);
nand U4405 (N_4405,N_3238,N_3494);
nand U4406 (N_4406,N_3808,N_3506);
and U4407 (N_4407,N_3326,N_3597);
xor U4408 (N_4408,N_3594,N_3228);
or U4409 (N_4409,N_3337,N_3424);
xnor U4410 (N_4410,N_3119,N_3053);
and U4411 (N_4411,N_3501,N_3455);
xor U4412 (N_4412,N_3156,N_3234);
and U4413 (N_4413,N_3339,N_3125);
or U4414 (N_4414,N_3782,N_3233);
nand U4415 (N_4415,N_3909,N_3215);
nor U4416 (N_4416,N_3711,N_3568);
and U4417 (N_4417,N_3470,N_3548);
and U4418 (N_4418,N_3116,N_3522);
nor U4419 (N_4419,N_3705,N_3373);
and U4420 (N_4420,N_3106,N_3590);
or U4421 (N_4421,N_3484,N_3266);
and U4422 (N_4422,N_3869,N_3946);
xor U4423 (N_4423,N_3582,N_3606);
or U4424 (N_4424,N_3310,N_3610);
and U4425 (N_4425,N_3159,N_3477);
nor U4426 (N_4426,N_3882,N_3195);
xor U4427 (N_4427,N_3933,N_3191);
and U4428 (N_4428,N_3394,N_3365);
or U4429 (N_4429,N_3462,N_3256);
nand U4430 (N_4430,N_3425,N_3342);
xnor U4431 (N_4431,N_3465,N_3817);
nand U4432 (N_4432,N_3643,N_3992);
xor U4433 (N_4433,N_3875,N_3070);
and U4434 (N_4434,N_3525,N_3085);
and U4435 (N_4435,N_3973,N_3837);
nand U4436 (N_4436,N_3130,N_3576);
nor U4437 (N_4437,N_3258,N_3174);
and U4438 (N_4438,N_3263,N_3064);
and U4439 (N_4439,N_3778,N_3900);
nor U4440 (N_4440,N_3617,N_3907);
and U4441 (N_4441,N_3049,N_3273);
nand U4442 (N_4442,N_3609,N_3781);
xnor U4443 (N_4443,N_3497,N_3948);
and U4444 (N_4444,N_3346,N_3981);
xnor U4445 (N_4445,N_3251,N_3566);
and U4446 (N_4446,N_3430,N_3641);
and U4447 (N_4447,N_3802,N_3182);
nor U4448 (N_4448,N_3375,N_3312);
nor U4449 (N_4449,N_3457,N_3585);
nor U4450 (N_4450,N_3652,N_3545);
nor U4451 (N_4451,N_3367,N_3583);
nor U4452 (N_4452,N_3439,N_3401);
nor U4453 (N_4453,N_3550,N_3704);
nor U4454 (N_4454,N_3051,N_3647);
nand U4455 (N_4455,N_3619,N_3268);
nor U4456 (N_4456,N_3164,N_3621);
nand U4457 (N_4457,N_3847,N_3448);
nand U4458 (N_4458,N_3804,N_3335);
or U4459 (N_4459,N_3812,N_3977);
xnor U4460 (N_4460,N_3672,N_3886);
nand U4461 (N_4461,N_3725,N_3447);
and U4462 (N_4462,N_3644,N_3358);
and U4463 (N_4463,N_3136,N_3092);
or U4464 (N_4464,N_3357,N_3833);
xor U4465 (N_4465,N_3402,N_3917);
nand U4466 (N_4466,N_3806,N_3629);
or U4467 (N_4467,N_3877,N_3077);
or U4468 (N_4468,N_3277,N_3437);
nor U4469 (N_4469,N_3696,N_3495);
nand U4470 (N_4470,N_3500,N_3021);
and U4471 (N_4471,N_3692,N_3890);
nand U4472 (N_4472,N_3851,N_3057);
nor U4473 (N_4473,N_3492,N_3832);
nand U4474 (N_4474,N_3006,N_3185);
xnor U4475 (N_4475,N_3243,N_3461);
and U4476 (N_4476,N_3355,N_3742);
xor U4477 (N_4477,N_3630,N_3733);
xor U4478 (N_4478,N_3471,N_3707);
nor U4479 (N_4479,N_3353,N_3252);
and U4480 (N_4480,N_3767,N_3756);
and U4481 (N_4481,N_3541,N_3632);
or U4482 (N_4482,N_3634,N_3272);
xor U4483 (N_4483,N_3818,N_3108);
or U4484 (N_4484,N_3059,N_3703);
nor U4485 (N_4485,N_3822,N_3336);
nor U4486 (N_4486,N_3934,N_3331);
nand U4487 (N_4487,N_3412,N_3803);
or U4488 (N_4488,N_3004,N_3181);
and U4489 (N_4489,N_3949,N_3450);
xnor U4490 (N_4490,N_3754,N_3511);
xnor U4491 (N_4491,N_3038,N_3577);
nand U4492 (N_4492,N_3751,N_3289);
nor U4493 (N_4493,N_3478,N_3616);
and U4494 (N_4494,N_3333,N_3912);
nand U4495 (N_4495,N_3764,N_3734);
and U4496 (N_4496,N_3037,N_3050);
nor U4497 (N_4497,N_3047,N_3955);
and U4498 (N_4498,N_3134,N_3007);
and U4499 (N_4499,N_3663,N_3356);
xnor U4500 (N_4500,N_3514,N_3570);
nand U4501 (N_4501,N_3011,N_3679);
xnor U4502 (N_4502,N_3272,N_3987);
nor U4503 (N_4503,N_3950,N_3945);
nor U4504 (N_4504,N_3248,N_3437);
nand U4505 (N_4505,N_3886,N_3242);
and U4506 (N_4506,N_3980,N_3913);
nor U4507 (N_4507,N_3185,N_3638);
and U4508 (N_4508,N_3413,N_3689);
and U4509 (N_4509,N_3696,N_3924);
or U4510 (N_4510,N_3413,N_3524);
and U4511 (N_4511,N_3708,N_3359);
and U4512 (N_4512,N_3373,N_3633);
and U4513 (N_4513,N_3838,N_3620);
nor U4514 (N_4514,N_3956,N_3017);
or U4515 (N_4515,N_3181,N_3936);
nor U4516 (N_4516,N_3901,N_3052);
xor U4517 (N_4517,N_3177,N_3716);
or U4518 (N_4518,N_3214,N_3752);
xnor U4519 (N_4519,N_3486,N_3206);
nand U4520 (N_4520,N_3716,N_3382);
or U4521 (N_4521,N_3161,N_3119);
nor U4522 (N_4522,N_3854,N_3222);
xor U4523 (N_4523,N_3904,N_3223);
or U4524 (N_4524,N_3020,N_3479);
nand U4525 (N_4525,N_3087,N_3323);
xor U4526 (N_4526,N_3528,N_3072);
nor U4527 (N_4527,N_3307,N_3267);
or U4528 (N_4528,N_3067,N_3888);
nor U4529 (N_4529,N_3914,N_3575);
or U4530 (N_4530,N_3736,N_3300);
nand U4531 (N_4531,N_3069,N_3015);
xor U4532 (N_4532,N_3429,N_3536);
nand U4533 (N_4533,N_3087,N_3818);
xnor U4534 (N_4534,N_3885,N_3752);
or U4535 (N_4535,N_3824,N_3821);
and U4536 (N_4536,N_3006,N_3864);
nand U4537 (N_4537,N_3300,N_3171);
and U4538 (N_4538,N_3317,N_3123);
or U4539 (N_4539,N_3273,N_3459);
xor U4540 (N_4540,N_3039,N_3803);
or U4541 (N_4541,N_3260,N_3598);
or U4542 (N_4542,N_3509,N_3628);
or U4543 (N_4543,N_3306,N_3249);
or U4544 (N_4544,N_3880,N_3594);
xnor U4545 (N_4545,N_3691,N_3835);
or U4546 (N_4546,N_3596,N_3572);
nand U4547 (N_4547,N_3548,N_3481);
and U4548 (N_4548,N_3657,N_3458);
nor U4549 (N_4549,N_3347,N_3069);
and U4550 (N_4550,N_3509,N_3861);
and U4551 (N_4551,N_3681,N_3302);
nand U4552 (N_4552,N_3612,N_3157);
and U4553 (N_4553,N_3400,N_3937);
and U4554 (N_4554,N_3228,N_3218);
xor U4555 (N_4555,N_3011,N_3407);
or U4556 (N_4556,N_3017,N_3190);
and U4557 (N_4557,N_3086,N_3064);
nor U4558 (N_4558,N_3438,N_3179);
and U4559 (N_4559,N_3489,N_3890);
and U4560 (N_4560,N_3699,N_3334);
or U4561 (N_4561,N_3968,N_3729);
or U4562 (N_4562,N_3521,N_3108);
and U4563 (N_4563,N_3208,N_3223);
or U4564 (N_4564,N_3470,N_3289);
nand U4565 (N_4565,N_3145,N_3341);
xor U4566 (N_4566,N_3901,N_3758);
and U4567 (N_4567,N_3705,N_3361);
or U4568 (N_4568,N_3698,N_3427);
nand U4569 (N_4569,N_3387,N_3542);
nor U4570 (N_4570,N_3449,N_3886);
xor U4571 (N_4571,N_3850,N_3465);
xor U4572 (N_4572,N_3394,N_3161);
xnor U4573 (N_4573,N_3878,N_3489);
nand U4574 (N_4574,N_3253,N_3633);
nand U4575 (N_4575,N_3106,N_3568);
xor U4576 (N_4576,N_3835,N_3951);
xor U4577 (N_4577,N_3398,N_3722);
xnor U4578 (N_4578,N_3679,N_3587);
nand U4579 (N_4579,N_3342,N_3357);
nor U4580 (N_4580,N_3216,N_3114);
nor U4581 (N_4581,N_3594,N_3460);
nand U4582 (N_4582,N_3920,N_3589);
or U4583 (N_4583,N_3313,N_3897);
nor U4584 (N_4584,N_3518,N_3509);
and U4585 (N_4585,N_3113,N_3233);
nor U4586 (N_4586,N_3742,N_3806);
nand U4587 (N_4587,N_3305,N_3531);
nand U4588 (N_4588,N_3810,N_3615);
and U4589 (N_4589,N_3166,N_3402);
nand U4590 (N_4590,N_3867,N_3362);
xnor U4591 (N_4591,N_3273,N_3842);
nand U4592 (N_4592,N_3707,N_3338);
xor U4593 (N_4593,N_3451,N_3645);
and U4594 (N_4594,N_3361,N_3588);
and U4595 (N_4595,N_3285,N_3988);
and U4596 (N_4596,N_3226,N_3342);
nor U4597 (N_4597,N_3901,N_3296);
nor U4598 (N_4598,N_3099,N_3386);
nand U4599 (N_4599,N_3561,N_3767);
or U4600 (N_4600,N_3127,N_3934);
and U4601 (N_4601,N_3824,N_3289);
xor U4602 (N_4602,N_3415,N_3224);
or U4603 (N_4603,N_3690,N_3337);
nor U4604 (N_4604,N_3404,N_3249);
nor U4605 (N_4605,N_3096,N_3785);
xnor U4606 (N_4606,N_3111,N_3932);
or U4607 (N_4607,N_3994,N_3770);
nor U4608 (N_4608,N_3856,N_3072);
nand U4609 (N_4609,N_3536,N_3161);
and U4610 (N_4610,N_3472,N_3123);
nand U4611 (N_4611,N_3243,N_3776);
nor U4612 (N_4612,N_3061,N_3980);
nand U4613 (N_4613,N_3081,N_3354);
nor U4614 (N_4614,N_3153,N_3974);
xnor U4615 (N_4615,N_3981,N_3616);
nor U4616 (N_4616,N_3212,N_3402);
xnor U4617 (N_4617,N_3182,N_3814);
or U4618 (N_4618,N_3528,N_3674);
nor U4619 (N_4619,N_3401,N_3453);
nand U4620 (N_4620,N_3612,N_3274);
or U4621 (N_4621,N_3219,N_3149);
nor U4622 (N_4622,N_3745,N_3672);
or U4623 (N_4623,N_3183,N_3857);
nand U4624 (N_4624,N_3435,N_3945);
and U4625 (N_4625,N_3359,N_3241);
or U4626 (N_4626,N_3639,N_3723);
or U4627 (N_4627,N_3983,N_3598);
nand U4628 (N_4628,N_3662,N_3898);
nand U4629 (N_4629,N_3011,N_3211);
xnor U4630 (N_4630,N_3883,N_3427);
nor U4631 (N_4631,N_3504,N_3207);
and U4632 (N_4632,N_3125,N_3874);
xnor U4633 (N_4633,N_3836,N_3306);
xnor U4634 (N_4634,N_3191,N_3073);
and U4635 (N_4635,N_3030,N_3357);
nor U4636 (N_4636,N_3721,N_3143);
nand U4637 (N_4637,N_3969,N_3949);
xnor U4638 (N_4638,N_3089,N_3779);
or U4639 (N_4639,N_3876,N_3029);
nand U4640 (N_4640,N_3648,N_3913);
nor U4641 (N_4641,N_3140,N_3105);
nor U4642 (N_4642,N_3385,N_3012);
xnor U4643 (N_4643,N_3559,N_3406);
or U4644 (N_4644,N_3906,N_3742);
and U4645 (N_4645,N_3867,N_3057);
or U4646 (N_4646,N_3930,N_3093);
xor U4647 (N_4647,N_3461,N_3812);
and U4648 (N_4648,N_3753,N_3383);
nand U4649 (N_4649,N_3946,N_3762);
nor U4650 (N_4650,N_3078,N_3792);
and U4651 (N_4651,N_3111,N_3952);
or U4652 (N_4652,N_3163,N_3796);
nor U4653 (N_4653,N_3557,N_3595);
xor U4654 (N_4654,N_3939,N_3326);
xor U4655 (N_4655,N_3045,N_3799);
xor U4656 (N_4656,N_3056,N_3569);
nor U4657 (N_4657,N_3064,N_3239);
or U4658 (N_4658,N_3166,N_3943);
or U4659 (N_4659,N_3936,N_3449);
nor U4660 (N_4660,N_3888,N_3947);
nor U4661 (N_4661,N_3558,N_3826);
and U4662 (N_4662,N_3523,N_3114);
or U4663 (N_4663,N_3862,N_3296);
and U4664 (N_4664,N_3329,N_3946);
nor U4665 (N_4665,N_3613,N_3966);
nor U4666 (N_4666,N_3545,N_3489);
nor U4667 (N_4667,N_3859,N_3840);
nor U4668 (N_4668,N_3560,N_3896);
xor U4669 (N_4669,N_3157,N_3416);
and U4670 (N_4670,N_3498,N_3426);
nand U4671 (N_4671,N_3916,N_3624);
xnor U4672 (N_4672,N_3601,N_3776);
xor U4673 (N_4673,N_3115,N_3584);
and U4674 (N_4674,N_3907,N_3198);
xor U4675 (N_4675,N_3324,N_3189);
xnor U4676 (N_4676,N_3552,N_3138);
and U4677 (N_4677,N_3399,N_3850);
nand U4678 (N_4678,N_3881,N_3094);
or U4679 (N_4679,N_3233,N_3414);
nand U4680 (N_4680,N_3232,N_3208);
or U4681 (N_4681,N_3463,N_3917);
or U4682 (N_4682,N_3949,N_3056);
and U4683 (N_4683,N_3120,N_3864);
or U4684 (N_4684,N_3598,N_3557);
xor U4685 (N_4685,N_3720,N_3317);
nor U4686 (N_4686,N_3199,N_3641);
nor U4687 (N_4687,N_3611,N_3931);
or U4688 (N_4688,N_3178,N_3308);
nand U4689 (N_4689,N_3989,N_3229);
or U4690 (N_4690,N_3916,N_3936);
or U4691 (N_4691,N_3551,N_3030);
nand U4692 (N_4692,N_3793,N_3606);
nor U4693 (N_4693,N_3847,N_3899);
xnor U4694 (N_4694,N_3074,N_3318);
xor U4695 (N_4695,N_3678,N_3478);
or U4696 (N_4696,N_3672,N_3931);
nand U4697 (N_4697,N_3845,N_3669);
nand U4698 (N_4698,N_3734,N_3469);
or U4699 (N_4699,N_3498,N_3545);
or U4700 (N_4700,N_3724,N_3632);
nor U4701 (N_4701,N_3982,N_3724);
nor U4702 (N_4702,N_3411,N_3899);
and U4703 (N_4703,N_3348,N_3140);
nand U4704 (N_4704,N_3143,N_3101);
or U4705 (N_4705,N_3580,N_3787);
nor U4706 (N_4706,N_3862,N_3018);
nor U4707 (N_4707,N_3774,N_3869);
and U4708 (N_4708,N_3882,N_3833);
or U4709 (N_4709,N_3018,N_3204);
nor U4710 (N_4710,N_3353,N_3806);
xnor U4711 (N_4711,N_3900,N_3750);
nand U4712 (N_4712,N_3277,N_3322);
xor U4713 (N_4713,N_3173,N_3162);
nor U4714 (N_4714,N_3540,N_3785);
nand U4715 (N_4715,N_3107,N_3940);
nand U4716 (N_4716,N_3693,N_3809);
nor U4717 (N_4717,N_3919,N_3372);
nand U4718 (N_4718,N_3242,N_3286);
xnor U4719 (N_4719,N_3076,N_3037);
nand U4720 (N_4720,N_3080,N_3598);
and U4721 (N_4721,N_3938,N_3234);
nor U4722 (N_4722,N_3802,N_3185);
xnor U4723 (N_4723,N_3022,N_3973);
nand U4724 (N_4724,N_3567,N_3891);
nand U4725 (N_4725,N_3087,N_3545);
xnor U4726 (N_4726,N_3955,N_3667);
xor U4727 (N_4727,N_3001,N_3108);
nand U4728 (N_4728,N_3860,N_3690);
and U4729 (N_4729,N_3556,N_3548);
nand U4730 (N_4730,N_3308,N_3858);
or U4731 (N_4731,N_3763,N_3270);
nor U4732 (N_4732,N_3043,N_3774);
or U4733 (N_4733,N_3050,N_3084);
xnor U4734 (N_4734,N_3640,N_3585);
nand U4735 (N_4735,N_3039,N_3306);
and U4736 (N_4736,N_3286,N_3597);
and U4737 (N_4737,N_3874,N_3097);
or U4738 (N_4738,N_3598,N_3920);
nor U4739 (N_4739,N_3620,N_3801);
nand U4740 (N_4740,N_3930,N_3386);
xor U4741 (N_4741,N_3768,N_3838);
and U4742 (N_4742,N_3516,N_3299);
nand U4743 (N_4743,N_3307,N_3873);
nor U4744 (N_4744,N_3579,N_3400);
xnor U4745 (N_4745,N_3027,N_3831);
nand U4746 (N_4746,N_3880,N_3424);
and U4747 (N_4747,N_3343,N_3058);
xor U4748 (N_4748,N_3945,N_3449);
or U4749 (N_4749,N_3157,N_3606);
nand U4750 (N_4750,N_3645,N_3193);
nand U4751 (N_4751,N_3453,N_3473);
nor U4752 (N_4752,N_3124,N_3446);
and U4753 (N_4753,N_3110,N_3391);
xor U4754 (N_4754,N_3611,N_3056);
nor U4755 (N_4755,N_3905,N_3458);
and U4756 (N_4756,N_3909,N_3324);
or U4757 (N_4757,N_3602,N_3322);
nor U4758 (N_4758,N_3101,N_3090);
nor U4759 (N_4759,N_3708,N_3536);
and U4760 (N_4760,N_3800,N_3280);
nand U4761 (N_4761,N_3744,N_3176);
or U4762 (N_4762,N_3963,N_3968);
nor U4763 (N_4763,N_3110,N_3496);
nand U4764 (N_4764,N_3446,N_3517);
nand U4765 (N_4765,N_3403,N_3747);
and U4766 (N_4766,N_3093,N_3595);
xor U4767 (N_4767,N_3195,N_3350);
nor U4768 (N_4768,N_3900,N_3867);
nand U4769 (N_4769,N_3429,N_3018);
xor U4770 (N_4770,N_3387,N_3226);
and U4771 (N_4771,N_3090,N_3338);
or U4772 (N_4772,N_3646,N_3471);
and U4773 (N_4773,N_3580,N_3027);
and U4774 (N_4774,N_3393,N_3037);
nor U4775 (N_4775,N_3972,N_3448);
and U4776 (N_4776,N_3161,N_3378);
nor U4777 (N_4777,N_3311,N_3297);
xnor U4778 (N_4778,N_3905,N_3866);
nor U4779 (N_4779,N_3142,N_3794);
nand U4780 (N_4780,N_3881,N_3426);
or U4781 (N_4781,N_3598,N_3144);
and U4782 (N_4782,N_3810,N_3535);
or U4783 (N_4783,N_3970,N_3199);
xnor U4784 (N_4784,N_3834,N_3958);
nand U4785 (N_4785,N_3637,N_3372);
nor U4786 (N_4786,N_3396,N_3116);
or U4787 (N_4787,N_3305,N_3772);
and U4788 (N_4788,N_3875,N_3679);
and U4789 (N_4789,N_3001,N_3663);
or U4790 (N_4790,N_3211,N_3805);
nand U4791 (N_4791,N_3408,N_3117);
or U4792 (N_4792,N_3916,N_3843);
nand U4793 (N_4793,N_3668,N_3370);
and U4794 (N_4794,N_3964,N_3415);
nor U4795 (N_4795,N_3553,N_3843);
and U4796 (N_4796,N_3465,N_3413);
xnor U4797 (N_4797,N_3561,N_3936);
nor U4798 (N_4798,N_3844,N_3533);
and U4799 (N_4799,N_3973,N_3255);
nand U4800 (N_4800,N_3405,N_3634);
nand U4801 (N_4801,N_3889,N_3981);
or U4802 (N_4802,N_3764,N_3686);
and U4803 (N_4803,N_3363,N_3154);
nor U4804 (N_4804,N_3041,N_3339);
or U4805 (N_4805,N_3325,N_3434);
xor U4806 (N_4806,N_3606,N_3756);
nor U4807 (N_4807,N_3917,N_3297);
or U4808 (N_4808,N_3981,N_3090);
nand U4809 (N_4809,N_3147,N_3211);
and U4810 (N_4810,N_3056,N_3625);
or U4811 (N_4811,N_3632,N_3390);
nand U4812 (N_4812,N_3159,N_3635);
nor U4813 (N_4813,N_3444,N_3566);
and U4814 (N_4814,N_3790,N_3314);
nand U4815 (N_4815,N_3057,N_3166);
nor U4816 (N_4816,N_3256,N_3743);
nor U4817 (N_4817,N_3953,N_3429);
or U4818 (N_4818,N_3410,N_3432);
nand U4819 (N_4819,N_3375,N_3948);
and U4820 (N_4820,N_3215,N_3811);
and U4821 (N_4821,N_3712,N_3459);
nor U4822 (N_4822,N_3071,N_3479);
or U4823 (N_4823,N_3165,N_3744);
or U4824 (N_4824,N_3273,N_3238);
nand U4825 (N_4825,N_3527,N_3647);
and U4826 (N_4826,N_3987,N_3423);
or U4827 (N_4827,N_3036,N_3697);
xnor U4828 (N_4828,N_3789,N_3696);
and U4829 (N_4829,N_3643,N_3360);
or U4830 (N_4830,N_3878,N_3349);
nor U4831 (N_4831,N_3308,N_3216);
nor U4832 (N_4832,N_3636,N_3578);
xor U4833 (N_4833,N_3135,N_3751);
xor U4834 (N_4834,N_3571,N_3819);
nor U4835 (N_4835,N_3583,N_3857);
nand U4836 (N_4836,N_3736,N_3481);
nor U4837 (N_4837,N_3725,N_3297);
xor U4838 (N_4838,N_3021,N_3418);
or U4839 (N_4839,N_3815,N_3928);
xnor U4840 (N_4840,N_3175,N_3795);
nand U4841 (N_4841,N_3053,N_3689);
nor U4842 (N_4842,N_3152,N_3642);
xor U4843 (N_4843,N_3708,N_3394);
nor U4844 (N_4844,N_3900,N_3958);
nand U4845 (N_4845,N_3794,N_3055);
nor U4846 (N_4846,N_3889,N_3924);
xnor U4847 (N_4847,N_3595,N_3262);
nor U4848 (N_4848,N_3871,N_3955);
and U4849 (N_4849,N_3957,N_3049);
nor U4850 (N_4850,N_3728,N_3531);
or U4851 (N_4851,N_3971,N_3055);
and U4852 (N_4852,N_3049,N_3366);
nand U4853 (N_4853,N_3406,N_3382);
nand U4854 (N_4854,N_3300,N_3581);
nor U4855 (N_4855,N_3940,N_3501);
and U4856 (N_4856,N_3596,N_3524);
xnor U4857 (N_4857,N_3300,N_3084);
or U4858 (N_4858,N_3688,N_3325);
xor U4859 (N_4859,N_3634,N_3722);
xnor U4860 (N_4860,N_3675,N_3678);
and U4861 (N_4861,N_3868,N_3857);
or U4862 (N_4862,N_3086,N_3526);
and U4863 (N_4863,N_3682,N_3405);
nor U4864 (N_4864,N_3399,N_3504);
nand U4865 (N_4865,N_3390,N_3872);
nand U4866 (N_4866,N_3398,N_3377);
and U4867 (N_4867,N_3207,N_3663);
and U4868 (N_4868,N_3392,N_3429);
or U4869 (N_4869,N_3269,N_3026);
xnor U4870 (N_4870,N_3805,N_3099);
xor U4871 (N_4871,N_3919,N_3369);
nor U4872 (N_4872,N_3833,N_3892);
and U4873 (N_4873,N_3575,N_3809);
or U4874 (N_4874,N_3412,N_3040);
and U4875 (N_4875,N_3173,N_3644);
xnor U4876 (N_4876,N_3071,N_3817);
xor U4877 (N_4877,N_3510,N_3412);
or U4878 (N_4878,N_3384,N_3211);
or U4879 (N_4879,N_3460,N_3770);
nand U4880 (N_4880,N_3119,N_3530);
and U4881 (N_4881,N_3498,N_3248);
nand U4882 (N_4882,N_3326,N_3501);
nor U4883 (N_4883,N_3819,N_3831);
or U4884 (N_4884,N_3305,N_3579);
nor U4885 (N_4885,N_3954,N_3740);
or U4886 (N_4886,N_3438,N_3105);
nand U4887 (N_4887,N_3106,N_3723);
or U4888 (N_4888,N_3237,N_3429);
xor U4889 (N_4889,N_3679,N_3878);
nand U4890 (N_4890,N_3554,N_3439);
or U4891 (N_4891,N_3775,N_3924);
nor U4892 (N_4892,N_3641,N_3876);
or U4893 (N_4893,N_3137,N_3831);
and U4894 (N_4894,N_3723,N_3705);
xnor U4895 (N_4895,N_3281,N_3217);
or U4896 (N_4896,N_3674,N_3826);
or U4897 (N_4897,N_3372,N_3739);
nor U4898 (N_4898,N_3651,N_3578);
or U4899 (N_4899,N_3710,N_3112);
nand U4900 (N_4900,N_3455,N_3391);
and U4901 (N_4901,N_3837,N_3410);
or U4902 (N_4902,N_3553,N_3103);
or U4903 (N_4903,N_3419,N_3827);
nand U4904 (N_4904,N_3329,N_3992);
or U4905 (N_4905,N_3031,N_3780);
nor U4906 (N_4906,N_3033,N_3836);
xor U4907 (N_4907,N_3281,N_3193);
nor U4908 (N_4908,N_3803,N_3275);
and U4909 (N_4909,N_3591,N_3600);
or U4910 (N_4910,N_3458,N_3800);
or U4911 (N_4911,N_3398,N_3277);
nand U4912 (N_4912,N_3158,N_3431);
or U4913 (N_4913,N_3318,N_3919);
and U4914 (N_4914,N_3201,N_3222);
nand U4915 (N_4915,N_3960,N_3130);
nand U4916 (N_4916,N_3978,N_3862);
and U4917 (N_4917,N_3468,N_3480);
and U4918 (N_4918,N_3742,N_3300);
or U4919 (N_4919,N_3752,N_3811);
nand U4920 (N_4920,N_3763,N_3744);
xnor U4921 (N_4921,N_3334,N_3727);
nor U4922 (N_4922,N_3643,N_3700);
and U4923 (N_4923,N_3805,N_3961);
nand U4924 (N_4924,N_3871,N_3841);
nor U4925 (N_4925,N_3200,N_3886);
and U4926 (N_4926,N_3945,N_3396);
and U4927 (N_4927,N_3494,N_3239);
and U4928 (N_4928,N_3929,N_3912);
nand U4929 (N_4929,N_3390,N_3623);
nor U4930 (N_4930,N_3554,N_3612);
nand U4931 (N_4931,N_3062,N_3311);
xor U4932 (N_4932,N_3207,N_3336);
nand U4933 (N_4933,N_3888,N_3446);
xnor U4934 (N_4934,N_3448,N_3362);
nand U4935 (N_4935,N_3550,N_3571);
or U4936 (N_4936,N_3374,N_3144);
xnor U4937 (N_4937,N_3397,N_3403);
nand U4938 (N_4938,N_3741,N_3438);
xnor U4939 (N_4939,N_3424,N_3786);
or U4940 (N_4940,N_3296,N_3628);
nor U4941 (N_4941,N_3948,N_3169);
xor U4942 (N_4942,N_3192,N_3118);
and U4943 (N_4943,N_3988,N_3659);
nor U4944 (N_4944,N_3754,N_3073);
xor U4945 (N_4945,N_3744,N_3316);
and U4946 (N_4946,N_3814,N_3605);
nand U4947 (N_4947,N_3427,N_3187);
nand U4948 (N_4948,N_3710,N_3073);
nand U4949 (N_4949,N_3959,N_3679);
nand U4950 (N_4950,N_3630,N_3529);
and U4951 (N_4951,N_3690,N_3523);
nand U4952 (N_4952,N_3957,N_3747);
nor U4953 (N_4953,N_3605,N_3397);
nor U4954 (N_4954,N_3082,N_3696);
nand U4955 (N_4955,N_3607,N_3176);
xor U4956 (N_4956,N_3024,N_3259);
xor U4957 (N_4957,N_3661,N_3730);
nand U4958 (N_4958,N_3249,N_3187);
xnor U4959 (N_4959,N_3551,N_3072);
and U4960 (N_4960,N_3285,N_3408);
xor U4961 (N_4961,N_3340,N_3188);
nor U4962 (N_4962,N_3354,N_3698);
or U4963 (N_4963,N_3731,N_3089);
or U4964 (N_4964,N_3289,N_3967);
xnor U4965 (N_4965,N_3568,N_3505);
xnor U4966 (N_4966,N_3469,N_3833);
nand U4967 (N_4967,N_3897,N_3584);
or U4968 (N_4968,N_3733,N_3648);
and U4969 (N_4969,N_3592,N_3475);
xor U4970 (N_4970,N_3853,N_3142);
or U4971 (N_4971,N_3168,N_3997);
nand U4972 (N_4972,N_3245,N_3066);
or U4973 (N_4973,N_3028,N_3293);
nor U4974 (N_4974,N_3617,N_3432);
and U4975 (N_4975,N_3941,N_3308);
or U4976 (N_4976,N_3537,N_3984);
nand U4977 (N_4977,N_3194,N_3260);
and U4978 (N_4978,N_3239,N_3128);
nand U4979 (N_4979,N_3568,N_3343);
or U4980 (N_4980,N_3913,N_3684);
or U4981 (N_4981,N_3021,N_3727);
or U4982 (N_4982,N_3052,N_3493);
xor U4983 (N_4983,N_3897,N_3630);
and U4984 (N_4984,N_3046,N_3611);
and U4985 (N_4985,N_3790,N_3442);
xnor U4986 (N_4986,N_3071,N_3506);
xor U4987 (N_4987,N_3424,N_3604);
xor U4988 (N_4988,N_3644,N_3899);
and U4989 (N_4989,N_3528,N_3773);
or U4990 (N_4990,N_3687,N_3012);
xor U4991 (N_4991,N_3111,N_3297);
xnor U4992 (N_4992,N_3067,N_3127);
or U4993 (N_4993,N_3907,N_3042);
nand U4994 (N_4994,N_3318,N_3681);
nand U4995 (N_4995,N_3706,N_3657);
nand U4996 (N_4996,N_3619,N_3040);
and U4997 (N_4997,N_3371,N_3448);
nand U4998 (N_4998,N_3722,N_3142);
and U4999 (N_4999,N_3190,N_3040);
xnor U5000 (N_5000,N_4801,N_4555);
or U5001 (N_5001,N_4293,N_4952);
nor U5002 (N_5002,N_4862,N_4027);
nand U5003 (N_5003,N_4846,N_4077);
nand U5004 (N_5004,N_4693,N_4354);
xnor U5005 (N_5005,N_4655,N_4026);
or U5006 (N_5006,N_4343,N_4116);
nand U5007 (N_5007,N_4521,N_4197);
nor U5008 (N_5008,N_4044,N_4134);
nor U5009 (N_5009,N_4471,N_4731);
nor U5010 (N_5010,N_4276,N_4468);
xnor U5011 (N_5011,N_4513,N_4737);
nor U5012 (N_5012,N_4664,N_4185);
and U5013 (N_5013,N_4921,N_4995);
xnor U5014 (N_5014,N_4297,N_4792);
or U5015 (N_5015,N_4182,N_4603);
nor U5016 (N_5016,N_4126,N_4873);
or U5017 (N_5017,N_4227,N_4331);
and U5018 (N_5018,N_4143,N_4071);
and U5019 (N_5019,N_4795,N_4807);
and U5020 (N_5020,N_4209,N_4761);
nand U5021 (N_5021,N_4606,N_4657);
or U5022 (N_5022,N_4759,N_4965);
and U5023 (N_5023,N_4022,N_4527);
xor U5024 (N_5024,N_4315,N_4696);
xnor U5025 (N_5025,N_4279,N_4475);
or U5026 (N_5026,N_4179,N_4740);
nor U5027 (N_5027,N_4100,N_4418);
nand U5028 (N_5028,N_4836,N_4734);
nand U5029 (N_5029,N_4887,N_4674);
nor U5030 (N_5030,N_4742,N_4114);
nor U5031 (N_5031,N_4955,N_4165);
or U5032 (N_5032,N_4913,N_4905);
nand U5033 (N_5033,N_4094,N_4281);
and U5034 (N_5034,N_4189,N_4849);
or U5035 (N_5035,N_4954,N_4081);
or U5036 (N_5036,N_4493,N_4469);
nand U5037 (N_5037,N_4098,N_4627);
nand U5038 (N_5038,N_4035,N_4864);
or U5039 (N_5039,N_4063,N_4308);
nand U5040 (N_5040,N_4250,N_4246);
nor U5041 (N_5041,N_4517,N_4167);
xnor U5042 (N_5042,N_4580,N_4534);
and U5043 (N_5043,N_4348,N_4973);
xor U5044 (N_5044,N_4295,N_4482);
nand U5045 (N_5045,N_4166,N_4728);
nand U5046 (N_5046,N_4856,N_4879);
nand U5047 (N_5047,N_4961,N_4816);
xnor U5048 (N_5048,N_4399,N_4918);
xnor U5049 (N_5049,N_4618,N_4249);
nor U5050 (N_5050,N_4712,N_4188);
and U5051 (N_5051,N_4679,N_4439);
nor U5052 (N_5052,N_4797,N_4611);
nor U5053 (N_5053,N_4200,N_4347);
and U5054 (N_5054,N_4813,N_4613);
nand U5055 (N_5055,N_4413,N_4902);
and U5056 (N_5056,N_4390,N_4445);
nor U5057 (N_5057,N_4457,N_4338);
or U5058 (N_5058,N_4421,N_4514);
nand U5059 (N_5059,N_4256,N_4144);
nand U5060 (N_5060,N_4097,N_4245);
nor U5061 (N_5061,N_4210,N_4670);
nor U5062 (N_5062,N_4556,N_4569);
nand U5063 (N_5063,N_4362,N_4841);
nor U5064 (N_5064,N_4205,N_4978);
and U5065 (N_5065,N_4560,N_4158);
nor U5066 (N_5066,N_4495,N_4830);
nand U5067 (N_5067,N_4812,N_4411);
or U5068 (N_5068,N_4883,N_4234);
xor U5069 (N_5069,N_4358,N_4191);
and U5070 (N_5070,N_4701,N_4275);
nand U5071 (N_5071,N_4659,N_4253);
nand U5072 (N_5072,N_4150,N_4003);
or U5073 (N_5073,N_4453,N_4239);
nor U5074 (N_5074,N_4298,N_4899);
or U5075 (N_5075,N_4401,N_4639);
or U5076 (N_5076,N_4083,N_4776);
or U5077 (N_5077,N_4842,N_4894);
xor U5078 (N_5078,N_4889,N_4643);
nor U5079 (N_5079,N_4435,N_4622);
and U5080 (N_5080,N_4199,N_4626);
and U5081 (N_5081,N_4156,N_4808);
or U5082 (N_5082,N_4079,N_4991);
or U5083 (N_5083,N_4443,N_4018);
nor U5084 (N_5084,N_4893,N_4789);
nor U5085 (N_5085,N_4703,N_4710);
nor U5086 (N_5086,N_4501,N_4406);
nand U5087 (N_5087,N_4178,N_4589);
nor U5088 (N_5088,N_4931,N_4715);
xnor U5089 (N_5089,N_4976,N_4845);
or U5090 (N_5090,N_4317,N_4516);
and U5091 (N_5091,N_4967,N_4168);
and U5092 (N_5092,N_4895,N_4775);
nand U5093 (N_5093,N_4780,N_4739);
xor U5094 (N_5094,N_4585,N_4290);
nand U5095 (N_5095,N_4711,N_4261);
xnor U5096 (N_5096,N_4029,N_4634);
and U5097 (N_5097,N_4751,N_4038);
or U5098 (N_5098,N_4650,N_4095);
xnor U5099 (N_5099,N_4070,N_4307);
xnor U5100 (N_5100,N_4654,N_4982);
xor U5101 (N_5101,N_4050,N_4912);
and U5102 (N_5102,N_4881,N_4184);
or U5103 (N_5103,N_4947,N_4053);
or U5104 (N_5104,N_4561,N_4377);
or U5105 (N_5105,N_4769,N_4535);
nand U5106 (N_5106,N_4624,N_4694);
nand U5107 (N_5107,N_4365,N_4272);
and U5108 (N_5108,N_4483,N_4638);
or U5109 (N_5109,N_4980,N_4882);
xor U5110 (N_5110,N_4481,N_4228);
or U5111 (N_5111,N_4571,N_4778);
nand U5112 (N_5112,N_4461,N_4419);
xnor U5113 (N_5113,N_4449,N_4758);
xnor U5114 (N_5114,N_4171,N_4202);
xnor U5115 (N_5115,N_4749,N_4819);
or U5116 (N_5116,N_4351,N_4215);
xor U5117 (N_5117,N_4875,N_4106);
nor U5118 (N_5118,N_4356,N_4099);
nor U5119 (N_5119,N_4832,N_4389);
xnor U5120 (N_5120,N_4366,N_4466);
xnor U5121 (N_5121,N_4426,N_4804);
nand U5122 (N_5122,N_4265,N_4970);
or U5123 (N_5123,N_4432,N_4262);
or U5124 (N_5124,N_4266,N_4798);
nand U5125 (N_5125,N_4594,N_4020);
and U5126 (N_5126,N_4423,N_4121);
nor U5127 (N_5127,N_4629,N_4251);
nor U5128 (N_5128,N_4174,N_4785);
or U5129 (N_5129,N_4897,N_4247);
and U5130 (N_5130,N_4718,N_4671);
nor U5131 (N_5131,N_4781,N_4147);
nand U5132 (N_5132,N_4031,N_4745);
and U5133 (N_5133,N_4672,N_4771);
or U5134 (N_5134,N_4645,N_4090);
xnor U5135 (N_5135,N_4312,N_4450);
or U5136 (N_5136,N_4487,N_4528);
and U5137 (N_5137,N_4680,N_4641);
and U5138 (N_5138,N_4698,N_4353);
xor U5139 (N_5139,N_4329,N_4592);
nor U5140 (N_5140,N_4911,N_4148);
nand U5141 (N_5141,N_4900,N_4990);
or U5142 (N_5142,N_4971,N_4013);
nand U5143 (N_5143,N_4361,N_4337);
or U5144 (N_5144,N_4107,N_4235);
nand U5145 (N_5145,N_4416,N_4690);
xor U5146 (N_5146,N_4975,N_4822);
xnor U5147 (N_5147,N_4566,N_4309);
or U5148 (N_5148,N_4120,N_4321);
nand U5149 (N_5149,N_4509,N_4524);
or U5150 (N_5150,N_4700,N_4499);
and U5151 (N_5151,N_4764,N_4162);
xnor U5152 (N_5152,N_4104,N_4019);
nand U5153 (N_5153,N_4824,N_4420);
and U5154 (N_5154,N_4551,N_4459);
nor U5155 (N_5155,N_4500,N_4851);
xnor U5156 (N_5156,N_4383,N_4056);
nand U5157 (N_5157,N_4997,N_4224);
and U5158 (N_5158,N_4244,N_4208);
xor U5159 (N_5159,N_4049,N_4896);
nand U5160 (N_5160,N_4030,N_4219);
or U5161 (N_5161,N_4962,N_4791);
nor U5162 (N_5162,N_4934,N_4024);
or U5163 (N_5163,N_4496,N_4204);
and U5164 (N_5164,N_4612,N_4440);
and U5165 (N_5165,N_4850,N_4958);
nor U5166 (N_5166,N_4059,N_4868);
xor U5167 (N_5167,N_4130,N_4273);
or U5168 (N_5168,N_4999,N_4969);
xnor U5169 (N_5169,N_4110,N_4225);
or U5170 (N_5170,N_4456,N_4311);
or U5171 (N_5171,N_4201,N_4325);
nor U5172 (N_5172,N_4753,N_4212);
and U5173 (N_5173,N_4048,N_4004);
nand U5174 (N_5174,N_4620,N_4588);
nand U5175 (N_5175,N_4310,N_4047);
and U5176 (N_5176,N_4576,N_4391);
xor U5177 (N_5177,N_4397,N_4869);
and U5178 (N_5178,N_4754,N_4447);
nor U5179 (N_5179,N_4800,N_4925);
nand U5180 (N_5180,N_4668,N_4374);
or U5181 (N_5181,N_4898,N_4408);
nand U5182 (N_5182,N_4259,N_4067);
or U5183 (N_5183,N_4916,N_4016);
and U5184 (N_5184,N_4448,N_4667);
nor U5185 (N_5185,N_4352,N_4438);
or U5186 (N_5186,N_4686,N_4405);
nand U5187 (N_5187,N_4324,N_4386);
and U5188 (N_5188,N_4708,N_4821);
and U5189 (N_5189,N_4927,N_4596);
xor U5190 (N_5190,N_4986,N_4089);
and U5191 (N_5191,N_4784,N_4779);
nor U5192 (N_5192,N_4519,N_4539);
xor U5193 (N_5193,N_4218,N_4434);
and U5194 (N_5194,N_4831,N_4621);
xor U5195 (N_5195,N_4268,N_4015);
xnor U5196 (N_5196,N_4033,N_4506);
nor U5197 (N_5197,N_4649,N_4531);
nand U5198 (N_5198,N_4075,N_4688);
and U5199 (N_5199,N_4609,N_4595);
xnor U5200 (N_5200,N_4230,N_4545);
nor U5201 (N_5201,N_4829,N_4867);
xor U5202 (N_5202,N_4537,N_4526);
nor U5203 (N_5203,N_4647,N_4633);
or U5204 (N_5204,N_4823,N_4190);
and U5205 (N_5205,N_4885,N_4313);
xnor U5206 (N_5206,N_4601,N_4623);
xnor U5207 (N_5207,N_4101,N_4260);
and U5208 (N_5208,N_4115,N_4766);
xor U5209 (N_5209,N_4857,N_4827);
xor U5210 (N_5210,N_4032,N_4145);
nor U5211 (N_5211,N_4203,N_4541);
nand U5212 (N_5212,N_4415,N_4722);
xor U5213 (N_5213,N_4180,N_4702);
xor U5214 (N_5214,N_4630,N_4451);
nand U5215 (N_5215,N_4135,N_4064);
nand U5216 (N_5216,N_4747,N_4828);
xor U5217 (N_5217,N_4052,N_4866);
or U5218 (N_5218,N_4505,N_4726);
nand U5219 (N_5219,N_4430,N_4364);
nor U5220 (N_5220,N_4085,N_4402);
nor U5221 (N_5221,N_4573,N_4730);
nor U5222 (N_5222,N_4051,N_4544);
nor U5223 (N_5223,N_4695,N_4291);
nor U5224 (N_5224,N_4172,N_4328);
xnor U5225 (N_5225,N_4304,N_4303);
or U5226 (N_5226,N_4904,N_4138);
xnor U5227 (N_5227,N_4716,N_4786);
or U5228 (N_5228,N_4678,N_4283);
nor U5229 (N_5229,N_4142,N_4124);
nand U5230 (N_5230,N_4131,N_4068);
nand U5231 (N_5231,N_4058,N_4211);
xor U5232 (N_5232,N_4939,N_4409);
nor U5233 (N_5233,N_4128,N_4723);
nor U5234 (N_5234,N_4546,N_4306);
xnor U5235 (N_5235,N_4177,N_4777);
or U5236 (N_5236,N_4946,N_4341);
and U5237 (N_5237,N_4750,N_4814);
xor U5238 (N_5238,N_4653,N_4915);
xor U5239 (N_5239,N_4733,N_4663);
nand U5240 (N_5240,N_4920,N_4959);
nor U5241 (N_5241,N_4614,N_4605);
or U5242 (N_5242,N_4562,N_4073);
xnor U5243 (N_5243,N_4575,N_4884);
nor U5244 (N_5244,N_4574,N_4604);
nor U5245 (N_5245,N_4799,N_4109);
xor U5246 (N_5246,N_4349,N_4125);
xnor U5247 (N_5247,N_4945,N_4292);
and U5248 (N_5248,N_4398,N_4590);
or U5249 (N_5249,N_4326,N_4746);
nand U5250 (N_5250,N_4242,N_4587);
or U5251 (N_5251,N_4372,N_4252);
xor U5252 (N_5252,N_4937,N_4673);
or U5253 (N_5253,N_4666,N_4511);
xor U5254 (N_5254,N_4835,N_4433);
and U5255 (N_5255,N_4660,N_4944);
xor U5256 (N_5256,N_4906,N_4642);
xnor U5257 (N_5257,N_4371,N_4631);
nand U5258 (N_5258,N_4093,N_4568);
and U5259 (N_5259,N_4082,N_4677);
nand U5260 (N_5260,N_4685,N_4988);
and U5261 (N_5261,N_4985,N_4772);
nand U5262 (N_5262,N_4520,N_4342);
nand U5263 (N_5263,N_4084,N_4992);
nor U5264 (N_5264,N_4334,N_4692);
nand U5265 (N_5265,N_4968,N_4284);
nor U5266 (N_5266,N_4652,N_4240);
xor U5267 (N_5267,N_4213,N_4817);
and U5268 (N_5268,N_4122,N_4422);
nor U5269 (N_5269,N_4229,N_4741);
nand U5270 (N_5270,N_4379,N_4427);
nor U5271 (N_5271,N_4484,N_4318);
xor U5272 (N_5272,N_4157,N_4238);
or U5273 (N_5273,N_4886,N_4512);
and U5274 (N_5274,N_4194,N_4796);
nor U5275 (N_5275,N_4974,N_4865);
nor U5276 (N_5276,N_4446,N_4600);
and U5277 (N_5277,N_4953,N_4045);
xor U5278 (N_5278,N_4206,N_4522);
and U5279 (N_5279,N_4146,N_4369);
nor U5280 (N_5280,N_4903,N_4441);
or U5281 (N_5281,N_4489,N_4810);
or U5282 (N_5282,N_4984,N_4625);
nand U5283 (N_5283,N_4930,N_4041);
nor U5284 (N_5284,N_4888,N_4287);
nand U5285 (N_5285,N_4078,N_4096);
or U5286 (N_5286,N_4062,N_4263);
or U5287 (N_5287,N_4891,N_4350);
nand U5288 (N_5288,N_4721,N_4488);
nand U5289 (N_5289,N_4586,N_4852);
nor U5290 (N_5290,N_4582,N_4597);
nor U5291 (N_5291,N_4581,N_4770);
nand U5292 (N_5292,N_4442,N_4910);
xor U5293 (N_5293,N_4762,N_4160);
or U5294 (N_5294,N_4464,N_4553);
or U5295 (N_5295,N_4359,N_4037);
or U5296 (N_5296,N_4296,N_4486);
nor U5297 (N_5297,N_4274,N_4523);
xnor U5298 (N_5298,N_4000,N_4302);
xnor U5299 (N_5299,N_4720,N_4755);
nand U5300 (N_5300,N_4989,N_4579);
xnor U5301 (N_5301,N_4602,N_4226);
or U5302 (N_5302,N_4139,N_4683);
or U5303 (N_5303,N_4387,N_4216);
or U5304 (N_5304,N_4844,N_4950);
xnor U5305 (N_5305,N_4155,N_4005);
or U5306 (N_5306,N_4957,N_4137);
xor U5307 (N_5307,N_4479,N_4322);
xnor U5308 (N_5308,N_4473,N_4258);
and U5309 (N_5309,N_4806,N_4141);
nor U5310 (N_5310,N_4923,N_4254);
and U5311 (N_5311,N_4963,N_4395);
or U5312 (N_5312,N_4729,N_4161);
and U5313 (N_5313,N_4598,N_4550);
xnor U5314 (N_5314,N_4577,N_4743);
and U5315 (N_5315,N_4567,N_4860);
or U5316 (N_5316,N_4518,N_4848);
and U5317 (N_5317,N_4023,N_4346);
nor U5318 (N_5318,N_4394,N_4393);
nor U5319 (N_5319,N_4724,N_4548);
and U5320 (N_5320,N_4237,N_4917);
or U5321 (N_5321,N_4593,N_4214);
nand U5322 (N_5322,N_4119,N_4102);
or U5323 (N_5323,N_4876,N_4658);
xor U5324 (N_5324,N_4707,N_4241);
and U5325 (N_5325,N_4267,N_4732);
or U5326 (N_5326,N_4936,N_4196);
and U5327 (N_5327,N_4648,N_4472);
xor U5328 (N_5328,N_4570,N_4286);
or U5329 (N_5329,N_4367,N_4748);
xnor U5330 (N_5330,N_4462,N_4530);
and U5331 (N_5331,N_4086,N_4388);
and U5332 (N_5332,N_4046,N_4651);
nor U5333 (N_5333,N_4264,N_4744);
nand U5334 (N_5334,N_4697,N_4820);
nand U5335 (N_5335,N_4176,N_4410);
nand U5336 (N_5336,N_4092,N_4173);
and U5337 (N_5337,N_4725,N_4681);
nor U5338 (N_5338,N_4502,N_4858);
xnor U5339 (N_5339,N_4012,N_4557);
xor U5340 (N_5340,N_4558,N_4826);
and U5341 (N_5341,N_4607,N_4403);
xnor U5342 (N_5342,N_4584,N_4076);
or U5343 (N_5343,N_4490,N_4536);
xor U5344 (N_5344,N_4554,N_4682);
and U5345 (N_5345,N_4951,N_4300);
and U5346 (N_5346,N_4508,N_4335);
or U5347 (N_5347,N_4080,N_4069);
nor U5348 (N_5348,N_4719,N_4669);
or U5349 (N_5349,N_4140,N_4485);
nand U5350 (N_5350,N_4540,N_4565);
and U5351 (N_5351,N_4344,N_4431);
or U5352 (N_5352,N_4914,N_4257);
nand U5353 (N_5353,N_4757,N_4170);
xnor U5354 (N_5354,N_4940,N_4428);
nand U5355 (N_5355,N_4332,N_4628);
nor U5356 (N_5356,N_4455,N_4735);
nor U5357 (N_5357,N_4932,N_4444);
and U5358 (N_5358,N_4507,N_4765);
nand U5359 (N_5359,N_4060,N_4552);
xor U5360 (N_5360,N_4007,N_4661);
nand U5361 (N_5361,N_4057,N_4153);
xor U5362 (N_5362,N_4691,N_4436);
xor U5363 (N_5363,N_4987,N_4042);
xnor U5364 (N_5364,N_4111,N_4221);
nand U5365 (N_5365,N_4705,N_4378);
nor U5366 (N_5366,N_4277,N_4195);
nor U5367 (N_5367,N_4738,N_4874);
xnor U5368 (N_5368,N_4055,N_4790);
nand U5369 (N_5369,N_4463,N_4504);
or U5370 (N_5370,N_4578,N_4034);
or U5371 (N_5371,N_4847,N_4615);
xnor U5372 (N_5372,N_4305,N_4465);
nand U5373 (N_5373,N_4815,N_4752);
nor U5374 (N_5374,N_4280,N_4793);
or U5375 (N_5375,N_4977,N_4949);
xnor U5376 (N_5376,N_4357,N_4803);
and U5377 (N_5377,N_4129,N_4943);
xor U5378 (N_5378,N_4543,N_4269);
and U5379 (N_5379,N_4118,N_4892);
xor U5380 (N_5380,N_4774,N_4983);
nand U5381 (N_5381,N_4704,N_4117);
or U5382 (N_5382,N_4207,N_4619);
nand U5383 (N_5383,N_4617,N_4198);
nand U5384 (N_5384,N_4236,N_4713);
xnor U5385 (N_5385,N_4859,N_4993);
and U5386 (N_5386,N_4065,N_4414);
nand U5387 (N_5387,N_4074,N_4717);
or U5388 (N_5388,N_4186,N_4470);
nand U5389 (N_5389,N_4088,N_4825);
xnor U5390 (N_5390,N_4255,N_4563);
nor U5391 (N_5391,N_4108,N_4760);
nor U5392 (N_5392,N_4529,N_4163);
nor U5393 (N_5393,N_4113,N_4025);
nor U5394 (N_5394,N_4956,N_4599);
nand U5395 (N_5395,N_4396,N_4043);
nand U5396 (N_5396,N_4382,N_4942);
nand U5397 (N_5397,N_4360,N_4271);
nand U5398 (N_5398,N_4091,N_4811);
nor U5399 (N_5399,N_4533,N_4183);
nor U5400 (N_5400,N_4187,N_4768);
or U5401 (N_5401,N_4908,N_4773);
xnor U5402 (N_5402,N_4355,N_4861);
or U5403 (N_5403,N_4837,N_4478);
nor U5404 (N_5404,N_4014,N_4452);
xor U5405 (N_5405,N_4010,N_4345);
nand U5406 (N_5406,N_4159,N_4294);
nor U5407 (N_5407,N_4756,N_4591);
and U5408 (N_5408,N_4564,N_4840);
or U5409 (N_5409,N_4223,N_4547);
nor U5410 (N_5410,N_4510,N_4404);
or U5411 (N_5411,N_4909,N_4400);
or U5412 (N_5412,N_4103,N_4285);
and U5413 (N_5413,N_4901,N_4981);
xnor U5414 (N_5414,N_4919,N_4736);
xor U5415 (N_5415,N_4843,N_4492);
or U5416 (N_5416,N_4996,N_4192);
nand U5417 (N_5417,N_4330,N_4549);
or U5418 (N_5418,N_4381,N_4676);
nor U5419 (N_5419,N_4333,N_4017);
and U5420 (N_5420,N_4480,N_4385);
nand U5421 (N_5421,N_4454,N_4714);
xnor U5422 (N_5422,N_4054,N_4960);
xor U5423 (N_5423,N_4288,N_4805);
nand U5424 (N_5424,N_4699,N_4572);
nor U5425 (N_5425,N_4863,N_4314);
and U5426 (N_5426,N_4689,N_4301);
nor U5427 (N_5427,N_4767,N_4870);
and U5428 (N_5428,N_4926,N_4392);
nand U5429 (N_5429,N_4327,N_4474);
or U5430 (N_5430,N_4154,N_4149);
or U5431 (N_5431,N_4656,N_4270);
nor U5432 (N_5432,N_4407,N_4072);
nor U5433 (N_5433,N_4181,N_4706);
or U5434 (N_5434,N_4193,N_4933);
xor U5435 (N_5435,N_4616,N_4425);
nand U5436 (N_5436,N_4127,N_4838);
xor U5437 (N_5437,N_4763,N_4818);
or U5438 (N_5438,N_4644,N_4880);
or U5439 (N_5439,N_4839,N_4872);
or U5440 (N_5440,N_4941,N_4998);
or U5441 (N_5441,N_4373,N_4662);
nor U5442 (N_5442,N_4542,N_4340);
xnor U5443 (N_5443,N_4935,N_4709);
and U5444 (N_5444,N_4532,N_4233);
nand U5445 (N_5445,N_4001,N_4610);
xor U5446 (N_5446,N_4282,N_4966);
and U5447 (N_5447,N_4964,N_4854);
nand U5448 (N_5448,N_4979,N_4972);
xnor U5449 (N_5449,N_4006,N_4924);
nor U5450 (N_5450,N_4278,N_4380);
xor U5451 (N_5451,N_4687,N_4665);
or U5452 (N_5452,N_4460,N_4684);
xor U5453 (N_5453,N_4429,N_4008);
xor U5454 (N_5454,N_4133,N_4727);
or U5455 (N_5455,N_4922,N_4809);
or U5456 (N_5456,N_4424,N_4336);
or U5457 (N_5457,N_4783,N_4833);
or U5458 (N_5458,N_4220,N_4476);
and U5459 (N_5459,N_4152,N_4497);
or U5460 (N_5460,N_4834,N_4175);
nor U5461 (N_5461,N_4319,N_4877);
or U5462 (N_5462,N_4123,N_4320);
nand U5463 (N_5463,N_4112,N_4538);
nor U5464 (N_5464,N_4494,N_4339);
xnor U5465 (N_5465,N_4376,N_4437);
nand U5466 (N_5466,N_4636,N_4151);
nand U5467 (N_5467,N_4498,N_4948);
and U5468 (N_5468,N_4040,N_4637);
nor U5469 (N_5469,N_4061,N_4608);
nand U5470 (N_5470,N_4217,N_4021);
or U5471 (N_5471,N_4039,N_4794);
or U5472 (N_5472,N_4491,N_4370);
or U5473 (N_5473,N_4368,N_4412);
xor U5474 (N_5474,N_4782,N_4994);
and U5475 (N_5475,N_4222,N_4316);
nor U5476 (N_5476,N_4515,N_4503);
and U5477 (N_5477,N_4640,N_4890);
and U5478 (N_5478,N_4559,N_4299);
or U5479 (N_5479,N_4675,N_4802);
and U5480 (N_5480,N_4002,N_4788);
xnor U5481 (N_5481,N_4938,N_4646);
and U5482 (N_5482,N_4635,N_4232);
nor U5483 (N_5483,N_4363,N_4525);
or U5484 (N_5484,N_4583,N_4477);
nor U5485 (N_5485,N_4066,N_4871);
nand U5486 (N_5486,N_4384,N_4467);
nand U5487 (N_5487,N_4009,N_4632);
xor U5488 (N_5488,N_4417,N_4132);
xor U5489 (N_5489,N_4853,N_4323);
and U5490 (N_5490,N_4878,N_4855);
and U5491 (N_5491,N_4164,N_4787);
nand U5492 (N_5492,N_4169,N_4458);
and U5493 (N_5493,N_4028,N_4375);
xor U5494 (N_5494,N_4929,N_4136);
nand U5495 (N_5495,N_4248,N_4011);
xnor U5496 (N_5496,N_4289,N_4087);
xnor U5497 (N_5497,N_4036,N_4907);
and U5498 (N_5498,N_4928,N_4231);
or U5499 (N_5499,N_4105,N_4243);
xor U5500 (N_5500,N_4292,N_4355);
xnor U5501 (N_5501,N_4943,N_4785);
nor U5502 (N_5502,N_4926,N_4713);
nor U5503 (N_5503,N_4810,N_4660);
xnor U5504 (N_5504,N_4687,N_4897);
and U5505 (N_5505,N_4861,N_4747);
and U5506 (N_5506,N_4730,N_4467);
and U5507 (N_5507,N_4702,N_4275);
nor U5508 (N_5508,N_4601,N_4944);
and U5509 (N_5509,N_4207,N_4323);
nor U5510 (N_5510,N_4002,N_4325);
nor U5511 (N_5511,N_4311,N_4832);
or U5512 (N_5512,N_4495,N_4481);
nor U5513 (N_5513,N_4891,N_4496);
nor U5514 (N_5514,N_4385,N_4498);
and U5515 (N_5515,N_4592,N_4719);
nand U5516 (N_5516,N_4470,N_4968);
or U5517 (N_5517,N_4051,N_4554);
and U5518 (N_5518,N_4535,N_4206);
or U5519 (N_5519,N_4688,N_4284);
xor U5520 (N_5520,N_4136,N_4755);
nor U5521 (N_5521,N_4260,N_4906);
nor U5522 (N_5522,N_4748,N_4654);
or U5523 (N_5523,N_4894,N_4883);
xor U5524 (N_5524,N_4978,N_4914);
xor U5525 (N_5525,N_4851,N_4866);
xnor U5526 (N_5526,N_4085,N_4032);
and U5527 (N_5527,N_4822,N_4894);
and U5528 (N_5528,N_4859,N_4652);
or U5529 (N_5529,N_4355,N_4840);
and U5530 (N_5530,N_4170,N_4813);
nand U5531 (N_5531,N_4700,N_4731);
nand U5532 (N_5532,N_4160,N_4124);
or U5533 (N_5533,N_4935,N_4192);
or U5534 (N_5534,N_4212,N_4084);
xor U5535 (N_5535,N_4026,N_4346);
nor U5536 (N_5536,N_4277,N_4608);
xnor U5537 (N_5537,N_4678,N_4219);
xor U5538 (N_5538,N_4033,N_4943);
or U5539 (N_5539,N_4128,N_4475);
xnor U5540 (N_5540,N_4162,N_4139);
nand U5541 (N_5541,N_4006,N_4325);
xnor U5542 (N_5542,N_4690,N_4005);
or U5543 (N_5543,N_4479,N_4110);
and U5544 (N_5544,N_4214,N_4824);
xor U5545 (N_5545,N_4840,N_4281);
nor U5546 (N_5546,N_4685,N_4752);
nand U5547 (N_5547,N_4468,N_4662);
and U5548 (N_5548,N_4026,N_4469);
and U5549 (N_5549,N_4077,N_4204);
nand U5550 (N_5550,N_4776,N_4003);
nand U5551 (N_5551,N_4667,N_4150);
xor U5552 (N_5552,N_4308,N_4565);
and U5553 (N_5553,N_4114,N_4142);
nor U5554 (N_5554,N_4431,N_4222);
or U5555 (N_5555,N_4519,N_4953);
xor U5556 (N_5556,N_4137,N_4490);
and U5557 (N_5557,N_4671,N_4567);
and U5558 (N_5558,N_4476,N_4391);
or U5559 (N_5559,N_4245,N_4824);
or U5560 (N_5560,N_4074,N_4340);
nor U5561 (N_5561,N_4634,N_4703);
nand U5562 (N_5562,N_4713,N_4440);
or U5563 (N_5563,N_4293,N_4145);
nand U5564 (N_5564,N_4451,N_4040);
xor U5565 (N_5565,N_4454,N_4237);
nor U5566 (N_5566,N_4504,N_4798);
nand U5567 (N_5567,N_4308,N_4485);
nand U5568 (N_5568,N_4550,N_4039);
and U5569 (N_5569,N_4544,N_4911);
or U5570 (N_5570,N_4413,N_4448);
nor U5571 (N_5571,N_4481,N_4764);
xnor U5572 (N_5572,N_4880,N_4287);
nand U5573 (N_5573,N_4181,N_4461);
and U5574 (N_5574,N_4507,N_4617);
nor U5575 (N_5575,N_4701,N_4666);
nand U5576 (N_5576,N_4370,N_4565);
xor U5577 (N_5577,N_4570,N_4632);
nor U5578 (N_5578,N_4237,N_4479);
nor U5579 (N_5579,N_4329,N_4154);
nand U5580 (N_5580,N_4812,N_4616);
nor U5581 (N_5581,N_4339,N_4006);
nand U5582 (N_5582,N_4425,N_4343);
and U5583 (N_5583,N_4030,N_4137);
nand U5584 (N_5584,N_4635,N_4984);
xnor U5585 (N_5585,N_4568,N_4210);
nand U5586 (N_5586,N_4215,N_4311);
nand U5587 (N_5587,N_4405,N_4036);
and U5588 (N_5588,N_4430,N_4513);
nor U5589 (N_5589,N_4338,N_4553);
nand U5590 (N_5590,N_4232,N_4589);
or U5591 (N_5591,N_4436,N_4319);
or U5592 (N_5592,N_4250,N_4596);
and U5593 (N_5593,N_4478,N_4555);
nor U5594 (N_5594,N_4323,N_4443);
or U5595 (N_5595,N_4539,N_4327);
xnor U5596 (N_5596,N_4021,N_4575);
nand U5597 (N_5597,N_4603,N_4599);
nor U5598 (N_5598,N_4992,N_4729);
or U5599 (N_5599,N_4217,N_4459);
or U5600 (N_5600,N_4496,N_4612);
nand U5601 (N_5601,N_4336,N_4903);
nor U5602 (N_5602,N_4939,N_4314);
nor U5603 (N_5603,N_4295,N_4142);
nand U5604 (N_5604,N_4684,N_4926);
xor U5605 (N_5605,N_4332,N_4570);
nor U5606 (N_5606,N_4423,N_4753);
nor U5607 (N_5607,N_4194,N_4415);
or U5608 (N_5608,N_4403,N_4955);
and U5609 (N_5609,N_4931,N_4886);
and U5610 (N_5610,N_4527,N_4728);
xor U5611 (N_5611,N_4880,N_4821);
nand U5612 (N_5612,N_4566,N_4501);
and U5613 (N_5613,N_4418,N_4096);
nor U5614 (N_5614,N_4132,N_4467);
nor U5615 (N_5615,N_4850,N_4024);
xor U5616 (N_5616,N_4846,N_4148);
or U5617 (N_5617,N_4903,N_4559);
xor U5618 (N_5618,N_4033,N_4124);
and U5619 (N_5619,N_4739,N_4795);
and U5620 (N_5620,N_4464,N_4974);
and U5621 (N_5621,N_4734,N_4470);
or U5622 (N_5622,N_4895,N_4847);
nor U5623 (N_5623,N_4170,N_4670);
xor U5624 (N_5624,N_4163,N_4927);
nand U5625 (N_5625,N_4326,N_4830);
nand U5626 (N_5626,N_4493,N_4880);
xor U5627 (N_5627,N_4025,N_4044);
or U5628 (N_5628,N_4390,N_4984);
xnor U5629 (N_5629,N_4848,N_4210);
nand U5630 (N_5630,N_4910,N_4613);
and U5631 (N_5631,N_4914,N_4043);
and U5632 (N_5632,N_4745,N_4386);
xor U5633 (N_5633,N_4324,N_4871);
and U5634 (N_5634,N_4411,N_4632);
nand U5635 (N_5635,N_4186,N_4738);
and U5636 (N_5636,N_4517,N_4425);
or U5637 (N_5637,N_4148,N_4748);
xnor U5638 (N_5638,N_4173,N_4664);
nor U5639 (N_5639,N_4139,N_4771);
nand U5640 (N_5640,N_4151,N_4558);
nor U5641 (N_5641,N_4802,N_4300);
and U5642 (N_5642,N_4356,N_4659);
or U5643 (N_5643,N_4505,N_4988);
nor U5644 (N_5644,N_4435,N_4122);
nor U5645 (N_5645,N_4972,N_4520);
or U5646 (N_5646,N_4560,N_4799);
xor U5647 (N_5647,N_4889,N_4808);
and U5648 (N_5648,N_4685,N_4018);
nor U5649 (N_5649,N_4731,N_4176);
nand U5650 (N_5650,N_4098,N_4716);
nor U5651 (N_5651,N_4379,N_4457);
and U5652 (N_5652,N_4112,N_4077);
nand U5653 (N_5653,N_4073,N_4371);
nand U5654 (N_5654,N_4724,N_4267);
and U5655 (N_5655,N_4147,N_4566);
and U5656 (N_5656,N_4710,N_4022);
nor U5657 (N_5657,N_4808,N_4069);
nand U5658 (N_5658,N_4172,N_4294);
nor U5659 (N_5659,N_4651,N_4570);
or U5660 (N_5660,N_4230,N_4194);
nand U5661 (N_5661,N_4961,N_4324);
or U5662 (N_5662,N_4891,N_4178);
or U5663 (N_5663,N_4051,N_4163);
xor U5664 (N_5664,N_4747,N_4043);
xnor U5665 (N_5665,N_4157,N_4664);
nand U5666 (N_5666,N_4285,N_4584);
and U5667 (N_5667,N_4991,N_4674);
xnor U5668 (N_5668,N_4155,N_4084);
or U5669 (N_5669,N_4043,N_4578);
or U5670 (N_5670,N_4837,N_4903);
and U5671 (N_5671,N_4528,N_4236);
xnor U5672 (N_5672,N_4628,N_4611);
nor U5673 (N_5673,N_4638,N_4501);
xnor U5674 (N_5674,N_4657,N_4426);
nor U5675 (N_5675,N_4162,N_4240);
and U5676 (N_5676,N_4249,N_4644);
nand U5677 (N_5677,N_4752,N_4985);
nand U5678 (N_5678,N_4743,N_4485);
or U5679 (N_5679,N_4172,N_4473);
and U5680 (N_5680,N_4001,N_4625);
nor U5681 (N_5681,N_4954,N_4139);
and U5682 (N_5682,N_4348,N_4600);
xor U5683 (N_5683,N_4341,N_4066);
nand U5684 (N_5684,N_4001,N_4476);
nand U5685 (N_5685,N_4128,N_4560);
or U5686 (N_5686,N_4040,N_4616);
or U5687 (N_5687,N_4997,N_4177);
and U5688 (N_5688,N_4628,N_4258);
xnor U5689 (N_5689,N_4277,N_4547);
or U5690 (N_5690,N_4196,N_4595);
xnor U5691 (N_5691,N_4022,N_4349);
or U5692 (N_5692,N_4538,N_4278);
nand U5693 (N_5693,N_4963,N_4983);
nand U5694 (N_5694,N_4420,N_4598);
nor U5695 (N_5695,N_4572,N_4084);
nor U5696 (N_5696,N_4530,N_4481);
nand U5697 (N_5697,N_4305,N_4853);
nand U5698 (N_5698,N_4865,N_4638);
or U5699 (N_5699,N_4024,N_4733);
nand U5700 (N_5700,N_4773,N_4511);
xor U5701 (N_5701,N_4868,N_4421);
or U5702 (N_5702,N_4646,N_4038);
or U5703 (N_5703,N_4848,N_4026);
and U5704 (N_5704,N_4165,N_4913);
xnor U5705 (N_5705,N_4279,N_4249);
nor U5706 (N_5706,N_4114,N_4914);
or U5707 (N_5707,N_4216,N_4961);
nand U5708 (N_5708,N_4678,N_4994);
nor U5709 (N_5709,N_4795,N_4922);
nand U5710 (N_5710,N_4484,N_4321);
and U5711 (N_5711,N_4031,N_4819);
or U5712 (N_5712,N_4848,N_4035);
nor U5713 (N_5713,N_4300,N_4792);
xor U5714 (N_5714,N_4553,N_4622);
or U5715 (N_5715,N_4564,N_4442);
nand U5716 (N_5716,N_4079,N_4589);
or U5717 (N_5717,N_4339,N_4814);
nor U5718 (N_5718,N_4080,N_4168);
nor U5719 (N_5719,N_4750,N_4166);
or U5720 (N_5720,N_4930,N_4202);
nand U5721 (N_5721,N_4458,N_4182);
nor U5722 (N_5722,N_4469,N_4125);
or U5723 (N_5723,N_4961,N_4600);
nor U5724 (N_5724,N_4052,N_4699);
or U5725 (N_5725,N_4957,N_4429);
nand U5726 (N_5726,N_4154,N_4115);
or U5727 (N_5727,N_4210,N_4843);
and U5728 (N_5728,N_4222,N_4368);
or U5729 (N_5729,N_4689,N_4260);
xnor U5730 (N_5730,N_4919,N_4904);
and U5731 (N_5731,N_4000,N_4676);
xor U5732 (N_5732,N_4711,N_4564);
xnor U5733 (N_5733,N_4081,N_4624);
nand U5734 (N_5734,N_4828,N_4033);
nand U5735 (N_5735,N_4175,N_4897);
xnor U5736 (N_5736,N_4955,N_4787);
or U5737 (N_5737,N_4405,N_4535);
nand U5738 (N_5738,N_4991,N_4269);
nor U5739 (N_5739,N_4689,N_4999);
or U5740 (N_5740,N_4601,N_4166);
and U5741 (N_5741,N_4371,N_4505);
and U5742 (N_5742,N_4266,N_4627);
or U5743 (N_5743,N_4853,N_4789);
xnor U5744 (N_5744,N_4572,N_4228);
or U5745 (N_5745,N_4450,N_4010);
xor U5746 (N_5746,N_4502,N_4247);
and U5747 (N_5747,N_4939,N_4253);
or U5748 (N_5748,N_4118,N_4570);
or U5749 (N_5749,N_4989,N_4876);
or U5750 (N_5750,N_4501,N_4591);
nor U5751 (N_5751,N_4072,N_4836);
xor U5752 (N_5752,N_4334,N_4010);
xor U5753 (N_5753,N_4763,N_4466);
xnor U5754 (N_5754,N_4853,N_4563);
xnor U5755 (N_5755,N_4164,N_4483);
nand U5756 (N_5756,N_4741,N_4799);
nand U5757 (N_5757,N_4327,N_4006);
nand U5758 (N_5758,N_4595,N_4499);
xnor U5759 (N_5759,N_4324,N_4547);
or U5760 (N_5760,N_4395,N_4733);
nor U5761 (N_5761,N_4284,N_4981);
xor U5762 (N_5762,N_4956,N_4264);
and U5763 (N_5763,N_4610,N_4974);
nor U5764 (N_5764,N_4111,N_4720);
xor U5765 (N_5765,N_4578,N_4020);
or U5766 (N_5766,N_4675,N_4305);
xor U5767 (N_5767,N_4164,N_4235);
and U5768 (N_5768,N_4791,N_4260);
and U5769 (N_5769,N_4262,N_4341);
and U5770 (N_5770,N_4938,N_4400);
nor U5771 (N_5771,N_4373,N_4804);
and U5772 (N_5772,N_4158,N_4701);
or U5773 (N_5773,N_4338,N_4657);
and U5774 (N_5774,N_4967,N_4837);
xnor U5775 (N_5775,N_4431,N_4910);
or U5776 (N_5776,N_4559,N_4317);
or U5777 (N_5777,N_4391,N_4990);
or U5778 (N_5778,N_4237,N_4981);
or U5779 (N_5779,N_4595,N_4369);
xnor U5780 (N_5780,N_4206,N_4294);
nor U5781 (N_5781,N_4803,N_4617);
nand U5782 (N_5782,N_4271,N_4541);
and U5783 (N_5783,N_4738,N_4483);
and U5784 (N_5784,N_4911,N_4256);
or U5785 (N_5785,N_4035,N_4160);
xor U5786 (N_5786,N_4363,N_4455);
nor U5787 (N_5787,N_4662,N_4803);
nand U5788 (N_5788,N_4324,N_4506);
or U5789 (N_5789,N_4936,N_4247);
nand U5790 (N_5790,N_4464,N_4203);
nor U5791 (N_5791,N_4574,N_4150);
xnor U5792 (N_5792,N_4425,N_4034);
and U5793 (N_5793,N_4857,N_4590);
nand U5794 (N_5794,N_4799,N_4378);
xor U5795 (N_5795,N_4459,N_4104);
nor U5796 (N_5796,N_4916,N_4377);
and U5797 (N_5797,N_4101,N_4186);
nor U5798 (N_5798,N_4815,N_4105);
nor U5799 (N_5799,N_4541,N_4647);
nor U5800 (N_5800,N_4463,N_4717);
nor U5801 (N_5801,N_4400,N_4088);
nand U5802 (N_5802,N_4343,N_4243);
or U5803 (N_5803,N_4063,N_4377);
or U5804 (N_5804,N_4188,N_4525);
nand U5805 (N_5805,N_4230,N_4466);
xor U5806 (N_5806,N_4574,N_4269);
nor U5807 (N_5807,N_4592,N_4985);
nand U5808 (N_5808,N_4427,N_4418);
nor U5809 (N_5809,N_4009,N_4169);
and U5810 (N_5810,N_4454,N_4346);
xnor U5811 (N_5811,N_4083,N_4801);
nand U5812 (N_5812,N_4072,N_4543);
or U5813 (N_5813,N_4502,N_4090);
or U5814 (N_5814,N_4493,N_4038);
xor U5815 (N_5815,N_4911,N_4484);
and U5816 (N_5816,N_4555,N_4259);
nand U5817 (N_5817,N_4079,N_4946);
nor U5818 (N_5818,N_4784,N_4704);
or U5819 (N_5819,N_4755,N_4019);
xnor U5820 (N_5820,N_4993,N_4408);
xnor U5821 (N_5821,N_4879,N_4513);
or U5822 (N_5822,N_4517,N_4688);
or U5823 (N_5823,N_4217,N_4303);
nor U5824 (N_5824,N_4241,N_4067);
or U5825 (N_5825,N_4013,N_4781);
xnor U5826 (N_5826,N_4648,N_4572);
nor U5827 (N_5827,N_4134,N_4875);
or U5828 (N_5828,N_4107,N_4459);
and U5829 (N_5829,N_4559,N_4583);
and U5830 (N_5830,N_4217,N_4171);
nand U5831 (N_5831,N_4973,N_4473);
and U5832 (N_5832,N_4667,N_4374);
xnor U5833 (N_5833,N_4030,N_4698);
nand U5834 (N_5834,N_4104,N_4428);
nand U5835 (N_5835,N_4473,N_4267);
or U5836 (N_5836,N_4517,N_4619);
and U5837 (N_5837,N_4929,N_4895);
nand U5838 (N_5838,N_4925,N_4856);
xor U5839 (N_5839,N_4627,N_4908);
nand U5840 (N_5840,N_4611,N_4699);
and U5841 (N_5841,N_4896,N_4540);
nor U5842 (N_5842,N_4945,N_4001);
or U5843 (N_5843,N_4492,N_4741);
or U5844 (N_5844,N_4399,N_4496);
nor U5845 (N_5845,N_4588,N_4360);
xor U5846 (N_5846,N_4884,N_4422);
xnor U5847 (N_5847,N_4909,N_4379);
nor U5848 (N_5848,N_4587,N_4071);
nand U5849 (N_5849,N_4540,N_4902);
or U5850 (N_5850,N_4115,N_4759);
nor U5851 (N_5851,N_4278,N_4815);
nor U5852 (N_5852,N_4577,N_4552);
xor U5853 (N_5853,N_4591,N_4657);
nor U5854 (N_5854,N_4217,N_4250);
or U5855 (N_5855,N_4090,N_4501);
nand U5856 (N_5856,N_4018,N_4878);
nand U5857 (N_5857,N_4300,N_4038);
nor U5858 (N_5858,N_4773,N_4877);
nand U5859 (N_5859,N_4201,N_4790);
and U5860 (N_5860,N_4857,N_4577);
xnor U5861 (N_5861,N_4465,N_4432);
xor U5862 (N_5862,N_4323,N_4570);
or U5863 (N_5863,N_4750,N_4775);
and U5864 (N_5864,N_4482,N_4135);
nor U5865 (N_5865,N_4077,N_4648);
xnor U5866 (N_5866,N_4622,N_4983);
xnor U5867 (N_5867,N_4631,N_4458);
and U5868 (N_5868,N_4566,N_4496);
or U5869 (N_5869,N_4960,N_4591);
xor U5870 (N_5870,N_4861,N_4225);
nand U5871 (N_5871,N_4352,N_4398);
xor U5872 (N_5872,N_4592,N_4399);
or U5873 (N_5873,N_4819,N_4301);
nand U5874 (N_5874,N_4669,N_4845);
nand U5875 (N_5875,N_4943,N_4401);
nand U5876 (N_5876,N_4047,N_4835);
nand U5877 (N_5877,N_4374,N_4448);
nor U5878 (N_5878,N_4260,N_4710);
nand U5879 (N_5879,N_4603,N_4577);
xor U5880 (N_5880,N_4726,N_4382);
nand U5881 (N_5881,N_4773,N_4745);
nand U5882 (N_5882,N_4254,N_4450);
nor U5883 (N_5883,N_4869,N_4916);
or U5884 (N_5884,N_4391,N_4181);
nor U5885 (N_5885,N_4695,N_4000);
nand U5886 (N_5886,N_4006,N_4502);
nor U5887 (N_5887,N_4684,N_4856);
or U5888 (N_5888,N_4034,N_4885);
or U5889 (N_5889,N_4569,N_4233);
or U5890 (N_5890,N_4608,N_4717);
and U5891 (N_5891,N_4782,N_4012);
nand U5892 (N_5892,N_4151,N_4086);
xor U5893 (N_5893,N_4833,N_4869);
and U5894 (N_5894,N_4485,N_4375);
xor U5895 (N_5895,N_4630,N_4288);
and U5896 (N_5896,N_4594,N_4739);
nand U5897 (N_5897,N_4674,N_4620);
and U5898 (N_5898,N_4817,N_4623);
nor U5899 (N_5899,N_4824,N_4305);
xnor U5900 (N_5900,N_4365,N_4426);
or U5901 (N_5901,N_4956,N_4201);
or U5902 (N_5902,N_4970,N_4877);
or U5903 (N_5903,N_4442,N_4689);
nor U5904 (N_5904,N_4712,N_4719);
xor U5905 (N_5905,N_4746,N_4406);
and U5906 (N_5906,N_4402,N_4417);
nor U5907 (N_5907,N_4333,N_4391);
and U5908 (N_5908,N_4595,N_4146);
or U5909 (N_5909,N_4409,N_4255);
xnor U5910 (N_5910,N_4522,N_4021);
and U5911 (N_5911,N_4036,N_4876);
nand U5912 (N_5912,N_4282,N_4829);
or U5913 (N_5913,N_4312,N_4246);
nor U5914 (N_5914,N_4891,N_4960);
nand U5915 (N_5915,N_4434,N_4360);
and U5916 (N_5916,N_4157,N_4471);
nand U5917 (N_5917,N_4912,N_4944);
xnor U5918 (N_5918,N_4100,N_4056);
and U5919 (N_5919,N_4872,N_4789);
or U5920 (N_5920,N_4966,N_4369);
nor U5921 (N_5921,N_4957,N_4174);
and U5922 (N_5922,N_4235,N_4033);
nor U5923 (N_5923,N_4383,N_4475);
or U5924 (N_5924,N_4135,N_4313);
and U5925 (N_5925,N_4796,N_4906);
xor U5926 (N_5926,N_4510,N_4321);
nor U5927 (N_5927,N_4063,N_4203);
nand U5928 (N_5928,N_4645,N_4503);
or U5929 (N_5929,N_4796,N_4095);
nor U5930 (N_5930,N_4229,N_4459);
nor U5931 (N_5931,N_4707,N_4011);
xor U5932 (N_5932,N_4435,N_4853);
and U5933 (N_5933,N_4120,N_4358);
or U5934 (N_5934,N_4974,N_4301);
nand U5935 (N_5935,N_4168,N_4113);
and U5936 (N_5936,N_4577,N_4484);
and U5937 (N_5937,N_4508,N_4660);
or U5938 (N_5938,N_4021,N_4483);
and U5939 (N_5939,N_4368,N_4626);
nor U5940 (N_5940,N_4089,N_4411);
nand U5941 (N_5941,N_4983,N_4163);
nor U5942 (N_5942,N_4304,N_4681);
xnor U5943 (N_5943,N_4981,N_4170);
nor U5944 (N_5944,N_4076,N_4821);
xor U5945 (N_5945,N_4325,N_4413);
and U5946 (N_5946,N_4771,N_4681);
nor U5947 (N_5947,N_4684,N_4141);
nor U5948 (N_5948,N_4171,N_4758);
nand U5949 (N_5949,N_4725,N_4231);
or U5950 (N_5950,N_4944,N_4832);
or U5951 (N_5951,N_4210,N_4891);
nand U5952 (N_5952,N_4940,N_4340);
nor U5953 (N_5953,N_4623,N_4124);
and U5954 (N_5954,N_4531,N_4614);
nand U5955 (N_5955,N_4903,N_4750);
or U5956 (N_5956,N_4273,N_4578);
or U5957 (N_5957,N_4191,N_4469);
nor U5958 (N_5958,N_4359,N_4994);
nand U5959 (N_5959,N_4717,N_4352);
nor U5960 (N_5960,N_4325,N_4712);
or U5961 (N_5961,N_4798,N_4745);
xor U5962 (N_5962,N_4861,N_4072);
or U5963 (N_5963,N_4112,N_4771);
or U5964 (N_5964,N_4413,N_4499);
xor U5965 (N_5965,N_4565,N_4179);
nor U5966 (N_5966,N_4299,N_4887);
and U5967 (N_5967,N_4690,N_4138);
and U5968 (N_5968,N_4919,N_4289);
nor U5969 (N_5969,N_4071,N_4229);
xor U5970 (N_5970,N_4664,N_4218);
xor U5971 (N_5971,N_4994,N_4060);
and U5972 (N_5972,N_4396,N_4130);
nand U5973 (N_5973,N_4166,N_4671);
and U5974 (N_5974,N_4609,N_4973);
or U5975 (N_5975,N_4029,N_4916);
or U5976 (N_5976,N_4363,N_4244);
nor U5977 (N_5977,N_4952,N_4429);
or U5978 (N_5978,N_4263,N_4341);
and U5979 (N_5979,N_4342,N_4288);
and U5980 (N_5980,N_4531,N_4527);
nand U5981 (N_5981,N_4502,N_4117);
or U5982 (N_5982,N_4382,N_4342);
nand U5983 (N_5983,N_4324,N_4747);
and U5984 (N_5984,N_4432,N_4754);
nand U5985 (N_5985,N_4210,N_4541);
xor U5986 (N_5986,N_4639,N_4015);
nand U5987 (N_5987,N_4288,N_4854);
nand U5988 (N_5988,N_4248,N_4753);
xor U5989 (N_5989,N_4745,N_4298);
xnor U5990 (N_5990,N_4325,N_4831);
or U5991 (N_5991,N_4078,N_4744);
xor U5992 (N_5992,N_4103,N_4958);
nor U5993 (N_5993,N_4702,N_4555);
nor U5994 (N_5994,N_4703,N_4890);
nand U5995 (N_5995,N_4164,N_4983);
and U5996 (N_5996,N_4093,N_4580);
nor U5997 (N_5997,N_4551,N_4115);
nor U5998 (N_5998,N_4582,N_4158);
nor U5999 (N_5999,N_4390,N_4498);
and U6000 (N_6000,N_5061,N_5845);
or U6001 (N_6001,N_5710,N_5414);
and U6002 (N_6002,N_5092,N_5546);
xor U6003 (N_6003,N_5064,N_5896);
or U6004 (N_6004,N_5374,N_5880);
nor U6005 (N_6005,N_5897,N_5813);
nand U6006 (N_6006,N_5233,N_5569);
or U6007 (N_6007,N_5679,N_5276);
nor U6008 (N_6008,N_5244,N_5672);
or U6009 (N_6009,N_5922,N_5465);
xor U6010 (N_6010,N_5657,N_5749);
and U6011 (N_6011,N_5885,N_5401);
or U6012 (N_6012,N_5622,N_5871);
or U6013 (N_6013,N_5119,N_5997);
and U6014 (N_6014,N_5778,N_5819);
or U6015 (N_6015,N_5416,N_5933);
nand U6016 (N_6016,N_5069,N_5865);
nand U6017 (N_6017,N_5089,N_5982);
nor U6018 (N_6018,N_5136,N_5166);
nor U6019 (N_6019,N_5388,N_5976);
or U6020 (N_6020,N_5516,N_5338);
or U6021 (N_6021,N_5826,N_5331);
or U6022 (N_6022,N_5683,N_5219);
xnor U6023 (N_6023,N_5355,N_5760);
and U6024 (N_6024,N_5725,N_5038);
or U6025 (N_6025,N_5654,N_5066);
or U6026 (N_6026,N_5999,N_5216);
xor U6027 (N_6027,N_5767,N_5030);
xor U6028 (N_6028,N_5434,N_5192);
or U6029 (N_6029,N_5727,N_5948);
nand U6030 (N_6030,N_5052,N_5911);
nand U6031 (N_6031,N_5169,N_5944);
and U6032 (N_6032,N_5353,N_5573);
or U6033 (N_6033,N_5724,N_5133);
and U6034 (N_6034,N_5577,N_5062);
and U6035 (N_6035,N_5613,N_5540);
nand U6036 (N_6036,N_5628,N_5261);
nor U6037 (N_6037,N_5691,N_5821);
or U6038 (N_6038,N_5506,N_5502);
and U6039 (N_6039,N_5698,N_5301);
and U6040 (N_6040,N_5489,N_5806);
nor U6041 (N_6041,N_5962,N_5914);
and U6042 (N_6042,N_5956,N_5775);
and U6043 (N_6043,N_5704,N_5637);
nor U6044 (N_6044,N_5118,N_5097);
xor U6045 (N_6045,N_5236,N_5448);
and U6046 (N_6046,N_5111,N_5605);
xor U6047 (N_6047,N_5482,N_5086);
and U6048 (N_6048,N_5838,N_5527);
or U6049 (N_6049,N_5277,N_5023);
xor U6050 (N_6050,N_5805,N_5928);
and U6051 (N_6051,N_5262,N_5931);
and U6052 (N_6052,N_5854,N_5837);
nor U6053 (N_6053,N_5708,N_5474);
and U6054 (N_6054,N_5311,N_5541);
xnor U6055 (N_6055,N_5321,N_5029);
xor U6056 (N_6056,N_5522,N_5239);
and U6057 (N_6057,N_5141,N_5494);
and U6058 (N_6058,N_5270,N_5598);
nand U6059 (N_6059,N_5512,N_5830);
and U6060 (N_6060,N_5732,N_5375);
nor U6061 (N_6061,N_5712,N_5651);
and U6062 (N_6062,N_5803,N_5579);
or U6063 (N_6063,N_5720,N_5951);
nand U6064 (N_6064,N_5452,N_5281);
xor U6065 (N_6065,N_5750,N_5115);
xor U6066 (N_6066,N_5013,N_5766);
nand U6067 (N_6067,N_5295,N_5793);
nor U6068 (N_6068,N_5246,N_5399);
nor U6069 (N_6069,N_5150,N_5503);
xor U6070 (N_6070,N_5581,N_5528);
nor U6071 (N_6071,N_5293,N_5299);
and U6072 (N_6072,N_5987,N_5396);
nand U6073 (N_6073,N_5004,N_5844);
and U6074 (N_6074,N_5393,N_5570);
and U6075 (N_6075,N_5218,N_5114);
or U6076 (N_6076,N_5970,N_5888);
or U6077 (N_6077,N_5080,N_5811);
xnor U6078 (N_6078,N_5113,N_5500);
nand U6079 (N_6079,N_5436,N_5268);
nor U6080 (N_6080,N_5034,N_5363);
nor U6081 (N_6081,N_5032,N_5106);
and U6082 (N_6082,N_5751,N_5128);
xnor U6083 (N_6083,N_5902,N_5279);
xnor U6084 (N_6084,N_5453,N_5792);
or U6085 (N_6085,N_5078,N_5209);
and U6086 (N_6086,N_5650,N_5343);
nor U6087 (N_6087,N_5054,N_5587);
nor U6088 (N_6088,N_5341,N_5170);
xor U6089 (N_6089,N_5709,N_5455);
nor U6090 (N_6090,N_5350,N_5125);
nor U6091 (N_6091,N_5196,N_5059);
xor U6092 (N_6092,N_5109,N_5186);
nand U6093 (N_6093,N_5467,N_5210);
nand U6094 (N_6094,N_5789,N_5237);
or U6095 (N_6095,N_5492,N_5222);
xor U6096 (N_6096,N_5110,N_5937);
nor U6097 (N_6097,N_5894,N_5861);
nand U6098 (N_6098,N_5665,N_5898);
and U6099 (N_6099,N_5135,N_5326);
xnor U6100 (N_6100,N_5238,N_5093);
xor U6101 (N_6101,N_5242,N_5060);
nand U6102 (N_6102,N_5212,N_5006);
and U6103 (N_6103,N_5535,N_5134);
or U6104 (N_6104,N_5200,N_5260);
nor U6105 (N_6105,N_5403,N_5905);
nand U6106 (N_6106,N_5839,N_5618);
nand U6107 (N_6107,N_5938,N_5204);
xor U6108 (N_6108,N_5638,N_5490);
nor U6109 (N_6109,N_5705,N_5368);
or U6110 (N_6110,N_5499,N_5958);
or U6111 (N_6111,N_5662,N_5907);
nand U6112 (N_6112,N_5784,N_5519);
or U6113 (N_6113,N_5788,N_5493);
nor U6114 (N_6114,N_5508,N_5526);
xnor U6115 (N_6115,N_5807,N_5913);
nor U6116 (N_6116,N_5926,N_5660);
xnor U6117 (N_6117,N_5158,N_5159);
or U6118 (N_6118,N_5247,N_5692);
nand U6119 (N_6119,N_5824,N_5787);
nor U6120 (N_6120,N_5206,N_5816);
nor U6121 (N_6121,N_5825,N_5791);
nand U6122 (N_6122,N_5347,N_5728);
or U6123 (N_6123,N_5700,N_5648);
or U6124 (N_6124,N_5875,N_5731);
nor U6125 (N_6125,N_5947,N_5998);
nand U6126 (N_6126,N_5142,N_5286);
or U6127 (N_6127,N_5904,N_5263);
xor U6128 (N_6128,N_5588,N_5328);
and U6129 (N_6129,N_5258,N_5822);
nand U6130 (N_6130,N_5475,N_5954);
nand U6131 (N_6131,N_5583,N_5757);
nor U6132 (N_6132,N_5847,N_5829);
xor U6133 (N_6133,N_5730,N_5674);
nor U6134 (N_6134,N_5877,N_5383);
and U6135 (N_6135,N_5977,N_5139);
nand U6136 (N_6136,N_5544,N_5804);
or U6137 (N_6137,N_5525,N_5213);
nor U6138 (N_6138,N_5386,N_5991);
and U6139 (N_6139,N_5123,N_5696);
or U6140 (N_6140,N_5217,N_5425);
nand U6141 (N_6141,N_5621,N_5870);
or U6142 (N_6142,N_5391,N_5164);
nand U6143 (N_6143,N_5056,N_5344);
nor U6144 (N_6144,N_5678,N_5339);
nand U6145 (N_6145,N_5671,N_5563);
or U6146 (N_6146,N_5382,N_5513);
or U6147 (N_6147,N_5862,N_5876);
xor U6148 (N_6148,N_5413,N_5384);
nor U6149 (N_6149,N_5424,N_5010);
or U6150 (N_6150,N_5138,N_5079);
nor U6151 (N_6151,N_5070,N_5183);
xnor U6152 (N_6152,N_5047,N_5445);
or U6153 (N_6153,N_5539,N_5867);
xor U6154 (N_6154,N_5140,N_5906);
xnor U6155 (N_6155,N_5002,N_5108);
nor U6156 (N_6156,N_5510,N_5753);
nand U6157 (N_6157,N_5738,N_5542);
nor U6158 (N_6158,N_5664,N_5304);
nor U6159 (N_6159,N_5144,N_5318);
or U6160 (N_6160,N_5883,N_5446);
and U6161 (N_6161,N_5485,N_5895);
or U6162 (N_6162,N_5466,N_5557);
or U6163 (N_6163,N_5882,N_5016);
or U6164 (N_6164,N_5227,N_5248);
nand U6165 (N_6165,N_5939,N_5087);
and U6166 (N_6166,N_5487,N_5547);
nor U6167 (N_6167,N_5182,N_5963);
and U6168 (N_6168,N_5294,N_5495);
xnor U6169 (N_6169,N_5076,N_5614);
or U6170 (N_6170,N_5392,N_5776);
or U6171 (N_6171,N_5945,N_5795);
or U6172 (N_6172,N_5156,N_5491);
xor U6173 (N_6173,N_5249,N_5846);
xor U6174 (N_6174,N_5723,N_5044);
and U6175 (N_6175,N_5315,N_5441);
and U6176 (N_6176,N_5381,N_5744);
nand U6177 (N_6177,N_5633,N_5940);
and U6178 (N_6178,N_5361,N_5120);
nor U6179 (N_6179,N_5713,N_5981);
nand U6180 (N_6180,N_5578,N_5759);
xnor U6181 (N_6181,N_5630,N_5084);
nand U6182 (N_6182,N_5360,N_5266);
xor U6183 (N_6183,N_5632,N_5562);
and U6184 (N_6184,N_5524,N_5185);
xor U6185 (N_6185,N_5559,N_5983);
and U6186 (N_6186,N_5680,N_5287);
xor U6187 (N_6187,N_5655,N_5719);
and U6188 (N_6188,N_5305,N_5194);
and U6189 (N_6189,N_5603,N_5693);
nand U6190 (N_6190,N_5716,N_5501);
and U6191 (N_6191,N_5160,N_5722);
and U6192 (N_6192,N_5003,N_5121);
and U6193 (N_6193,N_5561,N_5874);
and U6194 (N_6194,N_5129,N_5779);
nor U6195 (N_6195,N_5031,N_5370);
nand U6196 (N_6196,N_5726,N_5349);
xor U6197 (N_6197,N_5319,N_5993);
and U6198 (N_6198,N_5278,N_5197);
nor U6199 (N_6199,N_5697,N_5601);
or U6200 (N_6200,N_5042,N_5531);
and U6201 (N_6201,N_5151,N_5313);
nor U6202 (N_6202,N_5252,N_5476);
nor U6203 (N_6203,N_5624,N_5864);
xnor U6204 (N_6204,N_5105,N_5285);
nand U6205 (N_6205,N_5908,N_5053);
nor U6206 (N_6206,N_5715,N_5148);
and U6207 (N_6207,N_5828,N_5201);
and U6208 (N_6208,N_5916,N_5320);
or U6209 (N_6209,N_5163,N_5469);
nand U6210 (N_6210,N_5832,N_5505);
or U6211 (N_6211,N_5175,N_5254);
and U6212 (N_6212,N_5690,N_5127);
or U6213 (N_6213,N_5827,N_5428);
or U6214 (N_6214,N_5560,N_5666);
nor U6215 (N_6215,N_5373,N_5610);
nand U6216 (N_6216,N_5096,N_5955);
or U6217 (N_6217,N_5377,N_5193);
nand U6218 (N_6218,N_5507,N_5656);
nor U6219 (N_6219,N_5961,N_5835);
xor U6220 (N_6220,N_5564,N_5879);
or U6221 (N_6221,N_5202,N_5191);
xor U6222 (N_6222,N_5740,N_5636);
and U6223 (N_6223,N_5521,N_5498);
nand U6224 (N_6224,N_5585,N_5763);
and U6225 (N_6225,N_5429,N_5094);
and U6226 (N_6226,N_5761,N_5145);
nand U6227 (N_6227,N_5426,N_5941);
xnor U6228 (N_6228,N_5451,N_5647);
and U6229 (N_6229,N_5990,N_5812);
and U6230 (N_6230,N_5929,N_5903);
xor U6231 (N_6231,N_5780,N_5037);
xnor U6232 (N_6232,N_5171,N_5739);
nor U6233 (N_6233,N_5020,N_5411);
nor U6234 (N_6234,N_5790,N_5126);
nand U6235 (N_6235,N_5971,N_5214);
xnor U6236 (N_6236,N_5243,N_5817);
xnor U6237 (N_6237,N_5925,N_5178);
nand U6238 (N_6238,N_5387,N_5484);
xor U6239 (N_6239,N_5440,N_5303);
or U6240 (N_6240,N_5071,N_5019);
xnor U6241 (N_6241,N_5868,N_5851);
nor U6242 (N_6242,N_5366,N_5364);
or U6243 (N_6243,N_5554,N_5405);
nand U6244 (N_6244,N_5801,N_5550);
xor U6245 (N_6245,N_5863,N_5986);
nand U6246 (N_6246,N_5917,N_5641);
nor U6247 (N_6247,N_5878,N_5001);
nor U6248 (N_6248,N_5155,N_5566);
nand U6249 (N_6249,N_5427,N_5599);
and U6250 (N_6250,N_5886,N_5417);
and U6251 (N_6251,N_5257,N_5230);
or U6252 (N_6252,N_5966,N_5421);
and U6253 (N_6253,N_5274,N_5537);
nor U6254 (N_6254,N_5153,N_5702);
nor U6255 (N_6255,N_5221,N_5556);
xnor U6256 (N_6256,N_5686,N_5533);
or U6257 (N_6257,N_5369,N_5797);
xor U6258 (N_6258,N_5745,N_5290);
xor U6259 (N_6259,N_5187,N_5721);
and U6260 (N_6260,N_5900,N_5483);
nor U6261 (N_6261,N_5346,N_5478);
xnor U6262 (N_6262,N_5777,N_5132);
and U6263 (N_6263,N_5923,N_5600);
nor U6264 (N_6264,N_5644,N_5091);
and U6265 (N_6265,N_5122,N_5706);
nor U6266 (N_6266,N_5112,N_5284);
nand U6267 (N_6267,N_5420,N_5481);
and U6268 (N_6268,N_5629,N_5607);
xnor U6269 (N_6269,N_5359,N_5602);
xor U6270 (N_6270,N_5552,N_5984);
xor U6271 (N_6271,N_5978,N_5300);
xor U6272 (N_6272,N_5275,N_5703);
nor U6273 (N_6273,N_5593,N_5943);
xor U6274 (N_6274,N_5439,N_5298);
nand U6275 (N_6275,N_5088,N_5580);
xnor U6276 (N_6276,N_5551,N_5215);
or U6277 (N_6277,N_5283,N_5893);
nor U6278 (N_6278,N_5609,N_5927);
xor U6279 (N_6279,N_5265,N_5695);
nand U6280 (N_6280,N_5770,N_5575);
nor U6281 (N_6281,N_5571,N_5459);
and U6282 (N_6282,N_5470,N_5412);
nand U6283 (N_6283,N_5124,N_5652);
xnor U6284 (N_6284,N_5949,N_5174);
nand U6285 (N_6285,N_5815,N_5773);
and U6286 (N_6286,N_5404,N_5909);
nor U6287 (N_6287,N_5497,N_5594);
xnor U6288 (N_6288,N_5729,N_5082);
xor U6289 (N_6289,N_5619,N_5232);
and U6290 (N_6290,N_5184,N_5591);
and U6291 (N_6291,N_5199,N_5988);
or U6292 (N_6292,N_5235,N_5040);
nand U6293 (N_6293,N_5608,N_5334);
and U6294 (N_6294,N_5625,N_5309);
or U6295 (N_6295,N_5406,N_5771);
and U6296 (N_6296,N_5553,N_5548);
and U6297 (N_6297,N_5946,N_5921);
nor U6298 (N_6298,N_5932,N_5324);
or U6299 (N_6299,N_5910,N_5226);
or U6300 (N_6300,N_5468,N_5543);
and U6301 (N_6301,N_5969,N_5772);
or U6302 (N_6302,N_5408,N_5675);
and U6303 (N_6303,N_5365,N_5189);
nand U6304 (N_6304,N_5754,N_5635);
nand U6305 (N_6305,N_5464,N_5565);
nor U6306 (N_6306,N_5039,N_5985);
and U6307 (N_6307,N_5081,N_5677);
and U6308 (N_6308,N_5714,N_5130);
nand U6309 (N_6309,N_5960,N_5018);
xor U6310 (N_6310,N_5220,N_5131);
nand U6311 (N_6311,N_5959,N_5586);
nor U6312 (N_6312,N_5536,N_5058);
or U6313 (N_6313,N_5859,N_5848);
and U6314 (N_6314,N_5073,N_5462);
nor U6315 (N_6315,N_5994,N_5045);
nand U6316 (N_6316,N_5668,N_5041);
or U6317 (N_6317,N_5833,N_5154);
and U6318 (N_6318,N_5930,N_5335);
or U6319 (N_6319,N_5229,N_5746);
xor U6320 (N_6320,N_5649,N_5179);
and U6321 (N_6321,N_5435,N_5884);
nand U6322 (N_6322,N_5461,N_5241);
or U6323 (N_6323,N_5090,N_5592);
nor U6324 (N_6324,N_5534,N_5228);
nor U6325 (N_6325,N_5224,N_5597);
or U6326 (N_6326,N_5617,N_5008);
nor U6327 (N_6327,N_5322,N_5858);
nor U6328 (N_6328,N_5463,N_5853);
nand U6329 (N_6329,N_5251,N_5699);
and U6330 (N_6330,N_5176,N_5850);
xnor U6331 (N_6331,N_5965,N_5919);
nand U6332 (N_6332,N_5992,N_5670);
nand U6333 (N_6333,N_5025,N_5011);
nand U6334 (N_6334,N_5180,N_5327);
xnor U6335 (N_6335,N_5967,N_5188);
or U6336 (N_6336,N_5682,N_5634);
or U6337 (N_6337,N_5509,N_5758);
nand U6338 (N_6338,N_5074,N_5515);
and U6339 (N_6339,N_5529,N_5269);
xnor U6340 (N_6340,N_5028,N_5834);
xnor U6341 (N_6341,N_5046,N_5471);
or U6342 (N_6342,N_5245,N_5177);
nor U6343 (N_6343,N_5872,N_5794);
or U6344 (N_6344,N_5457,N_5576);
or U6345 (N_6345,N_5584,N_5015);
and U6346 (N_6346,N_5240,N_5989);
and U6347 (N_6347,N_5545,N_5167);
or U6348 (N_6348,N_5810,N_5325);
or U6349 (N_6349,N_5409,N_5336);
nand U6350 (N_6350,N_5667,N_5855);
and U6351 (N_6351,N_5371,N_5051);
xnor U6352 (N_6352,N_5024,N_5259);
nand U6353 (N_6353,N_5659,N_5149);
or U6354 (N_6354,N_5454,N_5116);
nor U6355 (N_6355,N_5748,N_5117);
xor U6356 (N_6356,N_5014,N_5768);
and U6357 (N_6357,N_5255,N_5107);
xnor U6358 (N_6358,N_5430,N_5645);
nand U6359 (N_6359,N_5101,N_5021);
or U6360 (N_6360,N_5918,N_5297);
nand U6361 (N_6361,N_5643,N_5972);
xor U6362 (N_6362,N_5733,N_5161);
xnor U6363 (N_6363,N_5511,N_5400);
or U6364 (N_6364,N_5272,N_5390);
nand U6365 (N_6365,N_5687,N_5694);
nor U6366 (N_6366,N_5857,N_5234);
nor U6367 (N_6367,N_5103,N_5362);
nand U6368 (N_6368,N_5843,N_5418);
nand U6369 (N_6369,N_5302,N_5422);
and U6370 (N_6370,N_5504,N_5572);
or U6371 (N_6371,N_5574,N_5323);
xnor U6372 (N_6372,N_5207,N_5808);
nor U6373 (N_6373,N_5743,N_5673);
and U6374 (N_6374,N_5157,N_5869);
nand U6375 (N_6375,N_5205,N_5068);
nand U6376 (N_6376,N_5357,N_5866);
and U6377 (N_6377,N_5172,N_5920);
and U6378 (N_6378,N_5292,N_5181);
or U6379 (N_6379,N_5842,N_5415);
nor U6380 (N_6380,N_5211,N_5231);
or U6381 (N_6381,N_5314,N_5549);
xor U6382 (N_6382,N_5168,N_5316);
nor U6383 (N_6383,N_5518,N_5083);
and U6384 (N_6384,N_5889,N_5437);
nand U6385 (N_6385,N_5684,N_5640);
xor U6386 (N_6386,N_5642,N_5000);
and U6387 (N_6387,N_5968,N_5849);
or U6388 (N_6388,N_5852,N_5996);
nand U6389 (N_6389,N_5376,N_5555);
and U6390 (N_6390,N_5653,N_5407);
xnor U6391 (N_6391,N_5799,N_5098);
nand U6392 (N_6392,N_5582,N_5433);
and U6393 (N_6393,N_5736,N_5841);
xor U6394 (N_6394,N_5823,N_5067);
xnor U6395 (N_6395,N_5280,N_5747);
nand U6396 (N_6396,N_5718,N_5306);
or U6397 (N_6397,N_5104,N_5049);
xnor U6398 (N_6398,N_5639,N_5057);
or U6399 (N_6399,N_5798,N_5785);
nor U6400 (N_6400,N_5378,N_5095);
nand U6401 (N_6401,N_5447,N_5394);
nor U6402 (N_6402,N_5443,N_5035);
xnor U6403 (N_6403,N_5836,N_5075);
xnor U6404 (N_6404,N_5173,N_5380);
or U6405 (N_6405,N_5831,N_5742);
or U6406 (N_6406,N_5820,N_5590);
xnor U6407 (N_6407,N_5558,N_5208);
or U6408 (N_6408,N_5707,N_5762);
nand U6409 (N_6409,N_5017,N_5048);
and U6410 (N_6410,N_5022,N_5312);
xnor U6411 (N_6411,N_5432,N_5310);
or U6412 (N_6412,N_5606,N_5329);
xor U6413 (N_6413,N_5538,N_5567);
and U6414 (N_6414,N_5317,N_5271);
and U6415 (N_6415,N_5419,N_5514);
or U6416 (N_6416,N_5782,N_5410);
nor U6417 (N_6417,N_5291,N_5289);
and U6418 (N_6418,N_5616,N_5063);
nand U6419 (N_6419,N_5005,N_5774);
nand U6420 (N_6420,N_5450,N_5137);
xor U6421 (N_6421,N_5395,N_5764);
and U6422 (N_6422,N_5952,N_5354);
nor U6423 (N_6423,N_5027,N_5072);
xnor U6424 (N_6424,N_5741,N_5974);
nand U6425 (N_6425,N_5102,N_5225);
nor U6426 (N_6426,N_5669,N_5438);
nor U6427 (N_6427,N_5737,N_5620);
xnor U6428 (N_6428,N_5887,N_5356);
and U6429 (N_6429,N_5701,N_5711);
nor U6430 (N_6430,N_5973,N_5934);
and U6431 (N_6431,N_5957,N_5717);
nor U6432 (N_6432,N_5007,N_5288);
or U6433 (N_6433,N_5488,N_5950);
nand U6434 (N_6434,N_5604,N_5460);
and U6435 (N_6435,N_5912,N_5351);
nor U6436 (N_6436,N_5342,N_5818);
xor U6437 (N_6437,N_5755,N_5924);
nor U6438 (N_6438,N_5661,N_5915);
and U6439 (N_6439,N_5203,N_5267);
xor U6440 (N_6440,N_5477,N_5486);
nand U6441 (N_6441,N_5352,N_5345);
xnor U6442 (N_6442,N_5379,N_5840);
xor U6443 (N_6443,N_5523,N_5626);
and U6444 (N_6444,N_5979,N_5253);
xnor U6445 (N_6445,N_5873,N_5337);
nand U6446 (N_6446,N_5308,N_5223);
and U6447 (N_6447,N_5881,N_5036);
and U6448 (N_6448,N_5611,N_5198);
and U6449 (N_6449,N_5596,N_5612);
nand U6450 (N_6450,N_5899,N_5689);
nand U6451 (N_6451,N_5307,N_5340);
or U6452 (N_6452,N_5273,N_5765);
xor U6453 (N_6453,N_5397,N_5190);
and U6454 (N_6454,N_5055,N_5472);
nor U6455 (N_6455,N_5479,N_5783);
xor U6456 (N_6456,N_5444,N_5814);
xor U6457 (N_6457,N_5860,N_5646);
nor U6458 (N_6458,N_5423,N_5398);
nand U6459 (N_6459,N_5623,N_5735);
nand U6460 (N_6460,N_5631,N_5077);
or U6461 (N_6461,N_5615,N_5935);
xnor U6462 (N_6462,N_5250,N_5473);
and U6463 (N_6463,N_5752,N_5012);
xor U6464 (N_6464,N_5595,N_5264);
or U6465 (N_6465,N_5162,N_5332);
nand U6466 (N_6466,N_5147,N_5449);
nor U6467 (N_6467,N_5099,N_5256);
or U6468 (N_6468,N_5781,N_5146);
or U6469 (N_6469,N_5496,N_5568);
and U6470 (N_6470,N_5372,N_5033);
xnor U6471 (N_6471,N_5796,N_5936);
xnor U6472 (N_6472,N_5681,N_5165);
nor U6473 (N_6473,N_5026,N_5348);
xnor U6474 (N_6474,N_5195,N_5456);
nand U6475 (N_6475,N_5892,N_5953);
or U6476 (N_6476,N_5532,N_5458);
nor U6477 (N_6477,N_5685,N_5330);
and U6478 (N_6478,N_5769,N_5627);
nand U6479 (N_6479,N_5589,N_5100);
and U6480 (N_6480,N_5282,N_5480);
nor U6481 (N_6481,N_5043,N_5995);
and U6482 (N_6482,N_5802,N_5389);
and U6483 (N_6483,N_5658,N_5809);
xor U6484 (N_6484,N_5358,N_5856);
nand U6485 (N_6485,N_5891,N_5942);
xor U6486 (N_6486,N_5009,N_5663);
xnor U6487 (N_6487,N_5385,N_5431);
xor U6488 (N_6488,N_5517,N_5800);
nor U6489 (N_6489,N_5676,N_5890);
or U6490 (N_6490,N_5688,N_5050);
nor U6491 (N_6491,N_5143,N_5296);
nand U6492 (N_6492,N_5980,N_5975);
and U6493 (N_6493,N_5734,N_5964);
or U6494 (N_6494,N_5402,N_5085);
nor U6495 (N_6495,N_5333,N_5520);
nor U6496 (N_6496,N_5756,N_5152);
nand U6497 (N_6497,N_5442,N_5065);
nand U6498 (N_6498,N_5367,N_5901);
nor U6499 (N_6499,N_5530,N_5786);
and U6500 (N_6500,N_5108,N_5104);
or U6501 (N_6501,N_5721,N_5460);
nor U6502 (N_6502,N_5448,N_5693);
nor U6503 (N_6503,N_5908,N_5631);
and U6504 (N_6504,N_5112,N_5138);
or U6505 (N_6505,N_5012,N_5810);
xnor U6506 (N_6506,N_5487,N_5123);
and U6507 (N_6507,N_5841,N_5096);
xnor U6508 (N_6508,N_5670,N_5739);
nand U6509 (N_6509,N_5439,N_5751);
and U6510 (N_6510,N_5542,N_5998);
nand U6511 (N_6511,N_5934,N_5551);
and U6512 (N_6512,N_5117,N_5543);
nand U6513 (N_6513,N_5470,N_5793);
xnor U6514 (N_6514,N_5493,N_5007);
nor U6515 (N_6515,N_5815,N_5928);
nor U6516 (N_6516,N_5224,N_5296);
and U6517 (N_6517,N_5156,N_5500);
nor U6518 (N_6518,N_5974,N_5182);
xnor U6519 (N_6519,N_5129,N_5460);
nor U6520 (N_6520,N_5619,N_5069);
or U6521 (N_6521,N_5704,N_5734);
xor U6522 (N_6522,N_5456,N_5136);
xor U6523 (N_6523,N_5798,N_5131);
nand U6524 (N_6524,N_5898,N_5428);
nor U6525 (N_6525,N_5311,N_5226);
xor U6526 (N_6526,N_5862,N_5562);
nor U6527 (N_6527,N_5873,N_5159);
and U6528 (N_6528,N_5340,N_5272);
nand U6529 (N_6529,N_5446,N_5458);
xor U6530 (N_6530,N_5627,N_5962);
nor U6531 (N_6531,N_5030,N_5032);
nand U6532 (N_6532,N_5828,N_5547);
or U6533 (N_6533,N_5055,N_5464);
and U6534 (N_6534,N_5657,N_5838);
or U6535 (N_6535,N_5917,N_5846);
and U6536 (N_6536,N_5854,N_5488);
or U6537 (N_6537,N_5425,N_5227);
nor U6538 (N_6538,N_5147,N_5831);
and U6539 (N_6539,N_5316,N_5519);
nor U6540 (N_6540,N_5160,N_5170);
xor U6541 (N_6541,N_5699,N_5688);
or U6542 (N_6542,N_5111,N_5413);
xnor U6543 (N_6543,N_5431,N_5324);
nor U6544 (N_6544,N_5319,N_5190);
or U6545 (N_6545,N_5141,N_5372);
nand U6546 (N_6546,N_5854,N_5168);
nor U6547 (N_6547,N_5246,N_5309);
xor U6548 (N_6548,N_5926,N_5841);
nand U6549 (N_6549,N_5927,N_5485);
nand U6550 (N_6550,N_5116,N_5976);
nand U6551 (N_6551,N_5004,N_5447);
and U6552 (N_6552,N_5125,N_5450);
xor U6553 (N_6553,N_5012,N_5436);
and U6554 (N_6554,N_5586,N_5641);
or U6555 (N_6555,N_5121,N_5790);
and U6556 (N_6556,N_5789,N_5739);
nor U6557 (N_6557,N_5594,N_5482);
and U6558 (N_6558,N_5638,N_5032);
or U6559 (N_6559,N_5711,N_5787);
xnor U6560 (N_6560,N_5725,N_5730);
and U6561 (N_6561,N_5841,N_5525);
nand U6562 (N_6562,N_5233,N_5920);
nand U6563 (N_6563,N_5598,N_5642);
or U6564 (N_6564,N_5815,N_5493);
nor U6565 (N_6565,N_5552,N_5000);
nand U6566 (N_6566,N_5497,N_5074);
nor U6567 (N_6567,N_5677,N_5738);
or U6568 (N_6568,N_5793,N_5388);
or U6569 (N_6569,N_5545,N_5697);
nand U6570 (N_6570,N_5305,N_5515);
nand U6571 (N_6571,N_5986,N_5370);
nand U6572 (N_6572,N_5998,N_5823);
or U6573 (N_6573,N_5522,N_5707);
nor U6574 (N_6574,N_5475,N_5992);
or U6575 (N_6575,N_5195,N_5076);
nor U6576 (N_6576,N_5847,N_5940);
nor U6577 (N_6577,N_5962,N_5204);
nand U6578 (N_6578,N_5568,N_5633);
and U6579 (N_6579,N_5136,N_5012);
nor U6580 (N_6580,N_5533,N_5653);
nand U6581 (N_6581,N_5904,N_5313);
nor U6582 (N_6582,N_5615,N_5854);
nand U6583 (N_6583,N_5977,N_5581);
nand U6584 (N_6584,N_5096,N_5381);
nor U6585 (N_6585,N_5971,N_5185);
nand U6586 (N_6586,N_5117,N_5532);
xnor U6587 (N_6587,N_5174,N_5357);
nor U6588 (N_6588,N_5394,N_5968);
and U6589 (N_6589,N_5381,N_5393);
and U6590 (N_6590,N_5168,N_5761);
nand U6591 (N_6591,N_5054,N_5062);
nor U6592 (N_6592,N_5555,N_5826);
xor U6593 (N_6593,N_5422,N_5190);
nand U6594 (N_6594,N_5180,N_5366);
nand U6595 (N_6595,N_5042,N_5021);
nor U6596 (N_6596,N_5173,N_5504);
nor U6597 (N_6597,N_5904,N_5752);
and U6598 (N_6598,N_5355,N_5795);
xnor U6599 (N_6599,N_5390,N_5787);
and U6600 (N_6600,N_5873,N_5992);
nand U6601 (N_6601,N_5230,N_5155);
nor U6602 (N_6602,N_5802,N_5148);
nand U6603 (N_6603,N_5245,N_5110);
xor U6604 (N_6604,N_5719,N_5531);
nor U6605 (N_6605,N_5834,N_5305);
xnor U6606 (N_6606,N_5484,N_5014);
or U6607 (N_6607,N_5482,N_5426);
or U6608 (N_6608,N_5365,N_5007);
nand U6609 (N_6609,N_5919,N_5531);
nand U6610 (N_6610,N_5756,N_5053);
nand U6611 (N_6611,N_5821,N_5852);
and U6612 (N_6612,N_5496,N_5659);
nor U6613 (N_6613,N_5061,N_5368);
and U6614 (N_6614,N_5810,N_5533);
nand U6615 (N_6615,N_5067,N_5694);
xor U6616 (N_6616,N_5234,N_5493);
or U6617 (N_6617,N_5732,N_5389);
xor U6618 (N_6618,N_5517,N_5677);
and U6619 (N_6619,N_5130,N_5400);
nand U6620 (N_6620,N_5302,N_5672);
nand U6621 (N_6621,N_5432,N_5829);
and U6622 (N_6622,N_5839,N_5403);
nand U6623 (N_6623,N_5072,N_5514);
nand U6624 (N_6624,N_5388,N_5301);
xnor U6625 (N_6625,N_5018,N_5901);
nand U6626 (N_6626,N_5808,N_5361);
or U6627 (N_6627,N_5751,N_5276);
or U6628 (N_6628,N_5014,N_5921);
and U6629 (N_6629,N_5280,N_5861);
and U6630 (N_6630,N_5357,N_5806);
nand U6631 (N_6631,N_5226,N_5274);
nor U6632 (N_6632,N_5154,N_5016);
nand U6633 (N_6633,N_5414,N_5510);
nor U6634 (N_6634,N_5864,N_5034);
xnor U6635 (N_6635,N_5904,N_5612);
or U6636 (N_6636,N_5288,N_5565);
and U6637 (N_6637,N_5843,N_5241);
and U6638 (N_6638,N_5359,N_5465);
nand U6639 (N_6639,N_5071,N_5413);
xor U6640 (N_6640,N_5619,N_5410);
xnor U6641 (N_6641,N_5847,N_5392);
or U6642 (N_6642,N_5566,N_5344);
nand U6643 (N_6643,N_5687,N_5430);
xnor U6644 (N_6644,N_5114,N_5549);
nor U6645 (N_6645,N_5373,N_5326);
xnor U6646 (N_6646,N_5618,N_5260);
and U6647 (N_6647,N_5261,N_5983);
or U6648 (N_6648,N_5366,N_5955);
xnor U6649 (N_6649,N_5305,N_5596);
nand U6650 (N_6650,N_5588,N_5719);
or U6651 (N_6651,N_5457,N_5630);
and U6652 (N_6652,N_5601,N_5930);
or U6653 (N_6653,N_5107,N_5316);
xor U6654 (N_6654,N_5469,N_5759);
nor U6655 (N_6655,N_5697,N_5350);
nor U6656 (N_6656,N_5002,N_5101);
and U6657 (N_6657,N_5952,N_5280);
nor U6658 (N_6658,N_5796,N_5675);
nand U6659 (N_6659,N_5197,N_5082);
and U6660 (N_6660,N_5684,N_5317);
and U6661 (N_6661,N_5574,N_5939);
or U6662 (N_6662,N_5796,N_5169);
and U6663 (N_6663,N_5948,N_5180);
and U6664 (N_6664,N_5221,N_5504);
and U6665 (N_6665,N_5756,N_5920);
or U6666 (N_6666,N_5090,N_5926);
and U6667 (N_6667,N_5085,N_5570);
nand U6668 (N_6668,N_5635,N_5638);
nand U6669 (N_6669,N_5997,N_5533);
nand U6670 (N_6670,N_5415,N_5069);
and U6671 (N_6671,N_5735,N_5761);
nor U6672 (N_6672,N_5356,N_5624);
or U6673 (N_6673,N_5953,N_5996);
and U6674 (N_6674,N_5065,N_5457);
or U6675 (N_6675,N_5190,N_5197);
nand U6676 (N_6676,N_5142,N_5262);
xnor U6677 (N_6677,N_5906,N_5636);
nand U6678 (N_6678,N_5189,N_5078);
and U6679 (N_6679,N_5129,N_5148);
or U6680 (N_6680,N_5168,N_5510);
nand U6681 (N_6681,N_5103,N_5508);
and U6682 (N_6682,N_5424,N_5521);
nor U6683 (N_6683,N_5226,N_5500);
and U6684 (N_6684,N_5786,N_5925);
and U6685 (N_6685,N_5741,N_5080);
nand U6686 (N_6686,N_5658,N_5232);
nand U6687 (N_6687,N_5390,N_5929);
nand U6688 (N_6688,N_5269,N_5824);
nand U6689 (N_6689,N_5783,N_5096);
nor U6690 (N_6690,N_5723,N_5351);
nand U6691 (N_6691,N_5747,N_5968);
nand U6692 (N_6692,N_5464,N_5296);
xnor U6693 (N_6693,N_5512,N_5745);
xnor U6694 (N_6694,N_5629,N_5626);
or U6695 (N_6695,N_5933,N_5258);
xnor U6696 (N_6696,N_5177,N_5093);
and U6697 (N_6697,N_5745,N_5805);
nor U6698 (N_6698,N_5386,N_5445);
nand U6699 (N_6699,N_5405,N_5378);
xor U6700 (N_6700,N_5611,N_5095);
nand U6701 (N_6701,N_5121,N_5926);
xor U6702 (N_6702,N_5453,N_5716);
nand U6703 (N_6703,N_5301,N_5783);
nor U6704 (N_6704,N_5322,N_5970);
nor U6705 (N_6705,N_5842,N_5957);
xor U6706 (N_6706,N_5571,N_5227);
nor U6707 (N_6707,N_5640,N_5965);
or U6708 (N_6708,N_5681,N_5888);
nand U6709 (N_6709,N_5906,N_5943);
and U6710 (N_6710,N_5216,N_5573);
and U6711 (N_6711,N_5120,N_5712);
nor U6712 (N_6712,N_5341,N_5876);
nor U6713 (N_6713,N_5531,N_5605);
or U6714 (N_6714,N_5658,N_5755);
xor U6715 (N_6715,N_5246,N_5674);
nand U6716 (N_6716,N_5356,N_5072);
xor U6717 (N_6717,N_5015,N_5387);
or U6718 (N_6718,N_5346,N_5092);
and U6719 (N_6719,N_5507,N_5707);
nor U6720 (N_6720,N_5165,N_5187);
and U6721 (N_6721,N_5323,N_5925);
or U6722 (N_6722,N_5724,N_5721);
nand U6723 (N_6723,N_5577,N_5602);
xnor U6724 (N_6724,N_5774,N_5792);
or U6725 (N_6725,N_5649,N_5660);
xnor U6726 (N_6726,N_5177,N_5195);
nand U6727 (N_6727,N_5937,N_5576);
nand U6728 (N_6728,N_5521,N_5005);
nand U6729 (N_6729,N_5447,N_5920);
or U6730 (N_6730,N_5205,N_5762);
xnor U6731 (N_6731,N_5366,N_5178);
and U6732 (N_6732,N_5412,N_5830);
xor U6733 (N_6733,N_5526,N_5761);
nand U6734 (N_6734,N_5199,N_5005);
and U6735 (N_6735,N_5320,N_5074);
and U6736 (N_6736,N_5866,N_5280);
xnor U6737 (N_6737,N_5775,N_5849);
nor U6738 (N_6738,N_5659,N_5037);
or U6739 (N_6739,N_5488,N_5323);
xor U6740 (N_6740,N_5174,N_5007);
xnor U6741 (N_6741,N_5099,N_5921);
or U6742 (N_6742,N_5871,N_5544);
nand U6743 (N_6743,N_5464,N_5762);
or U6744 (N_6744,N_5705,N_5889);
and U6745 (N_6745,N_5626,N_5846);
nor U6746 (N_6746,N_5780,N_5381);
xnor U6747 (N_6747,N_5535,N_5010);
nor U6748 (N_6748,N_5375,N_5086);
or U6749 (N_6749,N_5533,N_5999);
xor U6750 (N_6750,N_5621,N_5896);
nand U6751 (N_6751,N_5272,N_5900);
nor U6752 (N_6752,N_5826,N_5283);
or U6753 (N_6753,N_5985,N_5433);
xor U6754 (N_6754,N_5682,N_5484);
nand U6755 (N_6755,N_5690,N_5780);
nand U6756 (N_6756,N_5835,N_5920);
nor U6757 (N_6757,N_5713,N_5295);
nor U6758 (N_6758,N_5141,N_5107);
and U6759 (N_6759,N_5832,N_5162);
nand U6760 (N_6760,N_5651,N_5792);
nor U6761 (N_6761,N_5139,N_5634);
or U6762 (N_6762,N_5826,N_5388);
nor U6763 (N_6763,N_5229,N_5261);
xnor U6764 (N_6764,N_5933,N_5024);
nor U6765 (N_6765,N_5642,N_5215);
nand U6766 (N_6766,N_5884,N_5857);
nand U6767 (N_6767,N_5473,N_5877);
xor U6768 (N_6768,N_5668,N_5938);
or U6769 (N_6769,N_5269,N_5733);
or U6770 (N_6770,N_5076,N_5122);
xor U6771 (N_6771,N_5889,N_5346);
or U6772 (N_6772,N_5696,N_5625);
nand U6773 (N_6773,N_5104,N_5201);
nand U6774 (N_6774,N_5592,N_5323);
nand U6775 (N_6775,N_5707,N_5244);
or U6776 (N_6776,N_5555,N_5938);
and U6777 (N_6777,N_5789,N_5779);
and U6778 (N_6778,N_5346,N_5249);
nand U6779 (N_6779,N_5690,N_5946);
or U6780 (N_6780,N_5827,N_5050);
and U6781 (N_6781,N_5385,N_5163);
nor U6782 (N_6782,N_5200,N_5017);
or U6783 (N_6783,N_5348,N_5200);
or U6784 (N_6784,N_5835,N_5905);
and U6785 (N_6785,N_5167,N_5025);
or U6786 (N_6786,N_5335,N_5984);
nand U6787 (N_6787,N_5924,N_5407);
nor U6788 (N_6788,N_5953,N_5132);
and U6789 (N_6789,N_5017,N_5673);
xor U6790 (N_6790,N_5422,N_5407);
xnor U6791 (N_6791,N_5074,N_5829);
nand U6792 (N_6792,N_5366,N_5827);
nand U6793 (N_6793,N_5018,N_5936);
nor U6794 (N_6794,N_5775,N_5134);
and U6795 (N_6795,N_5897,N_5094);
and U6796 (N_6796,N_5547,N_5186);
nor U6797 (N_6797,N_5989,N_5112);
nor U6798 (N_6798,N_5312,N_5555);
and U6799 (N_6799,N_5837,N_5223);
and U6800 (N_6800,N_5686,N_5704);
xnor U6801 (N_6801,N_5393,N_5067);
nand U6802 (N_6802,N_5481,N_5071);
and U6803 (N_6803,N_5202,N_5450);
and U6804 (N_6804,N_5397,N_5012);
xor U6805 (N_6805,N_5608,N_5222);
xor U6806 (N_6806,N_5014,N_5057);
and U6807 (N_6807,N_5344,N_5826);
or U6808 (N_6808,N_5381,N_5497);
or U6809 (N_6809,N_5324,N_5797);
or U6810 (N_6810,N_5109,N_5087);
nor U6811 (N_6811,N_5936,N_5993);
and U6812 (N_6812,N_5478,N_5543);
nand U6813 (N_6813,N_5109,N_5700);
or U6814 (N_6814,N_5162,N_5151);
xnor U6815 (N_6815,N_5848,N_5429);
or U6816 (N_6816,N_5895,N_5387);
and U6817 (N_6817,N_5475,N_5431);
and U6818 (N_6818,N_5254,N_5382);
or U6819 (N_6819,N_5738,N_5823);
or U6820 (N_6820,N_5361,N_5909);
nand U6821 (N_6821,N_5287,N_5581);
nand U6822 (N_6822,N_5980,N_5525);
xor U6823 (N_6823,N_5867,N_5880);
nor U6824 (N_6824,N_5152,N_5718);
nor U6825 (N_6825,N_5359,N_5136);
xnor U6826 (N_6826,N_5140,N_5733);
and U6827 (N_6827,N_5398,N_5372);
nand U6828 (N_6828,N_5525,N_5937);
and U6829 (N_6829,N_5334,N_5929);
nor U6830 (N_6830,N_5702,N_5934);
nand U6831 (N_6831,N_5633,N_5657);
or U6832 (N_6832,N_5528,N_5456);
and U6833 (N_6833,N_5480,N_5125);
and U6834 (N_6834,N_5010,N_5883);
xnor U6835 (N_6835,N_5039,N_5234);
nor U6836 (N_6836,N_5570,N_5264);
or U6837 (N_6837,N_5972,N_5055);
and U6838 (N_6838,N_5777,N_5146);
xor U6839 (N_6839,N_5419,N_5610);
or U6840 (N_6840,N_5985,N_5439);
xnor U6841 (N_6841,N_5521,N_5034);
xnor U6842 (N_6842,N_5257,N_5937);
nor U6843 (N_6843,N_5032,N_5144);
nor U6844 (N_6844,N_5835,N_5492);
xor U6845 (N_6845,N_5495,N_5845);
or U6846 (N_6846,N_5868,N_5341);
or U6847 (N_6847,N_5456,N_5443);
nor U6848 (N_6848,N_5574,N_5234);
xor U6849 (N_6849,N_5563,N_5680);
xor U6850 (N_6850,N_5322,N_5386);
and U6851 (N_6851,N_5311,N_5691);
and U6852 (N_6852,N_5047,N_5363);
nand U6853 (N_6853,N_5298,N_5803);
nor U6854 (N_6854,N_5213,N_5093);
nor U6855 (N_6855,N_5568,N_5825);
nand U6856 (N_6856,N_5592,N_5238);
and U6857 (N_6857,N_5233,N_5558);
nor U6858 (N_6858,N_5600,N_5592);
xnor U6859 (N_6859,N_5960,N_5989);
or U6860 (N_6860,N_5295,N_5701);
xnor U6861 (N_6861,N_5015,N_5298);
nand U6862 (N_6862,N_5630,N_5824);
nand U6863 (N_6863,N_5099,N_5234);
nor U6864 (N_6864,N_5644,N_5525);
xor U6865 (N_6865,N_5988,N_5466);
or U6866 (N_6866,N_5065,N_5537);
nor U6867 (N_6867,N_5681,N_5475);
or U6868 (N_6868,N_5662,N_5842);
nor U6869 (N_6869,N_5251,N_5420);
xor U6870 (N_6870,N_5742,N_5202);
xor U6871 (N_6871,N_5077,N_5380);
and U6872 (N_6872,N_5234,N_5654);
or U6873 (N_6873,N_5061,N_5601);
xnor U6874 (N_6874,N_5234,N_5002);
and U6875 (N_6875,N_5895,N_5253);
nand U6876 (N_6876,N_5693,N_5190);
nand U6877 (N_6877,N_5936,N_5020);
or U6878 (N_6878,N_5817,N_5336);
xnor U6879 (N_6879,N_5869,N_5899);
xor U6880 (N_6880,N_5829,N_5547);
or U6881 (N_6881,N_5232,N_5596);
xnor U6882 (N_6882,N_5407,N_5836);
nor U6883 (N_6883,N_5920,N_5064);
or U6884 (N_6884,N_5093,N_5597);
nand U6885 (N_6885,N_5626,N_5855);
nor U6886 (N_6886,N_5406,N_5405);
nor U6887 (N_6887,N_5591,N_5011);
nand U6888 (N_6888,N_5551,N_5748);
or U6889 (N_6889,N_5983,N_5359);
nand U6890 (N_6890,N_5662,N_5889);
nand U6891 (N_6891,N_5911,N_5143);
xor U6892 (N_6892,N_5728,N_5426);
and U6893 (N_6893,N_5722,N_5275);
xor U6894 (N_6894,N_5506,N_5658);
or U6895 (N_6895,N_5381,N_5657);
xor U6896 (N_6896,N_5826,N_5357);
and U6897 (N_6897,N_5746,N_5834);
nor U6898 (N_6898,N_5377,N_5957);
nand U6899 (N_6899,N_5325,N_5757);
and U6900 (N_6900,N_5834,N_5506);
nand U6901 (N_6901,N_5719,N_5502);
and U6902 (N_6902,N_5926,N_5489);
or U6903 (N_6903,N_5012,N_5054);
and U6904 (N_6904,N_5541,N_5044);
xor U6905 (N_6905,N_5797,N_5827);
nor U6906 (N_6906,N_5440,N_5813);
and U6907 (N_6907,N_5448,N_5189);
nand U6908 (N_6908,N_5572,N_5630);
xnor U6909 (N_6909,N_5090,N_5315);
nor U6910 (N_6910,N_5406,N_5508);
or U6911 (N_6911,N_5291,N_5611);
nand U6912 (N_6912,N_5723,N_5229);
nand U6913 (N_6913,N_5155,N_5832);
nand U6914 (N_6914,N_5641,N_5510);
xor U6915 (N_6915,N_5339,N_5655);
nand U6916 (N_6916,N_5375,N_5760);
nand U6917 (N_6917,N_5276,N_5860);
nor U6918 (N_6918,N_5208,N_5531);
and U6919 (N_6919,N_5423,N_5863);
xnor U6920 (N_6920,N_5417,N_5976);
xor U6921 (N_6921,N_5754,N_5998);
nand U6922 (N_6922,N_5920,N_5825);
nand U6923 (N_6923,N_5381,N_5198);
nor U6924 (N_6924,N_5376,N_5995);
xor U6925 (N_6925,N_5798,N_5635);
or U6926 (N_6926,N_5291,N_5007);
or U6927 (N_6927,N_5112,N_5003);
and U6928 (N_6928,N_5755,N_5143);
nor U6929 (N_6929,N_5580,N_5756);
xnor U6930 (N_6930,N_5165,N_5644);
xor U6931 (N_6931,N_5780,N_5330);
or U6932 (N_6932,N_5100,N_5044);
and U6933 (N_6933,N_5071,N_5679);
xor U6934 (N_6934,N_5385,N_5991);
nor U6935 (N_6935,N_5163,N_5307);
nor U6936 (N_6936,N_5595,N_5883);
xor U6937 (N_6937,N_5547,N_5622);
xnor U6938 (N_6938,N_5000,N_5286);
nand U6939 (N_6939,N_5624,N_5780);
and U6940 (N_6940,N_5539,N_5819);
xor U6941 (N_6941,N_5109,N_5674);
xnor U6942 (N_6942,N_5534,N_5676);
nor U6943 (N_6943,N_5238,N_5099);
and U6944 (N_6944,N_5481,N_5337);
and U6945 (N_6945,N_5458,N_5037);
nand U6946 (N_6946,N_5476,N_5706);
xor U6947 (N_6947,N_5056,N_5842);
nor U6948 (N_6948,N_5628,N_5652);
or U6949 (N_6949,N_5160,N_5207);
or U6950 (N_6950,N_5309,N_5307);
and U6951 (N_6951,N_5685,N_5930);
or U6952 (N_6952,N_5109,N_5130);
nand U6953 (N_6953,N_5567,N_5311);
or U6954 (N_6954,N_5100,N_5351);
or U6955 (N_6955,N_5100,N_5359);
xor U6956 (N_6956,N_5935,N_5601);
and U6957 (N_6957,N_5218,N_5354);
and U6958 (N_6958,N_5760,N_5720);
and U6959 (N_6959,N_5700,N_5377);
or U6960 (N_6960,N_5385,N_5570);
nand U6961 (N_6961,N_5293,N_5019);
or U6962 (N_6962,N_5254,N_5701);
xnor U6963 (N_6963,N_5472,N_5876);
nand U6964 (N_6964,N_5088,N_5552);
nand U6965 (N_6965,N_5048,N_5938);
xnor U6966 (N_6966,N_5786,N_5959);
xnor U6967 (N_6967,N_5062,N_5235);
nor U6968 (N_6968,N_5009,N_5720);
xnor U6969 (N_6969,N_5441,N_5295);
nor U6970 (N_6970,N_5817,N_5257);
or U6971 (N_6971,N_5406,N_5750);
xnor U6972 (N_6972,N_5687,N_5711);
and U6973 (N_6973,N_5143,N_5715);
or U6974 (N_6974,N_5928,N_5932);
and U6975 (N_6975,N_5050,N_5934);
or U6976 (N_6976,N_5449,N_5234);
nor U6977 (N_6977,N_5906,N_5507);
or U6978 (N_6978,N_5273,N_5027);
nand U6979 (N_6979,N_5665,N_5440);
nor U6980 (N_6980,N_5803,N_5425);
and U6981 (N_6981,N_5290,N_5746);
nor U6982 (N_6982,N_5824,N_5083);
or U6983 (N_6983,N_5421,N_5350);
nand U6984 (N_6984,N_5833,N_5663);
nand U6985 (N_6985,N_5704,N_5332);
and U6986 (N_6986,N_5579,N_5033);
and U6987 (N_6987,N_5252,N_5524);
nand U6988 (N_6988,N_5069,N_5566);
xnor U6989 (N_6989,N_5909,N_5006);
and U6990 (N_6990,N_5613,N_5352);
xnor U6991 (N_6991,N_5575,N_5604);
nor U6992 (N_6992,N_5880,N_5069);
and U6993 (N_6993,N_5083,N_5366);
nand U6994 (N_6994,N_5755,N_5494);
or U6995 (N_6995,N_5060,N_5190);
xnor U6996 (N_6996,N_5951,N_5520);
nand U6997 (N_6997,N_5523,N_5669);
and U6998 (N_6998,N_5184,N_5023);
nor U6999 (N_6999,N_5395,N_5306);
or U7000 (N_7000,N_6838,N_6769);
nor U7001 (N_7001,N_6843,N_6228);
nand U7002 (N_7002,N_6363,N_6706);
and U7003 (N_7003,N_6752,N_6933);
or U7004 (N_7004,N_6627,N_6795);
or U7005 (N_7005,N_6175,N_6349);
xnor U7006 (N_7006,N_6165,N_6982);
nand U7007 (N_7007,N_6132,N_6648);
nand U7008 (N_7008,N_6857,N_6057);
xnor U7009 (N_7009,N_6343,N_6521);
and U7010 (N_7010,N_6341,N_6190);
and U7011 (N_7011,N_6764,N_6474);
nand U7012 (N_7012,N_6002,N_6261);
nand U7013 (N_7013,N_6911,N_6849);
nand U7014 (N_7014,N_6784,N_6288);
nand U7015 (N_7015,N_6802,N_6616);
and U7016 (N_7016,N_6400,N_6948);
and U7017 (N_7017,N_6763,N_6799);
xnor U7018 (N_7018,N_6021,N_6354);
xnor U7019 (N_7019,N_6301,N_6973);
nor U7020 (N_7020,N_6609,N_6456);
or U7021 (N_7021,N_6526,N_6153);
or U7022 (N_7022,N_6922,N_6086);
xnor U7023 (N_7023,N_6852,N_6280);
nor U7024 (N_7024,N_6307,N_6404);
xnor U7025 (N_7025,N_6437,N_6567);
or U7026 (N_7026,N_6104,N_6658);
xnor U7027 (N_7027,N_6940,N_6191);
and U7028 (N_7028,N_6846,N_6075);
or U7029 (N_7029,N_6388,N_6666);
xor U7030 (N_7030,N_6428,N_6408);
xnor U7031 (N_7031,N_6503,N_6826);
or U7032 (N_7032,N_6558,N_6957);
and U7033 (N_7033,N_6767,N_6020);
nor U7034 (N_7034,N_6461,N_6482);
and U7035 (N_7035,N_6485,N_6099);
xnor U7036 (N_7036,N_6705,N_6903);
xnor U7037 (N_7037,N_6087,N_6987);
nand U7038 (N_7038,N_6961,N_6779);
and U7039 (N_7039,N_6610,N_6675);
nand U7040 (N_7040,N_6007,N_6284);
and U7041 (N_7041,N_6774,N_6860);
xnor U7042 (N_7042,N_6770,N_6833);
nand U7043 (N_7043,N_6394,N_6986);
nor U7044 (N_7044,N_6757,N_6197);
nand U7045 (N_7045,N_6832,N_6152);
and U7046 (N_7046,N_6547,N_6629);
and U7047 (N_7047,N_6976,N_6006);
nor U7048 (N_7048,N_6393,N_6936);
and U7049 (N_7049,N_6595,N_6645);
xor U7050 (N_7050,N_6239,N_6525);
xor U7051 (N_7051,N_6513,N_6469);
xor U7052 (N_7052,N_6670,N_6907);
and U7053 (N_7053,N_6070,N_6088);
or U7054 (N_7054,N_6704,N_6192);
and U7055 (N_7055,N_6917,N_6946);
xnor U7056 (N_7056,N_6336,N_6359);
nand U7057 (N_7057,N_6156,N_6602);
or U7058 (N_7058,N_6108,N_6722);
xnor U7059 (N_7059,N_6096,N_6800);
or U7060 (N_7060,N_6279,N_6494);
nor U7061 (N_7061,N_6150,N_6155);
and U7062 (N_7062,N_6443,N_6240);
nand U7063 (N_7063,N_6095,N_6506);
nand U7064 (N_7064,N_6939,N_6992);
nor U7065 (N_7065,N_6980,N_6822);
nor U7066 (N_7066,N_6138,N_6326);
xnor U7067 (N_7067,N_6141,N_6251);
and U7068 (N_7068,N_6131,N_6264);
and U7069 (N_7069,N_6032,N_6081);
or U7070 (N_7070,N_6355,N_6632);
nand U7071 (N_7071,N_6956,N_6908);
and U7072 (N_7072,N_6058,N_6783);
nand U7073 (N_7073,N_6805,N_6452);
nor U7074 (N_7074,N_6013,N_6944);
nor U7075 (N_7075,N_6290,N_6892);
and U7076 (N_7076,N_6089,N_6630);
xor U7077 (N_7077,N_6129,N_6215);
or U7078 (N_7078,N_6734,N_6615);
nand U7079 (N_7079,N_6820,N_6738);
or U7080 (N_7080,N_6473,N_6386);
nor U7081 (N_7081,N_6119,N_6247);
xnor U7082 (N_7082,N_6528,N_6694);
nor U7083 (N_7083,N_6827,N_6662);
nand U7084 (N_7084,N_6835,N_6342);
nand U7085 (N_7085,N_6146,N_6222);
nor U7086 (N_7086,N_6829,N_6367);
xor U7087 (N_7087,N_6901,N_6399);
or U7088 (N_7088,N_6902,N_6000);
nand U7089 (N_7089,N_6049,N_6125);
or U7090 (N_7090,N_6894,N_6193);
nor U7091 (N_7091,N_6453,N_6847);
nor U7092 (N_7092,N_6999,N_6967);
nor U7093 (N_7093,N_6597,N_6082);
and U7094 (N_7094,N_6330,N_6929);
nand U7095 (N_7095,N_6712,N_6899);
nand U7096 (N_7096,N_6954,N_6268);
or U7097 (N_7097,N_6504,N_6586);
or U7098 (N_7098,N_6210,N_6126);
nor U7099 (N_7099,N_6373,N_6711);
nor U7100 (N_7100,N_6876,N_6390);
nand U7101 (N_7101,N_6703,N_6733);
xor U7102 (N_7102,N_6566,N_6025);
and U7103 (N_7103,N_6942,N_6411);
and U7104 (N_7104,N_6989,N_6376);
xnor U7105 (N_7105,N_6867,N_6242);
nor U7106 (N_7106,N_6368,N_6008);
and U7107 (N_7107,N_6549,N_6172);
xnor U7108 (N_7108,N_6497,N_6934);
nand U7109 (N_7109,N_6671,N_6766);
and U7110 (N_7110,N_6270,N_6551);
and U7111 (N_7111,N_6366,N_6231);
nor U7112 (N_7112,N_6890,N_6729);
xnor U7113 (N_7113,N_6979,N_6932);
nor U7114 (N_7114,N_6457,N_6718);
nand U7115 (N_7115,N_6338,N_6224);
or U7116 (N_7116,N_6971,N_6323);
nor U7117 (N_7117,N_6825,N_6953);
nand U7118 (N_7118,N_6183,N_6962);
and U7119 (N_7119,N_6026,N_6604);
and U7120 (N_7120,N_6797,N_6077);
nand U7121 (N_7121,N_6518,N_6047);
xor U7122 (N_7122,N_6362,N_6332);
or U7123 (N_7123,N_6158,N_6448);
nand U7124 (N_7124,N_6421,N_6552);
or U7125 (N_7125,N_6765,N_6990);
or U7126 (N_7126,N_6195,N_6855);
or U7127 (N_7127,N_6599,N_6257);
nor U7128 (N_7128,N_6955,N_6885);
and U7129 (N_7129,N_6993,N_6382);
xnor U7130 (N_7130,N_6776,N_6164);
xor U7131 (N_7131,N_6003,N_6378);
and U7132 (N_7132,N_6441,N_6161);
nand U7133 (N_7133,N_6643,N_6294);
and U7134 (N_7134,N_6888,N_6500);
or U7135 (N_7135,N_6947,N_6751);
or U7136 (N_7136,N_6277,N_6364);
nor U7137 (N_7137,N_6546,N_6012);
nor U7138 (N_7138,N_6325,N_6842);
nand U7139 (N_7139,N_6344,N_6634);
or U7140 (N_7140,N_6199,N_6848);
xor U7141 (N_7141,N_6068,N_6550);
xor U7142 (N_7142,N_6964,N_6311);
and U7143 (N_7143,N_6501,N_6432);
nand U7144 (N_7144,N_6059,N_6837);
and U7145 (N_7145,N_6928,N_6109);
or U7146 (N_7146,N_6435,N_6185);
nor U7147 (N_7147,N_6879,N_6154);
xnor U7148 (N_7148,N_6203,N_6022);
and U7149 (N_7149,N_6010,N_6238);
nand U7150 (N_7150,N_6085,N_6561);
nand U7151 (N_7151,N_6935,N_6815);
nor U7152 (N_7152,N_6173,N_6710);
and U7153 (N_7153,N_6789,N_6969);
or U7154 (N_7154,N_6282,N_6673);
or U7155 (N_7155,N_6912,N_6353);
and U7156 (N_7156,N_6530,N_6786);
or U7157 (N_7157,N_6650,N_6202);
nor U7158 (N_7158,N_6465,N_6061);
and U7159 (N_7159,N_6794,N_6396);
xor U7160 (N_7160,N_6346,N_6103);
or U7161 (N_7161,N_6620,N_6681);
xor U7162 (N_7162,N_6592,N_6920);
nor U7163 (N_7163,N_6896,N_6758);
xnor U7164 (N_7164,N_6591,N_6853);
nor U7165 (N_7165,N_6340,N_6925);
xor U7166 (N_7166,N_6237,N_6479);
or U7167 (N_7167,N_6747,N_6335);
xnor U7168 (N_7168,N_6106,N_6813);
or U7169 (N_7169,N_6196,N_6149);
nand U7170 (N_7170,N_6863,N_6029);
or U7171 (N_7171,N_6123,N_6413);
nand U7172 (N_7172,N_6223,N_6900);
and U7173 (N_7173,N_6112,N_6559);
and U7174 (N_7174,N_6931,N_6182);
nor U7175 (N_7175,N_6255,N_6537);
or U7176 (N_7176,N_6523,N_6339);
xor U7177 (N_7177,N_6484,N_6717);
nand U7178 (N_7178,N_6489,N_6889);
nand U7179 (N_7179,N_6587,N_6520);
nor U7180 (N_7180,N_6067,N_6785);
xor U7181 (N_7181,N_6248,N_6039);
nand U7182 (N_7182,N_6701,N_6881);
or U7183 (N_7183,N_6180,N_6229);
nand U7184 (N_7184,N_6572,N_6157);
nor U7185 (N_7185,N_6069,N_6854);
nand U7186 (N_7186,N_6601,N_6514);
nand U7187 (N_7187,N_6403,N_6177);
xnor U7188 (N_7188,N_6563,N_6118);
nor U7189 (N_7189,N_6291,N_6914);
and U7190 (N_7190,N_6950,N_6628);
xnor U7191 (N_7191,N_6972,N_6236);
and U7192 (N_7192,N_6416,N_6578);
nor U7193 (N_7193,N_6759,N_6593);
or U7194 (N_7194,N_6674,N_6545);
nor U7195 (N_7195,N_6166,N_6415);
or U7196 (N_7196,N_6100,N_6619);
nor U7197 (N_7197,N_6467,N_6678);
or U7198 (N_7198,N_6211,N_6318);
nor U7199 (N_7199,N_6997,N_6614);
and U7200 (N_7200,N_6137,N_6806);
nor U7201 (N_7201,N_6517,N_6535);
xor U7202 (N_7202,N_6205,N_6577);
nand U7203 (N_7203,N_6027,N_6996);
or U7204 (N_7204,N_6375,N_6269);
xnor U7205 (N_7205,N_6680,N_6808);
and U7206 (N_7206,N_6834,N_6234);
nand U7207 (N_7207,N_6637,N_6055);
xnor U7208 (N_7208,N_6913,N_6796);
xor U7209 (N_7209,N_6389,N_6543);
nor U7210 (N_7210,N_6062,N_6760);
xnor U7211 (N_7211,N_6444,N_6975);
nor U7212 (N_7212,N_6212,N_6791);
xor U7213 (N_7213,N_6033,N_6668);
nand U7214 (N_7214,N_6427,N_6720);
nor U7215 (N_7215,N_6723,N_6730);
xnor U7216 (N_7216,N_6357,N_6244);
xor U7217 (N_7217,N_6669,N_6691);
xnor U7218 (N_7218,N_6893,N_6046);
nor U7219 (N_7219,N_6207,N_6097);
and U7220 (N_7220,N_6447,N_6748);
nor U7221 (N_7221,N_6065,N_6882);
xor U7222 (N_7222,N_6927,N_6746);
nand U7223 (N_7223,N_6721,N_6449);
or U7224 (N_7224,N_6001,N_6557);
or U7225 (N_7225,N_6869,N_6135);
nor U7226 (N_7226,N_6371,N_6841);
nor U7227 (N_7227,N_6657,N_6206);
xnor U7228 (N_7228,N_6387,N_6700);
nand U7229 (N_7229,N_6483,N_6582);
nor U7230 (N_7230,N_6866,N_6218);
xnor U7231 (N_7231,N_6468,N_6436);
xnor U7232 (N_7232,N_6128,N_6225);
or U7233 (N_7233,N_6380,N_6804);
or U7234 (N_7234,N_6873,N_6639);
xnor U7235 (N_7235,N_6807,N_6686);
or U7236 (N_7236,N_6877,N_6454);
nor U7237 (N_7237,N_6644,N_6677);
and U7238 (N_7238,N_6810,N_6124);
and U7239 (N_7239,N_6665,N_6633);
nand U7240 (N_7240,N_6379,N_6308);
or U7241 (N_7241,N_6423,N_6726);
xnor U7242 (N_7242,N_6781,N_6170);
or U7243 (N_7243,N_6310,N_6048);
or U7244 (N_7244,N_6606,N_6725);
nand U7245 (N_7245,N_6286,N_6926);
or U7246 (N_7246,N_6740,N_6798);
xnor U7247 (N_7247,N_6272,N_6213);
or U7248 (N_7248,N_6130,N_6856);
and U7249 (N_7249,N_6419,N_6351);
nor U7250 (N_7250,N_6188,N_6060);
and U7251 (N_7251,N_6392,N_6475);
xor U7252 (N_7252,N_6836,N_6121);
nand U7253 (N_7253,N_6816,N_6564);
and U7254 (N_7254,N_6983,N_6439);
or U7255 (N_7255,N_6037,N_6023);
and U7256 (N_7256,N_6412,N_6470);
or U7257 (N_7257,N_6043,N_6898);
nor U7258 (N_7258,N_6556,N_6050);
nand U7259 (N_7259,N_6744,N_6515);
or U7260 (N_7260,N_6731,N_6451);
and U7261 (N_7261,N_6107,N_6005);
and U7262 (N_7262,N_6642,N_6321);
or U7263 (N_7263,N_6576,N_6736);
or U7264 (N_7264,N_6245,N_6555);
nand U7265 (N_7265,N_6117,N_6656);
nor U7266 (N_7266,N_6937,N_6793);
or U7267 (N_7267,N_6148,N_6063);
and U7268 (N_7268,N_6554,N_6274);
xnor U7269 (N_7269,N_6493,N_6790);
or U7270 (N_7270,N_6072,N_6951);
and U7271 (N_7271,N_6184,N_6178);
nor U7272 (N_7272,N_6529,N_6612);
nor U7273 (N_7273,N_6622,N_6455);
or U7274 (N_7274,N_6750,N_6312);
nand U7275 (N_7275,N_6350,N_6187);
nor U7276 (N_7276,N_6011,N_6424);
and U7277 (N_7277,N_6028,N_6963);
or U7278 (N_7278,N_6418,N_6036);
nand U7279 (N_7279,N_6462,N_6374);
nor U7280 (N_7280,N_6271,N_6683);
or U7281 (N_7281,N_6626,N_6256);
or U7282 (N_7282,N_6004,N_6709);
xnor U7283 (N_7283,N_6625,N_6544);
nand U7284 (N_7284,N_6923,N_6283);
nand U7285 (N_7285,N_6801,N_6053);
or U7286 (N_7286,N_6079,N_6263);
nor U7287 (N_7287,N_6676,N_6016);
xor U7288 (N_7288,N_6646,N_6233);
or U7289 (N_7289,N_6243,N_6420);
nand U7290 (N_7290,N_6631,N_6538);
nor U7291 (N_7291,N_6753,N_6333);
nor U7292 (N_7292,N_6814,N_6787);
xnor U7293 (N_7293,N_6488,N_6120);
or U7294 (N_7294,N_6111,N_6699);
nand U7295 (N_7295,N_6741,N_6431);
and U7296 (N_7296,N_6293,N_6071);
or U7297 (N_7297,N_6830,N_6450);
or U7298 (N_7298,N_6041,N_6425);
or U7299 (N_7299,N_6246,N_6573);
nor U7300 (N_7300,N_6414,N_6078);
nor U7301 (N_7301,N_6695,N_6635);
xnor U7302 (N_7302,N_6162,N_6970);
or U7303 (N_7303,N_6780,N_6383);
nand U7304 (N_7304,N_6275,N_6958);
nand U7305 (N_7305,N_6285,N_6044);
and U7306 (N_7306,N_6697,N_6916);
or U7307 (N_7307,N_6636,N_6875);
nor U7308 (N_7308,N_6745,N_6689);
or U7309 (N_7309,N_6426,N_6306);
xor U7310 (N_7310,N_6859,N_6490);
xor U7311 (N_7311,N_6713,N_6788);
and U7312 (N_7312,N_6904,N_6941);
or U7313 (N_7313,N_6527,N_6994);
and U7314 (N_7314,N_6698,N_6569);
and U7315 (N_7315,N_6589,N_6874);
and U7316 (N_7316,N_6562,N_6507);
xor U7317 (N_7317,N_6724,N_6080);
and U7318 (N_7318,N_6716,N_6254);
or U7319 (N_7319,N_6897,N_6661);
xnor U7320 (N_7320,N_6019,N_6819);
or U7321 (N_7321,N_6623,N_6133);
xnor U7322 (N_7322,N_6664,N_6030);
nor U7323 (N_7323,N_6358,N_6433);
and U7324 (N_7324,N_6370,N_6812);
nand U7325 (N_7325,N_6943,N_6289);
xnor U7326 (N_7326,N_6887,N_6434);
nand U7327 (N_7327,N_6985,N_6319);
or U7328 (N_7328,N_6266,N_6959);
nand U7329 (N_7329,N_6792,N_6762);
and U7330 (N_7330,N_6653,N_6042);
nand U7331 (N_7331,N_6861,N_6252);
nor U7332 (N_7332,N_6851,N_6297);
or U7333 (N_7333,N_6324,N_6594);
nand U7334 (N_7334,N_6647,N_6803);
and U7335 (N_7335,N_6142,N_6052);
and U7336 (N_7336,N_6105,N_6534);
xor U7337 (N_7337,N_6145,N_6110);
nand U7338 (N_7338,N_6458,N_6998);
xnor U7339 (N_7339,N_6064,N_6018);
nand U7340 (N_7340,N_6034,N_6977);
and U7341 (N_7341,N_6915,N_6608);
and U7342 (N_7342,N_6056,N_6607);
nand U7343 (N_7343,N_6539,N_6391);
nor U7344 (N_7344,N_6696,N_6965);
nand U7345 (N_7345,N_6208,N_6621);
nor U7346 (N_7346,N_6442,N_6966);
and U7347 (N_7347,N_6739,N_6114);
or U7348 (N_7348,N_6728,N_6585);
nand U7349 (N_7349,N_6667,N_6113);
or U7350 (N_7350,N_6575,N_6580);
nand U7351 (N_7351,N_6176,N_6250);
xnor U7352 (N_7352,N_6761,N_6584);
nor U7353 (N_7353,N_6652,N_6115);
nand U7354 (N_7354,N_6360,N_6320);
xor U7355 (N_7355,N_6579,N_6519);
or U7356 (N_7356,N_6014,N_6317);
nand U7357 (N_7357,N_6895,N_6329);
and U7358 (N_7358,N_6660,N_6051);
nand U7359 (N_7359,N_6905,N_6476);
xnor U7360 (N_7360,N_6159,N_6204);
nand U7361 (N_7361,N_6267,N_6771);
and U7362 (N_7362,N_6693,N_6276);
nand U7363 (N_7363,N_6533,N_6066);
or U7364 (N_7364,N_6296,N_6921);
xor U7365 (N_7365,N_6565,N_6384);
and U7366 (N_7366,N_6491,N_6327);
or U7367 (N_7367,N_6169,N_6281);
xnor U7368 (N_7368,N_6464,N_6405);
and U7369 (N_7369,N_6777,N_6219);
xor U7370 (N_7370,N_6230,N_6641);
or U7371 (N_7371,N_6074,N_6850);
nand U7372 (N_7372,N_6516,N_6596);
nand U7373 (N_7373,N_6611,N_6574);
xnor U7374 (N_7374,N_6140,N_6988);
or U7375 (N_7375,N_6924,N_6466);
nand U7376 (N_7376,N_6083,N_6499);
and U7377 (N_7377,N_6531,N_6328);
and U7378 (N_7378,N_6446,N_6496);
or U7379 (N_7379,N_6707,N_6708);
nor U7380 (N_7380,N_6568,N_6235);
xnor U7381 (N_7381,N_6365,N_6163);
or U7382 (N_7382,N_6952,N_6823);
and U7383 (N_7383,N_6638,N_6868);
nand U7384 (N_7384,N_6870,N_6262);
nand U7385 (N_7385,N_6727,N_6486);
nor U7386 (N_7386,N_6831,N_6605);
xor U7387 (N_7387,N_6093,N_6278);
or U7388 (N_7388,N_6809,N_6845);
and U7389 (N_7389,N_6828,N_6512);
and U7390 (N_7390,N_6968,N_6509);
nand U7391 (N_7391,N_6754,N_6991);
xnor U7392 (N_7392,N_6429,N_6938);
nand U7393 (N_7393,N_6460,N_6076);
nand U7394 (N_7394,N_6352,N_6571);
and U7395 (N_7395,N_6598,N_6663);
nor U7396 (N_7396,N_6295,N_6811);
xor U7397 (N_7397,N_6910,N_6054);
nand U7398 (N_7398,N_6654,N_6316);
xnor U7399 (N_7399,N_6265,N_6618);
and U7400 (N_7400,N_6524,N_6603);
nor U7401 (N_7401,N_6749,N_6287);
or U7402 (N_7402,N_6541,N_6151);
xnor U7403 (N_7403,N_6143,N_6144);
nand U7404 (N_7404,N_6570,N_6756);
nor U7405 (N_7405,N_6302,N_6430);
or U7406 (N_7406,N_6492,N_6818);
nand U7407 (N_7407,N_6214,N_6017);
nand U7408 (N_7408,N_6583,N_6715);
and U7409 (N_7409,N_6305,N_6221);
nor U7410 (N_7410,N_6369,N_6737);
xnor U7411 (N_7411,N_6981,N_6960);
xnor U7412 (N_7412,N_6102,N_6672);
nor U7413 (N_7413,N_6732,N_6168);
nor U7414 (N_7414,N_6147,N_6755);
xor U7415 (N_7415,N_6772,N_6398);
nand U7416 (N_7416,N_6502,N_6407);
nor U7417 (N_7417,N_6226,N_6073);
nand U7418 (N_7418,N_6995,N_6167);
nor U7419 (N_7419,N_6560,N_6345);
nand U7420 (N_7420,N_6134,N_6045);
and U7421 (N_7421,N_6397,N_6865);
or U7422 (N_7422,N_6682,N_6858);
or U7423 (N_7423,N_6844,N_6258);
xor U7424 (N_7424,N_6372,N_6768);
or U7425 (N_7425,N_6878,N_6945);
nor U7426 (N_7426,N_6778,N_6919);
xor U7427 (N_7427,N_6684,N_6782);
nand U7428 (N_7428,N_6495,N_6510);
xor U7429 (N_7429,N_6891,N_6445);
xnor U7430 (N_7430,N_6122,N_6314);
nand U7431 (N_7431,N_6649,N_6385);
or U7432 (N_7432,N_6459,N_6216);
or U7433 (N_7433,N_6227,N_6498);
nand U7434 (N_7434,N_6440,N_6918);
and U7435 (N_7435,N_6347,N_6232);
nor U7436 (N_7436,N_6659,N_6679);
and U7437 (N_7437,N_6309,N_6817);
and U7438 (N_7438,N_6690,N_6884);
and U7439 (N_7439,N_6617,N_6548);
xor U7440 (N_7440,N_6655,N_6090);
or U7441 (N_7441,N_6098,N_6880);
or U7442 (N_7442,N_6839,N_6356);
nor U7443 (N_7443,N_6038,N_6949);
nor U7444 (N_7444,N_6409,N_6687);
nand U7445 (N_7445,N_6298,N_6181);
xor U7446 (N_7446,N_6862,N_6101);
xnor U7447 (N_7447,N_6337,N_6930);
or U7448 (N_7448,N_6031,N_6422);
nor U7449 (N_7449,N_6313,N_6186);
nor U7450 (N_7450,N_6978,N_6438);
and U7451 (N_7451,N_6209,N_6463);
or U7452 (N_7452,N_6714,N_6864);
xor U7453 (N_7453,N_6260,N_6241);
and U7454 (N_7454,N_6094,N_6909);
nand U7455 (N_7455,N_6477,N_6361);
nor U7456 (N_7456,N_6505,N_6719);
nand U7457 (N_7457,N_6273,N_6872);
xor U7458 (N_7458,N_6259,N_6410);
or U7459 (N_7459,N_6478,N_6600);
nor U7460 (N_7460,N_6417,N_6395);
or U7461 (N_7461,N_6542,N_6536);
and U7462 (N_7462,N_6773,N_6300);
xor U7463 (N_7463,N_6009,N_6472);
and U7464 (N_7464,N_6613,N_6035);
or U7465 (N_7465,N_6377,N_6742);
nand U7466 (N_7466,N_6299,N_6171);
or U7467 (N_7467,N_6702,N_6315);
xor U7468 (N_7468,N_6334,N_6253);
nor U7469 (N_7469,N_6532,N_6401);
and U7470 (N_7470,N_6198,N_6024);
nor U7471 (N_7471,N_6348,N_6139);
and U7472 (N_7472,N_6381,N_6040);
and U7473 (N_7473,N_6194,N_6136);
nand U7474 (N_7474,N_6974,N_6127);
xor U7475 (N_7475,N_6116,N_6402);
and U7476 (N_7476,N_6160,N_6331);
or U7477 (N_7477,N_6249,N_6179);
or U7478 (N_7478,N_6883,N_6217);
nand U7479 (N_7479,N_6481,N_6015);
nand U7480 (N_7480,N_6590,N_6220);
nor U7481 (N_7481,N_6624,N_6824);
nand U7482 (N_7482,N_6743,N_6200);
or U7483 (N_7483,N_6304,N_6821);
and U7484 (N_7484,N_6735,N_6540);
nand U7485 (N_7485,N_6553,N_6508);
nor U7486 (N_7486,N_6688,N_6651);
or U7487 (N_7487,N_6406,N_6174);
xor U7488 (N_7488,N_6588,N_6692);
or U7489 (N_7489,N_6303,N_6092);
xor U7490 (N_7490,N_6522,N_6640);
xor U7491 (N_7491,N_6775,N_6084);
and U7492 (N_7492,N_6480,N_6091);
xnor U7493 (N_7493,N_6840,N_6322);
xor U7494 (N_7494,N_6685,N_6984);
xnor U7495 (N_7495,N_6511,N_6189);
and U7496 (N_7496,N_6906,N_6201);
nor U7497 (N_7497,N_6886,N_6487);
nand U7498 (N_7498,N_6581,N_6471);
nand U7499 (N_7499,N_6871,N_6292);
xnor U7500 (N_7500,N_6872,N_6409);
or U7501 (N_7501,N_6185,N_6293);
or U7502 (N_7502,N_6166,N_6362);
or U7503 (N_7503,N_6517,N_6398);
and U7504 (N_7504,N_6295,N_6985);
nor U7505 (N_7505,N_6825,N_6363);
or U7506 (N_7506,N_6201,N_6512);
nor U7507 (N_7507,N_6352,N_6834);
and U7508 (N_7508,N_6628,N_6691);
xnor U7509 (N_7509,N_6074,N_6118);
xnor U7510 (N_7510,N_6926,N_6717);
nand U7511 (N_7511,N_6479,N_6836);
xnor U7512 (N_7512,N_6642,N_6202);
or U7513 (N_7513,N_6183,N_6490);
xor U7514 (N_7514,N_6175,N_6003);
nand U7515 (N_7515,N_6139,N_6121);
and U7516 (N_7516,N_6324,N_6622);
or U7517 (N_7517,N_6759,N_6664);
or U7518 (N_7518,N_6904,N_6582);
and U7519 (N_7519,N_6289,N_6972);
and U7520 (N_7520,N_6135,N_6371);
xnor U7521 (N_7521,N_6155,N_6098);
and U7522 (N_7522,N_6059,N_6568);
or U7523 (N_7523,N_6931,N_6391);
nor U7524 (N_7524,N_6155,N_6183);
xnor U7525 (N_7525,N_6703,N_6934);
nor U7526 (N_7526,N_6306,N_6501);
or U7527 (N_7527,N_6524,N_6615);
nand U7528 (N_7528,N_6615,N_6185);
or U7529 (N_7529,N_6359,N_6386);
xnor U7530 (N_7530,N_6011,N_6846);
nor U7531 (N_7531,N_6533,N_6736);
or U7532 (N_7532,N_6295,N_6140);
nand U7533 (N_7533,N_6495,N_6898);
xor U7534 (N_7534,N_6422,N_6288);
and U7535 (N_7535,N_6156,N_6212);
xnor U7536 (N_7536,N_6779,N_6397);
nor U7537 (N_7537,N_6230,N_6967);
nand U7538 (N_7538,N_6134,N_6639);
or U7539 (N_7539,N_6711,N_6622);
nand U7540 (N_7540,N_6563,N_6293);
xnor U7541 (N_7541,N_6641,N_6664);
nor U7542 (N_7542,N_6208,N_6530);
or U7543 (N_7543,N_6191,N_6769);
or U7544 (N_7544,N_6988,N_6410);
nand U7545 (N_7545,N_6810,N_6438);
nand U7546 (N_7546,N_6850,N_6655);
and U7547 (N_7547,N_6183,N_6166);
or U7548 (N_7548,N_6295,N_6988);
nand U7549 (N_7549,N_6343,N_6082);
xor U7550 (N_7550,N_6704,N_6844);
or U7551 (N_7551,N_6839,N_6821);
nor U7552 (N_7552,N_6251,N_6042);
nor U7553 (N_7553,N_6880,N_6929);
nor U7554 (N_7554,N_6636,N_6071);
nand U7555 (N_7555,N_6405,N_6417);
nand U7556 (N_7556,N_6106,N_6728);
and U7557 (N_7557,N_6425,N_6820);
xnor U7558 (N_7558,N_6078,N_6758);
and U7559 (N_7559,N_6327,N_6853);
or U7560 (N_7560,N_6976,N_6855);
nor U7561 (N_7561,N_6948,N_6211);
nand U7562 (N_7562,N_6146,N_6583);
and U7563 (N_7563,N_6166,N_6909);
nor U7564 (N_7564,N_6815,N_6793);
xnor U7565 (N_7565,N_6646,N_6141);
xnor U7566 (N_7566,N_6450,N_6946);
and U7567 (N_7567,N_6821,N_6604);
nand U7568 (N_7568,N_6627,N_6996);
nand U7569 (N_7569,N_6399,N_6148);
or U7570 (N_7570,N_6517,N_6974);
nor U7571 (N_7571,N_6929,N_6849);
nand U7572 (N_7572,N_6962,N_6551);
nor U7573 (N_7573,N_6126,N_6784);
and U7574 (N_7574,N_6990,N_6321);
nor U7575 (N_7575,N_6936,N_6424);
and U7576 (N_7576,N_6114,N_6449);
and U7577 (N_7577,N_6792,N_6262);
nand U7578 (N_7578,N_6493,N_6855);
nor U7579 (N_7579,N_6117,N_6894);
nor U7580 (N_7580,N_6377,N_6370);
and U7581 (N_7581,N_6149,N_6819);
xor U7582 (N_7582,N_6175,N_6338);
and U7583 (N_7583,N_6567,N_6229);
nor U7584 (N_7584,N_6571,N_6790);
or U7585 (N_7585,N_6840,N_6138);
or U7586 (N_7586,N_6586,N_6489);
or U7587 (N_7587,N_6172,N_6472);
nor U7588 (N_7588,N_6298,N_6091);
nand U7589 (N_7589,N_6621,N_6226);
and U7590 (N_7590,N_6601,N_6166);
and U7591 (N_7591,N_6927,N_6626);
or U7592 (N_7592,N_6159,N_6735);
and U7593 (N_7593,N_6818,N_6049);
nand U7594 (N_7594,N_6300,N_6438);
xor U7595 (N_7595,N_6567,N_6265);
xnor U7596 (N_7596,N_6576,N_6563);
xnor U7597 (N_7597,N_6576,N_6210);
and U7598 (N_7598,N_6490,N_6124);
nand U7599 (N_7599,N_6549,N_6743);
xnor U7600 (N_7600,N_6215,N_6798);
nor U7601 (N_7601,N_6518,N_6316);
nand U7602 (N_7602,N_6322,N_6430);
xnor U7603 (N_7603,N_6000,N_6830);
or U7604 (N_7604,N_6261,N_6471);
and U7605 (N_7605,N_6319,N_6986);
xnor U7606 (N_7606,N_6769,N_6797);
nand U7607 (N_7607,N_6032,N_6885);
and U7608 (N_7608,N_6281,N_6402);
or U7609 (N_7609,N_6490,N_6888);
or U7610 (N_7610,N_6866,N_6049);
xnor U7611 (N_7611,N_6442,N_6302);
and U7612 (N_7612,N_6648,N_6143);
nor U7613 (N_7613,N_6797,N_6858);
and U7614 (N_7614,N_6889,N_6323);
nand U7615 (N_7615,N_6460,N_6391);
nand U7616 (N_7616,N_6689,N_6772);
nor U7617 (N_7617,N_6300,N_6891);
nand U7618 (N_7618,N_6600,N_6472);
nor U7619 (N_7619,N_6316,N_6090);
nor U7620 (N_7620,N_6870,N_6434);
nor U7621 (N_7621,N_6945,N_6026);
nor U7622 (N_7622,N_6685,N_6484);
nand U7623 (N_7623,N_6643,N_6502);
nand U7624 (N_7624,N_6182,N_6069);
xnor U7625 (N_7625,N_6142,N_6265);
xnor U7626 (N_7626,N_6333,N_6116);
nand U7627 (N_7627,N_6465,N_6196);
nor U7628 (N_7628,N_6719,N_6091);
and U7629 (N_7629,N_6326,N_6944);
and U7630 (N_7630,N_6947,N_6614);
xnor U7631 (N_7631,N_6210,N_6198);
nor U7632 (N_7632,N_6591,N_6339);
xor U7633 (N_7633,N_6274,N_6187);
or U7634 (N_7634,N_6994,N_6453);
or U7635 (N_7635,N_6584,N_6160);
nand U7636 (N_7636,N_6832,N_6521);
and U7637 (N_7637,N_6746,N_6697);
or U7638 (N_7638,N_6445,N_6456);
and U7639 (N_7639,N_6386,N_6571);
or U7640 (N_7640,N_6905,N_6072);
and U7641 (N_7641,N_6043,N_6524);
xnor U7642 (N_7642,N_6114,N_6531);
nand U7643 (N_7643,N_6813,N_6425);
xor U7644 (N_7644,N_6934,N_6349);
and U7645 (N_7645,N_6744,N_6129);
nand U7646 (N_7646,N_6767,N_6244);
nand U7647 (N_7647,N_6832,N_6312);
nand U7648 (N_7648,N_6246,N_6690);
and U7649 (N_7649,N_6996,N_6955);
or U7650 (N_7650,N_6529,N_6272);
nor U7651 (N_7651,N_6329,N_6584);
and U7652 (N_7652,N_6380,N_6590);
xnor U7653 (N_7653,N_6798,N_6163);
nor U7654 (N_7654,N_6393,N_6530);
nor U7655 (N_7655,N_6224,N_6127);
or U7656 (N_7656,N_6077,N_6672);
nand U7657 (N_7657,N_6749,N_6746);
nor U7658 (N_7658,N_6179,N_6069);
nand U7659 (N_7659,N_6780,N_6174);
and U7660 (N_7660,N_6438,N_6642);
or U7661 (N_7661,N_6737,N_6185);
xnor U7662 (N_7662,N_6070,N_6778);
nor U7663 (N_7663,N_6575,N_6870);
or U7664 (N_7664,N_6028,N_6013);
and U7665 (N_7665,N_6107,N_6122);
xnor U7666 (N_7666,N_6319,N_6563);
nand U7667 (N_7667,N_6592,N_6556);
nand U7668 (N_7668,N_6641,N_6973);
nor U7669 (N_7669,N_6091,N_6132);
nand U7670 (N_7670,N_6196,N_6993);
and U7671 (N_7671,N_6660,N_6219);
and U7672 (N_7672,N_6693,N_6293);
and U7673 (N_7673,N_6935,N_6254);
and U7674 (N_7674,N_6884,N_6357);
and U7675 (N_7675,N_6194,N_6295);
and U7676 (N_7676,N_6085,N_6271);
and U7677 (N_7677,N_6781,N_6323);
and U7678 (N_7678,N_6236,N_6312);
nand U7679 (N_7679,N_6377,N_6115);
nor U7680 (N_7680,N_6711,N_6924);
nor U7681 (N_7681,N_6525,N_6855);
and U7682 (N_7682,N_6179,N_6578);
xor U7683 (N_7683,N_6398,N_6899);
xnor U7684 (N_7684,N_6091,N_6628);
nand U7685 (N_7685,N_6140,N_6630);
or U7686 (N_7686,N_6975,N_6000);
and U7687 (N_7687,N_6303,N_6977);
nand U7688 (N_7688,N_6543,N_6950);
and U7689 (N_7689,N_6268,N_6943);
xor U7690 (N_7690,N_6286,N_6933);
and U7691 (N_7691,N_6401,N_6607);
and U7692 (N_7692,N_6979,N_6779);
or U7693 (N_7693,N_6792,N_6297);
nor U7694 (N_7694,N_6565,N_6385);
nor U7695 (N_7695,N_6125,N_6256);
or U7696 (N_7696,N_6081,N_6855);
xnor U7697 (N_7697,N_6460,N_6323);
nand U7698 (N_7698,N_6270,N_6046);
nand U7699 (N_7699,N_6144,N_6104);
or U7700 (N_7700,N_6822,N_6930);
nor U7701 (N_7701,N_6818,N_6674);
or U7702 (N_7702,N_6508,N_6319);
nand U7703 (N_7703,N_6706,N_6584);
nand U7704 (N_7704,N_6335,N_6799);
nor U7705 (N_7705,N_6413,N_6722);
nand U7706 (N_7706,N_6912,N_6605);
xor U7707 (N_7707,N_6926,N_6344);
nor U7708 (N_7708,N_6333,N_6332);
nand U7709 (N_7709,N_6335,N_6869);
xnor U7710 (N_7710,N_6977,N_6365);
nand U7711 (N_7711,N_6229,N_6711);
or U7712 (N_7712,N_6893,N_6620);
nor U7713 (N_7713,N_6905,N_6689);
nor U7714 (N_7714,N_6204,N_6683);
and U7715 (N_7715,N_6725,N_6956);
nand U7716 (N_7716,N_6692,N_6124);
or U7717 (N_7717,N_6522,N_6398);
xor U7718 (N_7718,N_6891,N_6163);
and U7719 (N_7719,N_6409,N_6675);
nor U7720 (N_7720,N_6202,N_6893);
xnor U7721 (N_7721,N_6027,N_6019);
and U7722 (N_7722,N_6948,N_6419);
and U7723 (N_7723,N_6051,N_6174);
nor U7724 (N_7724,N_6428,N_6914);
nor U7725 (N_7725,N_6237,N_6096);
xor U7726 (N_7726,N_6570,N_6601);
nor U7727 (N_7727,N_6957,N_6092);
nor U7728 (N_7728,N_6238,N_6521);
nand U7729 (N_7729,N_6977,N_6491);
or U7730 (N_7730,N_6938,N_6758);
xor U7731 (N_7731,N_6004,N_6996);
nand U7732 (N_7732,N_6875,N_6340);
or U7733 (N_7733,N_6658,N_6557);
nor U7734 (N_7734,N_6861,N_6352);
nand U7735 (N_7735,N_6914,N_6383);
or U7736 (N_7736,N_6984,N_6210);
or U7737 (N_7737,N_6865,N_6076);
and U7738 (N_7738,N_6109,N_6639);
or U7739 (N_7739,N_6445,N_6227);
or U7740 (N_7740,N_6198,N_6974);
and U7741 (N_7741,N_6511,N_6011);
or U7742 (N_7742,N_6937,N_6974);
nor U7743 (N_7743,N_6670,N_6044);
and U7744 (N_7744,N_6484,N_6822);
xnor U7745 (N_7745,N_6481,N_6662);
xor U7746 (N_7746,N_6337,N_6987);
or U7747 (N_7747,N_6818,N_6411);
nand U7748 (N_7748,N_6069,N_6888);
or U7749 (N_7749,N_6789,N_6402);
or U7750 (N_7750,N_6938,N_6024);
or U7751 (N_7751,N_6629,N_6239);
nor U7752 (N_7752,N_6354,N_6280);
and U7753 (N_7753,N_6968,N_6255);
xor U7754 (N_7754,N_6504,N_6054);
or U7755 (N_7755,N_6443,N_6932);
or U7756 (N_7756,N_6785,N_6721);
nand U7757 (N_7757,N_6159,N_6059);
nor U7758 (N_7758,N_6053,N_6341);
nor U7759 (N_7759,N_6625,N_6848);
nand U7760 (N_7760,N_6302,N_6433);
xor U7761 (N_7761,N_6606,N_6589);
or U7762 (N_7762,N_6179,N_6920);
xnor U7763 (N_7763,N_6715,N_6766);
and U7764 (N_7764,N_6504,N_6991);
nor U7765 (N_7765,N_6921,N_6334);
and U7766 (N_7766,N_6030,N_6921);
xor U7767 (N_7767,N_6234,N_6929);
xnor U7768 (N_7768,N_6839,N_6664);
nand U7769 (N_7769,N_6593,N_6574);
xor U7770 (N_7770,N_6323,N_6164);
or U7771 (N_7771,N_6725,N_6689);
xor U7772 (N_7772,N_6426,N_6076);
or U7773 (N_7773,N_6966,N_6159);
or U7774 (N_7774,N_6452,N_6256);
nor U7775 (N_7775,N_6318,N_6026);
nand U7776 (N_7776,N_6920,N_6900);
xor U7777 (N_7777,N_6685,N_6074);
nand U7778 (N_7778,N_6926,N_6783);
nor U7779 (N_7779,N_6843,N_6771);
xnor U7780 (N_7780,N_6106,N_6249);
xnor U7781 (N_7781,N_6846,N_6183);
or U7782 (N_7782,N_6174,N_6338);
nand U7783 (N_7783,N_6373,N_6012);
nand U7784 (N_7784,N_6688,N_6303);
nor U7785 (N_7785,N_6432,N_6793);
nor U7786 (N_7786,N_6477,N_6113);
nor U7787 (N_7787,N_6722,N_6215);
and U7788 (N_7788,N_6682,N_6281);
nand U7789 (N_7789,N_6008,N_6986);
nand U7790 (N_7790,N_6770,N_6459);
and U7791 (N_7791,N_6845,N_6790);
nand U7792 (N_7792,N_6876,N_6603);
xor U7793 (N_7793,N_6513,N_6316);
or U7794 (N_7794,N_6552,N_6218);
nand U7795 (N_7795,N_6993,N_6926);
nand U7796 (N_7796,N_6602,N_6220);
and U7797 (N_7797,N_6620,N_6451);
nand U7798 (N_7798,N_6532,N_6537);
and U7799 (N_7799,N_6398,N_6876);
nor U7800 (N_7800,N_6210,N_6888);
xnor U7801 (N_7801,N_6080,N_6188);
xor U7802 (N_7802,N_6103,N_6403);
nor U7803 (N_7803,N_6583,N_6745);
xnor U7804 (N_7804,N_6707,N_6212);
and U7805 (N_7805,N_6252,N_6027);
or U7806 (N_7806,N_6281,N_6233);
and U7807 (N_7807,N_6416,N_6214);
or U7808 (N_7808,N_6704,N_6957);
xor U7809 (N_7809,N_6481,N_6781);
or U7810 (N_7810,N_6496,N_6287);
nor U7811 (N_7811,N_6616,N_6194);
xor U7812 (N_7812,N_6886,N_6052);
nand U7813 (N_7813,N_6048,N_6609);
or U7814 (N_7814,N_6219,N_6283);
nor U7815 (N_7815,N_6065,N_6334);
and U7816 (N_7816,N_6404,N_6536);
or U7817 (N_7817,N_6418,N_6584);
xor U7818 (N_7818,N_6621,N_6882);
or U7819 (N_7819,N_6824,N_6108);
nand U7820 (N_7820,N_6420,N_6212);
xnor U7821 (N_7821,N_6122,N_6300);
or U7822 (N_7822,N_6494,N_6069);
xnor U7823 (N_7823,N_6647,N_6861);
nand U7824 (N_7824,N_6932,N_6916);
xor U7825 (N_7825,N_6495,N_6446);
nand U7826 (N_7826,N_6196,N_6814);
nor U7827 (N_7827,N_6145,N_6118);
nand U7828 (N_7828,N_6606,N_6511);
nor U7829 (N_7829,N_6560,N_6374);
and U7830 (N_7830,N_6323,N_6120);
or U7831 (N_7831,N_6711,N_6510);
xnor U7832 (N_7832,N_6376,N_6250);
or U7833 (N_7833,N_6251,N_6641);
nand U7834 (N_7834,N_6888,N_6326);
or U7835 (N_7835,N_6423,N_6289);
nor U7836 (N_7836,N_6211,N_6535);
nor U7837 (N_7837,N_6861,N_6447);
or U7838 (N_7838,N_6679,N_6286);
xor U7839 (N_7839,N_6541,N_6681);
and U7840 (N_7840,N_6726,N_6677);
and U7841 (N_7841,N_6761,N_6336);
and U7842 (N_7842,N_6661,N_6690);
and U7843 (N_7843,N_6791,N_6367);
or U7844 (N_7844,N_6896,N_6895);
nand U7845 (N_7845,N_6231,N_6711);
and U7846 (N_7846,N_6017,N_6794);
and U7847 (N_7847,N_6368,N_6396);
nor U7848 (N_7848,N_6143,N_6076);
or U7849 (N_7849,N_6615,N_6331);
nand U7850 (N_7850,N_6659,N_6578);
xnor U7851 (N_7851,N_6739,N_6448);
xnor U7852 (N_7852,N_6159,N_6675);
nor U7853 (N_7853,N_6846,N_6919);
nand U7854 (N_7854,N_6166,N_6122);
nor U7855 (N_7855,N_6449,N_6530);
xor U7856 (N_7856,N_6664,N_6120);
nor U7857 (N_7857,N_6708,N_6018);
and U7858 (N_7858,N_6679,N_6360);
or U7859 (N_7859,N_6198,N_6098);
and U7860 (N_7860,N_6311,N_6493);
nor U7861 (N_7861,N_6485,N_6039);
or U7862 (N_7862,N_6154,N_6706);
nor U7863 (N_7863,N_6126,N_6814);
xor U7864 (N_7864,N_6893,N_6302);
and U7865 (N_7865,N_6482,N_6976);
or U7866 (N_7866,N_6241,N_6812);
xor U7867 (N_7867,N_6176,N_6841);
xor U7868 (N_7868,N_6394,N_6389);
or U7869 (N_7869,N_6861,N_6899);
xnor U7870 (N_7870,N_6805,N_6537);
nand U7871 (N_7871,N_6512,N_6806);
nor U7872 (N_7872,N_6897,N_6018);
and U7873 (N_7873,N_6419,N_6293);
or U7874 (N_7874,N_6203,N_6858);
nor U7875 (N_7875,N_6288,N_6820);
and U7876 (N_7876,N_6215,N_6547);
nand U7877 (N_7877,N_6719,N_6066);
xor U7878 (N_7878,N_6341,N_6493);
or U7879 (N_7879,N_6214,N_6413);
xnor U7880 (N_7880,N_6926,N_6434);
or U7881 (N_7881,N_6640,N_6770);
nand U7882 (N_7882,N_6178,N_6708);
and U7883 (N_7883,N_6381,N_6285);
xor U7884 (N_7884,N_6776,N_6897);
nand U7885 (N_7885,N_6302,N_6351);
nand U7886 (N_7886,N_6426,N_6122);
and U7887 (N_7887,N_6835,N_6337);
or U7888 (N_7888,N_6769,N_6530);
nand U7889 (N_7889,N_6260,N_6015);
nor U7890 (N_7890,N_6782,N_6941);
nor U7891 (N_7891,N_6808,N_6702);
nor U7892 (N_7892,N_6318,N_6964);
and U7893 (N_7893,N_6035,N_6741);
xnor U7894 (N_7894,N_6148,N_6942);
nand U7895 (N_7895,N_6422,N_6964);
and U7896 (N_7896,N_6922,N_6211);
nor U7897 (N_7897,N_6233,N_6759);
and U7898 (N_7898,N_6500,N_6750);
nand U7899 (N_7899,N_6948,N_6034);
xor U7900 (N_7900,N_6455,N_6513);
and U7901 (N_7901,N_6550,N_6913);
nand U7902 (N_7902,N_6901,N_6933);
or U7903 (N_7903,N_6919,N_6850);
nor U7904 (N_7904,N_6885,N_6076);
nor U7905 (N_7905,N_6414,N_6495);
nand U7906 (N_7906,N_6823,N_6732);
xor U7907 (N_7907,N_6181,N_6828);
nor U7908 (N_7908,N_6103,N_6320);
or U7909 (N_7909,N_6500,N_6026);
and U7910 (N_7910,N_6528,N_6690);
xor U7911 (N_7911,N_6509,N_6737);
and U7912 (N_7912,N_6469,N_6720);
nand U7913 (N_7913,N_6357,N_6553);
or U7914 (N_7914,N_6032,N_6302);
nand U7915 (N_7915,N_6917,N_6292);
nor U7916 (N_7916,N_6817,N_6218);
or U7917 (N_7917,N_6547,N_6233);
nand U7918 (N_7918,N_6482,N_6215);
nor U7919 (N_7919,N_6512,N_6697);
nand U7920 (N_7920,N_6408,N_6827);
nand U7921 (N_7921,N_6929,N_6151);
and U7922 (N_7922,N_6005,N_6266);
xnor U7923 (N_7923,N_6238,N_6122);
or U7924 (N_7924,N_6247,N_6609);
or U7925 (N_7925,N_6965,N_6471);
or U7926 (N_7926,N_6054,N_6897);
and U7927 (N_7927,N_6724,N_6535);
and U7928 (N_7928,N_6651,N_6609);
nand U7929 (N_7929,N_6554,N_6898);
nor U7930 (N_7930,N_6391,N_6156);
or U7931 (N_7931,N_6766,N_6948);
xor U7932 (N_7932,N_6874,N_6816);
xnor U7933 (N_7933,N_6683,N_6468);
xnor U7934 (N_7934,N_6597,N_6377);
and U7935 (N_7935,N_6143,N_6742);
nand U7936 (N_7936,N_6147,N_6253);
and U7937 (N_7937,N_6626,N_6803);
or U7938 (N_7938,N_6142,N_6388);
xor U7939 (N_7939,N_6871,N_6971);
and U7940 (N_7940,N_6236,N_6525);
nor U7941 (N_7941,N_6649,N_6568);
nand U7942 (N_7942,N_6542,N_6217);
nor U7943 (N_7943,N_6652,N_6926);
and U7944 (N_7944,N_6868,N_6946);
and U7945 (N_7945,N_6833,N_6663);
nand U7946 (N_7946,N_6473,N_6950);
and U7947 (N_7947,N_6574,N_6244);
or U7948 (N_7948,N_6848,N_6204);
or U7949 (N_7949,N_6934,N_6055);
xnor U7950 (N_7950,N_6354,N_6752);
and U7951 (N_7951,N_6823,N_6529);
and U7952 (N_7952,N_6507,N_6326);
or U7953 (N_7953,N_6696,N_6998);
and U7954 (N_7954,N_6994,N_6118);
nand U7955 (N_7955,N_6715,N_6759);
or U7956 (N_7956,N_6352,N_6074);
nand U7957 (N_7957,N_6354,N_6231);
nand U7958 (N_7958,N_6573,N_6728);
xnor U7959 (N_7959,N_6121,N_6407);
nor U7960 (N_7960,N_6247,N_6648);
nor U7961 (N_7961,N_6939,N_6181);
and U7962 (N_7962,N_6825,N_6761);
nor U7963 (N_7963,N_6966,N_6533);
or U7964 (N_7964,N_6263,N_6057);
xnor U7965 (N_7965,N_6799,N_6049);
xnor U7966 (N_7966,N_6035,N_6763);
nor U7967 (N_7967,N_6728,N_6470);
and U7968 (N_7968,N_6648,N_6925);
xnor U7969 (N_7969,N_6235,N_6089);
or U7970 (N_7970,N_6110,N_6027);
nor U7971 (N_7971,N_6899,N_6791);
xnor U7972 (N_7972,N_6400,N_6662);
and U7973 (N_7973,N_6107,N_6479);
nand U7974 (N_7974,N_6147,N_6347);
nand U7975 (N_7975,N_6946,N_6285);
nand U7976 (N_7976,N_6097,N_6413);
or U7977 (N_7977,N_6750,N_6631);
or U7978 (N_7978,N_6634,N_6876);
nor U7979 (N_7979,N_6661,N_6792);
xor U7980 (N_7980,N_6633,N_6647);
and U7981 (N_7981,N_6668,N_6577);
nor U7982 (N_7982,N_6224,N_6804);
and U7983 (N_7983,N_6424,N_6300);
xnor U7984 (N_7984,N_6605,N_6954);
and U7985 (N_7985,N_6983,N_6202);
or U7986 (N_7986,N_6284,N_6206);
and U7987 (N_7987,N_6813,N_6851);
and U7988 (N_7988,N_6897,N_6804);
nand U7989 (N_7989,N_6161,N_6549);
and U7990 (N_7990,N_6150,N_6983);
or U7991 (N_7991,N_6170,N_6159);
nor U7992 (N_7992,N_6561,N_6648);
or U7993 (N_7993,N_6354,N_6162);
nor U7994 (N_7994,N_6847,N_6334);
nor U7995 (N_7995,N_6547,N_6669);
xnor U7996 (N_7996,N_6895,N_6044);
or U7997 (N_7997,N_6768,N_6055);
or U7998 (N_7998,N_6705,N_6906);
nor U7999 (N_7999,N_6895,N_6477);
and U8000 (N_8000,N_7969,N_7617);
nand U8001 (N_8001,N_7217,N_7001);
xor U8002 (N_8002,N_7642,N_7694);
and U8003 (N_8003,N_7065,N_7026);
nand U8004 (N_8004,N_7941,N_7376);
or U8005 (N_8005,N_7700,N_7182);
or U8006 (N_8006,N_7504,N_7111);
nand U8007 (N_8007,N_7965,N_7168);
or U8008 (N_8008,N_7777,N_7519);
or U8009 (N_8009,N_7103,N_7881);
xnor U8010 (N_8010,N_7463,N_7833);
nor U8011 (N_8011,N_7944,N_7566);
nor U8012 (N_8012,N_7922,N_7392);
xnor U8013 (N_8013,N_7767,N_7604);
nor U8014 (N_8014,N_7279,N_7013);
and U8015 (N_8015,N_7015,N_7095);
and U8016 (N_8016,N_7336,N_7876);
or U8017 (N_8017,N_7543,N_7363);
nand U8018 (N_8018,N_7780,N_7695);
nand U8019 (N_8019,N_7704,N_7819);
nand U8020 (N_8020,N_7326,N_7439);
xor U8021 (N_8021,N_7536,N_7926);
or U8022 (N_8022,N_7594,N_7334);
xor U8023 (N_8023,N_7154,N_7874);
nor U8024 (N_8024,N_7238,N_7775);
and U8025 (N_8025,N_7714,N_7323);
xnor U8026 (N_8026,N_7955,N_7356);
xor U8027 (N_8027,N_7362,N_7974);
or U8028 (N_8028,N_7079,N_7825);
xor U8029 (N_8029,N_7468,N_7585);
or U8030 (N_8030,N_7913,N_7502);
nand U8031 (N_8031,N_7533,N_7273);
or U8032 (N_8032,N_7124,N_7216);
and U8033 (N_8033,N_7265,N_7126);
nand U8034 (N_8034,N_7612,N_7441);
and U8035 (N_8035,N_7956,N_7868);
nand U8036 (N_8036,N_7781,N_7343);
nand U8037 (N_8037,N_7359,N_7198);
or U8038 (N_8038,N_7559,N_7471);
nor U8039 (N_8039,N_7107,N_7232);
and U8040 (N_8040,N_7480,N_7218);
or U8041 (N_8041,N_7078,N_7607);
and U8042 (N_8042,N_7771,N_7651);
xor U8043 (N_8043,N_7951,N_7779);
nand U8044 (N_8044,N_7658,N_7177);
xnor U8045 (N_8045,N_7138,N_7341);
and U8046 (N_8046,N_7640,N_7598);
xor U8047 (N_8047,N_7398,N_7059);
and U8048 (N_8048,N_7142,N_7481);
and U8049 (N_8049,N_7277,N_7121);
or U8050 (N_8050,N_7828,N_7464);
and U8051 (N_8051,N_7952,N_7222);
nand U8052 (N_8052,N_7417,N_7758);
xor U8053 (N_8053,N_7386,N_7385);
and U8054 (N_8054,N_7603,N_7950);
xor U8055 (N_8055,N_7094,N_7170);
nor U8056 (N_8056,N_7520,N_7432);
or U8057 (N_8057,N_7048,N_7637);
nor U8058 (N_8058,N_7497,N_7804);
and U8059 (N_8059,N_7482,N_7584);
nor U8060 (N_8060,N_7228,N_7477);
xor U8061 (N_8061,N_7389,N_7146);
and U8062 (N_8062,N_7155,N_7797);
nor U8063 (N_8063,N_7555,N_7761);
xnor U8064 (N_8064,N_7050,N_7940);
xor U8065 (N_8065,N_7233,N_7012);
xnor U8066 (N_8066,N_7425,N_7418);
nor U8067 (N_8067,N_7041,N_7304);
nand U8068 (N_8068,N_7203,N_7259);
and U8069 (N_8069,N_7794,N_7800);
xor U8070 (N_8070,N_7656,N_7062);
xnor U8071 (N_8071,N_7366,N_7237);
and U8072 (N_8072,N_7629,N_7615);
or U8073 (N_8073,N_7229,N_7889);
or U8074 (N_8074,N_7856,N_7479);
nand U8075 (N_8075,N_7759,N_7474);
and U8076 (N_8076,N_7899,N_7581);
or U8077 (N_8077,N_7085,N_7354);
nand U8078 (N_8078,N_7410,N_7141);
xor U8079 (N_8079,N_7632,N_7673);
and U8080 (N_8080,N_7263,N_7434);
nand U8081 (N_8081,N_7503,N_7647);
nand U8082 (N_8082,N_7236,N_7115);
xnor U8083 (N_8083,N_7671,N_7374);
nand U8084 (N_8084,N_7145,N_7312);
nor U8085 (N_8085,N_7290,N_7002);
xor U8086 (N_8086,N_7949,N_7678);
nand U8087 (N_8087,N_7301,N_7046);
and U8088 (N_8088,N_7143,N_7407);
nand U8089 (N_8089,N_7877,N_7871);
nor U8090 (N_8090,N_7136,N_7090);
nor U8091 (N_8091,N_7730,N_7753);
and U8092 (N_8092,N_7882,N_7246);
and U8093 (N_8093,N_7208,N_7674);
nand U8094 (N_8094,N_7980,N_7708);
or U8095 (N_8095,N_7370,N_7644);
nor U8096 (N_8096,N_7861,N_7494);
xor U8097 (N_8097,N_7883,N_7823);
xor U8098 (N_8098,N_7358,N_7500);
or U8099 (N_8099,N_7774,N_7827);
xnor U8100 (N_8100,N_7666,N_7844);
and U8101 (N_8101,N_7628,N_7812);
xnor U8102 (N_8102,N_7611,N_7660);
nand U8103 (N_8103,N_7082,N_7716);
nand U8104 (N_8104,N_7925,N_7687);
and U8105 (N_8105,N_7428,N_7419);
xnor U8106 (N_8106,N_7089,N_7932);
nor U8107 (N_8107,N_7315,N_7108);
nand U8108 (N_8108,N_7507,N_7788);
xnor U8109 (N_8109,N_7933,N_7515);
nand U8110 (N_8110,N_7183,N_7711);
nand U8111 (N_8111,N_7728,N_7506);
or U8112 (N_8112,N_7006,N_7158);
and U8113 (N_8113,N_7721,N_7175);
nor U8114 (N_8114,N_7302,N_7467);
and U8115 (N_8115,N_7226,N_7976);
nor U8116 (N_8116,N_7499,N_7454);
and U8117 (N_8117,N_7029,N_7060);
nor U8118 (N_8118,N_7484,N_7361);
xor U8119 (N_8119,N_7395,N_7030);
or U8120 (N_8120,N_7857,N_7406);
xor U8121 (N_8121,N_7377,N_7998);
nand U8122 (N_8122,N_7038,N_7578);
xnor U8123 (N_8123,N_7818,N_7099);
xnor U8124 (N_8124,N_7133,N_7490);
nor U8125 (N_8125,N_7928,N_7938);
or U8126 (N_8126,N_7817,N_7387);
and U8127 (N_8127,N_7491,N_7963);
nor U8128 (N_8128,N_7973,N_7076);
nand U8129 (N_8129,N_7970,N_7591);
nand U8130 (N_8130,N_7747,N_7193);
nor U8131 (N_8131,N_7764,N_7908);
nand U8132 (N_8132,N_7547,N_7548);
nand U8133 (N_8133,N_7967,N_7664);
nor U8134 (N_8134,N_7894,N_7074);
and U8135 (N_8135,N_7219,N_7285);
nand U8136 (N_8136,N_7296,N_7117);
or U8137 (N_8137,N_7227,N_7652);
xor U8138 (N_8138,N_7348,N_7453);
nor U8139 (N_8139,N_7532,N_7028);
nor U8140 (N_8140,N_7648,N_7033);
and U8141 (N_8141,N_7744,N_7100);
or U8142 (N_8142,N_7590,N_7424);
nor U8143 (N_8143,N_7902,N_7247);
or U8144 (N_8144,N_7318,N_7586);
xor U8145 (N_8145,N_7564,N_7081);
xor U8146 (N_8146,N_7668,N_7654);
and U8147 (N_8147,N_7895,N_7396);
xnor U8148 (N_8148,N_7054,N_7561);
xnor U8149 (N_8149,N_7959,N_7313);
or U8150 (N_8150,N_7866,N_7413);
nor U8151 (N_8151,N_7712,N_7862);
xnor U8152 (N_8152,N_7689,N_7286);
or U8153 (N_8153,N_7717,N_7443);
nor U8154 (N_8154,N_7526,N_7901);
and U8155 (N_8155,N_7845,N_7197);
nand U8156 (N_8156,N_7920,N_7863);
and U8157 (N_8157,N_7870,N_7679);
and U8158 (N_8158,N_7421,N_7171);
or U8159 (N_8159,N_7683,N_7806);
and U8160 (N_8160,N_7791,N_7268);
xnor U8161 (N_8161,N_7577,N_7667);
nand U8162 (N_8162,N_7609,N_7159);
and U8163 (N_8163,N_7641,N_7657);
nor U8164 (N_8164,N_7905,N_7676);
or U8165 (N_8165,N_7291,N_7743);
nor U8166 (N_8166,N_7442,N_7707);
or U8167 (N_8167,N_7537,N_7622);
and U8168 (N_8168,N_7776,N_7670);
xor U8169 (N_8169,N_7997,N_7045);
and U8170 (N_8170,N_7025,N_7073);
xnor U8171 (N_8171,N_7858,N_7663);
nor U8172 (N_8172,N_7992,N_7732);
nand U8173 (N_8173,N_7461,N_7596);
nor U8174 (N_8174,N_7587,N_7662);
nand U8175 (N_8175,N_7961,N_7098);
and U8176 (N_8176,N_7253,N_7623);
nand U8177 (N_8177,N_7986,N_7049);
xor U8178 (N_8178,N_7665,N_7202);
nor U8179 (N_8179,N_7729,N_7795);
nand U8180 (N_8180,N_7738,N_7692);
or U8181 (N_8181,N_7207,N_7703);
and U8182 (N_8182,N_7355,N_7210);
nor U8183 (N_8183,N_7064,N_7262);
or U8184 (N_8184,N_7782,N_7364);
nand U8185 (N_8185,N_7378,N_7842);
nand U8186 (N_8186,N_7245,N_7600);
nand U8187 (N_8187,N_7869,N_7373);
nor U8188 (N_8188,N_7958,N_7523);
xnor U8189 (N_8189,N_7996,N_7524);
and U8190 (N_8190,N_7750,N_7096);
and U8191 (N_8191,N_7725,N_7251);
nand U8192 (N_8192,N_7860,N_7031);
nand U8193 (N_8193,N_7787,N_7472);
xor U8194 (N_8194,N_7852,N_7016);
and U8195 (N_8195,N_7904,N_7139);
nand U8196 (N_8196,N_7039,N_7538);
and U8197 (N_8197,N_7166,N_7552);
and U8198 (N_8198,N_7324,N_7911);
nor U8199 (N_8199,N_7003,N_7971);
xnor U8200 (N_8200,N_7267,N_7435);
and U8201 (N_8201,N_7269,N_7789);
nor U8202 (N_8202,N_7426,N_7128);
and U8203 (N_8203,N_7231,N_7365);
and U8204 (N_8204,N_7448,N_7786);
and U8205 (N_8205,N_7769,N_7368);
xnor U8206 (N_8206,N_7184,N_7037);
nand U8207 (N_8207,N_7826,N_7962);
xnor U8208 (N_8208,N_7731,N_7397);
nor U8209 (N_8209,N_7568,N_7748);
and U8210 (N_8210,N_7019,N_7772);
and U8211 (N_8211,N_7293,N_7760);
nor U8212 (N_8212,N_7040,N_7943);
nand U8213 (N_8213,N_7196,N_7129);
xnor U8214 (N_8214,N_7488,N_7636);
nor U8215 (N_8215,N_7405,N_7101);
xor U8216 (N_8216,N_7067,N_7720);
and U8217 (N_8217,N_7541,N_7420);
nand U8218 (N_8218,N_7854,N_7211);
or U8219 (N_8219,N_7906,N_7008);
nand U8220 (N_8220,N_7686,N_7885);
and U8221 (N_8221,N_7314,N_7773);
or U8222 (N_8222,N_7476,N_7283);
nor U8223 (N_8223,N_7093,N_7379);
or U8224 (N_8224,N_7544,N_7887);
and U8225 (N_8225,N_7485,N_7599);
nor U8226 (N_8226,N_7930,N_7560);
or U8227 (N_8227,N_7465,N_7597);
nand U8228 (N_8228,N_7778,N_7853);
and U8229 (N_8229,N_7706,N_7610);
and U8230 (N_8230,N_7529,N_7102);
nor U8231 (N_8231,N_7814,N_7022);
or U8232 (N_8232,N_7917,N_7939);
xnor U8233 (N_8233,N_7957,N_7630);
or U8234 (N_8234,N_7966,N_7272);
nand U8235 (N_8235,N_7595,N_7191);
nor U8236 (N_8236,N_7745,N_7572);
and U8237 (N_8237,N_7785,N_7625);
nor U8238 (N_8238,N_7433,N_7140);
and U8239 (N_8239,N_7077,N_7498);
or U8240 (N_8240,N_7204,N_7075);
nand U8241 (N_8241,N_7762,N_7255);
nor U8242 (N_8242,N_7492,N_7810);
and U8243 (N_8243,N_7346,N_7214);
or U8244 (N_8244,N_7114,N_7440);
and U8245 (N_8245,N_7352,N_7979);
nand U8246 (N_8246,N_7052,N_7816);
or U8247 (N_8247,N_7068,N_7134);
nand U8248 (N_8248,N_7327,N_7811);
nand U8249 (N_8249,N_7691,N_7535);
nand U8250 (N_8250,N_7638,N_7650);
nand U8251 (N_8251,N_7338,N_7382);
or U8252 (N_8252,N_7614,N_7280);
or U8253 (N_8253,N_7174,N_7257);
and U8254 (N_8254,N_7509,N_7297);
and U8255 (N_8255,N_7912,N_7088);
nor U8256 (N_8256,N_7035,N_7206);
nand U8257 (N_8257,N_7284,N_7380);
or U8258 (N_8258,N_7501,N_7161);
nor U8259 (N_8259,N_7188,N_7162);
and U8260 (N_8260,N_7332,N_7669);
nand U8261 (N_8261,N_7575,N_7999);
nor U8262 (N_8262,N_7294,N_7287);
and U8263 (N_8263,N_7243,N_7968);
and U8264 (N_8264,N_7110,N_7401);
nor U8265 (N_8265,N_7260,N_7403);
and U8266 (N_8266,N_7157,N_7224);
or U8267 (N_8267,N_7807,N_7859);
nor U8268 (N_8268,N_7808,N_7256);
nand U8269 (N_8269,N_7903,N_7009);
nand U8270 (N_8270,N_7713,N_7550);
and U8271 (N_8271,N_7875,N_7493);
nor U8272 (N_8272,N_7011,N_7872);
nand U8273 (N_8273,N_7489,N_7528);
or U8274 (N_8274,N_7946,N_7832);
and U8275 (N_8275,N_7371,N_7696);
or U8276 (N_8276,N_7890,N_7987);
nor U8277 (N_8277,N_7539,N_7106);
xor U8278 (N_8278,N_7582,N_7593);
xnor U8279 (N_8279,N_7179,N_7835);
or U8280 (N_8280,N_7847,N_7137);
nor U8281 (N_8281,N_7840,N_7557);
or U8282 (N_8282,N_7508,N_7404);
or U8283 (N_8283,N_7556,N_7056);
or U8284 (N_8284,N_7014,N_7281);
or U8285 (N_8285,N_7333,N_7086);
and U8286 (N_8286,N_7736,N_7573);
xor U8287 (N_8287,N_7851,N_7672);
nor U8288 (N_8288,N_7900,N_7153);
and U8289 (N_8289,N_7415,N_7292);
and U8290 (N_8290,N_7682,N_7225);
nor U8291 (N_8291,N_7530,N_7347);
xor U8292 (N_8292,N_7402,N_7083);
nor U8293 (N_8293,N_7715,N_7514);
nor U8294 (N_8294,N_7620,N_7105);
nand U8295 (N_8295,N_7613,N_7000);
xor U8296 (N_8296,N_7274,N_7349);
nor U8297 (N_8297,N_7919,N_7144);
and U8298 (N_8298,N_7653,N_7450);
xor U8299 (N_8299,N_7699,N_7414);
and U8300 (N_8300,N_7512,N_7131);
or U8301 (N_8301,N_7892,N_7722);
and U8302 (N_8302,N_7734,N_7792);
xnor U8303 (N_8303,N_7702,N_7199);
nand U8304 (N_8304,N_7991,N_7619);
and U8305 (N_8305,N_7937,N_7462);
and U8306 (N_8306,N_7055,N_7718);
xor U8307 (N_8307,N_7815,N_7391);
or U8308 (N_8308,N_7570,N_7558);
xor U8309 (N_8309,N_7384,N_7757);
nand U8310 (N_8310,N_7375,N_7646);
nor U8311 (N_8311,N_7626,N_7879);
xnor U8312 (N_8312,N_7864,N_7122);
xor U8313 (N_8313,N_7034,N_7452);
and U8314 (N_8314,N_7988,N_7163);
and U8315 (N_8315,N_7553,N_7698);
or U8316 (N_8316,N_7360,N_7240);
and U8317 (N_8317,N_7187,N_7931);
and U8318 (N_8318,N_7330,N_7972);
xor U8319 (N_8319,N_7063,N_7149);
nand U8320 (N_8320,N_7487,N_7846);
nor U8321 (N_8321,N_7803,N_7213);
or U8322 (N_8322,N_7351,N_7793);
nand U8323 (N_8323,N_7205,N_7680);
or U8324 (N_8324,N_7618,N_7156);
nor U8325 (N_8325,N_7466,N_7212);
and U8326 (N_8326,N_7549,N_7770);
and U8327 (N_8327,N_7180,N_7200);
or U8328 (N_8328,N_7763,N_7634);
xnor U8329 (N_8329,N_7147,N_7091);
and U8330 (N_8330,N_7469,N_7021);
nor U8331 (N_8331,N_7735,N_7339);
and U8332 (N_8332,N_7266,N_7565);
or U8333 (N_8333,N_7221,N_7898);
nor U8334 (N_8334,N_7319,N_7914);
xnor U8335 (N_8335,N_7005,N_7423);
xor U8336 (N_8336,N_7724,N_7574);
and U8337 (N_8337,N_7709,N_7893);
xnor U8338 (N_8338,N_7563,N_7813);
nor U8339 (N_8339,N_7891,N_7545);
nand U8340 (N_8340,N_7645,N_7152);
nor U8341 (N_8341,N_7446,N_7185);
nor U8342 (N_8342,N_7020,N_7317);
or U8343 (N_8343,N_7719,N_7909);
nand U8344 (N_8344,N_7223,N_7195);
xnor U8345 (N_8345,N_7978,N_7416);
or U8346 (N_8346,N_7130,N_7878);
or U8347 (N_8347,N_7066,N_7181);
xor U8348 (N_8348,N_7948,N_7119);
nor U8349 (N_8349,N_7436,N_7655);
nand U8350 (N_8350,N_7325,N_7173);
nand U8351 (N_8351,N_7990,N_7084);
or U8352 (N_8352,N_7985,N_7455);
nor U8353 (N_8353,N_7017,N_7639);
nor U8354 (N_8354,N_7701,N_7150);
nor U8355 (N_8355,N_7132,N_7880);
or U8356 (N_8356,N_7726,N_7710);
nand U8357 (N_8357,N_7104,N_7412);
or U8358 (N_8358,N_7337,N_7120);
nor U8359 (N_8359,N_7831,N_7867);
nor U8360 (N_8360,N_7282,N_7822);
or U8361 (N_8361,N_7690,N_7510);
nor U8362 (N_8362,N_7907,N_7176);
and U8363 (N_8363,N_7043,N_7186);
or U8364 (N_8364,N_7608,N_7071);
nor U8365 (N_8365,N_7896,N_7733);
xor U8366 (N_8366,N_7824,N_7602);
or U8367 (N_8367,N_7527,N_7850);
nand U8368 (N_8368,N_7836,N_7756);
nand U8369 (N_8369,N_7123,N_7357);
xnor U8370 (N_8370,N_7004,N_7505);
nor U8371 (N_8371,N_7576,N_7449);
xor U8372 (N_8372,N_7927,N_7821);
xnor U8373 (N_8373,N_7087,N_7571);
nor U8374 (N_8374,N_7685,N_7621);
nand U8375 (N_8375,N_7569,N_7244);
or U8376 (N_8376,N_7234,N_7254);
nand U8377 (N_8377,N_7947,N_7784);
or U8378 (N_8378,N_7982,N_7849);
nand U8379 (N_8379,N_7042,N_7798);
xor U8380 (N_8380,N_7092,N_7809);
nor U8381 (N_8381,N_7353,N_7746);
xor U8382 (N_8382,N_7737,N_7329);
or U8383 (N_8383,N_7606,N_7061);
and U8384 (N_8384,N_7194,N_7230);
nand U8385 (N_8385,N_7264,N_7542);
nor U8386 (N_8386,N_7295,N_7661);
nand U8387 (N_8387,N_7693,N_7799);
or U8388 (N_8388,N_7945,N_7942);
xor U8389 (N_8389,N_7024,N_7289);
xnor U8390 (N_8390,N_7215,N_7496);
or U8391 (N_8391,N_7242,N_7047);
nor U8392 (N_8392,N_7345,N_7855);
nand U8393 (N_8393,N_7116,N_7865);
and U8394 (N_8394,N_7381,N_7768);
nand U8395 (N_8395,N_7148,N_7023);
or U8396 (N_8396,N_7923,N_7677);
xnor U8397 (N_8397,N_7517,N_7635);
nand U8398 (N_8398,N_7579,N_7921);
nand U8399 (N_8399,N_7838,N_7367);
xor U8400 (N_8400,N_7470,N_7178);
xor U8401 (N_8401,N_7303,N_7456);
nand U8402 (N_8402,N_7801,N_7511);
and U8403 (N_8403,N_7430,N_7080);
xnor U8404 (N_8404,N_7681,N_7688);
and U8405 (N_8405,N_7390,N_7451);
nor U8406 (N_8406,N_7649,N_7109);
or U8407 (N_8407,N_7918,N_7627);
xnor U8408 (N_8408,N_7172,N_7834);
and U8409 (N_8409,N_7984,N_7534);
and U8410 (N_8410,N_7910,N_7447);
xor U8411 (N_8411,N_7749,N_7383);
nand U8412 (N_8412,N_7036,N_7460);
nand U8413 (N_8413,N_7475,N_7190);
and U8414 (N_8414,N_7960,N_7342);
or U8415 (N_8415,N_7306,N_7589);
and U8416 (N_8416,N_7675,N_7754);
or U8417 (N_8417,N_7624,N_7429);
nand U8418 (N_8418,N_7135,N_7751);
and U8419 (N_8419,N_7934,N_7220);
or U8420 (N_8420,N_7007,N_7445);
xor U8421 (N_8421,N_7705,N_7328);
nor U8422 (N_8422,N_7954,N_7981);
and U8423 (N_8423,N_7989,N_7010);
nand U8424 (N_8424,N_7495,N_7044);
or U8425 (N_8425,N_7309,N_7409);
or U8426 (N_8426,N_7311,N_7457);
nand U8427 (N_8427,N_7058,N_7740);
nand U8428 (N_8428,N_7884,N_7340);
nand U8429 (N_8429,N_7422,N_7752);
or U8430 (N_8430,N_7209,N_7616);
and U8431 (N_8431,N_7766,N_7189);
nor U8432 (N_8432,N_7032,N_7805);
xnor U8433 (N_8433,N_7531,N_7388);
and U8434 (N_8434,N_7953,N_7936);
nor U8435 (N_8435,N_7127,N_7562);
or U8436 (N_8436,N_7316,N_7841);
xnor U8437 (N_8437,N_7697,N_7235);
nand U8438 (N_8438,N_7118,N_7331);
nor U8439 (N_8439,N_7112,N_7113);
nand U8440 (N_8440,N_7473,N_7796);
and U8441 (N_8441,N_7522,N_7444);
xnor U8442 (N_8442,N_7897,N_7848);
and U8443 (N_8443,N_7916,N_7915);
nor U8444 (N_8444,N_7321,N_7241);
or U8445 (N_8445,N_7070,N_7431);
and U8446 (N_8446,N_7888,N_7873);
or U8447 (N_8447,N_7053,N_7830);
nor U8448 (N_8448,N_7742,N_7097);
or U8449 (N_8449,N_7164,N_7546);
nand U8450 (N_8450,N_7567,N_7270);
nand U8451 (N_8451,N_7459,N_7300);
and U8452 (N_8452,N_7583,N_7540);
or U8453 (N_8453,N_7437,N_7483);
or U8454 (N_8454,N_7739,N_7802);
or U8455 (N_8455,N_7399,N_7169);
and U8456 (N_8456,N_7394,N_7320);
or U8457 (N_8457,N_7322,N_7151);
and U8458 (N_8458,N_7977,N_7057);
nor U8459 (N_8459,N_7755,N_7829);
or U8460 (N_8460,N_7727,N_7633);
nand U8461 (N_8461,N_7310,N_7165);
or U8462 (N_8462,N_7741,N_7308);
nor U8463 (N_8463,N_7486,N_7631);
and U8464 (N_8464,N_7335,N_7438);
nand U8465 (N_8465,N_7261,N_7601);
xor U8466 (N_8466,N_7554,N_7249);
or U8467 (N_8467,N_7643,N_7278);
and U8468 (N_8468,N_7288,N_7027);
or U8469 (N_8469,N_7521,N_7372);
xor U8470 (N_8470,N_7201,N_7837);
nand U8471 (N_8471,N_7993,N_7160);
and U8472 (N_8472,N_7307,N_7250);
and U8473 (N_8473,N_7393,N_7072);
nand U8474 (N_8474,N_7275,N_7605);
xnor U8475 (N_8475,N_7125,N_7271);
nand U8476 (N_8476,N_7344,N_7843);
nor U8477 (N_8477,N_7723,N_7516);
nand U8478 (N_8478,N_7427,N_7935);
nor U8479 (N_8479,N_7684,N_7820);
or U8480 (N_8480,N_7983,N_7525);
nand U8481 (N_8481,N_7478,N_7069);
and U8482 (N_8482,N_7458,N_7051);
nor U8483 (N_8483,N_7258,N_7924);
and U8484 (N_8484,N_7580,N_7018);
and U8485 (N_8485,N_7659,N_7551);
nor U8486 (N_8486,N_7299,N_7839);
and U8487 (N_8487,N_7513,N_7276);
or U8488 (N_8488,N_7350,N_7305);
or U8489 (N_8489,N_7408,N_7975);
xor U8490 (N_8490,N_7518,N_7765);
xnor U8491 (N_8491,N_7588,N_7167);
nor U8492 (N_8492,N_7964,N_7252);
nor U8493 (N_8493,N_7886,N_7783);
xnor U8494 (N_8494,N_7592,N_7239);
nand U8495 (N_8495,N_7994,N_7929);
and U8496 (N_8496,N_7400,N_7248);
xnor U8497 (N_8497,N_7995,N_7411);
xnor U8498 (N_8498,N_7192,N_7298);
or U8499 (N_8499,N_7790,N_7369);
nor U8500 (N_8500,N_7164,N_7706);
nor U8501 (N_8501,N_7110,N_7341);
xnor U8502 (N_8502,N_7391,N_7818);
nor U8503 (N_8503,N_7676,N_7013);
or U8504 (N_8504,N_7707,N_7676);
nand U8505 (N_8505,N_7436,N_7557);
xnor U8506 (N_8506,N_7708,N_7190);
or U8507 (N_8507,N_7664,N_7536);
or U8508 (N_8508,N_7487,N_7067);
xor U8509 (N_8509,N_7440,N_7933);
nand U8510 (N_8510,N_7312,N_7463);
and U8511 (N_8511,N_7042,N_7895);
xor U8512 (N_8512,N_7227,N_7555);
and U8513 (N_8513,N_7688,N_7581);
xor U8514 (N_8514,N_7121,N_7212);
nand U8515 (N_8515,N_7015,N_7294);
and U8516 (N_8516,N_7557,N_7360);
nand U8517 (N_8517,N_7329,N_7490);
xor U8518 (N_8518,N_7356,N_7722);
nor U8519 (N_8519,N_7949,N_7221);
and U8520 (N_8520,N_7485,N_7832);
nor U8521 (N_8521,N_7389,N_7945);
and U8522 (N_8522,N_7033,N_7397);
xor U8523 (N_8523,N_7891,N_7838);
and U8524 (N_8524,N_7650,N_7370);
or U8525 (N_8525,N_7856,N_7579);
nor U8526 (N_8526,N_7140,N_7137);
or U8527 (N_8527,N_7826,N_7017);
nand U8528 (N_8528,N_7307,N_7892);
nor U8529 (N_8529,N_7901,N_7168);
and U8530 (N_8530,N_7140,N_7772);
and U8531 (N_8531,N_7615,N_7088);
nor U8532 (N_8532,N_7288,N_7415);
nor U8533 (N_8533,N_7919,N_7623);
xnor U8534 (N_8534,N_7995,N_7245);
xor U8535 (N_8535,N_7063,N_7224);
nor U8536 (N_8536,N_7081,N_7868);
nor U8537 (N_8537,N_7476,N_7181);
nand U8538 (N_8538,N_7293,N_7688);
and U8539 (N_8539,N_7414,N_7750);
and U8540 (N_8540,N_7041,N_7965);
nor U8541 (N_8541,N_7071,N_7134);
nor U8542 (N_8542,N_7108,N_7889);
or U8543 (N_8543,N_7376,N_7921);
nor U8544 (N_8544,N_7270,N_7481);
xor U8545 (N_8545,N_7631,N_7221);
nor U8546 (N_8546,N_7751,N_7182);
and U8547 (N_8547,N_7963,N_7302);
xor U8548 (N_8548,N_7271,N_7558);
or U8549 (N_8549,N_7178,N_7894);
xor U8550 (N_8550,N_7166,N_7319);
nand U8551 (N_8551,N_7844,N_7234);
or U8552 (N_8552,N_7322,N_7763);
nand U8553 (N_8553,N_7481,N_7487);
and U8554 (N_8554,N_7813,N_7696);
xor U8555 (N_8555,N_7943,N_7014);
xor U8556 (N_8556,N_7651,N_7097);
xnor U8557 (N_8557,N_7755,N_7900);
and U8558 (N_8558,N_7850,N_7439);
xor U8559 (N_8559,N_7247,N_7461);
nand U8560 (N_8560,N_7835,N_7167);
nand U8561 (N_8561,N_7322,N_7284);
and U8562 (N_8562,N_7546,N_7517);
nor U8563 (N_8563,N_7443,N_7600);
nor U8564 (N_8564,N_7473,N_7161);
or U8565 (N_8565,N_7215,N_7040);
nand U8566 (N_8566,N_7538,N_7937);
xnor U8567 (N_8567,N_7766,N_7378);
nor U8568 (N_8568,N_7997,N_7373);
xor U8569 (N_8569,N_7015,N_7342);
and U8570 (N_8570,N_7248,N_7835);
and U8571 (N_8571,N_7671,N_7687);
nor U8572 (N_8572,N_7923,N_7660);
and U8573 (N_8573,N_7375,N_7449);
or U8574 (N_8574,N_7863,N_7396);
or U8575 (N_8575,N_7368,N_7439);
xor U8576 (N_8576,N_7231,N_7300);
and U8577 (N_8577,N_7536,N_7745);
xor U8578 (N_8578,N_7798,N_7696);
xnor U8579 (N_8579,N_7667,N_7768);
and U8580 (N_8580,N_7155,N_7275);
and U8581 (N_8581,N_7926,N_7927);
nor U8582 (N_8582,N_7727,N_7105);
and U8583 (N_8583,N_7723,N_7162);
and U8584 (N_8584,N_7459,N_7742);
and U8585 (N_8585,N_7021,N_7217);
nand U8586 (N_8586,N_7501,N_7332);
or U8587 (N_8587,N_7237,N_7343);
nand U8588 (N_8588,N_7346,N_7627);
xor U8589 (N_8589,N_7682,N_7757);
xor U8590 (N_8590,N_7722,N_7050);
xnor U8591 (N_8591,N_7201,N_7573);
nand U8592 (N_8592,N_7398,N_7314);
nor U8593 (N_8593,N_7585,N_7878);
and U8594 (N_8594,N_7899,N_7790);
or U8595 (N_8595,N_7040,N_7173);
nor U8596 (N_8596,N_7848,N_7971);
and U8597 (N_8597,N_7976,N_7098);
or U8598 (N_8598,N_7048,N_7576);
and U8599 (N_8599,N_7351,N_7700);
nor U8600 (N_8600,N_7944,N_7463);
or U8601 (N_8601,N_7471,N_7527);
nor U8602 (N_8602,N_7273,N_7368);
or U8603 (N_8603,N_7696,N_7627);
nand U8604 (N_8604,N_7903,N_7269);
xnor U8605 (N_8605,N_7292,N_7601);
xor U8606 (N_8606,N_7985,N_7286);
and U8607 (N_8607,N_7106,N_7519);
xnor U8608 (N_8608,N_7310,N_7947);
nand U8609 (N_8609,N_7270,N_7259);
and U8610 (N_8610,N_7812,N_7639);
nand U8611 (N_8611,N_7988,N_7860);
nor U8612 (N_8612,N_7837,N_7760);
xor U8613 (N_8613,N_7368,N_7894);
xor U8614 (N_8614,N_7836,N_7153);
and U8615 (N_8615,N_7030,N_7437);
xnor U8616 (N_8616,N_7464,N_7620);
xnor U8617 (N_8617,N_7530,N_7769);
nor U8618 (N_8618,N_7084,N_7698);
nand U8619 (N_8619,N_7526,N_7618);
and U8620 (N_8620,N_7670,N_7163);
and U8621 (N_8621,N_7106,N_7617);
nand U8622 (N_8622,N_7969,N_7395);
nand U8623 (N_8623,N_7636,N_7118);
and U8624 (N_8624,N_7772,N_7291);
and U8625 (N_8625,N_7337,N_7493);
xnor U8626 (N_8626,N_7510,N_7200);
nand U8627 (N_8627,N_7944,N_7662);
nor U8628 (N_8628,N_7179,N_7330);
or U8629 (N_8629,N_7676,N_7102);
nor U8630 (N_8630,N_7830,N_7603);
nor U8631 (N_8631,N_7158,N_7808);
or U8632 (N_8632,N_7009,N_7466);
or U8633 (N_8633,N_7314,N_7723);
nand U8634 (N_8634,N_7796,N_7776);
nand U8635 (N_8635,N_7242,N_7930);
and U8636 (N_8636,N_7802,N_7568);
xnor U8637 (N_8637,N_7274,N_7457);
nand U8638 (N_8638,N_7383,N_7605);
nand U8639 (N_8639,N_7539,N_7134);
or U8640 (N_8640,N_7857,N_7975);
nand U8641 (N_8641,N_7298,N_7797);
or U8642 (N_8642,N_7292,N_7066);
nor U8643 (N_8643,N_7920,N_7029);
nand U8644 (N_8644,N_7149,N_7088);
and U8645 (N_8645,N_7326,N_7689);
and U8646 (N_8646,N_7985,N_7204);
nor U8647 (N_8647,N_7574,N_7967);
and U8648 (N_8648,N_7622,N_7383);
nand U8649 (N_8649,N_7140,N_7343);
nand U8650 (N_8650,N_7542,N_7683);
and U8651 (N_8651,N_7967,N_7640);
and U8652 (N_8652,N_7175,N_7306);
nor U8653 (N_8653,N_7897,N_7939);
and U8654 (N_8654,N_7412,N_7061);
nand U8655 (N_8655,N_7662,N_7443);
nand U8656 (N_8656,N_7085,N_7844);
or U8657 (N_8657,N_7726,N_7580);
xor U8658 (N_8658,N_7849,N_7661);
nor U8659 (N_8659,N_7626,N_7834);
nand U8660 (N_8660,N_7627,N_7014);
nor U8661 (N_8661,N_7627,N_7380);
and U8662 (N_8662,N_7345,N_7567);
nand U8663 (N_8663,N_7950,N_7427);
nand U8664 (N_8664,N_7342,N_7139);
nor U8665 (N_8665,N_7643,N_7046);
nand U8666 (N_8666,N_7636,N_7648);
and U8667 (N_8667,N_7957,N_7509);
nand U8668 (N_8668,N_7879,N_7732);
xor U8669 (N_8669,N_7395,N_7449);
nor U8670 (N_8670,N_7449,N_7770);
xor U8671 (N_8671,N_7656,N_7079);
nand U8672 (N_8672,N_7170,N_7376);
nor U8673 (N_8673,N_7161,N_7214);
or U8674 (N_8674,N_7975,N_7244);
nor U8675 (N_8675,N_7224,N_7015);
xnor U8676 (N_8676,N_7106,N_7431);
and U8677 (N_8677,N_7406,N_7663);
or U8678 (N_8678,N_7302,N_7426);
nand U8679 (N_8679,N_7021,N_7538);
xnor U8680 (N_8680,N_7670,N_7212);
or U8681 (N_8681,N_7005,N_7304);
or U8682 (N_8682,N_7847,N_7896);
xor U8683 (N_8683,N_7120,N_7631);
and U8684 (N_8684,N_7584,N_7371);
nand U8685 (N_8685,N_7185,N_7712);
or U8686 (N_8686,N_7875,N_7720);
and U8687 (N_8687,N_7913,N_7185);
nor U8688 (N_8688,N_7028,N_7177);
nand U8689 (N_8689,N_7282,N_7976);
and U8690 (N_8690,N_7576,N_7688);
nand U8691 (N_8691,N_7751,N_7451);
or U8692 (N_8692,N_7245,N_7013);
xnor U8693 (N_8693,N_7662,N_7180);
or U8694 (N_8694,N_7516,N_7310);
nor U8695 (N_8695,N_7612,N_7864);
nand U8696 (N_8696,N_7453,N_7484);
nand U8697 (N_8697,N_7120,N_7432);
and U8698 (N_8698,N_7143,N_7921);
and U8699 (N_8699,N_7582,N_7594);
nand U8700 (N_8700,N_7684,N_7903);
or U8701 (N_8701,N_7302,N_7865);
and U8702 (N_8702,N_7631,N_7877);
or U8703 (N_8703,N_7927,N_7941);
nand U8704 (N_8704,N_7128,N_7680);
nand U8705 (N_8705,N_7467,N_7017);
xor U8706 (N_8706,N_7770,N_7946);
nand U8707 (N_8707,N_7668,N_7990);
nand U8708 (N_8708,N_7240,N_7106);
or U8709 (N_8709,N_7742,N_7664);
xor U8710 (N_8710,N_7002,N_7934);
or U8711 (N_8711,N_7517,N_7385);
and U8712 (N_8712,N_7743,N_7348);
xor U8713 (N_8713,N_7646,N_7633);
or U8714 (N_8714,N_7348,N_7991);
or U8715 (N_8715,N_7930,N_7074);
nor U8716 (N_8716,N_7431,N_7657);
or U8717 (N_8717,N_7076,N_7406);
nor U8718 (N_8718,N_7276,N_7079);
xnor U8719 (N_8719,N_7536,N_7710);
nor U8720 (N_8720,N_7543,N_7894);
xnor U8721 (N_8721,N_7178,N_7053);
nand U8722 (N_8722,N_7151,N_7453);
nand U8723 (N_8723,N_7124,N_7397);
nand U8724 (N_8724,N_7199,N_7736);
xor U8725 (N_8725,N_7580,N_7524);
and U8726 (N_8726,N_7941,N_7986);
xnor U8727 (N_8727,N_7973,N_7480);
and U8728 (N_8728,N_7736,N_7525);
and U8729 (N_8729,N_7997,N_7425);
xor U8730 (N_8730,N_7685,N_7566);
and U8731 (N_8731,N_7447,N_7220);
and U8732 (N_8732,N_7493,N_7664);
nor U8733 (N_8733,N_7046,N_7195);
xor U8734 (N_8734,N_7243,N_7902);
nand U8735 (N_8735,N_7809,N_7554);
nor U8736 (N_8736,N_7572,N_7206);
nand U8737 (N_8737,N_7694,N_7632);
nor U8738 (N_8738,N_7981,N_7707);
and U8739 (N_8739,N_7287,N_7231);
nor U8740 (N_8740,N_7126,N_7996);
xnor U8741 (N_8741,N_7065,N_7981);
nor U8742 (N_8742,N_7370,N_7523);
nor U8743 (N_8743,N_7818,N_7446);
xor U8744 (N_8744,N_7013,N_7326);
nor U8745 (N_8745,N_7143,N_7449);
xnor U8746 (N_8746,N_7100,N_7061);
or U8747 (N_8747,N_7316,N_7929);
nor U8748 (N_8748,N_7575,N_7743);
and U8749 (N_8749,N_7685,N_7968);
or U8750 (N_8750,N_7207,N_7736);
or U8751 (N_8751,N_7964,N_7562);
xor U8752 (N_8752,N_7628,N_7745);
nand U8753 (N_8753,N_7103,N_7936);
or U8754 (N_8754,N_7366,N_7413);
or U8755 (N_8755,N_7240,N_7237);
nand U8756 (N_8756,N_7207,N_7471);
and U8757 (N_8757,N_7869,N_7867);
xnor U8758 (N_8758,N_7755,N_7460);
nand U8759 (N_8759,N_7920,N_7153);
xor U8760 (N_8760,N_7641,N_7939);
nor U8761 (N_8761,N_7820,N_7260);
xor U8762 (N_8762,N_7226,N_7903);
nor U8763 (N_8763,N_7304,N_7256);
xnor U8764 (N_8764,N_7202,N_7538);
nand U8765 (N_8765,N_7247,N_7554);
nand U8766 (N_8766,N_7087,N_7546);
xnor U8767 (N_8767,N_7178,N_7844);
or U8768 (N_8768,N_7981,N_7317);
nor U8769 (N_8769,N_7705,N_7108);
xor U8770 (N_8770,N_7465,N_7767);
or U8771 (N_8771,N_7474,N_7785);
and U8772 (N_8772,N_7033,N_7584);
or U8773 (N_8773,N_7806,N_7197);
nor U8774 (N_8774,N_7693,N_7875);
and U8775 (N_8775,N_7878,N_7189);
nand U8776 (N_8776,N_7008,N_7252);
and U8777 (N_8777,N_7634,N_7713);
and U8778 (N_8778,N_7835,N_7244);
nand U8779 (N_8779,N_7983,N_7033);
xnor U8780 (N_8780,N_7959,N_7151);
xnor U8781 (N_8781,N_7699,N_7538);
nand U8782 (N_8782,N_7258,N_7313);
and U8783 (N_8783,N_7421,N_7802);
or U8784 (N_8784,N_7167,N_7586);
xor U8785 (N_8785,N_7099,N_7792);
nand U8786 (N_8786,N_7519,N_7921);
nor U8787 (N_8787,N_7012,N_7924);
nand U8788 (N_8788,N_7382,N_7480);
nand U8789 (N_8789,N_7437,N_7789);
xor U8790 (N_8790,N_7687,N_7376);
xnor U8791 (N_8791,N_7642,N_7629);
nor U8792 (N_8792,N_7901,N_7935);
and U8793 (N_8793,N_7813,N_7944);
nor U8794 (N_8794,N_7561,N_7632);
and U8795 (N_8795,N_7871,N_7561);
nor U8796 (N_8796,N_7374,N_7697);
and U8797 (N_8797,N_7612,N_7349);
nand U8798 (N_8798,N_7838,N_7973);
nand U8799 (N_8799,N_7620,N_7837);
or U8800 (N_8800,N_7916,N_7495);
nor U8801 (N_8801,N_7174,N_7927);
xnor U8802 (N_8802,N_7226,N_7689);
xor U8803 (N_8803,N_7195,N_7045);
or U8804 (N_8804,N_7592,N_7036);
or U8805 (N_8805,N_7613,N_7508);
or U8806 (N_8806,N_7122,N_7050);
nand U8807 (N_8807,N_7817,N_7251);
and U8808 (N_8808,N_7878,N_7781);
nand U8809 (N_8809,N_7323,N_7121);
or U8810 (N_8810,N_7990,N_7687);
nand U8811 (N_8811,N_7744,N_7567);
nand U8812 (N_8812,N_7630,N_7215);
xor U8813 (N_8813,N_7690,N_7697);
nand U8814 (N_8814,N_7366,N_7097);
xor U8815 (N_8815,N_7642,N_7278);
nor U8816 (N_8816,N_7808,N_7955);
or U8817 (N_8817,N_7490,N_7849);
xor U8818 (N_8818,N_7742,N_7405);
nand U8819 (N_8819,N_7501,N_7834);
nor U8820 (N_8820,N_7281,N_7323);
xor U8821 (N_8821,N_7360,N_7317);
and U8822 (N_8822,N_7403,N_7197);
or U8823 (N_8823,N_7484,N_7822);
xnor U8824 (N_8824,N_7475,N_7814);
nor U8825 (N_8825,N_7140,N_7129);
and U8826 (N_8826,N_7379,N_7294);
xnor U8827 (N_8827,N_7844,N_7741);
nand U8828 (N_8828,N_7362,N_7651);
and U8829 (N_8829,N_7782,N_7660);
nor U8830 (N_8830,N_7721,N_7026);
or U8831 (N_8831,N_7733,N_7947);
xor U8832 (N_8832,N_7569,N_7723);
and U8833 (N_8833,N_7768,N_7811);
and U8834 (N_8834,N_7153,N_7743);
xor U8835 (N_8835,N_7080,N_7774);
and U8836 (N_8836,N_7841,N_7313);
xnor U8837 (N_8837,N_7665,N_7074);
xor U8838 (N_8838,N_7228,N_7880);
or U8839 (N_8839,N_7353,N_7552);
nand U8840 (N_8840,N_7615,N_7166);
or U8841 (N_8841,N_7101,N_7630);
nor U8842 (N_8842,N_7227,N_7456);
nand U8843 (N_8843,N_7470,N_7369);
nor U8844 (N_8844,N_7216,N_7361);
or U8845 (N_8845,N_7771,N_7148);
or U8846 (N_8846,N_7603,N_7964);
or U8847 (N_8847,N_7386,N_7504);
and U8848 (N_8848,N_7108,N_7142);
and U8849 (N_8849,N_7376,N_7616);
nand U8850 (N_8850,N_7623,N_7566);
xor U8851 (N_8851,N_7309,N_7631);
nor U8852 (N_8852,N_7053,N_7704);
nand U8853 (N_8853,N_7763,N_7959);
nor U8854 (N_8854,N_7932,N_7056);
nor U8855 (N_8855,N_7085,N_7349);
xor U8856 (N_8856,N_7335,N_7683);
nor U8857 (N_8857,N_7318,N_7003);
xnor U8858 (N_8858,N_7471,N_7142);
nand U8859 (N_8859,N_7346,N_7849);
nand U8860 (N_8860,N_7350,N_7240);
xnor U8861 (N_8861,N_7407,N_7344);
xnor U8862 (N_8862,N_7652,N_7346);
and U8863 (N_8863,N_7762,N_7460);
or U8864 (N_8864,N_7541,N_7854);
nor U8865 (N_8865,N_7683,N_7234);
xor U8866 (N_8866,N_7798,N_7353);
and U8867 (N_8867,N_7506,N_7598);
nand U8868 (N_8868,N_7210,N_7443);
and U8869 (N_8869,N_7032,N_7886);
and U8870 (N_8870,N_7668,N_7611);
or U8871 (N_8871,N_7518,N_7752);
xor U8872 (N_8872,N_7291,N_7754);
xor U8873 (N_8873,N_7225,N_7415);
nor U8874 (N_8874,N_7908,N_7329);
nor U8875 (N_8875,N_7745,N_7741);
or U8876 (N_8876,N_7995,N_7724);
or U8877 (N_8877,N_7296,N_7661);
xor U8878 (N_8878,N_7783,N_7929);
xor U8879 (N_8879,N_7881,N_7772);
xnor U8880 (N_8880,N_7628,N_7150);
nand U8881 (N_8881,N_7416,N_7049);
xnor U8882 (N_8882,N_7576,N_7341);
nand U8883 (N_8883,N_7934,N_7819);
nor U8884 (N_8884,N_7953,N_7753);
nor U8885 (N_8885,N_7540,N_7140);
and U8886 (N_8886,N_7554,N_7791);
and U8887 (N_8887,N_7333,N_7072);
nand U8888 (N_8888,N_7698,N_7269);
nand U8889 (N_8889,N_7591,N_7953);
and U8890 (N_8890,N_7976,N_7743);
or U8891 (N_8891,N_7249,N_7704);
nor U8892 (N_8892,N_7416,N_7803);
nor U8893 (N_8893,N_7416,N_7678);
xor U8894 (N_8894,N_7700,N_7491);
nand U8895 (N_8895,N_7834,N_7893);
nand U8896 (N_8896,N_7667,N_7431);
or U8897 (N_8897,N_7079,N_7596);
xnor U8898 (N_8898,N_7712,N_7150);
or U8899 (N_8899,N_7326,N_7857);
and U8900 (N_8900,N_7898,N_7283);
nand U8901 (N_8901,N_7757,N_7978);
nand U8902 (N_8902,N_7475,N_7355);
xnor U8903 (N_8903,N_7043,N_7210);
nand U8904 (N_8904,N_7732,N_7994);
nand U8905 (N_8905,N_7221,N_7908);
or U8906 (N_8906,N_7957,N_7949);
xor U8907 (N_8907,N_7708,N_7587);
and U8908 (N_8908,N_7491,N_7734);
nor U8909 (N_8909,N_7208,N_7523);
or U8910 (N_8910,N_7087,N_7405);
nand U8911 (N_8911,N_7272,N_7689);
or U8912 (N_8912,N_7278,N_7354);
and U8913 (N_8913,N_7035,N_7186);
nand U8914 (N_8914,N_7418,N_7293);
nand U8915 (N_8915,N_7508,N_7524);
nor U8916 (N_8916,N_7026,N_7931);
and U8917 (N_8917,N_7656,N_7878);
nor U8918 (N_8918,N_7770,N_7697);
and U8919 (N_8919,N_7696,N_7397);
and U8920 (N_8920,N_7256,N_7387);
xnor U8921 (N_8921,N_7431,N_7883);
xor U8922 (N_8922,N_7078,N_7179);
nand U8923 (N_8923,N_7698,N_7174);
xnor U8924 (N_8924,N_7315,N_7204);
nand U8925 (N_8925,N_7945,N_7895);
nand U8926 (N_8926,N_7059,N_7483);
xnor U8927 (N_8927,N_7429,N_7899);
nand U8928 (N_8928,N_7092,N_7629);
nand U8929 (N_8929,N_7057,N_7520);
or U8930 (N_8930,N_7590,N_7677);
xor U8931 (N_8931,N_7988,N_7973);
and U8932 (N_8932,N_7202,N_7227);
nor U8933 (N_8933,N_7356,N_7125);
xnor U8934 (N_8934,N_7779,N_7429);
nor U8935 (N_8935,N_7214,N_7898);
xor U8936 (N_8936,N_7227,N_7681);
nor U8937 (N_8937,N_7445,N_7109);
nor U8938 (N_8938,N_7962,N_7722);
nand U8939 (N_8939,N_7519,N_7597);
xnor U8940 (N_8940,N_7172,N_7812);
xor U8941 (N_8941,N_7878,N_7847);
nor U8942 (N_8942,N_7061,N_7256);
nand U8943 (N_8943,N_7609,N_7095);
nand U8944 (N_8944,N_7268,N_7588);
and U8945 (N_8945,N_7197,N_7499);
nor U8946 (N_8946,N_7537,N_7672);
nor U8947 (N_8947,N_7842,N_7958);
nand U8948 (N_8948,N_7128,N_7099);
nand U8949 (N_8949,N_7873,N_7173);
xnor U8950 (N_8950,N_7508,N_7101);
xnor U8951 (N_8951,N_7883,N_7086);
nor U8952 (N_8952,N_7850,N_7697);
xor U8953 (N_8953,N_7220,N_7471);
or U8954 (N_8954,N_7636,N_7225);
and U8955 (N_8955,N_7473,N_7842);
nand U8956 (N_8956,N_7414,N_7093);
or U8957 (N_8957,N_7340,N_7838);
and U8958 (N_8958,N_7502,N_7869);
nor U8959 (N_8959,N_7140,N_7767);
nor U8960 (N_8960,N_7986,N_7624);
or U8961 (N_8961,N_7499,N_7064);
nor U8962 (N_8962,N_7175,N_7254);
and U8963 (N_8963,N_7882,N_7385);
xor U8964 (N_8964,N_7445,N_7158);
and U8965 (N_8965,N_7609,N_7006);
nand U8966 (N_8966,N_7364,N_7207);
and U8967 (N_8967,N_7340,N_7133);
nand U8968 (N_8968,N_7476,N_7505);
xor U8969 (N_8969,N_7576,N_7816);
nand U8970 (N_8970,N_7859,N_7263);
nor U8971 (N_8971,N_7295,N_7077);
or U8972 (N_8972,N_7454,N_7461);
nand U8973 (N_8973,N_7868,N_7056);
nand U8974 (N_8974,N_7428,N_7088);
xnor U8975 (N_8975,N_7658,N_7733);
and U8976 (N_8976,N_7053,N_7976);
and U8977 (N_8977,N_7089,N_7194);
xnor U8978 (N_8978,N_7272,N_7902);
and U8979 (N_8979,N_7084,N_7614);
and U8980 (N_8980,N_7286,N_7704);
or U8981 (N_8981,N_7493,N_7155);
nand U8982 (N_8982,N_7063,N_7807);
nor U8983 (N_8983,N_7766,N_7109);
or U8984 (N_8984,N_7765,N_7137);
xor U8985 (N_8985,N_7061,N_7108);
xor U8986 (N_8986,N_7886,N_7845);
and U8987 (N_8987,N_7767,N_7614);
xor U8988 (N_8988,N_7340,N_7103);
and U8989 (N_8989,N_7641,N_7467);
nand U8990 (N_8990,N_7948,N_7689);
and U8991 (N_8991,N_7446,N_7742);
or U8992 (N_8992,N_7573,N_7971);
nor U8993 (N_8993,N_7055,N_7516);
nand U8994 (N_8994,N_7835,N_7617);
nand U8995 (N_8995,N_7508,N_7980);
nor U8996 (N_8996,N_7856,N_7487);
or U8997 (N_8997,N_7182,N_7759);
nand U8998 (N_8998,N_7365,N_7679);
nand U8999 (N_8999,N_7770,N_7002);
and U9000 (N_9000,N_8988,N_8523);
xor U9001 (N_9001,N_8023,N_8227);
nor U9002 (N_9002,N_8973,N_8424);
nand U9003 (N_9003,N_8977,N_8197);
xor U9004 (N_9004,N_8806,N_8836);
and U9005 (N_9005,N_8264,N_8166);
nor U9006 (N_9006,N_8490,N_8519);
xnor U9007 (N_9007,N_8212,N_8408);
and U9008 (N_9008,N_8110,N_8935);
nor U9009 (N_9009,N_8232,N_8449);
or U9010 (N_9010,N_8575,N_8145);
nor U9011 (N_9011,N_8284,N_8390);
xor U9012 (N_9012,N_8036,N_8272);
xnor U9013 (N_9013,N_8526,N_8769);
nor U9014 (N_9014,N_8505,N_8719);
and U9015 (N_9015,N_8962,N_8684);
xor U9016 (N_9016,N_8326,N_8996);
nand U9017 (N_9017,N_8661,N_8017);
xnor U9018 (N_9018,N_8394,N_8693);
nor U9019 (N_9019,N_8368,N_8225);
xor U9020 (N_9020,N_8095,N_8667);
xnor U9021 (N_9021,N_8196,N_8990);
xnor U9022 (N_9022,N_8048,N_8933);
nand U9023 (N_9023,N_8369,N_8847);
nand U9024 (N_9024,N_8177,N_8537);
or U9025 (N_9025,N_8294,N_8772);
nand U9026 (N_9026,N_8218,N_8361);
and U9027 (N_9027,N_8556,N_8783);
xor U9028 (N_9028,N_8463,N_8222);
and U9029 (N_9029,N_8793,N_8649);
xor U9030 (N_9030,N_8509,N_8100);
or U9031 (N_9031,N_8090,N_8834);
nor U9032 (N_9032,N_8426,N_8487);
xnor U9033 (N_9033,N_8280,N_8897);
and U9034 (N_9034,N_8478,N_8946);
and U9035 (N_9035,N_8815,N_8479);
xnor U9036 (N_9036,N_8091,N_8502);
or U9037 (N_9037,N_8276,N_8186);
nor U9038 (N_9038,N_8053,N_8169);
and U9039 (N_9039,N_8328,N_8830);
xnor U9040 (N_9040,N_8738,N_8752);
nand U9041 (N_9041,N_8200,N_8436);
nand U9042 (N_9042,N_8160,N_8944);
nand U9043 (N_9043,N_8228,N_8079);
nand U9044 (N_9044,N_8253,N_8414);
nand U9045 (N_9045,N_8949,N_8235);
xor U9046 (N_9046,N_8746,N_8252);
or U9047 (N_9047,N_8455,N_8901);
or U9048 (N_9048,N_8675,N_8690);
nand U9049 (N_9049,N_8002,N_8388);
nand U9050 (N_9050,N_8628,N_8040);
or U9051 (N_9051,N_8979,N_8231);
and U9052 (N_9052,N_8476,N_8356);
nor U9053 (N_9053,N_8648,N_8874);
xor U9054 (N_9054,N_8810,N_8199);
nand U9055 (N_9055,N_8150,N_8754);
nand U9056 (N_9056,N_8192,N_8380);
or U9057 (N_9057,N_8560,N_8659);
xnor U9058 (N_9058,N_8640,N_8441);
nor U9059 (N_9059,N_8698,N_8484);
and U9060 (N_9060,N_8205,N_8960);
xnor U9061 (N_9061,N_8006,N_8578);
nor U9062 (N_9062,N_8886,N_8613);
nor U9063 (N_9063,N_8364,N_8113);
nor U9064 (N_9064,N_8384,N_8327);
xnor U9065 (N_9065,N_8561,N_8921);
and U9066 (N_9066,N_8518,N_8085);
and U9067 (N_9067,N_8211,N_8319);
xnor U9068 (N_9068,N_8304,N_8050);
or U9069 (N_9069,N_8516,N_8097);
and U9070 (N_9070,N_8273,N_8315);
xor U9071 (N_9071,N_8459,N_8725);
nand U9072 (N_9072,N_8337,N_8181);
nand U9073 (N_9073,N_8662,N_8279);
and U9074 (N_9074,N_8934,N_8701);
nand U9075 (N_9075,N_8501,N_8498);
nand U9076 (N_9076,N_8541,N_8907);
or U9077 (N_9077,N_8545,N_8358);
xor U9078 (N_9078,N_8872,N_8204);
and U9079 (N_9079,N_8413,N_8587);
nand U9080 (N_9080,N_8795,N_8668);
nand U9081 (N_9081,N_8548,N_8296);
and U9082 (N_9082,N_8396,N_8580);
and U9083 (N_9083,N_8103,N_8001);
nor U9084 (N_9084,N_8345,N_8832);
or U9085 (N_9085,N_8052,N_8187);
or U9086 (N_9086,N_8482,N_8905);
nand U9087 (N_9087,N_8522,N_8767);
xor U9088 (N_9088,N_8081,N_8618);
nand U9089 (N_9089,N_8465,N_8664);
nor U9090 (N_9090,N_8077,N_8722);
or U9091 (N_9091,N_8771,N_8510);
nor U9092 (N_9092,N_8061,N_8507);
xor U9093 (N_9093,N_8665,N_8194);
or U9094 (N_9094,N_8993,N_8234);
nand U9095 (N_9095,N_8534,N_8736);
or U9096 (N_9096,N_8822,N_8098);
or U9097 (N_9097,N_8965,N_8670);
nand U9098 (N_9098,N_8131,N_8566);
xnor U9099 (N_9099,N_8473,N_8481);
or U9100 (N_9100,N_8381,N_8467);
xnor U9101 (N_9101,N_8775,N_8055);
or U9102 (N_9102,N_8343,N_8549);
nand U9103 (N_9103,N_8593,N_8819);
or U9104 (N_9104,N_8309,N_8056);
or U9105 (N_9105,N_8718,N_8342);
nor U9106 (N_9106,N_8334,N_8773);
xnor U9107 (N_9107,N_8401,N_8242);
nor U9108 (N_9108,N_8639,N_8692);
nand U9109 (N_9109,N_8835,N_8683);
xnor U9110 (N_9110,N_8416,N_8951);
nand U9111 (N_9111,N_8729,N_8174);
nor U9112 (N_9112,N_8405,N_8986);
nor U9113 (N_9113,N_8877,N_8215);
nand U9114 (N_9114,N_8604,N_8976);
and U9115 (N_9115,N_8844,N_8622);
and U9116 (N_9116,N_8839,N_8130);
nor U9117 (N_9117,N_8290,N_8353);
nand U9118 (N_9118,N_8882,N_8804);
nor U9119 (N_9119,N_8720,N_8805);
and U9120 (N_9120,N_8258,N_8182);
xnor U9121 (N_9121,N_8803,N_8883);
nor U9122 (N_9122,N_8774,N_8520);
nand U9123 (N_9123,N_8954,N_8313);
or U9124 (N_9124,N_8579,N_8493);
xor U9125 (N_9125,N_8407,N_8306);
xnor U9126 (N_9126,N_8645,N_8428);
and U9127 (N_9127,N_8755,N_8359);
nand U9128 (N_9128,N_8788,N_8321);
nor U9129 (N_9129,N_8293,N_8303);
or U9130 (N_9130,N_8109,N_8539);
xor U9131 (N_9131,N_8101,N_8828);
and U9132 (N_9132,N_8992,N_8959);
nand U9133 (N_9133,N_8574,N_8991);
or U9134 (N_9134,N_8302,N_8014);
and U9135 (N_9135,N_8766,N_8240);
or U9136 (N_9136,N_8923,N_8653);
xnor U9137 (N_9137,N_8311,N_8360);
xnor U9138 (N_9138,N_8325,N_8477);
nand U9139 (N_9139,N_8386,N_8288);
xnor U9140 (N_9140,N_8525,N_8717);
nor U9141 (N_9141,N_8589,N_8600);
and U9142 (N_9142,N_8324,N_8474);
xor U9143 (N_9143,N_8393,N_8121);
nor U9144 (N_9144,N_8597,N_8873);
xnor U9145 (N_9145,N_8444,N_8089);
or U9146 (N_9146,N_8282,N_8320);
nor U9147 (N_9147,N_8590,N_8348);
xnor U9148 (N_9148,N_8535,N_8943);
xor U9149 (N_9149,N_8987,N_8869);
and U9150 (N_9150,N_8049,N_8246);
or U9151 (N_9151,N_8144,N_8123);
or U9152 (N_9152,N_8093,N_8536);
and U9153 (N_9153,N_8676,N_8953);
nor U9154 (N_9154,N_8721,N_8267);
and U9155 (N_9155,N_8281,N_8763);
xnor U9156 (N_9156,N_8112,N_8908);
xor U9157 (N_9157,N_8571,N_8111);
or U9158 (N_9158,N_8796,N_8789);
xnor U9159 (N_9159,N_8982,N_8057);
and U9160 (N_9160,N_8292,N_8856);
or U9161 (N_9161,N_8432,N_8012);
or U9162 (N_9162,N_8642,N_8129);
or U9163 (N_9163,N_8475,N_8924);
and U9164 (N_9164,N_8878,N_8925);
nand U9165 (N_9165,N_8938,N_8157);
nor U9166 (N_9166,N_8894,N_8811);
or U9167 (N_9167,N_8163,N_8028);
nor U9168 (N_9168,N_8714,N_8974);
or U9169 (N_9169,N_8739,N_8703);
xnor U9170 (N_9170,N_8486,N_8786);
xor U9171 (N_9171,N_8608,N_8453);
xnor U9172 (N_9172,N_8699,N_8915);
or U9173 (N_9173,N_8802,N_8004);
nand U9174 (N_9174,N_8623,N_8148);
or U9175 (N_9175,N_8823,N_8415);
or U9176 (N_9176,N_8213,N_8909);
nor U9177 (N_9177,N_8673,N_8896);
or U9178 (N_9178,N_8679,N_8753);
and U9179 (N_9179,N_8619,N_8078);
or U9180 (N_9180,N_8355,N_8708);
and U9181 (N_9181,N_8567,N_8759);
and U9182 (N_9182,N_8239,N_8378);
nor U9183 (N_9183,N_8434,N_8814);
nor U9184 (N_9184,N_8351,N_8377);
or U9185 (N_9185,N_8480,N_8059);
nor U9186 (N_9186,N_8126,N_8691);
or U9187 (N_9187,N_8762,N_8115);
nor U9188 (N_9188,N_8395,N_8149);
and U9189 (N_9189,N_8297,N_8956);
and U9190 (N_9190,N_8451,N_8015);
or U9191 (N_9191,N_8249,N_8241);
xnor U9192 (N_9192,N_8930,N_8626);
xor U9193 (N_9193,N_8372,N_8185);
nand U9194 (N_9194,N_8884,N_8244);
nor U9195 (N_9195,N_8289,N_8968);
and U9196 (N_9196,N_8584,N_8880);
nand U9197 (N_9197,N_8782,N_8462);
nor U9198 (N_9198,N_8072,N_8527);
xnor U9199 (N_9199,N_8120,N_8054);
nand U9200 (N_9200,N_8494,N_8605);
or U9201 (N_9201,N_8207,N_8045);
nand U9202 (N_9202,N_8599,N_8660);
nor U9203 (N_9203,N_8821,N_8411);
nor U9204 (N_9204,N_8517,N_8316);
and U9205 (N_9205,N_8346,N_8403);
nand U9206 (N_9206,N_8562,N_8850);
nand U9207 (N_9207,N_8452,N_8132);
xnor U9208 (N_9208,N_8270,N_8751);
or U9209 (N_9209,N_8601,N_8219);
nor U9210 (N_9210,N_8347,N_8568);
nor U9211 (N_9211,N_8859,N_8866);
and U9212 (N_9212,N_8427,N_8164);
and U9213 (N_9213,N_8891,N_8062);
xnor U9214 (N_9214,N_8175,N_8748);
nand U9215 (N_9215,N_8153,N_8606);
or U9216 (N_9216,N_8170,N_8382);
xor U9217 (N_9217,N_8443,N_8362);
xor U9218 (N_9218,N_8603,N_8269);
or U9219 (N_9219,N_8585,N_8464);
nor U9220 (N_9220,N_8871,N_8615);
nand U9221 (N_9221,N_8696,N_8438);
and U9222 (N_9222,N_8610,N_8939);
nand U9223 (N_9223,N_8245,N_8011);
nor U9224 (N_9224,N_8421,N_8948);
or U9225 (N_9225,N_8142,N_8020);
nand U9226 (N_9226,N_8942,N_8899);
or U9227 (N_9227,N_8955,N_8283);
or U9228 (N_9228,N_8895,N_8067);
nand U9229 (N_9229,N_8543,N_8125);
and U9230 (N_9230,N_8940,N_8581);
and U9231 (N_9231,N_8073,N_8515);
nand U9232 (N_9232,N_8506,N_8741);
nor U9233 (N_9233,N_8391,N_8151);
nand U9234 (N_9234,N_8532,N_8807);
nand U9235 (N_9235,N_8122,N_8663);
nand U9236 (N_9236,N_8423,N_8707);
and U9237 (N_9237,N_8217,N_8224);
or U9238 (N_9238,N_8500,N_8417);
nand U9239 (N_9239,N_8375,N_8134);
xor U9240 (N_9240,N_8461,N_8201);
or U9241 (N_9241,N_8024,N_8614);
and U9242 (N_9242,N_8445,N_8504);
and U9243 (N_9243,N_8140,N_8216);
or U9244 (N_9244,N_8508,N_8027);
and U9245 (N_9245,N_8889,N_8794);
nor U9246 (N_9246,N_8800,N_8879);
nor U9247 (N_9247,N_8226,N_8576);
nor U9248 (N_9248,N_8770,N_8700);
and U9249 (N_9249,N_8529,N_8338);
xnor U9250 (N_9250,N_8229,N_8765);
xnor U9251 (N_9251,N_8641,N_8888);
nor U9252 (N_9252,N_8367,N_8491);
xor U9253 (N_9253,N_8998,N_8105);
nand U9254 (N_9254,N_8638,N_8984);
xnor U9255 (N_9255,N_8650,N_8787);
nand U9256 (N_9256,N_8885,N_8032);
nand U9257 (N_9257,N_8733,N_8096);
xnor U9258 (N_9258,N_8503,N_8277);
nor U9259 (N_9259,N_8980,N_8392);
nand U9260 (N_9260,N_8577,N_8981);
nand U9261 (N_9261,N_8617,N_8627);
or U9262 (N_9262,N_8176,N_8730);
and U9263 (N_9263,N_8634,N_8747);
nand U9264 (N_9264,N_8009,N_8827);
or U9265 (N_9265,N_8159,N_8791);
nor U9266 (N_9266,N_8760,N_8088);
and U9267 (N_9267,N_8195,N_8727);
or U9268 (N_9268,N_8329,N_8983);
and U9269 (N_9269,N_8582,N_8333);
xnor U9270 (N_9270,N_8087,N_8551);
or U9271 (N_9271,N_8420,N_8595);
or U9272 (N_9272,N_8454,N_8687);
nor U9273 (N_9273,N_8573,N_8521);
nand U9274 (N_9274,N_8128,N_8124);
nor U9275 (N_9275,N_8435,N_8547);
and U9276 (N_9276,N_8488,N_8928);
or U9277 (N_9277,N_8060,N_8354);
nor U9278 (N_9278,N_8929,N_8404);
xor U9279 (N_9279,N_8654,N_8624);
nand U9280 (N_9280,N_8588,N_8075);
nor U9281 (N_9281,N_8855,N_8094);
and U9282 (N_9282,N_8625,N_8511);
and U9283 (N_9283,N_8937,N_8076);
or U9284 (N_9284,N_8322,N_8133);
nor U9285 (N_9285,N_8412,N_8189);
xnor U9286 (N_9286,N_8868,N_8630);
nor U9287 (N_9287,N_8188,N_8307);
and U9288 (N_9288,N_8167,N_8039);
nand U9289 (N_9289,N_8643,N_8887);
xnor U9290 (N_9290,N_8236,N_8496);
xor U9291 (N_9291,N_8745,N_8171);
nand U9292 (N_9292,N_8447,N_8742);
xnor U9293 (N_9293,N_8564,N_8682);
and U9294 (N_9294,N_8472,N_8410);
nor U9295 (N_9295,N_8591,N_8021);
nand U9296 (N_9296,N_8402,N_8495);
or U9297 (N_9297,N_8947,N_8931);
and U9298 (N_9298,N_8489,N_8265);
nand U9299 (N_9299,N_8070,N_8812);
and U9300 (N_9300,N_8744,N_8713);
and U9301 (N_9301,N_8371,N_8310);
nor U9302 (N_9302,N_8499,N_8813);
or U9303 (N_9303,N_8042,N_8620);
nand U9304 (N_9304,N_8243,N_8251);
nor U9305 (N_9305,N_8260,N_8165);
and U9306 (N_9306,N_8612,N_8340);
or U9307 (N_9307,N_8433,N_8764);
nor U9308 (N_9308,N_8332,N_8958);
and U9309 (N_9309,N_8155,N_8865);
and U9310 (N_9310,N_8308,N_8971);
xnor U9311 (N_9311,N_8798,N_8530);
and U9312 (N_9312,N_8671,N_8695);
nand U9313 (N_9313,N_8035,N_8826);
nand U9314 (N_9314,N_8680,N_8287);
or U9315 (N_9315,N_8425,N_8557);
nand U9316 (N_9316,N_8256,N_8734);
nand U9317 (N_9317,N_8468,N_8689);
nand U9318 (N_9318,N_8756,N_8092);
or U9319 (N_9319,N_8154,N_8046);
xor U9320 (N_9320,N_8349,N_8598);
nor U9321 (N_9321,N_8350,N_8817);
xor U9322 (N_9322,N_8191,N_8596);
nor U9323 (N_9323,N_8570,N_8758);
or U9324 (N_9324,N_8779,N_8672);
or U9325 (N_9325,N_8274,N_8084);
nor U9326 (N_9326,N_8331,N_8305);
xnor U9327 (N_9327,N_8824,N_8852);
xor U9328 (N_9328,N_8278,N_8065);
xor U9329 (N_9329,N_8193,N_8694);
nand U9330 (N_9330,N_8621,N_8632);
nor U9331 (N_9331,N_8261,N_8026);
nand U9332 (N_9332,N_8941,N_8291);
nor U9333 (N_9333,N_8792,N_8178);
and U9334 (N_9334,N_8848,N_8460);
and U9335 (N_9335,N_8183,N_8172);
and U9336 (N_9336,N_8715,N_8554);
and U9337 (N_9337,N_8969,N_8285);
xor U9338 (N_9338,N_8711,N_8858);
and U9339 (N_9339,N_8903,N_8458);
nor U9340 (N_9340,N_8034,N_8341);
nor U9341 (N_9341,N_8259,N_8063);
xnor U9342 (N_9342,N_8920,N_8318);
and U9343 (N_9343,N_8400,N_8857);
and U9344 (N_9344,N_8190,N_8854);
nor U9345 (N_9345,N_8141,N_8558);
nand U9346 (N_9346,N_8064,N_8569);
nand U9347 (N_9347,N_8656,N_8846);
or U9348 (N_9348,N_8801,N_8083);
or U9349 (N_9349,N_8723,N_8471);
or U9350 (N_9350,N_8208,N_8037);
xnor U9351 (N_9351,N_8952,N_8840);
nor U9352 (N_9352,N_8250,N_8651);
and U9353 (N_9353,N_8336,N_8898);
or U9354 (N_9354,N_8118,N_8446);
nor U9355 (N_9355,N_8106,N_8710);
or U9356 (N_9356,N_8071,N_8180);
nor U9357 (N_9357,N_8247,N_8179);
and U9358 (N_9358,N_8728,N_8030);
and U9359 (N_9359,N_8268,N_8743);
or U9360 (N_9360,N_8022,N_8559);
nand U9361 (N_9361,N_8003,N_8709);
or U9362 (N_9362,N_8785,N_8594);
xor U9363 (N_9363,N_8143,N_8849);
and U9364 (N_9364,N_8550,N_8540);
nand U9365 (N_9365,N_8555,N_8528);
nor U9366 (N_9366,N_8221,N_8373);
xor U9367 (N_9367,N_8317,N_8902);
and U9368 (N_9368,N_8398,N_8114);
and U9369 (N_9369,N_8932,N_8790);
nor U9370 (N_9370,N_8138,N_8860);
nand U9371 (N_9371,N_8851,N_8162);
and U9372 (N_9372,N_8917,N_8892);
nor U9373 (N_9373,N_8616,N_8300);
nand U9374 (N_9374,N_8387,N_8966);
xnor U9375 (N_9375,N_8677,N_8314);
or U9376 (N_9376,N_8116,N_8636);
and U9377 (N_9377,N_8950,N_8047);
and U9378 (N_9378,N_8999,N_8963);
nand U9379 (N_9379,N_8043,N_8688);
or U9380 (N_9380,N_8019,N_8437);
nand U9381 (N_9381,N_8910,N_8409);
nor U9382 (N_9382,N_8286,N_8156);
and U9383 (N_9383,N_8013,N_8018);
nor U9384 (N_9384,N_8784,N_8818);
xnor U9385 (N_9385,N_8041,N_8146);
nand U9386 (N_9386,N_8439,N_8911);
and U9387 (N_9387,N_8829,N_8861);
or U9388 (N_9388,N_8135,N_8629);
nand U9389 (N_9389,N_8538,N_8633);
nand U9390 (N_9390,N_8657,N_8658);
nand U9391 (N_9391,N_8137,N_8470);
or U9392 (N_9392,N_8893,N_8716);
xnor U9393 (N_9393,N_8237,N_8586);
or U9394 (N_9394,N_8644,N_8964);
and U9395 (N_9395,N_8702,N_8731);
nand U9396 (N_9396,N_8842,N_8352);
and U9397 (N_9397,N_8737,N_8961);
or U9398 (N_9398,N_8419,N_8257);
xor U9399 (N_9399,N_8972,N_8970);
and U9400 (N_9400,N_8647,N_8271);
or U9401 (N_9401,N_8635,N_8357);
xnor U9402 (N_9402,N_8086,N_8863);
and U9403 (N_9403,N_8099,N_8678);
nand U9404 (N_9404,N_8853,N_8080);
or U9405 (N_9405,N_8202,N_8312);
and U9406 (N_9406,N_8389,N_8609);
xor U9407 (N_9407,N_8295,N_8000);
and U9408 (N_9408,N_8210,N_8147);
and U9409 (N_9409,N_8117,N_8666);
xor U9410 (N_9410,N_8542,N_8833);
xor U9411 (N_9411,N_8108,N_8706);
nor U9412 (N_9412,N_8565,N_8127);
and U9413 (N_9413,N_8563,N_8652);
nand U9414 (N_9414,N_8919,N_8168);
nor U9415 (N_9415,N_8366,N_8385);
nand U9416 (N_9416,N_8139,N_8330);
xor U9417 (N_9417,N_8524,N_8967);
xor U9418 (N_9418,N_8881,N_8497);
or U9419 (N_9419,N_8927,N_8780);
nor U9420 (N_9420,N_8301,N_8450);
nor U9421 (N_9421,N_8740,N_8102);
nor U9422 (N_9422,N_8862,N_8379);
xor U9423 (N_9423,N_8867,N_8044);
and U9424 (N_9424,N_8033,N_8422);
and U9425 (N_9425,N_8916,N_8906);
nor U9426 (N_9426,N_8370,N_8238);
nor U9427 (N_9427,N_8631,N_8038);
nor U9428 (N_9428,N_8875,N_8255);
xor U9429 (N_9429,N_8989,N_8429);
and U9430 (N_9430,N_8797,N_8323);
and U9431 (N_9431,N_8456,N_8206);
or U9432 (N_9432,N_8029,N_8592);
and U9433 (N_9433,N_8781,N_8732);
nand U9434 (N_9434,N_8025,N_8173);
or U9435 (N_9435,N_8749,N_8104);
nand U9436 (N_9436,N_8010,N_8512);
nand U9437 (N_9437,N_8985,N_8082);
and U9438 (N_9438,N_8997,N_8681);
nand U9439 (N_9439,N_8344,N_8669);
xnor U9440 (N_9440,N_8837,N_8607);
xor U9441 (N_9441,N_8418,N_8777);
nand U9442 (N_9442,N_8339,N_8058);
xnor U9443 (N_9443,N_8799,N_8704);
nor U9444 (N_9444,N_8119,N_8158);
xor U9445 (N_9445,N_8904,N_8492);
or U9446 (N_9446,N_8843,N_8263);
nand U9447 (N_9447,N_8203,N_8994);
nor U9448 (N_9448,N_8831,N_8485);
and U9449 (N_9449,N_8220,N_8957);
and U9450 (N_9450,N_8074,N_8890);
xor U9451 (N_9451,N_8900,N_8066);
xor U9452 (N_9452,N_8514,N_8876);
or U9453 (N_9453,N_8583,N_8864);
nor U9454 (N_9454,N_8553,N_8069);
nor U9455 (N_9455,N_8262,N_8572);
xor U9456 (N_9456,N_8724,N_8778);
nor U9457 (N_9457,N_8533,N_8397);
xnor U9458 (N_9458,N_8936,N_8298);
or U9459 (N_9459,N_8735,N_8825);
nor U9460 (N_9460,N_8685,N_8431);
nor U9461 (N_9461,N_8299,N_8383);
and U9462 (N_9462,N_8726,N_8430);
and U9463 (N_9463,N_8016,N_8816);
xor U9464 (N_9464,N_8152,N_8674);
xor U9465 (N_9465,N_8602,N_8808);
and U9466 (N_9466,N_8442,N_8913);
and U9467 (N_9467,N_8161,N_8448);
or U9468 (N_9468,N_8230,N_8544);
nor U9469 (N_9469,N_8761,N_8483);
or U9470 (N_9470,N_8406,N_8198);
and U9471 (N_9471,N_8978,N_8845);
and U9472 (N_9472,N_8637,N_8757);
or U9473 (N_9473,N_8552,N_8051);
and U9474 (N_9474,N_8209,N_8809);
nand U9475 (N_9475,N_8214,N_8248);
nand U9476 (N_9476,N_8686,N_8184);
and U9477 (N_9477,N_8031,N_8870);
and U9478 (N_9478,N_8922,N_8750);
or U9479 (N_9479,N_8466,N_8469);
and U9480 (N_9480,N_8546,N_8926);
and U9481 (N_9481,N_8440,N_8697);
nor U9482 (N_9482,N_8399,N_8975);
or U9483 (N_9483,N_8820,N_8457);
or U9484 (N_9484,N_8914,N_8513);
xnor U9485 (N_9485,N_8531,N_8611);
or U9486 (N_9486,N_8912,N_8655);
xnor U9487 (N_9487,N_8335,N_8376);
and U9488 (N_9488,N_8918,N_8136);
nand U9489 (N_9489,N_8838,N_8275);
nor U9490 (N_9490,N_8705,N_8995);
and U9491 (N_9491,N_8945,N_8007);
or U9492 (N_9492,N_8365,N_8768);
nand U9493 (N_9493,N_8068,N_8254);
nand U9494 (N_9494,N_8646,N_8107);
or U9495 (N_9495,N_8266,N_8233);
and U9496 (N_9496,N_8008,N_8005);
nor U9497 (N_9497,N_8841,N_8374);
xor U9498 (N_9498,N_8363,N_8776);
nand U9499 (N_9499,N_8712,N_8223);
or U9500 (N_9500,N_8303,N_8171);
nand U9501 (N_9501,N_8252,N_8273);
xor U9502 (N_9502,N_8888,N_8715);
xnor U9503 (N_9503,N_8983,N_8108);
nor U9504 (N_9504,N_8167,N_8395);
nor U9505 (N_9505,N_8526,N_8260);
xnor U9506 (N_9506,N_8749,N_8677);
and U9507 (N_9507,N_8188,N_8887);
or U9508 (N_9508,N_8384,N_8617);
or U9509 (N_9509,N_8094,N_8763);
or U9510 (N_9510,N_8035,N_8572);
nand U9511 (N_9511,N_8323,N_8154);
or U9512 (N_9512,N_8764,N_8378);
or U9513 (N_9513,N_8381,N_8723);
or U9514 (N_9514,N_8799,N_8279);
or U9515 (N_9515,N_8702,N_8664);
nor U9516 (N_9516,N_8878,N_8119);
nand U9517 (N_9517,N_8625,N_8992);
nand U9518 (N_9518,N_8007,N_8887);
nand U9519 (N_9519,N_8428,N_8060);
nand U9520 (N_9520,N_8959,N_8195);
nand U9521 (N_9521,N_8889,N_8857);
and U9522 (N_9522,N_8157,N_8129);
nand U9523 (N_9523,N_8223,N_8196);
xor U9524 (N_9524,N_8559,N_8455);
xor U9525 (N_9525,N_8799,N_8012);
nand U9526 (N_9526,N_8031,N_8254);
nor U9527 (N_9527,N_8213,N_8116);
nand U9528 (N_9528,N_8415,N_8920);
or U9529 (N_9529,N_8016,N_8167);
or U9530 (N_9530,N_8626,N_8269);
nand U9531 (N_9531,N_8801,N_8917);
xnor U9532 (N_9532,N_8309,N_8492);
nand U9533 (N_9533,N_8976,N_8624);
and U9534 (N_9534,N_8583,N_8445);
nand U9535 (N_9535,N_8061,N_8876);
and U9536 (N_9536,N_8357,N_8066);
nand U9537 (N_9537,N_8182,N_8670);
nand U9538 (N_9538,N_8972,N_8058);
or U9539 (N_9539,N_8815,N_8677);
nor U9540 (N_9540,N_8029,N_8761);
nand U9541 (N_9541,N_8382,N_8417);
and U9542 (N_9542,N_8237,N_8917);
or U9543 (N_9543,N_8577,N_8300);
and U9544 (N_9544,N_8979,N_8629);
nand U9545 (N_9545,N_8060,N_8679);
or U9546 (N_9546,N_8201,N_8444);
xnor U9547 (N_9547,N_8605,N_8701);
nand U9548 (N_9548,N_8746,N_8344);
or U9549 (N_9549,N_8060,N_8534);
and U9550 (N_9550,N_8846,N_8172);
or U9551 (N_9551,N_8559,N_8258);
nor U9552 (N_9552,N_8803,N_8827);
nor U9553 (N_9553,N_8103,N_8474);
nor U9554 (N_9554,N_8579,N_8669);
nor U9555 (N_9555,N_8144,N_8469);
or U9556 (N_9556,N_8895,N_8748);
and U9557 (N_9557,N_8929,N_8596);
nor U9558 (N_9558,N_8334,N_8957);
or U9559 (N_9559,N_8814,N_8973);
or U9560 (N_9560,N_8342,N_8445);
nand U9561 (N_9561,N_8528,N_8040);
and U9562 (N_9562,N_8535,N_8176);
xnor U9563 (N_9563,N_8886,N_8199);
and U9564 (N_9564,N_8621,N_8076);
xor U9565 (N_9565,N_8824,N_8883);
nor U9566 (N_9566,N_8594,N_8320);
nor U9567 (N_9567,N_8963,N_8660);
or U9568 (N_9568,N_8317,N_8156);
nand U9569 (N_9569,N_8699,N_8922);
xor U9570 (N_9570,N_8280,N_8261);
xor U9571 (N_9571,N_8274,N_8347);
or U9572 (N_9572,N_8426,N_8984);
or U9573 (N_9573,N_8438,N_8992);
nand U9574 (N_9574,N_8488,N_8791);
nor U9575 (N_9575,N_8959,N_8567);
nor U9576 (N_9576,N_8099,N_8174);
nand U9577 (N_9577,N_8127,N_8144);
or U9578 (N_9578,N_8268,N_8094);
nor U9579 (N_9579,N_8012,N_8994);
xor U9580 (N_9580,N_8077,N_8528);
xor U9581 (N_9581,N_8734,N_8864);
nor U9582 (N_9582,N_8330,N_8862);
nor U9583 (N_9583,N_8849,N_8421);
nand U9584 (N_9584,N_8279,N_8419);
and U9585 (N_9585,N_8798,N_8191);
xnor U9586 (N_9586,N_8173,N_8316);
nand U9587 (N_9587,N_8673,N_8305);
nor U9588 (N_9588,N_8418,N_8325);
nor U9589 (N_9589,N_8038,N_8294);
nor U9590 (N_9590,N_8130,N_8175);
or U9591 (N_9591,N_8663,N_8744);
xnor U9592 (N_9592,N_8667,N_8551);
nor U9593 (N_9593,N_8118,N_8077);
or U9594 (N_9594,N_8649,N_8189);
or U9595 (N_9595,N_8358,N_8027);
and U9596 (N_9596,N_8649,N_8819);
xnor U9597 (N_9597,N_8899,N_8898);
and U9598 (N_9598,N_8723,N_8662);
xor U9599 (N_9599,N_8898,N_8756);
nand U9600 (N_9600,N_8875,N_8289);
and U9601 (N_9601,N_8132,N_8430);
and U9602 (N_9602,N_8212,N_8546);
or U9603 (N_9603,N_8411,N_8194);
xnor U9604 (N_9604,N_8839,N_8024);
nor U9605 (N_9605,N_8859,N_8267);
xnor U9606 (N_9606,N_8536,N_8512);
nand U9607 (N_9607,N_8853,N_8838);
or U9608 (N_9608,N_8407,N_8262);
and U9609 (N_9609,N_8005,N_8038);
and U9610 (N_9610,N_8719,N_8402);
and U9611 (N_9611,N_8284,N_8549);
nand U9612 (N_9612,N_8045,N_8258);
and U9613 (N_9613,N_8783,N_8563);
and U9614 (N_9614,N_8728,N_8801);
and U9615 (N_9615,N_8628,N_8145);
nor U9616 (N_9616,N_8593,N_8212);
nand U9617 (N_9617,N_8062,N_8574);
xnor U9618 (N_9618,N_8876,N_8308);
nor U9619 (N_9619,N_8533,N_8037);
or U9620 (N_9620,N_8000,N_8047);
or U9621 (N_9621,N_8300,N_8731);
or U9622 (N_9622,N_8249,N_8386);
nand U9623 (N_9623,N_8212,N_8613);
xor U9624 (N_9624,N_8757,N_8850);
xnor U9625 (N_9625,N_8294,N_8407);
nand U9626 (N_9626,N_8239,N_8966);
or U9627 (N_9627,N_8751,N_8976);
nand U9628 (N_9628,N_8072,N_8146);
nor U9629 (N_9629,N_8178,N_8875);
and U9630 (N_9630,N_8834,N_8777);
or U9631 (N_9631,N_8572,N_8911);
and U9632 (N_9632,N_8770,N_8467);
nor U9633 (N_9633,N_8679,N_8097);
xor U9634 (N_9634,N_8545,N_8648);
nand U9635 (N_9635,N_8632,N_8407);
nand U9636 (N_9636,N_8102,N_8600);
xnor U9637 (N_9637,N_8981,N_8423);
nand U9638 (N_9638,N_8278,N_8019);
and U9639 (N_9639,N_8000,N_8435);
nand U9640 (N_9640,N_8394,N_8256);
nor U9641 (N_9641,N_8726,N_8620);
and U9642 (N_9642,N_8220,N_8011);
or U9643 (N_9643,N_8523,N_8020);
nand U9644 (N_9644,N_8822,N_8589);
nand U9645 (N_9645,N_8407,N_8383);
nor U9646 (N_9646,N_8589,N_8476);
xor U9647 (N_9647,N_8541,N_8172);
nand U9648 (N_9648,N_8279,N_8935);
nor U9649 (N_9649,N_8097,N_8588);
or U9650 (N_9650,N_8664,N_8198);
or U9651 (N_9651,N_8084,N_8330);
nor U9652 (N_9652,N_8363,N_8356);
xnor U9653 (N_9653,N_8827,N_8269);
xnor U9654 (N_9654,N_8608,N_8569);
or U9655 (N_9655,N_8346,N_8216);
and U9656 (N_9656,N_8607,N_8512);
nor U9657 (N_9657,N_8984,N_8756);
xnor U9658 (N_9658,N_8831,N_8253);
nor U9659 (N_9659,N_8807,N_8445);
xnor U9660 (N_9660,N_8246,N_8673);
and U9661 (N_9661,N_8476,N_8620);
and U9662 (N_9662,N_8791,N_8523);
nor U9663 (N_9663,N_8140,N_8982);
nor U9664 (N_9664,N_8827,N_8457);
nor U9665 (N_9665,N_8082,N_8923);
or U9666 (N_9666,N_8942,N_8268);
xor U9667 (N_9667,N_8490,N_8495);
nand U9668 (N_9668,N_8806,N_8296);
nand U9669 (N_9669,N_8607,N_8271);
nand U9670 (N_9670,N_8909,N_8879);
nand U9671 (N_9671,N_8662,N_8186);
or U9672 (N_9672,N_8151,N_8192);
nor U9673 (N_9673,N_8183,N_8698);
nor U9674 (N_9674,N_8448,N_8581);
and U9675 (N_9675,N_8795,N_8430);
and U9676 (N_9676,N_8007,N_8148);
nand U9677 (N_9677,N_8242,N_8129);
or U9678 (N_9678,N_8278,N_8220);
nand U9679 (N_9679,N_8284,N_8917);
nor U9680 (N_9680,N_8608,N_8741);
or U9681 (N_9681,N_8940,N_8390);
xnor U9682 (N_9682,N_8337,N_8473);
xor U9683 (N_9683,N_8039,N_8064);
nand U9684 (N_9684,N_8219,N_8623);
or U9685 (N_9685,N_8469,N_8895);
and U9686 (N_9686,N_8387,N_8506);
nor U9687 (N_9687,N_8520,N_8326);
or U9688 (N_9688,N_8091,N_8616);
or U9689 (N_9689,N_8352,N_8164);
nand U9690 (N_9690,N_8035,N_8414);
nand U9691 (N_9691,N_8607,N_8084);
or U9692 (N_9692,N_8987,N_8752);
nand U9693 (N_9693,N_8546,N_8771);
xor U9694 (N_9694,N_8290,N_8889);
nand U9695 (N_9695,N_8968,N_8108);
xnor U9696 (N_9696,N_8317,N_8131);
and U9697 (N_9697,N_8219,N_8339);
or U9698 (N_9698,N_8305,N_8459);
nor U9699 (N_9699,N_8557,N_8908);
nor U9700 (N_9700,N_8443,N_8736);
or U9701 (N_9701,N_8995,N_8146);
nand U9702 (N_9702,N_8424,N_8425);
nor U9703 (N_9703,N_8947,N_8479);
and U9704 (N_9704,N_8464,N_8690);
or U9705 (N_9705,N_8971,N_8633);
nor U9706 (N_9706,N_8479,N_8302);
nand U9707 (N_9707,N_8065,N_8545);
xor U9708 (N_9708,N_8401,N_8088);
nor U9709 (N_9709,N_8820,N_8418);
or U9710 (N_9710,N_8251,N_8116);
xor U9711 (N_9711,N_8432,N_8245);
xnor U9712 (N_9712,N_8198,N_8492);
and U9713 (N_9713,N_8364,N_8021);
or U9714 (N_9714,N_8494,N_8202);
nand U9715 (N_9715,N_8659,N_8073);
xor U9716 (N_9716,N_8791,N_8069);
or U9717 (N_9717,N_8997,N_8035);
and U9718 (N_9718,N_8706,N_8132);
and U9719 (N_9719,N_8769,N_8130);
or U9720 (N_9720,N_8185,N_8478);
and U9721 (N_9721,N_8851,N_8181);
xnor U9722 (N_9722,N_8185,N_8573);
or U9723 (N_9723,N_8996,N_8618);
and U9724 (N_9724,N_8705,N_8082);
or U9725 (N_9725,N_8694,N_8500);
nand U9726 (N_9726,N_8805,N_8328);
or U9727 (N_9727,N_8833,N_8480);
or U9728 (N_9728,N_8051,N_8769);
and U9729 (N_9729,N_8218,N_8465);
nand U9730 (N_9730,N_8828,N_8063);
nand U9731 (N_9731,N_8080,N_8768);
xor U9732 (N_9732,N_8264,N_8430);
nand U9733 (N_9733,N_8068,N_8413);
xor U9734 (N_9734,N_8152,N_8763);
and U9735 (N_9735,N_8879,N_8087);
or U9736 (N_9736,N_8408,N_8205);
nor U9737 (N_9737,N_8550,N_8999);
and U9738 (N_9738,N_8865,N_8673);
nor U9739 (N_9739,N_8114,N_8189);
nand U9740 (N_9740,N_8484,N_8130);
nand U9741 (N_9741,N_8629,N_8611);
xor U9742 (N_9742,N_8945,N_8559);
nor U9743 (N_9743,N_8270,N_8162);
or U9744 (N_9744,N_8640,N_8215);
nand U9745 (N_9745,N_8698,N_8731);
or U9746 (N_9746,N_8330,N_8110);
and U9747 (N_9747,N_8127,N_8381);
nor U9748 (N_9748,N_8868,N_8295);
nand U9749 (N_9749,N_8613,N_8539);
or U9750 (N_9750,N_8721,N_8610);
and U9751 (N_9751,N_8555,N_8549);
nor U9752 (N_9752,N_8670,N_8916);
nand U9753 (N_9753,N_8032,N_8008);
and U9754 (N_9754,N_8104,N_8671);
nand U9755 (N_9755,N_8478,N_8369);
nor U9756 (N_9756,N_8408,N_8927);
nor U9757 (N_9757,N_8545,N_8689);
and U9758 (N_9758,N_8942,N_8861);
nand U9759 (N_9759,N_8183,N_8256);
and U9760 (N_9760,N_8144,N_8266);
nor U9761 (N_9761,N_8840,N_8798);
and U9762 (N_9762,N_8820,N_8673);
xor U9763 (N_9763,N_8400,N_8748);
xor U9764 (N_9764,N_8389,N_8303);
or U9765 (N_9765,N_8072,N_8107);
nand U9766 (N_9766,N_8536,N_8911);
nor U9767 (N_9767,N_8855,N_8598);
or U9768 (N_9768,N_8169,N_8995);
nor U9769 (N_9769,N_8594,N_8060);
xnor U9770 (N_9770,N_8307,N_8589);
or U9771 (N_9771,N_8884,N_8478);
or U9772 (N_9772,N_8771,N_8999);
nor U9773 (N_9773,N_8248,N_8896);
and U9774 (N_9774,N_8452,N_8312);
and U9775 (N_9775,N_8302,N_8576);
and U9776 (N_9776,N_8763,N_8148);
and U9777 (N_9777,N_8757,N_8756);
xnor U9778 (N_9778,N_8565,N_8415);
xnor U9779 (N_9779,N_8150,N_8584);
xnor U9780 (N_9780,N_8068,N_8019);
nor U9781 (N_9781,N_8245,N_8072);
xnor U9782 (N_9782,N_8517,N_8684);
xnor U9783 (N_9783,N_8780,N_8672);
nand U9784 (N_9784,N_8826,N_8266);
nor U9785 (N_9785,N_8744,N_8982);
or U9786 (N_9786,N_8923,N_8250);
and U9787 (N_9787,N_8309,N_8124);
nor U9788 (N_9788,N_8862,N_8109);
nor U9789 (N_9789,N_8122,N_8276);
or U9790 (N_9790,N_8884,N_8412);
and U9791 (N_9791,N_8271,N_8425);
and U9792 (N_9792,N_8697,N_8853);
nor U9793 (N_9793,N_8356,N_8291);
xnor U9794 (N_9794,N_8716,N_8529);
xnor U9795 (N_9795,N_8004,N_8528);
nand U9796 (N_9796,N_8731,N_8900);
xor U9797 (N_9797,N_8986,N_8042);
xnor U9798 (N_9798,N_8026,N_8497);
or U9799 (N_9799,N_8906,N_8797);
and U9800 (N_9800,N_8616,N_8918);
and U9801 (N_9801,N_8235,N_8034);
nor U9802 (N_9802,N_8539,N_8831);
and U9803 (N_9803,N_8217,N_8177);
or U9804 (N_9804,N_8309,N_8452);
nor U9805 (N_9805,N_8509,N_8161);
and U9806 (N_9806,N_8834,N_8408);
nand U9807 (N_9807,N_8791,N_8411);
and U9808 (N_9808,N_8010,N_8664);
nor U9809 (N_9809,N_8646,N_8625);
nand U9810 (N_9810,N_8949,N_8774);
or U9811 (N_9811,N_8518,N_8414);
or U9812 (N_9812,N_8432,N_8406);
xor U9813 (N_9813,N_8901,N_8070);
and U9814 (N_9814,N_8201,N_8835);
nor U9815 (N_9815,N_8997,N_8226);
or U9816 (N_9816,N_8893,N_8718);
and U9817 (N_9817,N_8551,N_8425);
or U9818 (N_9818,N_8126,N_8084);
and U9819 (N_9819,N_8378,N_8203);
nand U9820 (N_9820,N_8557,N_8124);
nor U9821 (N_9821,N_8592,N_8478);
xor U9822 (N_9822,N_8115,N_8012);
or U9823 (N_9823,N_8471,N_8763);
nor U9824 (N_9824,N_8527,N_8963);
or U9825 (N_9825,N_8840,N_8856);
nand U9826 (N_9826,N_8396,N_8614);
and U9827 (N_9827,N_8099,N_8645);
nor U9828 (N_9828,N_8819,N_8915);
xnor U9829 (N_9829,N_8954,N_8983);
nor U9830 (N_9830,N_8365,N_8043);
or U9831 (N_9831,N_8955,N_8415);
nand U9832 (N_9832,N_8793,N_8029);
xnor U9833 (N_9833,N_8096,N_8907);
nand U9834 (N_9834,N_8938,N_8963);
or U9835 (N_9835,N_8740,N_8636);
or U9836 (N_9836,N_8237,N_8404);
nand U9837 (N_9837,N_8750,N_8588);
xor U9838 (N_9838,N_8995,N_8221);
nor U9839 (N_9839,N_8017,N_8634);
and U9840 (N_9840,N_8171,N_8968);
nor U9841 (N_9841,N_8417,N_8771);
and U9842 (N_9842,N_8464,N_8207);
nand U9843 (N_9843,N_8586,N_8454);
or U9844 (N_9844,N_8663,N_8955);
xnor U9845 (N_9845,N_8282,N_8608);
nand U9846 (N_9846,N_8856,N_8071);
and U9847 (N_9847,N_8179,N_8235);
nand U9848 (N_9848,N_8291,N_8110);
nand U9849 (N_9849,N_8219,N_8513);
nor U9850 (N_9850,N_8128,N_8896);
or U9851 (N_9851,N_8502,N_8064);
and U9852 (N_9852,N_8268,N_8324);
nand U9853 (N_9853,N_8521,N_8301);
nor U9854 (N_9854,N_8921,N_8651);
nor U9855 (N_9855,N_8598,N_8773);
nand U9856 (N_9856,N_8821,N_8626);
nand U9857 (N_9857,N_8419,N_8743);
nor U9858 (N_9858,N_8803,N_8598);
xor U9859 (N_9859,N_8884,N_8808);
or U9860 (N_9860,N_8065,N_8676);
or U9861 (N_9861,N_8627,N_8007);
nor U9862 (N_9862,N_8993,N_8765);
and U9863 (N_9863,N_8276,N_8639);
nand U9864 (N_9864,N_8409,N_8202);
nor U9865 (N_9865,N_8981,N_8155);
or U9866 (N_9866,N_8853,N_8911);
or U9867 (N_9867,N_8802,N_8038);
and U9868 (N_9868,N_8642,N_8215);
nor U9869 (N_9869,N_8801,N_8103);
nand U9870 (N_9870,N_8307,N_8146);
nand U9871 (N_9871,N_8105,N_8229);
xor U9872 (N_9872,N_8602,N_8247);
and U9873 (N_9873,N_8074,N_8797);
and U9874 (N_9874,N_8957,N_8285);
nand U9875 (N_9875,N_8918,N_8931);
nor U9876 (N_9876,N_8590,N_8683);
and U9877 (N_9877,N_8390,N_8500);
and U9878 (N_9878,N_8391,N_8419);
xnor U9879 (N_9879,N_8431,N_8681);
and U9880 (N_9880,N_8757,N_8146);
nand U9881 (N_9881,N_8545,N_8718);
or U9882 (N_9882,N_8860,N_8389);
nand U9883 (N_9883,N_8418,N_8433);
nor U9884 (N_9884,N_8405,N_8088);
nand U9885 (N_9885,N_8389,N_8428);
xnor U9886 (N_9886,N_8788,N_8512);
xor U9887 (N_9887,N_8284,N_8827);
nor U9888 (N_9888,N_8484,N_8687);
nor U9889 (N_9889,N_8030,N_8065);
and U9890 (N_9890,N_8082,N_8842);
and U9891 (N_9891,N_8101,N_8854);
or U9892 (N_9892,N_8035,N_8037);
xnor U9893 (N_9893,N_8396,N_8399);
xnor U9894 (N_9894,N_8232,N_8384);
nor U9895 (N_9895,N_8728,N_8511);
nand U9896 (N_9896,N_8449,N_8261);
nand U9897 (N_9897,N_8173,N_8635);
and U9898 (N_9898,N_8550,N_8661);
xor U9899 (N_9899,N_8564,N_8267);
nor U9900 (N_9900,N_8992,N_8528);
or U9901 (N_9901,N_8289,N_8228);
xnor U9902 (N_9902,N_8561,N_8349);
nor U9903 (N_9903,N_8718,N_8475);
nand U9904 (N_9904,N_8427,N_8671);
xnor U9905 (N_9905,N_8434,N_8217);
nor U9906 (N_9906,N_8844,N_8518);
and U9907 (N_9907,N_8081,N_8116);
nand U9908 (N_9908,N_8342,N_8613);
nand U9909 (N_9909,N_8355,N_8865);
or U9910 (N_9910,N_8110,N_8531);
nor U9911 (N_9911,N_8976,N_8049);
nor U9912 (N_9912,N_8262,N_8132);
and U9913 (N_9913,N_8115,N_8352);
and U9914 (N_9914,N_8579,N_8778);
nand U9915 (N_9915,N_8872,N_8993);
xnor U9916 (N_9916,N_8751,N_8372);
nor U9917 (N_9917,N_8676,N_8551);
nand U9918 (N_9918,N_8051,N_8818);
nor U9919 (N_9919,N_8298,N_8171);
nor U9920 (N_9920,N_8954,N_8093);
or U9921 (N_9921,N_8667,N_8103);
xor U9922 (N_9922,N_8047,N_8093);
or U9923 (N_9923,N_8384,N_8899);
or U9924 (N_9924,N_8427,N_8499);
and U9925 (N_9925,N_8098,N_8631);
nand U9926 (N_9926,N_8114,N_8428);
or U9927 (N_9927,N_8110,N_8256);
nor U9928 (N_9928,N_8762,N_8214);
xor U9929 (N_9929,N_8212,N_8076);
or U9930 (N_9930,N_8934,N_8693);
xor U9931 (N_9931,N_8503,N_8622);
nor U9932 (N_9932,N_8502,N_8368);
or U9933 (N_9933,N_8034,N_8105);
nand U9934 (N_9934,N_8809,N_8675);
xnor U9935 (N_9935,N_8109,N_8894);
xnor U9936 (N_9936,N_8981,N_8909);
xnor U9937 (N_9937,N_8159,N_8463);
nand U9938 (N_9938,N_8632,N_8571);
and U9939 (N_9939,N_8061,N_8645);
nand U9940 (N_9940,N_8095,N_8411);
nand U9941 (N_9941,N_8522,N_8476);
xor U9942 (N_9942,N_8123,N_8127);
or U9943 (N_9943,N_8587,N_8913);
or U9944 (N_9944,N_8005,N_8237);
xor U9945 (N_9945,N_8399,N_8477);
or U9946 (N_9946,N_8211,N_8601);
nor U9947 (N_9947,N_8649,N_8883);
xnor U9948 (N_9948,N_8501,N_8544);
nor U9949 (N_9949,N_8492,N_8349);
nor U9950 (N_9950,N_8632,N_8869);
nand U9951 (N_9951,N_8487,N_8175);
nor U9952 (N_9952,N_8257,N_8631);
nand U9953 (N_9953,N_8102,N_8711);
or U9954 (N_9954,N_8989,N_8649);
xor U9955 (N_9955,N_8446,N_8225);
nor U9956 (N_9956,N_8076,N_8280);
nand U9957 (N_9957,N_8855,N_8379);
or U9958 (N_9958,N_8778,N_8455);
or U9959 (N_9959,N_8223,N_8526);
xnor U9960 (N_9960,N_8874,N_8475);
nor U9961 (N_9961,N_8000,N_8579);
nor U9962 (N_9962,N_8145,N_8988);
or U9963 (N_9963,N_8427,N_8868);
or U9964 (N_9964,N_8489,N_8000);
nand U9965 (N_9965,N_8303,N_8272);
xor U9966 (N_9966,N_8026,N_8191);
or U9967 (N_9967,N_8116,N_8073);
nor U9968 (N_9968,N_8091,N_8630);
xor U9969 (N_9969,N_8113,N_8188);
nor U9970 (N_9970,N_8429,N_8438);
nor U9971 (N_9971,N_8197,N_8983);
and U9972 (N_9972,N_8733,N_8156);
or U9973 (N_9973,N_8024,N_8481);
and U9974 (N_9974,N_8741,N_8442);
or U9975 (N_9975,N_8837,N_8445);
nor U9976 (N_9976,N_8204,N_8845);
nor U9977 (N_9977,N_8875,N_8967);
nor U9978 (N_9978,N_8369,N_8458);
nand U9979 (N_9979,N_8895,N_8650);
nand U9980 (N_9980,N_8527,N_8279);
and U9981 (N_9981,N_8572,N_8426);
xor U9982 (N_9982,N_8157,N_8133);
and U9983 (N_9983,N_8019,N_8292);
or U9984 (N_9984,N_8471,N_8424);
and U9985 (N_9985,N_8164,N_8152);
or U9986 (N_9986,N_8474,N_8714);
xnor U9987 (N_9987,N_8778,N_8543);
xnor U9988 (N_9988,N_8967,N_8047);
xor U9989 (N_9989,N_8962,N_8633);
xor U9990 (N_9990,N_8033,N_8529);
nand U9991 (N_9991,N_8633,N_8592);
nor U9992 (N_9992,N_8580,N_8190);
nand U9993 (N_9993,N_8562,N_8209);
nor U9994 (N_9994,N_8750,N_8890);
nand U9995 (N_9995,N_8544,N_8847);
nor U9996 (N_9996,N_8895,N_8435);
nor U9997 (N_9997,N_8187,N_8563);
nand U9998 (N_9998,N_8257,N_8518);
nor U9999 (N_9999,N_8033,N_8706);
nor U10000 (N_10000,N_9955,N_9645);
nand U10001 (N_10001,N_9095,N_9952);
xor U10002 (N_10002,N_9533,N_9627);
or U10003 (N_10003,N_9144,N_9240);
xnor U10004 (N_10004,N_9807,N_9739);
or U10005 (N_10005,N_9719,N_9972);
nor U10006 (N_10006,N_9389,N_9520);
nand U10007 (N_10007,N_9163,N_9990);
or U10008 (N_10008,N_9505,N_9850);
nand U10009 (N_10009,N_9040,N_9843);
or U10010 (N_10010,N_9672,N_9416);
nor U10011 (N_10011,N_9727,N_9072);
and U10012 (N_10012,N_9999,N_9029);
and U10013 (N_10013,N_9272,N_9610);
xor U10014 (N_10014,N_9615,N_9816);
nand U10015 (N_10015,N_9134,N_9530);
xnor U10016 (N_10016,N_9124,N_9766);
or U10017 (N_10017,N_9537,N_9074);
nand U10018 (N_10018,N_9171,N_9662);
nor U10019 (N_10019,N_9818,N_9049);
xor U10020 (N_10020,N_9892,N_9617);
xnor U10021 (N_10021,N_9552,N_9265);
xnor U10022 (N_10022,N_9569,N_9117);
nand U10023 (N_10023,N_9464,N_9126);
nand U10024 (N_10024,N_9623,N_9877);
or U10025 (N_10025,N_9934,N_9957);
and U10026 (N_10026,N_9798,N_9660);
nand U10027 (N_10027,N_9279,N_9979);
nor U10028 (N_10028,N_9842,N_9891);
nand U10029 (N_10029,N_9304,N_9907);
xnor U10030 (N_10030,N_9933,N_9069);
nand U10031 (N_10031,N_9702,N_9806);
nor U10032 (N_10032,N_9027,N_9313);
xnor U10033 (N_10033,N_9954,N_9000);
xnor U10034 (N_10034,N_9102,N_9001);
nor U10035 (N_10035,N_9162,N_9371);
xor U10036 (N_10036,N_9889,N_9318);
xor U10037 (N_10037,N_9961,N_9646);
nand U10038 (N_10038,N_9918,N_9708);
nand U10039 (N_10039,N_9786,N_9777);
nand U10040 (N_10040,N_9032,N_9688);
or U10041 (N_10041,N_9607,N_9622);
and U10042 (N_10042,N_9586,N_9120);
and U10043 (N_10043,N_9384,N_9060);
nand U10044 (N_10044,N_9975,N_9055);
and U10045 (N_10045,N_9742,N_9613);
nor U10046 (N_10046,N_9061,N_9020);
and U10047 (N_10047,N_9355,N_9704);
or U10048 (N_10048,N_9349,N_9902);
nand U10049 (N_10049,N_9939,N_9148);
xor U10050 (N_10050,N_9222,N_9916);
xor U10051 (N_10051,N_9506,N_9044);
and U10052 (N_10052,N_9486,N_9502);
and U10053 (N_10053,N_9085,N_9017);
xnor U10054 (N_10054,N_9577,N_9861);
nand U10055 (N_10055,N_9251,N_9185);
or U10056 (N_10056,N_9181,N_9387);
xnor U10057 (N_10057,N_9446,N_9465);
or U10058 (N_10058,N_9811,N_9199);
and U10059 (N_10059,N_9320,N_9532);
xor U10060 (N_10060,N_9686,N_9024);
nand U10061 (N_10061,N_9982,N_9542);
xor U10062 (N_10062,N_9278,N_9734);
nand U10063 (N_10063,N_9255,N_9913);
xnor U10064 (N_10064,N_9353,N_9883);
xnor U10065 (N_10065,N_9504,N_9854);
xnor U10066 (N_10066,N_9395,N_9637);
nand U10067 (N_10067,N_9523,N_9980);
and U10068 (N_10068,N_9959,N_9812);
nor U10069 (N_10069,N_9308,N_9492);
nand U10070 (N_10070,N_9815,N_9721);
nor U10071 (N_10071,N_9300,N_9706);
nor U10072 (N_10072,N_9795,N_9946);
nand U10073 (N_10073,N_9476,N_9670);
xor U10074 (N_10074,N_9083,N_9213);
or U10075 (N_10075,N_9346,N_9516);
nand U10076 (N_10076,N_9399,N_9664);
or U10077 (N_10077,N_9249,N_9335);
nor U10078 (N_10078,N_9796,N_9316);
nand U10079 (N_10079,N_9819,N_9543);
nor U10080 (N_10080,N_9137,N_9746);
xnor U10081 (N_10081,N_9431,N_9479);
or U10082 (N_10082,N_9657,N_9332);
or U10083 (N_10083,N_9451,N_9014);
and U10084 (N_10084,N_9432,N_9182);
nand U10085 (N_10085,N_9025,N_9472);
and U10086 (N_10086,N_9601,N_9123);
and U10087 (N_10087,N_9602,N_9944);
nand U10088 (N_10088,N_9781,N_9914);
and U10089 (N_10089,N_9857,N_9823);
and U10090 (N_10090,N_9666,N_9941);
or U10091 (N_10091,N_9453,N_9653);
and U10092 (N_10092,N_9831,N_9554);
nand U10093 (N_10093,N_9738,N_9636);
or U10094 (N_10094,N_9714,N_9274);
and U10095 (N_10095,N_9107,N_9398);
or U10096 (N_10096,N_9367,N_9896);
xor U10097 (N_10097,N_9940,N_9401);
and U10098 (N_10098,N_9986,N_9232);
and U10099 (N_10099,N_9234,N_9491);
nand U10100 (N_10100,N_9603,N_9226);
and U10101 (N_10101,N_9847,N_9976);
and U10102 (N_10102,N_9551,N_9498);
nor U10103 (N_10103,N_9503,N_9559);
nand U10104 (N_10104,N_9175,N_9204);
or U10105 (N_10105,N_9462,N_9494);
xor U10106 (N_10106,N_9632,N_9733);
nand U10107 (N_10107,N_9690,N_9236);
xor U10108 (N_10108,N_9325,N_9059);
xor U10109 (N_10109,N_9712,N_9583);
or U10110 (N_10110,N_9879,N_9418);
or U10111 (N_10111,N_9435,N_9848);
and U10112 (N_10112,N_9930,N_9103);
or U10113 (N_10113,N_9745,N_9997);
and U10114 (N_10114,N_9549,N_9403);
nand U10115 (N_10115,N_9114,N_9836);
xnor U10116 (N_10116,N_9339,N_9390);
nand U10117 (N_10117,N_9484,N_9150);
nand U10118 (N_10118,N_9826,N_9876);
or U10119 (N_10119,N_9077,N_9748);
nor U10120 (N_10120,N_9598,N_9866);
or U10121 (N_10121,N_9051,N_9856);
xor U10122 (N_10122,N_9419,N_9245);
or U10123 (N_10123,N_9197,N_9612);
nand U10124 (N_10124,N_9611,N_9352);
and U10125 (N_10125,N_9297,N_9840);
nor U10126 (N_10126,N_9334,N_9167);
nand U10127 (N_10127,N_9317,N_9264);
nand U10128 (N_10128,N_9604,N_9835);
nand U10129 (N_10129,N_9276,N_9450);
or U10130 (N_10130,N_9109,N_9832);
and U10131 (N_10131,N_9321,N_9887);
xor U10132 (N_10132,N_9932,N_9113);
or U10133 (N_10133,N_9562,N_9104);
nand U10134 (N_10134,N_9269,N_9271);
nor U10135 (N_10135,N_9100,N_9374);
nor U10136 (N_10136,N_9391,N_9629);
or U10137 (N_10137,N_9493,N_9337);
and U10138 (N_10138,N_9179,N_9046);
and U10139 (N_10139,N_9501,N_9436);
nand U10140 (N_10140,N_9684,N_9923);
xnor U10141 (N_10141,N_9071,N_9441);
nor U10142 (N_10142,N_9878,N_9732);
and U10143 (N_10143,N_9490,N_9289);
nand U10144 (N_10144,N_9153,N_9978);
and U10145 (N_10145,N_9749,N_9780);
nor U10146 (N_10146,N_9863,N_9205);
nor U10147 (N_10147,N_9016,N_9262);
nor U10148 (N_10148,N_9063,N_9691);
or U10149 (N_10149,N_9969,N_9368);
and U10150 (N_10150,N_9075,N_9377);
xnor U10151 (N_10151,N_9568,N_9217);
xnor U10152 (N_10152,N_9512,N_9483);
nand U10153 (N_10153,N_9964,N_9201);
nand U10154 (N_10154,N_9618,N_9594);
xnor U10155 (N_10155,N_9149,N_9814);
and U10156 (N_10156,N_9676,N_9008);
or U10157 (N_10157,N_9002,N_9853);
nand U10158 (N_10158,N_9965,N_9214);
nand U10159 (N_10159,N_9736,N_9301);
nand U10160 (N_10160,N_9310,N_9718);
or U10161 (N_10161,N_9424,N_9396);
nor U10162 (N_10162,N_9340,N_9038);
nand U10163 (N_10163,N_9026,N_9326);
xor U10164 (N_10164,N_9259,N_9903);
nand U10165 (N_10165,N_9078,N_9936);
or U10166 (N_10166,N_9915,N_9286);
xnor U10167 (N_10167,N_9130,N_9985);
or U10168 (N_10168,N_9942,N_9128);
nor U10169 (N_10169,N_9053,N_9388);
xnor U10170 (N_10170,N_9342,N_9101);
and U10171 (N_10171,N_9929,N_9871);
xor U10172 (N_10172,N_9164,N_9184);
or U10173 (N_10173,N_9140,N_9227);
or U10174 (N_10174,N_9680,N_9671);
xnor U10175 (N_10175,N_9679,N_9567);
xnor U10176 (N_10176,N_9018,N_9021);
xor U10177 (N_10177,N_9967,N_9689);
and U10178 (N_10178,N_9288,N_9455);
xor U10179 (N_10179,N_9073,N_9722);
nor U10180 (N_10180,N_9378,N_9663);
or U10181 (N_10181,N_9145,N_9463);
nand U10182 (N_10182,N_9302,N_9135);
nand U10183 (N_10183,N_9769,N_9729);
nor U10184 (N_10184,N_9634,N_9723);
nor U10185 (N_10185,N_9440,N_9365);
or U10186 (N_10186,N_9880,N_9009);
or U10187 (N_10187,N_9700,N_9758);
or U10188 (N_10188,N_9280,N_9136);
or U10189 (N_10189,N_9299,N_9086);
xor U10190 (N_10190,N_9229,N_9968);
nor U10191 (N_10191,N_9359,N_9513);
or U10192 (N_10192,N_9548,N_9587);
nand U10193 (N_10193,N_9413,N_9564);
xnor U10194 (N_10194,N_9652,N_9635);
or U10195 (N_10195,N_9709,N_9481);
nor U10196 (N_10196,N_9720,N_9508);
xor U10197 (N_10197,N_9905,N_9973);
xor U10198 (N_10198,N_9698,N_9138);
and U10199 (N_10199,N_9731,N_9995);
and U10200 (N_10200,N_9345,N_9425);
nand U10201 (N_10201,N_9058,N_9667);
and U10202 (N_10202,N_9458,N_9785);
nand U10203 (N_10203,N_9282,N_9035);
and U10204 (N_10204,N_9323,N_9560);
nand U10205 (N_10205,N_9146,N_9022);
xnor U10206 (N_10206,N_9216,N_9169);
nor U10207 (N_10207,N_9628,N_9687);
or U10208 (N_10208,N_9407,N_9141);
or U10209 (N_10209,N_9070,N_9890);
nand U10210 (N_10210,N_9574,N_9273);
nand U10211 (N_10211,N_9324,N_9090);
and U10212 (N_10212,N_9319,N_9166);
and U10213 (N_10213,N_9057,N_9015);
and U10214 (N_10214,N_9996,N_9593);
nor U10215 (N_10215,N_9752,N_9755);
xnor U10216 (N_10216,N_9747,N_9971);
nor U10217 (N_10217,N_9616,N_9091);
xnor U10218 (N_10218,N_9219,N_9127);
nand U10219 (N_10219,N_9949,N_9496);
xor U10220 (N_10220,N_9290,N_9098);
nor U10221 (N_10221,N_9168,N_9960);
xnor U10222 (N_10222,N_9697,N_9261);
xnor U10223 (N_10223,N_9488,N_9950);
nor U10224 (N_10224,N_9247,N_9094);
nand U10225 (N_10225,N_9336,N_9005);
or U10226 (N_10226,N_9047,N_9206);
nor U10227 (N_10227,N_9068,N_9155);
or U10228 (N_10228,N_9829,N_9683);
and U10229 (N_10229,N_9445,N_9845);
xor U10230 (N_10230,N_9953,N_9544);
nor U10231 (N_10231,N_9408,N_9354);
and U10232 (N_10232,N_9042,N_9237);
and U10233 (N_10233,N_9189,N_9202);
and U10234 (N_10234,N_9099,N_9443);
and U10235 (N_10235,N_9173,N_9703);
xnor U10236 (N_10236,N_9036,N_9284);
or U10237 (N_10237,N_9888,N_9421);
nor U10238 (N_10238,N_9322,N_9315);
nand U10239 (N_10239,N_9433,N_9281);
xor U10240 (N_10240,N_9793,N_9893);
or U10241 (N_10241,N_9248,N_9115);
nor U10242 (N_10242,N_9254,N_9935);
nor U10243 (N_10243,N_9619,N_9152);
and U10244 (N_10244,N_9386,N_9647);
and U10245 (N_10245,N_9531,N_9415);
and U10246 (N_10246,N_9655,N_9351);
or U10247 (N_10247,N_9019,N_9156);
nor U10248 (N_10248,N_9195,N_9790);
nand U10249 (N_10249,N_9442,N_9238);
or U10250 (N_10250,N_9350,N_9258);
and U10251 (N_10251,N_9011,N_9087);
and U10252 (N_10252,N_9224,N_9203);
nor U10253 (N_10253,N_9735,N_9989);
or U10254 (N_10254,N_9926,N_9599);
xor U10255 (N_10255,N_9792,N_9244);
and U10256 (N_10256,N_9595,N_9329);
nor U10257 (N_10257,N_9917,N_9469);
and U10258 (N_10258,N_9713,N_9707);
nand U10259 (N_10259,N_9454,N_9437);
xor U10260 (N_10260,N_9050,N_9715);
and U10261 (N_10261,N_9404,N_9885);
or U10262 (N_10262,N_9088,N_9775);
and U10263 (N_10263,N_9759,N_9539);
nor U10264 (N_10264,N_9535,N_9466);
nand U10265 (N_10265,N_9106,N_9639);
nor U10266 (N_10266,N_9056,N_9174);
nor U10267 (N_10267,N_9994,N_9439);
nand U10268 (N_10268,N_9827,N_9430);
or U10269 (N_10269,N_9522,N_9860);
nor U10270 (N_10270,N_9343,N_9682);
xnor U10271 (N_10271,N_9406,N_9865);
nor U10272 (N_10272,N_9624,N_9789);
or U10273 (N_10273,N_9631,N_9669);
nor U10274 (N_10274,N_9048,N_9509);
xnor U10275 (N_10275,N_9782,N_9212);
nor U10276 (N_10276,N_9331,N_9741);
nand U10277 (N_10277,N_9394,N_9724);
xor U10278 (N_10278,N_9383,N_9405);
or U10279 (N_10279,N_9154,N_9546);
and U10280 (N_10280,N_9253,N_9794);
xnor U10281 (N_10281,N_9716,N_9641);
nand U10282 (N_10282,N_9561,N_9218);
xor U10283 (N_10283,N_9750,N_9041);
xor U10284 (N_10284,N_9411,N_9366);
or U10285 (N_10285,N_9821,N_9473);
or U10286 (N_10286,N_9118,N_9638);
or U10287 (N_10287,N_9196,N_9423);
and U10288 (N_10288,N_9881,N_9012);
nor U10289 (N_10289,N_9580,N_9373);
nor U10290 (N_10290,N_9448,N_9525);
and U10291 (N_10291,N_9570,N_9572);
xor U10292 (N_10292,N_9305,N_9007);
nand U10293 (N_10293,N_9370,N_9283);
nand U10294 (N_10294,N_9685,N_9487);
and U10295 (N_10295,N_9897,N_9859);
nor U10296 (N_10296,N_9550,N_9030);
and U10297 (N_10297,N_9545,N_9194);
nand U10298 (N_10298,N_9527,N_9763);
xnor U10299 (N_10299,N_9906,N_9193);
and U10300 (N_10300,N_9563,N_9894);
and U10301 (N_10301,N_9043,N_9787);
xnor U10302 (N_10302,N_9882,N_9221);
xor U10303 (N_10303,N_9605,N_9161);
nand U10304 (N_10304,N_9924,N_9737);
nand U10305 (N_10305,N_9591,N_9470);
and U10306 (N_10306,N_9110,N_9757);
nand U10307 (N_10307,N_9648,N_9298);
and U10308 (N_10308,N_9803,N_9770);
xnor U10309 (N_10309,N_9922,N_9402);
or U10310 (N_10310,N_9067,N_9344);
and U10311 (N_10311,N_9079,N_9357);
xor U10312 (N_10312,N_9963,N_9369);
nor U10313 (N_10313,N_9825,N_9267);
or U10314 (N_10314,N_9133,N_9725);
xnor U10315 (N_10315,N_9293,N_9180);
nand U10316 (N_10316,N_9519,N_9447);
xor U10317 (N_10317,N_9081,N_9275);
nor U10318 (N_10318,N_9231,N_9006);
nor U10319 (N_10319,N_9867,N_9987);
nand U10320 (N_10320,N_9830,N_9837);
xnor U10321 (N_10321,N_9330,N_9207);
or U10322 (N_10322,N_9565,N_9291);
xnor U10323 (N_10323,N_9263,N_9951);
and U10324 (N_10324,N_9529,N_9250);
nor U10325 (N_10325,N_9921,N_9460);
and U10326 (N_10326,N_9270,N_9928);
or U10327 (N_10327,N_9268,N_9361);
nand U10328 (N_10328,N_9003,N_9870);
or U10329 (N_10329,N_9467,N_9696);
nand U10330 (N_10330,N_9191,N_9555);
or U10331 (N_10331,N_9558,N_9356);
nand U10332 (N_10332,N_9328,N_9147);
xnor U10333 (N_10333,N_9158,N_9675);
and U10334 (N_10334,N_9129,N_9111);
nor U10335 (N_10335,N_9364,N_9991);
nand U10336 (N_10336,N_9710,N_9277);
and U10337 (N_10337,N_9287,N_9459);
and U10338 (N_10338,N_9242,N_9434);
and U10339 (N_10339,N_9241,N_9105);
and U10340 (N_10340,N_9170,N_9693);
and U10341 (N_10341,N_9589,N_9210);
and U10342 (N_10342,N_9309,N_9651);
xor U10343 (N_10343,N_9478,N_9644);
nor U10344 (N_10344,N_9065,N_9977);
nor U10345 (N_10345,N_9223,N_9515);
nor U10346 (N_10346,N_9575,N_9838);
and U10347 (N_10347,N_9116,N_9849);
nand U10348 (N_10348,N_9510,N_9076);
xnor U10349 (N_10349,N_9937,N_9983);
nand U10350 (N_10350,N_9761,N_9521);
and U10351 (N_10351,N_9919,N_9358);
nor U10352 (N_10352,N_9314,N_9547);
nor U10353 (N_10353,N_9159,N_9142);
nor U10354 (N_10354,N_9382,N_9868);
xnor U10355 (N_10355,N_9341,N_9186);
and U10356 (N_10356,N_9165,N_9380);
xnor U10357 (N_10357,N_9412,N_9220);
or U10358 (N_10358,N_9958,N_9661);
nor U10359 (N_10359,N_9809,N_9066);
or U10360 (N_10360,N_9855,N_9235);
nor U10361 (N_10361,N_9157,N_9536);
or U10362 (N_10362,N_9600,N_9872);
and U10363 (N_10363,N_9779,N_9379);
nand U10364 (N_10364,N_9208,N_9228);
xor U10365 (N_10365,N_9797,N_9846);
or U10366 (N_10366,N_9311,N_9064);
nand U10367 (N_10367,N_9392,N_9172);
nand U10368 (N_10368,N_9132,N_9970);
xnor U10369 (N_10369,N_9654,N_9517);
and U10370 (N_10370,N_9783,N_9895);
nand U10371 (N_10371,N_9744,N_9471);
or U10372 (N_10372,N_9642,N_9851);
nand U10373 (N_10373,N_9678,N_9904);
nor U10374 (N_10374,N_9673,N_9187);
xor U10375 (N_10375,N_9820,N_9338);
or U10376 (N_10376,N_9920,N_9625);
and U10377 (N_10377,N_9397,N_9348);
and U10378 (N_10378,N_9938,N_9312);
nand U10379 (N_10379,N_9160,N_9768);
and U10380 (N_10380,N_9692,N_9092);
nor U10381 (N_10381,N_9898,N_9514);
nor U10382 (N_10382,N_9592,N_9584);
nor U10383 (N_10383,N_9489,N_9717);
and U10384 (N_10384,N_9844,N_9534);
or U10385 (N_10385,N_9966,N_9381);
xor U10386 (N_10386,N_9659,N_9511);
nor U10387 (N_10387,N_9256,N_9909);
xnor U10388 (N_10388,N_9699,N_9762);
nand U10389 (N_10389,N_9385,N_9215);
nand U10390 (N_10390,N_9993,N_9557);
and U10391 (N_10391,N_9760,N_9927);
and U10392 (N_10392,N_9556,N_9767);
or U10393 (N_10393,N_9908,N_9200);
nand U10394 (N_10394,N_9571,N_9774);
or U10395 (N_10395,N_9778,N_9566);
xnor U10396 (N_10396,N_9576,N_9925);
xor U10397 (N_10397,N_9884,N_9608);
or U10398 (N_10398,N_9956,N_9139);
nand U10399 (N_10399,N_9307,N_9198);
xor U10400 (N_10400,N_9694,N_9773);
and U10401 (N_10401,N_9711,N_9728);
or U10402 (N_10402,N_9784,N_9943);
xor U10403 (N_10403,N_9410,N_9246);
nand U10404 (N_10404,N_9633,N_9869);
nand U10405 (N_10405,N_9864,N_9034);
or U10406 (N_10406,N_9010,N_9681);
nor U10407 (N_10407,N_9452,N_9852);
and U10408 (N_10408,N_9886,N_9497);
nand U10409 (N_10409,N_9910,N_9426);
and U10410 (N_10410,N_9225,N_9230);
nor U10411 (N_10411,N_9873,N_9438);
nand U10412 (N_10412,N_9500,N_9658);
and U10413 (N_10413,N_9084,N_9363);
nor U10414 (N_10414,N_9033,N_9573);
xnor U10415 (N_10415,N_9800,N_9776);
xor U10416 (N_10416,N_9062,N_9037);
and U10417 (N_10417,N_9266,N_9597);
nor U10418 (N_10418,N_9257,N_9962);
nand U10419 (N_10419,N_9526,N_9630);
and U10420 (N_10420,N_9119,N_9039);
or U10421 (N_10421,N_9911,N_9801);
nor U10422 (N_10422,N_9121,N_9640);
nor U10423 (N_10423,N_9992,N_9808);
or U10424 (N_10424,N_9643,N_9393);
and U10425 (N_10425,N_9528,N_9756);
xor U10426 (N_10426,N_9901,N_9125);
xor U10427 (N_10427,N_9414,N_9292);
nor U10428 (N_10428,N_9178,N_9813);
nor U10429 (N_10429,N_9327,N_9998);
nor U10430 (N_10430,N_9824,N_9495);
and U10431 (N_10431,N_9754,N_9400);
nand U10432 (N_10432,N_9499,N_9449);
and U10433 (N_10433,N_9296,N_9306);
xor U10434 (N_10434,N_9585,N_9122);
and U10435 (N_10435,N_9701,N_9772);
and U10436 (N_10436,N_9805,N_9948);
xnor U10437 (N_10437,N_9677,N_9751);
xnor U10438 (N_10438,N_9054,N_9862);
xor U10439 (N_10439,N_9606,N_9372);
nand U10440 (N_10440,N_9620,N_9730);
or U10441 (N_10441,N_9822,N_9839);
or U10442 (N_10442,N_9581,N_9052);
xor U10443 (N_10443,N_9578,N_9649);
nand U10444 (N_10444,N_9428,N_9858);
and U10445 (N_10445,N_9112,N_9031);
nand U10446 (N_10446,N_9834,N_9841);
and U10447 (N_10447,N_9444,N_9461);
xor U10448 (N_10448,N_9828,N_9726);
or U10449 (N_10449,N_9541,N_9013);
nor U10450 (N_10450,N_9151,N_9507);
or U10451 (N_10451,N_9650,N_9875);
xor U10452 (N_10452,N_9656,N_9376);
or U10453 (N_10453,N_9417,N_9740);
nor U10454 (N_10454,N_9108,N_9260);
xor U10455 (N_10455,N_9540,N_9674);
nand U10456 (N_10456,N_9482,N_9233);
xor U10457 (N_10457,N_9468,N_9553);
or U10458 (N_10458,N_9285,N_9981);
and U10459 (N_10459,N_9802,N_9833);
or U10460 (N_10460,N_9420,N_9294);
or U10461 (N_10461,N_9538,N_9765);
nand U10462 (N_10462,N_9422,N_9360);
and U10463 (N_10463,N_9303,N_9028);
xor U10464 (N_10464,N_9045,N_9900);
nor U10465 (N_10465,N_9668,N_9614);
or U10466 (N_10466,N_9082,N_9804);
nand U10467 (N_10467,N_9945,N_9988);
and U10468 (N_10468,N_9096,N_9362);
or U10469 (N_10469,N_9188,N_9695);
and U10470 (N_10470,N_9004,N_9474);
and U10471 (N_10471,N_9743,N_9974);
or U10472 (N_10472,N_9931,N_9791);
xor U10473 (N_10473,N_9192,N_9524);
or U10474 (N_10474,N_9582,N_9131);
or U10475 (N_10475,N_9177,N_9243);
nor U10476 (N_10476,N_9211,N_9621);
nand U10477 (N_10477,N_9190,N_9176);
and U10478 (N_10478,N_9375,N_9579);
xor U10479 (N_10479,N_9143,N_9295);
xnor U10480 (N_10480,N_9874,N_9810);
or U10481 (N_10481,N_9899,N_9753);
nand U10482 (N_10482,N_9485,N_9477);
or U10483 (N_10483,N_9764,N_9705);
xnor U10484 (N_10484,N_9183,N_9409);
xor U10485 (N_10485,N_9799,N_9209);
or U10486 (N_10486,N_9912,N_9457);
or U10487 (N_10487,N_9097,N_9588);
xor U10488 (N_10488,N_9590,N_9475);
nor U10489 (N_10489,N_9456,N_9609);
xnor U10490 (N_10490,N_9333,N_9596);
and U10491 (N_10491,N_9771,N_9817);
xor U10492 (N_10492,N_9252,N_9984);
or U10493 (N_10493,N_9480,N_9427);
and U10494 (N_10494,N_9089,N_9788);
and U10495 (N_10495,N_9665,N_9518);
or U10496 (N_10496,N_9626,N_9080);
and U10497 (N_10497,N_9239,N_9947);
xnor U10498 (N_10498,N_9023,N_9347);
xnor U10499 (N_10499,N_9093,N_9429);
nand U10500 (N_10500,N_9693,N_9670);
xor U10501 (N_10501,N_9652,N_9950);
nor U10502 (N_10502,N_9757,N_9542);
or U10503 (N_10503,N_9846,N_9808);
xnor U10504 (N_10504,N_9142,N_9371);
and U10505 (N_10505,N_9081,N_9804);
nand U10506 (N_10506,N_9997,N_9268);
nor U10507 (N_10507,N_9983,N_9322);
nand U10508 (N_10508,N_9764,N_9885);
nand U10509 (N_10509,N_9941,N_9908);
xor U10510 (N_10510,N_9271,N_9293);
nand U10511 (N_10511,N_9894,N_9064);
or U10512 (N_10512,N_9116,N_9451);
xnor U10513 (N_10513,N_9067,N_9142);
xnor U10514 (N_10514,N_9837,N_9265);
xor U10515 (N_10515,N_9987,N_9308);
and U10516 (N_10516,N_9457,N_9817);
nand U10517 (N_10517,N_9612,N_9619);
xor U10518 (N_10518,N_9560,N_9747);
or U10519 (N_10519,N_9171,N_9114);
or U10520 (N_10520,N_9357,N_9941);
nor U10521 (N_10521,N_9642,N_9266);
nor U10522 (N_10522,N_9290,N_9983);
or U10523 (N_10523,N_9623,N_9723);
and U10524 (N_10524,N_9667,N_9741);
and U10525 (N_10525,N_9499,N_9261);
and U10526 (N_10526,N_9191,N_9465);
nor U10527 (N_10527,N_9147,N_9324);
and U10528 (N_10528,N_9452,N_9461);
nor U10529 (N_10529,N_9134,N_9259);
nor U10530 (N_10530,N_9552,N_9349);
and U10531 (N_10531,N_9393,N_9166);
xnor U10532 (N_10532,N_9584,N_9993);
nor U10533 (N_10533,N_9479,N_9459);
or U10534 (N_10534,N_9897,N_9058);
nand U10535 (N_10535,N_9480,N_9191);
nand U10536 (N_10536,N_9265,N_9291);
or U10537 (N_10537,N_9595,N_9899);
or U10538 (N_10538,N_9995,N_9334);
and U10539 (N_10539,N_9825,N_9405);
nor U10540 (N_10540,N_9938,N_9085);
xnor U10541 (N_10541,N_9048,N_9696);
xnor U10542 (N_10542,N_9496,N_9225);
nor U10543 (N_10543,N_9580,N_9855);
and U10544 (N_10544,N_9610,N_9701);
and U10545 (N_10545,N_9715,N_9947);
nand U10546 (N_10546,N_9355,N_9225);
and U10547 (N_10547,N_9761,N_9075);
nand U10548 (N_10548,N_9553,N_9141);
and U10549 (N_10549,N_9813,N_9045);
nand U10550 (N_10550,N_9863,N_9710);
nor U10551 (N_10551,N_9997,N_9431);
nand U10552 (N_10552,N_9516,N_9437);
or U10553 (N_10553,N_9890,N_9650);
and U10554 (N_10554,N_9784,N_9869);
and U10555 (N_10555,N_9382,N_9924);
or U10556 (N_10556,N_9489,N_9510);
or U10557 (N_10557,N_9166,N_9296);
nand U10558 (N_10558,N_9022,N_9225);
or U10559 (N_10559,N_9896,N_9977);
xor U10560 (N_10560,N_9812,N_9405);
nand U10561 (N_10561,N_9622,N_9768);
and U10562 (N_10562,N_9873,N_9879);
xnor U10563 (N_10563,N_9284,N_9821);
xor U10564 (N_10564,N_9421,N_9689);
xor U10565 (N_10565,N_9384,N_9414);
and U10566 (N_10566,N_9437,N_9027);
nor U10567 (N_10567,N_9424,N_9716);
or U10568 (N_10568,N_9534,N_9395);
nand U10569 (N_10569,N_9661,N_9063);
nand U10570 (N_10570,N_9368,N_9117);
nand U10571 (N_10571,N_9892,N_9327);
or U10572 (N_10572,N_9409,N_9796);
and U10573 (N_10573,N_9521,N_9286);
nand U10574 (N_10574,N_9261,N_9652);
nor U10575 (N_10575,N_9203,N_9783);
xor U10576 (N_10576,N_9355,N_9382);
and U10577 (N_10577,N_9943,N_9684);
and U10578 (N_10578,N_9778,N_9915);
xor U10579 (N_10579,N_9298,N_9390);
nand U10580 (N_10580,N_9168,N_9867);
nand U10581 (N_10581,N_9115,N_9691);
nor U10582 (N_10582,N_9720,N_9168);
nand U10583 (N_10583,N_9038,N_9974);
and U10584 (N_10584,N_9573,N_9854);
and U10585 (N_10585,N_9838,N_9110);
nand U10586 (N_10586,N_9391,N_9171);
and U10587 (N_10587,N_9871,N_9720);
xor U10588 (N_10588,N_9062,N_9740);
nand U10589 (N_10589,N_9953,N_9297);
nor U10590 (N_10590,N_9966,N_9053);
or U10591 (N_10591,N_9218,N_9760);
xor U10592 (N_10592,N_9760,N_9807);
or U10593 (N_10593,N_9088,N_9830);
or U10594 (N_10594,N_9695,N_9256);
xnor U10595 (N_10595,N_9298,N_9942);
and U10596 (N_10596,N_9045,N_9596);
xor U10597 (N_10597,N_9700,N_9038);
and U10598 (N_10598,N_9470,N_9714);
nor U10599 (N_10599,N_9003,N_9851);
xnor U10600 (N_10600,N_9938,N_9642);
xor U10601 (N_10601,N_9604,N_9101);
nor U10602 (N_10602,N_9157,N_9624);
nor U10603 (N_10603,N_9482,N_9595);
or U10604 (N_10604,N_9449,N_9780);
or U10605 (N_10605,N_9347,N_9463);
nor U10606 (N_10606,N_9640,N_9971);
nand U10607 (N_10607,N_9529,N_9228);
xnor U10608 (N_10608,N_9299,N_9339);
nor U10609 (N_10609,N_9539,N_9959);
or U10610 (N_10610,N_9021,N_9999);
nand U10611 (N_10611,N_9305,N_9234);
xor U10612 (N_10612,N_9370,N_9891);
or U10613 (N_10613,N_9324,N_9738);
and U10614 (N_10614,N_9708,N_9977);
xnor U10615 (N_10615,N_9002,N_9419);
and U10616 (N_10616,N_9279,N_9332);
xor U10617 (N_10617,N_9519,N_9563);
and U10618 (N_10618,N_9982,N_9471);
and U10619 (N_10619,N_9797,N_9215);
and U10620 (N_10620,N_9039,N_9111);
xor U10621 (N_10621,N_9749,N_9310);
nor U10622 (N_10622,N_9074,N_9104);
nand U10623 (N_10623,N_9996,N_9741);
xnor U10624 (N_10624,N_9811,N_9711);
and U10625 (N_10625,N_9773,N_9896);
and U10626 (N_10626,N_9594,N_9577);
or U10627 (N_10627,N_9204,N_9532);
nor U10628 (N_10628,N_9356,N_9196);
xor U10629 (N_10629,N_9158,N_9096);
nand U10630 (N_10630,N_9075,N_9222);
xor U10631 (N_10631,N_9798,N_9973);
nor U10632 (N_10632,N_9327,N_9603);
xor U10633 (N_10633,N_9386,N_9745);
nand U10634 (N_10634,N_9103,N_9751);
or U10635 (N_10635,N_9111,N_9215);
nor U10636 (N_10636,N_9786,N_9942);
nor U10637 (N_10637,N_9903,N_9325);
and U10638 (N_10638,N_9597,N_9200);
and U10639 (N_10639,N_9902,N_9591);
nand U10640 (N_10640,N_9485,N_9005);
xnor U10641 (N_10641,N_9914,N_9250);
xor U10642 (N_10642,N_9333,N_9412);
nand U10643 (N_10643,N_9691,N_9147);
or U10644 (N_10644,N_9906,N_9385);
or U10645 (N_10645,N_9121,N_9997);
nor U10646 (N_10646,N_9290,N_9980);
nand U10647 (N_10647,N_9973,N_9449);
xnor U10648 (N_10648,N_9012,N_9998);
nand U10649 (N_10649,N_9721,N_9433);
or U10650 (N_10650,N_9134,N_9079);
xor U10651 (N_10651,N_9883,N_9241);
xor U10652 (N_10652,N_9190,N_9505);
xor U10653 (N_10653,N_9491,N_9489);
nand U10654 (N_10654,N_9004,N_9560);
and U10655 (N_10655,N_9428,N_9215);
xor U10656 (N_10656,N_9361,N_9945);
and U10657 (N_10657,N_9957,N_9686);
nand U10658 (N_10658,N_9126,N_9288);
or U10659 (N_10659,N_9426,N_9214);
xnor U10660 (N_10660,N_9727,N_9897);
nor U10661 (N_10661,N_9564,N_9468);
xnor U10662 (N_10662,N_9450,N_9070);
or U10663 (N_10663,N_9910,N_9879);
xor U10664 (N_10664,N_9560,N_9823);
and U10665 (N_10665,N_9617,N_9543);
nand U10666 (N_10666,N_9831,N_9419);
xor U10667 (N_10667,N_9597,N_9803);
xnor U10668 (N_10668,N_9719,N_9299);
xnor U10669 (N_10669,N_9111,N_9280);
nor U10670 (N_10670,N_9989,N_9285);
nand U10671 (N_10671,N_9922,N_9649);
nand U10672 (N_10672,N_9261,N_9722);
xor U10673 (N_10673,N_9709,N_9393);
and U10674 (N_10674,N_9834,N_9999);
xnor U10675 (N_10675,N_9598,N_9241);
nor U10676 (N_10676,N_9487,N_9308);
and U10677 (N_10677,N_9909,N_9520);
nand U10678 (N_10678,N_9946,N_9423);
xor U10679 (N_10679,N_9957,N_9305);
or U10680 (N_10680,N_9649,N_9624);
xnor U10681 (N_10681,N_9434,N_9848);
or U10682 (N_10682,N_9978,N_9547);
and U10683 (N_10683,N_9813,N_9612);
nand U10684 (N_10684,N_9198,N_9464);
nand U10685 (N_10685,N_9141,N_9541);
and U10686 (N_10686,N_9627,N_9098);
or U10687 (N_10687,N_9885,N_9591);
or U10688 (N_10688,N_9241,N_9311);
nor U10689 (N_10689,N_9139,N_9099);
or U10690 (N_10690,N_9385,N_9212);
nand U10691 (N_10691,N_9750,N_9433);
xor U10692 (N_10692,N_9488,N_9397);
or U10693 (N_10693,N_9599,N_9675);
nor U10694 (N_10694,N_9700,N_9336);
xor U10695 (N_10695,N_9615,N_9501);
nand U10696 (N_10696,N_9857,N_9404);
xor U10697 (N_10697,N_9248,N_9388);
nor U10698 (N_10698,N_9567,N_9667);
or U10699 (N_10699,N_9392,N_9272);
and U10700 (N_10700,N_9481,N_9275);
and U10701 (N_10701,N_9495,N_9620);
and U10702 (N_10702,N_9612,N_9679);
or U10703 (N_10703,N_9026,N_9290);
xnor U10704 (N_10704,N_9402,N_9014);
or U10705 (N_10705,N_9107,N_9850);
and U10706 (N_10706,N_9114,N_9645);
xor U10707 (N_10707,N_9744,N_9677);
or U10708 (N_10708,N_9764,N_9756);
xnor U10709 (N_10709,N_9377,N_9512);
xor U10710 (N_10710,N_9023,N_9743);
and U10711 (N_10711,N_9371,N_9028);
nand U10712 (N_10712,N_9627,N_9618);
nor U10713 (N_10713,N_9568,N_9397);
nor U10714 (N_10714,N_9373,N_9610);
and U10715 (N_10715,N_9477,N_9377);
and U10716 (N_10716,N_9637,N_9881);
and U10717 (N_10717,N_9594,N_9569);
nand U10718 (N_10718,N_9080,N_9707);
nor U10719 (N_10719,N_9779,N_9196);
nand U10720 (N_10720,N_9164,N_9109);
xor U10721 (N_10721,N_9853,N_9587);
or U10722 (N_10722,N_9777,N_9192);
nand U10723 (N_10723,N_9452,N_9630);
nand U10724 (N_10724,N_9054,N_9303);
xor U10725 (N_10725,N_9699,N_9536);
and U10726 (N_10726,N_9986,N_9006);
nand U10727 (N_10727,N_9070,N_9264);
nor U10728 (N_10728,N_9898,N_9020);
or U10729 (N_10729,N_9642,N_9450);
and U10730 (N_10730,N_9517,N_9004);
nor U10731 (N_10731,N_9764,N_9447);
xnor U10732 (N_10732,N_9346,N_9861);
or U10733 (N_10733,N_9916,N_9462);
nor U10734 (N_10734,N_9218,N_9661);
or U10735 (N_10735,N_9683,N_9787);
nand U10736 (N_10736,N_9797,N_9443);
nor U10737 (N_10737,N_9546,N_9632);
xnor U10738 (N_10738,N_9149,N_9761);
nor U10739 (N_10739,N_9464,N_9224);
nor U10740 (N_10740,N_9283,N_9631);
and U10741 (N_10741,N_9273,N_9025);
nand U10742 (N_10742,N_9576,N_9787);
and U10743 (N_10743,N_9314,N_9629);
nor U10744 (N_10744,N_9504,N_9248);
or U10745 (N_10745,N_9624,N_9866);
or U10746 (N_10746,N_9818,N_9246);
nor U10747 (N_10747,N_9178,N_9362);
and U10748 (N_10748,N_9155,N_9033);
and U10749 (N_10749,N_9702,N_9801);
or U10750 (N_10750,N_9063,N_9245);
or U10751 (N_10751,N_9236,N_9589);
and U10752 (N_10752,N_9157,N_9294);
xnor U10753 (N_10753,N_9793,N_9330);
nor U10754 (N_10754,N_9585,N_9035);
nor U10755 (N_10755,N_9871,N_9446);
or U10756 (N_10756,N_9914,N_9155);
or U10757 (N_10757,N_9143,N_9487);
or U10758 (N_10758,N_9907,N_9291);
nor U10759 (N_10759,N_9502,N_9484);
nand U10760 (N_10760,N_9379,N_9985);
nand U10761 (N_10761,N_9806,N_9780);
and U10762 (N_10762,N_9165,N_9320);
nor U10763 (N_10763,N_9563,N_9985);
xor U10764 (N_10764,N_9624,N_9805);
and U10765 (N_10765,N_9565,N_9781);
and U10766 (N_10766,N_9259,N_9239);
nand U10767 (N_10767,N_9221,N_9775);
and U10768 (N_10768,N_9449,N_9792);
or U10769 (N_10769,N_9373,N_9862);
nor U10770 (N_10770,N_9568,N_9511);
and U10771 (N_10771,N_9374,N_9821);
nand U10772 (N_10772,N_9253,N_9702);
xnor U10773 (N_10773,N_9933,N_9703);
nand U10774 (N_10774,N_9986,N_9088);
or U10775 (N_10775,N_9880,N_9337);
nor U10776 (N_10776,N_9015,N_9228);
nand U10777 (N_10777,N_9258,N_9099);
nor U10778 (N_10778,N_9075,N_9481);
or U10779 (N_10779,N_9803,N_9754);
xor U10780 (N_10780,N_9218,N_9442);
nand U10781 (N_10781,N_9781,N_9243);
and U10782 (N_10782,N_9382,N_9622);
nor U10783 (N_10783,N_9014,N_9759);
xnor U10784 (N_10784,N_9219,N_9058);
and U10785 (N_10785,N_9706,N_9799);
nor U10786 (N_10786,N_9920,N_9025);
and U10787 (N_10787,N_9746,N_9295);
xor U10788 (N_10788,N_9148,N_9928);
nand U10789 (N_10789,N_9860,N_9813);
nor U10790 (N_10790,N_9479,N_9829);
xnor U10791 (N_10791,N_9379,N_9724);
nor U10792 (N_10792,N_9455,N_9837);
nand U10793 (N_10793,N_9327,N_9635);
nor U10794 (N_10794,N_9713,N_9910);
nand U10795 (N_10795,N_9149,N_9461);
nand U10796 (N_10796,N_9188,N_9668);
nor U10797 (N_10797,N_9173,N_9933);
xnor U10798 (N_10798,N_9415,N_9731);
nor U10799 (N_10799,N_9416,N_9949);
nand U10800 (N_10800,N_9564,N_9815);
xnor U10801 (N_10801,N_9586,N_9523);
nor U10802 (N_10802,N_9255,N_9022);
nand U10803 (N_10803,N_9916,N_9047);
and U10804 (N_10804,N_9363,N_9651);
and U10805 (N_10805,N_9087,N_9999);
nor U10806 (N_10806,N_9702,N_9054);
nand U10807 (N_10807,N_9251,N_9170);
xnor U10808 (N_10808,N_9907,N_9630);
nor U10809 (N_10809,N_9582,N_9759);
xor U10810 (N_10810,N_9842,N_9943);
or U10811 (N_10811,N_9155,N_9472);
nand U10812 (N_10812,N_9027,N_9723);
xnor U10813 (N_10813,N_9900,N_9716);
xnor U10814 (N_10814,N_9899,N_9625);
and U10815 (N_10815,N_9692,N_9314);
nor U10816 (N_10816,N_9293,N_9670);
nand U10817 (N_10817,N_9951,N_9682);
and U10818 (N_10818,N_9432,N_9223);
nand U10819 (N_10819,N_9596,N_9738);
or U10820 (N_10820,N_9186,N_9168);
or U10821 (N_10821,N_9401,N_9952);
or U10822 (N_10822,N_9948,N_9090);
or U10823 (N_10823,N_9047,N_9960);
xnor U10824 (N_10824,N_9333,N_9581);
and U10825 (N_10825,N_9220,N_9414);
and U10826 (N_10826,N_9399,N_9110);
and U10827 (N_10827,N_9338,N_9069);
nor U10828 (N_10828,N_9295,N_9614);
nand U10829 (N_10829,N_9267,N_9531);
and U10830 (N_10830,N_9678,N_9901);
or U10831 (N_10831,N_9382,N_9515);
xnor U10832 (N_10832,N_9050,N_9148);
and U10833 (N_10833,N_9896,N_9051);
nand U10834 (N_10834,N_9329,N_9176);
nor U10835 (N_10835,N_9974,N_9884);
xnor U10836 (N_10836,N_9221,N_9403);
nand U10837 (N_10837,N_9706,N_9803);
nand U10838 (N_10838,N_9337,N_9628);
xnor U10839 (N_10839,N_9985,N_9724);
nor U10840 (N_10840,N_9872,N_9185);
nor U10841 (N_10841,N_9996,N_9507);
nor U10842 (N_10842,N_9766,N_9282);
nand U10843 (N_10843,N_9345,N_9440);
xor U10844 (N_10844,N_9940,N_9982);
nor U10845 (N_10845,N_9815,N_9870);
nor U10846 (N_10846,N_9923,N_9040);
nor U10847 (N_10847,N_9904,N_9605);
nand U10848 (N_10848,N_9442,N_9384);
and U10849 (N_10849,N_9095,N_9937);
and U10850 (N_10850,N_9060,N_9603);
nor U10851 (N_10851,N_9871,N_9188);
or U10852 (N_10852,N_9172,N_9294);
and U10853 (N_10853,N_9523,N_9156);
nor U10854 (N_10854,N_9027,N_9327);
or U10855 (N_10855,N_9459,N_9579);
or U10856 (N_10856,N_9545,N_9211);
nor U10857 (N_10857,N_9116,N_9376);
xor U10858 (N_10858,N_9163,N_9422);
and U10859 (N_10859,N_9660,N_9785);
nand U10860 (N_10860,N_9061,N_9984);
xor U10861 (N_10861,N_9740,N_9790);
xor U10862 (N_10862,N_9403,N_9809);
nor U10863 (N_10863,N_9675,N_9344);
nand U10864 (N_10864,N_9793,N_9716);
or U10865 (N_10865,N_9924,N_9555);
or U10866 (N_10866,N_9469,N_9213);
xor U10867 (N_10867,N_9724,N_9729);
xnor U10868 (N_10868,N_9488,N_9892);
nand U10869 (N_10869,N_9044,N_9103);
nand U10870 (N_10870,N_9086,N_9215);
nor U10871 (N_10871,N_9693,N_9226);
nor U10872 (N_10872,N_9081,N_9241);
nor U10873 (N_10873,N_9374,N_9281);
xor U10874 (N_10874,N_9435,N_9977);
or U10875 (N_10875,N_9161,N_9860);
nor U10876 (N_10876,N_9747,N_9854);
nor U10877 (N_10877,N_9310,N_9887);
nand U10878 (N_10878,N_9649,N_9122);
xor U10879 (N_10879,N_9089,N_9274);
nand U10880 (N_10880,N_9585,N_9000);
nand U10881 (N_10881,N_9612,N_9273);
nor U10882 (N_10882,N_9031,N_9074);
nand U10883 (N_10883,N_9411,N_9643);
nand U10884 (N_10884,N_9888,N_9491);
nor U10885 (N_10885,N_9749,N_9891);
or U10886 (N_10886,N_9344,N_9736);
xor U10887 (N_10887,N_9901,N_9512);
and U10888 (N_10888,N_9787,N_9491);
or U10889 (N_10889,N_9614,N_9519);
nor U10890 (N_10890,N_9320,N_9474);
or U10891 (N_10891,N_9965,N_9889);
or U10892 (N_10892,N_9002,N_9014);
nand U10893 (N_10893,N_9404,N_9891);
nand U10894 (N_10894,N_9203,N_9513);
and U10895 (N_10895,N_9928,N_9612);
nor U10896 (N_10896,N_9567,N_9935);
or U10897 (N_10897,N_9278,N_9656);
nand U10898 (N_10898,N_9924,N_9996);
nor U10899 (N_10899,N_9703,N_9189);
nor U10900 (N_10900,N_9343,N_9400);
xnor U10901 (N_10901,N_9967,N_9877);
xor U10902 (N_10902,N_9986,N_9390);
xor U10903 (N_10903,N_9293,N_9537);
and U10904 (N_10904,N_9779,N_9805);
nor U10905 (N_10905,N_9685,N_9991);
or U10906 (N_10906,N_9970,N_9101);
xor U10907 (N_10907,N_9342,N_9294);
nor U10908 (N_10908,N_9461,N_9586);
nor U10909 (N_10909,N_9061,N_9721);
nand U10910 (N_10910,N_9692,N_9452);
nand U10911 (N_10911,N_9974,N_9028);
nor U10912 (N_10912,N_9787,N_9066);
or U10913 (N_10913,N_9937,N_9857);
nand U10914 (N_10914,N_9128,N_9672);
nor U10915 (N_10915,N_9718,N_9953);
nand U10916 (N_10916,N_9972,N_9821);
or U10917 (N_10917,N_9563,N_9950);
and U10918 (N_10918,N_9939,N_9070);
and U10919 (N_10919,N_9801,N_9821);
nor U10920 (N_10920,N_9873,N_9493);
and U10921 (N_10921,N_9082,N_9433);
xnor U10922 (N_10922,N_9783,N_9440);
and U10923 (N_10923,N_9095,N_9166);
xor U10924 (N_10924,N_9133,N_9634);
xnor U10925 (N_10925,N_9350,N_9520);
xnor U10926 (N_10926,N_9222,N_9894);
xor U10927 (N_10927,N_9659,N_9412);
xnor U10928 (N_10928,N_9360,N_9020);
or U10929 (N_10929,N_9144,N_9971);
or U10930 (N_10930,N_9941,N_9566);
xnor U10931 (N_10931,N_9788,N_9133);
nand U10932 (N_10932,N_9130,N_9132);
and U10933 (N_10933,N_9534,N_9133);
or U10934 (N_10934,N_9902,N_9885);
and U10935 (N_10935,N_9799,N_9460);
or U10936 (N_10936,N_9878,N_9856);
and U10937 (N_10937,N_9772,N_9615);
and U10938 (N_10938,N_9214,N_9847);
nor U10939 (N_10939,N_9392,N_9929);
xor U10940 (N_10940,N_9225,N_9495);
xor U10941 (N_10941,N_9500,N_9282);
nor U10942 (N_10942,N_9777,N_9621);
or U10943 (N_10943,N_9529,N_9594);
nor U10944 (N_10944,N_9219,N_9513);
or U10945 (N_10945,N_9746,N_9473);
and U10946 (N_10946,N_9656,N_9949);
nand U10947 (N_10947,N_9222,N_9509);
nor U10948 (N_10948,N_9189,N_9713);
or U10949 (N_10949,N_9886,N_9989);
nor U10950 (N_10950,N_9954,N_9022);
nor U10951 (N_10951,N_9618,N_9939);
nor U10952 (N_10952,N_9041,N_9392);
nor U10953 (N_10953,N_9594,N_9671);
nor U10954 (N_10954,N_9340,N_9005);
or U10955 (N_10955,N_9740,N_9989);
or U10956 (N_10956,N_9391,N_9987);
and U10957 (N_10957,N_9920,N_9137);
nor U10958 (N_10958,N_9220,N_9804);
xnor U10959 (N_10959,N_9763,N_9707);
nand U10960 (N_10960,N_9915,N_9226);
nand U10961 (N_10961,N_9236,N_9555);
xor U10962 (N_10962,N_9052,N_9505);
nor U10963 (N_10963,N_9609,N_9486);
and U10964 (N_10964,N_9118,N_9493);
nand U10965 (N_10965,N_9660,N_9500);
or U10966 (N_10966,N_9469,N_9872);
or U10967 (N_10967,N_9495,N_9750);
nand U10968 (N_10968,N_9271,N_9632);
or U10969 (N_10969,N_9824,N_9966);
nor U10970 (N_10970,N_9529,N_9352);
xor U10971 (N_10971,N_9277,N_9079);
and U10972 (N_10972,N_9194,N_9564);
and U10973 (N_10973,N_9917,N_9142);
and U10974 (N_10974,N_9473,N_9263);
or U10975 (N_10975,N_9959,N_9839);
and U10976 (N_10976,N_9828,N_9231);
or U10977 (N_10977,N_9174,N_9596);
and U10978 (N_10978,N_9332,N_9029);
nand U10979 (N_10979,N_9487,N_9927);
and U10980 (N_10980,N_9338,N_9349);
and U10981 (N_10981,N_9270,N_9313);
and U10982 (N_10982,N_9576,N_9545);
and U10983 (N_10983,N_9876,N_9652);
nand U10984 (N_10984,N_9332,N_9378);
xnor U10985 (N_10985,N_9446,N_9175);
xnor U10986 (N_10986,N_9725,N_9633);
or U10987 (N_10987,N_9715,N_9774);
nor U10988 (N_10988,N_9258,N_9583);
nand U10989 (N_10989,N_9505,N_9163);
nand U10990 (N_10990,N_9397,N_9960);
and U10991 (N_10991,N_9452,N_9103);
nand U10992 (N_10992,N_9857,N_9282);
nor U10993 (N_10993,N_9935,N_9812);
xor U10994 (N_10994,N_9910,N_9415);
and U10995 (N_10995,N_9461,N_9286);
and U10996 (N_10996,N_9993,N_9564);
nor U10997 (N_10997,N_9383,N_9713);
nand U10998 (N_10998,N_9826,N_9370);
or U10999 (N_10999,N_9110,N_9519);
nor U11000 (N_11000,N_10236,N_10186);
xnor U11001 (N_11001,N_10091,N_10679);
nand U11002 (N_11002,N_10213,N_10732);
or U11003 (N_11003,N_10767,N_10579);
xor U11004 (N_11004,N_10333,N_10825);
nand U11005 (N_11005,N_10136,N_10821);
nor U11006 (N_11006,N_10835,N_10603);
nor U11007 (N_11007,N_10640,N_10100);
and U11008 (N_11008,N_10770,N_10085);
xnor U11009 (N_11009,N_10406,N_10991);
or U11010 (N_11010,N_10250,N_10626);
and U11011 (N_11011,N_10853,N_10096);
nor U11012 (N_11012,N_10785,N_10231);
nand U11013 (N_11013,N_10432,N_10163);
or U11014 (N_11014,N_10536,N_10866);
nand U11015 (N_11015,N_10869,N_10147);
and U11016 (N_11016,N_10949,N_10989);
and U11017 (N_11017,N_10562,N_10824);
nand U11018 (N_11018,N_10534,N_10707);
nor U11019 (N_11019,N_10962,N_10245);
or U11020 (N_11020,N_10628,N_10295);
xnor U11021 (N_11021,N_10296,N_10129);
nand U11022 (N_11022,N_10248,N_10590);
nor U11023 (N_11023,N_10179,N_10318);
nand U11024 (N_11024,N_10609,N_10778);
or U11025 (N_11025,N_10905,N_10385);
or U11026 (N_11026,N_10342,N_10030);
or U11027 (N_11027,N_10440,N_10274);
or U11028 (N_11028,N_10014,N_10366);
and U11029 (N_11029,N_10346,N_10126);
nand U11030 (N_11030,N_10202,N_10069);
nor U11031 (N_11031,N_10508,N_10933);
nor U11032 (N_11032,N_10697,N_10336);
nor U11033 (N_11033,N_10084,N_10010);
nor U11034 (N_11034,N_10783,N_10430);
nor U11035 (N_11035,N_10545,N_10565);
nand U11036 (N_11036,N_10715,N_10407);
nand U11037 (N_11037,N_10196,N_10944);
xnor U11038 (N_11038,N_10374,N_10125);
nor U11039 (N_11039,N_10303,N_10742);
or U11040 (N_11040,N_10329,N_10643);
nand U11041 (N_11041,N_10919,N_10714);
nand U11042 (N_11042,N_10820,N_10513);
nand U11043 (N_11043,N_10674,N_10755);
or U11044 (N_11044,N_10034,N_10752);
xnor U11045 (N_11045,N_10491,N_10849);
and U11046 (N_11046,N_10401,N_10909);
and U11047 (N_11047,N_10768,N_10546);
nor U11048 (N_11048,N_10867,N_10376);
and U11049 (N_11049,N_10394,N_10036);
xnor U11050 (N_11050,N_10544,N_10288);
nor U11051 (N_11051,N_10223,N_10306);
or U11052 (N_11052,N_10352,N_10542);
or U11053 (N_11053,N_10387,N_10984);
xor U11054 (N_11054,N_10819,N_10335);
nor U11055 (N_11055,N_10008,N_10927);
nor U11056 (N_11056,N_10974,N_10311);
nor U11057 (N_11057,N_10973,N_10167);
and U11058 (N_11058,N_10852,N_10595);
xor U11059 (N_11059,N_10165,N_10698);
xnor U11060 (N_11060,N_10533,N_10593);
or U11061 (N_11061,N_10415,N_10906);
or U11062 (N_11062,N_10171,N_10522);
xnor U11063 (N_11063,N_10591,N_10629);
nand U11064 (N_11064,N_10003,N_10161);
xnor U11065 (N_11065,N_10656,N_10130);
nor U11066 (N_11066,N_10627,N_10718);
or U11067 (N_11067,N_10257,N_10775);
nand U11068 (N_11068,N_10605,N_10964);
nor U11069 (N_11069,N_10841,N_10281);
nand U11070 (N_11070,N_10511,N_10237);
nor U11071 (N_11071,N_10174,N_10235);
nand U11072 (N_11072,N_10453,N_10361);
nor U11073 (N_11073,N_10576,N_10194);
or U11074 (N_11074,N_10381,N_10134);
xnor U11075 (N_11075,N_10398,N_10239);
or U11076 (N_11076,N_10816,N_10804);
nor U11077 (N_11077,N_10782,N_10462);
or U11078 (N_11078,N_10688,N_10308);
or U11079 (N_11079,N_10280,N_10947);
nor U11080 (N_11080,N_10332,N_10547);
or U11081 (N_11081,N_10243,N_10753);
nor U11082 (N_11082,N_10710,N_10878);
nor U11083 (N_11083,N_10363,N_10300);
or U11084 (N_11084,N_10327,N_10203);
xnor U11085 (N_11085,N_10713,N_10302);
xor U11086 (N_11086,N_10903,N_10813);
and U11087 (N_11087,N_10173,N_10960);
nor U11088 (N_11088,N_10514,N_10086);
nand U11089 (N_11089,N_10611,N_10420);
or U11090 (N_11090,N_10341,N_10001);
or U11091 (N_11091,N_10264,N_10836);
nand U11092 (N_11092,N_10178,N_10959);
or U11093 (N_11093,N_10505,N_10166);
xor U11094 (N_11094,N_10695,N_10693);
nor U11095 (N_11095,N_10393,N_10487);
and U11096 (N_11096,N_10224,N_10429);
nand U11097 (N_11097,N_10645,N_10655);
and U11098 (N_11098,N_10523,N_10340);
nor U11099 (N_11099,N_10484,N_10143);
nand U11100 (N_11100,N_10868,N_10317);
xor U11101 (N_11101,N_10833,N_10578);
and U11102 (N_11102,N_10798,N_10496);
xor U11103 (N_11103,N_10653,N_10081);
and U11104 (N_11104,N_10470,N_10048);
or U11105 (N_11105,N_10249,N_10399);
nor U11106 (N_11106,N_10856,N_10677);
or U11107 (N_11107,N_10071,N_10610);
nand U11108 (N_11108,N_10559,N_10145);
nand U11109 (N_11109,N_10663,N_10594);
xnor U11110 (N_11110,N_10386,N_10598);
nand U11111 (N_11111,N_10185,N_10552);
nor U11112 (N_11112,N_10826,N_10620);
xnor U11113 (N_11113,N_10774,N_10551);
and U11114 (N_11114,N_10097,N_10073);
nand U11115 (N_11115,N_10712,N_10560);
xnor U11116 (N_11116,N_10809,N_10894);
and U11117 (N_11117,N_10686,N_10692);
and U11118 (N_11118,N_10467,N_10460);
or U11119 (N_11119,N_10419,N_10823);
or U11120 (N_11120,N_10937,N_10006);
nor U11121 (N_11121,N_10606,N_10735);
xor U11122 (N_11122,N_10017,N_10337);
and U11123 (N_11123,N_10998,N_10951);
or U11124 (N_11124,N_10221,N_10180);
nand U11125 (N_11125,N_10876,N_10209);
and U11126 (N_11126,N_10910,N_10635);
nor U11127 (N_11127,N_10204,N_10094);
nor U11128 (N_11128,N_10259,N_10210);
or U11129 (N_11129,N_10769,N_10586);
xnor U11130 (N_11130,N_10763,N_10472);
and U11131 (N_11131,N_10344,N_10963);
nor U11132 (N_11132,N_10276,N_10811);
nor U11133 (N_11133,N_10900,N_10928);
and U11134 (N_11134,N_10189,N_10696);
nand U11135 (N_11135,N_10284,N_10675);
or U11136 (N_11136,N_10741,N_10338);
xnor U11137 (N_11137,N_10761,N_10700);
xnor U11138 (N_11138,N_10754,N_10382);
or U11139 (N_11139,N_10499,N_10654);
nand U11140 (N_11140,N_10260,N_10349);
nor U11141 (N_11141,N_10877,N_10583);
nand U11142 (N_11142,N_10050,N_10557);
or U11143 (N_11143,N_10685,N_10132);
or U11144 (N_11144,N_10142,N_10988);
or U11145 (N_11145,N_10657,N_10026);
and U11146 (N_11146,N_10681,N_10212);
nand U11147 (N_11147,N_10254,N_10834);
nand U11148 (N_11148,N_10116,N_10446);
and U11149 (N_11149,N_10294,N_10445);
and U11150 (N_11150,N_10854,N_10351);
nand U11151 (N_11151,N_10018,N_10885);
or U11152 (N_11152,N_10241,N_10584);
or U11153 (N_11153,N_10322,N_10131);
nand U11154 (N_11154,N_10067,N_10007);
nand U11155 (N_11155,N_10531,N_10155);
nand U11156 (N_11156,N_10301,N_10678);
and U11157 (N_11157,N_10055,N_10745);
xor U11158 (N_11158,N_10737,N_10566);
nand U11159 (N_11159,N_10307,N_10286);
or U11160 (N_11160,N_10490,N_10493);
and U11161 (N_11161,N_10582,N_10451);
nand U11162 (N_11162,N_10345,N_10730);
nand U11163 (N_11163,N_10787,N_10799);
nor U11164 (N_11164,N_10230,N_10765);
nor U11165 (N_11165,N_10733,N_10556);
xnor U11166 (N_11166,N_10158,N_10780);
and U11167 (N_11167,N_10646,N_10183);
or U11168 (N_11168,N_10672,N_10516);
nor U11169 (N_11169,N_10413,N_10454);
and U11170 (N_11170,N_10795,N_10471);
xor U11171 (N_11171,N_10388,N_10265);
nand U11172 (N_11172,N_10734,N_10012);
nand U11173 (N_11173,N_10256,N_10831);
nor U11174 (N_11174,N_10309,N_10882);
nor U11175 (N_11175,N_10450,N_10773);
xnor U11176 (N_11176,N_10104,N_10115);
and U11177 (N_11177,N_10297,N_10358);
or U11178 (N_11178,N_10503,N_10364);
and U11179 (N_11179,N_10362,N_10673);
nor U11180 (N_11180,N_10431,N_10561);
xor U11181 (N_11181,N_10328,N_10624);
xor U11182 (N_11182,N_10187,N_10711);
and U11183 (N_11183,N_10671,N_10918);
xnor U11184 (N_11184,N_10205,N_10893);
xor U11185 (N_11185,N_10433,N_10781);
nand U11186 (N_11186,N_10400,N_10383);
xor U11187 (N_11187,N_10121,N_10033);
or U11188 (N_11188,N_10438,N_10901);
or U11189 (N_11189,N_10888,N_10936);
xor U11190 (N_11190,N_10389,N_10886);
nand U11191 (N_11191,N_10043,N_10028);
or U11192 (N_11192,N_10577,N_10418);
and U11193 (N_11193,N_10762,N_10666);
nor U11194 (N_11194,N_10153,N_10786);
xor U11195 (N_11195,N_10234,N_10779);
nor U11196 (N_11196,N_10720,N_10156);
and U11197 (N_11197,N_10792,N_10887);
and U11198 (N_11198,N_10979,N_10573);
and U11199 (N_11199,N_10558,N_10169);
or U11200 (N_11200,N_10473,N_10575);
and U11201 (N_11201,N_10099,N_10537);
or U11202 (N_11202,N_10079,N_10638);
and U11203 (N_11203,N_10520,N_10022);
or U11204 (N_11204,N_10943,N_10369);
xor U11205 (N_11205,N_10980,N_10992);
xnor U11206 (N_11206,N_10676,N_10421);
xnor U11207 (N_11207,N_10863,N_10495);
xnor U11208 (N_11208,N_10188,N_10585);
xnor U11209 (N_11209,N_10312,N_10310);
or U11210 (N_11210,N_10649,N_10216);
nor U11211 (N_11211,N_10228,N_10667);
or U11212 (N_11212,N_10981,N_10412);
nand U11213 (N_11213,N_10957,N_10739);
nand U11214 (N_11214,N_10873,N_10444);
nor U11215 (N_11215,N_10896,N_10011);
xor U11216 (N_11216,N_10347,N_10160);
and U11217 (N_11217,N_10539,N_10409);
nand U11218 (N_11218,N_10892,N_10760);
xor U11219 (N_11219,N_10941,N_10904);
nor U11220 (N_11220,N_10808,N_10634);
nand U11221 (N_11221,N_10191,N_10285);
or U11222 (N_11222,N_10612,N_10047);
xnor U11223 (N_11223,N_10706,N_10855);
and U11224 (N_11224,N_10946,N_10016);
xor U11225 (N_11225,N_10651,N_10682);
and U11226 (N_11226,N_10837,N_10112);
xnor U11227 (N_11227,N_10497,N_10320);
xnor U11228 (N_11228,N_10278,N_10506);
xor U11229 (N_11229,N_10743,N_10987);
xnor U11230 (N_11230,N_10997,N_10481);
xor U11231 (N_11231,N_10217,N_10891);
and U11232 (N_11232,N_10436,N_10832);
nand U11233 (N_11233,N_10330,N_10670);
nor U11234 (N_11234,N_10072,N_10690);
xnor U11235 (N_11235,N_10299,N_10907);
or U11236 (N_11236,N_10262,N_10291);
or U11237 (N_11237,N_10902,N_10990);
and U11238 (N_11238,N_10468,N_10923);
nor U11239 (N_11239,N_10077,N_10550);
nand U11240 (N_11240,N_10717,N_10190);
nor U11241 (N_11241,N_10592,N_10353);
nor U11242 (N_11242,N_10095,N_10922);
nand U11243 (N_11243,N_10540,N_10969);
nand U11244 (N_11244,N_10865,N_10405);
or U11245 (N_11245,N_10372,N_10159);
or U11246 (N_11246,N_10749,N_10459);
and U11247 (N_11247,N_10838,N_10553);
or U11248 (N_11248,N_10647,N_10709);
xor U11249 (N_11249,N_10268,N_10524);
and U11250 (N_11250,N_10045,N_10040);
xor U11251 (N_11251,N_10983,N_10510);
or U11252 (N_11252,N_10059,N_10958);
nand U11253 (N_11253,N_10122,N_10083);
xnor U11254 (N_11254,N_10633,N_10541);
and U11255 (N_11255,N_10478,N_10689);
nor U11256 (N_11256,N_10965,N_10035);
nand U11257 (N_11257,N_10642,N_10365);
nand U11258 (N_11258,N_10426,N_10207);
and U11259 (N_11259,N_10177,N_10051);
nor U11260 (N_11260,N_10092,N_10683);
or U11261 (N_11261,N_10117,N_10597);
and U11262 (N_11262,N_10273,N_10476);
and U11263 (N_11263,N_10859,N_10277);
nor U11264 (N_11264,N_10144,N_10538);
nand U11265 (N_11265,N_10848,N_10384);
xnor U11266 (N_11266,N_10261,N_10925);
and U11267 (N_11267,N_10985,N_10747);
xor U11268 (N_11268,N_10915,N_10049);
nor U11269 (N_11269,N_10549,N_10862);
nand U11270 (N_11270,N_10800,N_10818);
nand U11271 (N_11271,N_10064,N_10618);
nand U11272 (N_11272,N_10660,N_10750);
nor U11273 (N_11273,N_10563,N_10282);
nor U11274 (N_11274,N_10184,N_10982);
nor U11275 (N_11275,N_10266,N_10108);
or U11276 (N_11276,N_10827,N_10176);
and U11277 (N_11277,N_10395,N_10000);
nand U11278 (N_11278,N_10098,N_10736);
xnor U11279 (N_11279,N_10815,N_10746);
xor U11280 (N_11280,N_10680,N_10764);
nand U11281 (N_11281,N_10864,N_10323);
nand U11282 (N_11282,N_10846,N_10843);
nand U11283 (N_11283,N_10967,N_10860);
and U11284 (N_11284,N_10350,N_10242);
nor U11285 (N_11285,N_10020,N_10465);
and U11286 (N_11286,N_10154,N_10914);
or U11287 (N_11287,N_10410,N_10287);
nand U11288 (N_11288,N_10926,N_10319);
nor U11289 (N_11289,N_10464,N_10615);
nor U11290 (N_11290,N_10251,N_10326);
nor U11291 (N_11291,N_10367,N_10954);
nand U11292 (N_11292,N_10812,N_10845);
xor U11293 (N_11293,N_10390,N_10201);
nand U11294 (N_11294,N_10917,N_10805);
nand U11295 (N_11295,N_10519,N_10023);
or U11296 (N_11296,N_10956,N_10621);
or U11297 (N_11297,N_10298,N_10727);
and U11298 (N_11298,N_10684,N_10146);
and U11299 (N_11299,N_10716,N_10911);
nand U11300 (N_11300,N_10950,N_10200);
xor U11301 (N_11301,N_10314,N_10482);
xnor U11302 (N_11302,N_10939,N_10172);
nand U11303 (N_11303,N_10279,N_10758);
or U11304 (N_11304,N_10622,N_10839);
or U11305 (N_11305,N_10568,N_10423);
or U11306 (N_11306,N_10613,N_10428);
nand U11307 (N_11307,N_10057,N_10292);
or U11308 (N_11308,N_10123,N_10373);
nand U11309 (N_11309,N_10124,N_10009);
nand U11310 (N_11310,N_10313,N_10567);
nand U11311 (N_11311,N_10507,N_10535);
and U11312 (N_11312,N_10502,N_10107);
or U11313 (N_11313,N_10652,N_10461);
xor U11314 (N_11314,N_10271,N_10181);
or U11315 (N_11315,N_10731,N_10881);
xor U11316 (N_11316,N_10641,N_10149);
or U11317 (N_11317,N_10801,N_10422);
xnor U11318 (N_11318,N_10058,N_10002);
or U11319 (N_11319,N_10870,N_10486);
xor U11320 (N_11320,N_10872,N_10466);
xnor U11321 (N_11321,N_10788,N_10581);
xnor U11322 (N_11322,N_10614,N_10305);
and U11323 (N_11323,N_10443,N_10293);
nor U11324 (N_11324,N_10599,N_10480);
nor U11325 (N_11325,N_10935,N_10425);
or U11326 (N_11326,N_10380,N_10222);
nor U11327 (N_11327,N_10041,N_10483);
xnor U11328 (N_11328,N_10402,N_10708);
and U11329 (N_11329,N_10119,N_10477);
nor U11330 (N_11330,N_10601,N_10790);
and U11331 (N_11331,N_10150,N_10528);
nor U11332 (N_11332,N_10370,N_10494);
and U11333 (N_11333,N_10705,N_10884);
or U11334 (N_11334,N_10110,N_10101);
nand U11335 (N_11335,N_10971,N_10932);
xor U11336 (N_11336,N_10501,N_10238);
xor U11337 (N_11337,N_10206,N_10648);
xor U11338 (N_11338,N_10475,N_10162);
nor U11339 (N_11339,N_10548,N_10424);
nand U11340 (N_11340,N_10220,N_10368);
xor U11341 (N_11341,N_10784,N_10439);
nor U11342 (N_11342,N_10192,N_10109);
nand U11343 (N_11343,N_10088,N_10074);
and U11344 (N_11344,N_10847,N_10199);
or U11345 (N_11345,N_10840,N_10521);
or U11346 (N_11346,N_10701,N_10090);
xnor U11347 (N_11347,N_10258,N_10725);
and U11348 (N_11348,N_10817,N_10526);
nor U11349 (N_11349,N_10343,N_10024);
or U11350 (N_11350,N_10334,N_10569);
or U11351 (N_11351,N_10953,N_10793);
xnor U11352 (N_11352,N_10791,N_10252);
and U11353 (N_11353,N_10411,N_10227);
or U11354 (N_11354,N_10899,N_10916);
or U11355 (N_11355,N_10458,N_10851);
nor U11356 (N_11356,N_10908,N_10029);
nand U11357 (N_11357,N_10065,N_10408);
nor U11358 (N_11358,N_10993,N_10702);
or U11359 (N_11359,N_10135,N_10617);
xor U11360 (N_11360,N_10093,N_10543);
nor U11361 (N_11361,N_10175,N_10729);
xnor U11362 (N_11362,N_10080,N_10229);
nor U11363 (N_11363,N_10504,N_10636);
or U11364 (N_11364,N_10321,N_10062);
xnor U11365 (N_11365,N_10442,N_10457);
nand U11366 (N_11366,N_10756,N_10005);
nand U11367 (N_11367,N_10874,N_10525);
and U11368 (N_11368,N_10527,N_10637);
and U11369 (N_11369,N_10738,N_10529);
or U11370 (N_11370,N_10331,N_10039);
xor U11371 (N_11371,N_10066,N_10105);
or U11372 (N_11372,N_10325,N_10972);
and U11373 (N_11373,N_10500,N_10722);
nor U11374 (N_11374,N_10232,N_10356);
xor U11375 (N_11375,N_10397,N_10269);
or U11376 (N_11376,N_10046,N_10924);
and U11377 (N_11377,N_10283,N_10449);
nor U11378 (N_11378,N_10607,N_10518);
and U11379 (N_11379,N_10377,N_10133);
and U11380 (N_11380,N_10512,N_10659);
nand U11381 (N_11381,N_10940,N_10802);
or U11382 (N_11382,N_10290,N_10076);
and U11383 (N_11383,N_10704,N_10148);
or U11384 (N_11384,N_10078,N_10572);
and U11385 (N_11385,N_10263,N_10244);
and U11386 (N_11386,N_10978,N_10912);
xnor U11387 (N_11387,N_10441,N_10070);
xor U11388 (N_11388,N_10138,N_10976);
and U11389 (N_11389,N_10719,N_10530);
and U11390 (N_11390,N_10632,N_10757);
nor U11391 (N_11391,N_10895,N_10118);
nor U11392 (N_11392,N_10897,N_10102);
and U11393 (N_11393,N_10930,N_10517);
xnor U11394 (N_11394,N_10360,N_10726);
nor U11395 (N_11395,N_10883,N_10255);
nor U11396 (N_11396,N_10644,N_10089);
and U11397 (N_11397,N_10602,N_10455);
or U11398 (N_11398,N_10211,N_10996);
and U11399 (N_11399,N_10316,N_10359);
nor U11400 (N_11400,N_10748,N_10215);
and U11401 (N_11401,N_10564,N_10060);
nand U11402 (N_11402,N_10934,N_10371);
or U11403 (N_11403,N_10587,N_10828);
nor U11404 (N_11404,N_10650,N_10253);
and U11405 (N_11405,N_10015,N_10289);
nand U11406 (N_11406,N_10474,N_10054);
or U11407 (N_11407,N_10921,N_10772);
and U11408 (N_11408,N_10348,N_10631);
nor U11409 (N_11409,N_10616,N_10931);
nand U11410 (N_11410,N_10378,N_10082);
nor U11411 (N_11411,N_10103,N_10723);
xnor U11412 (N_11412,N_10053,N_10994);
and U11413 (N_11413,N_10829,N_10664);
nand U11414 (N_11414,N_10031,N_10830);
nand U11415 (N_11415,N_10304,N_10198);
or U11416 (N_11416,N_10469,N_10063);
xor U11417 (N_11417,N_10699,N_10339);
or U11418 (N_11418,N_10844,N_10986);
nor U11419 (N_11419,N_10789,N_10447);
and U11420 (N_11420,N_10087,N_10068);
or U11421 (N_11421,N_10247,N_10379);
or U11422 (N_11422,N_10488,N_10889);
nor U11423 (N_11423,N_10751,N_10796);
nand U11424 (N_11424,N_10661,N_10152);
xnor U11425 (N_11425,N_10759,N_10662);
nor U11426 (N_11426,N_10120,N_10197);
nor U11427 (N_11427,N_10452,N_10037);
or U11428 (N_11428,N_10938,N_10219);
xnor U11429 (N_11429,N_10021,N_10822);
and U11430 (N_11430,N_10027,N_10728);
nor U11431 (N_11431,N_10056,N_10061);
nor U11432 (N_11432,N_10771,N_10776);
nor U11433 (N_11433,N_10724,N_10164);
xor U11434 (N_11434,N_10485,N_10208);
nand U11435 (N_11435,N_10141,N_10945);
nor U11436 (N_11436,N_10275,N_10111);
nor U11437 (N_11437,N_10803,N_10137);
nand U11438 (N_11438,N_10324,N_10214);
or U11439 (N_11439,N_10391,N_10668);
xor U11440 (N_11440,N_10463,N_10004);
nand U11441 (N_11441,N_10479,N_10375);
nor U11442 (N_11442,N_10970,N_10555);
nand U11443 (N_11443,N_10456,N_10920);
nor U11444 (N_11444,N_10170,N_10600);
or U11445 (N_11445,N_10955,N_10625);
nor U11446 (N_11446,N_10913,N_10113);
and U11447 (N_11447,N_10875,N_10703);
or U11448 (N_11448,N_10157,N_10691);
xor U11449 (N_11449,N_10272,N_10554);
and U11450 (N_11450,N_10128,N_10588);
nand U11451 (N_11451,N_10797,N_10571);
xnor U11452 (N_11452,N_10850,N_10354);
nand U11453 (N_11453,N_10403,N_10968);
or U11454 (N_11454,N_10042,N_10858);
or U11455 (N_11455,N_10766,N_10168);
nand U11456 (N_11456,N_10630,N_10929);
nor U11457 (N_11457,N_10139,N_10396);
or U11458 (N_11458,N_10515,N_10740);
or U11459 (N_11459,N_10193,N_10948);
and U11460 (N_11460,N_10596,N_10226);
nor U11461 (N_11461,N_10075,N_10871);
xor U11462 (N_11462,N_10842,N_10861);
and U11463 (N_11463,N_10879,N_10580);
and U11464 (N_11464,N_10810,N_10140);
or U11465 (N_11465,N_10814,N_10721);
nor U11466 (N_11466,N_10777,N_10604);
or U11467 (N_11467,N_10995,N_10687);
nor U11468 (N_11468,N_10052,N_10744);
xor U11469 (N_11469,N_10857,N_10665);
xor U11470 (N_11470,N_10890,N_10437);
and U11471 (N_11471,N_10807,N_10417);
nand U11472 (N_11472,N_10038,N_10570);
and U11473 (N_11473,N_10127,N_10416);
or U11474 (N_11474,N_10589,N_10013);
and U11475 (N_11475,N_10270,N_10942);
or U11476 (N_11476,N_10435,N_10448);
nand U11477 (N_11477,N_10623,N_10574);
or U11478 (N_11478,N_10608,N_10315);
or U11479 (N_11479,N_10880,N_10233);
nand U11480 (N_11480,N_10794,N_10267);
nand U11481 (N_11481,N_10961,N_10694);
nor U11482 (N_11482,N_10532,N_10025);
nand U11483 (N_11483,N_10658,N_10032);
and U11484 (N_11484,N_10898,N_10044);
xor U11485 (N_11485,N_10246,N_10182);
and U11486 (N_11486,N_10952,N_10498);
or U11487 (N_11487,N_10639,N_10492);
nor U11488 (N_11488,N_10225,N_10355);
or U11489 (N_11489,N_10151,N_10669);
nor U11490 (N_11490,N_10509,N_10427);
xor U11491 (N_11491,N_10489,N_10195);
and U11492 (N_11492,N_10404,N_10434);
and U11493 (N_11493,N_10999,N_10357);
nor U11494 (N_11494,N_10414,N_10975);
xnor U11495 (N_11495,N_10392,N_10019);
xnor U11496 (N_11496,N_10106,N_10977);
nor U11497 (N_11497,N_10114,N_10218);
or U11498 (N_11498,N_10240,N_10619);
and U11499 (N_11499,N_10966,N_10806);
xnor U11500 (N_11500,N_10018,N_10436);
and U11501 (N_11501,N_10631,N_10156);
xor U11502 (N_11502,N_10774,N_10893);
or U11503 (N_11503,N_10979,N_10198);
nand U11504 (N_11504,N_10612,N_10975);
nor U11505 (N_11505,N_10254,N_10283);
nand U11506 (N_11506,N_10751,N_10036);
nor U11507 (N_11507,N_10360,N_10106);
and U11508 (N_11508,N_10940,N_10641);
and U11509 (N_11509,N_10655,N_10857);
xor U11510 (N_11510,N_10058,N_10727);
and U11511 (N_11511,N_10382,N_10133);
nand U11512 (N_11512,N_10560,N_10495);
or U11513 (N_11513,N_10306,N_10668);
or U11514 (N_11514,N_10464,N_10531);
nor U11515 (N_11515,N_10221,N_10753);
nor U11516 (N_11516,N_10611,N_10940);
or U11517 (N_11517,N_10131,N_10920);
nand U11518 (N_11518,N_10066,N_10026);
and U11519 (N_11519,N_10488,N_10197);
and U11520 (N_11520,N_10361,N_10624);
nand U11521 (N_11521,N_10722,N_10937);
nor U11522 (N_11522,N_10761,N_10832);
nor U11523 (N_11523,N_10444,N_10369);
nand U11524 (N_11524,N_10435,N_10251);
xor U11525 (N_11525,N_10556,N_10601);
xnor U11526 (N_11526,N_10441,N_10577);
nor U11527 (N_11527,N_10395,N_10835);
nand U11528 (N_11528,N_10280,N_10670);
and U11529 (N_11529,N_10321,N_10013);
nand U11530 (N_11530,N_10047,N_10909);
and U11531 (N_11531,N_10424,N_10453);
and U11532 (N_11532,N_10708,N_10699);
nor U11533 (N_11533,N_10731,N_10648);
nand U11534 (N_11534,N_10168,N_10147);
xor U11535 (N_11535,N_10062,N_10414);
nand U11536 (N_11536,N_10128,N_10063);
xnor U11537 (N_11537,N_10987,N_10686);
xnor U11538 (N_11538,N_10209,N_10467);
and U11539 (N_11539,N_10362,N_10326);
and U11540 (N_11540,N_10881,N_10045);
xor U11541 (N_11541,N_10370,N_10805);
or U11542 (N_11542,N_10901,N_10061);
xor U11543 (N_11543,N_10318,N_10024);
nor U11544 (N_11544,N_10095,N_10674);
xnor U11545 (N_11545,N_10271,N_10865);
and U11546 (N_11546,N_10758,N_10801);
xnor U11547 (N_11547,N_10865,N_10371);
xor U11548 (N_11548,N_10170,N_10647);
nand U11549 (N_11549,N_10963,N_10328);
nor U11550 (N_11550,N_10074,N_10865);
nand U11551 (N_11551,N_10572,N_10363);
nand U11552 (N_11552,N_10966,N_10454);
nor U11553 (N_11553,N_10354,N_10285);
nand U11554 (N_11554,N_10973,N_10570);
or U11555 (N_11555,N_10966,N_10046);
nor U11556 (N_11556,N_10476,N_10693);
nor U11557 (N_11557,N_10916,N_10674);
and U11558 (N_11558,N_10961,N_10925);
nand U11559 (N_11559,N_10387,N_10049);
and U11560 (N_11560,N_10131,N_10345);
and U11561 (N_11561,N_10830,N_10589);
nor U11562 (N_11562,N_10913,N_10914);
xnor U11563 (N_11563,N_10374,N_10534);
and U11564 (N_11564,N_10076,N_10573);
or U11565 (N_11565,N_10466,N_10890);
nor U11566 (N_11566,N_10723,N_10923);
nand U11567 (N_11567,N_10433,N_10249);
or U11568 (N_11568,N_10331,N_10263);
or U11569 (N_11569,N_10430,N_10121);
nor U11570 (N_11570,N_10730,N_10981);
nor U11571 (N_11571,N_10308,N_10973);
and U11572 (N_11572,N_10109,N_10110);
xnor U11573 (N_11573,N_10933,N_10124);
xor U11574 (N_11574,N_10731,N_10094);
xor U11575 (N_11575,N_10241,N_10975);
and U11576 (N_11576,N_10124,N_10449);
and U11577 (N_11577,N_10976,N_10501);
nor U11578 (N_11578,N_10485,N_10851);
xor U11579 (N_11579,N_10712,N_10419);
nor U11580 (N_11580,N_10308,N_10536);
and U11581 (N_11581,N_10325,N_10824);
or U11582 (N_11582,N_10775,N_10758);
nand U11583 (N_11583,N_10436,N_10414);
or U11584 (N_11584,N_10202,N_10491);
nor U11585 (N_11585,N_10760,N_10958);
and U11586 (N_11586,N_10930,N_10724);
nor U11587 (N_11587,N_10355,N_10703);
or U11588 (N_11588,N_10777,N_10504);
nor U11589 (N_11589,N_10243,N_10369);
nand U11590 (N_11590,N_10234,N_10883);
xnor U11591 (N_11591,N_10985,N_10138);
xnor U11592 (N_11592,N_10573,N_10911);
and U11593 (N_11593,N_10799,N_10185);
xnor U11594 (N_11594,N_10916,N_10929);
nor U11595 (N_11595,N_10484,N_10064);
or U11596 (N_11596,N_10944,N_10086);
nor U11597 (N_11597,N_10719,N_10116);
and U11598 (N_11598,N_10134,N_10349);
or U11599 (N_11599,N_10838,N_10869);
or U11600 (N_11600,N_10265,N_10369);
or U11601 (N_11601,N_10481,N_10170);
and U11602 (N_11602,N_10678,N_10238);
nor U11603 (N_11603,N_10056,N_10184);
xor U11604 (N_11604,N_10880,N_10742);
or U11605 (N_11605,N_10019,N_10105);
nand U11606 (N_11606,N_10466,N_10812);
nand U11607 (N_11607,N_10203,N_10258);
or U11608 (N_11608,N_10730,N_10266);
or U11609 (N_11609,N_10340,N_10015);
or U11610 (N_11610,N_10829,N_10133);
nand U11611 (N_11611,N_10989,N_10119);
xnor U11612 (N_11612,N_10542,N_10057);
or U11613 (N_11613,N_10842,N_10426);
and U11614 (N_11614,N_10118,N_10109);
and U11615 (N_11615,N_10869,N_10612);
and U11616 (N_11616,N_10581,N_10922);
nand U11617 (N_11617,N_10089,N_10843);
xnor U11618 (N_11618,N_10621,N_10383);
nor U11619 (N_11619,N_10602,N_10932);
or U11620 (N_11620,N_10830,N_10166);
nand U11621 (N_11621,N_10136,N_10290);
nand U11622 (N_11622,N_10157,N_10550);
xor U11623 (N_11623,N_10960,N_10328);
xnor U11624 (N_11624,N_10596,N_10449);
and U11625 (N_11625,N_10929,N_10396);
or U11626 (N_11626,N_10909,N_10540);
nor U11627 (N_11627,N_10472,N_10023);
and U11628 (N_11628,N_10330,N_10198);
and U11629 (N_11629,N_10206,N_10929);
nor U11630 (N_11630,N_10615,N_10771);
nor U11631 (N_11631,N_10395,N_10694);
xnor U11632 (N_11632,N_10357,N_10560);
xnor U11633 (N_11633,N_10190,N_10896);
nor U11634 (N_11634,N_10163,N_10874);
nand U11635 (N_11635,N_10188,N_10231);
nand U11636 (N_11636,N_10447,N_10699);
or U11637 (N_11637,N_10964,N_10050);
nand U11638 (N_11638,N_10109,N_10513);
or U11639 (N_11639,N_10823,N_10410);
and U11640 (N_11640,N_10592,N_10705);
and U11641 (N_11641,N_10004,N_10084);
or U11642 (N_11642,N_10623,N_10794);
and U11643 (N_11643,N_10477,N_10994);
xor U11644 (N_11644,N_10816,N_10053);
xnor U11645 (N_11645,N_10471,N_10200);
nand U11646 (N_11646,N_10186,N_10181);
and U11647 (N_11647,N_10449,N_10631);
nor U11648 (N_11648,N_10695,N_10903);
nand U11649 (N_11649,N_10481,N_10526);
nor U11650 (N_11650,N_10634,N_10860);
and U11651 (N_11651,N_10721,N_10574);
or U11652 (N_11652,N_10647,N_10341);
nand U11653 (N_11653,N_10809,N_10975);
and U11654 (N_11654,N_10785,N_10330);
xnor U11655 (N_11655,N_10687,N_10307);
or U11656 (N_11656,N_10235,N_10038);
xor U11657 (N_11657,N_10937,N_10592);
xnor U11658 (N_11658,N_10578,N_10291);
xor U11659 (N_11659,N_10982,N_10848);
nor U11660 (N_11660,N_10956,N_10791);
nor U11661 (N_11661,N_10029,N_10352);
xnor U11662 (N_11662,N_10139,N_10003);
nand U11663 (N_11663,N_10065,N_10559);
nor U11664 (N_11664,N_10249,N_10127);
and U11665 (N_11665,N_10395,N_10649);
and U11666 (N_11666,N_10781,N_10307);
xor U11667 (N_11667,N_10081,N_10091);
nand U11668 (N_11668,N_10593,N_10470);
nand U11669 (N_11669,N_10075,N_10910);
xor U11670 (N_11670,N_10160,N_10721);
xor U11671 (N_11671,N_10725,N_10854);
xor U11672 (N_11672,N_10985,N_10304);
nor U11673 (N_11673,N_10238,N_10067);
nand U11674 (N_11674,N_10093,N_10049);
nor U11675 (N_11675,N_10024,N_10465);
xor U11676 (N_11676,N_10448,N_10335);
xor U11677 (N_11677,N_10287,N_10394);
xnor U11678 (N_11678,N_10857,N_10996);
or U11679 (N_11679,N_10044,N_10419);
and U11680 (N_11680,N_10233,N_10279);
nor U11681 (N_11681,N_10788,N_10662);
nor U11682 (N_11682,N_10379,N_10673);
nand U11683 (N_11683,N_10209,N_10099);
and U11684 (N_11684,N_10545,N_10665);
and U11685 (N_11685,N_10837,N_10787);
nor U11686 (N_11686,N_10458,N_10704);
xor U11687 (N_11687,N_10671,N_10990);
and U11688 (N_11688,N_10871,N_10669);
and U11689 (N_11689,N_10022,N_10155);
nand U11690 (N_11690,N_10834,N_10600);
nand U11691 (N_11691,N_10110,N_10246);
and U11692 (N_11692,N_10708,N_10454);
and U11693 (N_11693,N_10308,N_10149);
and U11694 (N_11694,N_10976,N_10565);
and U11695 (N_11695,N_10368,N_10420);
nor U11696 (N_11696,N_10061,N_10894);
and U11697 (N_11697,N_10728,N_10558);
nor U11698 (N_11698,N_10425,N_10006);
nand U11699 (N_11699,N_10883,N_10412);
nor U11700 (N_11700,N_10243,N_10331);
xor U11701 (N_11701,N_10063,N_10575);
nor U11702 (N_11702,N_10898,N_10834);
nand U11703 (N_11703,N_10912,N_10598);
xnor U11704 (N_11704,N_10834,N_10948);
xor U11705 (N_11705,N_10582,N_10014);
xor U11706 (N_11706,N_10651,N_10981);
or U11707 (N_11707,N_10692,N_10016);
and U11708 (N_11708,N_10397,N_10076);
nor U11709 (N_11709,N_10421,N_10204);
and U11710 (N_11710,N_10220,N_10695);
or U11711 (N_11711,N_10188,N_10266);
and U11712 (N_11712,N_10147,N_10183);
nor U11713 (N_11713,N_10375,N_10844);
xor U11714 (N_11714,N_10441,N_10868);
and U11715 (N_11715,N_10162,N_10558);
nor U11716 (N_11716,N_10126,N_10158);
or U11717 (N_11717,N_10689,N_10401);
or U11718 (N_11718,N_10586,N_10433);
nor U11719 (N_11719,N_10622,N_10237);
xor U11720 (N_11720,N_10423,N_10375);
xnor U11721 (N_11721,N_10401,N_10713);
nor U11722 (N_11722,N_10253,N_10256);
or U11723 (N_11723,N_10021,N_10250);
nor U11724 (N_11724,N_10492,N_10975);
nor U11725 (N_11725,N_10379,N_10466);
and U11726 (N_11726,N_10497,N_10568);
xor U11727 (N_11727,N_10338,N_10313);
nand U11728 (N_11728,N_10823,N_10761);
xnor U11729 (N_11729,N_10425,N_10651);
nand U11730 (N_11730,N_10022,N_10935);
nand U11731 (N_11731,N_10018,N_10963);
nand U11732 (N_11732,N_10382,N_10474);
nor U11733 (N_11733,N_10165,N_10420);
or U11734 (N_11734,N_10208,N_10025);
nor U11735 (N_11735,N_10639,N_10419);
nor U11736 (N_11736,N_10976,N_10891);
nor U11737 (N_11737,N_10446,N_10865);
nor U11738 (N_11738,N_10818,N_10300);
nand U11739 (N_11739,N_10517,N_10095);
and U11740 (N_11740,N_10737,N_10661);
and U11741 (N_11741,N_10819,N_10803);
nor U11742 (N_11742,N_10400,N_10791);
nor U11743 (N_11743,N_10030,N_10198);
nand U11744 (N_11744,N_10742,N_10719);
and U11745 (N_11745,N_10533,N_10034);
or U11746 (N_11746,N_10105,N_10713);
or U11747 (N_11747,N_10164,N_10430);
nor U11748 (N_11748,N_10357,N_10832);
xnor U11749 (N_11749,N_10372,N_10306);
nor U11750 (N_11750,N_10734,N_10490);
nand U11751 (N_11751,N_10398,N_10900);
nor U11752 (N_11752,N_10940,N_10400);
nand U11753 (N_11753,N_10936,N_10166);
and U11754 (N_11754,N_10929,N_10000);
nand U11755 (N_11755,N_10086,N_10003);
or U11756 (N_11756,N_10528,N_10518);
xnor U11757 (N_11757,N_10588,N_10858);
nor U11758 (N_11758,N_10254,N_10739);
xor U11759 (N_11759,N_10397,N_10684);
nand U11760 (N_11760,N_10855,N_10845);
nand U11761 (N_11761,N_10272,N_10103);
nand U11762 (N_11762,N_10549,N_10761);
and U11763 (N_11763,N_10310,N_10015);
and U11764 (N_11764,N_10979,N_10850);
nand U11765 (N_11765,N_10102,N_10356);
nand U11766 (N_11766,N_10884,N_10835);
nand U11767 (N_11767,N_10909,N_10892);
or U11768 (N_11768,N_10583,N_10517);
or U11769 (N_11769,N_10086,N_10215);
or U11770 (N_11770,N_10095,N_10629);
nor U11771 (N_11771,N_10692,N_10227);
nor U11772 (N_11772,N_10940,N_10627);
xor U11773 (N_11773,N_10159,N_10953);
xor U11774 (N_11774,N_10403,N_10856);
nor U11775 (N_11775,N_10653,N_10851);
nand U11776 (N_11776,N_10799,N_10488);
and U11777 (N_11777,N_10161,N_10650);
or U11778 (N_11778,N_10252,N_10420);
nor U11779 (N_11779,N_10386,N_10527);
nand U11780 (N_11780,N_10688,N_10785);
and U11781 (N_11781,N_10309,N_10143);
xor U11782 (N_11782,N_10136,N_10949);
and U11783 (N_11783,N_10296,N_10470);
xor U11784 (N_11784,N_10279,N_10781);
xnor U11785 (N_11785,N_10829,N_10419);
nand U11786 (N_11786,N_10881,N_10266);
xnor U11787 (N_11787,N_10994,N_10050);
nor U11788 (N_11788,N_10463,N_10129);
xnor U11789 (N_11789,N_10137,N_10673);
nor U11790 (N_11790,N_10909,N_10577);
or U11791 (N_11791,N_10012,N_10154);
and U11792 (N_11792,N_10773,N_10220);
nor U11793 (N_11793,N_10308,N_10311);
xor U11794 (N_11794,N_10603,N_10982);
nand U11795 (N_11795,N_10160,N_10668);
nand U11796 (N_11796,N_10232,N_10281);
nor U11797 (N_11797,N_10601,N_10399);
nor U11798 (N_11798,N_10839,N_10945);
or U11799 (N_11799,N_10131,N_10589);
and U11800 (N_11800,N_10870,N_10928);
nand U11801 (N_11801,N_10573,N_10225);
nand U11802 (N_11802,N_10177,N_10264);
nand U11803 (N_11803,N_10481,N_10784);
xor U11804 (N_11804,N_10591,N_10244);
nand U11805 (N_11805,N_10797,N_10632);
or U11806 (N_11806,N_10488,N_10727);
and U11807 (N_11807,N_10320,N_10261);
nand U11808 (N_11808,N_10699,N_10052);
and U11809 (N_11809,N_10925,N_10811);
xor U11810 (N_11810,N_10083,N_10505);
or U11811 (N_11811,N_10041,N_10484);
xnor U11812 (N_11812,N_10176,N_10107);
nand U11813 (N_11813,N_10361,N_10993);
nor U11814 (N_11814,N_10654,N_10736);
xnor U11815 (N_11815,N_10610,N_10287);
or U11816 (N_11816,N_10693,N_10859);
and U11817 (N_11817,N_10535,N_10852);
xor U11818 (N_11818,N_10226,N_10327);
and U11819 (N_11819,N_10699,N_10509);
nand U11820 (N_11820,N_10726,N_10933);
and U11821 (N_11821,N_10595,N_10745);
xnor U11822 (N_11822,N_10938,N_10155);
and U11823 (N_11823,N_10708,N_10713);
and U11824 (N_11824,N_10376,N_10369);
nor U11825 (N_11825,N_10024,N_10346);
nand U11826 (N_11826,N_10283,N_10382);
and U11827 (N_11827,N_10101,N_10940);
or U11828 (N_11828,N_10891,N_10419);
xor U11829 (N_11829,N_10529,N_10931);
nor U11830 (N_11830,N_10583,N_10892);
nor U11831 (N_11831,N_10707,N_10597);
and U11832 (N_11832,N_10069,N_10024);
or U11833 (N_11833,N_10185,N_10213);
nand U11834 (N_11834,N_10923,N_10007);
and U11835 (N_11835,N_10448,N_10366);
nand U11836 (N_11836,N_10303,N_10018);
nand U11837 (N_11837,N_10773,N_10208);
nor U11838 (N_11838,N_10880,N_10419);
xor U11839 (N_11839,N_10133,N_10074);
nor U11840 (N_11840,N_10374,N_10642);
and U11841 (N_11841,N_10584,N_10558);
and U11842 (N_11842,N_10413,N_10329);
nand U11843 (N_11843,N_10496,N_10307);
or U11844 (N_11844,N_10237,N_10342);
and U11845 (N_11845,N_10243,N_10277);
or U11846 (N_11846,N_10377,N_10190);
or U11847 (N_11847,N_10471,N_10586);
nand U11848 (N_11848,N_10162,N_10205);
xnor U11849 (N_11849,N_10433,N_10684);
xnor U11850 (N_11850,N_10664,N_10928);
and U11851 (N_11851,N_10052,N_10852);
nand U11852 (N_11852,N_10252,N_10686);
and U11853 (N_11853,N_10315,N_10658);
and U11854 (N_11854,N_10929,N_10578);
and U11855 (N_11855,N_10822,N_10279);
nor U11856 (N_11856,N_10376,N_10694);
nand U11857 (N_11857,N_10694,N_10472);
xnor U11858 (N_11858,N_10046,N_10883);
nand U11859 (N_11859,N_10496,N_10581);
or U11860 (N_11860,N_10999,N_10046);
xor U11861 (N_11861,N_10509,N_10263);
xor U11862 (N_11862,N_10426,N_10047);
and U11863 (N_11863,N_10659,N_10617);
nor U11864 (N_11864,N_10183,N_10201);
nor U11865 (N_11865,N_10074,N_10560);
nor U11866 (N_11866,N_10495,N_10549);
nand U11867 (N_11867,N_10551,N_10614);
nand U11868 (N_11868,N_10561,N_10394);
xnor U11869 (N_11869,N_10808,N_10891);
xor U11870 (N_11870,N_10897,N_10615);
nor U11871 (N_11871,N_10669,N_10623);
nand U11872 (N_11872,N_10856,N_10939);
nand U11873 (N_11873,N_10365,N_10669);
nand U11874 (N_11874,N_10944,N_10397);
nor U11875 (N_11875,N_10674,N_10322);
and U11876 (N_11876,N_10441,N_10873);
and U11877 (N_11877,N_10586,N_10796);
or U11878 (N_11878,N_10793,N_10152);
nor U11879 (N_11879,N_10733,N_10059);
and U11880 (N_11880,N_10370,N_10995);
and U11881 (N_11881,N_10476,N_10456);
nor U11882 (N_11882,N_10472,N_10952);
and U11883 (N_11883,N_10360,N_10787);
and U11884 (N_11884,N_10988,N_10862);
nor U11885 (N_11885,N_10626,N_10898);
xor U11886 (N_11886,N_10137,N_10152);
xor U11887 (N_11887,N_10686,N_10272);
xnor U11888 (N_11888,N_10000,N_10593);
and U11889 (N_11889,N_10121,N_10174);
and U11890 (N_11890,N_10877,N_10411);
or U11891 (N_11891,N_10454,N_10535);
or U11892 (N_11892,N_10526,N_10527);
or U11893 (N_11893,N_10011,N_10115);
or U11894 (N_11894,N_10876,N_10019);
nand U11895 (N_11895,N_10854,N_10163);
and U11896 (N_11896,N_10039,N_10494);
or U11897 (N_11897,N_10988,N_10520);
xnor U11898 (N_11898,N_10827,N_10547);
xnor U11899 (N_11899,N_10854,N_10843);
nand U11900 (N_11900,N_10621,N_10045);
or U11901 (N_11901,N_10405,N_10980);
xor U11902 (N_11902,N_10360,N_10412);
nor U11903 (N_11903,N_10559,N_10119);
xor U11904 (N_11904,N_10521,N_10059);
or U11905 (N_11905,N_10603,N_10541);
nand U11906 (N_11906,N_10658,N_10596);
or U11907 (N_11907,N_10410,N_10079);
nand U11908 (N_11908,N_10102,N_10836);
and U11909 (N_11909,N_10728,N_10555);
and U11910 (N_11910,N_10432,N_10499);
nor U11911 (N_11911,N_10349,N_10051);
and U11912 (N_11912,N_10959,N_10422);
or U11913 (N_11913,N_10638,N_10702);
or U11914 (N_11914,N_10149,N_10073);
nand U11915 (N_11915,N_10047,N_10462);
nor U11916 (N_11916,N_10288,N_10512);
xor U11917 (N_11917,N_10027,N_10076);
and U11918 (N_11918,N_10238,N_10815);
and U11919 (N_11919,N_10358,N_10969);
or U11920 (N_11920,N_10870,N_10802);
and U11921 (N_11921,N_10880,N_10267);
and U11922 (N_11922,N_10085,N_10987);
nand U11923 (N_11923,N_10600,N_10351);
and U11924 (N_11924,N_10129,N_10782);
xnor U11925 (N_11925,N_10210,N_10637);
xor U11926 (N_11926,N_10319,N_10699);
or U11927 (N_11927,N_10560,N_10009);
xnor U11928 (N_11928,N_10165,N_10221);
and U11929 (N_11929,N_10015,N_10720);
nand U11930 (N_11930,N_10343,N_10666);
nand U11931 (N_11931,N_10724,N_10211);
xor U11932 (N_11932,N_10874,N_10403);
xor U11933 (N_11933,N_10088,N_10434);
nor U11934 (N_11934,N_10541,N_10804);
nor U11935 (N_11935,N_10866,N_10763);
or U11936 (N_11936,N_10649,N_10166);
xor U11937 (N_11937,N_10724,N_10955);
xnor U11938 (N_11938,N_10174,N_10291);
nand U11939 (N_11939,N_10687,N_10672);
or U11940 (N_11940,N_10710,N_10101);
xor U11941 (N_11941,N_10356,N_10247);
and U11942 (N_11942,N_10631,N_10900);
nor U11943 (N_11943,N_10558,N_10709);
and U11944 (N_11944,N_10510,N_10222);
or U11945 (N_11945,N_10095,N_10483);
and U11946 (N_11946,N_10845,N_10282);
nor U11947 (N_11947,N_10192,N_10865);
nand U11948 (N_11948,N_10181,N_10711);
and U11949 (N_11949,N_10352,N_10834);
xor U11950 (N_11950,N_10290,N_10851);
nand U11951 (N_11951,N_10123,N_10604);
nor U11952 (N_11952,N_10991,N_10964);
nand U11953 (N_11953,N_10168,N_10673);
and U11954 (N_11954,N_10736,N_10120);
nand U11955 (N_11955,N_10576,N_10261);
and U11956 (N_11956,N_10746,N_10061);
or U11957 (N_11957,N_10893,N_10560);
or U11958 (N_11958,N_10775,N_10048);
or U11959 (N_11959,N_10298,N_10674);
nor U11960 (N_11960,N_10462,N_10510);
nor U11961 (N_11961,N_10917,N_10459);
and U11962 (N_11962,N_10560,N_10218);
and U11963 (N_11963,N_10097,N_10252);
xor U11964 (N_11964,N_10427,N_10807);
or U11965 (N_11965,N_10636,N_10199);
and U11966 (N_11966,N_10688,N_10708);
or U11967 (N_11967,N_10056,N_10169);
nand U11968 (N_11968,N_10232,N_10229);
nand U11969 (N_11969,N_10593,N_10116);
nor U11970 (N_11970,N_10419,N_10389);
nand U11971 (N_11971,N_10891,N_10210);
or U11972 (N_11972,N_10605,N_10451);
nand U11973 (N_11973,N_10657,N_10271);
or U11974 (N_11974,N_10456,N_10460);
and U11975 (N_11975,N_10554,N_10813);
and U11976 (N_11976,N_10733,N_10827);
or U11977 (N_11977,N_10477,N_10239);
xor U11978 (N_11978,N_10774,N_10366);
and U11979 (N_11979,N_10087,N_10631);
nand U11980 (N_11980,N_10847,N_10125);
nor U11981 (N_11981,N_10565,N_10080);
nor U11982 (N_11982,N_10018,N_10257);
nand U11983 (N_11983,N_10484,N_10805);
xor U11984 (N_11984,N_10828,N_10372);
nand U11985 (N_11985,N_10933,N_10688);
xor U11986 (N_11986,N_10951,N_10957);
or U11987 (N_11987,N_10500,N_10188);
or U11988 (N_11988,N_10173,N_10917);
nand U11989 (N_11989,N_10031,N_10953);
or U11990 (N_11990,N_10153,N_10074);
nor U11991 (N_11991,N_10515,N_10159);
nand U11992 (N_11992,N_10033,N_10446);
nor U11993 (N_11993,N_10520,N_10222);
and U11994 (N_11994,N_10649,N_10908);
or U11995 (N_11995,N_10984,N_10165);
or U11996 (N_11996,N_10419,N_10232);
nand U11997 (N_11997,N_10096,N_10086);
or U11998 (N_11998,N_10538,N_10056);
and U11999 (N_11999,N_10341,N_10044);
and U12000 (N_12000,N_11872,N_11244);
nand U12001 (N_12001,N_11590,N_11008);
and U12002 (N_12002,N_11723,N_11205);
or U12003 (N_12003,N_11851,N_11349);
xor U12004 (N_12004,N_11203,N_11280);
and U12005 (N_12005,N_11673,N_11603);
nand U12006 (N_12006,N_11272,N_11730);
or U12007 (N_12007,N_11391,N_11961);
or U12008 (N_12008,N_11147,N_11599);
nand U12009 (N_12009,N_11046,N_11839);
nor U12010 (N_12010,N_11773,N_11345);
nand U12011 (N_12011,N_11464,N_11485);
nand U12012 (N_12012,N_11386,N_11920);
nor U12013 (N_12013,N_11856,N_11829);
and U12014 (N_12014,N_11021,N_11363);
and U12015 (N_12015,N_11939,N_11517);
xor U12016 (N_12016,N_11911,N_11245);
or U12017 (N_12017,N_11806,N_11564);
and U12018 (N_12018,N_11357,N_11395);
nor U12019 (N_12019,N_11107,N_11061);
and U12020 (N_12020,N_11389,N_11569);
or U12021 (N_12021,N_11028,N_11265);
nand U12022 (N_12022,N_11136,N_11071);
nand U12023 (N_12023,N_11956,N_11185);
xnor U12024 (N_12024,N_11001,N_11493);
nor U12025 (N_12025,N_11047,N_11945);
nand U12026 (N_12026,N_11695,N_11063);
nor U12027 (N_12027,N_11354,N_11819);
and U12028 (N_12028,N_11528,N_11159);
nand U12029 (N_12029,N_11764,N_11955);
and U12030 (N_12030,N_11650,N_11216);
and U12031 (N_12031,N_11250,N_11805);
nand U12032 (N_12032,N_11651,N_11770);
nand U12033 (N_12033,N_11288,N_11328);
nand U12034 (N_12034,N_11337,N_11519);
xnor U12035 (N_12035,N_11356,N_11266);
and U12036 (N_12036,N_11030,N_11069);
and U12037 (N_12037,N_11752,N_11290);
nor U12038 (N_12038,N_11885,N_11767);
or U12039 (N_12039,N_11538,N_11375);
or U12040 (N_12040,N_11152,N_11537);
and U12041 (N_12041,N_11463,N_11511);
nor U12042 (N_12042,N_11840,N_11029);
or U12043 (N_12043,N_11551,N_11059);
and U12044 (N_12044,N_11253,N_11714);
xor U12045 (N_12045,N_11527,N_11434);
or U12046 (N_12046,N_11532,N_11378);
xor U12047 (N_12047,N_11148,N_11134);
nand U12048 (N_12048,N_11713,N_11313);
nor U12049 (N_12049,N_11425,N_11957);
or U12050 (N_12050,N_11922,N_11403);
xnor U12051 (N_12051,N_11847,N_11369);
or U12052 (N_12052,N_11346,N_11355);
nor U12053 (N_12053,N_11672,N_11818);
and U12054 (N_12054,N_11643,N_11077);
nand U12055 (N_12055,N_11771,N_11367);
or U12056 (N_12056,N_11499,N_11424);
and U12057 (N_12057,N_11993,N_11645);
nor U12058 (N_12058,N_11082,N_11091);
and U12059 (N_12059,N_11273,N_11379);
xnor U12060 (N_12060,N_11717,N_11814);
xor U12061 (N_12061,N_11711,N_11133);
xor U12062 (N_12062,N_11417,N_11274);
or U12063 (N_12063,N_11854,N_11816);
nor U12064 (N_12064,N_11746,N_11659);
nor U12065 (N_12065,N_11085,N_11325);
nor U12066 (N_12066,N_11906,N_11812);
or U12067 (N_12067,N_11104,N_11276);
or U12068 (N_12068,N_11308,N_11666);
nor U12069 (N_12069,N_11097,N_11687);
nor U12070 (N_12070,N_11234,N_11667);
nand U12071 (N_12071,N_11755,N_11503);
nand U12072 (N_12072,N_11384,N_11896);
and U12073 (N_12073,N_11545,N_11968);
xor U12074 (N_12074,N_11977,N_11583);
xnor U12075 (N_12075,N_11632,N_11292);
and U12076 (N_12076,N_11910,N_11083);
nor U12077 (N_12077,N_11800,N_11581);
and U12078 (N_12078,N_11399,N_11056);
nor U12079 (N_12079,N_11454,N_11963);
xnor U12080 (N_12080,N_11943,N_11795);
xor U12081 (N_12081,N_11743,N_11699);
and U12082 (N_12082,N_11624,N_11033);
or U12083 (N_12083,N_11067,N_11787);
nand U12084 (N_12084,N_11330,N_11591);
and U12085 (N_12085,N_11373,N_11285);
or U12086 (N_12086,N_11988,N_11750);
nand U12087 (N_12087,N_11648,N_11921);
nand U12088 (N_12088,N_11984,N_11326);
xnor U12089 (N_12089,N_11287,N_11210);
xnor U12090 (N_12090,N_11825,N_11408);
and U12091 (N_12091,N_11789,N_11011);
or U12092 (N_12092,N_11846,N_11320);
and U12093 (N_12093,N_11034,N_11735);
nor U12094 (N_12094,N_11170,N_11561);
nor U12095 (N_12095,N_11305,N_11893);
and U12096 (N_12096,N_11683,N_11066);
xnor U12097 (N_12097,N_11641,N_11201);
nor U12098 (N_12098,N_11032,N_11300);
or U12099 (N_12099,N_11881,N_11207);
or U12100 (N_12100,N_11693,N_11451);
and U12101 (N_12101,N_11845,N_11700);
nor U12102 (N_12102,N_11989,N_11453);
and U12103 (N_12103,N_11248,N_11584);
nor U12104 (N_12104,N_11157,N_11677);
nand U12105 (N_12105,N_11361,N_11937);
nand U12106 (N_12106,N_11721,N_11577);
nor U12107 (N_12107,N_11718,N_11169);
xor U12108 (N_12108,N_11226,N_11720);
xnor U12109 (N_12109,N_11359,N_11293);
nand U12110 (N_12110,N_11897,N_11710);
xnor U12111 (N_12111,N_11926,N_11694);
and U12112 (N_12112,N_11663,N_11178);
nor U12113 (N_12113,N_11410,N_11515);
and U12114 (N_12114,N_11394,N_11158);
xnor U12115 (N_12115,N_11332,N_11243);
nand U12116 (N_12116,N_11415,N_11068);
xnor U12117 (N_12117,N_11127,N_11277);
nor U12118 (N_12118,N_11049,N_11540);
or U12119 (N_12119,N_11035,N_11189);
nand U12120 (N_12120,N_11060,N_11702);
xor U12121 (N_12121,N_11242,N_11647);
nor U12122 (N_12122,N_11976,N_11598);
or U12123 (N_12123,N_11882,N_11461);
nor U12124 (N_12124,N_11574,N_11801);
xor U12125 (N_12125,N_11970,N_11421);
and U12126 (N_12126,N_11878,N_11376);
nor U12127 (N_12127,N_11680,N_11655);
nor U12128 (N_12128,N_11283,N_11638);
and U12129 (N_12129,N_11501,N_11240);
and U12130 (N_12130,N_11368,N_11592);
xnor U12131 (N_12131,N_11790,N_11225);
nor U12132 (N_12132,N_11467,N_11270);
xnor U12133 (N_12133,N_11890,N_11826);
nor U12134 (N_12134,N_11558,N_11496);
or U12135 (N_12135,N_11617,N_11549);
nand U12136 (N_12136,N_11252,N_11128);
nor U12137 (N_12137,N_11726,N_11912);
nor U12138 (N_12138,N_11715,N_11324);
or U12139 (N_12139,N_11524,N_11745);
or U12140 (N_12140,N_11102,N_11281);
or U12141 (N_12141,N_11002,N_11442);
nor U12142 (N_12142,N_11748,N_11753);
nand U12143 (N_12143,N_11132,N_11982);
nor U12144 (N_12144,N_11484,N_11843);
nor U12145 (N_12145,N_11015,N_11366);
or U12146 (N_12146,N_11535,N_11181);
and U12147 (N_12147,N_11810,N_11406);
or U12148 (N_12148,N_11541,N_11724);
and U12149 (N_12149,N_11180,N_11914);
or U12150 (N_12150,N_11595,N_11879);
nand U12151 (N_12151,N_11756,N_11975);
nor U12152 (N_12152,N_11448,N_11626);
or U12153 (N_12153,N_11064,N_11803);
nand U12154 (N_12154,N_11338,N_11629);
nand U12155 (N_12155,N_11393,N_11858);
xnor U12156 (N_12156,N_11195,N_11550);
and U12157 (N_12157,N_11855,N_11435);
nor U12158 (N_12158,N_11678,N_11763);
or U12159 (N_12159,N_11747,N_11802);
or U12160 (N_12160,N_11191,N_11336);
or U12161 (N_12161,N_11208,N_11725);
and U12162 (N_12162,N_11352,N_11414);
xor U12163 (N_12163,N_11575,N_11940);
and U12164 (N_12164,N_11076,N_11036);
xnor U12165 (N_12165,N_11705,N_11321);
or U12166 (N_12166,N_11760,N_11960);
or U12167 (N_12167,N_11627,N_11597);
nand U12168 (N_12168,N_11994,N_11441);
xnor U12169 (N_12169,N_11874,N_11062);
nand U12170 (N_12170,N_11606,N_11862);
and U12171 (N_12171,N_11915,N_11864);
nand U12172 (N_12172,N_11635,N_11923);
nand U12173 (N_12173,N_11873,N_11168);
xor U12174 (N_12174,N_11849,N_11539);
xnor U12175 (N_12175,N_11419,N_11155);
nand U12176 (N_12176,N_11114,N_11709);
nor U12177 (N_12177,N_11209,N_11115);
nor U12178 (N_12178,N_11491,N_11218);
nand U12179 (N_12179,N_11072,N_11162);
nand U12180 (N_12180,N_11727,N_11486);
nand U12181 (N_12181,N_11460,N_11222);
nand U12182 (N_12182,N_11190,N_11733);
nor U12183 (N_12183,N_11782,N_11174);
xor U12184 (N_12184,N_11509,N_11712);
and U12185 (N_12185,N_11502,N_11125);
xor U12186 (N_12186,N_11140,N_11654);
nand U12187 (N_12187,N_11951,N_11804);
and U12188 (N_12188,N_11870,N_11224);
nand U12189 (N_12189,N_11553,N_11869);
and U12190 (N_12190,N_11794,N_11098);
and U12191 (N_12191,N_11704,N_11876);
nor U12192 (N_12192,N_11228,N_11738);
nor U12193 (N_12193,N_11172,N_11808);
xnor U12194 (N_12194,N_11865,N_11202);
nand U12195 (N_12195,N_11331,N_11950);
nand U12196 (N_12196,N_11227,N_11311);
nor U12197 (N_12197,N_11439,N_11786);
xor U12198 (N_12198,N_11294,N_11314);
nand U12199 (N_12199,N_11322,N_11859);
and U12200 (N_12200,N_11660,N_11490);
xor U12201 (N_12201,N_11757,N_11057);
and U12202 (N_12202,N_11543,N_11495);
and U12203 (N_12203,N_11684,N_11991);
nor U12204 (N_12204,N_11065,N_11284);
and U12205 (N_12205,N_11883,N_11935);
xnor U12206 (N_12206,N_11165,N_11934);
nor U12207 (N_12207,N_11037,N_11930);
and U12208 (N_12208,N_11438,N_11775);
nand U12209 (N_12209,N_11401,N_11692);
xor U12210 (N_12210,N_11658,N_11100);
and U12211 (N_12211,N_11000,N_11917);
xor U12212 (N_12212,N_11507,N_11898);
and U12213 (N_12213,N_11981,N_11124);
xnor U12214 (N_12214,N_11405,N_11706);
nor U12215 (N_12215,N_11447,N_11536);
xnor U12216 (N_12216,N_11565,N_11618);
nor U12217 (N_12217,N_11488,N_11150);
xnor U12218 (N_12218,N_11559,N_11372);
xnor U12219 (N_12219,N_11520,N_11749);
nor U12220 (N_12220,N_11877,N_11120);
and U12221 (N_12221,N_11580,N_11719);
nand U12222 (N_12222,N_11109,N_11038);
nor U12223 (N_12223,N_11547,N_11867);
and U12224 (N_12224,N_11220,N_11610);
or U12225 (N_12225,N_11099,N_11619);
nor U12226 (N_12226,N_11385,N_11197);
and U12227 (N_12227,N_11026,N_11139);
xnor U12228 (N_12228,N_11301,N_11506);
nand U12229 (N_12229,N_11455,N_11018);
nor U12230 (N_12230,N_11661,N_11716);
xnor U12231 (N_12231,N_11309,N_11237);
or U12232 (N_12232,N_11908,N_11916);
xnor U12233 (N_12233,N_11769,N_11298);
nand U12234 (N_12234,N_11374,N_11249);
xor U12235 (N_12235,N_11048,N_11286);
and U12236 (N_12236,N_11998,N_11531);
and U12237 (N_12237,N_11254,N_11997);
and U12238 (N_12238,N_11430,N_11260);
or U12239 (N_12239,N_11834,N_11831);
xor U12240 (N_12240,N_11974,N_11126);
or U12241 (N_12241,N_11895,N_11668);
nand U12242 (N_12242,N_11087,N_11271);
xnor U12243 (N_12243,N_11089,N_11119);
xnor U12244 (N_12244,N_11918,N_11903);
and U12245 (N_12245,N_11781,N_11303);
nor U12246 (N_12246,N_11341,N_11848);
or U12247 (N_12247,N_11335,N_11798);
nand U12248 (N_12248,N_11353,N_11836);
xnor U12249 (N_12249,N_11010,N_11123);
xnor U12250 (N_12250,N_11154,N_11785);
and U12251 (N_12251,N_11529,N_11871);
or U12252 (N_12252,N_11729,N_11307);
or U12253 (N_12253,N_11736,N_11105);
nand U12254 (N_12254,N_11211,N_11480);
and U12255 (N_12255,N_11092,N_11217);
xor U12256 (N_12256,N_11462,N_11766);
xor U12257 (N_12257,N_11055,N_11156);
and U12258 (N_12258,N_11609,N_11835);
nor U12259 (N_12259,N_11247,N_11508);
xor U12260 (N_12260,N_11437,N_11223);
nand U12261 (N_12261,N_11443,N_11952);
or U12262 (N_12262,N_11116,N_11978);
or U12263 (N_12263,N_11788,N_11143);
or U12264 (N_12264,N_11844,N_11186);
xnor U12265 (N_12265,N_11832,N_11924);
xor U12266 (N_12266,N_11949,N_11929);
nand U12267 (N_12267,N_11996,N_11576);
nand U12268 (N_12268,N_11891,N_11731);
and U12269 (N_12269,N_11296,N_11688);
or U12270 (N_12270,N_11685,N_11167);
xor U12271 (N_12271,N_11212,N_11350);
nand U12272 (N_12272,N_11634,N_11653);
xnor U12273 (N_12273,N_11620,N_11481);
or U12274 (N_12274,N_11809,N_11118);
xor U12275 (N_12275,N_11475,N_11964);
xnor U12276 (N_12276,N_11941,N_11504);
and U12277 (N_12277,N_11090,N_11302);
and U12278 (N_12278,N_11075,N_11039);
nor U12279 (N_12279,N_11566,N_11103);
and U12280 (N_12280,N_11432,N_11518);
xnor U12281 (N_12281,N_11382,N_11639);
or U12282 (N_12282,N_11830,N_11416);
xnor U12283 (N_12283,N_11214,N_11774);
nand U12284 (N_12284,N_11777,N_11776);
and U12285 (N_12285,N_11404,N_11426);
xnor U12286 (N_12286,N_11476,N_11841);
nand U12287 (N_12287,N_11004,N_11675);
nand U12288 (N_12288,N_11458,N_11027);
nand U12289 (N_12289,N_11446,N_11636);
nor U12290 (N_12290,N_11081,N_11479);
or U12291 (N_12291,N_11999,N_11135);
and U12292 (N_12292,N_11608,N_11691);
nand U12293 (N_12293,N_11070,N_11884);
or U12294 (N_12294,N_11698,N_11602);
or U12295 (N_12295,N_11852,N_11122);
and U12296 (N_12296,N_11477,N_11947);
nand U12297 (N_12297,N_11074,N_11837);
nor U12298 (N_12298,N_11986,N_11251);
or U12299 (N_12299,N_11728,N_11433);
nand U12300 (N_12300,N_11958,N_11969);
or U12301 (N_12301,N_11907,N_11182);
or U12302 (N_12302,N_11235,N_11542);
and U12303 (N_12303,N_11058,N_11739);
nand U12304 (N_12304,N_11701,N_11533);
and U12305 (N_12305,N_11633,N_11187);
xnor U12306 (N_12306,N_11622,N_11875);
or U12307 (N_12307,N_11390,N_11343);
xnor U12308 (N_12308,N_11315,N_11412);
and U12309 (N_12309,N_11567,N_11452);
nor U12310 (N_12310,N_11646,N_11319);
nor U12311 (N_12311,N_11498,N_11887);
and U12312 (N_12312,N_11005,N_11556);
or U12313 (N_12313,N_11588,N_11006);
nand U12314 (N_12314,N_11664,N_11409);
or U12315 (N_12315,N_11101,N_11644);
xnor U12316 (N_12316,N_11175,N_11177);
nand U12317 (N_12317,N_11465,N_11990);
and U12318 (N_12318,N_11073,N_11823);
xnor U12319 (N_12319,N_11557,N_11043);
nor U12320 (N_12320,N_11258,N_11050);
nor U12321 (N_12321,N_11817,N_11649);
xnor U12322 (N_12322,N_11051,N_11526);
and U12323 (N_12323,N_11094,N_11045);
xor U12324 (N_12324,N_11267,N_11793);
and U12325 (N_12325,N_11861,N_11933);
nor U12326 (N_12326,N_11340,N_11173);
nor U12327 (N_12327,N_11612,N_11522);
and U12328 (N_12328,N_11899,N_11842);
xnor U12329 (N_12329,N_11967,N_11402);
nor U12330 (N_12330,N_11546,N_11054);
or U12331 (N_12331,N_11973,N_11192);
or U12332 (N_12332,N_11144,N_11261);
and U12333 (N_12333,N_11052,N_11780);
and U12334 (N_12334,N_11820,N_11388);
nand U12335 (N_12335,N_11257,N_11894);
nand U12336 (N_12336,N_11469,N_11722);
nor U12337 (N_12337,N_11450,N_11329);
nor U12338 (N_12338,N_11003,N_11176);
nand U12339 (N_12339,N_11928,N_11640);
xor U12340 (N_12340,N_11734,N_11482);
nor U12341 (N_12341,N_11523,N_11605);
nor U12342 (N_12342,N_11231,N_11980);
and U12343 (N_12343,N_11679,N_11936);
nor U12344 (N_12344,N_11621,N_11505);
or U12345 (N_12345,N_11512,N_11637);
xor U12346 (N_12346,N_11901,N_11616);
or U12347 (N_12347,N_11615,N_11886);
or U12348 (N_12348,N_11164,N_11431);
or U12349 (N_12349,N_11611,N_11323);
nor U12350 (N_12350,N_11084,N_11457);
or U12351 (N_12351,N_11239,N_11444);
xor U12352 (N_12352,N_11111,N_11470);
or U12353 (N_12353,N_11765,N_11579);
or U12354 (N_12354,N_11241,N_11304);
or U12355 (N_12355,N_11860,N_11044);
xor U12356 (N_12356,N_11657,N_11909);
nor U12357 (N_12357,N_11427,N_11117);
or U12358 (N_12358,N_11573,N_11696);
nor U12359 (N_12359,N_11088,N_11925);
and U12360 (N_12360,N_11863,N_11166);
nand U12361 (N_12361,N_11282,N_11138);
or U12362 (N_12362,N_11630,N_11510);
or U12363 (N_12363,N_11295,N_11853);
and U12364 (N_12364,N_11703,N_11024);
xor U12365 (N_12365,N_11113,N_11671);
or U12366 (N_12366,N_11022,N_11797);
and U12367 (N_12367,N_11179,N_11656);
nand U12368 (N_12368,N_11291,N_11857);
nand U12369 (N_12369,N_11023,N_11779);
or U12370 (N_12370,N_11472,N_11578);
xor U12371 (N_12371,N_11613,N_11707);
nand U12372 (N_12372,N_11585,N_11279);
xor U12373 (N_12373,N_11108,N_11146);
and U12374 (N_12374,N_11262,N_11031);
xnor U12375 (N_12375,N_11530,N_11310);
xor U12376 (N_12376,N_11106,N_11318);
nor U12377 (N_12377,N_11697,N_11768);
nand U12378 (N_12378,N_11130,N_11041);
nand U12379 (N_12379,N_11783,N_11161);
nand U12380 (N_12380,N_11880,N_11708);
nand U12381 (N_12381,N_11327,N_11900);
nand U12382 (N_12382,N_11418,N_11784);
and U12383 (N_12383,N_11778,N_11473);
nor U12384 (N_12384,N_11468,N_11459);
and U12385 (N_12385,N_11607,N_11919);
and U12386 (N_12386,N_11387,N_11948);
nand U12387 (N_12387,N_11555,N_11669);
nand U12388 (N_12388,N_11944,N_11121);
nand U12389 (N_12389,N_11759,N_11019);
nand U12390 (N_12390,N_11625,N_11850);
xor U12391 (N_12391,N_11219,N_11489);
and U12392 (N_12392,N_11312,N_11815);
xor U12393 (N_12393,N_11079,N_11586);
xor U12394 (N_12394,N_11020,N_11892);
or U12395 (N_12395,N_11392,N_11971);
nor U12396 (N_12396,N_11601,N_11364);
nor U12397 (N_12397,N_11306,N_11396);
xnor U12398 (N_12398,N_11013,N_11194);
or U12399 (N_12399,N_11381,N_11487);
nand U12400 (N_12400,N_11563,N_11631);
nand U12401 (N_12401,N_11799,N_11268);
nand U12402 (N_12402,N_11946,N_11992);
and U12403 (N_12403,N_11256,N_11571);
nor U12404 (N_12404,N_11966,N_11959);
nor U12405 (N_12405,N_11428,N_11772);
xnor U12406 (N_12406,N_11979,N_11289);
xor U12407 (N_12407,N_11149,N_11525);
nand U12408 (N_12408,N_11398,N_11492);
or U12409 (N_12409,N_11362,N_11741);
xor U12410 (N_12410,N_11014,N_11017);
nand U12411 (N_12411,N_11686,N_11811);
or U12412 (N_12412,N_11927,N_11889);
nor U12413 (N_12413,N_11316,N_11552);
nand U12414 (N_12414,N_11954,N_11593);
xnor U12415 (N_12415,N_11429,N_11131);
or U12416 (N_12416,N_11740,N_11995);
or U12417 (N_12417,N_11371,N_11317);
xor U12418 (N_12418,N_11744,N_11652);
nor U12419 (N_12419,N_11297,N_11278);
and U12420 (N_12420,N_11184,N_11230);
nand U12421 (N_12421,N_11568,N_11931);
nand U12422 (N_12422,N_11737,N_11813);
or U12423 (N_12423,N_11348,N_11436);
xnor U12424 (N_12424,N_11093,N_11440);
or U12425 (N_12425,N_11080,N_11344);
and U12426 (N_12426,N_11095,N_11497);
and U12427 (N_12427,N_11420,N_11534);
nor U12428 (N_12428,N_11333,N_11681);
xnor U12429 (N_12429,N_11263,N_11690);
nor U12430 (N_12430,N_11662,N_11141);
or U12431 (N_12431,N_11380,N_11972);
nand U12432 (N_12432,N_11942,N_11423);
nor U12433 (N_12433,N_11962,N_11953);
xor U12434 (N_12434,N_11642,N_11232);
or U12435 (N_12435,N_11163,N_11902);
nand U12436 (N_12436,N_11792,N_11255);
xor U12437 (N_12437,N_11665,N_11078);
nor U12438 (N_12438,N_11670,N_11236);
xor U12439 (N_12439,N_11012,N_11449);
and U12440 (N_12440,N_11360,N_11516);
or U12441 (N_12441,N_11456,N_11086);
nor U12442 (N_12442,N_11246,N_11965);
or U12443 (N_12443,N_11016,N_11594);
and U12444 (N_12444,N_11833,N_11985);
or U12445 (N_12445,N_11151,N_11042);
xor U12446 (N_12446,N_11758,N_11587);
and U12447 (N_12447,N_11838,N_11200);
nor U12448 (N_12448,N_11589,N_11269);
or U12449 (N_12449,N_11213,N_11562);
nor U12450 (N_12450,N_11025,N_11888);
nor U12451 (N_12451,N_11938,N_11183);
and U12452 (N_12452,N_11521,N_11275);
nand U12453 (N_12453,N_11761,N_11827);
nor U12454 (N_12454,N_11824,N_11142);
xnor U12455 (N_12455,N_11623,N_11342);
nand U12456 (N_12456,N_11264,N_11596);
nor U12457 (N_12457,N_11198,N_11233);
nor U12458 (N_12458,N_11370,N_11096);
or U12459 (N_12459,N_11751,N_11299);
xor U12460 (N_12460,N_11193,N_11110);
or U12461 (N_12461,N_11215,N_11600);
nor U12462 (N_12462,N_11196,N_11732);
xor U12463 (N_12463,N_11572,N_11238);
nor U12464 (N_12464,N_11112,N_11137);
nand U12465 (N_12465,N_11494,N_11483);
and U12466 (N_12466,N_11500,N_11007);
xnor U12467 (N_12467,N_11221,N_11513);
nand U12468 (N_12468,N_11474,N_11570);
and U12469 (N_12469,N_11614,N_11742);
or U12470 (N_12470,N_11791,N_11868);
and U12471 (N_12471,N_11628,N_11822);
nand U12472 (N_12472,N_11582,N_11204);
and U12473 (N_12473,N_11471,N_11411);
or U12474 (N_12474,N_11905,N_11754);
nor U12475 (N_12475,N_11548,N_11674);
and U12476 (N_12476,N_11229,N_11358);
or U12477 (N_12477,N_11383,N_11604);
xor U12478 (N_12478,N_11544,N_11554);
nor U12479 (N_12479,N_11009,N_11807);
or U12480 (N_12480,N_11259,N_11206);
and U12481 (N_12481,N_11478,N_11040);
or U12482 (N_12482,N_11377,N_11400);
and U12483 (N_12483,N_11560,N_11983);
nor U12484 (N_12484,N_11689,N_11351);
or U12485 (N_12485,N_11413,N_11129);
xnor U12486 (N_12486,N_11199,N_11762);
nor U12487 (N_12487,N_11188,N_11407);
or U12488 (N_12488,N_11365,N_11913);
xnor U12489 (N_12489,N_11682,N_11466);
or U12490 (N_12490,N_11866,N_11987);
or U12491 (N_12491,N_11153,N_11904);
nor U12492 (N_12492,N_11397,N_11160);
and U12493 (N_12493,N_11828,N_11676);
nor U12494 (N_12494,N_11422,N_11514);
nor U12495 (N_12495,N_11821,N_11334);
nand U12496 (N_12496,N_11171,N_11347);
or U12497 (N_12497,N_11932,N_11053);
xor U12498 (N_12498,N_11145,N_11339);
nand U12499 (N_12499,N_11445,N_11796);
or U12500 (N_12500,N_11673,N_11554);
xnor U12501 (N_12501,N_11873,N_11867);
or U12502 (N_12502,N_11196,N_11014);
xor U12503 (N_12503,N_11206,N_11433);
or U12504 (N_12504,N_11505,N_11813);
and U12505 (N_12505,N_11489,N_11539);
nor U12506 (N_12506,N_11626,N_11949);
nand U12507 (N_12507,N_11800,N_11773);
nand U12508 (N_12508,N_11779,N_11529);
and U12509 (N_12509,N_11704,N_11384);
or U12510 (N_12510,N_11988,N_11809);
and U12511 (N_12511,N_11078,N_11800);
or U12512 (N_12512,N_11352,N_11308);
or U12513 (N_12513,N_11825,N_11945);
xnor U12514 (N_12514,N_11541,N_11885);
nor U12515 (N_12515,N_11141,N_11925);
nor U12516 (N_12516,N_11740,N_11874);
or U12517 (N_12517,N_11730,N_11858);
xor U12518 (N_12518,N_11179,N_11852);
or U12519 (N_12519,N_11774,N_11014);
nor U12520 (N_12520,N_11199,N_11951);
xnor U12521 (N_12521,N_11342,N_11445);
nor U12522 (N_12522,N_11252,N_11464);
and U12523 (N_12523,N_11414,N_11695);
or U12524 (N_12524,N_11698,N_11907);
nand U12525 (N_12525,N_11125,N_11371);
or U12526 (N_12526,N_11742,N_11404);
xor U12527 (N_12527,N_11783,N_11326);
nor U12528 (N_12528,N_11345,N_11916);
or U12529 (N_12529,N_11872,N_11854);
nand U12530 (N_12530,N_11308,N_11529);
nor U12531 (N_12531,N_11691,N_11578);
nand U12532 (N_12532,N_11760,N_11284);
and U12533 (N_12533,N_11456,N_11297);
or U12534 (N_12534,N_11242,N_11562);
nand U12535 (N_12535,N_11763,N_11975);
or U12536 (N_12536,N_11942,N_11438);
nand U12537 (N_12537,N_11528,N_11185);
and U12538 (N_12538,N_11526,N_11264);
nor U12539 (N_12539,N_11161,N_11490);
or U12540 (N_12540,N_11177,N_11016);
nand U12541 (N_12541,N_11687,N_11406);
xor U12542 (N_12542,N_11489,N_11977);
and U12543 (N_12543,N_11776,N_11486);
and U12544 (N_12544,N_11605,N_11220);
nand U12545 (N_12545,N_11781,N_11871);
nand U12546 (N_12546,N_11463,N_11352);
and U12547 (N_12547,N_11049,N_11581);
and U12548 (N_12548,N_11065,N_11210);
nand U12549 (N_12549,N_11633,N_11049);
nor U12550 (N_12550,N_11833,N_11265);
xor U12551 (N_12551,N_11770,N_11631);
nand U12552 (N_12552,N_11679,N_11881);
xnor U12553 (N_12553,N_11694,N_11155);
xor U12554 (N_12554,N_11280,N_11644);
nor U12555 (N_12555,N_11153,N_11099);
nor U12556 (N_12556,N_11239,N_11866);
xnor U12557 (N_12557,N_11373,N_11081);
nand U12558 (N_12558,N_11118,N_11973);
and U12559 (N_12559,N_11419,N_11963);
and U12560 (N_12560,N_11081,N_11228);
nand U12561 (N_12561,N_11921,N_11238);
nand U12562 (N_12562,N_11250,N_11133);
xnor U12563 (N_12563,N_11908,N_11628);
nand U12564 (N_12564,N_11163,N_11314);
nand U12565 (N_12565,N_11140,N_11583);
nand U12566 (N_12566,N_11377,N_11569);
nor U12567 (N_12567,N_11208,N_11660);
nand U12568 (N_12568,N_11147,N_11503);
or U12569 (N_12569,N_11668,N_11922);
nand U12570 (N_12570,N_11559,N_11622);
nand U12571 (N_12571,N_11184,N_11905);
xnor U12572 (N_12572,N_11553,N_11852);
nand U12573 (N_12573,N_11458,N_11804);
and U12574 (N_12574,N_11218,N_11527);
nor U12575 (N_12575,N_11057,N_11006);
xor U12576 (N_12576,N_11373,N_11087);
and U12577 (N_12577,N_11911,N_11235);
xor U12578 (N_12578,N_11175,N_11499);
and U12579 (N_12579,N_11291,N_11333);
and U12580 (N_12580,N_11113,N_11726);
nor U12581 (N_12581,N_11998,N_11804);
and U12582 (N_12582,N_11017,N_11565);
nand U12583 (N_12583,N_11965,N_11432);
nor U12584 (N_12584,N_11638,N_11440);
or U12585 (N_12585,N_11794,N_11904);
and U12586 (N_12586,N_11008,N_11030);
xor U12587 (N_12587,N_11324,N_11714);
and U12588 (N_12588,N_11844,N_11660);
and U12589 (N_12589,N_11958,N_11598);
nor U12590 (N_12590,N_11940,N_11450);
or U12591 (N_12591,N_11997,N_11571);
xor U12592 (N_12592,N_11705,N_11741);
nor U12593 (N_12593,N_11264,N_11927);
or U12594 (N_12594,N_11245,N_11243);
nand U12595 (N_12595,N_11798,N_11877);
nand U12596 (N_12596,N_11698,N_11010);
or U12597 (N_12597,N_11057,N_11026);
and U12598 (N_12598,N_11667,N_11826);
xnor U12599 (N_12599,N_11050,N_11971);
or U12600 (N_12600,N_11923,N_11273);
or U12601 (N_12601,N_11770,N_11152);
nand U12602 (N_12602,N_11559,N_11146);
or U12603 (N_12603,N_11757,N_11471);
nand U12604 (N_12604,N_11755,N_11361);
or U12605 (N_12605,N_11050,N_11466);
and U12606 (N_12606,N_11700,N_11685);
nand U12607 (N_12607,N_11125,N_11192);
and U12608 (N_12608,N_11536,N_11020);
or U12609 (N_12609,N_11867,N_11866);
nand U12610 (N_12610,N_11374,N_11719);
nand U12611 (N_12611,N_11126,N_11021);
and U12612 (N_12612,N_11750,N_11164);
nand U12613 (N_12613,N_11078,N_11140);
nand U12614 (N_12614,N_11102,N_11341);
xnor U12615 (N_12615,N_11574,N_11670);
xor U12616 (N_12616,N_11294,N_11714);
and U12617 (N_12617,N_11541,N_11550);
nand U12618 (N_12618,N_11237,N_11842);
and U12619 (N_12619,N_11956,N_11443);
xnor U12620 (N_12620,N_11050,N_11485);
or U12621 (N_12621,N_11674,N_11157);
nand U12622 (N_12622,N_11671,N_11555);
nor U12623 (N_12623,N_11816,N_11788);
xor U12624 (N_12624,N_11170,N_11891);
nor U12625 (N_12625,N_11026,N_11849);
nor U12626 (N_12626,N_11408,N_11744);
or U12627 (N_12627,N_11739,N_11391);
or U12628 (N_12628,N_11624,N_11752);
nand U12629 (N_12629,N_11522,N_11693);
nand U12630 (N_12630,N_11000,N_11939);
xor U12631 (N_12631,N_11516,N_11839);
xnor U12632 (N_12632,N_11964,N_11713);
or U12633 (N_12633,N_11983,N_11442);
xnor U12634 (N_12634,N_11776,N_11915);
or U12635 (N_12635,N_11356,N_11749);
or U12636 (N_12636,N_11118,N_11327);
xnor U12637 (N_12637,N_11752,N_11394);
or U12638 (N_12638,N_11300,N_11067);
xnor U12639 (N_12639,N_11931,N_11574);
xnor U12640 (N_12640,N_11897,N_11589);
nor U12641 (N_12641,N_11885,N_11817);
and U12642 (N_12642,N_11228,N_11213);
nor U12643 (N_12643,N_11360,N_11159);
nor U12644 (N_12644,N_11221,N_11726);
nor U12645 (N_12645,N_11693,N_11564);
nor U12646 (N_12646,N_11486,N_11711);
nor U12647 (N_12647,N_11202,N_11150);
or U12648 (N_12648,N_11730,N_11560);
nand U12649 (N_12649,N_11643,N_11900);
or U12650 (N_12650,N_11212,N_11279);
xnor U12651 (N_12651,N_11821,N_11288);
or U12652 (N_12652,N_11230,N_11180);
nand U12653 (N_12653,N_11746,N_11965);
xnor U12654 (N_12654,N_11881,N_11393);
and U12655 (N_12655,N_11389,N_11442);
or U12656 (N_12656,N_11377,N_11592);
or U12657 (N_12657,N_11382,N_11795);
nand U12658 (N_12658,N_11295,N_11815);
xor U12659 (N_12659,N_11495,N_11316);
or U12660 (N_12660,N_11172,N_11099);
or U12661 (N_12661,N_11540,N_11521);
xnor U12662 (N_12662,N_11452,N_11088);
xor U12663 (N_12663,N_11083,N_11232);
xnor U12664 (N_12664,N_11830,N_11797);
xor U12665 (N_12665,N_11204,N_11626);
xnor U12666 (N_12666,N_11562,N_11472);
and U12667 (N_12667,N_11927,N_11342);
or U12668 (N_12668,N_11025,N_11208);
xnor U12669 (N_12669,N_11871,N_11055);
or U12670 (N_12670,N_11351,N_11253);
nand U12671 (N_12671,N_11922,N_11690);
and U12672 (N_12672,N_11681,N_11215);
nand U12673 (N_12673,N_11426,N_11548);
or U12674 (N_12674,N_11867,N_11362);
nand U12675 (N_12675,N_11346,N_11070);
and U12676 (N_12676,N_11933,N_11182);
and U12677 (N_12677,N_11841,N_11496);
xor U12678 (N_12678,N_11280,N_11212);
nand U12679 (N_12679,N_11861,N_11896);
or U12680 (N_12680,N_11321,N_11367);
nor U12681 (N_12681,N_11644,N_11844);
and U12682 (N_12682,N_11558,N_11822);
xnor U12683 (N_12683,N_11238,N_11114);
or U12684 (N_12684,N_11974,N_11666);
nor U12685 (N_12685,N_11513,N_11422);
or U12686 (N_12686,N_11010,N_11306);
xor U12687 (N_12687,N_11425,N_11833);
nor U12688 (N_12688,N_11303,N_11125);
xor U12689 (N_12689,N_11378,N_11660);
and U12690 (N_12690,N_11873,N_11063);
nand U12691 (N_12691,N_11258,N_11715);
nor U12692 (N_12692,N_11615,N_11839);
nand U12693 (N_12693,N_11364,N_11411);
xor U12694 (N_12694,N_11070,N_11851);
and U12695 (N_12695,N_11437,N_11828);
nand U12696 (N_12696,N_11602,N_11610);
xor U12697 (N_12697,N_11367,N_11981);
and U12698 (N_12698,N_11325,N_11987);
and U12699 (N_12699,N_11084,N_11802);
and U12700 (N_12700,N_11163,N_11524);
xor U12701 (N_12701,N_11350,N_11494);
xnor U12702 (N_12702,N_11945,N_11401);
nand U12703 (N_12703,N_11527,N_11859);
or U12704 (N_12704,N_11890,N_11717);
xnor U12705 (N_12705,N_11652,N_11906);
nor U12706 (N_12706,N_11076,N_11349);
or U12707 (N_12707,N_11771,N_11745);
nand U12708 (N_12708,N_11285,N_11275);
and U12709 (N_12709,N_11672,N_11355);
nor U12710 (N_12710,N_11165,N_11249);
nand U12711 (N_12711,N_11889,N_11084);
xor U12712 (N_12712,N_11769,N_11936);
nand U12713 (N_12713,N_11530,N_11250);
or U12714 (N_12714,N_11386,N_11108);
or U12715 (N_12715,N_11500,N_11290);
and U12716 (N_12716,N_11772,N_11781);
nor U12717 (N_12717,N_11572,N_11321);
xor U12718 (N_12718,N_11345,N_11870);
xnor U12719 (N_12719,N_11044,N_11859);
nor U12720 (N_12720,N_11418,N_11765);
or U12721 (N_12721,N_11126,N_11206);
nand U12722 (N_12722,N_11341,N_11277);
and U12723 (N_12723,N_11151,N_11870);
xnor U12724 (N_12724,N_11544,N_11337);
xnor U12725 (N_12725,N_11723,N_11683);
xor U12726 (N_12726,N_11068,N_11302);
nand U12727 (N_12727,N_11843,N_11381);
nand U12728 (N_12728,N_11822,N_11409);
xnor U12729 (N_12729,N_11758,N_11473);
or U12730 (N_12730,N_11860,N_11322);
xnor U12731 (N_12731,N_11416,N_11716);
or U12732 (N_12732,N_11436,N_11468);
and U12733 (N_12733,N_11366,N_11170);
xnor U12734 (N_12734,N_11395,N_11946);
or U12735 (N_12735,N_11425,N_11826);
nand U12736 (N_12736,N_11266,N_11668);
nand U12737 (N_12737,N_11466,N_11699);
and U12738 (N_12738,N_11885,N_11594);
nand U12739 (N_12739,N_11068,N_11175);
nand U12740 (N_12740,N_11106,N_11039);
nand U12741 (N_12741,N_11967,N_11613);
nor U12742 (N_12742,N_11144,N_11609);
nor U12743 (N_12743,N_11507,N_11310);
nor U12744 (N_12744,N_11370,N_11134);
or U12745 (N_12745,N_11030,N_11501);
and U12746 (N_12746,N_11759,N_11760);
and U12747 (N_12747,N_11255,N_11171);
xnor U12748 (N_12748,N_11209,N_11977);
xnor U12749 (N_12749,N_11884,N_11663);
xor U12750 (N_12750,N_11987,N_11944);
and U12751 (N_12751,N_11561,N_11798);
nand U12752 (N_12752,N_11758,N_11491);
nor U12753 (N_12753,N_11522,N_11361);
xnor U12754 (N_12754,N_11402,N_11516);
nand U12755 (N_12755,N_11287,N_11897);
nor U12756 (N_12756,N_11931,N_11915);
nand U12757 (N_12757,N_11730,N_11105);
nor U12758 (N_12758,N_11392,N_11110);
xnor U12759 (N_12759,N_11149,N_11493);
and U12760 (N_12760,N_11597,N_11853);
xor U12761 (N_12761,N_11805,N_11241);
nand U12762 (N_12762,N_11378,N_11548);
nand U12763 (N_12763,N_11028,N_11494);
nor U12764 (N_12764,N_11712,N_11627);
xor U12765 (N_12765,N_11048,N_11161);
xor U12766 (N_12766,N_11429,N_11243);
and U12767 (N_12767,N_11023,N_11657);
xnor U12768 (N_12768,N_11697,N_11948);
nor U12769 (N_12769,N_11047,N_11701);
xor U12770 (N_12770,N_11855,N_11119);
nor U12771 (N_12771,N_11779,N_11950);
nand U12772 (N_12772,N_11273,N_11478);
nand U12773 (N_12773,N_11820,N_11095);
nand U12774 (N_12774,N_11212,N_11592);
nor U12775 (N_12775,N_11908,N_11324);
xnor U12776 (N_12776,N_11099,N_11395);
nand U12777 (N_12777,N_11603,N_11695);
xnor U12778 (N_12778,N_11052,N_11194);
nor U12779 (N_12779,N_11090,N_11537);
nor U12780 (N_12780,N_11709,N_11175);
nand U12781 (N_12781,N_11198,N_11427);
and U12782 (N_12782,N_11521,N_11084);
or U12783 (N_12783,N_11963,N_11733);
nand U12784 (N_12784,N_11773,N_11842);
xor U12785 (N_12785,N_11898,N_11618);
or U12786 (N_12786,N_11193,N_11257);
nor U12787 (N_12787,N_11527,N_11946);
and U12788 (N_12788,N_11698,N_11898);
nand U12789 (N_12789,N_11295,N_11086);
nor U12790 (N_12790,N_11689,N_11743);
xnor U12791 (N_12791,N_11757,N_11193);
xor U12792 (N_12792,N_11716,N_11288);
nand U12793 (N_12793,N_11452,N_11476);
or U12794 (N_12794,N_11663,N_11945);
nor U12795 (N_12795,N_11795,N_11836);
xor U12796 (N_12796,N_11252,N_11763);
or U12797 (N_12797,N_11549,N_11357);
and U12798 (N_12798,N_11915,N_11817);
and U12799 (N_12799,N_11895,N_11216);
and U12800 (N_12800,N_11442,N_11780);
nor U12801 (N_12801,N_11211,N_11200);
nand U12802 (N_12802,N_11789,N_11367);
nor U12803 (N_12803,N_11089,N_11298);
or U12804 (N_12804,N_11777,N_11444);
nand U12805 (N_12805,N_11844,N_11892);
and U12806 (N_12806,N_11850,N_11484);
and U12807 (N_12807,N_11003,N_11450);
nor U12808 (N_12808,N_11394,N_11478);
xnor U12809 (N_12809,N_11286,N_11431);
nor U12810 (N_12810,N_11302,N_11607);
and U12811 (N_12811,N_11208,N_11195);
nand U12812 (N_12812,N_11132,N_11189);
nand U12813 (N_12813,N_11059,N_11508);
or U12814 (N_12814,N_11645,N_11041);
nand U12815 (N_12815,N_11031,N_11329);
nor U12816 (N_12816,N_11510,N_11956);
and U12817 (N_12817,N_11005,N_11331);
nor U12818 (N_12818,N_11591,N_11220);
xnor U12819 (N_12819,N_11852,N_11487);
nor U12820 (N_12820,N_11911,N_11593);
xnor U12821 (N_12821,N_11777,N_11787);
nor U12822 (N_12822,N_11811,N_11172);
nand U12823 (N_12823,N_11187,N_11190);
or U12824 (N_12824,N_11298,N_11627);
xor U12825 (N_12825,N_11520,N_11668);
or U12826 (N_12826,N_11973,N_11255);
or U12827 (N_12827,N_11984,N_11423);
nor U12828 (N_12828,N_11112,N_11735);
or U12829 (N_12829,N_11597,N_11100);
or U12830 (N_12830,N_11237,N_11890);
or U12831 (N_12831,N_11042,N_11706);
nor U12832 (N_12832,N_11635,N_11019);
and U12833 (N_12833,N_11625,N_11931);
xor U12834 (N_12834,N_11148,N_11654);
nand U12835 (N_12835,N_11805,N_11029);
nor U12836 (N_12836,N_11287,N_11718);
nand U12837 (N_12837,N_11013,N_11275);
and U12838 (N_12838,N_11775,N_11204);
nand U12839 (N_12839,N_11650,N_11053);
nand U12840 (N_12840,N_11209,N_11009);
nand U12841 (N_12841,N_11968,N_11012);
nand U12842 (N_12842,N_11651,N_11647);
xor U12843 (N_12843,N_11400,N_11139);
or U12844 (N_12844,N_11163,N_11081);
nor U12845 (N_12845,N_11432,N_11722);
or U12846 (N_12846,N_11322,N_11892);
nor U12847 (N_12847,N_11216,N_11451);
nor U12848 (N_12848,N_11801,N_11475);
nor U12849 (N_12849,N_11176,N_11533);
or U12850 (N_12850,N_11472,N_11227);
or U12851 (N_12851,N_11717,N_11045);
nor U12852 (N_12852,N_11676,N_11183);
nand U12853 (N_12853,N_11478,N_11289);
xnor U12854 (N_12854,N_11077,N_11480);
nand U12855 (N_12855,N_11927,N_11430);
xor U12856 (N_12856,N_11478,N_11783);
and U12857 (N_12857,N_11128,N_11679);
nor U12858 (N_12858,N_11553,N_11227);
or U12859 (N_12859,N_11974,N_11431);
nand U12860 (N_12860,N_11575,N_11620);
xnor U12861 (N_12861,N_11324,N_11606);
and U12862 (N_12862,N_11484,N_11609);
xnor U12863 (N_12863,N_11324,N_11602);
xnor U12864 (N_12864,N_11798,N_11411);
or U12865 (N_12865,N_11562,N_11325);
and U12866 (N_12866,N_11760,N_11698);
and U12867 (N_12867,N_11877,N_11573);
nor U12868 (N_12868,N_11863,N_11140);
xor U12869 (N_12869,N_11752,N_11882);
and U12870 (N_12870,N_11067,N_11897);
nand U12871 (N_12871,N_11707,N_11573);
nand U12872 (N_12872,N_11841,N_11956);
xor U12873 (N_12873,N_11264,N_11220);
or U12874 (N_12874,N_11398,N_11953);
xnor U12875 (N_12875,N_11743,N_11460);
and U12876 (N_12876,N_11069,N_11814);
and U12877 (N_12877,N_11240,N_11285);
and U12878 (N_12878,N_11003,N_11188);
nor U12879 (N_12879,N_11742,N_11069);
and U12880 (N_12880,N_11472,N_11633);
nand U12881 (N_12881,N_11332,N_11234);
xor U12882 (N_12882,N_11779,N_11640);
nor U12883 (N_12883,N_11812,N_11031);
and U12884 (N_12884,N_11338,N_11871);
or U12885 (N_12885,N_11237,N_11581);
nor U12886 (N_12886,N_11029,N_11672);
and U12887 (N_12887,N_11732,N_11662);
and U12888 (N_12888,N_11310,N_11639);
or U12889 (N_12889,N_11778,N_11044);
or U12890 (N_12890,N_11133,N_11417);
nor U12891 (N_12891,N_11408,N_11458);
nor U12892 (N_12892,N_11972,N_11227);
and U12893 (N_12893,N_11612,N_11932);
xnor U12894 (N_12894,N_11106,N_11822);
and U12895 (N_12895,N_11630,N_11662);
xor U12896 (N_12896,N_11375,N_11797);
or U12897 (N_12897,N_11109,N_11523);
and U12898 (N_12898,N_11297,N_11204);
nand U12899 (N_12899,N_11366,N_11511);
or U12900 (N_12900,N_11258,N_11496);
nor U12901 (N_12901,N_11561,N_11369);
or U12902 (N_12902,N_11679,N_11550);
xor U12903 (N_12903,N_11469,N_11003);
and U12904 (N_12904,N_11868,N_11850);
nand U12905 (N_12905,N_11246,N_11552);
nand U12906 (N_12906,N_11866,N_11530);
and U12907 (N_12907,N_11485,N_11368);
xnor U12908 (N_12908,N_11532,N_11262);
and U12909 (N_12909,N_11943,N_11202);
and U12910 (N_12910,N_11225,N_11723);
or U12911 (N_12911,N_11816,N_11933);
nand U12912 (N_12912,N_11470,N_11129);
and U12913 (N_12913,N_11615,N_11591);
or U12914 (N_12914,N_11032,N_11403);
xnor U12915 (N_12915,N_11201,N_11660);
nand U12916 (N_12916,N_11449,N_11812);
or U12917 (N_12917,N_11873,N_11329);
xor U12918 (N_12918,N_11823,N_11513);
nand U12919 (N_12919,N_11690,N_11123);
nand U12920 (N_12920,N_11747,N_11818);
or U12921 (N_12921,N_11691,N_11001);
or U12922 (N_12922,N_11926,N_11953);
nor U12923 (N_12923,N_11279,N_11580);
nor U12924 (N_12924,N_11882,N_11807);
and U12925 (N_12925,N_11016,N_11834);
and U12926 (N_12926,N_11357,N_11771);
nor U12927 (N_12927,N_11604,N_11446);
nor U12928 (N_12928,N_11675,N_11828);
nand U12929 (N_12929,N_11117,N_11719);
xor U12930 (N_12930,N_11817,N_11229);
nor U12931 (N_12931,N_11943,N_11718);
and U12932 (N_12932,N_11113,N_11001);
and U12933 (N_12933,N_11120,N_11379);
nor U12934 (N_12934,N_11983,N_11948);
or U12935 (N_12935,N_11555,N_11019);
and U12936 (N_12936,N_11558,N_11650);
or U12937 (N_12937,N_11429,N_11275);
nor U12938 (N_12938,N_11339,N_11066);
or U12939 (N_12939,N_11009,N_11150);
nor U12940 (N_12940,N_11045,N_11938);
or U12941 (N_12941,N_11454,N_11096);
or U12942 (N_12942,N_11309,N_11052);
nand U12943 (N_12943,N_11110,N_11016);
and U12944 (N_12944,N_11227,N_11168);
nor U12945 (N_12945,N_11591,N_11286);
or U12946 (N_12946,N_11913,N_11900);
and U12947 (N_12947,N_11727,N_11455);
or U12948 (N_12948,N_11513,N_11387);
nand U12949 (N_12949,N_11395,N_11622);
nand U12950 (N_12950,N_11150,N_11867);
nor U12951 (N_12951,N_11076,N_11116);
xnor U12952 (N_12952,N_11012,N_11700);
and U12953 (N_12953,N_11981,N_11254);
nand U12954 (N_12954,N_11416,N_11412);
xor U12955 (N_12955,N_11240,N_11932);
xnor U12956 (N_12956,N_11246,N_11261);
nor U12957 (N_12957,N_11891,N_11359);
and U12958 (N_12958,N_11737,N_11772);
or U12959 (N_12959,N_11043,N_11765);
xnor U12960 (N_12960,N_11602,N_11441);
xnor U12961 (N_12961,N_11775,N_11720);
nand U12962 (N_12962,N_11340,N_11246);
nor U12963 (N_12963,N_11805,N_11967);
nand U12964 (N_12964,N_11865,N_11837);
or U12965 (N_12965,N_11270,N_11707);
nor U12966 (N_12966,N_11317,N_11357);
xnor U12967 (N_12967,N_11422,N_11064);
or U12968 (N_12968,N_11142,N_11291);
and U12969 (N_12969,N_11046,N_11088);
and U12970 (N_12970,N_11102,N_11649);
xnor U12971 (N_12971,N_11517,N_11884);
and U12972 (N_12972,N_11355,N_11413);
xnor U12973 (N_12973,N_11019,N_11941);
or U12974 (N_12974,N_11120,N_11808);
or U12975 (N_12975,N_11300,N_11499);
nor U12976 (N_12976,N_11799,N_11313);
and U12977 (N_12977,N_11233,N_11824);
xor U12978 (N_12978,N_11910,N_11957);
nand U12979 (N_12979,N_11837,N_11642);
and U12980 (N_12980,N_11055,N_11302);
nor U12981 (N_12981,N_11237,N_11537);
or U12982 (N_12982,N_11419,N_11761);
xor U12983 (N_12983,N_11438,N_11983);
xor U12984 (N_12984,N_11429,N_11139);
xor U12985 (N_12985,N_11726,N_11404);
nand U12986 (N_12986,N_11503,N_11872);
nor U12987 (N_12987,N_11819,N_11371);
and U12988 (N_12988,N_11764,N_11861);
nand U12989 (N_12989,N_11493,N_11576);
and U12990 (N_12990,N_11136,N_11201);
or U12991 (N_12991,N_11143,N_11214);
or U12992 (N_12992,N_11123,N_11533);
or U12993 (N_12993,N_11269,N_11080);
or U12994 (N_12994,N_11495,N_11642);
nor U12995 (N_12995,N_11421,N_11376);
xnor U12996 (N_12996,N_11910,N_11936);
xnor U12997 (N_12997,N_11388,N_11390);
xnor U12998 (N_12998,N_11400,N_11351);
xnor U12999 (N_12999,N_11836,N_11926);
nor U13000 (N_13000,N_12443,N_12869);
and U13001 (N_13001,N_12233,N_12172);
xor U13002 (N_13002,N_12738,N_12886);
nand U13003 (N_13003,N_12573,N_12097);
and U13004 (N_13004,N_12594,N_12433);
and U13005 (N_13005,N_12446,N_12916);
or U13006 (N_13006,N_12863,N_12460);
nor U13007 (N_13007,N_12153,N_12262);
xnor U13008 (N_13008,N_12119,N_12611);
or U13009 (N_13009,N_12899,N_12568);
and U13010 (N_13010,N_12223,N_12282);
nand U13011 (N_13011,N_12324,N_12205);
or U13012 (N_13012,N_12931,N_12803);
nor U13013 (N_13013,N_12691,N_12947);
and U13014 (N_13014,N_12855,N_12212);
or U13015 (N_13015,N_12378,N_12111);
nor U13016 (N_13016,N_12686,N_12471);
xor U13017 (N_13017,N_12071,N_12929);
nand U13018 (N_13018,N_12708,N_12839);
nand U13019 (N_13019,N_12046,N_12984);
and U13020 (N_13020,N_12250,N_12320);
xnor U13021 (N_13021,N_12346,N_12570);
xnor U13022 (N_13022,N_12149,N_12240);
nor U13023 (N_13023,N_12315,N_12844);
xnor U13024 (N_13024,N_12652,N_12575);
and U13025 (N_13025,N_12644,N_12053);
or U13026 (N_13026,N_12184,N_12749);
and U13027 (N_13027,N_12058,N_12163);
nor U13028 (N_13028,N_12330,N_12779);
nand U13029 (N_13029,N_12655,N_12638);
xnor U13030 (N_13030,N_12525,N_12624);
or U13031 (N_13031,N_12906,N_12273);
nand U13032 (N_13032,N_12334,N_12550);
nand U13033 (N_13033,N_12439,N_12634);
and U13034 (N_13034,N_12455,N_12487);
nor U13035 (N_13035,N_12410,N_12619);
nor U13036 (N_13036,N_12123,N_12880);
nand U13037 (N_13037,N_12989,N_12909);
and U13038 (N_13038,N_12354,N_12201);
nand U13039 (N_13039,N_12635,N_12539);
or U13040 (N_13040,N_12725,N_12962);
nand U13041 (N_13041,N_12679,N_12741);
xor U13042 (N_13042,N_12774,N_12535);
or U13043 (N_13043,N_12778,N_12585);
xnor U13044 (N_13044,N_12672,N_12292);
xor U13045 (N_13045,N_12753,N_12599);
xnor U13046 (N_13046,N_12811,N_12829);
or U13047 (N_13047,N_12561,N_12579);
or U13048 (N_13048,N_12077,N_12249);
nor U13049 (N_13049,N_12166,N_12875);
and U13050 (N_13050,N_12593,N_12505);
nor U13051 (N_13051,N_12372,N_12332);
xnor U13052 (N_13052,N_12073,N_12082);
xor U13053 (N_13053,N_12995,N_12059);
xnor U13054 (N_13054,N_12609,N_12588);
nor U13055 (N_13055,N_12202,N_12854);
nand U13056 (N_13056,N_12701,N_12414);
or U13057 (N_13057,N_12050,N_12998);
nand U13058 (N_13058,N_12402,N_12775);
nand U13059 (N_13059,N_12030,N_12274);
nand U13060 (N_13060,N_12789,N_12727);
and U13061 (N_13061,N_12801,N_12280);
or U13062 (N_13062,N_12057,N_12940);
nand U13063 (N_13063,N_12807,N_12232);
xnor U13064 (N_13064,N_12013,N_12662);
nor U13065 (N_13065,N_12895,N_12698);
and U13066 (N_13066,N_12120,N_12098);
nand U13067 (N_13067,N_12628,N_12583);
xor U13068 (N_13068,N_12196,N_12467);
or U13069 (N_13069,N_12648,N_12362);
xnor U13070 (N_13070,N_12721,N_12355);
nand U13071 (N_13071,N_12840,N_12667);
nand U13072 (N_13072,N_12608,N_12828);
or U13073 (N_13073,N_12926,N_12382);
and U13074 (N_13074,N_12215,N_12183);
xnor U13075 (N_13075,N_12289,N_12833);
and U13076 (N_13076,N_12952,N_12331);
nor U13077 (N_13077,N_12818,N_12411);
nand U13078 (N_13078,N_12534,N_12470);
and U13079 (N_13079,N_12421,N_12804);
or U13080 (N_13080,N_12258,N_12546);
and U13081 (N_13081,N_12156,N_12649);
or U13082 (N_13082,N_12650,N_12036);
or U13083 (N_13083,N_12752,N_12415);
and U13084 (N_13084,N_12269,N_12155);
and U13085 (N_13085,N_12620,N_12285);
or U13086 (N_13086,N_12566,N_12560);
nand U13087 (N_13087,N_12519,N_12238);
nor U13088 (N_13088,N_12496,N_12316);
and U13089 (N_13089,N_12671,N_12515);
or U13090 (N_13090,N_12279,N_12365);
and U13091 (N_13091,N_12857,N_12220);
nand U13092 (N_13092,N_12657,N_12264);
or U13093 (N_13093,N_12625,N_12217);
nor U13094 (N_13094,N_12230,N_12049);
or U13095 (N_13095,N_12255,N_12006);
or U13096 (N_13096,N_12819,N_12179);
and U13097 (N_13097,N_12602,N_12261);
nand U13098 (N_13098,N_12040,N_12437);
or U13099 (N_13099,N_12958,N_12208);
xnor U13100 (N_13100,N_12994,N_12802);
nor U13101 (N_13101,N_12557,N_12533);
and U13102 (N_13102,N_12696,N_12390);
nor U13103 (N_13103,N_12787,N_12419);
nand U13104 (N_13104,N_12214,N_12921);
nand U13105 (N_13105,N_12490,N_12225);
or U13106 (N_13106,N_12095,N_12963);
nand U13107 (N_13107,N_12675,N_12764);
nand U13108 (N_13108,N_12707,N_12981);
and U13109 (N_13109,N_12061,N_12878);
or U13110 (N_13110,N_12480,N_12834);
nand U13111 (N_13111,N_12506,N_12595);
nor U13112 (N_13112,N_12888,N_12861);
nor U13113 (N_13113,N_12047,N_12937);
and U13114 (N_13114,N_12345,N_12511);
or U13115 (N_13115,N_12706,N_12141);
nor U13116 (N_13116,N_12942,N_12128);
or U13117 (N_13117,N_12536,N_12814);
and U13118 (N_13118,N_12216,N_12526);
xnor U13119 (N_13119,N_12389,N_12021);
nand U13120 (N_13120,N_12008,N_12224);
or U13121 (N_13121,N_12112,N_12150);
nor U13122 (N_13122,N_12710,N_12288);
nand U13123 (N_13123,N_12969,N_12837);
and U13124 (N_13124,N_12482,N_12483);
nor U13125 (N_13125,N_12584,N_12661);
nor U13126 (N_13126,N_12842,N_12676);
nor U13127 (N_13127,N_12422,N_12134);
xnor U13128 (N_13128,N_12266,N_12883);
and U13129 (N_13129,N_12604,N_12800);
nor U13130 (N_13130,N_12398,N_12824);
and U13131 (N_13131,N_12291,N_12178);
nand U13132 (N_13132,N_12328,N_12659);
and U13133 (N_13133,N_12125,N_12256);
nand U13134 (N_13134,N_12094,N_12849);
xor U13135 (N_13135,N_12502,N_12528);
or U13136 (N_13136,N_12297,N_12394);
or U13137 (N_13137,N_12581,N_12722);
xnor U13138 (N_13138,N_12531,N_12106);
xor U13139 (N_13139,N_12514,N_12379);
nor U13140 (N_13140,N_12322,N_12333);
and U13141 (N_13141,N_12976,N_12758);
xor U13142 (N_13142,N_12780,N_12086);
or U13143 (N_13143,N_12554,N_12312);
nand U13144 (N_13144,N_12750,N_12089);
nand U13145 (N_13145,N_12180,N_12041);
nand U13146 (N_13146,N_12173,N_12518);
or U13147 (N_13147,N_12397,N_12812);
nand U13148 (N_13148,N_12306,N_12713);
or U13149 (N_13149,N_12973,N_12001);
and U13150 (N_13150,N_12567,N_12191);
xnor U13151 (N_13151,N_12275,N_12896);
xnor U13152 (N_13152,N_12504,N_12508);
nand U13153 (N_13153,N_12831,N_12339);
and U13154 (N_13154,N_12427,N_12733);
nor U13155 (N_13155,N_12712,N_12856);
nor U13156 (N_13156,N_12610,N_12772);
xor U13157 (N_13157,N_12847,N_12965);
or U13158 (N_13158,N_12574,N_12352);
nand U13159 (N_13159,N_12907,N_12616);
and U13160 (N_13160,N_12336,N_12598);
xnor U13161 (N_13161,N_12431,N_12497);
and U13162 (N_13162,N_12674,N_12080);
or U13163 (N_13163,N_12243,N_12793);
xnor U13164 (N_13164,N_12950,N_12293);
nand U13165 (N_13165,N_12582,N_12190);
and U13166 (N_13166,N_12517,N_12085);
xor U13167 (N_13167,N_12865,N_12299);
xor U13168 (N_13168,N_12129,N_12537);
nor U13169 (N_13169,N_12023,N_12777);
and U13170 (N_13170,N_12359,N_12991);
or U13171 (N_13171,N_12392,N_12783);
nor U13172 (N_13172,N_12016,N_12720);
nor U13173 (N_13173,N_12034,N_12067);
or U13174 (N_13174,N_12795,N_12375);
xnor U13175 (N_13175,N_12118,N_12409);
and U13176 (N_13176,N_12136,N_12520);
or U13177 (N_13177,N_12360,N_12386);
and U13178 (N_13178,N_12350,N_12673);
or U13179 (N_13179,N_12003,N_12709);
and U13180 (N_13180,N_12719,N_12088);
nand U13181 (N_13181,N_12270,N_12908);
xor U13182 (N_13182,N_12724,N_12396);
nor U13183 (N_13183,N_12157,N_12992);
or U13184 (N_13184,N_12479,N_12423);
and U13185 (N_13185,N_12209,N_12596);
nand U13186 (N_13186,N_12254,N_12944);
nand U13187 (N_13187,N_12914,N_12318);
nand U13188 (N_13188,N_12187,N_12476);
and U13189 (N_13189,N_12668,N_12426);
nor U13190 (N_13190,N_12559,N_12226);
nand U13191 (N_13191,N_12821,N_12605);
nor U13192 (N_13192,N_12744,N_12391);
xnor U13193 (N_13193,N_12660,N_12083);
and U13194 (N_13194,N_12435,N_12064);
nor U13195 (N_13195,N_12501,N_12472);
or U13196 (N_13196,N_12323,N_12406);
nor U13197 (N_13197,N_12503,N_12101);
xor U13198 (N_13198,N_12843,N_12445);
xor U13199 (N_13199,N_12314,N_12177);
xnor U13200 (N_13200,N_12798,N_12056);
and U13201 (N_13201,N_12924,N_12489);
nor U13202 (N_13202,N_12257,N_12882);
xnor U13203 (N_13203,N_12934,N_12160);
xor U13204 (N_13204,N_12158,N_12116);
nor U13205 (N_13205,N_12678,N_12465);
xnor U13206 (N_13206,N_12769,N_12010);
nand U13207 (N_13207,N_12690,N_12137);
and U13208 (N_13208,N_12731,N_12076);
and U13209 (N_13209,N_12577,N_12632);
or U13210 (N_13210,N_12495,N_12627);
nand U13211 (N_13211,N_12797,N_12523);
xor U13212 (N_13212,N_12565,N_12167);
xnor U13213 (N_13213,N_12151,N_12728);
nor U13214 (N_13214,N_12052,N_12681);
nand U13215 (N_13215,N_12213,N_12613);
xnor U13216 (N_13216,N_12004,N_12239);
nand U13217 (N_13217,N_12009,N_12222);
nor U13218 (N_13218,N_12296,N_12308);
nor U13219 (N_13219,N_12968,N_12425);
nand U13220 (N_13220,N_12327,N_12986);
nor U13221 (N_13221,N_12453,N_12735);
xnor U13222 (N_13222,N_12541,N_12927);
nor U13223 (N_13223,N_12913,N_12461);
xor U13224 (N_13224,N_12571,N_12260);
nor U13225 (N_13225,N_12353,N_12867);
and U13226 (N_13226,N_12715,N_12317);
or U13227 (N_13227,N_12766,N_12960);
and U13228 (N_13228,N_12990,N_12408);
nand U13229 (N_13229,N_12377,N_12956);
or U13230 (N_13230,N_12663,N_12538);
and U13231 (N_13231,N_12848,N_12692);
and U13232 (N_13232,N_12716,N_12945);
xor U13233 (N_13233,N_12093,N_12303);
xor U13234 (N_13234,N_12351,N_12259);
and U13235 (N_13235,N_12890,N_12458);
nand U13236 (N_13236,N_12033,N_12817);
or U13237 (N_13237,N_12621,N_12265);
nor U13238 (N_13238,N_12176,N_12108);
nor U13239 (N_13239,N_12245,N_12302);
xnor U13240 (N_13240,N_12794,N_12979);
nor U13241 (N_13241,N_12953,N_12161);
nor U13242 (N_13242,N_12169,N_12898);
or U13243 (N_13243,N_12450,N_12197);
xor U13244 (N_13244,N_12236,N_12174);
nor U13245 (N_13245,N_12054,N_12615);
nand U13246 (N_13246,N_12796,N_12131);
nor U13247 (N_13247,N_12547,N_12060);
or U13248 (N_13248,N_12640,N_12670);
or U13249 (N_13249,N_12893,N_12987);
or U13250 (N_13250,N_12955,N_12109);
or U13251 (N_13251,N_12494,N_12486);
or U13252 (N_13252,N_12019,N_12743);
nor U13253 (N_13253,N_12488,N_12031);
and U13254 (N_13254,N_12403,N_12910);
or U13255 (N_13255,N_12922,N_12832);
and U13256 (N_13256,N_12186,N_12204);
nor U13257 (N_13257,N_12048,N_12911);
or U13258 (N_13258,N_12734,N_12768);
nor U13259 (N_13259,N_12072,N_12607);
xor U13260 (N_13260,N_12231,N_12932);
nand U13261 (N_13261,N_12773,N_12879);
or U13262 (N_13262,N_12203,N_12871);
xor U13263 (N_13263,N_12551,N_12841);
or U13264 (N_13264,N_12124,N_12020);
and U13265 (N_13265,N_12835,N_12498);
nor U13266 (N_13266,N_12874,N_12127);
and U13267 (N_13267,N_12281,N_12558);
nand U13268 (N_13268,N_12105,N_12977);
and U13269 (N_13269,N_12027,N_12918);
nor U13270 (N_13270,N_12466,N_12144);
xor U13271 (N_13271,N_12162,N_12925);
or U13272 (N_13272,N_12740,N_12873);
nor U13273 (N_13273,N_12272,N_12263);
xor U13274 (N_13274,N_12694,N_12170);
and U13275 (N_13275,N_12530,N_12711);
nor U13276 (N_13276,N_12387,N_12074);
nand U13277 (N_13277,N_12007,N_12478);
and U13278 (N_13278,N_12597,N_12756);
xnor U13279 (N_13279,N_12442,N_12147);
and U13280 (N_13280,N_12348,N_12666);
or U13281 (N_13281,N_12693,N_12456);
xor U13282 (N_13282,N_12894,N_12714);
or U13283 (N_13283,N_12363,N_12358);
xor U13284 (N_13284,N_12846,N_12737);
nand U13285 (N_13285,N_12117,N_12527);
or U13286 (N_13286,N_12943,N_12126);
or U13287 (N_13287,N_12189,N_12276);
nand U13288 (N_13288,N_12685,N_12286);
or U13289 (N_13289,N_12904,N_12669);
nor U13290 (N_13290,N_12747,N_12081);
xnor U13291 (N_13291,N_12905,N_12540);
or U13292 (N_13292,N_12370,N_12891);
xor U13293 (N_13293,N_12481,N_12298);
or U13294 (N_13294,N_12100,N_12055);
nor U13295 (N_13295,N_12246,N_12374);
nor U13296 (N_13296,N_12110,N_12405);
nand U13297 (N_13297,N_12569,N_12484);
or U13298 (N_13298,N_12881,N_12107);
or U13299 (N_13299,N_12785,N_12967);
nand U13300 (N_13300,N_12211,N_12463);
nor U13301 (N_13301,N_12809,N_12664);
or U13302 (N_13302,N_12210,N_12996);
nor U13303 (N_13303,N_12510,N_12552);
or U13304 (N_13304,N_12251,N_12622);
and U13305 (N_13305,N_12234,N_12920);
nand U13306 (N_13306,N_12959,N_12626);
or U13307 (N_13307,N_12658,N_12133);
or U13308 (N_13308,N_12782,N_12578);
nand U13309 (N_13309,N_12207,N_12325);
xor U13310 (N_13310,N_12014,N_12175);
nand U13311 (N_13311,N_12140,N_12200);
and U13312 (N_13312,N_12786,N_12139);
nor U13313 (N_13313,N_12680,N_12278);
xor U13314 (N_13314,N_12545,N_12424);
nor U13315 (N_13315,N_12970,N_12826);
nand U13316 (N_13316,N_12459,N_12342);
nand U13317 (N_13317,N_12677,N_12454);
nand U13318 (N_13318,N_12618,N_12182);
xor U13319 (N_13319,N_12654,N_12978);
nand U13320 (N_13320,N_12114,N_12765);
xor U13321 (N_13321,N_12294,N_12037);
or U13322 (N_13322,N_12930,N_12132);
or U13323 (N_13323,N_12941,N_12688);
or U13324 (N_13324,N_12042,N_12165);
nand U13325 (N_13325,N_12065,N_12235);
xnor U13326 (N_13326,N_12113,N_12935);
or U13327 (N_13327,N_12684,N_12002);
nand U13328 (N_13328,N_12748,N_12326);
nor U13329 (N_13329,N_12623,N_12647);
xor U13330 (N_13330,N_12589,N_12521);
and U13331 (N_13331,N_12268,N_12993);
nand U13332 (N_13332,N_12115,N_12705);
xor U13333 (N_13333,N_12473,N_12889);
or U13334 (N_13334,N_12901,N_12404);
nor U13335 (N_13335,N_12369,N_12591);
xnor U13336 (N_13336,N_12553,N_12951);
nor U13337 (N_13337,N_12335,N_12492);
xnor U13338 (N_13338,N_12143,N_12781);
and U13339 (N_13339,N_12972,N_12474);
nor U13340 (N_13340,N_12078,N_12860);
nor U13341 (N_13341,N_12877,N_12399);
nand U13342 (N_13342,N_12689,N_12079);
nor U13343 (N_13343,N_12122,N_12395);
or U13344 (N_13344,N_12154,N_12024);
or U13345 (N_13345,N_12321,N_12227);
and U13346 (N_13346,N_12838,N_12413);
and U13347 (N_13347,N_12954,N_12026);
xnor U13348 (N_13348,N_12902,N_12305);
nor U13349 (N_13349,N_12641,N_12063);
nor U13350 (N_13350,N_12767,N_12859);
and U13351 (N_13351,N_12416,N_12499);
xor U13352 (N_13352,N_12313,N_12146);
xnor U13353 (N_13353,N_12636,N_12702);
and U13354 (N_13354,N_12475,N_12185);
or U13355 (N_13355,N_12820,N_12357);
nand U13356 (N_13356,N_12919,N_12915);
nor U13357 (N_13357,N_12237,N_12851);
nor U13358 (N_13358,N_12181,N_12917);
nor U13359 (N_13359,N_12300,N_12606);
and U13360 (N_13360,N_12700,N_12412);
nand U13361 (N_13361,N_12938,N_12436);
and U13362 (N_13362,N_12500,N_12897);
or U13363 (N_13363,N_12928,N_12364);
nor U13364 (N_13364,N_12017,N_12988);
or U13365 (N_13365,N_12633,N_12509);
xnor U13366 (N_13366,N_12444,N_12563);
xor U13367 (N_13367,N_12068,N_12104);
and U13368 (N_13368,N_12903,N_12337);
and U13369 (N_13369,N_12029,N_12892);
xnor U13370 (N_13370,N_12142,N_12248);
nor U13371 (N_13371,N_12310,N_12939);
xor U13372 (N_13372,N_12761,N_12228);
or U13373 (N_13373,N_12617,N_12949);
or U13374 (N_13374,N_12152,N_12736);
nor U13375 (N_13375,N_12946,N_12576);
xnor U13376 (N_13376,N_12066,N_12742);
or U13377 (N_13377,N_12440,N_12221);
and U13378 (N_13378,N_12420,N_12580);
xor U13379 (N_13379,N_12816,N_12542);
or U13380 (N_13380,N_12092,N_12380);
and U13381 (N_13381,N_12643,N_12825);
xor U13382 (N_13382,N_12381,N_12776);
xor U13383 (N_13383,N_12192,N_12367);
and U13384 (N_13384,N_12687,N_12069);
and U13385 (N_13385,N_12980,N_12513);
or U13386 (N_13386,N_12754,N_12287);
xnor U13387 (N_13387,N_12507,N_12823);
and U13388 (N_13388,N_12600,N_12799);
and U13389 (N_13389,N_12544,N_12341);
nand U13390 (N_13390,N_12301,N_12319);
nand U13391 (N_13391,N_12198,N_12028);
or U13392 (N_13392,N_12683,N_12726);
nand U13393 (N_13393,N_12253,N_12193);
nand U13394 (N_13394,N_12639,N_12241);
or U13395 (N_13395,N_12271,N_12864);
xor U13396 (N_13396,N_12850,N_12784);
nand U13397 (N_13397,N_12805,N_12732);
or U13398 (N_13398,N_12462,N_12592);
or U13399 (N_13399,N_12770,N_12751);
or U13400 (N_13400,N_12304,N_12642);
nor U13401 (N_13401,N_12145,N_12051);
or U13402 (N_13402,N_12656,N_12813);
nor U13403 (N_13403,N_12830,N_12457);
xor U13404 (N_13404,N_12148,N_12791);
and U13405 (N_13405,N_12384,N_12090);
nor U13406 (N_13406,N_12651,N_12697);
and U13407 (N_13407,N_12356,N_12448);
or U13408 (N_13408,N_12637,N_12091);
nand U13409 (N_13409,N_12997,N_12385);
and U13410 (N_13410,N_12344,N_12792);
nor U13411 (N_13411,N_12159,N_12745);
and U13412 (N_13412,N_12070,N_12022);
and U13413 (N_13413,N_12038,N_12366);
nand U13414 (N_13414,N_12788,N_12469);
xor U13415 (N_13415,N_12603,N_12295);
nand U13416 (N_13416,N_12532,N_12340);
or U13417 (N_13417,N_12999,N_12522);
or U13418 (N_13418,N_12555,N_12005);
or U13419 (N_13419,N_12062,N_12884);
and U13420 (N_13420,N_12827,N_12746);
xor U13421 (N_13421,N_12477,N_12099);
nor U13422 (N_13422,N_12376,N_12371);
nand U13423 (N_13423,N_12631,N_12218);
xor U13424 (N_13424,N_12524,N_12548);
nor U13425 (N_13425,N_12485,N_12964);
nand U13426 (N_13426,N_12373,N_12933);
nor U13427 (N_13427,N_12000,N_12252);
and U13428 (N_13428,N_12887,N_12957);
xor U13429 (N_13429,N_12866,N_12590);
or U13430 (N_13430,N_12572,N_12307);
nand U13431 (N_13431,N_12138,N_12730);
xnor U13432 (N_13432,N_12368,N_12277);
nor U13433 (N_13433,N_12464,N_12361);
xor U13434 (N_13434,N_12451,N_12452);
or U13435 (N_13435,N_12032,N_12836);
nand U13436 (N_13436,N_12432,N_12206);
nor U13437 (N_13437,N_12418,N_12815);
xnor U13438 (N_13438,N_12103,N_12188);
nand U13439 (N_13439,N_12195,N_12974);
nor U13440 (N_13440,N_12018,N_12309);
or U13441 (N_13441,N_12630,N_12739);
or U13442 (N_13442,N_12948,N_12587);
nor U13443 (N_13443,N_12199,N_12755);
or U13444 (N_13444,N_12283,N_12075);
nor U13445 (N_13445,N_12512,N_12025);
xor U13446 (N_13446,N_12493,N_12383);
nand U13447 (N_13447,N_12703,N_12876);
and U13448 (N_13448,N_12975,N_12808);
or U13449 (N_13449,N_12044,N_12760);
xor U13450 (N_13450,N_12982,N_12718);
and U13451 (N_13451,N_12194,N_12084);
or U13452 (N_13452,N_12845,N_12564);
and U13453 (N_13453,N_12966,N_12247);
nor U13454 (N_13454,N_12983,N_12900);
or U13455 (N_13455,N_12400,N_12810);
nor U13456 (N_13456,N_12438,N_12759);
nand U13457 (N_13457,N_12311,N_12338);
or U13458 (N_13458,N_12468,N_12612);
xnor U13459 (N_13459,N_12015,N_12549);
and U13460 (N_13460,N_12586,N_12923);
nand U13461 (N_13461,N_12035,N_12853);
or U13462 (N_13462,N_12601,N_12762);
nand U13463 (N_13463,N_12529,N_12646);
or U13464 (N_13464,N_12087,N_12102);
xor U13465 (N_13465,N_12429,N_12858);
or U13466 (N_13466,N_12562,N_12343);
nor U13467 (N_13467,N_12244,N_12790);
or U13468 (N_13468,N_12267,N_12012);
nand U13469 (N_13469,N_12695,N_12862);
xor U13470 (N_13470,N_12614,N_12516);
and U13471 (N_13471,N_12822,N_12870);
nand U13472 (N_13472,N_12757,N_12699);
nor U13473 (N_13473,N_12096,N_12043);
xnor U13474 (N_13474,N_12682,N_12936);
or U13475 (N_13475,N_12430,N_12852);
nand U13476 (N_13476,N_12729,N_12388);
or U13477 (N_13477,N_12242,N_12704);
nor U13478 (N_13478,N_12543,N_12771);
nand U13479 (N_13479,N_12961,N_12045);
or U13480 (N_13480,N_12349,N_12971);
nor U13481 (N_13481,N_12229,N_12164);
and U13482 (N_13482,N_12449,N_12401);
and U13483 (N_13483,N_12135,N_12491);
and U13484 (N_13484,N_12219,N_12665);
nand U13485 (N_13485,N_12653,N_12407);
and U13486 (N_13486,N_12393,N_12447);
or U13487 (N_13487,N_12428,N_12130);
nor U13488 (N_13488,N_12329,N_12039);
or U13489 (N_13489,N_12121,N_12168);
nand U13490 (N_13490,N_12556,N_12011);
and U13491 (N_13491,N_12629,N_12763);
nand U13492 (N_13492,N_12806,N_12434);
xnor U13493 (N_13493,N_12171,N_12717);
nor U13494 (N_13494,N_12868,N_12347);
nand U13495 (N_13495,N_12985,N_12885);
xor U13496 (N_13496,N_12645,N_12417);
nand U13497 (N_13497,N_12290,N_12284);
or U13498 (N_13498,N_12441,N_12912);
nor U13499 (N_13499,N_12723,N_12872);
or U13500 (N_13500,N_12215,N_12612);
xor U13501 (N_13501,N_12873,N_12227);
nand U13502 (N_13502,N_12810,N_12021);
nand U13503 (N_13503,N_12137,N_12106);
nand U13504 (N_13504,N_12887,N_12330);
nor U13505 (N_13505,N_12490,N_12890);
nor U13506 (N_13506,N_12279,N_12482);
nor U13507 (N_13507,N_12350,N_12730);
nor U13508 (N_13508,N_12223,N_12154);
nor U13509 (N_13509,N_12078,N_12070);
and U13510 (N_13510,N_12368,N_12560);
or U13511 (N_13511,N_12765,N_12674);
nand U13512 (N_13512,N_12130,N_12397);
nor U13513 (N_13513,N_12537,N_12197);
or U13514 (N_13514,N_12567,N_12398);
nand U13515 (N_13515,N_12635,N_12833);
xor U13516 (N_13516,N_12293,N_12221);
or U13517 (N_13517,N_12944,N_12522);
or U13518 (N_13518,N_12885,N_12524);
nor U13519 (N_13519,N_12087,N_12780);
or U13520 (N_13520,N_12612,N_12157);
nor U13521 (N_13521,N_12145,N_12974);
nand U13522 (N_13522,N_12505,N_12327);
nand U13523 (N_13523,N_12092,N_12402);
or U13524 (N_13524,N_12249,N_12813);
xnor U13525 (N_13525,N_12063,N_12804);
nor U13526 (N_13526,N_12352,N_12656);
nand U13527 (N_13527,N_12445,N_12134);
xor U13528 (N_13528,N_12335,N_12890);
nand U13529 (N_13529,N_12010,N_12514);
and U13530 (N_13530,N_12556,N_12706);
nand U13531 (N_13531,N_12397,N_12227);
nor U13532 (N_13532,N_12265,N_12558);
nand U13533 (N_13533,N_12139,N_12432);
nand U13534 (N_13534,N_12800,N_12506);
nand U13535 (N_13535,N_12630,N_12266);
and U13536 (N_13536,N_12271,N_12360);
and U13537 (N_13537,N_12787,N_12335);
and U13538 (N_13538,N_12276,N_12348);
nor U13539 (N_13539,N_12981,N_12535);
nand U13540 (N_13540,N_12555,N_12162);
nor U13541 (N_13541,N_12967,N_12924);
or U13542 (N_13542,N_12174,N_12534);
and U13543 (N_13543,N_12570,N_12246);
or U13544 (N_13544,N_12220,N_12717);
nor U13545 (N_13545,N_12390,N_12153);
and U13546 (N_13546,N_12779,N_12625);
nand U13547 (N_13547,N_12535,N_12337);
nor U13548 (N_13548,N_12806,N_12457);
nand U13549 (N_13549,N_12532,N_12079);
nor U13550 (N_13550,N_12571,N_12618);
xor U13551 (N_13551,N_12248,N_12442);
or U13552 (N_13552,N_12723,N_12188);
nand U13553 (N_13553,N_12989,N_12169);
nor U13554 (N_13554,N_12097,N_12067);
or U13555 (N_13555,N_12503,N_12937);
or U13556 (N_13556,N_12145,N_12687);
nand U13557 (N_13557,N_12909,N_12021);
nor U13558 (N_13558,N_12713,N_12937);
or U13559 (N_13559,N_12429,N_12819);
nand U13560 (N_13560,N_12117,N_12086);
nor U13561 (N_13561,N_12090,N_12757);
nand U13562 (N_13562,N_12274,N_12428);
xnor U13563 (N_13563,N_12024,N_12676);
xnor U13564 (N_13564,N_12779,N_12646);
nor U13565 (N_13565,N_12477,N_12285);
nor U13566 (N_13566,N_12563,N_12309);
nand U13567 (N_13567,N_12215,N_12143);
or U13568 (N_13568,N_12736,N_12327);
xnor U13569 (N_13569,N_12994,N_12602);
or U13570 (N_13570,N_12678,N_12191);
xor U13571 (N_13571,N_12441,N_12745);
nor U13572 (N_13572,N_12311,N_12099);
nor U13573 (N_13573,N_12935,N_12839);
nand U13574 (N_13574,N_12875,N_12691);
nand U13575 (N_13575,N_12996,N_12181);
nand U13576 (N_13576,N_12909,N_12523);
nor U13577 (N_13577,N_12539,N_12289);
or U13578 (N_13578,N_12586,N_12038);
and U13579 (N_13579,N_12621,N_12567);
xnor U13580 (N_13580,N_12496,N_12339);
and U13581 (N_13581,N_12019,N_12402);
or U13582 (N_13582,N_12675,N_12986);
nor U13583 (N_13583,N_12498,N_12136);
nand U13584 (N_13584,N_12454,N_12991);
or U13585 (N_13585,N_12619,N_12465);
xnor U13586 (N_13586,N_12110,N_12846);
xor U13587 (N_13587,N_12226,N_12724);
xor U13588 (N_13588,N_12885,N_12157);
nor U13589 (N_13589,N_12693,N_12859);
and U13590 (N_13590,N_12965,N_12321);
nand U13591 (N_13591,N_12748,N_12760);
xnor U13592 (N_13592,N_12011,N_12674);
and U13593 (N_13593,N_12616,N_12432);
xor U13594 (N_13594,N_12971,N_12907);
nor U13595 (N_13595,N_12729,N_12122);
and U13596 (N_13596,N_12424,N_12447);
xor U13597 (N_13597,N_12815,N_12782);
nand U13598 (N_13598,N_12484,N_12378);
xor U13599 (N_13599,N_12946,N_12496);
nor U13600 (N_13600,N_12359,N_12720);
nand U13601 (N_13601,N_12933,N_12685);
nand U13602 (N_13602,N_12575,N_12440);
xor U13603 (N_13603,N_12964,N_12729);
nor U13604 (N_13604,N_12407,N_12403);
xor U13605 (N_13605,N_12028,N_12575);
nand U13606 (N_13606,N_12595,N_12123);
nor U13607 (N_13607,N_12481,N_12812);
and U13608 (N_13608,N_12932,N_12865);
or U13609 (N_13609,N_12223,N_12928);
nand U13610 (N_13610,N_12474,N_12229);
nor U13611 (N_13611,N_12074,N_12658);
xor U13612 (N_13612,N_12476,N_12513);
or U13613 (N_13613,N_12759,N_12670);
nor U13614 (N_13614,N_12558,N_12234);
xor U13615 (N_13615,N_12522,N_12873);
xnor U13616 (N_13616,N_12302,N_12798);
nand U13617 (N_13617,N_12319,N_12831);
xnor U13618 (N_13618,N_12963,N_12274);
nand U13619 (N_13619,N_12880,N_12645);
nand U13620 (N_13620,N_12064,N_12005);
nor U13621 (N_13621,N_12727,N_12559);
or U13622 (N_13622,N_12092,N_12452);
or U13623 (N_13623,N_12062,N_12061);
or U13624 (N_13624,N_12833,N_12820);
xor U13625 (N_13625,N_12444,N_12274);
nor U13626 (N_13626,N_12520,N_12942);
and U13627 (N_13627,N_12280,N_12555);
xor U13628 (N_13628,N_12372,N_12436);
nand U13629 (N_13629,N_12529,N_12554);
or U13630 (N_13630,N_12226,N_12955);
nand U13631 (N_13631,N_12272,N_12283);
nand U13632 (N_13632,N_12296,N_12694);
xnor U13633 (N_13633,N_12467,N_12593);
and U13634 (N_13634,N_12763,N_12582);
and U13635 (N_13635,N_12356,N_12594);
and U13636 (N_13636,N_12610,N_12203);
xor U13637 (N_13637,N_12881,N_12261);
nor U13638 (N_13638,N_12274,N_12193);
nor U13639 (N_13639,N_12547,N_12043);
and U13640 (N_13640,N_12295,N_12723);
and U13641 (N_13641,N_12709,N_12442);
nor U13642 (N_13642,N_12972,N_12977);
or U13643 (N_13643,N_12763,N_12685);
xor U13644 (N_13644,N_12699,N_12559);
xor U13645 (N_13645,N_12207,N_12809);
nor U13646 (N_13646,N_12085,N_12531);
nor U13647 (N_13647,N_12786,N_12373);
xnor U13648 (N_13648,N_12597,N_12728);
nand U13649 (N_13649,N_12183,N_12719);
nor U13650 (N_13650,N_12649,N_12777);
nand U13651 (N_13651,N_12997,N_12894);
nand U13652 (N_13652,N_12975,N_12079);
nand U13653 (N_13653,N_12376,N_12933);
xnor U13654 (N_13654,N_12286,N_12833);
nand U13655 (N_13655,N_12077,N_12056);
nand U13656 (N_13656,N_12087,N_12285);
nand U13657 (N_13657,N_12748,N_12812);
xnor U13658 (N_13658,N_12971,N_12584);
nor U13659 (N_13659,N_12475,N_12983);
or U13660 (N_13660,N_12930,N_12414);
nor U13661 (N_13661,N_12736,N_12268);
xor U13662 (N_13662,N_12650,N_12695);
xnor U13663 (N_13663,N_12326,N_12891);
nand U13664 (N_13664,N_12950,N_12628);
xnor U13665 (N_13665,N_12530,N_12010);
xnor U13666 (N_13666,N_12169,N_12724);
or U13667 (N_13667,N_12708,N_12032);
or U13668 (N_13668,N_12021,N_12242);
or U13669 (N_13669,N_12712,N_12004);
nor U13670 (N_13670,N_12646,N_12063);
nand U13671 (N_13671,N_12502,N_12854);
xor U13672 (N_13672,N_12028,N_12345);
or U13673 (N_13673,N_12539,N_12954);
and U13674 (N_13674,N_12894,N_12301);
and U13675 (N_13675,N_12353,N_12953);
or U13676 (N_13676,N_12029,N_12632);
or U13677 (N_13677,N_12529,N_12108);
nand U13678 (N_13678,N_12097,N_12968);
or U13679 (N_13679,N_12469,N_12744);
nand U13680 (N_13680,N_12265,N_12308);
nand U13681 (N_13681,N_12479,N_12370);
or U13682 (N_13682,N_12768,N_12397);
and U13683 (N_13683,N_12474,N_12273);
and U13684 (N_13684,N_12946,N_12095);
or U13685 (N_13685,N_12658,N_12169);
or U13686 (N_13686,N_12309,N_12698);
nand U13687 (N_13687,N_12402,N_12910);
nor U13688 (N_13688,N_12875,N_12260);
or U13689 (N_13689,N_12627,N_12371);
and U13690 (N_13690,N_12691,N_12771);
xnor U13691 (N_13691,N_12046,N_12075);
nor U13692 (N_13692,N_12700,N_12049);
and U13693 (N_13693,N_12876,N_12651);
nand U13694 (N_13694,N_12983,N_12756);
and U13695 (N_13695,N_12229,N_12342);
and U13696 (N_13696,N_12089,N_12485);
and U13697 (N_13697,N_12688,N_12207);
and U13698 (N_13698,N_12464,N_12011);
or U13699 (N_13699,N_12609,N_12830);
nand U13700 (N_13700,N_12567,N_12060);
and U13701 (N_13701,N_12256,N_12009);
or U13702 (N_13702,N_12849,N_12997);
and U13703 (N_13703,N_12412,N_12418);
xor U13704 (N_13704,N_12906,N_12416);
nor U13705 (N_13705,N_12785,N_12612);
and U13706 (N_13706,N_12233,N_12236);
and U13707 (N_13707,N_12339,N_12429);
and U13708 (N_13708,N_12443,N_12185);
nand U13709 (N_13709,N_12407,N_12114);
or U13710 (N_13710,N_12270,N_12532);
or U13711 (N_13711,N_12557,N_12278);
or U13712 (N_13712,N_12241,N_12063);
or U13713 (N_13713,N_12874,N_12756);
xnor U13714 (N_13714,N_12823,N_12142);
xor U13715 (N_13715,N_12874,N_12255);
xor U13716 (N_13716,N_12088,N_12229);
or U13717 (N_13717,N_12551,N_12244);
nor U13718 (N_13718,N_12446,N_12911);
or U13719 (N_13719,N_12466,N_12709);
nor U13720 (N_13720,N_12916,N_12309);
xor U13721 (N_13721,N_12782,N_12166);
nor U13722 (N_13722,N_12269,N_12704);
nand U13723 (N_13723,N_12524,N_12088);
nand U13724 (N_13724,N_12243,N_12871);
nor U13725 (N_13725,N_12323,N_12822);
nand U13726 (N_13726,N_12266,N_12087);
and U13727 (N_13727,N_12337,N_12023);
or U13728 (N_13728,N_12720,N_12756);
xnor U13729 (N_13729,N_12638,N_12183);
or U13730 (N_13730,N_12023,N_12369);
xor U13731 (N_13731,N_12758,N_12004);
or U13732 (N_13732,N_12303,N_12797);
and U13733 (N_13733,N_12215,N_12122);
nor U13734 (N_13734,N_12820,N_12857);
xor U13735 (N_13735,N_12211,N_12278);
xnor U13736 (N_13736,N_12449,N_12188);
or U13737 (N_13737,N_12824,N_12597);
nand U13738 (N_13738,N_12211,N_12580);
nand U13739 (N_13739,N_12953,N_12474);
nand U13740 (N_13740,N_12285,N_12438);
nor U13741 (N_13741,N_12592,N_12359);
or U13742 (N_13742,N_12998,N_12069);
xor U13743 (N_13743,N_12612,N_12772);
and U13744 (N_13744,N_12904,N_12743);
xnor U13745 (N_13745,N_12092,N_12638);
or U13746 (N_13746,N_12639,N_12867);
nand U13747 (N_13747,N_12403,N_12593);
or U13748 (N_13748,N_12725,N_12223);
nor U13749 (N_13749,N_12831,N_12557);
xnor U13750 (N_13750,N_12499,N_12399);
and U13751 (N_13751,N_12037,N_12699);
nor U13752 (N_13752,N_12165,N_12750);
nand U13753 (N_13753,N_12573,N_12107);
and U13754 (N_13754,N_12581,N_12462);
or U13755 (N_13755,N_12377,N_12863);
nand U13756 (N_13756,N_12574,N_12139);
nand U13757 (N_13757,N_12923,N_12435);
or U13758 (N_13758,N_12013,N_12288);
or U13759 (N_13759,N_12430,N_12570);
or U13760 (N_13760,N_12233,N_12357);
nand U13761 (N_13761,N_12870,N_12090);
nand U13762 (N_13762,N_12695,N_12487);
nor U13763 (N_13763,N_12001,N_12331);
xor U13764 (N_13764,N_12766,N_12568);
xor U13765 (N_13765,N_12710,N_12356);
xnor U13766 (N_13766,N_12545,N_12586);
and U13767 (N_13767,N_12405,N_12755);
and U13768 (N_13768,N_12040,N_12514);
and U13769 (N_13769,N_12715,N_12625);
or U13770 (N_13770,N_12887,N_12161);
nand U13771 (N_13771,N_12837,N_12054);
nor U13772 (N_13772,N_12295,N_12201);
xor U13773 (N_13773,N_12247,N_12111);
or U13774 (N_13774,N_12486,N_12207);
or U13775 (N_13775,N_12046,N_12422);
nand U13776 (N_13776,N_12882,N_12099);
xor U13777 (N_13777,N_12836,N_12128);
or U13778 (N_13778,N_12868,N_12708);
nor U13779 (N_13779,N_12190,N_12139);
and U13780 (N_13780,N_12558,N_12349);
xnor U13781 (N_13781,N_12370,N_12405);
nand U13782 (N_13782,N_12639,N_12888);
nor U13783 (N_13783,N_12019,N_12493);
nand U13784 (N_13784,N_12054,N_12354);
and U13785 (N_13785,N_12429,N_12382);
or U13786 (N_13786,N_12156,N_12539);
xnor U13787 (N_13787,N_12334,N_12676);
nor U13788 (N_13788,N_12274,N_12833);
xor U13789 (N_13789,N_12406,N_12723);
nor U13790 (N_13790,N_12071,N_12379);
nand U13791 (N_13791,N_12933,N_12676);
xnor U13792 (N_13792,N_12367,N_12691);
or U13793 (N_13793,N_12017,N_12415);
nor U13794 (N_13794,N_12040,N_12853);
nand U13795 (N_13795,N_12254,N_12857);
xnor U13796 (N_13796,N_12640,N_12570);
nor U13797 (N_13797,N_12261,N_12898);
and U13798 (N_13798,N_12287,N_12182);
nand U13799 (N_13799,N_12132,N_12767);
nand U13800 (N_13800,N_12713,N_12317);
nand U13801 (N_13801,N_12615,N_12949);
nand U13802 (N_13802,N_12616,N_12961);
xor U13803 (N_13803,N_12731,N_12290);
nand U13804 (N_13804,N_12604,N_12972);
nand U13805 (N_13805,N_12671,N_12923);
nand U13806 (N_13806,N_12227,N_12352);
nand U13807 (N_13807,N_12620,N_12642);
nand U13808 (N_13808,N_12957,N_12662);
xor U13809 (N_13809,N_12007,N_12494);
and U13810 (N_13810,N_12024,N_12696);
nor U13811 (N_13811,N_12355,N_12801);
nand U13812 (N_13812,N_12263,N_12026);
nor U13813 (N_13813,N_12649,N_12192);
or U13814 (N_13814,N_12266,N_12649);
nor U13815 (N_13815,N_12206,N_12006);
xor U13816 (N_13816,N_12798,N_12929);
xnor U13817 (N_13817,N_12830,N_12118);
and U13818 (N_13818,N_12890,N_12975);
nor U13819 (N_13819,N_12838,N_12314);
and U13820 (N_13820,N_12716,N_12929);
nor U13821 (N_13821,N_12031,N_12713);
nand U13822 (N_13822,N_12521,N_12178);
and U13823 (N_13823,N_12120,N_12675);
nor U13824 (N_13824,N_12631,N_12284);
xnor U13825 (N_13825,N_12048,N_12029);
xnor U13826 (N_13826,N_12958,N_12756);
and U13827 (N_13827,N_12406,N_12708);
nor U13828 (N_13828,N_12650,N_12321);
and U13829 (N_13829,N_12053,N_12077);
nor U13830 (N_13830,N_12288,N_12034);
or U13831 (N_13831,N_12991,N_12621);
nand U13832 (N_13832,N_12933,N_12406);
nor U13833 (N_13833,N_12091,N_12095);
or U13834 (N_13834,N_12005,N_12177);
nand U13835 (N_13835,N_12129,N_12436);
xor U13836 (N_13836,N_12354,N_12266);
and U13837 (N_13837,N_12553,N_12839);
nand U13838 (N_13838,N_12706,N_12648);
or U13839 (N_13839,N_12945,N_12920);
xnor U13840 (N_13840,N_12749,N_12406);
nor U13841 (N_13841,N_12623,N_12961);
xnor U13842 (N_13842,N_12889,N_12444);
nor U13843 (N_13843,N_12240,N_12233);
or U13844 (N_13844,N_12792,N_12339);
nor U13845 (N_13845,N_12647,N_12611);
and U13846 (N_13846,N_12599,N_12127);
or U13847 (N_13847,N_12603,N_12199);
nor U13848 (N_13848,N_12100,N_12485);
and U13849 (N_13849,N_12246,N_12874);
nand U13850 (N_13850,N_12125,N_12639);
nor U13851 (N_13851,N_12088,N_12126);
nor U13852 (N_13852,N_12190,N_12952);
and U13853 (N_13853,N_12822,N_12633);
and U13854 (N_13854,N_12009,N_12781);
and U13855 (N_13855,N_12311,N_12483);
and U13856 (N_13856,N_12289,N_12436);
nand U13857 (N_13857,N_12976,N_12889);
and U13858 (N_13858,N_12295,N_12240);
xor U13859 (N_13859,N_12237,N_12957);
xor U13860 (N_13860,N_12974,N_12970);
xor U13861 (N_13861,N_12387,N_12230);
nor U13862 (N_13862,N_12253,N_12949);
nand U13863 (N_13863,N_12188,N_12363);
nor U13864 (N_13864,N_12115,N_12084);
nand U13865 (N_13865,N_12196,N_12947);
and U13866 (N_13866,N_12384,N_12820);
and U13867 (N_13867,N_12741,N_12823);
and U13868 (N_13868,N_12783,N_12305);
or U13869 (N_13869,N_12933,N_12912);
xnor U13870 (N_13870,N_12149,N_12251);
and U13871 (N_13871,N_12522,N_12537);
and U13872 (N_13872,N_12993,N_12185);
xor U13873 (N_13873,N_12431,N_12637);
nor U13874 (N_13874,N_12926,N_12284);
nor U13875 (N_13875,N_12971,N_12138);
or U13876 (N_13876,N_12833,N_12185);
or U13877 (N_13877,N_12762,N_12218);
and U13878 (N_13878,N_12851,N_12957);
and U13879 (N_13879,N_12870,N_12558);
nor U13880 (N_13880,N_12698,N_12464);
or U13881 (N_13881,N_12669,N_12558);
and U13882 (N_13882,N_12686,N_12921);
nor U13883 (N_13883,N_12499,N_12952);
xor U13884 (N_13884,N_12308,N_12356);
nand U13885 (N_13885,N_12073,N_12993);
and U13886 (N_13886,N_12307,N_12795);
xor U13887 (N_13887,N_12126,N_12968);
nand U13888 (N_13888,N_12377,N_12131);
xnor U13889 (N_13889,N_12246,N_12846);
or U13890 (N_13890,N_12984,N_12468);
nor U13891 (N_13891,N_12185,N_12086);
and U13892 (N_13892,N_12578,N_12352);
nor U13893 (N_13893,N_12106,N_12573);
xor U13894 (N_13894,N_12726,N_12091);
or U13895 (N_13895,N_12818,N_12121);
nand U13896 (N_13896,N_12131,N_12263);
nand U13897 (N_13897,N_12600,N_12487);
nand U13898 (N_13898,N_12439,N_12551);
xor U13899 (N_13899,N_12741,N_12531);
or U13900 (N_13900,N_12692,N_12509);
xor U13901 (N_13901,N_12779,N_12696);
or U13902 (N_13902,N_12030,N_12555);
nand U13903 (N_13903,N_12564,N_12314);
xnor U13904 (N_13904,N_12189,N_12659);
nor U13905 (N_13905,N_12699,N_12364);
nand U13906 (N_13906,N_12009,N_12037);
or U13907 (N_13907,N_12708,N_12655);
and U13908 (N_13908,N_12832,N_12596);
and U13909 (N_13909,N_12705,N_12897);
and U13910 (N_13910,N_12064,N_12045);
nand U13911 (N_13911,N_12693,N_12937);
nor U13912 (N_13912,N_12871,N_12889);
nor U13913 (N_13913,N_12219,N_12472);
nand U13914 (N_13914,N_12321,N_12206);
nor U13915 (N_13915,N_12205,N_12254);
xor U13916 (N_13916,N_12652,N_12592);
nand U13917 (N_13917,N_12849,N_12839);
xnor U13918 (N_13918,N_12147,N_12895);
xor U13919 (N_13919,N_12404,N_12146);
nor U13920 (N_13920,N_12559,N_12994);
or U13921 (N_13921,N_12499,N_12037);
or U13922 (N_13922,N_12848,N_12755);
nor U13923 (N_13923,N_12896,N_12711);
nor U13924 (N_13924,N_12732,N_12240);
xor U13925 (N_13925,N_12920,N_12087);
and U13926 (N_13926,N_12343,N_12915);
nor U13927 (N_13927,N_12428,N_12408);
nor U13928 (N_13928,N_12859,N_12397);
and U13929 (N_13929,N_12808,N_12212);
or U13930 (N_13930,N_12008,N_12616);
nand U13931 (N_13931,N_12574,N_12396);
and U13932 (N_13932,N_12443,N_12544);
xor U13933 (N_13933,N_12939,N_12609);
and U13934 (N_13934,N_12290,N_12427);
nand U13935 (N_13935,N_12693,N_12803);
xnor U13936 (N_13936,N_12297,N_12351);
nand U13937 (N_13937,N_12009,N_12250);
nor U13938 (N_13938,N_12513,N_12564);
nand U13939 (N_13939,N_12611,N_12083);
or U13940 (N_13940,N_12814,N_12477);
xor U13941 (N_13941,N_12811,N_12826);
nand U13942 (N_13942,N_12231,N_12949);
or U13943 (N_13943,N_12606,N_12548);
nand U13944 (N_13944,N_12700,N_12047);
or U13945 (N_13945,N_12089,N_12761);
or U13946 (N_13946,N_12277,N_12284);
or U13947 (N_13947,N_12734,N_12704);
xor U13948 (N_13948,N_12655,N_12646);
nor U13949 (N_13949,N_12257,N_12797);
nor U13950 (N_13950,N_12053,N_12385);
xor U13951 (N_13951,N_12437,N_12864);
and U13952 (N_13952,N_12645,N_12261);
nor U13953 (N_13953,N_12422,N_12502);
and U13954 (N_13954,N_12364,N_12916);
or U13955 (N_13955,N_12346,N_12241);
and U13956 (N_13956,N_12531,N_12176);
or U13957 (N_13957,N_12096,N_12396);
nand U13958 (N_13958,N_12777,N_12925);
nand U13959 (N_13959,N_12257,N_12438);
xnor U13960 (N_13960,N_12849,N_12038);
or U13961 (N_13961,N_12060,N_12812);
xnor U13962 (N_13962,N_12402,N_12041);
or U13963 (N_13963,N_12546,N_12257);
xor U13964 (N_13964,N_12627,N_12854);
and U13965 (N_13965,N_12614,N_12561);
nor U13966 (N_13966,N_12000,N_12155);
nor U13967 (N_13967,N_12081,N_12687);
xnor U13968 (N_13968,N_12637,N_12094);
nand U13969 (N_13969,N_12542,N_12845);
or U13970 (N_13970,N_12352,N_12958);
xor U13971 (N_13971,N_12026,N_12720);
nor U13972 (N_13972,N_12824,N_12002);
nand U13973 (N_13973,N_12032,N_12351);
or U13974 (N_13974,N_12967,N_12652);
xor U13975 (N_13975,N_12097,N_12032);
and U13976 (N_13976,N_12382,N_12802);
nor U13977 (N_13977,N_12378,N_12579);
nand U13978 (N_13978,N_12097,N_12978);
nand U13979 (N_13979,N_12040,N_12900);
nor U13980 (N_13980,N_12911,N_12117);
nor U13981 (N_13981,N_12465,N_12249);
and U13982 (N_13982,N_12242,N_12581);
nand U13983 (N_13983,N_12928,N_12061);
xnor U13984 (N_13984,N_12808,N_12307);
nand U13985 (N_13985,N_12128,N_12598);
and U13986 (N_13986,N_12644,N_12725);
and U13987 (N_13987,N_12007,N_12305);
xnor U13988 (N_13988,N_12314,N_12539);
and U13989 (N_13989,N_12466,N_12247);
nand U13990 (N_13990,N_12024,N_12595);
and U13991 (N_13991,N_12845,N_12124);
xor U13992 (N_13992,N_12582,N_12309);
or U13993 (N_13993,N_12951,N_12922);
nand U13994 (N_13994,N_12452,N_12304);
nand U13995 (N_13995,N_12798,N_12248);
xor U13996 (N_13996,N_12511,N_12175);
and U13997 (N_13997,N_12843,N_12989);
and U13998 (N_13998,N_12761,N_12093);
and U13999 (N_13999,N_12725,N_12041);
nor U14000 (N_14000,N_13121,N_13258);
nand U14001 (N_14001,N_13534,N_13846);
and U14002 (N_14002,N_13508,N_13942);
and U14003 (N_14003,N_13557,N_13022);
or U14004 (N_14004,N_13003,N_13189);
nor U14005 (N_14005,N_13608,N_13728);
nand U14006 (N_14006,N_13758,N_13722);
and U14007 (N_14007,N_13068,N_13230);
and U14008 (N_14008,N_13856,N_13625);
nor U14009 (N_14009,N_13226,N_13990);
nor U14010 (N_14010,N_13658,N_13998);
nor U14011 (N_14011,N_13347,N_13025);
nand U14012 (N_14012,N_13436,N_13523);
nand U14013 (N_14013,N_13339,N_13151);
or U14014 (N_14014,N_13575,N_13082);
nor U14015 (N_14015,N_13460,N_13772);
and U14016 (N_14016,N_13117,N_13449);
xor U14017 (N_14017,N_13703,N_13131);
nor U14018 (N_14018,N_13697,N_13964);
nor U14019 (N_14019,N_13743,N_13585);
or U14020 (N_14020,N_13317,N_13039);
and U14021 (N_14021,N_13096,N_13170);
nor U14022 (N_14022,N_13007,N_13443);
nor U14023 (N_14023,N_13052,N_13417);
xor U14024 (N_14024,N_13393,N_13564);
nand U14025 (N_14025,N_13403,N_13665);
nand U14026 (N_14026,N_13821,N_13828);
and U14027 (N_14027,N_13810,N_13362);
or U14028 (N_14028,N_13825,N_13934);
nor U14029 (N_14029,N_13136,N_13601);
nor U14030 (N_14030,N_13452,N_13023);
and U14031 (N_14031,N_13357,N_13955);
nor U14032 (N_14032,N_13962,N_13609);
nor U14033 (N_14033,N_13332,N_13373);
and U14034 (N_14034,N_13811,N_13526);
nand U14035 (N_14035,N_13192,N_13187);
or U14036 (N_14036,N_13790,N_13632);
xor U14037 (N_14037,N_13634,N_13866);
and U14038 (N_14038,N_13745,N_13066);
nand U14039 (N_14039,N_13574,N_13806);
or U14040 (N_14040,N_13454,N_13135);
xnor U14041 (N_14041,N_13392,N_13026);
nor U14042 (N_14042,N_13313,N_13893);
xnor U14043 (N_14043,N_13272,N_13252);
nor U14044 (N_14044,N_13982,N_13549);
nor U14045 (N_14045,N_13502,N_13820);
or U14046 (N_14046,N_13303,N_13276);
nor U14047 (N_14047,N_13660,N_13035);
and U14048 (N_14048,N_13544,N_13168);
xor U14049 (N_14049,N_13320,N_13232);
nor U14050 (N_14050,N_13986,N_13246);
xnor U14051 (N_14051,N_13744,N_13908);
and U14052 (N_14052,N_13217,N_13579);
and U14053 (N_14053,N_13591,N_13500);
xor U14054 (N_14054,N_13118,N_13006);
nor U14055 (N_14055,N_13331,N_13848);
or U14056 (N_14056,N_13756,N_13424);
nor U14057 (N_14057,N_13211,N_13802);
or U14058 (N_14058,N_13103,N_13376);
or U14059 (N_14059,N_13571,N_13905);
or U14060 (N_14060,N_13321,N_13953);
and U14061 (N_14061,N_13183,N_13688);
and U14062 (N_14062,N_13651,N_13568);
nand U14063 (N_14063,N_13817,N_13679);
nor U14064 (N_14064,N_13429,N_13140);
xor U14065 (N_14065,N_13027,N_13446);
or U14066 (N_14066,N_13784,N_13970);
nand U14067 (N_14067,N_13030,N_13778);
or U14068 (N_14068,N_13199,N_13723);
and U14069 (N_14069,N_13588,N_13713);
or U14070 (N_14070,N_13012,N_13130);
nand U14071 (N_14071,N_13898,N_13150);
xor U14072 (N_14072,N_13004,N_13092);
xor U14073 (N_14073,N_13350,N_13235);
and U14074 (N_14074,N_13620,N_13128);
or U14075 (N_14075,N_13786,N_13157);
xnor U14076 (N_14076,N_13611,N_13223);
or U14077 (N_14077,N_13663,N_13041);
xnor U14078 (N_14078,N_13038,N_13299);
and U14079 (N_14079,N_13268,N_13528);
and U14080 (N_14080,N_13408,N_13674);
nand U14081 (N_14081,N_13107,N_13553);
and U14082 (N_14082,N_13036,N_13055);
nor U14083 (N_14083,N_13203,N_13843);
or U14084 (N_14084,N_13971,N_13442);
nor U14085 (N_14085,N_13212,N_13421);
xor U14086 (N_14086,N_13488,N_13366);
nor U14087 (N_14087,N_13419,N_13180);
or U14088 (N_14088,N_13670,N_13532);
or U14089 (N_14089,N_13300,N_13239);
and U14090 (N_14090,N_13294,N_13716);
nand U14091 (N_14091,N_13434,N_13525);
nor U14092 (N_14092,N_13586,N_13791);
and U14093 (N_14093,N_13485,N_13682);
nor U14094 (N_14094,N_13943,N_13218);
or U14095 (N_14095,N_13542,N_13209);
and U14096 (N_14096,N_13378,N_13717);
xnor U14097 (N_14097,N_13928,N_13046);
xnor U14098 (N_14098,N_13512,N_13999);
nand U14099 (N_14099,N_13899,N_13067);
nor U14100 (N_14100,N_13139,N_13886);
nor U14101 (N_14101,N_13098,N_13750);
nand U14102 (N_14102,N_13636,N_13916);
or U14103 (N_14103,N_13288,N_13345);
nor U14104 (N_14104,N_13335,N_13177);
and U14105 (N_14105,N_13463,N_13677);
nor U14106 (N_14106,N_13584,N_13261);
or U14107 (N_14107,N_13946,N_13947);
and U14108 (N_14108,N_13680,N_13926);
nor U14109 (N_14109,N_13629,N_13324);
or U14110 (N_14110,N_13286,N_13256);
and U14111 (N_14111,N_13219,N_13240);
or U14112 (N_14112,N_13330,N_13543);
nor U14113 (N_14113,N_13097,N_13281);
nor U14114 (N_14114,N_13400,N_13872);
and U14115 (N_14115,N_13120,N_13237);
nor U14116 (N_14116,N_13101,N_13504);
or U14117 (N_14117,N_13334,N_13468);
or U14118 (N_14118,N_13126,N_13869);
nand U14119 (N_14119,N_13657,N_13250);
nor U14120 (N_14120,N_13667,N_13621);
or U14121 (N_14121,N_13381,N_13462);
xnor U14122 (N_14122,N_13989,N_13975);
or U14123 (N_14123,N_13257,N_13058);
or U14124 (N_14124,N_13389,N_13929);
or U14125 (N_14125,N_13056,N_13940);
nand U14126 (N_14126,N_13263,N_13777);
nand U14127 (N_14127,N_13995,N_13490);
nand U14128 (N_14128,N_13708,N_13640);
and U14129 (N_14129,N_13382,N_13517);
and U14130 (N_14130,N_13656,N_13262);
and U14131 (N_14131,N_13701,N_13086);
xnor U14132 (N_14132,N_13450,N_13984);
or U14133 (N_14133,N_13764,N_13896);
and U14134 (N_14134,N_13622,N_13844);
nor U14135 (N_14135,N_13433,N_13072);
nor U14136 (N_14136,N_13234,N_13838);
nor U14137 (N_14137,N_13789,N_13099);
or U14138 (N_14138,N_13581,N_13205);
xnor U14139 (N_14139,N_13228,N_13597);
nor U14140 (N_14140,N_13633,N_13312);
xnor U14141 (N_14141,N_13912,N_13141);
or U14142 (N_14142,N_13801,N_13319);
nand U14143 (N_14143,N_13705,N_13116);
xnor U14144 (N_14144,N_13457,N_13973);
or U14145 (N_14145,N_13236,N_13779);
xnor U14146 (N_14146,N_13043,N_13951);
xnor U14147 (N_14147,N_13618,N_13333);
nor U14148 (N_14148,N_13000,N_13143);
and U14149 (N_14149,N_13095,N_13418);
nor U14150 (N_14150,N_13184,N_13133);
xnor U14151 (N_14151,N_13994,N_13010);
xnor U14152 (N_14152,N_13650,N_13692);
and U14153 (N_14153,N_13461,N_13686);
and U14154 (N_14154,N_13241,N_13159);
or U14155 (N_14155,N_13675,N_13496);
or U14156 (N_14156,N_13985,N_13215);
xor U14157 (N_14157,N_13751,N_13522);
xor U14158 (N_14158,N_13198,N_13638);
and U14159 (N_14159,N_13882,N_13507);
and U14160 (N_14160,N_13037,N_13351);
or U14161 (N_14161,N_13933,N_13914);
xor U14162 (N_14162,N_13011,N_13693);
or U14163 (N_14163,N_13439,N_13747);
and U14164 (N_14164,N_13001,N_13570);
nand U14165 (N_14165,N_13200,N_13405);
and U14166 (N_14166,N_13616,N_13935);
or U14167 (N_14167,N_13009,N_13605);
nand U14168 (N_14168,N_13353,N_13997);
nor U14169 (N_14169,N_13280,N_13029);
nand U14170 (N_14170,N_13706,N_13541);
and U14171 (N_14171,N_13832,N_13370);
xor U14172 (N_14172,N_13254,N_13104);
or U14173 (N_14173,N_13737,N_13840);
xnor U14174 (N_14174,N_13194,N_13475);
xor U14175 (N_14175,N_13152,N_13146);
xnor U14176 (N_14176,N_13440,N_13260);
or U14177 (N_14177,N_13163,N_13432);
or U14178 (N_14178,N_13923,N_13020);
or U14179 (N_14179,N_13878,N_13155);
nand U14180 (N_14180,N_13578,N_13941);
and U14181 (N_14181,N_13494,N_13814);
nor U14182 (N_14182,N_13782,N_13719);
nand U14183 (N_14183,N_13191,N_13111);
or U14184 (N_14184,N_13057,N_13799);
and U14185 (N_14185,N_13438,N_13593);
xor U14186 (N_14186,N_13944,N_13253);
xnor U14187 (N_14187,N_13694,N_13304);
nand U14188 (N_14188,N_13493,N_13404);
nor U14189 (N_14189,N_13380,N_13561);
nand U14190 (N_14190,N_13078,N_13792);
and U14191 (N_14191,N_13961,N_13486);
or U14192 (N_14192,N_13042,N_13277);
or U14193 (N_14193,N_13793,N_13920);
and U14194 (N_14194,N_13283,N_13064);
nor U14195 (N_14195,N_13375,N_13388);
xor U14196 (N_14196,N_13904,N_13599);
xnor U14197 (N_14197,N_13800,N_13510);
xnor U14198 (N_14198,N_13562,N_13374);
nand U14199 (N_14199,N_13453,N_13148);
and U14200 (N_14200,N_13501,N_13604);
or U14201 (N_14201,N_13641,N_13652);
nor U14202 (N_14202,N_13063,N_13515);
or U14203 (N_14203,N_13711,N_13887);
and U14204 (N_14204,N_13024,N_13348);
xor U14205 (N_14205,N_13478,N_13114);
nand U14206 (N_14206,N_13760,N_13013);
and U14207 (N_14207,N_13213,N_13295);
nor U14208 (N_14208,N_13214,N_13090);
xnor U14209 (N_14209,N_13119,N_13169);
nor U14210 (N_14210,N_13748,N_13470);
and U14211 (N_14211,N_13956,N_13019);
xor U14212 (N_14212,N_13612,N_13459);
xnor U14213 (N_14213,N_13482,N_13144);
or U14214 (N_14214,N_13134,N_13977);
nand U14215 (N_14215,N_13885,N_13165);
xor U14216 (N_14216,N_13091,N_13726);
xor U14217 (N_14217,N_13979,N_13361);
or U14218 (N_14218,N_13922,N_13520);
xnor U14219 (N_14219,N_13505,N_13852);
and U14220 (N_14220,N_13524,N_13040);
and U14221 (N_14221,N_13769,N_13336);
nor U14222 (N_14222,N_13857,N_13600);
or U14223 (N_14223,N_13383,N_13603);
nor U14224 (N_14224,N_13506,N_13385);
nor U14225 (N_14225,N_13771,N_13664);
nand U14226 (N_14226,N_13907,N_13306);
or U14227 (N_14227,N_13059,N_13645);
and U14228 (N_14228,N_13499,N_13826);
xnor U14229 (N_14229,N_13630,N_13161);
nand U14230 (N_14230,N_13685,N_13873);
xnor U14231 (N_14231,N_13687,N_13394);
nor U14232 (N_14232,N_13053,N_13412);
nor U14233 (N_14233,N_13842,N_13164);
or U14234 (N_14234,N_13270,N_13195);
and U14235 (N_14235,N_13476,N_13572);
nor U14236 (N_14236,N_13206,N_13867);
and U14237 (N_14237,N_13709,N_13302);
xnor U14238 (N_14238,N_13619,N_13550);
nand U14239 (N_14239,N_13487,N_13837);
or U14240 (N_14240,N_13396,N_13070);
nor U14241 (N_14241,N_13647,N_13427);
nand U14242 (N_14242,N_13365,N_13316);
nand U14243 (N_14243,N_13113,N_13906);
xor U14244 (N_14244,N_13950,N_13305);
nand U14245 (N_14245,N_13736,N_13558);
and U14246 (N_14246,N_13227,N_13346);
xor U14247 (N_14247,N_13759,N_13624);
xor U14248 (N_14248,N_13435,N_13340);
xnor U14249 (N_14249,N_13202,N_13422);
nor U14250 (N_14250,N_13224,N_13749);
nand U14251 (N_14251,N_13819,N_13479);
xor U14252 (N_14252,N_13871,N_13993);
and U14253 (N_14253,N_13939,N_13966);
and U14254 (N_14254,N_13513,N_13077);
nand U14255 (N_14255,N_13798,N_13530);
xnor U14256 (N_14256,N_13691,N_13822);
xor U14257 (N_14257,N_13690,N_13655);
xnor U14258 (N_14258,N_13560,N_13216);
nor U14259 (N_14259,N_13718,N_13061);
and U14260 (N_14260,N_13102,N_13518);
or U14261 (N_14261,N_13326,N_13160);
nor U14262 (N_14262,N_13293,N_13841);
nand U14263 (N_14263,N_13124,N_13387);
or U14264 (N_14264,N_13983,N_13492);
nor U14265 (N_14265,N_13894,N_13839);
and U14266 (N_14266,N_13830,N_13631);
nand U14267 (N_14267,N_13654,N_13472);
xnor U14268 (N_14268,N_13770,N_13967);
nand U14269 (N_14269,N_13936,N_13712);
or U14270 (N_14270,N_13426,N_13125);
nand U14271 (N_14271,N_13238,N_13005);
nor U14272 (N_14272,N_13489,N_13372);
nand U14273 (N_14273,N_13423,N_13746);
nor U14274 (N_14274,N_13643,N_13661);
xor U14275 (N_14275,N_13519,N_13430);
nor U14276 (N_14276,N_13264,N_13509);
or U14277 (N_14277,N_13108,N_13795);
and U14278 (N_14278,N_13364,N_13291);
nand U14279 (N_14279,N_13269,N_13755);
nand U14280 (N_14280,N_13444,N_13411);
or U14281 (N_14281,N_13610,N_13642);
xor U14282 (N_14282,N_13399,N_13740);
xnor U14283 (N_14283,N_13473,N_13699);
or U14284 (N_14284,N_13456,N_13106);
xor U14285 (N_14285,N_13329,N_13352);
nor U14286 (N_14286,N_13721,N_13927);
and U14287 (N_14287,N_13285,N_13780);
or U14288 (N_14288,N_13368,N_13458);
and U14289 (N_14289,N_13613,N_13002);
xnor U14290 (N_14290,N_13915,N_13049);
or U14291 (N_14291,N_13868,N_13583);
nand U14292 (N_14292,N_13021,N_13308);
and U14293 (N_14293,N_13958,N_13358);
nand U14294 (N_14294,N_13765,N_13676);
nand U14295 (N_14295,N_13715,N_13949);
xnor U14296 (N_14296,N_13018,N_13930);
or U14297 (N_14297,N_13384,N_13259);
or U14298 (N_14298,N_13137,N_13084);
or U14299 (N_14299,N_13531,N_13757);
nor U14300 (N_14300,N_13807,N_13957);
and U14301 (N_14301,N_13328,N_13987);
nand U14302 (N_14302,N_13210,N_13356);
xor U14303 (N_14303,N_13533,N_13537);
nor U14304 (N_14304,N_13729,N_13555);
or U14305 (N_14305,N_13589,N_13242);
and U14306 (N_14306,N_13190,N_13379);
nor U14307 (N_14307,N_13733,N_13919);
and U14308 (N_14308,N_13441,N_13794);
xor U14309 (N_14309,N_13592,N_13309);
and U14310 (N_14310,N_13698,N_13323);
nor U14311 (N_14311,N_13892,N_13292);
or U14312 (N_14312,N_13415,N_13535);
xor U14313 (N_14313,N_13051,N_13607);
xor U14314 (N_14314,N_13017,N_13902);
nor U14315 (N_14315,N_13925,N_13074);
xor U14316 (N_14316,N_13414,N_13428);
nand U14317 (N_14317,N_13753,N_13363);
nor U14318 (N_14318,N_13796,N_13731);
nor U14319 (N_14319,N_13179,N_13673);
xor U14320 (N_14320,N_13244,N_13204);
nand U14321 (N_14321,N_13644,N_13559);
or U14322 (N_14322,N_13273,N_13813);
or U14323 (N_14323,N_13781,N_13766);
xor U14324 (N_14324,N_13833,N_13797);
and U14325 (N_14325,N_13044,N_13367);
nor U14326 (N_14326,N_13890,N_13371);
xnor U14327 (N_14327,N_13884,N_13511);
nand U14328 (N_14328,N_13845,N_13808);
xor U14329 (N_14329,N_13249,N_13596);
or U14330 (N_14330,N_13752,N_13567);
or U14331 (N_14331,N_13566,N_13425);
nand U14332 (N_14332,N_13287,N_13901);
or U14333 (N_14333,N_13094,N_13071);
or U14334 (N_14334,N_13700,N_13980);
and U14335 (N_14335,N_13937,N_13594);
xnor U14336 (N_14336,N_13623,N_13344);
xor U14337 (N_14337,N_13318,N_13521);
xnor U14338 (N_14338,N_13762,N_13938);
or U14339 (N_14339,N_13341,N_13627);
and U14340 (N_14340,N_13034,N_13684);
xnor U14341 (N_14341,N_13854,N_13327);
nor U14342 (N_14342,N_13342,N_13181);
and U14343 (N_14343,N_13858,N_13727);
xnor U14344 (N_14344,N_13863,N_13577);
or U14345 (N_14345,N_13835,N_13590);
or U14346 (N_14346,N_13420,N_13875);
xor U14347 (N_14347,N_13477,N_13451);
xnor U14348 (N_14348,N_13231,N_13805);
nand U14349 (N_14349,N_13491,N_13818);
nand U14350 (N_14350,N_13208,N_13307);
or U14351 (N_14351,N_13255,N_13836);
xor U14352 (N_14352,N_13127,N_13816);
and U14353 (N_14353,N_13666,N_13669);
xor U14354 (N_14354,N_13156,N_13891);
or U14355 (N_14355,N_13062,N_13773);
and U14356 (N_14356,N_13474,N_13761);
nand U14357 (N_14357,N_13547,N_13881);
and U14358 (N_14358,N_13297,N_13917);
or U14359 (N_14359,N_13483,N_13138);
nor U14360 (N_14360,N_13088,N_13573);
nor U14361 (N_14361,N_13960,N_13909);
nand U14362 (N_14362,N_13724,N_13267);
nor U14363 (N_14363,N_13710,N_13870);
nor U14364 (N_14364,N_13683,N_13552);
nand U14365 (N_14365,N_13668,N_13048);
or U14366 (N_14366,N_13447,N_13734);
nor U14367 (N_14367,N_13681,N_13377);
and U14368 (N_14368,N_13851,N_13355);
xor U14369 (N_14369,N_13471,N_13431);
nor U14370 (N_14370,N_13824,N_13275);
nor U14371 (N_14371,N_13315,N_13991);
and U14372 (N_14372,N_13158,N_13981);
or U14373 (N_14373,N_13188,N_13900);
and U14374 (N_14374,N_13672,N_13847);
or U14375 (N_14375,N_13274,N_13085);
nor U14376 (N_14376,N_13783,N_13897);
nor U14377 (N_14377,N_13110,N_13207);
and U14378 (N_14378,N_13338,N_13948);
xor U14379 (N_14379,N_13033,N_13812);
and U14380 (N_14380,N_13696,N_13735);
and U14381 (N_14381,N_13154,N_13831);
nand U14382 (N_14382,N_13069,N_13083);
nor U14383 (N_14383,N_13322,N_13678);
nand U14384 (N_14384,N_13861,N_13081);
xor U14385 (N_14385,N_13360,N_13529);
and U14386 (N_14386,N_13289,N_13464);
xor U14387 (N_14387,N_13193,N_13173);
nand U14388 (N_14388,N_13266,N_13182);
nand U14389 (N_14389,N_13437,N_13284);
nand U14390 (N_14390,N_13538,N_13197);
and U14391 (N_14391,N_13162,N_13112);
or U14392 (N_14392,N_13093,N_13409);
and U14393 (N_14393,N_13637,N_13580);
and U14394 (N_14394,N_13167,N_13815);
or U14395 (N_14395,N_13546,N_13123);
nor U14396 (N_14396,N_13480,N_13185);
and U14397 (N_14397,N_13540,N_13498);
or U14398 (N_14398,N_13245,N_13413);
or U14399 (N_14399,N_13497,N_13369);
xor U14400 (N_14400,N_13662,N_13763);
nand U14401 (N_14401,N_13271,N_13115);
nand U14402 (N_14402,N_13576,N_13298);
or U14403 (N_14403,N_13563,N_13787);
nand U14404 (N_14404,N_13877,N_13626);
nor U14405 (N_14405,N_13100,N_13406);
xor U14406 (N_14406,N_13996,N_13073);
and U14407 (N_14407,N_13864,N_13767);
xnor U14408 (N_14408,N_13014,N_13895);
nor U14409 (N_14409,N_13391,N_13602);
xor U14410 (N_14410,N_13968,N_13648);
xnor U14411 (N_14411,N_13466,N_13495);
and U14412 (N_14412,N_13467,N_13876);
nand U14413 (N_14413,N_13883,N_13075);
nand U14414 (N_14414,N_13754,N_13774);
nor U14415 (N_14415,N_13028,N_13978);
nand U14416 (N_14416,N_13397,N_13880);
nor U14417 (N_14417,N_13176,N_13296);
or U14418 (N_14418,N_13888,N_13527);
nor U14419 (N_14419,N_13079,N_13015);
nor U14420 (N_14420,N_13065,N_13974);
nand U14421 (N_14421,N_13448,N_13775);
and U14422 (N_14422,N_13776,N_13704);
nand U14423 (N_14423,N_13233,N_13416);
xor U14424 (N_14424,N_13145,N_13702);
xnor U14425 (N_14425,N_13398,N_13243);
nor U14426 (N_14426,N_13972,N_13465);
and U14427 (N_14427,N_13301,N_13646);
xnor U14428 (N_14428,N_13337,N_13325);
or U14429 (N_14429,N_13860,N_13707);
xor U14430 (N_14430,N_13889,N_13865);
xnor U14431 (N_14431,N_13080,N_13788);
and U14432 (N_14432,N_13032,N_13314);
or U14433 (N_14433,N_13615,N_13829);
and U14434 (N_14434,N_13122,N_13768);
or U14435 (N_14435,N_13407,N_13689);
or U14436 (N_14436,N_13220,N_13595);
or U14437 (N_14437,N_13859,N_13175);
or U14438 (N_14438,N_13047,N_13222);
xor U14439 (N_14439,N_13171,N_13988);
nand U14440 (N_14440,N_13054,N_13952);
nand U14441 (N_14441,N_13401,N_13551);
nand U14442 (N_14442,N_13201,N_13910);
and U14443 (N_14443,N_13045,N_13834);
and U14444 (N_14444,N_13554,N_13849);
xor U14445 (N_14445,N_13390,N_13142);
nor U14446 (N_14446,N_13963,N_13539);
or U14447 (N_14447,N_13251,N_13247);
or U14448 (N_14448,N_13969,N_13395);
and U14449 (N_14449,N_13178,N_13659);
xnor U14450 (N_14450,N_13265,N_13714);
nand U14451 (N_14451,N_13153,N_13921);
nor U14452 (N_14452,N_13639,N_13862);
xnor U14453 (N_14453,N_13536,N_13653);
xnor U14454 (N_14454,N_13671,N_13924);
nand U14455 (N_14455,N_13730,N_13785);
and U14456 (N_14456,N_13410,N_13565);
and U14457 (N_14457,N_13354,N_13087);
xnor U14458 (N_14458,N_13076,N_13455);
xnor U14459 (N_14459,N_13548,N_13649);
xnor U14460 (N_14460,N_13050,N_13628);
nor U14461 (N_14461,N_13614,N_13598);
nor U14462 (N_14462,N_13976,N_13959);
or U14463 (N_14463,N_13514,N_13359);
and U14464 (N_14464,N_13732,N_13954);
xnor U14465 (N_14465,N_13918,N_13343);
and U14466 (N_14466,N_13469,N_13809);
xnor U14467 (N_14467,N_13008,N_13932);
xnor U14468 (N_14468,N_13016,N_13349);
nand U14469 (N_14469,N_13742,N_13248);
or U14470 (N_14470,N_13481,N_13725);
nand U14471 (N_14471,N_13186,N_13804);
and U14472 (N_14472,N_13617,N_13166);
xnor U14473 (N_14473,N_13503,N_13738);
nor U14474 (N_14474,N_13229,N_13402);
xor U14475 (N_14475,N_13720,N_13741);
nor U14476 (N_14476,N_13911,N_13582);
nand U14477 (N_14477,N_13635,N_13132);
xor U14478 (N_14478,N_13445,N_13282);
or U14479 (N_14479,N_13739,N_13903);
and U14480 (N_14480,N_13105,N_13129);
nor U14481 (N_14481,N_13879,N_13278);
nand U14482 (N_14482,N_13587,N_13089);
xor U14483 (N_14483,N_13569,N_13109);
xnor U14484 (N_14484,N_13221,N_13545);
and U14485 (N_14485,N_13031,N_13174);
or U14486 (N_14486,N_13225,N_13149);
or U14487 (N_14487,N_13855,N_13853);
and U14488 (N_14488,N_13606,N_13945);
nor U14489 (N_14489,N_13992,N_13310);
or U14490 (N_14490,N_13147,N_13516);
xnor U14491 (N_14491,N_13823,N_13827);
nor U14492 (N_14492,N_13279,N_13196);
nor U14493 (N_14493,N_13386,N_13556);
xor U14494 (N_14494,N_13311,N_13803);
nand U14495 (N_14495,N_13874,N_13965);
xor U14496 (N_14496,N_13060,N_13931);
nand U14497 (N_14497,N_13695,N_13172);
and U14498 (N_14498,N_13850,N_13913);
nand U14499 (N_14499,N_13484,N_13290);
xor U14500 (N_14500,N_13813,N_13900);
and U14501 (N_14501,N_13072,N_13695);
nor U14502 (N_14502,N_13998,N_13027);
and U14503 (N_14503,N_13699,N_13370);
xnor U14504 (N_14504,N_13254,N_13898);
nor U14505 (N_14505,N_13445,N_13609);
and U14506 (N_14506,N_13501,N_13463);
xor U14507 (N_14507,N_13939,N_13594);
and U14508 (N_14508,N_13426,N_13334);
xnor U14509 (N_14509,N_13558,N_13125);
and U14510 (N_14510,N_13646,N_13481);
xor U14511 (N_14511,N_13718,N_13406);
xnor U14512 (N_14512,N_13545,N_13790);
or U14513 (N_14513,N_13681,N_13726);
and U14514 (N_14514,N_13718,N_13470);
or U14515 (N_14515,N_13858,N_13706);
xnor U14516 (N_14516,N_13850,N_13955);
xor U14517 (N_14517,N_13824,N_13924);
and U14518 (N_14518,N_13474,N_13599);
and U14519 (N_14519,N_13483,N_13215);
xnor U14520 (N_14520,N_13606,N_13532);
nor U14521 (N_14521,N_13782,N_13838);
nor U14522 (N_14522,N_13411,N_13275);
nand U14523 (N_14523,N_13665,N_13998);
and U14524 (N_14524,N_13849,N_13947);
or U14525 (N_14525,N_13060,N_13795);
xor U14526 (N_14526,N_13174,N_13438);
or U14527 (N_14527,N_13950,N_13149);
or U14528 (N_14528,N_13986,N_13952);
or U14529 (N_14529,N_13993,N_13228);
nand U14530 (N_14530,N_13771,N_13638);
and U14531 (N_14531,N_13316,N_13039);
or U14532 (N_14532,N_13499,N_13500);
nand U14533 (N_14533,N_13522,N_13511);
xor U14534 (N_14534,N_13587,N_13221);
and U14535 (N_14535,N_13513,N_13315);
nand U14536 (N_14536,N_13302,N_13079);
nand U14537 (N_14537,N_13199,N_13932);
and U14538 (N_14538,N_13316,N_13768);
nand U14539 (N_14539,N_13952,N_13572);
and U14540 (N_14540,N_13147,N_13370);
nand U14541 (N_14541,N_13635,N_13539);
xor U14542 (N_14542,N_13783,N_13633);
xnor U14543 (N_14543,N_13752,N_13732);
or U14544 (N_14544,N_13752,N_13709);
or U14545 (N_14545,N_13670,N_13239);
and U14546 (N_14546,N_13175,N_13949);
or U14547 (N_14547,N_13313,N_13702);
xor U14548 (N_14548,N_13766,N_13017);
and U14549 (N_14549,N_13475,N_13985);
nor U14550 (N_14550,N_13140,N_13251);
xor U14551 (N_14551,N_13000,N_13911);
nor U14552 (N_14552,N_13670,N_13350);
nand U14553 (N_14553,N_13683,N_13169);
nand U14554 (N_14554,N_13313,N_13552);
nand U14555 (N_14555,N_13654,N_13784);
or U14556 (N_14556,N_13381,N_13606);
and U14557 (N_14557,N_13678,N_13828);
or U14558 (N_14558,N_13076,N_13530);
xnor U14559 (N_14559,N_13629,N_13864);
or U14560 (N_14560,N_13465,N_13757);
or U14561 (N_14561,N_13057,N_13263);
or U14562 (N_14562,N_13954,N_13045);
xor U14563 (N_14563,N_13273,N_13118);
xnor U14564 (N_14564,N_13846,N_13528);
nor U14565 (N_14565,N_13792,N_13157);
nand U14566 (N_14566,N_13868,N_13760);
nor U14567 (N_14567,N_13029,N_13605);
and U14568 (N_14568,N_13238,N_13415);
and U14569 (N_14569,N_13457,N_13603);
and U14570 (N_14570,N_13541,N_13191);
nor U14571 (N_14571,N_13008,N_13246);
nor U14572 (N_14572,N_13654,N_13918);
and U14573 (N_14573,N_13653,N_13172);
or U14574 (N_14574,N_13886,N_13649);
xnor U14575 (N_14575,N_13098,N_13192);
nand U14576 (N_14576,N_13715,N_13052);
and U14577 (N_14577,N_13897,N_13179);
nand U14578 (N_14578,N_13538,N_13474);
or U14579 (N_14579,N_13552,N_13252);
or U14580 (N_14580,N_13027,N_13865);
nor U14581 (N_14581,N_13539,N_13103);
and U14582 (N_14582,N_13012,N_13975);
nand U14583 (N_14583,N_13690,N_13842);
xnor U14584 (N_14584,N_13645,N_13988);
xnor U14585 (N_14585,N_13488,N_13729);
and U14586 (N_14586,N_13783,N_13112);
or U14587 (N_14587,N_13919,N_13687);
or U14588 (N_14588,N_13193,N_13309);
and U14589 (N_14589,N_13668,N_13654);
nand U14590 (N_14590,N_13934,N_13445);
and U14591 (N_14591,N_13294,N_13544);
or U14592 (N_14592,N_13975,N_13593);
xor U14593 (N_14593,N_13517,N_13635);
or U14594 (N_14594,N_13185,N_13093);
nor U14595 (N_14595,N_13815,N_13371);
nand U14596 (N_14596,N_13213,N_13952);
or U14597 (N_14597,N_13284,N_13640);
nor U14598 (N_14598,N_13932,N_13803);
nor U14599 (N_14599,N_13856,N_13983);
xor U14600 (N_14600,N_13259,N_13711);
xnor U14601 (N_14601,N_13763,N_13821);
and U14602 (N_14602,N_13510,N_13180);
nand U14603 (N_14603,N_13645,N_13202);
nand U14604 (N_14604,N_13527,N_13253);
and U14605 (N_14605,N_13141,N_13941);
nand U14606 (N_14606,N_13056,N_13899);
xnor U14607 (N_14607,N_13080,N_13228);
nand U14608 (N_14608,N_13564,N_13804);
and U14609 (N_14609,N_13640,N_13516);
xnor U14610 (N_14610,N_13346,N_13827);
nor U14611 (N_14611,N_13739,N_13128);
nor U14612 (N_14612,N_13504,N_13659);
xor U14613 (N_14613,N_13271,N_13122);
and U14614 (N_14614,N_13252,N_13897);
xnor U14615 (N_14615,N_13868,N_13844);
or U14616 (N_14616,N_13928,N_13366);
and U14617 (N_14617,N_13319,N_13008);
nand U14618 (N_14618,N_13171,N_13533);
and U14619 (N_14619,N_13108,N_13695);
or U14620 (N_14620,N_13831,N_13854);
and U14621 (N_14621,N_13825,N_13210);
nand U14622 (N_14622,N_13578,N_13820);
nand U14623 (N_14623,N_13308,N_13919);
nand U14624 (N_14624,N_13431,N_13953);
nand U14625 (N_14625,N_13232,N_13426);
nand U14626 (N_14626,N_13236,N_13264);
and U14627 (N_14627,N_13892,N_13118);
xor U14628 (N_14628,N_13628,N_13521);
xnor U14629 (N_14629,N_13270,N_13392);
nand U14630 (N_14630,N_13384,N_13753);
and U14631 (N_14631,N_13879,N_13011);
xnor U14632 (N_14632,N_13584,N_13044);
xor U14633 (N_14633,N_13788,N_13621);
nor U14634 (N_14634,N_13397,N_13679);
or U14635 (N_14635,N_13561,N_13693);
nor U14636 (N_14636,N_13392,N_13028);
nor U14637 (N_14637,N_13697,N_13071);
or U14638 (N_14638,N_13898,N_13850);
nand U14639 (N_14639,N_13514,N_13616);
xor U14640 (N_14640,N_13876,N_13533);
or U14641 (N_14641,N_13238,N_13186);
and U14642 (N_14642,N_13719,N_13237);
or U14643 (N_14643,N_13218,N_13572);
or U14644 (N_14644,N_13336,N_13238);
and U14645 (N_14645,N_13703,N_13369);
or U14646 (N_14646,N_13714,N_13503);
or U14647 (N_14647,N_13034,N_13891);
nand U14648 (N_14648,N_13745,N_13855);
or U14649 (N_14649,N_13731,N_13153);
or U14650 (N_14650,N_13374,N_13307);
nor U14651 (N_14651,N_13077,N_13849);
and U14652 (N_14652,N_13238,N_13795);
xnor U14653 (N_14653,N_13468,N_13785);
and U14654 (N_14654,N_13785,N_13461);
xnor U14655 (N_14655,N_13928,N_13779);
or U14656 (N_14656,N_13331,N_13515);
nand U14657 (N_14657,N_13949,N_13218);
or U14658 (N_14658,N_13507,N_13982);
nor U14659 (N_14659,N_13505,N_13798);
or U14660 (N_14660,N_13188,N_13654);
xnor U14661 (N_14661,N_13758,N_13274);
nand U14662 (N_14662,N_13559,N_13377);
nor U14663 (N_14663,N_13596,N_13062);
xor U14664 (N_14664,N_13195,N_13929);
and U14665 (N_14665,N_13186,N_13827);
nor U14666 (N_14666,N_13985,N_13548);
xor U14667 (N_14667,N_13399,N_13255);
and U14668 (N_14668,N_13831,N_13581);
nand U14669 (N_14669,N_13448,N_13484);
or U14670 (N_14670,N_13802,N_13461);
nand U14671 (N_14671,N_13156,N_13294);
nor U14672 (N_14672,N_13250,N_13880);
xnor U14673 (N_14673,N_13497,N_13561);
nor U14674 (N_14674,N_13842,N_13371);
and U14675 (N_14675,N_13738,N_13336);
nand U14676 (N_14676,N_13080,N_13166);
xnor U14677 (N_14677,N_13276,N_13548);
nor U14678 (N_14678,N_13680,N_13280);
or U14679 (N_14679,N_13655,N_13971);
and U14680 (N_14680,N_13596,N_13842);
nor U14681 (N_14681,N_13602,N_13927);
nand U14682 (N_14682,N_13282,N_13249);
or U14683 (N_14683,N_13298,N_13879);
and U14684 (N_14684,N_13993,N_13755);
nor U14685 (N_14685,N_13357,N_13901);
nor U14686 (N_14686,N_13516,N_13597);
or U14687 (N_14687,N_13580,N_13888);
nor U14688 (N_14688,N_13081,N_13020);
or U14689 (N_14689,N_13614,N_13242);
and U14690 (N_14690,N_13567,N_13993);
nand U14691 (N_14691,N_13273,N_13357);
or U14692 (N_14692,N_13384,N_13437);
nor U14693 (N_14693,N_13703,N_13315);
xnor U14694 (N_14694,N_13336,N_13791);
and U14695 (N_14695,N_13205,N_13412);
and U14696 (N_14696,N_13892,N_13929);
xor U14697 (N_14697,N_13012,N_13913);
xor U14698 (N_14698,N_13225,N_13831);
xor U14699 (N_14699,N_13950,N_13279);
nand U14700 (N_14700,N_13749,N_13047);
nor U14701 (N_14701,N_13904,N_13168);
nor U14702 (N_14702,N_13915,N_13586);
and U14703 (N_14703,N_13634,N_13454);
and U14704 (N_14704,N_13924,N_13118);
and U14705 (N_14705,N_13285,N_13255);
nor U14706 (N_14706,N_13532,N_13123);
xnor U14707 (N_14707,N_13310,N_13584);
nand U14708 (N_14708,N_13192,N_13180);
xor U14709 (N_14709,N_13880,N_13802);
nor U14710 (N_14710,N_13541,N_13088);
nand U14711 (N_14711,N_13774,N_13354);
and U14712 (N_14712,N_13535,N_13706);
or U14713 (N_14713,N_13778,N_13122);
nor U14714 (N_14714,N_13411,N_13216);
nand U14715 (N_14715,N_13222,N_13085);
xnor U14716 (N_14716,N_13398,N_13106);
nor U14717 (N_14717,N_13320,N_13056);
and U14718 (N_14718,N_13037,N_13779);
nand U14719 (N_14719,N_13563,N_13102);
nor U14720 (N_14720,N_13232,N_13675);
and U14721 (N_14721,N_13394,N_13615);
and U14722 (N_14722,N_13931,N_13209);
nand U14723 (N_14723,N_13123,N_13976);
xnor U14724 (N_14724,N_13284,N_13917);
and U14725 (N_14725,N_13669,N_13920);
nand U14726 (N_14726,N_13496,N_13186);
nand U14727 (N_14727,N_13683,N_13455);
or U14728 (N_14728,N_13195,N_13180);
xor U14729 (N_14729,N_13414,N_13830);
nand U14730 (N_14730,N_13698,N_13884);
xnor U14731 (N_14731,N_13389,N_13317);
nor U14732 (N_14732,N_13363,N_13142);
xor U14733 (N_14733,N_13052,N_13460);
nand U14734 (N_14734,N_13107,N_13886);
nor U14735 (N_14735,N_13923,N_13322);
nor U14736 (N_14736,N_13599,N_13109);
nand U14737 (N_14737,N_13397,N_13945);
xnor U14738 (N_14738,N_13893,N_13842);
xnor U14739 (N_14739,N_13133,N_13900);
nand U14740 (N_14740,N_13790,N_13860);
nand U14741 (N_14741,N_13396,N_13507);
or U14742 (N_14742,N_13608,N_13059);
nor U14743 (N_14743,N_13903,N_13896);
and U14744 (N_14744,N_13381,N_13306);
or U14745 (N_14745,N_13397,N_13421);
xor U14746 (N_14746,N_13359,N_13449);
or U14747 (N_14747,N_13564,N_13459);
or U14748 (N_14748,N_13433,N_13638);
or U14749 (N_14749,N_13965,N_13807);
or U14750 (N_14750,N_13538,N_13139);
and U14751 (N_14751,N_13389,N_13813);
xor U14752 (N_14752,N_13547,N_13298);
or U14753 (N_14753,N_13420,N_13033);
xor U14754 (N_14754,N_13815,N_13753);
and U14755 (N_14755,N_13571,N_13903);
xor U14756 (N_14756,N_13289,N_13389);
or U14757 (N_14757,N_13466,N_13164);
nand U14758 (N_14758,N_13005,N_13202);
and U14759 (N_14759,N_13407,N_13260);
xor U14760 (N_14760,N_13647,N_13749);
or U14761 (N_14761,N_13271,N_13365);
nor U14762 (N_14762,N_13584,N_13512);
nand U14763 (N_14763,N_13850,N_13885);
nand U14764 (N_14764,N_13923,N_13888);
or U14765 (N_14765,N_13038,N_13194);
nor U14766 (N_14766,N_13364,N_13843);
nor U14767 (N_14767,N_13314,N_13436);
nand U14768 (N_14768,N_13557,N_13121);
nand U14769 (N_14769,N_13393,N_13436);
or U14770 (N_14770,N_13178,N_13708);
nor U14771 (N_14771,N_13547,N_13879);
xnor U14772 (N_14772,N_13993,N_13307);
nand U14773 (N_14773,N_13921,N_13641);
and U14774 (N_14774,N_13580,N_13256);
nor U14775 (N_14775,N_13315,N_13454);
and U14776 (N_14776,N_13766,N_13997);
and U14777 (N_14777,N_13253,N_13554);
nor U14778 (N_14778,N_13342,N_13751);
or U14779 (N_14779,N_13402,N_13676);
or U14780 (N_14780,N_13982,N_13856);
nor U14781 (N_14781,N_13493,N_13281);
nand U14782 (N_14782,N_13974,N_13791);
xnor U14783 (N_14783,N_13500,N_13960);
or U14784 (N_14784,N_13605,N_13181);
xor U14785 (N_14785,N_13420,N_13761);
or U14786 (N_14786,N_13541,N_13958);
nand U14787 (N_14787,N_13881,N_13389);
or U14788 (N_14788,N_13420,N_13069);
nor U14789 (N_14789,N_13245,N_13818);
nand U14790 (N_14790,N_13551,N_13247);
and U14791 (N_14791,N_13160,N_13599);
or U14792 (N_14792,N_13901,N_13376);
and U14793 (N_14793,N_13950,N_13811);
or U14794 (N_14794,N_13094,N_13516);
nor U14795 (N_14795,N_13516,N_13730);
or U14796 (N_14796,N_13721,N_13562);
and U14797 (N_14797,N_13196,N_13134);
xor U14798 (N_14798,N_13266,N_13132);
and U14799 (N_14799,N_13595,N_13235);
nor U14800 (N_14800,N_13667,N_13809);
nand U14801 (N_14801,N_13705,N_13381);
nand U14802 (N_14802,N_13916,N_13461);
or U14803 (N_14803,N_13424,N_13873);
nand U14804 (N_14804,N_13203,N_13592);
and U14805 (N_14805,N_13426,N_13510);
nand U14806 (N_14806,N_13084,N_13972);
nand U14807 (N_14807,N_13530,N_13927);
and U14808 (N_14808,N_13828,N_13838);
nand U14809 (N_14809,N_13831,N_13754);
or U14810 (N_14810,N_13074,N_13433);
xor U14811 (N_14811,N_13456,N_13022);
or U14812 (N_14812,N_13634,N_13455);
nand U14813 (N_14813,N_13144,N_13109);
xor U14814 (N_14814,N_13833,N_13298);
xnor U14815 (N_14815,N_13819,N_13292);
or U14816 (N_14816,N_13227,N_13170);
xnor U14817 (N_14817,N_13263,N_13932);
xnor U14818 (N_14818,N_13171,N_13033);
nor U14819 (N_14819,N_13897,N_13810);
and U14820 (N_14820,N_13009,N_13159);
and U14821 (N_14821,N_13094,N_13739);
nand U14822 (N_14822,N_13960,N_13951);
and U14823 (N_14823,N_13866,N_13265);
nand U14824 (N_14824,N_13666,N_13396);
and U14825 (N_14825,N_13020,N_13503);
nand U14826 (N_14826,N_13288,N_13737);
nor U14827 (N_14827,N_13767,N_13429);
and U14828 (N_14828,N_13242,N_13994);
nand U14829 (N_14829,N_13657,N_13596);
and U14830 (N_14830,N_13934,N_13201);
nor U14831 (N_14831,N_13294,N_13962);
or U14832 (N_14832,N_13138,N_13822);
nor U14833 (N_14833,N_13563,N_13019);
xnor U14834 (N_14834,N_13122,N_13085);
nand U14835 (N_14835,N_13782,N_13166);
xor U14836 (N_14836,N_13519,N_13392);
xnor U14837 (N_14837,N_13381,N_13966);
and U14838 (N_14838,N_13935,N_13856);
and U14839 (N_14839,N_13254,N_13350);
and U14840 (N_14840,N_13059,N_13485);
nor U14841 (N_14841,N_13484,N_13029);
and U14842 (N_14842,N_13232,N_13526);
nor U14843 (N_14843,N_13970,N_13796);
xor U14844 (N_14844,N_13699,N_13125);
or U14845 (N_14845,N_13940,N_13018);
nand U14846 (N_14846,N_13282,N_13368);
or U14847 (N_14847,N_13236,N_13731);
xor U14848 (N_14848,N_13821,N_13664);
xor U14849 (N_14849,N_13313,N_13080);
xor U14850 (N_14850,N_13246,N_13312);
nand U14851 (N_14851,N_13272,N_13690);
nor U14852 (N_14852,N_13443,N_13387);
nand U14853 (N_14853,N_13860,N_13830);
nand U14854 (N_14854,N_13190,N_13385);
or U14855 (N_14855,N_13445,N_13294);
or U14856 (N_14856,N_13258,N_13648);
xor U14857 (N_14857,N_13707,N_13926);
and U14858 (N_14858,N_13019,N_13055);
xor U14859 (N_14859,N_13343,N_13352);
nor U14860 (N_14860,N_13920,N_13910);
nor U14861 (N_14861,N_13142,N_13218);
nand U14862 (N_14862,N_13382,N_13642);
nand U14863 (N_14863,N_13682,N_13799);
xnor U14864 (N_14864,N_13808,N_13849);
nor U14865 (N_14865,N_13015,N_13782);
and U14866 (N_14866,N_13832,N_13330);
and U14867 (N_14867,N_13629,N_13696);
or U14868 (N_14868,N_13683,N_13532);
xor U14869 (N_14869,N_13516,N_13010);
nor U14870 (N_14870,N_13455,N_13414);
and U14871 (N_14871,N_13819,N_13144);
or U14872 (N_14872,N_13455,N_13364);
and U14873 (N_14873,N_13132,N_13768);
and U14874 (N_14874,N_13285,N_13581);
nand U14875 (N_14875,N_13911,N_13282);
nand U14876 (N_14876,N_13600,N_13831);
nor U14877 (N_14877,N_13820,N_13241);
or U14878 (N_14878,N_13444,N_13044);
or U14879 (N_14879,N_13688,N_13140);
nor U14880 (N_14880,N_13399,N_13782);
and U14881 (N_14881,N_13549,N_13701);
xor U14882 (N_14882,N_13056,N_13257);
or U14883 (N_14883,N_13936,N_13969);
xnor U14884 (N_14884,N_13930,N_13760);
nand U14885 (N_14885,N_13970,N_13551);
nor U14886 (N_14886,N_13240,N_13741);
and U14887 (N_14887,N_13675,N_13528);
nand U14888 (N_14888,N_13727,N_13782);
nand U14889 (N_14889,N_13596,N_13834);
nor U14890 (N_14890,N_13538,N_13916);
xor U14891 (N_14891,N_13769,N_13679);
or U14892 (N_14892,N_13025,N_13813);
nor U14893 (N_14893,N_13679,N_13068);
nand U14894 (N_14894,N_13102,N_13764);
or U14895 (N_14895,N_13671,N_13808);
nor U14896 (N_14896,N_13045,N_13753);
xor U14897 (N_14897,N_13885,N_13220);
or U14898 (N_14898,N_13047,N_13579);
and U14899 (N_14899,N_13872,N_13325);
or U14900 (N_14900,N_13922,N_13282);
nor U14901 (N_14901,N_13929,N_13561);
nand U14902 (N_14902,N_13204,N_13614);
xor U14903 (N_14903,N_13731,N_13286);
nor U14904 (N_14904,N_13653,N_13732);
nor U14905 (N_14905,N_13735,N_13138);
nand U14906 (N_14906,N_13187,N_13220);
xor U14907 (N_14907,N_13259,N_13962);
or U14908 (N_14908,N_13444,N_13901);
or U14909 (N_14909,N_13119,N_13505);
or U14910 (N_14910,N_13846,N_13407);
nand U14911 (N_14911,N_13245,N_13597);
or U14912 (N_14912,N_13966,N_13076);
or U14913 (N_14913,N_13013,N_13025);
nor U14914 (N_14914,N_13543,N_13748);
nor U14915 (N_14915,N_13270,N_13874);
nor U14916 (N_14916,N_13785,N_13701);
nor U14917 (N_14917,N_13266,N_13931);
nor U14918 (N_14918,N_13408,N_13132);
xnor U14919 (N_14919,N_13206,N_13597);
or U14920 (N_14920,N_13461,N_13157);
nand U14921 (N_14921,N_13333,N_13332);
and U14922 (N_14922,N_13246,N_13761);
nor U14923 (N_14923,N_13361,N_13575);
or U14924 (N_14924,N_13437,N_13858);
nand U14925 (N_14925,N_13697,N_13498);
and U14926 (N_14926,N_13597,N_13786);
and U14927 (N_14927,N_13744,N_13715);
nor U14928 (N_14928,N_13520,N_13818);
or U14929 (N_14929,N_13055,N_13605);
nand U14930 (N_14930,N_13268,N_13871);
nand U14931 (N_14931,N_13792,N_13030);
and U14932 (N_14932,N_13866,N_13606);
nor U14933 (N_14933,N_13940,N_13737);
and U14934 (N_14934,N_13689,N_13989);
or U14935 (N_14935,N_13462,N_13484);
and U14936 (N_14936,N_13952,N_13466);
xor U14937 (N_14937,N_13810,N_13398);
xor U14938 (N_14938,N_13199,N_13882);
nand U14939 (N_14939,N_13760,N_13694);
nor U14940 (N_14940,N_13202,N_13599);
and U14941 (N_14941,N_13890,N_13655);
nor U14942 (N_14942,N_13662,N_13520);
or U14943 (N_14943,N_13460,N_13222);
and U14944 (N_14944,N_13930,N_13372);
xor U14945 (N_14945,N_13677,N_13955);
or U14946 (N_14946,N_13569,N_13275);
or U14947 (N_14947,N_13847,N_13221);
nand U14948 (N_14948,N_13878,N_13097);
nand U14949 (N_14949,N_13685,N_13149);
nor U14950 (N_14950,N_13867,N_13784);
nand U14951 (N_14951,N_13165,N_13573);
or U14952 (N_14952,N_13536,N_13523);
nor U14953 (N_14953,N_13069,N_13158);
nor U14954 (N_14954,N_13404,N_13410);
or U14955 (N_14955,N_13539,N_13007);
nand U14956 (N_14956,N_13125,N_13880);
nand U14957 (N_14957,N_13384,N_13581);
and U14958 (N_14958,N_13201,N_13326);
nor U14959 (N_14959,N_13334,N_13950);
nor U14960 (N_14960,N_13346,N_13556);
xor U14961 (N_14961,N_13572,N_13190);
nand U14962 (N_14962,N_13044,N_13767);
nand U14963 (N_14963,N_13717,N_13198);
nand U14964 (N_14964,N_13663,N_13017);
and U14965 (N_14965,N_13433,N_13240);
nor U14966 (N_14966,N_13294,N_13342);
and U14967 (N_14967,N_13671,N_13529);
nand U14968 (N_14968,N_13254,N_13622);
xnor U14969 (N_14969,N_13004,N_13358);
nand U14970 (N_14970,N_13453,N_13263);
nand U14971 (N_14971,N_13810,N_13176);
nand U14972 (N_14972,N_13685,N_13852);
or U14973 (N_14973,N_13200,N_13477);
nor U14974 (N_14974,N_13455,N_13058);
or U14975 (N_14975,N_13288,N_13153);
nor U14976 (N_14976,N_13638,N_13233);
or U14977 (N_14977,N_13374,N_13938);
or U14978 (N_14978,N_13186,N_13107);
xor U14979 (N_14979,N_13934,N_13229);
xor U14980 (N_14980,N_13713,N_13914);
nand U14981 (N_14981,N_13192,N_13737);
nand U14982 (N_14982,N_13063,N_13056);
nor U14983 (N_14983,N_13824,N_13820);
xnor U14984 (N_14984,N_13377,N_13856);
nand U14985 (N_14985,N_13947,N_13532);
nand U14986 (N_14986,N_13731,N_13542);
nor U14987 (N_14987,N_13313,N_13342);
and U14988 (N_14988,N_13049,N_13242);
and U14989 (N_14989,N_13402,N_13199);
nor U14990 (N_14990,N_13778,N_13849);
xnor U14991 (N_14991,N_13110,N_13930);
or U14992 (N_14992,N_13310,N_13146);
nand U14993 (N_14993,N_13085,N_13939);
and U14994 (N_14994,N_13258,N_13327);
or U14995 (N_14995,N_13070,N_13291);
nand U14996 (N_14996,N_13335,N_13383);
nand U14997 (N_14997,N_13626,N_13318);
nor U14998 (N_14998,N_13281,N_13138);
nor U14999 (N_14999,N_13077,N_13466);
and U15000 (N_15000,N_14230,N_14298);
or U15001 (N_15001,N_14995,N_14149);
xor U15002 (N_15002,N_14943,N_14426);
or U15003 (N_15003,N_14145,N_14847);
and U15004 (N_15004,N_14515,N_14337);
and U15005 (N_15005,N_14090,N_14841);
xor U15006 (N_15006,N_14002,N_14566);
xnor U15007 (N_15007,N_14915,N_14194);
or U15008 (N_15008,N_14126,N_14445);
nor U15009 (N_15009,N_14049,N_14466);
or U15010 (N_15010,N_14027,N_14758);
nand U15011 (N_15011,N_14356,N_14241);
nand U15012 (N_15012,N_14406,N_14292);
and U15013 (N_15013,N_14155,N_14615);
xnor U15014 (N_15014,N_14717,N_14349);
nand U15015 (N_15015,N_14626,N_14037);
and U15016 (N_15016,N_14346,N_14117);
nand U15017 (N_15017,N_14201,N_14586);
nor U15018 (N_15018,N_14727,N_14297);
xor U15019 (N_15019,N_14517,N_14701);
nand U15020 (N_15020,N_14955,N_14369);
and U15021 (N_15021,N_14964,N_14577);
nand U15022 (N_15022,N_14216,N_14110);
and U15023 (N_15023,N_14776,N_14303);
or U15024 (N_15024,N_14203,N_14066);
xnor U15025 (N_15025,N_14116,N_14190);
or U15026 (N_15026,N_14111,N_14138);
or U15027 (N_15027,N_14900,N_14227);
or U15028 (N_15028,N_14759,N_14869);
and U15029 (N_15029,N_14164,N_14512);
xnor U15030 (N_15030,N_14183,N_14098);
and U15031 (N_15031,N_14153,N_14826);
xnor U15032 (N_15032,N_14679,N_14625);
nand U15033 (N_15033,N_14248,N_14485);
and U15034 (N_15034,N_14197,N_14715);
xor U15035 (N_15035,N_14889,N_14109);
xor U15036 (N_15036,N_14797,N_14747);
nand U15037 (N_15037,N_14206,N_14592);
nand U15038 (N_15038,N_14225,N_14779);
or U15039 (N_15039,N_14607,N_14749);
or U15040 (N_15040,N_14627,N_14556);
or U15041 (N_15041,N_14524,N_14004);
or U15042 (N_15042,N_14214,N_14718);
or U15043 (N_15043,N_14233,N_14383);
and U15044 (N_15044,N_14600,N_14585);
nor U15045 (N_15045,N_14065,N_14804);
xnor U15046 (N_15046,N_14144,N_14091);
xor U15047 (N_15047,N_14856,N_14481);
and U15048 (N_15048,N_14534,N_14911);
nor U15049 (N_15049,N_14008,N_14532);
xor U15050 (N_15050,N_14536,N_14444);
and U15051 (N_15051,N_14809,N_14215);
nand U15052 (N_15052,N_14909,N_14198);
nand U15053 (N_15053,N_14307,N_14500);
nor U15054 (N_15054,N_14119,N_14754);
or U15055 (N_15055,N_14450,N_14275);
or U15056 (N_15056,N_14937,N_14786);
and U15057 (N_15057,N_14016,N_14345);
nor U15058 (N_15058,N_14694,N_14609);
or U15059 (N_15059,N_14533,N_14781);
nand U15060 (N_15060,N_14720,N_14589);
nor U15061 (N_15061,N_14036,N_14716);
xor U15062 (N_15062,N_14866,N_14259);
xnor U15063 (N_15063,N_14744,N_14833);
nor U15064 (N_15064,N_14010,N_14505);
xor U15065 (N_15065,N_14125,N_14906);
xnor U15066 (N_15066,N_14163,N_14315);
or U15067 (N_15067,N_14761,N_14687);
and U15068 (N_15068,N_14122,N_14174);
nand U15069 (N_15069,N_14564,N_14099);
xor U15070 (N_15070,N_14622,N_14608);
nand U15071 (N_15071,N_14658,N_14612);
nand U15072 (N_15072,N_14985,N_14410);
nand U15073 (N_15073,N_14721,N_14428);
and U15074 (N_15074,N_14782,N_14342);
or U15075 (N_15075,N_14790,N_14278);
or U15076 (N_15076,N_14028,N_14492);
nand U15077 (N_15077,N_14921,N_14686);
nand U15078 (N_15078,N_14838,N_14488);
xor U15079 (N_15079,N_14223,N_14039);
nor U15080 (N_15080,N_14907,N_14367);
xnor U15081 (N_15081,N_14530,N_14771);
and U15082 (N_15082,N_14285,N_14070);
and U15083 (N_15083,N_14919,N_14055);
and U15084 (N_15084,N_14571,N_14076);
or U15085 (N_15085,N_14325,N_14266);
or U15086 (N_15086,N_14237,N_14128);
or U15087 (N_15087,N_14504,N_14879);
xor U15088 (N_15088,N_14817,N_14798);
xnor U15089 (N_15089,N_14708,N_14540);
nor U15090 (N_15090,N_14881,N_14335);
or U15091 (N_15091,N_14897,N_14801);
nor U15092 (N_15092,N_14180,N_14252);
nand U15093 (N_15093,N_14478,N_14118);
nor U15094 (N_15094,N_14281,N_14343);
nor U15095 (N_15095,N_14186,N_14825);
nor U15096 (N_15096,N_14330,N_14989);
or U15097 (N_15097,N_14063,N_14350);
and U15098 (N_15098,N_14148,N_14461);
xor U15099 (N_15099,N_14666,N_14685);
xor U15100 (N_15100,N_14613,N_14896);
nand U15101 (N_15101,N_14147,N_14291);
xnor U15102 (N_15102,N_14333,N_14068);
nor U15103 (N_15103,N_14871,N_14332);
or U15104 (N_15104,N_14736,N_14582);
or U15105 (N_15105,N_14965,N_14290);
nand U15106 (N_15106,N_14100,N_14618);
xor U15107 (N_15107,N_14531,N_14047);
xnor U15108 (N_15108,N_14997,N_14501);
or U15109 (N_15109,N_14173,N_14092);
or U15110 (N_15110,N_14944,N_14509);
xnor U15111 (N_15111,N_14046,N_14756);
nand U15112 (N_15112,N_14816,N_14599);
and U15113 (N_15113,N_14860,N_14418);
nor U15114 (N_15114,N_14941,N_14348);
nor U15115 (N_15115,N_14384,N_14684);
nand U15116 (N_15116,N_14220,N_14014);
xnor U15117 (N_15117,N_14210,N_14712);
xnor U15118 (N_15118,N_14802,N_14024);
nand U15119 (N_15119,N_14570,N_14904);
or U15120 (N_15120,N_14677,N_14226);
nor U15121 (N_15121,N_14419,N_14352);
and U15122 (N_15122,N_14537,N_14732);
xnor U15123 (N_15123,N_14260,N_14641);
and U15124 (N_15124,N_14837,N_14886);
nor U15125 (N_15125,N_14412,N_14903);
xnor U15126 (N_15126,N_14025,N_14660);
nand U15127 (N_15127,N_14218,N_14709);
or U15128 (N_15128,N_14925,N_14001);
or U15129 (N_15129,N_14486,N_14420);
or U15130 (N_15130,N_14242,N_14603);
and U15131 (N_15131,N_14982,N_14849);
nand U15132 (N_15132,N_14820,N_14652);
nor U15133 (N_15133,N_14150,N_14397);
xnor U15134 (N_15134,N_14541,N_14288);
nand U15135 (N_15135,N_14045,N_14722);
xnor U15136 (N_15136,N_14396,N_14213);
and U15137 (N_15137,N_14044,N_14967);
nand U15138 (N_15138,N_14587,N_14473);
or U15139 (N_15139,N_14211,N_14018);
and U15140 (N_15140,N_14772,N_14729);
xnor U15141 (N_15141,N_14395,N_14651);
and U15142 (N_15142,N_14441,N_14760);
nor U15143 (N_15143,N_14806,N_14535);
and U15144 (N_15144,N_14678,N_14401);
or U15145 (N_15145,N_14452,N_14740);
nor U15146 (N_15146,N_14638,N_14482);
nand U15147 (N_15147,N_14883,N_14040);
xnor U15148 (N_15148,N_14236,N_14158);
xor U15149 (N_15149,N_14026,N_14200);
nor U15150 (N_15150,N_14699,N_14151);
xor U15151 (N_15151,N_14232,N_14591);
nand U15152 (N_15152,N_14707,N_14393);
and U15153 (N_15153,N_14606,N_14217);
nor U15154 (N_15154,N_14360,N_14526);
xnor U15155 (N_15155,N_14936,N_14750);
or U15156 (N_15156,N_14354,N_14457);
xor U15157 (N_15157,N_14762,N_14280);
xnor U15158 (N_15158,N_14518,N_14133);
nand U15159 (N_15159,N_14484,N_14377);
nand U15160 (N_15160,N_14499,N_14446);
or U15161 (N_15161,N_14489,N_14435);
xor U15162 (N_15162,N_14204,N_14135);
nand U15163 (N_15163,N_14690,N_14495);
xnor U15164 (N_15164,N_14752,N_14703);
and U15165 (N_15165,N_14874,N_14075);
nand U15166 (N_15166,N_14506,N_14081);
xor U15167 (N_15167,N_14391,N_14934);
and U15168 (N_15168,N_14256,N_14705);
or U15169 (N_15169,N_14726,N_14598);
nand U15170 (N_15170,N_14812,N_14120);
nor U15171 (N_15171,N_14831,N_14558);
nor U15172 (N_15172,N_14981,N_14277);
and U15173 (N_15173,N_14191,N_14430);
or U15174 (N_15174,N_14807,N_14742);
or U15175 (N_15175,N_14822,N_14873);
nand U15176 (N_15176,N_14913,N_14364);
or U15177 (N_15177,N_14379,N_14328);
or U15178 (N_15178,N_14132,N_14828);
nand U15179 (N_15179,N_14502,N_14319);
or U15180 (N_15180,N_14424,N_14623);
nand U15181 (N_15181,N_14697,N_14258);
xor U15182 (N_15182,N_14926,N_14311);
xor U15183 (N_15183,N_14818,N_14422);
nand U15184 (N_15184,N_14057,N_14184);
or U15185 (N_15185,N_14273,N_14574);
nand U15186 (N_15186,N_14855,N_14601);
nand U15187 (N_15187,N_14443,N_14082);
and U15188 (N_15188,N_14240,N_14719);
and U15189 (N_15189,N_14178,N_14308);
xnor U15190 (N_15190,N_14770,N_14956);
nor U15191 (N_15191,N_14262,N_14875);
xor U15192 (N_15192,N_14610,N_14235);
or U15193 (N_15193,N_14508,N_14867);
nor U15194 (N_15194,N_14939,N_14511);
xnor U15195 (N_15195,N_14372,N_14813);
xnor U15196 (N_15196,N_14324,N_14166);
nor U15197 (N_15197,N_14803,N_14853);
nor U15198 (N_15198,N_14267,N_14338);
nor U15199 (N_15199,N_14131,N_14918);
xnor U15200 (N_15200,N_14632,N_14269);
or U15201 (N_15201,N_14968,N_14789);
or U15202 (N_15202,N_14305,N_14105);
xor U15203 (N_15203,N_14403,N_14734);
or U15204 (N_15204,N_14862,N_14279);
or U15205 (N_15205,N_14013,N_14972);
and U15206 (N_15206,N_14991,N_14318);
nand U15207 (N_15207,N_14629,N_14954);
and U15208 (N_15208,N_14246,N_14894);
or U15209 (N_15209,N_14108,N_14695);
xor U15210 (N_15210,N_14030,N_14407);
or U15211 (N_15211,N_14331,N_14633);
nor U15212 (N_15212,N_14041,N_14783);
nor U15213 (N_15213,N_14035,N_14080);
and U15214 (N_15214,N_14669,N_14614);
and U15215 (N_15215,N_14336,N_14547);
or U15216 (N_15216,N_14265,N_14253);
and U15217 (N_15217,N_14159,N_14673);
nand U15218 (N_15218,N_14073,N_14192);
nand U15219 (N_15219,N_14661,N_14086);
xnor U15220 (N_15220,N_14576,N_14519);
xnor U15221 (N_15221,N_14078,N_14800);
nand U15222 (N_15222,N_14827,N_14850);
and U15223 (N_15223,N_14560,N_14142);
nor U15224 (N_15224,N_14094,N_14584);
nor U15225 (N_15225,N_14101,N_14573);
nand U15226 (N_15226,N_14739,N_14844);
nor U15227 (N_15227,N_14983,N_14980);
or U15228 (N_15228,N_14552,N_14548);
nor U15229 (N_15229,N_14129,N_14572);
nor U15230 (N_15230,N_14808,N_14411);
and U15231 (N_15231,N_14193,N_14923);
xnor U15232 (N_15232,N_14402,N_14984);
or U15233 (N_15233,N_14616,N_14583);
or U15234 (N_15234,N_14433,N_14229);
or U15235 (N_15235,N_14079,N_14042);
or U15236 (N_15236,N_14969,N_14427);
and U15237 (N_15237,N_14971,N_14152);
or U15238 (N_15238,N_14554,N_14205);
nor U15239 (N_15239,N_14239,N_14301);
nand U15240 (N_15240,N_14743,N_14636);
or U15241 (N_15241,N_14528,N_14999);
or U15242 (N_15242,N_14745,N_14104);
and U15243 (N_15243,N_14725,N_14463);
nor U15244 (N_15244,N_14413,N_14876);
nand U15245 (N_15245,N_14780,N_14891);
and U15246 (N_15246,N_14966,N_14208);
and U15247 (N_15247,N_14946,N_14851);
or U15248 (N_15248,N_14032,N_14674);
nand U15249 (N_15249,N_14711,N_14713);
xnor U15250 (N_15250,N_14767,N_14656);
or U15251 (N_15251,N_14832,N_14340);
or U15252 (N_15252,N_14575,N_14029);
xnor U15253 (N_15253,N_14649,N_14320);
and U15254 (N_15254,N_14839,N_14255);
nand U15255 (N_15255,N_14257,N_14243);
and U15256 (N_15256,N_14753,N_14670);
nand U15257 (N_15257,N_14814,N_14887);
nor U15258 (N_15258,N_14637,N_14738);
nand U15259 (N_15259,N_14438,N_14475);
nor U15260 (N_15260,N_14858,N_14640);
and U15261 (N_15261,N_14154,N_14527);
nand U15262 (N_15262,N_14312,N_14347);
nand U15263 (N_15263,N_14978,N_14012);
nor U15264 (N_15264,N_14642,N_14176);
nand U15265 (N_15265,N_14351,N_14702);
or U15266 (N_15266,N_14514,N_14022);
xor U15267 (N_15267,N_14112,N_14525);
or U15268 (N_15268,N_14134,N_14497);
and U15269 (N_15269,N_14456,N_14949);
nor U15270 (N_15270,N_14408,N_14052);
or U15271 (N_15271,N_14810,N_14177);
nand U15272 (N_15272,N_14620,N_14960);
and U15273 (N_15273,N_14878,N_14924);
nor U15274 (N_15274,N_14365,N_14787);
or U15275 (N_15275,N_14970,N_14893);
and U15276 (N_15276,N_14380,N_14121);
xor U15277 (N_15277,N_14023,N_14160);
xor U15278 (N_15278,N_14635,N_14852);
xnor U15279 (N_15279,N_14439,N_14619);
and U15280 (N_15280,N_14181,N_14339);
and U15281 (N_15281,N_14731,N_14487);
or U15282 (N_15282,N_14510,N_14961);
nor U15283 (N_15283,N_14162,N_14821);
or U15284 (N_15284,N_14795,N_14902);
or U15285 (N_15285,N_14421,N_14938);
nor U15286 (N_15286,N_14387,N_14043);
nor U15287 (N_15287,N_14910,N_14058);
and U15288 (N_15288,N_14363,N_14429);
or U15289 (N_15289,N_14423,N_14631);
nand U15290 (N_15290,N_14139,N_14017);
or U15291 (N_15291,N_14053,N_14920);
xnor U15292 (N_15292,N_14644,N_14565);
nand U15293 (N_15293,N_14778,N_14491);
xor U15294 (N_15294,N_14317,N_14544);
xnor U15295 (N_15295,N_14003,N_14060);
xnor U15296 (N_15296,N_14048,N_14170);
nand U15297 (N_15297,N_14683,N_14639);
and U15298 (N_15298,N_14169,N_14579);
or U15299 (N_15299,N_14388,N_14792);
nor U15300 (N_15300,N_14621,N_14474);
nand U15301 (N_15301,N_14447,N_14442);
xnor U15302 (N_15302,N_14766,N_14299);
or U15303 (N_15303,N_14358,N_14681);
or U15304 (N_15304,N_14179,N_14663);
nor U15305 (N_15305,N_14249,N_14137);
and U15306 (N_15306,N_14261,N_14769);
nor U15307 (N_15307,N_14882,N_14355);
and U15308 (N_15308,N_14819,N_14643);
or U15309 (N_15309,N_14436,N_14187);
nor U15310 (N_15310,N_14464,N_14189);
and U15311 (N_15311,N_14823,N_14951);
or U15312 (N_15312,N_14945,N_14378);
nand U15313 (N_15313,N_14359,N_14529);
or U15314 (N_15314,N_14286,N_14908);
nor U15315 (N_15315,N_14634,N_14448);
xnor U15316 (N_15316,N_14254,N_14932);
nor U15317 (N_15317,N_14006,N_14723);
and U15318 (N_15318,N_14597,N_14561);
and U15319 (N_15319,N_14682,N_14513);
nor U15320 (N_15320,N_14977,N_14796);
nand U15321 (N_15321,N_14453,N_14196);
xor U15322 (N_15322,N_14161,N_14064);
xor U15323 (N_15323,N_14293,N_14399);
xor U15324 (N_15324,N_14788,N_14313);
and U15325 (N_15325,N_14588,N_14095);
nor U15326 (N_15326,N_14768,N_14664);
and U15327 (N_15327,N_14829,N_14757);
nand U15328 (N_15328,N_14763,N_14973);
and U15329 (N_15329,N_14947,N_14115);
nor U15330 (N_15330,N_14884,N_14628);
nor U15331 (N_15331,N_14523,N_14268);
xor U15332 (N_15332,N_14988,N_14195);
xnor U15333 (N_15333,N_14563,N_14569);
and U15334 (N_15334,N_14594,N_14454);
nor U15335 (N_15335,N_14156,N_14276);
nand U15336 (N_15336,N_14596,N_14329);
nand U15337 (N_15337,N_14546,N_14551);
nand U15338 (N_15338,N_14764,N_14019);
or U15339 (N_15339,N_14021,N_14958);
nor U15340 (N_15340,N_14244,N_14437);
xnor U15341 (N_15341,N_14264,N_14050);
nor U15342 (N_15342,N_14199,N_14692);
xnor U15343 (N_15343,N_14704,N_14948);
and U15344 (N_15344,N_14927,N_14219);
nand U15345 (N_15345,N_14034,N_14791);
or U15346 (N_15346,N_14326,N_14357);
or U15347 (N_15347,N_14710,N_14993);
and U15348 (N_15348,N_14794,N_14458);
nand U15349 (N_15349,N_14931,N_14899);
and U15350 (N_15350,N_14316,N_14735);
xnor U15351 (N_15351,N_14289,N_14167);
xnor U15352 (N_15352,N_14842,N_14088);
nor U15353 (N_15353,N_14835,N_14657);
xor U15354 (N_15354,N_14294,N_14659);
nor U15355 (N_15355,N_14415,N_14785);
or U15356 (N_15356,N_14274,N_14493);
and U15357 (N_15357,N_14471,N_14974);
and U15358 (N_15358,N_14870,N_14748);
and U15359 (N_15359,N_14698,N_14270);
nand U15360 (N_15360,N_14959,N_14469);
nand U15361 (N_15361,N_14476,N_14127);
nor U15362 (N_15362,N_14568,N_14093);
nor U15363 (N_15363,N_14550,N_14238);
nor U15364 (N_15364,N_14590,N_14084);
nand U15365 (N_15365,N_14845,N_14917);
nor U15366 (N_15366,N_14113,N_14662);
and U15367 (N_15367,N_14775,N_14602);
and U15368 (N_15368,N_14398,N_14087);
nor U15369 (N_15369,N_14414,N_14287);
or U15370 (N_15370,N_14467,N_14263);
nor U15371 (N_15371,N_14400,N_14353);
nand U15372 (N_15372,N_14344,N_14930);
nand U15373 (N_15373,N_14733,N_14462);
or U15374 (N_15374,N_14171,N_14503);
or U15375 (N_15375,N_14103,N_14470);
nor U15376 (N_15376,N_14667,N_14507);
nor U15377 (N_15377,N_14067,N_14054);
nand U15378 (N_15378,N_14432,N_14859);
nor U15379 (N_15379,N_14124,N_14872);
nor U15380 (N_15380,N_14304,N_14188);
xor U15381 (N_15381,N_14207,N_14604);
xnor U15382 (N_15382,N_14382,N_14668);
or U15383 (N_15383,N_14953,N_14477);
and U15384 (N_15384,N_14371,N_14892);
or U15385 (N_15385,N_14895,N_14490);
nand U15386 (N_15386,N_14077,N_14957);
or U15387 (N_15387,N_14251,N_14221);
xnor U15388 (N_15388,N_14730,N_14848);
or U15389 (N_15389,N_14898,N_14373);
nand U15390 (N_15390,N_14815,N_14861);
xor U15391 (N_15391,N_14309,N_14394);
nand U15392 (N_15392,N_14865,N_14114);
nor U15393 (N_15393,N_14843,N_14392);
nand U15394 (N_15394,N_14942,N_14366);
nor U15395 (N_15395,N_14940,N_14630);
or U15396 (N_15396,N_14645,N_14283);
nor U15397 (N_15397,N_14617,N_14976);
and U15398 (N_15398,N_14557,N_14250);
nand U15399 (N_15399,N_14480,N_14009);
or U15400 (N_15400,N_14846,N_14987);
nor U15401 (N_15401,N_14496,N_14321);
nor U15402 (N_15402,N_14714,N_14693);
nand U15403 (N_15403,N_14905,N_14996);
nor U15404 (N_15404,N_14986,N_14741);
nor U15405 (N_15405,N_14033,N_14375);
nor U15406 (N_15406,N_14655,N_14784);
nand U15407 (N_15407,N_14130,N_14696);
and U15408 (N_15408,N_14417,N_14578);
xnor U15409 (N_15409,N_14062,N_14834);
xor U15410 (N_15410,N_14059,N_14755);
nand U15411 (N_15411,N_14654,N_14774);
nand U15412 (N_15412,N_14777,N_14868);
or U15413 (N_15413,N_14950,N_14224);
nor U15414 (N_15414,N_14830,N_14885);
nand U15415 (N_15415,N_14011,N_14793);
xnor U15416 (N_15416,N_14314,N_14020);
or U15417 (N_15417,N_14172,N_14168);
nand U15418 (N_15418,N_14521,N_14724);
and U15419 (N_15419,N_14000,N_14864);
and U15420 (N_15420,N_14549,N_14370);
nand U15421 (N_15421,N_14580,N_14520);
or U15422 (N_15422,N_14451,N_14545);
nor U15423 (N_15423,N_14157,N_14465);
nand U15424 (N_15424,N_14146,N_14007);
xor U15425 (N_15425,N_14680,N_14840);
and U15426 (N_15426,N_14097,N_14689);
xnor U15427 (N_15427,N_14031,N_14479);
and U15428 (N_15428,N_14998,N_14306);
and U15429 (N_15429,N_14543,N_14675);
xnor U15430 (N_15430,N_14555,N_14890);
nand U15431 (N_15431,N_14854,N_14691);
xor U15432 (N_15432,N_14282,N_14051);
and U15433 (N_15433,N_14605,N_14405);
nor U15434 (N_15434,N_14061,N_14038);
nand U15435 (N_15435,N_14888,N_14005);
or U15436 (N_15436,N_14389,N_14368);
nor U15437 (N_15437,N_14361,N_14624);
xor U15438 (N_15438,N_14863,N_14914);
and U15439 (N_15439,N_14322,N_14449);
and U15440 (N_15440,N_14671,N_14234);
or U15441 (N_15441,N_14522,N_14746);
nor U15442 (N_15442,N_14647,N_14302);
or U15443 (N_15443,N_14665,N_14362);
or U15444 (N_15444,N_14074,N_14212);
nor U15445 (N_15445,N_14425,N_14737);
nor U15446 (N_15446,N_14979,N_14468);
xnor U15447 (N_15447,N_14434,N_14089);
nor U15448 (N_15448,N_14992,N_14390);
nor U15449 (N_15449,N_14209,N_14805);
and U15450 (N_15450,N_14271,N_14494);
nor U15451 (N_15451,N_14611,N_14676);
or U15452 (N_15452,N_14107,N_14341);
or U15453 (N_15453,N_14334,N_14928);
xor U15454 (N_15454,N_14646,N_14516);
nand U15455 (N_15455,N_14409,N_14952);
or U15456 (N_15456,N_14083,N_14182);
xor U15457 (N_15457,N_14799,N_14653);
and U15458 (N_15458,N_14202,N_14085);
nor U15459 (N_15459,N_14143,N_14165);
and U15460 (N_15460,N_14175,N_14539);
and U15461 (N_15461,N_14728,N_14562);
xnor U15462 (N_15462,N_14272,N_14381);
and U15463 (N_15463,N_14935,N_14141);
and U15464 (N_15464,N_14404,N_14385);
and U15465 (N_15465,N_14374,N_14300);
nor U15466 (N_15466,N_14096,N_14975);
nand U15467 (N_15467,N_14990,N_14072);
nand U15468 (N_15468,N_14567,N_14542);
and U15469 (N_15469,N_14559,N_14228);
nor U15470 (N_15470,N_14553,N_14460);
nor U15471 (N_15471,N_14310,N_14963);
or U15472 (N_15472,N_14912,N_14140);
or U15473 (N_15473,N_14231,N_14773);
nand U15474 (N_15474,N_14877,N_14498);
nand U15475 (N_15475,N_14376,N_14581);
nand U15476 (N_15476,N_14901,N_14386);
xor U15477 (N_15477,N_14811,N_14069);
nand U15478 (N_15478,N_14593,N_14071);
nor U15479 (N_15479,N_14765,N_14650);
nand U15480 (N_15480,N_14751,N_14472);
nand U15481 (N_15481,N_14136,N_14962);
or U15482 (N_15482,N_14222,N_14296);
xnor U15483 (N_15483,N_14483,N_14295);
nor U15484 (N_15484,N_14648,N_14459);
or U15485 (N_15485,N_14857,N_14327);
and U15486 (N_15486,N_14672,N_14916);
or U15487 (N_15487,N_14824,N_14836);
nand U15488 (N_15488,N_14455,N_14323);
xor U15489 (N_15489,N_14123,N_14015);
or U15490 (N_15490,N_14922,N_14245);
nor U15491 (N_15491,N_14102,N_14994);
nor U15492 (N_15492,N_14929,N_14416);
nand U15493 (N_15493,N_14538,N_14595);
and U15494 (N_15494,N_14700,N_14688);
nand U15495 (N_15495,N_14706,N_14185);
nand U15496 (N_15496,N_14880,N_14933);
nor U15497 (N_15497,N_14106,N_14056);
or U15498 (N_15498,N_14431,N_14440);
xnor U15499 (N_15499,N_14284,N_14247);
xnor U15500 (N_15500,N_14280,N_14525);
xor U15501 (N_15501,N_14967,N_14162);
nand U15502 (N_15502,N_14248,N_14311);
nor U15503 (N_15503,N_14375,N_14691);
xor U15504 (N_15504,N_14482,N_14561);
nand U15505 (N_15505,N_14914,N_14844);
nor U15506 (N_15506,N_14420,N_14335);
nand U15507 (N_15507,N_14719,N_14002);
nor U15508 (N_15508,N_14438,N_14726);
nand U15509 (N_15509,N_14894,N_14032);
or U15510 (N_15510,N_14112,N_14211);
nor U15511 (N_15511,N_14273,N_14719);
nor U15512 (N_15512,N_14642,N_14033);
nor U15513 (N_15513,N_14521,N_14456);
or U15514 (N_15514,N_14483,N_14558);
nor U15515 (N_15515,N_14856,N_14313);
and U15516 (N_15516,N_14173,N_14788);
nand U15517 (N_15517,N_14139,N_14843);
xnor U15518 (N_15518,N_14534,N_14677);
and U15519 (N_15519,N_14431,N_14581);
nor U15520 (N_15520,N_14070,N_14929);
nand U15521 (N_15521,N_14600,N_14930);
nor U15522 (N_15522,N_14258,N_14229);
nor U15523 (N_15523,N_14730,N_14693);
xnor U15524 (N_15524,N_14495,N_14460);
nand U15525 (N_15525,N_14431,N_14293);
and U15526 (N_15526,N_14431,N_14359);
and U15527 (N_15527,N_14041,N_14181);
or U15528 (N_15528,N_14691,N_14915);
nand U15529 (N_15529,N_14486,N_14543);
nand U15530 (N_15530,N_14491,N_14842);
or U15531 (N_15531,N_14992,N_14384);
or U15532 (N_15532,N_14009,N_14163);
nor U15533 (N_15533,N_14632,N_14383);
nand U15534 (N_15534,N_14242,N_14412);
nor U15535 (N_15535,N_14788,N_14011);
or U15536 (N_15536,N_14064,N_14206);
and U15537 (N_15537,N_14289,N_14072);
or U15538 (N_15538,N_14100,N_14884);
xnor U15539 (N_15539,N_14547,N_14799);
and U15540 (N_15540,N_14937,N_14774);
or U15541 (N_15541,N_14185,N_14427);
nor U15542 (N_15542,N_14247,N_14392);
and U15543 (N_15543,N_14665,N_14877);
nor U15544 (N_15544,N_14708,N_14616);
xor U15545 (N_15545,N_14095,N_14822);
and U15546 (N_15546,N_14154,N_14843);
xnor U15547 (N_15547,N_14789,N_14943);
nor U15548 (N_15548,N_14495,N_14776);
and U15549 (N_15549,N_14391,N_14671);
nor U15550 (N_15550,N_14591,N_14358);
and U15551 (N_15551,N_14728,N_14471);
and U15552 (N_15552,N_14012,N_14256);
or U15553 (N_15553,N_14017,N_14162);
or U15554 (N_15554,N_14641,N_14493);
nor U15555 (N_15555,N_14664,N_14785);
nor U15556 (N_15556,N_14027,N_14473);
nand U15557 (N_15557,N_14835,N_14096);
xor U15558 (N_15558,N_14763,N_14569);
and U15559 (N_15559,N_14171,N_14706);
or U15560 (N_15560,N_14983,N_14578);
or U15561 (N_15561,N_14527,N_14568);
nand U15562 (N_15562,N_14411,N_14092);
xor U15563 (N_15563,N_14795,N_14886);
xor U15564 (N_15564,N_14901,N_14898);
nor U15565 (N_15565,N_14846,N_14870);
nand U15566 (N_15566,N_14992,N_14449);
xnor U15567 (N_15567,N_14452,N_14682);
and U15568 (N_15568,N_14943,N_14377);
xor U15569 (N_15569,N_14565,N_14822);
xor U15570 (N_15570,N_14921,N_14320);
or U15571 (N_15571,N_14830,N_14873);
nor U15572 (N_15572,N_14935,N_14801);
nand U15573 (N_15573,N_14526,N_14341);
xnor U15574 (N_15574,N_14296,N_14154);
and U15575 (N_15575,N_14328,N_14684);
nand U15576 (N_15576,N_14640,N_14501);
nand U15577 (N_15577,N_14693,N_14868);
xor U15578 (N_15578,N_14923,N_14294);
nand U15579 (N_15579,N_14217,N_14960);
nand U15580 (N_15580,N_14497,N_14830);
nand U15581 (N_15581,N_14723,N_14848);
and U15582 (N_15582,N_14174,N_14757);
and U15583 (N_15583,N_14632,N_14567);
nand U15584 (N_15584,N_14199,N_14004);
and U15585 (N_15585,N_14152,N_14104);
and U15586 (N_15586,N_14447,N_14071);
nand U15587 (N_15587,N_14769,N_14994);
nor U15588 (N_15588,N_14199,N_14297);
xnor U15589 (N_15589,N_14822,N_14257);
or U15590 (N_15590,N_14032,N_14576);
and U15591 (N_15591,N_14966,N_14280);
or U15592 (N_15592,N_14154,N_14545);
and U15593 (N_15593,N_14291,N_14000);
nor U15594 (N_15594,N_14885,N_14921);
and U15595 (N_15595,N_14748,N_14067);
nor U15596 (N_15596,N_14287,N_14225);
xnor U15597 (N_15597,N_14684,N_14453);
or U15598 (N_15598,N_14519,N_14302);
and U15599 (N_15599,N_14937,N_14028);
or U15600 (N_15600,N_14953,N_14907);
and U15601 (N_15601,N_14862,N_14390);
and U15602 (N_15602,N_14753,N_14776);
xnor U15603 (N_15603,N_14577,N_14646);
and U15604 (N_15604,N_14377,N_14106);
and U15605 (N_15605,N_14321,N_14304);
xnor U15606 (N_15606,N_14851,N_14203);
nand U15607 (N_15607,N_14394,N_14074);
nand U15608 (N_15608,N_14721,N_14418);
nor U15609 (N_15609,N_14393,N_14388);
or U15610 (N_15610,N_14632,N_14909);
or U15611 (N_15611,N_14999,N_14090);
xnor U15612 (N_15612,N_14155,N_14314);
or U15613 (N_15613,N_14209,N_14416);
and U15614 (N_15614,N_14801,N_14429);
xor U15615 (N_15615,N_14386,N_14794);
or U15616 (N_15616,N_14914,N_14258);
xnor U15617 (N_15617,N_14632,N_14601);
nand U15618 (N_15618,N_14996,N_14511);
or U15619 (N_15619,N_14969,N_14589);
nand U15620 (N_15620,N_14396,N_14770);
xor U15621 (N_15621,N_14938,N_14463);
or U15622 (N_15622,N_14915,N_14980);
and U15623 (N_15623,N_14353,N_14957);
nand U15624 (N_15624,N_14022,N_14056);
nand U15625 (N_15625,N_14965,N_14611);
nand U15626 (N_15626,N_14803,N_14587);
or U15627 (N_15627,N_14880,N_14945);
nand U15628 (N_15628,N_14200,N_14195);
nor U15629 (N_15629,N_14947,N_14292);
or U15630 (N_15630,N_14318,N_14634);
nand U15631 (N_15631,N_14554,N_14508);
xnor U15632 (N_15632,N_14243,N_14351);
nand U15633 (N_15633,N_14416,N_14351);
nor U15634 (N_15634,N_14711,N_14663);
and U15635 (N_15635,N_14615,N_14228);
nand U15636 (N_15636,N_14993,N_14450);
or U15637 (N_15637,N_14196,N_14190);
xor U15638 (N_15638,N_14032,N_14151);
xor U15639 (N_15639,N_14605,N_14814);
nor U15640 (N_15640,N_14847,N_14031);
nor U15641 (N_15641,N_14772,N_14018);
and U15642 (N_15642,N_14609,N_14458);
and U15643 (N_15643,N_14908,N_14992);
or U15644 (N_15644,N_14585,N_14283);
nor U15645 (N_15645,N_14487,N_14374);
and U15646 (N_15646,N_14642,N_14676);
nor U15647 (N_15647,N_14557,N_14818);
or U15648 (N_15648,N_14935,N_14328);
nor U15649 (N_15649,N_14632,N_14833);
and U15650 (N_15650,N_14013,N_14171);
or U15651 (N_15651,N_14467,N_14968);
nand U15652 (N_15652,N_14589,N_14800);
nand U15653 (N_15653,N_14073,N_14530);
xnor U15654 (N_15654,N_14005,N_14155);
nor U15655 (N_15655,N_14598,N_14350);
xnor U15656 (N_15656,N_14764,N_14024);
or U15657 (N_15657,N_14182,N_14902);
or U15658 (N_15658,N_14454,N_14152);
nor U15659 (N_15659,N_14835,N_14069);
xnor U15660 (N_15660,N_14149,N_14623);
or U15661 (N_15661,N_14352,N_14748);
and U15662 (N_15662,N_14554,N_14334);
nand U15663 (N_15663,N_14247,N_14964);
nor U15664 (N_15664,N_14484,N_14299);
nor U15665 (N_15665,N_14098,N_14997);
nor U15666 (N_15666,N_14134,N_14084);
nor U15667 (N_15667,N_14940,N_14816);
nand U15668 (N_15668,N_14277,N_14738);
and U15669 (N_15669,N_14275,N_14189);
or U15670 (N_15670,N_14739,N_14994);
xor U15671 (N_15671,N_14392,N_14196);
and U15672 (N_15672,N_14720,N_14577);
nor U15673 (N_15673,N_14419,N_14679);
nor U15674 (N_15674,N_14931,N_14050);
xnor U15675 (N_15675,N_14377,N_14030);
or U15676 (N_15676,N_14951,N_14609);
or U15677 (N_15677,N_14160,N_14251);
and U15678 (N_15678,N_14431,N_14869);
or U15679 (N_15679,N_14967,N_14137);
xnor U15680 (N_15680,N_14231,N_14238);
nor U15681 (N_15681,N_14434,N_14694);
xor U15682 (N_15682,N_14128,N_14271);
xor U15683 (N_15683,N_14110,N_14634);
nand U15684 (N_15684,N_14112,N_14500);
nand U15685 (N_15685,N_14967,N_14663);
nor U15686 (N_15686,N_14512,N_14782);
nand U15687 (N_15687,N_14868,N_14269);
and U15688 (N_15688,N_14222,N_14887);
nor U15689 (N_15689,N_14820,N_14310);
nand U15690 (N_15690,N_14507,N_14052);
nand U15691 (N_15691,N_14584,N_14446);
xor U15692 (N_15692,N_14867,N_14103);
and U15693 (N_15693,N_14615,N_14775);
nor U15694 (N_15694,N_14808,N_14577);
xor U15695 (N_15695,N_14137,N_14817);
or U15696 (N_15696,N_14865,N_14853);
nor U15697 (N_15697,N_14828,N_14091);
nand U15698 (N_15698,N_14965,N_14195);
nor U15699 (N_15699,N_14393,N_14652);
and U15700 (N_15700,N_14187,N_14994);
and U15701 (N_15701,N_14126,N_14076);
nand U15702 (N_15702,N_14511,N_14411);
xor U15703 (N_15703,N_14425,N_14901);
nand U15704 (N_15704,N_14218,N_14486);
nor U15705 (N_15705,N_14303,N_14929);
nor U15706 (N_15706,N_14355,N_14233);
nor U15707 (N_15707,N_14570,N_14117);
and U15708 (N_15708,N_14475,N_14347);
nand U15709 (N_15709,N_14498,N_14555);
and U15710 (N_15710,N_14598,N_14331);
nor U15711 (N_15711,N_14328,N_14030);
or U15712 (N_15712,N_14044,N_14017);
or U15713 (N_15713,N_14899,N_14715);
nor U15714 (N_15714,N_14079,N_14096);
nor U15715 (N_15715,N_14524,N_14452);
xor U15716 (N_15716,N_14182,N_14700);
nor U15717 (N_15717,N_14236,N_14543);
nor U15718 (N_15718,N_14123,N_14149);
xor U15719 (N_15719,N_14913,N_14846);
xor U15720 (N_15720,N_14566,N_14258);
nand U15721 (N_15721,N_14802,N_14760);
or U15722 (N_15722,N_14188,N_14031);
or U15723 (N_15723,N_14497,N_14887);
nor U15724 (N_15724,N_14847,N_14526);
nor U15725 (N_15725,N_14552,N_14814);
nand U15726 (N_15726,N_14431,N_14664);
or U15727 (N_15727,N_14637,N_14190);
nor U15728 (N_15728,N_14941,N_14605);
nor U15729 (N_15729,N_14087,N_14939);
nand U15730 (N_15730,N_14602,N_14560);
and U15731 (N_15731,N_14090,N_14869);
nor U15732 (N_15732,N_14979,N_14824);
or U15733 (N_15733,N_14129,N_14693);
nand U15734 (N_15734,N_14168,N_14877);
and U15735 (N_15735,N_14086,N_14591);
nand U15736 (N_15736,N_14186,N_14341);
xnor U15737 (N_15737,N_14587,N_14858);
or U15738 (N_15738,N_14544,N_14541);
or U15739 (N_15739,N_14284,N_14297);
xnor U15740 (N_15740,N_14188,N_14203);
and U15741 (N_15741,N_14437,N_14289);
or U15742 (N_15742,N_14147,N_14512);
or U15743 (N_15743,N_14050,N_14231);
or U15744 (N_15744,N_14219,N_14802);
and U15745 (N_15745,N_14105,N_14846);
or U15746 (N_15746,N_14328,N_14900);
xor U15747 (N_15747,N_14309,N_14013);
nand U15748 (N_15748,N_14938,N_14610);
and U15749 (N_15749,N_14236,N_14170);
xnor U15750 (N_15750,N_14389,N_14865);
xnor U15751 (N_15751,N_14901,N_14752);
or U15752 (N_15752,N_14801,N_14250);
and U15753 (N_15753,N_14881,N_14314);
nor U15754 (N_15754,N_14947,N_14539);
nand U15755 (N_15755,N_14059,N_14871);
or U15756 (N_15756,N_14888,N_14868);
xor U15757 (N_15757,N_14418,N_14313);
or U15758 (N_15758,N_14578,N_14665);
nor U15759 (N_15759,N_14495,N_14333);
nor U15760 (N_15760,N_14696,N_14656);
nor U15761 (N_15761,N_14805,N_14478);
nor U15762 (N_15762,N_14402,N_14030);
and U15763 (N_15763,N_14296,N_14361);
or U15764 (N_15764,N_14293,N_14924);
or U15765 (N_15765,N_14018,N_14982);
and U15766 (N_15766,N_14485,N_14944);
nor U15767 (N_15767,N_14775,N_14973);
xor U15768 (N_15768,N_14364,N_14806);
and U15769 (N_15769,N_14096,N_14010);
or U15770 (N_15770,N_14999,N_14143);
nand U15771 (N_15771,N_14297,N_14287);
nor U15772 (N_15772,N_14287,N_14882);
nand U15773 (N_15773,N_14481,N_14540);
xor U15774 (N_15774,N_14505,N_14751);
or U15775 (N_15775,N_14905,N_14980);
or U15776 (N_15776,N_14625,N_14573);
xor U15777 (N_15777,N_14881,N_14198);
xnor U15778 (N_15778,N_14906,N_14642);
nor U15779 (N_15779,N_14506,N_14516);
nand U15780 (N_15780,N_14105,N_14708);
nor U15781 (N_15781,N_14871,N_14973);
nor U15782 (N_15782,N_14605,N_14544);
nor U15783 (N_15783,N_14971,N_14681);
nor U15784 (N_15784,N_14718,N_14971);
xnor U15785 (N_15785,N_14700,N_14517);
nor U15786 (N_15786,N_14123,N_14357);
nor U15787 (N_15787,N_14014,N_14622);
nand U15788 (N_15788,N_14800,N_14947);
xor U15789 (N_15789,N_14934,N_14862);
nand U15790 (N_15790,N_14758,N_14652);
nand U15791 (N_15791,N_14591,N_14387);
nand U15792 (N_15792,N_14506,N_14519);
nand U15793 (N_15793,N_14379,N_14466);
xnor U15794 (N_15794,N_14840,N_14942);
or U15795 (N_15795,N_14170,N_14025);
xor U15796 (N_15796,N_14737,N_14991);
nor U15797 (N_15797,N_14535,N_14272);
nor U15798 (N_15798,N_14430,N_14714);
nor U15799 (N_15799,N_14646,N_14035);
nand U15800 (N_15800,N_14007,N_14564);
nor U15801 (N_15801,N_14347,N_14573);
and U15802 (N_15802,N_14902,N_14161);
xnor U15803 (N_15803,N_14420,N_14464);
xor U15804 (N_15804,N_14427,N_14636);
xor U15805 (N_15805,N_14853,N_14156);
nand U15806 (N_15806,N_14574,N_14031);
and U15807 (N_15807,N_14016,N_14421);
or U15808 (N_15808,N_14192,N_14014);
and U15809 (N_15809,N_14681,N_14566);
nor U15810 (N_15810,N_14969,N_14865);
xnor U15811 (N_15811,N_14091,N_14467);
xnor U15812 (N_15812,N_14920,N_14365);
nor U15813 (N_15813,N_14351,N_14790);
or U15814 (N_15814,N_14786,N_14329);
or U15815 (N_15815,N_14089,N_14055);
or U15816 (N_15816,N_14821,N_14534);
or U15817 (N_15817,N_14937,N_14293);
and U15818 (N_15818,N_14842,N_14312);
and U15819 (N_15819,N_14365,N_14320);
and U15820 (N_15820,N_14745,N_14348);
and U15821 (N_15821,N_14492,N_14189);
or U15822 (N_15822,N_14927,N_14902);
xnor U15823 (N_15823,N_14897,N_14690);
xnor U15824 (N_15824,N_14465,N_14627);
nand U15825 (N_15825,N_14616,N_14503);
or U15826 (N_15826,N_14517,N_14662);
nand U15827 (N_15827,N_14613,N_14871);
nor U15828 (N_15828,N_14016,N_14069);
or U15829 (N_15829,N_14858,N_14641);
and U15830 (N_15830,N_14241,N_14444);
nor U15831 (N_15831,N_14827,N_14330);
and U15832 (N_15832,N_14428,N_14937);
or U15833 (N_15833,N_14590,N_14702);
and U15834 (N_15834,N_14832,N_14058);
nor U15835 (N_15835,N_14360,N_14058);
xor U15836 (N_15836,N_14825,N_14055);
nand U15837 (N_15837,N_14656,N_14812);
and U15838 (N_15838,N_14664,N_14420);
xor U15839 (N_15839,N_14206,N_14822);
nor U15840 (N_15840,N_14779,N_14983);
nor U15841 (N_15841,N_14960,N_14555);
nor U15842 (N_15842,N_14615,N_14317);
and U15843 (N_15843,N_14206,N_14261);
xnor U15844 (N_15844,N_14379,N_14091);
nand U15845 (N_15845,N_14408,N_14815);
xor U15846 (N_15846,N_14405,N_14209);
or U15847 (N_15847,N_14635,N_14305);
nand U15848 (N_15848,N_14279,N_14400);
or U15849 (N_15849,N_14375,N_14225);
and U15850 (N_15850,N_14000,N_14973);
xor U15851 (N_15851,N_14163,N_14257);
or U15852 (N_15852,N_14251,N_14204);
xor U15853 (N_15853,N_14783,N_14234);
nor U15854 (N_15854,N_14628,N_14471);
and U15855 (N_15855,N_14034,N_14261);
xor U15856 (N_15856,N_14228,N_14504);
xnor U15857 (N_15857,N_14095,N_14414);
nand U15858 (N_15858,N_14796,N_14138);
nand U15859 (N_15859,N_14341,N_14661);
xnor U15860 (N_15860,N_14426,N_14381);
and U15861 (N_15861,N_14580,N_14915);
xnor U15862 (N_15862,N_14721,N_14811);
nand U15863 (N_15863,N_14349,N_14924);
and U15864 (N_15864,N_14743,N_14679);
and U15865 (N_15865,N_14969,N_14249);
nor U15866 (N_15866,N_14066,N_14888);
nor U15867 (N_15867,N_14469,N_14283);
nor U15868 (N_15868,N_14874,N_14153);
nand U15869 (N_15869,N_14737,N_14398);
and U15870 (N_15870,N_14563,N_14237);
or U15871 (N_15871,N_14988,N_14252);
and U15872 (N_15872,N_14513,N_14135);
nor U15873 (N_15873,N_14865,N_14927);
or U15874 (N_15874,N_14465,N_14962);
xnor U15875 (N_15875,N_14887,N_14972);
nor U15876 (N_15876,N_14253,N_14766);
and U15877 (N_15877,N_14314,N_14889);
or U15878 (N_15878,N_14689,N_14106);
or U15879 (N_15879,N_14223,N_14317);
nor U15880 (N_15880,N_14608,N_14189);
xor U15881 (N_15881,N_14041,N_14282);
nor U15882 (N_15882,N_14738,N_14125);
and U15883 (N_15883,N_14355,N_14431);
nand U15884 (N_15884,N_14920,N_14117);
nand U15885 (N_15885,N_14665,N_14316);
xor U15886 (N_15886,N_14713,N_14898);
or U15887 (N_15887,N_14025,N_14500);
nand U15888 (N_15888,N_14559,N_14383);
xnor U15889 (N_15889,N_14026,N_14687);
or U15890 (N_15890,N_14646,N_14665);
or U15891 (N_15891,N_14729,N_14785);
nand U15892 (N_15892,N_14041,N_14945);
nand U15893 (N_15893,N_14976,N_14052);
xnor U15894 (N_15894,N_14241,N_14266);
nor U15895 (N_15895,N_14862,N_14933);
nand U15896 (N_15896,N_14475,N_14607);
or U15897 (N_15897,N_14454,N_14739);
or U15898 (N_15898,N_14088,N_14885);
nand U15899 (N_15899,N_14846,N_14983);
nor U15900 (N_15900,N_14380,N_14494);
or U15901 (N_15901,N_14341,N_14996);
or U15902 (N_15902,N_14875,N_14395);
or U15903 (N_15903,N_14012,N_14917);
nor U15904 (N_15904,N_14047,N_14399);
nor U15905 (N_15905,N_14848,N_14724);
nand U15906 (N_15906,N_14254,N_14291);
nand U15907 (N_15907,N_14953,N_14048);
or U15908 (N_15908,N_14731,N_14007);
or U15909 (N_15909,N_14998,N_14469);
and U15910 (N_15910,N_14317,N_14021);
nand U15911 (N_15911,N_14973,N_14662);
and U15912 (N_15912,N_14025,N_14097);
or U15913 (N_15913,N_14352,N_14623);
and U15914 (N_15914,N_14783,N_14976);
nor U15915 (N_15915,N_14402,N_14755);
nand U15916 (N_15916,N_14633,N_14043);
nor U15917 (N_15917,N_14300,N_14022);
or U15918 (N_15918,N_14650,N_14667);
nand U15919 (N_15919,N_14719,N_14375);
nand U15920 (N_15920,N_14881,N_14911);
and U15921 (N_15921,N_14647,N_14001);
xnor U15922 (N_15922,N_14168,N_14092);
or U15923 (N_15923,N_14459,N_14709);
nor U15924 (N_15924,N_14703,N_14490);
or U15925 (N_15925,N_14682,N_14366);
nand U15926 (N_15926,N_14508,N_14405);
nor U15927 (N_15927,N_14038,N_14970);
xor U15928 (N_15928,N_14547,N_14238);
xor U15929 (N_15929,N_14181,N_14648);
or U15930 (N_15930,N_14915,N_14278);
or U15931 (N_15931,N_14025,N_14153);
xor U15932 (N_15932,N_14139,N_14983);
nand U15933 (N_15933,N_14691,N_14169);
or U15934 (N_15934,N_14606,N_14415);
or U15935 (N_15935,N_14190,N_14306);
xnor U15936 (N_15936,N_14367,N_14440);
xor U15937 (N_15937,N_14547,N_14693);
nor U15938 (N_15938,N_14670,N_14553);
xor U15939 (N_15939,N_14512,N_14447);
nor U15940 (N_15940,N_14939,N_14966);
nor U15941 (N_15941,N_14750,N_14006);
nand U15942 (N_15942,N_14773,N_14575);
xnor U15943 (N_15943,N_14765,N_14182);
xor U15944 (N_15944,N_14057,N_14286);
xnor U15945 (N_15945,N_14026,N_14968);
or U15946 (N_15946,N_14498,N_14994);
nand U15947 (N_15947,N_14447,N_14784);
or U15948 (N_15948,N_14216,N_14725);
xnor U15949 (N_15949,N_14685,N_14227);
or U15950 (N_15950,N_14191,N_14193);
nand U15951 (N_15951,N_14817,N_14801);
xor U15952 (N_15952,N_14415,N_14235);
or U15953 (N_15953,N_14480,N_14163);
or U15954 (N_15954,N_14700,N_14003);
and U15955 (N_15955,N_14097,N_14955);
and U15956 (N_15956,N_14442,N_14501);
xnor U15957 (N_15957,N_14458,N_14097);
and U15958 (N_15958,N_14686,N_14095);
xnor U15959 (N_15959,N_14505,N_14803);
nand U15960 (N_15960,N_14913,N_14569);
and U15961 (N_15961,N_14919,N_14233);
nor U15962 (N_15962,N_14476,N_14086);
and U15963 (N_15963,N_14817,N_14768);
xnor U15964 (N_15964,N_14154,N_14226);
xnor U15965 (N_15965,N_14390,N_14476);
nor U15966 (N_15966,N_14204,N_14840);
and U15967 (N_15967,N_14080,N_14613);
and U15968 (N_15968,N_14600,N_14339);
nand U15969 (N_15969,N_14207,N_14975);
nor U15970 (N_15970,N_14246,N_14983);
nor U15971 (N_15971,N_14522,N_14053);
nor U15972 (N_15972,N_14251,N_14075);
or U15973 (N_15973,N_14255,N_14906);
or U15974 (N_15974,N_14000,N_14112);
nand U15975 (N_15975,N_14001,N_14970);
xor U15976 (N_15976,N_14064,N_14542);
nand U15977 (N_15977,N_14604,N_14230);
xnor U15978 (N_15978,N_14869,N_14467);
nand U15979 (N_15979,N_14937,N_14319);
nor U15980 (N_15980,N_14168,N_14920);
nand U15981 (N_15981,N_14426,N_14441);
nand U15982 (N_15982,N_14429,N_14587);
or U15983 (N_15983,N_14120,N_14649);
or U15984 (N_15984,N_14780,N_14428);
nor U15985 (N_15985,N_14040,N_14224);
and U15986 (N_15986,N_14492,N_14609);
or U15987 (N_15987,N_14778,N_14649);
xor U15988 (N_15988,N_14753,N_14421);
nor U15989 (N_15989,N_14979,N_14285);
and U15990 (N_15990,N_14804,N_14570);
or U15991 (N_15991,N_14720,N_14189);
nand U15992 (N_15992,N_14693,N_14633);
nand U15993 (N_15993,N_14888,N_14168);
and U15994 (N_15994,N_14480,N_14754);
xor U15995 (N_15995,N_14105,N_14838);
nor U15996 (N_15996,N_14153,N_14381);
and U15997 (N_15997,N_14371,N_14523);
xor U15998 (N_15998,N_14376,N_14112);
or U15999 (N_15999,N_14075,N_14385);
nor U16000 (N_16000,N_15218,N_15895);
xor U16001 (N_16001,N_15153,N_15745);
nand U16002 (N_16002,N_15064,N_15051);
nand U16003 (N_16003,N_15105,N_15724);
or U16004 (N_16004,N_15033,N_15622);
xor U16005 (N_16005,N_15385,N_15569);
or U16006 (N_16006,N_15847,N_15369);
and U16007 (N_16007,N_15907,N_15130);
and U16008 (N_16008,N_15615,N_15241);
and U16009 (N_16009,N_15499,N_15705);
nand U16010 (N_16010,N_15662,N_15640);
and U16011 (N_16011,N_15787,N_15276);
xor U16012 (N_16012,N_15523,N_15478);
nor U16013 (N_16013,N_15347,N_15883);
nor U16014 (N_16014,N_15498,N_15419);
xnor U16015 (N_16015,N_15901,N_15744);
nand U16016 (N_16016,N_15576,N_15384);
or U16017 (N_16017,N_15877,N_15976);
and U16018 (N_16018,N_15169,N_15422);
nand U16019 (N_16019,N_15725,N_15028);
and U16020 (N_16020,N_15626,N_15191);
and U16021 (N_16021,N_15958,N_15920);
or U16022 (N_16022,N_15565,N_15238);
or U16023 (N_16023,N_15339,N_15852);
nand U16024 (N_16024,N_15971,N_15819);
or U16025 (N_16025,N_15212,N_15860);
nand U16026 (N_16026,N_15167,N_15670);
nor U16027 (N_16027,N_15551,N_15287);
and U16028 (N_16028,N_15373,N_15991);
nor U16029 (N_16029,N_15682,N_15942);
nand U16030 (N_16030,N_15000,N_15442);
nand U16031 (N_16031,N_15633,N_15196);
nor U16032 (N_16032,N_15467,N_15572);
nand U16033 (N_16033,N_15372,N_15862);
xor U16034 (N_16034,N_15675,N_15468);
and U16035 (N_16035,N_15613,N_15823);
nand U16036 (N_16036,N_15150,N_15732);
nand U16037 (N_16037,N_15328,N_15597);
nand U16038 (N_16038,N_15762,N_15412);
xnor U16039 (N_16039,N_15588,N_15709);
xor U16040 (N_16040,N_15959,N_15790);
nand U16041 (N_16041,N_15444,N_15506);
xor U16042 (N_16042,N_15277,N_15164);
nor U16043 (N_16043,N_15261,N_15343);
xnor U16044 (N_16044,N_15786,N_15262);
xnor U16045 (N_16045,N_15831,N_15798);
or U16046 (N_16046,N_15059,N_15485);
nor U16047 (N_16047,N_15625,N_15249);
xor U16048 (N_16048,N_15538,N_15233);
xor U16049 (N_16049,N_15096,N_15101);
xnor U16050 (N_16050,N_15543,N_15484);
or U16051 (N_16051,N_15637,N_15294);
and U16052 (N_16052,N_15913,N_15402);
and U16053 (N_16053,N_15522,N_15863);
nor U16054 (N_16054,N_15309,N_15515);
nor U16055 (N_16055,N_15380,N_15307);
xor U16056 (N_16056,N_15691,N_15956);
or U16057 (N_16057,N_15677,N_15616);
nand U16058 (N_16058,N_15094,N_15184);
nand U16059 (N_16059,N_15041,N_15447);
nor U16060 (N_16060,N_15106,N_15519);
xor U16061 (N_16061,N_15200,N_15617);
or U16062 (N_16062,N_15337,N_15687);
nor U16063 (N_16063,N_15941,N_15301);
and U16064 (N_16064,N_15269,N_15175);
xor U16065 (N_16065,N_15793,N_15885);
xnor U16066 (N_16066,N_15118,N_15221);
or U16067 (N_16067,N_15076,N_15501);
xnor U16068 (N_16068,N_15610,N_15993);
and U16069 (N_16069,N_15162,N_15122);
or U16070 (N_16070,N_15336,N_15240);
xnor U16071 (N_16071,N_15836,N_15739);
nor U16072 (N_16072,N_15359,N_15205);
xor U16073 (N_16073,N_15231,N_15089);
or U16074 (N_16074,N_15654,N_15513);
and U16075 (N_16075,N_15652,N_15119);
xnor U16076 (N_16076,N_15393,N_15379);
nor U16077 (N_16077,N_15636,N_15356);
nor U16078 (N_16078,N_15845,N_15401);
nand U16079 (N_16079,N_15382,N_15018);
and U16080 (N_16080,N_15720,N_15248);
nor U16081 (N_16081,N_15701,N_15824);
nand U16082 (N_16082,N_15573,N_15367);
and U16083 (N_16083,N_15146,N_15607);
or U16084 (N_16084,N_15765,N_15110);
or U16085 (N_16085,N_15867,N_15230);
nor U16086 (N_16086,N_15044,N_15987);
and U16087 (N_16087,N_15002,N_15935);
xnor U16088 (N_16088,N_15896,N_15842);
nor U16089 (N_16089,N_15043,N_15158);
nor U16090 (N_16090,N_15776,N_15058);
nand U16091 (N_16091,N_15090,N_15788);
nand U16092 (N_16092,N_15255,N_15733);
or U16093 (N_16093,N_15143,N_15600);
xor U16094 (N_16094,N_15792,N_15668);
nand U16095 (N_16095,N_15156,N_15772);
and U16096 (N_16096,N_15360,N_15142);
and U16097 (N_16097,N_15536,N_15134);
and U16098 (N_16098,N_15507,N_15278);
nand U16099 (N_16099,N_15855,N_15562);
nand U16100 (N_16100,N_15057,N_15432);
or U16101 (N_16101,N_15243,N_15387);
nand U16102 (N_16102,N_15389,N_15570);
nand U16103 (N_16103,N_15390,N_15194);
and U16104 (N_16104,N_15838,N_15815);
nor U16105 (N_16105,N_15237,N_15025);
nor U16106 (N_16106,N_15296,N_15563);
and U16107 (N_16107,N_15921,N_15281);
xnor U16108 (N_16108,N_15868,N_15073);
nor U16109 (N_16109,N_15549,N_15056);
or U16110 (N_16110,N_15365,N_15049);
and U16111 (N_16111,N_15398,N_15446);
xor U16112 (N_16112,N_15348,N_15535);
or U16113 (N_16113,N_15140,N_15803);
and U16114 (N_16114,N_15689,N_15039);
xnor U16115 (N_16115,N_15545,N_15960);
xnor U16116 (N_16116,N_15195,N_15177);
xnor U16117 (N_16117,N_15334,N_15638);
xor U16118 (N_16118,N_15332,N_15108);
nor U16119 (N_16119,N_15310,N_15232);
nand U16120 (N_16120,N_15400,N_15857);
nand U16121 (N_16121,N_15813,N_15575);
nor U16122 (N_16122,N_15584,N_15273);
and U16123 (N_16123,N_15735,N_15804);
xnor U16124 (N_16124,N_15320,N_15297);
xnor U16125 (N_16125,N_15381,N_15411);
xnor U16126 (N_16126,N_15890,N_15554);
nor U16127 (N_16127,N_15770,N_15678);
nand U16128 (N_16128,N_15526,N_15290);
xor U16129 (N_16129,N_15247,N_15629);
and U16130 (N_16130,N_15107,N_15982);
or U16131 (N_16131,N_15875,N_15394);
nor U16132 (N_16132,N_15011,N_15567);
nor U16133 (N_16133,N_15820,N_15302);
and U16134 (N_16134,N_15954,N_15022);
or U16135 (N_16135,N_15590,N_15925);
or U16136 (N_16136,N_15013,N_15807);
or U16137 (N_16137,N_15985,N_15112);
or U16138 (N_16138,N_15226,N_15035);
and U16139 (N_16139,N_15173,N_15646);
nor U16140 (N_16140,N_15698,N_15727);
xor U16141 (N_16141,N_15658,N_15708);
or U16142 (N_16142,N_15561,N_15566);
and U16143 (N_16143,N_15653,N_15973);
or U16144 (N_16144,N_15253,N_15438);
or U16145 (N_16145,N_15854,N_15943);
and U16146 (N_16146,N_15785,N_15274);
xnor U16147 (N_16147,N_15746,N_15034);
xor U16148 (N_16148,N_15060,N_15126);
or U16149 (N_16149,N_15641,N_15665);
nand U16150 (N_16150,N_15496,N_15970);
xor U16151 (N_16151,N_15780,N_15109);
nand U16152 (N_16152,N_15583,N_15228);
xor U16153 (N_16153,N_15856,N_15601);
or U16154 (N_16154,N_15693,N_15783);
and U16155 (N_16155,N_15679,N_15703);
xnor U16156 (N_16156,N_15267,N_15796);
or U16157 (N_16157,N_15070,N_15279);
nor U16158 (N_16158,N_15455,N_15759);
nand U16159 (N_16159,N_15214,N_15898);
nand U16160 (N_16160,N_15266,N_15078);
or U16161 (N_16161,N_15087,N_15830);
nand U16162 (N_16162,N_15462,N_15222);
xor U16163 (N_16163,N_15858,N_15546);
or U16164 (N_16164,N_15475,N_15494);
nor U16165 (N_16165,N_15429,N_15292);
or U16166 (N_16166,N_15915,N_15331);
and U16167 (N_16167,N_15618,N_15789);
nand U16168 (N_16168,N_15069,N_15763);
and U16169 (N_16169,N_15283,N_15539);
nand U16170 (N_16170,N_15995,N_15428);
xor U16171 (N_16171,N_15316,N_15851);
and U16172 (N_16172,N_15964,N_15295);
nand U16173 (N_16173,N_15647,N_15782);
or U16174 (N_16174,N_15967,N_15225);
and U16175 (N_16175,N_15818,N_15312);
nand U16176 (N_16176,N_15902,N_15784);
nand U16177 (N_16177,N_15171,N_15945);
and U16178 (N_16178,N_15151,N_15514);
nand U16179 (N_16179,N_15293,N_15834);
and U16180 (N_16180,N_15799,N_15910);
and U16181 (N_16181,N_15377,N_15026);
or U16182 (N_16182,N_15254,N_15939);
nand U16183 (N_16183,N_15550,N_15046);
xnor U16184 (N_16184,N_15574,N_15651);
or U16185 (N_16185,N_15611,N_15750);
and U16186 (N_16186,N_15603,N_15947);
and U16187 (N_16187,N_15027,N_15932);
and U16188 (N_16188,N_15125,N_15085);
xor U16189 (N_16189,N_15702,N_15216);
and U16190 (N_16190,N_15355,N_15189);
or U16191 (N_16191,N_15628,N_15479);
xor U16192 (N_16192,N_15489,N_15155);
xor U16193 (N_16193,N_15362,N_15642);
and U16194 (N_16194,N_15716,N_15886);
nor U16195 (N_16195,N_15704,N_15751);
nor U16196 (N_16196,N_15366,N_15656);
nand U16197 (N_16197,N_15516,N_15361);
or U16198 (N_16198,N_15333,N_15257);
nand U16199 (N_16199,N_15869,N_15345);
nand U16200 (N_16200,N_15966,N_15053);
and U16201 (N_16201,N_15165,N_15284);
nand U16202 (N_16202,N_15614,N_15874);
or U16203 (N_16203,N_15001,N_15342);
xnor U16204 (N_16204,N_15508,N_15023);
and U16205 (N_16205,N_15850,N_15540);
nand U16206 (N_16206,N_15979,N_15975);
and U16207 (N_16207,N_15198,N_15029);
nand U16208 (N_16208,N_15463,N_15421);
xor U16209 (N_16209,N_15795,N_15676);
and U16210 (N_16210,N_15172,N_15871);
or U16211 (N_16211,N_15086,N_15594);
nor U16212 (N_16212,N_15884,N_15812);
xnor U16213 (N_16213,N_15929,N_15451);
or U16214 (N_16214,N_15048,N_15835);
xor U16215 (N_16215,N_15998,N_15912);
and U16216 (N_16216,N_15760,N_15344);
or U16217 (N_16217,N_15477,N_15694);
and U16218 (N_16218,N_15931,N_15256);
or U16219 (N_16219,N_15145,N_15435);
and U16220 (N_16220,N_15188,N_15800);
and U16221 (N_16221,N_15683,N_15341);
or U16222 (N_16222,N_15439,N_15873);
and U16223 (N_16223,N_15648,N_15075);
nand U16224 (N_16224,N_15473,N_15627);
nor U16225 (N_16225,N_15681,N_15436);
or U16226 (N_16226,N_15525,N_15826);
xor U16227 (N_16227,N_15892,N_15557);
nand U16228 (N_16228,N_15897,N_15923);
nor U16229 (N_16229,N_15120,N_15441);
nor U16230 (N_16230,N_15062,N_15327);
nand U16231 (N_16231,N_15181,N_15399);
nor U16232 (N_16232,N_15608,N_15488);
xor U16233 (N_16233,N_15459,N_15185);
nand U16234 (N_16234,N_15045,N_15391);
nand U16235 (N_16235,N_15992,N_15092);
or U16236 (N_16236,N_15866,N_15378);
nor U16237 (N_16237,N_15768,N_15580);
and U16238 (N_16238,N_15220,N_15215);
nand U16239 (N_16239,N_15012,N_15457);
or U16240 (N_16240,N_15055,N_15454);
xor U16241 (N_16241,N_15245,N_15286);
and U16242 (N_16242,N_15364,N_15493);
or U16243 (N_16243,N_15889,N_15458);
xnor U16244 (N_16244,N_15936,N_15685);
xor U16245 (N_16245,N_15953,N_15197);
or U16246 (N_16246,N_15081,N_15204);
nand U16247 (N_16247,N_15511,N_15052);
or U16248 (N_16248,N_15392,N_15100);
and U16249 (N_16249,N_15020,N_15133);
or U16250 (N_16250,N_15680,N_15406);
and U16251 (N_16251,N_15577,N_15427);
or U16252 (N_16252,N_15980,N_15235);
xnor U16253 (N_16253,N_15692,N_15848);
and U16254 (N_16254,N_15938,N_15994);
and U16255 (N_16255,N_15779,N_15955);
nand U16256 (N_16256,N_15909,N_15349);
and U16257 (N_16257,N_15265,N_15275);
nand U16258 (N_16258,N_15753,N_15797);
nor U16259 (N_16259,N_15403,N_15946);
nand U16260 (N_16260,N_15849,N_15911);
nand U16261 (N_16261,N_15778,N_15008);
or U16262 (N_16262,N_15542,N_15674);
xnor U16263 (N_16263,N_15322,N_15903);
and U16264 (N_16264,N_15121,N_15986);
xor U16265 (N_16265,N_15754,N_15844);
nand U16266 (N_16266,N_15031,N_15141);
nor U16267 (N_16267,N_15631,N_15099);
nand U16268 (N_16268,N_15213,N_15461);
or U16269 (N_16269,N_15717,N_15755);
xor U16270 (N_16270,N_15752,N_15553);
nand U16271 (N_16271,N_15258,N_15904);
xor U16272 (N_16272,N_15358,N_15019);
nor U16273 (N_16273,N_15635,N_15305);
and U16274 (N_16274,N_15906,N_15311);
nor U16275 (N_16275,N_15351,N_15015);
nor U16276 (N_16276,N_15518,N_15211);
nor U16277 (N_16277,N_15690,N_15729);
xnor U16278 (N_16278,N_15202,N_15127);
or U16279 (N_16279,N_15063,N_15456);
nand U16280 (N_16280,N_15919,N_15559);
nand U16281 (N_16281,N_15531,N_15529);
or U16282 (N_16282,N_15148,N_15227);
and U16283 (N_16283,N_15926,N_15916);
xnor U16284 (N_16284,N_15224,N_15123);
nand U16285 (N_16285,N_15252,N_15880);
and U16286 (N_16286,N_15131,N_15632);
or U16287 (N_16287,N_15952,N_15649);
or U16288 (N_16288,N_15758,N_15497);
xnor U16289 (N_16289,N_15908,N_15465);
xnor U16290 (N_16290,N_15132,N_15777);
or U16291 (N_16291,N_15605,N_15138);
and U16292 (N_16292,N_15180,N_15371);
or U16293 (N_16293,N_15599,N_15408);
nand U16294 (N_16294,N_15192,N_15304);
xor U16295 (N_16295,N_15009,N_15083);
nor U16296 (N_16296,N_15272,N_15114);
and U16297 (N_16297,N_15710,N_15289);
or U16298 (N_16298,N_15989,N_15639);
or U16299 (N_16299,N_15974,N_15537);
and U16300 (N_16300,N_15068,N_15071);
nor U16301 (N_16301,N_15407,N_15490);
or U16302 (N_16302,N_15541,N_15353);
nor U16303 (N_16303,N_15007,N_15756);
and U16304 (N_16304,N_15581,N_15509);
nor U16305 (N_16305,N_15630,N_15791);
and U16306 (N_16306,N_15282,N_15937);
and U16307 (N_16307,N_15452,N_15010);
xor U16308 (N_16308,N_15091,N_15234);
or U16309 (N_16309,N_15983,N_15821);
xnor U16310 (N_16310,N_15111,N_15667);
or U16311 (N_16311,N_15077,N_15891);
or U16312 (N_16312,N_15832,N_15259);
and U16313 (N_16313,N_15924,N_15969);
nand U16314 (N_16314,N_15288,N_15203);
nor U16315 (N_16315,N_15074,N_15718);
or U16316 (N_16316,N_15839,N_15104);
nand U16317 (N_16317,N_15161,N_15264);
nand U16318 (N_16318,N_15193,N_15723);
or U16319 (N_16319,N_15115,N_15655);
xor U16320 (N_16320,N_15659,N_15900);
or U16321 (N_16321,N_15159,N_15503);
or U16322 (N_16322,N_15715,N_15303);
or U16323 (N_16323,N_15579,N_15949);
xor U16324 (N_16324,N_15244,N_15491);
and U16325 (N_16325,N_15426,N_15928);
nor U16326 (N_16326,N_15298,N_15619);
and U16327 (N_16327,N_15775,N_15731);
or U16328 (N_16328,N_15673,N_15696);
and U16329 (N_16329,N_15449,N_15088);
or U16330 (N_16330,N_15314,N_15006);
nor U16331 (N_16331,N_15876,N_15250);
xnor U16332 (N_16332,N_15346,N_15829);
nand U16333 (N_16333,N_15512,N_15005);
or U16334 (N_16334,N_15672,N_15460);
nand U16335 (N_16335,N_15423,N_15740);
nand U16336 (N_16336,N_15853,N_15037);
xnor U16337 (N_16337,N_15781,N_15965);
or U16338 (N_16338,N_15065,N_15748);
xnor U16339 (N_16339,N_15922,N_15533);
and U16340 (N_16340,N_15340,N_15657);
xor U16341 (N_16341,N_15623,N_15067);
or U16342 (N_16342,N_15017,N_15808);
or U16343 (N_16343,N_15882,N_15410);
nor U16344 (N_16344,N_15480,N_15521);
nor U16345 (N_16345,N_15453,N_15219);
or U16346 (N_16346,N_15263,N_15395);
xnor U16347 (N_16347,N_15445,N_15040);
nand U16348 (N_16348,N_15814,N_15116);
nor U16349 (N_16349,N_15918,N_15388);
nor U16350 (N_16350,N_15981,N_15664);
xor U16351 (N_16351,N_15103,N_15686);
or U16352 (N_16352,N_15174,N_15734);
xor U16353 (N_16353,N_15036,N_15502);
nand U16354 (N_16354,N_15242,N_15944);
nor U16355 (N_16355,N_15139,N_15699);
xor U16356 (N_16356,N_15879,N_15749);
nor U16357 (N_16357,N_15236,N_15578);
or U16358 (N_16358,N_15082,N_15524);
nand U16359 (N_16359,N_15050,N_15547);
nand U16360 (N_16360,N_15738,N_15591);
and U16361 (N_16361,N_15335,N_15084);
nand U16362 (N_16362,N_15927,N_15977);
and U16363 (N_16363,N_15500,N_15968);
nand U16364 (N_16364,N_15021,N_15621);
or U16365 (N_16365,N_15285,N_15505);
xor U16366 (N_16366,N_15433,N_15766);
nand U16367 (N_16367,N_15471,N_15833);
or U16368 (N_16368,N_15246,N_15961);
xor U16369 (N_16369,N_15383,N_15963);
and U16370 (N_16370,N_15318,N_15870);
nand U16371 (N_16371,N_15650,N_15405);
and U16372 (N_16372,N_15917,N_15352);
or U16373 (N_16373,N_15510,N_15154);
xnor U16374 (N_16374,N_15129,N_15802);
nor U16375 (N_16375,N_15024,N_15308);
and U16376 (N_16376,N_15363,N_15135);
nor U16377 (N_16377,N_15859,N_15532);
or U16378 (N_16378,N_15984,N_15487);
and U16379 (N_16379,N_15595,N_15270);
nand U16380 (N_16380,N_15999,N_15714);
and U16381 (N_16381,N_15016,N_15737);
xor U16382 (N_16382,N_15157,N_15806);
nand U16383 (N_16383,N_15593,N_15558);
nor U16384 (N_16384,N_15817,N_15747);
xor U16385 (N_16385,N_15495,N_15801);
and U16386 (N_16386,N_15472,N_15688);
and U16387 (N_16387,N_15430,N_15773);
or U16388 (N_16388,N_15846,N_15014);
xnor U16389 (N_16389,N_15972,N_15329);
and U16390 (N_16390,N_15047,N_15606);
or U16391 (N_16391,N_15988,N_15396);
and U16392 (N_16392,N_15201,N_15386);
and U16393 (N_16393,N_15663,N_15571);
xor U16394 (N_16394,N_15431,N_15466);
or U16395 (N_16395,N_15742,N_15251);
nand U16396 (N_16396,N_15038,N_15093);
nand U16397 (N_16397,N_15186,N_15170);
nor U16398 (N_16398,N_15030,N_15684);
or U16399 (N_16399,N_15598,N_15416);
xor U16400 (N_16400,N_15713,N_15437);
xor U16401 (N_16401,N_15434,N_15997);
nor U16402 (N_16402,N_15179,N_15492);
xnor U16403 (N_16403,N_15774,N_15223);
xnor U16404 (N_16404,N_15424,N_15217);
nand U16405 (N_16405,N_15117,N_15210);
or U16406 (N_16406,N_15736,N_15767);
nor U16407 (N_16407,N_15888,N_15624);
and U16408 (N_16408,N_15299,N_15707);
nand U16409 (N_16409,N_15042,N_15079);
and U16410 (N_16410,N_15840,N_15899);
nor U16411 (N_16411,N_15761,N_15166);
or U16412 (N_16412,N_15003,N_15556);
or U16413 (N_16413,N_15951,N_15414);
nor U16414 (N_16414,N_15528,N_15990);
nand U16415 (N_16415,N_15054,N_15404);
and U16416 (N_16416,N_15661,N_15350);
xnor U16417 (N_16417,N_15602,N_15644);
nand U16418 (N_16418,N_15300,N_15881);
nor U16419 (N_16419,N_15124,N_15809);
nand U16420 (N_16420,N_15671,N_15147);
nor U16421 (N_16421,N_15187,N_15816);
nand U16422 (N_16422,N_15560,N_15905);
nand U16423 (N_16423,N_15319,N_15711);
nor U16424 (N_16424,N_15669,N_15828);
xnor U16425 (N_16425,N_15317,N_15530);
or U16426 (N_16426,N_15476,N_15004);
or U16427 (N_16427,N_15948,N_15837);
nand U16428 (N_16428,N_15183,N_15764);
nor U16429 (N_16429,N_15822,N_15861);
nand U16430 (N_16430,N_15587,N_15564);
or U16431 (N_16431,N_15470,N_15483);
nand U16432 (N_16432,N_15864,N_15592);
or U16433 (N_16433,N_15805,N_15719);
xnor U16434 (N_16434,N_15306,N_15865);
and U16435 (N_16435,N_15825,N_15374);
and U16436 (N_16436,N_15080,N_15527);
xor U16437 (N_16437,N_15113,N_15728);
xnor U16438 (N_16438,N_15418,N_15417);
and U16439 (N_16439,N_15137,N_15568);
nor U16440 (N_16440,N_15325,N_15887);
nand U16441 (N_16441,N_15596,N_15548);
and U16442 (N_16442,N_15324,N_15957);
or U16443 (N_16443,N_15190,N_15330);
nand U16444 (N_16444,N_15534,N_15695);
xor U16445 (N_16445,N_15586,N_15136);
nand U16446 (N_16446,N_15152,N_15271);
or U16447 (N_16447,N_15420,N_15811);
xor U16448 (N_16448,N_15095,N_15582);
or U16449 (N_16449,N_15409,N_15634);
or U16450 (N_16450,N_15930,N_15425);
nor U16451 (N_16451,N_15229,N_15712);
nor U16452 (N_16452,N_15149,N_15066);
or U16453 (N_16453,N_15097,N_15504);
or U16454 (N_16454,N_15643,N_15940);
nor U16455 (N_16455,N_15178,N_15326);
xnor U16456 (N_16456,N_15589,N_15260);
xor U16457 (N_16457,N_15168,N_15239);
or U16458 (N_16458,N_15950,N_15280);
and U16459 (N_16459,N_15552,N_15894);
and U16460 (N_16460,N_15102,N_15206);
and U16461 (N_16461,N_15722,N_15741);
nand U16462 (N_16462,N_15376,N_15323);
xnor U16463 (N_16463,N_15933,N_15827);
nand U16464 (N_16464,N_15448,N_15878);
and U16465 (N_16465,N_15207,N_15375);
xnor U16466 (N_16466,N_15486,N_15321);
nor U16467 (N_16467,N_15469,N_15128);
and U16468 (N_16468,N_15666,N_15700);
nand U16469 (N_16469,N_15338,N_15315);
and U16470 (N_16470,N_15368,N_15609);
or U16471 (N_16471,N_15706,N_15757);
or U16472 (N_16472,N_15585,N_15726);
and U16473 (N_16473,N_15464,N_15413);
xnor U16474 (N_16474,N_15199,N_15440);
and U16475 (N_16475,N_15841,N_15160);
or U16476 (N_16476,N_15697,N_15520);
xor U16477 (N_16477,N_15481,N_15604);
nand U16478 (N_16478,N_15357,N_15660);
nand U16479 (N_16479,N_15144,N_15645);
or U16480 (N_16480,N_15743,N_15354);
and U16481 (N_16481,N_15934,N_15313);
nand U16482 (N_16482,N_15443,N_15482);
and U16483 (N_16483,N_15370,N_15072);
nand U16484 (N_16484,N_15517,N_15996);
or U16485 (N_16485,N_15209,N_15032);
or U16486 (N_16486,N_15893,N_15978);
and U16487 (N_16487,N_15721,N_15163);
or U16488 (N_16488,N_15612,N_15415);
nor U16489 (N_16489,N_15182,N_15555);
or U16490 (N_16490,N_15098,N_15544);
and U16491 (N_16491,N_15176,N_15794);
nand U16492 (N_16492,N_15291,N_15843);
xnor U16493 (N_16493,N_15730,N_15771);
nand U16494 (N_16494,N_15061,N_15769);
and U16495 (N_16495,N_15914,N_15397);
nor U16496 (N_16496,N_15450,N_15872);
and U16497 (N_16497,N_15474,N_15620);
xor U16498 (N_16498,N_15810,N_15208);
nor U16499 (N_16499,N_15268,N_15962);
or U16500 (N_16500,N_15645,N_15400);
nor U16501 (N_16501,N_15289,N_15148);
and U16502 (N_16502,N_15381,N_15148);
nor U16503 (N_16503,N_15537,N_15165);
nor U16504 (N_16504,N_15877,N_15716);
xnor U16505 (N_16505,N_15693,N_15650);
or U16506 (N_16506,N_15083,N_15984);
nand U16507 (N_16507,N_15217,N_15076);
nand U16508 (N_16508,N_15556,N_15643);
nand U16509 (N_16509,N_15384,N_15843);
xor U16510 (N_16510,N_15373,N_15594);
nand U16511 (N_16511,N_15041,N_15066);
and U16512 (N_16512,N_15790,N_15047);
xor U16513 (N_16513,N_15598,N_15746);
nor U16514 (N_16514,N_15181,N_15901);
xor U16515 (N_16515,N_15088,N_15622);
and U16516 (N_16516,N_15473,N_15317);
nor U16517 (N_16517,N_15357,N_15975);
nor U16518 (N_16518,N_15883,N_15922);
xor U16519 (N_16519,N_15205,N_15884);
and U16520 (N_16520,N_15923,N_15908);
and U16521 (N_16521,N_15665,N_15820);
nor U16522 (N_16522,N_15778,N_15463);
nor U16523 (N_16523,N_15434,N_15328);
nand U16524 (N_16524,N_15817,N_15560);
or U16525 (N_16525,N_15188,N_15972);
xnor U16526 (N_16526,N_15969,N_15565);
or U16527 (N_16527,N_15777,N_15272);
nor U16528 (N_16528,N_15923,N_15215);
xnor U16529 (N_16529,N_15356,N_15740);
nor U16530 (N_16530,N_15759,N_15107);
nor U16531 (N_16531,N_15297,N_15243);
and U16532 (N_16532,N_15888,N_15871);
nand U16533 (N_16533,N_15707,N_15795);
and U16534 (N_16534,N_15828,N_15468);
xor U16535 (N_16535,N_15158,N_15568);
xnor U16536 (N_16536,N_15772,N_15645);
or U16537 (N_16537,N_15733,N_15855);
nand U16538 (N_16538,N_15765,N_15532);
or U16539 (N_16539,N_15129,N_15626);
nand U16540 (N_16540,N_15407,N_15561);
or U16541 (N_16541,N_15190,N_15084);
xor U16542 (N_16542,N_15360,N_15078);
or U16543 (N_16543,N_15068,N_15453);
or U16544 (N_16544,N_15145,N_15424);
xnor U16545 (N_16545,N_15615,N_15473);
or U16546 (N_16546,N_15137,N_15141);
xnor U16547 (N_16547,N_15372,N_15991);
nor U16548 (N_16548,N_15402,N_15974);
xor U16549 (N_16549,N_15816,N_15325);
nand U16550 (N_16550,N_15510,N_15503);
or U16551 (N_16551,N_15774,N_15494);
xnor U16552 (N_16552,N_15070,N_15002);
nand U16553 (N_16553,N_15011,N_15787);
nand U16554 (N_16554,N_15723,N_15624);
and U16555 (N_16555,N_15157,N_15889);
or U16556 (N_16556,N_15279,N_15927);
and U16557 (N_16557,N_15793,N_15873);
or U16558 (N_16558,N_15805,N_15312);
nor U16559 (N_16559,N_15571,N_15057);
xnor U16560 (N_16560,N_15821,N_15680);
nor U16561 (N_16561,N_15291,N_15922);
xor U16562 (N_16562,N_15259,N_15137);
or U16563 (N_16563,N_15546,N_15809);
xor U16564 (N_16564,N_15513,N_15738);
nor U16565 (N_16565,N_15746,N_15826);
nand U16566 (N_16566,N_15861,N_15650);
and U16567 (N_16567,N_15085,N_15258);
xnor U16568 (N_16568,N_15510,N_15301);
or U16569 (N_16569,N_15178,N_15983);
and U16570 (N_16570,N_15773,N_15781);
nor U16571 (N_16571,N_15981,N_15678);
nor U16572 (N_16572,N_15316,N_15798);
and U16573 (N_16573,N_15313,N_15686);
or U16574 (N_16574,N_15494,N_15305);
nand U16575 (N_16575,N_15428,N_15598);
xor U16576 (N_16576,N_15371,N_15576);
nand U16577 (N_16577,N_15632,N_15227);
or U16578 (N_16578,N_15822,N_15572);
nor U16579 (N_16579,N_15025,N_15648);
or U16580 (N_16580,N_15487,N_15792);
nor U16581 (N_16581,N_15361,N_15382);
nand U16582 (N_16582,N_15583,N_15380);
nor U16583 (N_16583,N_15587,N_15678);
and U16584 (N_16584,N_15310,N_15050);
nor U16585 (N_16585,N_15886,N_15457);
or U16586 (N_16586,N_15504,N_15955);
or U16587 (N_16587,N_15555,N_15081);
nor U16588 (N_16588,N_15426,N_15296);
or U16589 (N_16589,N_15395,N_15587);
nor U16590 (N_16590,N_15773,N_15242);
xor U16591 (N_16591,N_15830,N_15517);
xnor U16592 (N_16592,N_15490,N_15395);
nand U16593 (N_16593,N_15255,N_15524);
or U16594 (N_16594,N_15174,N_15468);
nor U16595 (N_16595,N_15573,N_15683);
nor U16596 (N_16596,N_15747,N_15506);
or U16597 (N_16597,N_15414,N_15421);
nor U16598 (N_16598,N_15597,N_15389);
nand U16599 (N_16599,N_15853,N_15774);
nand U16600 (N_16600,N_15895,N_15026);
xnor U16601 (N_16601,N_15335,N_15131);
and U16602 (N_16602,N_15341,N_15358);
or U16603 (N_16603,N_15161,N_15637);
nor U16604 (N_16604,N_15134,N_15843);
nand U16605 (N_16605,N_15882,N_15029);
nand U16606 (N_16606,N_15241,N_15969);
xor U16607 (N_16607,N_15220,N_15274);
nand U16608 (N_16608,N_15342,N_15145);
xnor U16609 (N_16609,N_15062,N_15526);
xor U16610 (N_16610,N_15848,N_15105);
and U16611 (N_16611,N_15317,N_15056);
or U16612 (N_16612,N_15809,N_15034);
nand U16613 (N_16613,N_15573,N_15359);
nand U16614 (N_16614,N_15930,N_15805);
nand U16615 (N_16615,N_15705,N_15628);
and U16616 (N_16616,N_15094,N_15318);
or U16617 (N_16617,N_15435,N_15808);
xor U16618 (N_16618,N_15504,N_15228);
nand U16619 (N_16619,N_15270,N_15179);
xnor U16620 (N_16620,N_15059,N_15654);
or U16621 (N_16621,N_15950,N_15161);
xor U16622 (N_16622,N_15619,N_15375);
nor U16623 (N_16623,N_15380,N_15425);
xnor U16624 (N_16624,N_15396,N_15266);
or U16625 (N_16625,N_15475,N_15570);
nand U16626 (N_16626,N_15978,N_15650);
nand U16627 (N_16627,N_15373,N_15469);
or U16628 (N_16628,N_15893,N_15662);
nor U16629 (N_16629,N_15220,N_15998);
or U16630 (N_16630,N_15848,N_15925);
or U16631 (N_16631,N_15777,N_15771);
xnor U16632 (N_16632,N_15759,N_15190);
or U16633 (N_16633,N_15777,N_15737);
nor U16634 (N_16634,N_15925,N_15751);
or U16635 (N_16635,N_15879,N_15364);
and U16636 (N_16636,N_15916,N_15584);
and U16637 (N_16637,N_15971,N_15149);
xor U16638 (N_16638,N_15963,N_15796);
or U16639 (N_16639,N_15733,N_15148);
and U16640 (N_16640,N_15704,N_15508);
nand U16641 (N_16641,N_15708,N_15837);
or U16642 (N_16642,N_15253,N_15357);
and U16643 (N_16643,N_15757,N_15250);
or U16644 (N_16644,N_15921,N_15258);
nand U16645 (N_16645,N_15912,N_15898);
nor U16646 (N_16646,N_15943,N_15539);
or U16647 (N_16647,N_15658,N_15282);
and U16648 (N_16648,N_15636,N_15175);
xnor U16649 (N_16649,N_15971,N_15153);
and U16650 (N_16650,N_15382,N_15509);
and U16651 (N_16651,N_15853,N_15596);
nand U16652 (N_16652,N_15130,N_15812);
and U16653 (N_16653,N_15311,N_15513);
or U16654 (N_16654,N_15332,N_15291);
or U16655 (N_16655,N_15866,N_15680);
nand U16656 (N_16656,N_15246,N_15369);
or U16657 (N_16657,N_15399,N_15558);
nor U16658 (N_16658,N_15644,N_15584);
nor U16659 (N_16659,N_15124,N_15219);
nor U16660 (N_16660,N_15156,N_15216);
nor U16661 (N_16661,N_15407,N_15601);
xor U16662 (N_16662,N_15755,N_15380);
and U16663 (N_16663,N_15977,N_15563);
nand U16664 (N_16664,N_15920,N_15969);
and U16665 (N_16665,N_15328,N_15430);
xnor U16666 (N_16666,N_15634,N_15725);
or U16667 (N_16667,N_15727,N_15118);
nor U16668 (N_16668,N_15977,N_15519);
or U16669 (N_16669,N_15633,N_15249);
nor U16670 (N_16670,N_15018,N_15338);
nand U16671 (N_16671,N_15286,N_15188);
nand U16672 (N_16672,N_15315,N_15163);
nor U16673 (N_16673,N_15475,N_15477);
or U16674 (N_16674,N_15182,N_15492);
nand U16675 (N_16675,N_15638,N_15530);
or U16676 (N_16676,N_15197,N_15300);
and U16677 (N_16677,N_15319,N_15998);
xnor U16678 (N_16678,N_15093,N_15112);
or U16679 (N_16679,N_15540,N_15914);
and U16680 (N_16680,N_15537,N_15375);
nor U16681 (N_16681,N_15437,N_15200);
nor U16682 (N_16682,N_15468,N_15489);
nor U16683 (N_16683,N_15441,N_15981);
nand U16684 (N_16684,N_15001,N_15435);
nand U16685 (N_16685,N_15440,N_15461);
nor U16686 (N_16686,N_15656,N_15851);
nand U16687 (N_16687,N_15352,N_15383);
or U16688 (N_16688,N_15444,N_15571);
nand U16689 (N_16689,N_15306,N_15678);
nor U16690 (N_16690,N_15597,N_15669);
and U16691 (N_16691,N_15461,N_15559);
nor U16692 (N_16692,N_15891,N_15948);
nand U16693 (N_16693,N_15030,N_15371);
nor U16694 (N_16694,N_15845,N_15697);
nand U16695 (N_16695,N_15574,N_15913);
xor U16696 (N_16696,N_15695,N_15956);
nor U16697 (N_16697,N_15142,N_15737);
and U16698 (N_16698,N_15035,N_15222);
nand U16699 (N_16699,N_15118,N_15845);
nor U16700 (N_16700,N_15526,N_15982);
nor U16701 (N_16701,N_15947,N_15940);
and U16702 (N_16702,N_15808,N_15057);
nor U16703 (N_16703,N_15518,N_15406);
xor U16704 (N_16704,N_15161,N_15101);
or U16705 (N_16705,N_15425,N_15938);
xor U16706 (N_16706,N_15659,N_15987);
xnor U16707 (N_16707,N_15499,N_15806);
or U16708 (N_16708,N_15139,N_15033);
nand U16709 (N_16709,N_15229,N_15527);
nand U16710 (N_16710,N_15375,N_15600);
or U16711 (N_16711,N_15597,N_15011);
nand U16712 (N_16712,N_15467,N_15318);
xnor U16713 (N_16713,N_15691,N_15312);
nor U16714 (N_16714,N_15896,N_15634);
or U16715 (N_16715,N_15259,N_15484);
nor U16716 (N_16716,N_15505,N_15902);
nor U16717 (N_16717,N_15360,N_15805);
nand U16718 (N_16718,N_15772,N_15273);
nor U16719 (N_16719,N_15168,N_15463);
or U16720 (N_16720,N_15398,N_15692);
xnor U16721 (N_16721,N_15267,N_15293);
nor U16722 (N_16722,N_15912,N_15805);
nor U16723 (N_16723,N_15944,N_15542);
and U16724 (N_16724,N_15966,N_15961);
nand U16725 (N_16725,N_15761,N_15087);
xnor U16726 (N_16726,N_15509,N_15167);
nor U16727 (N_16727,N_15564,N_15710);
nand U16728 (N_16728,N_15999,N_15013);
or U16729 (N_16729,N_15939,N_15103);
xnor U16730 (N_16730,N_15703,N_15503);
nand U16731 (N_16731,N_15846,N_15439);
and U16732 (N_16732,N_15557,N_15917);
xnor U16733 (N_16733,N_15902,N_15292);
nand U16734 (N_16734,N_15785,N_15465);
or U16735 (N_16735,N_15361,N_15581);
or U16736 (N_16736,N_15105,N_15081);
nor U16737 (N_16737,N_15470,N_15711);
or U16738 (N_16738,N_15446,N_15418);
and U16739 (N_16739,N_15493,N_15043);
xor U16740 (N_16740,N_15414,N_15678);
xor U16741 (N_16741,N_15915,N_15541);
nor U16742 (N_16742,N_15088,N_15284);
or U16743 (N_16743,N_15478,N_15485);
or U16744 (N_16744,N_15765,N_15017);
nor U16745 (N_16745,N_15285,N_15182);
xor U16746 (N_16746,N_15458,N_15872);
nand U16747 (N_16747,N_15014,N_15485);
nand U16748 (N_16748,N_15392,N_15639);
xor U16749 (N_16749,N_15655,N_15475);
and U16750 (N_16750,N_15939,N_15388);
or U16751 (N_16751,N_15670,N_15475);
nand U16752 (N_16752,N_15631,N_15492);
and U16753 (N_16753,N_15375,N_15377);
or U16754 (N_16754,N_15992,N_15994);
nand U16755 (N_16755,N_15343,N_15435);
and U16756 (N_16756,N_15604,N_15971);
or U16757 (N_16757,N_15741,N_15870);
or U16758 (N_16758,N_15039,N_15316);
nor U16759 (N_16759,N_15471,N_15858);
xor U16760 (N_16760,N_15439,N_15912);
xnor U16761 (N_16761,N_15567,N_15475);
or U16762 (N_16762,N_15546,N_15163);
nor U16763 (N_16763,N_15923,N_15730);
and U16764 (N_16764,N_15924,N_15063);
or U16765 (N_16765,N_15941,N_15369);
nand U16766 (N_16766,N_15633,N_15394);
and U16767 (N_16767,N_15017,N_15366);
nor U16768 (N_16768,N_15437,N_15359);
xor U16769 (N_16769,N_15569,N_15652);
and U16770 (N_16770,N_15819,N_15304);
xnor U16771 (N_16771,N_15263,N_15667);
xnor U16772 (N_16772,N_15955,N_15717);
and U16773 (N_16773,N_15954,N_15546);
and U16774 (N_16774,N_15499,N_15335);
nor U16775 (N_16775,N_15597,N_15876);
or U16776 (N_16776,N_15932,N_15429);
or U16777 (N_16777,N_15291,N_15585);
nor U16778 (N_16778,N_15373,N_15092);
nand U16779 (N_16779,N_15032,N_15104);
nand U16780 (N_16780,N_15460,N_15057);
or U16781 (N_16781,N_15538,N_15254);
and U16782 (N_16782,N_15840,N_15087);
and U16783 (N_16783,N_15621,N_15023);
or U16784 (N_16784,N_15474,N_15217);
nor U16785 (N_16785,N_15649,N_15573);
nand U16786 (N_16786,N_15918,N_15387);
nand U16787 (N_16787,N_15981,N_15748);
or U16788 (N_16788,N_15555,N_15451);
nor U16789 (N_16789,N_15763,N_15578);
nand U16790 (N_16790,N_15848,N_15481);
nand U16791 (N_16791,N_15164,N_15834);
xnor U16792 (N_16792,N_15697,N_15774);
nand U16793 (N_16793,N_15862,N_15423);
xor U16794 (N_16794,N_15064,N_15020);
or U16795 (N_16795,N_15179,N_15821);
nor U16796 (N_16796,N_15678,N_15787);
xnor U16797 (N_16797,N_15543,N_15968);
nor U16798 (N_16798,N_15913,N_15754);
nor U16799 (N_16799,N_15544,N_15466);
nand U16800 (N_16800,N_15250,N_15470);
or U16801 (N_16801,N_15159,N_15743);
xnor U16802 (N_16802,N_15618,N_15165);
xor U16803 (N_16803,N_15609,N_15082);
or U16804 (N_16804,N_15318,N_15606);
or U16805 (N_16805,N_15087,N_15096);
nand U16806 (N_16806,N_15627,N_15858);
nand U16807 (N_16807,N_15638,N_15751);
nand U16808 (N_16808,N_15150,N_15355);
xnor U16809 (N_16809,N_15228,N_15864);
nor U16810 (N_16810,N_15857,N_15101);
or U16811 (N_16811,N_15122,N_15936);
xor U16812 (N_16812,N_15986,N_15087);
xnor U16813 (N_16813,N_15444,N_15157);
or U16814 (N_16814,N_15546,N_15146);
and U16815 (N_16815,N_15177,N_15964);
or U16816 (N_16816,N_15753,N_15008);
nand U16817 (N_16817,N_15003,N_15633);
nor U16818 (N_16818,N_15606,N_15182);
and U16819 (N_16819,N_15953,N_15387);
nand U16820 (N_16820,N_15854,N_15810);
or U16821 (N_16821,N_15002,N_15178);
and U16822 (N_16822,N_15688,N_15692);
nand U16823 (N_16823,N_15032,N_15066);
nor U16824 (N_16824,N_15879,N_15939);
or U16825 (N_16825,N_15874,N_15680);
and U16826 (N_16826,N_15130,N_15984);
and U16827 (N_16827,N_15324,N_15500);
nand U16828 (N_16828,N_15651,N_15961);
or U16829 (N_16829,N_15451,N_15419);
and U16830 (N_16830,N_15383,N_15471);
xnor U16831 (N_16831,N_15004,N_15087);
and U16832 (N_16832,N_15536,N_15689);
nor U16833 (N_16833,N_15988,N_15127);
nand U16834 (N_16834,N_15709,N_15316);
and U16835 (N_16835,N_15059,N_15942);
nor U16836 (N_16836,N_15070,N_15182);
and U16837 (N_16837,N_15865,N_15741);
nand U16838 (N_16838,N_15692,N_15469);
nand U16839 (N_16839,N_15658,N_15474);
and U16840 (N_16840,N_15299,N_15644);
nor U16841 (N_16841,N_15655,N_15328);
xor U16842 (N_16842,N_15278,N_15122);
nor U16843 (N_16843,N_15610,N_15976);
xor U16844 (N_16844,N_15203,N_15072);
xnor U16845 (N_16845,N_15383,N_15593);
nand U16846 (N_16846,N_15371,N_15109);
nor U16847 (N_16847,N_15151,N_15073);
xor U16848 (N_16848,N_15869,N_15579);
and U16849 (N_16849,N_15207,N_15576);
nand U16850 (N_16850,N_15210,N_15721);
nor U16851 (N_16851,N_15168,N_15627);
and U16852 (N_16852,N_15692,N_15424);
nand U16853 (N_16853,N_15570,N_15990);
or U16854 (N_16854,N_15946,N_15710);
xnor U16855 (N_16855,N_15157,N_15640);
or U16856 (N_16856,N_15173,N_15923);
nand U16857 (N_16857,N_15272,N_15478);
xnor U16858 (N_16858,N_15143,N_15458);
nor U16859 (N_16859,N_15088,N_15061);
xor U16860 (N_16860,N_15205,N_15949);
xor U16861 (N_16861,N_15723,N_15183);
xnor U16862 (N_16862,N_15295,N_15700);
xor U16863 (N_16863,N_15411,N_15835);
nand U16864 (N_16864,N_15085,N_15008);
xor U16865 (N_16865,N_15416,N_15807);
and U16866 (N_16866,N_15762,N_15928);
and U16867 (N_16867,N_15104,N_15760);
xnor U16868 (N_16868,N_15510,N_15570);
and U16869 (N_16869,N_15045,N_15993);
and U16870 (N_16870,N_15366,N_15891);
nor U16871 (N_16871,N_15434,N_15198);
and U16872 (N_16872,N_15630,N_15185);
xnor U16873 (N_16873,N_15380,N_15699);
xnor U16874 (N_16874,N_15865,N_15442);
xor U16875 (N_16875,N_15476,N_15387);
nand U16876 (N_16876,N_15883,N_15665);
nor U16877 (N_16877,N_15659,N_15652);
xor U16878 (N_16878,N_15485,N_15129);
xor U16879 (N_16879,N_15551,N_15014);
or U16880 (N_16880,N_15660,N_15935);
nor U16881 (N_16881,N_15428,N_15469);
and U16882 (N_16882,N_15179,N_15683);
or U16883 (N_16883,N_15806,N_15325);
and U16884 (N_16884,N_15823,N_15429);
and U16885 (N_16885,N_15439,N_15671);
and U16886 (N_16886,N_15729,N_15699);
xor U16887 (N_16887,N_15148,N_15493);
or U16888 (N_16888,N_15698,N_15770);
nand U16889 (N_16889,N_15600,N_15544);
xor U16890 (N_16890,N_15422,N_15746);
or U16891 (N_16891,N_15537,N_15339);
nor U16892 (N_16892,N_15259,N_15232);
nor U16893 (N_16893,N_15529,N_15411);
nand U16894 (N_16894,N_15689,N_15031);
or U16895 (N_16895,N_15840,N_15143);
and U16896 (N_16896,N_15113,N_15076);
or U16897 (N_16897,N_15334,N_15864);
nand U16898 (N_16898,N_15832,N_15428);
xor U16899 (N_16899,N_15508,N_15150);
or U16900 (N_16900,N_15860,N_15312);
nor U16901 (N_16901,N_15910,N_15117);
nor U16902 (N_16902,N_15481,N_15412);
nand U16903 (N_16903,N_15256,N_15077);
nand U16904 (N_16904,N_15549,N_15979);
xor U16905 (N_16905,N_15872,N_15524);
or U16906 (N_16906,N_15741,N_15145);
nand U16907 (N_16907,N_15751,N_15029);
xnor U16908 (N_16908,N_15398,N_15480);
xnor U16909 (N_16909,N_15887,N_15011);
and U16910 (N_16910,N_15326,N_15670);
nand U16911 (N_16911,N_15165,N_15603);
nand U16912 (N_16912,N_15902,N_15227);
and U16913 (N_16913,N_15577,N_15629);
xor U16914 (N_16914,N_15960,N_15143);
xnor U16915 (N_16915,N_15419,N_15641);
xnor U16916 (N_16916,N_15126,N_15241);
nor U16917 (N_16917,N_15795,N_15291);
xnor U16918 (N_16918,N_15989,N_15614);
xor U16919 (N_16919,N_15453,N_15475);
or U16920 (N_16920,N_15444,N_15676);
nand U16921 (N_16921,N_15546,N_15378);
xnor U16922 (N_16922,N_15779,N_15231);
and U16923 (N_16923,N_15406,N_15165);
and U16924 (N_16924,N_15843,N_15074);
xnor U16925 (N_16925,N_15264,N_15441);
and U16926 (N_16926,N_15284,N_15398);
nor U16927 (N_16927,N_15615,N_15675);
or U16928 (N_16928,N_15854,N_15507);
xor U16929 (N_16929,N_15926,N_15197);
or U16930 (N_16930,N_15314,N_15606);
nand U16931 (N_16931,N_15354,N_15649);
or U16932 (N_16932,N_15359,N_15785);
xnor U16933 (N_16933,N_15030,N_15707);
or U16934 (N_16934,N_15996,N_15935);
nor U16935 (N_16935,N_15997,N_15708);
xnor U16936 (N_16936,N_15388,N_15724);
xor U16937 (N_16937,N_15900,N_15337);
and U16938 (N_16938,N_15499,N_15412);
and U16939 (N_16939,N_15298,N_15412);
and U16940 (N_16940,N_15221,N_15031);
or U16941 (N_16941,N_15124,N_15053);
xor U16942 (N_16942,N_15689,N_15103);
or U16943 (N_16943,N_15299,N_15030);
or U16944 (N_16944,N_15009,N_15431);
nor U16945 (N_16945,N_15265,N_15008);
and U16946 (N_16946,N_15379,N_15693);
nand U16947 (N_16947,N_15649,N_15219);
xor U16948 (N_16948,N_15190,N_15166);
nand U16949 (N_16949,N_15160,N_15743);
xnor U16950 (N_16950,N_15258,N_15597);
and U16951 (N_16951,N_15802,N_15961);
xor U16952 (N_16952,N_15910,N_15284);
or U16953 (N_16953,N_15356,N_15690);
and U16954 (N_16954,N_15148,N_15394);
nor U16955 (N_16955,N_15616,N_15924);
or U16956 (N_16956,N_15836,N_15011);
nor U16957 (N_16957,N_15497,N_15592);
nor U16958 (N_16958,N_15557,N_15263);
or U16959 (N_16959,N_15951,N_15620);
or U16960 (N_16960,N_15688,N_15305);
xor U16961 (N_16961,N_15991,N_15538);
nand U16962 (N_16962,N_15979,N_15097);
or U16963 (N_16963,N_15400,N_15203);
nand U16964 (N_16964,N_15334,N_15233);
nor U16965 (N_16965,N_15469,N_15347);
nor U16966 (N_16966,N_15812,N_15180);
nor U16967 (N_16967,N_15494,N_15920);
nor U16968 (N_16968,N_15303,N_15434);
nor U16969 (N_16969,N_15162,N_15013);
nor U16970 (N_16970,N_15452,N_15070);
and U16971 (N_16971,N_15170,N_15631);
nor U16972 (N_16972,N_15968,N_15265);
and U16973 (N_16973,N_15912,N_15223);
xor U16974 (N_16974,N_15036,N_15483);
or U16975 (N_16975,N_15481,N_15158);
xor U16976 (N_16976,N_15276,N_15002);
or U16977 (N_16977,N_15145,N_15679);
xnor U16978 (N_16978,N_15925,N_15473);
nand U16979 (N_16979,N_15400,N_15098);
xnor U16980 (N_16980,N_15945,N_15179);
nand U16981 (N_16981,N_15446,N_15675);
nor U16982 (N_16982,N_15082,N_15383);
nand U16983 (N_16983,N_15636,N_15791);
and U16984 (N_16984,N_15712,N_15210);
and U16985 (N_16985,N_15496,N_15191);
and U16986 (N_16986,N_15338,N_15562);
and U16987 (N_16987,N_15235,N_15825);
nand U16988 (N_16988,N_15792,N_15566);
or U16989 (N_16989,N_15741,N_15727);
xnor U16990 (N_16990,N_15593,N_15489);
nor U16991 (N_16991,N_15264,N_15035);
nor U16992 (N_16992,N_15228,N_15818);
nand U16993 (N_16993,N_15243,N_15682);
nor U16994 (N_16994,N_15621,N_15465);
and U16995 (N_16995,N_15446,N_15927);
nor U16996 (N_16996,N_15195,N_15947);
nor U16997 (N_16997,N_15361,N_15131);
nor U16998 (N_16998,N_15500,N_15353);
and U16999 (N_16999,N_15409,N_15960);
nor U17000 (N_17000,N_16209,N_16869);
nor U17001 (N_17001,N_16492,N_16483);
nor U17002 (N_17002,N_16373,N_16232);
and U17003 (N_17003,N_16047,N_16838);
nand U17004 (N_17004,N_16762,N_16225);
nand U17005 (N_17005,N_16545,N_16823);
nand U17006 (N_17006,N_16464,N_16247);
or U17007 (N_17007,N_16864,N_16158);
xor U17008 (N_17008,N_16773,N_16202);
xor U17009 (N_17009,N_16485,N_16767);
nand U17010 (N_17010,N_16587,N_16080);
nand U17011 (N_17011,N_16768,N_16295);
nand U17012 (N_17012,N_16913,N_16234);
nand U17013 (N_17013,N_16365,N_16652);
nand U17014 (N_17014,N_16064,N_16764);
nor U17015 (N_17015,N_16037,N_16125);
nand U17016 (N_17016,N_16650,N_16299);
nor U17017 (N_17017,N_16458,N_16572);
nor U17018 (N_17018,N_16756,N_16059);
or U17019 (N_17019,N_16834,N_16555);
nand U17020 (N_17020,N_16244,N_16355);
nand U17021 (N_17021,N_16251,N_16704);
nand U17022 (N_17022,N_16662,N_16521);
and U17023 (N_17023,N_16107,N_16894);
and U17024 (N_17024,N_16314,N_16766);
xnor U17025 (N_17025,N_16453,N_16473);
nor U17026 (N_17026,N_16312,N_16554);
or U17027 (N_17027,N_16613,N_16809);
nand U17028 (N_17028,N_16278,N_16745);
and U17029 (N_17029,N_16185,N_16364);
or U17030 (N_17030,N_16850,N_16290);
nand U17031 (N_17031,N_16504,N_16142);
and U17032 (N_17032,N_16403,N_16248);
nor U17033 (N_17033,N_16942,N_16702);
xnor U17034 (N_17034,N_16874,N_16088);
or U17035 (N_17035,N_16619,N_16741);
nor U17036 (N_17036,N_16992,N_16904);
nor U17037 (N_17037,N_16563,N_16176);
or U17038 (N_17038,N_16359,N_16285);
or U17039 (N_17039,N_16082,N_16535);
xor U17040 (N_17040,N_16186,N_16391);
nand U17041 (N_17041,N_16500,N_16437);
xor U17042 (N_17042,N_16581,N_16887);
or U17043 (N_17043,N_16468,N_16471);
and U17044 (N_17044,N_16306,N_16332);
nand U17045 (N_17045,N_16262,N_16148);
nand U17046 (N_17046,N_16716,N_16028);
xnor U17047 (N_17047,N_16608,N_16384);
nor U17048 (N_17048,N_16656,N_16197);
nor U17049 (N_17049,N_16970,N_16641);
xor U17050 (N_17050,N_16639,N_16812);
nor U17051 (N_17051,N_16164,N_16646);
and U17052 (N_17052,N_16114,N_16177);
and U17053 (N_17053,N_16549,N_16099);
nand U17054 (N_17054,N_16979,N_16456);
nand U17055 (N_17055,N_16091,N_16634);
nor U17056 (N_17056,N_16936,N_16924);
and U17057 (N_17057,N_16275,N_16053);
xnor U17058 (N_17058,N_16517,N_16246);
nor U17059 (N_17059,N_16018,N_16096);
nor U17060 (N_17060,N_16415,N_16873);
xor U17061 (N_17061,N_16982,N_16024);
and U17062 (N_17062,N_16112,N_16543);
nor U17063 (N_17063,N_16727,N_16329);
nand U17064 (N_17064,N_16862,N_16980);
xnor U17065 (N_17065,N_16577,N_16014);
nor U17066 (N_17066,N_16932,N_16733);
and U17067 (N_17067,N_16732,N_16371);
nor U17068 (N_17068,N_16801,N_16782);
and U17069 (N_17069,N_16792,N_16145);
nor U17070 (N_17070,N_16796,N_16911);
and U17071 (N_17071,N_16304,N_16965);
nor U17072 (N_17072,N_16358,N_16692);
nand U17073 (N_17073,N_16455,N_16695);
or U17074 (N_17074,N_16751,N_16627);
and U17075 (N_17075,N_16070,N_16218);
xor U17076 (N_17076,N_16914,N_16986);
nand U17077 (N_17077,N_16405,N_16419);
nand U17078 (N_17078,N_16859,N_16445);
nor U17079 (N_17079,N_16896,N_16508);
or U17080 (N_17080,N_16241,N_16638);
xnor U17081 (N_17081,N_16677,N_16921);
xnor U17082 (N_17082,N_16159,N_16220);
nor U17083 (N_17083,N_16253,N_16795);
xnor U17084 (N_17084,N_16893,N_16509);
and U17085 (N_17085,N_16073,N_16211);
nor U17086 (N_17086,N_16085,N_16075);
xor U17087 (N_17087,N_16589,N_16518);
nand U17088 (N_17088,N_16196,N_16780);
nand U17089 (N_17089,N_16360,N_16151);
nor U17090 (N_17090,N_16660,N_16827);
nand U17091 (N_17091,N_16217,N_16595);
nand U17092 (N_17092,N_16322,N_16341);
nand U17093 (N_17093,N_16038,N_16738);
nand U17094 (N_17094,N_16644,N_16268);
and U17095 (N_17095,N_16394,N_16943);
or U17096 (N_17096,N_16486,N_16976);
xor U17097 (N_17097,N_16072,N_16212);
or U17098 (N_17098,N_16567,N_16906);
nand U17099 (N_17099,N_16269,N_16342);
and U17100 (N_17100,N_16353,N_16242);
xor U17101 (N_17101,N_16006,N_16436);
and U17102 (N_17102,N_16205,N_16841);
or U17103 (N_17103,N_16956,N_16866);
xnor U17104 (N_17104,N_16614,N_16691);
nand U17105 (N_17105,N_16407,N_16654);
or U17106 (N_17106,N_16389,N_16422);
or U17107 (N_17107,N_16195,N_16811);
xnor U17108 (N_17108,N_16883,N_16513);
or U17109 (N_17109,N_16915,N_16477);
nand U17110 (N_17110,N_16502,N_16356);
nand U17111 (N_17111,N_16446,N_16640);
nand U17112 (N_17112,N_16750,N_16266);
xor U17113 (N_17113,N_16687,N_16372);
nand U17114 (N_17114,N_16206,N_16908);
or U17115 (N_17115,N_16566,N_16267);
nand U17116 (N_17116,N_16669,N_16167);
nand U17117 (N_17117,N_16201,N_16032);
nor U17118 (N_17118,N_16519,N_16568);
nand U17119 (N_17119,N_16190,N_16770);
nand U17120 (N_17120,N_16319,N_16607);
or U17121 (N_17121,N_16447,N_16296);
or U17122 (N_17122,N_16802,N_16001);
nor U17123 (N_17123,N_16544,N_16532);
nand U17124 (N_17124,N_16785,N_16065);
or U17125 (N_17125,N_16487,N_16665);
nor U17126 (N_17126,N_16111,N_16818);
or U17127 (N_17127,N_16536,N_16622);
nor U17128 (N_17128,N_16842,N_16821);
nor U17129 (N_17129,N_16993,N_16127);
and U17130 (N_17130,N_16124,N_16819);
nand U17131 (N_17131,N_16408,N_16240);
or U17132 (N_17132,N_16971,N_16012);
and U17133 (N_17133,N_16840,N_16664);
xor U17134 (N_17134,N_16865,N_16347);
xor U17135 (N_17135,N_16410,N_16263);
or U17136 (N_17136,N_16128,N_16081);
or U17137 (N_17137,N_16880,N_16706);
nand U17138 (N_17138,N_16760,N_16666);
nor U17139 (N_17139,N_16828,N_16907);
nor U17140 (N_17140,N_16889,N_16039);
xor U17141 (N_17141,N_16063,N_16033);
nand U17142 (N_17142,N_16441,N_16835);
nand U17143 (N_17143,N_16917,N_16960);
xnor U17144 (N_17144,N_16313,N_16041);
xor U17145 (N_17145,N_16839,N_16433);
xnor U17146 (N_17146,N_16576,N_16175);
and U17147 (N_17147,N_16188,N_16144);
nor U17148 (N_17148,N_16621,N_16854);
xnor U17149 (N_17149,N_16129,N_16141);
xor U17150 (N_17150,N_16042,N_16130);
nor U17151 (N_17151,N_16606,N_16946);
xor U17152 (N_17152,N_16310,N_16478);
xnor U17153 (N_17153,N_16352,N_16138);
and U17154 (N_17154,N_16071,N_16737);
xor U17155 (N_17155,N_16569,N_16222);
xor U17156 (N_17156,N_16857,N_16121);
xor U17157 (N_17157,N_16705,N_16119);
or U17158 (N_17158,N_16474,N_16095);
or U17159 (N_17159,N_16564,N_16414);
or U17160 (N_17160,N_16916,N_16385);
and U17161 (N_17161,N_16459,N_16600);
nor U17162 (N_17162,N_16155,N_16100);
nor U17163 (N_17163,N_16962,N_16772);
xor U17164 (N_17164,N_16747,N_16400);
or U17165 (N_17165,N_16531,N_16254);
xnor U17166 (N_17166,N_16542,N_16224);
and U17167 (N_17167,N_16602,N_16259);
nand U17168 (N_17168,N_16899,N_16448);
and U17169 (N_17169,N_16061,N_16113);
and U17170 (N_17170,N_16725,N_16689);
xnor U17171 (N_17171,N_16872,N_16470);
nor U17172 (N_17172,N_16901,N_16628);
nand U17173 (N_17173,N_16961,N_16270);
nand U17174 (N_17174,N_16324,N_16878);
xor U17175 (N_17175,N_16788,N_16787);
nor U17176 (N_17176,N_16632,N_16629);
nor U17177 (N_17177,N_16199,N_16397);
xor U17178 (N_17178,N_16328,N_16699);
nand U17179 (N_17179,N_16147,N_16925);
nand U17180 (N_17180,N_16580,N_16588);
or U17181 (N_17181,N_16590,N_16786);
nor U17182 (N_17182,N_16680,N_16803);
or U17183 (N_17183,N_16316,N_16236);
nor U17184 (N_17184,N_16713,N_16340);
nand U17185 (N_17185,N_16777,N_16046);
nor U17186 (N_17186,N_16090,N_16714);
xnor U17187 (N_17187,N_16069,N_16514);
xor U17188 (N_17188,N_16635,N_16800);
nor U17189 (N_17189,N_16981,N_16198);
nor U17190 (N_17190,N_16528,N_16510);
and U17191 (N_17191,N_16829,N_16948);
and U17192 (N_17192,N_16748,N_16152);
nor U17193 (N_17193,N_16977,N_16243);
or U17194 (N_17194,N_16898,N_16912);
and U17195 (N_17195,N_16848,N_16905);
nor U17196 (N_17196,N_16623,N_16781);
and U17197 (N_17197,N_16552,N_16420);
xnor U17198 (N_17198,N_16031,N_16661);
nand U17199 (N_17199,N_16845,N_16048);
and U17200 (N_17200,N_16430,N_16833);
or U17201 (N_17201,N_16375,N_16374);
or U17202 (N_17202,N_16994,N_16663);
xnor U17203 (N_17203,N_16227,N_16672);
or U17204 (N_17204,N_16931,N_16999);
nor U17205 (N_17205,N_16276,N_16363);
xnor U17206 (N_17206,N_16007,N_16890);
and U17207 (N_17207,N_16902,N_16945);
nand U17208 (N_17208,N_16463,N_16444);
nand U17209 (N_17209,N_16626,N_16710);
xor U17210 (N_17210,N_16655,N_16527);
nand U17211 (N_17211,N_16529,N_16192);
nor U17212 (N_17212,N_16200,N_16434);
and U17213 (N_17213,N_16438,N_16413);
and U17214 (N_17214,N_16280,N_16219);
nand U17215 (N_17215,N_16271,N_16029);
nor U17216 (N_17216,N_16068,N_16283);
nand U17217 (N_17217,N_16616,N_16743);
and U17218 (N_17218,N_16362,N_16411);
nor U17219 (N_17219,N_16941,N_16055);
nand U17220 (N_17220,N_16491,N_16618);
nor U17221 (N_17221,N_16861,N_16017);
nor U17222 (N_17222,N_16126,N_16368);
nand U17223 (N_17223,N_16076,N_16490);
nand U17224 (N_17224,N_16084,N_16256);
nand U17225 (N_17225,N_16900,N_16011);
nand U17226 (N_17226,N_16265,N_16670);
xnor U17227 (N_17227,N_16944,N_16284);
xnor U17228 (N_17228,N_16277,N_16550);
or U17229 (N_17229,N_16746,N_16435);
xor U17230 (N_17230,N_16493,N_16382);
and U17231 (N_17231,N_16798,N_16035);
xnor U17232 (N_17232,N_16831,N_16707);
and U17233 (N_17233,N_16189,N_16668);
or U17234 (N_17234,N_16150,N_16272);
nand U17235 (N_17235,N_16309,N_16547);
or U17236 (N_17236,N_16282,N_16257);
xor U17237 (N_17237,N_16708,N_16876);
and U17238 (N_17238,N_16557,N_16273);
xor U17239 (N_17239,N_16043,N_16334);
nor U17240 (N_17240,N_16625,N_16735);
nor U17241 (N_17241,N_16213,N_16136);
or U17242 (N_17242,N_16074,N_16494);
xor U17243 (N_17243,N_16230,N_16123);
nor U17244 (N_17244,N_16860,N_16884);
and U17245 (N_17245,N_16671,N_16891);
and U17246 (N_17246,N_16754,N_16496);
xor U17247 (N_17247,N_16958,N_16424);
or U17248 (N_17248,N_16003,N_16953);
and U17249 (N_17249,N_16933,N_16013);
or U17250 (N_17250,N_16631,N_16879);
nor U17251 (N_17251,N_16331,N_16548);
nor U17252 (N_17252,N_16909,N_16178);
xnor U17253 (N_17253,N_16228,N_16797);
nor U17254 (N_17254,N_16815,N_16758);
and U17255 (N_17255,N_16968,N_16886);
nor U17256 (N_17256,N_16822,N_16005);
and U17257 (N_17257,N_16367,N_16034);
xor U17258 (N_17258,N_16657,N_16810);
xnor U17259 (N_17259,N_16120,N_16852);
nor U17260 (N_17260,N_16469,N_16297);
and U17261 (N_17261,N_16252,N_16103);
and U17262 (N_17262,N_16794,N_16700);
and U17263 (N_17263,N_16867,N_16534);
xor U17264 (N_17264,N_16172,N_16685);
xnor U17265 (N_17265,N_16805,N_16472);
or U17266 (N_17266,N_16643,N_16769);
or U17267 (N_17267,N_16843,N_16022);
and U17268 (N_17268,N_16651,N_16421);
xor U17269 (N_17269,N_16134,N_16044);
nor U17270 (N_17270,N_16816,N_16281);
or U17271 (N_17271,N_16615,N_16369);
or U17272 (N_17272,N_16578,N_16877);
and U17273 (N_17273,N_16895,N_16963);
xnor U17274 (N_17274,N_16255,N_16882);
and U17275 (N_17275,N_16573,N_16855);
nor U17276 (N_17276,N_16723,N_16985);
xor U17277 (N_17277,N_16778,N_16765);
or U17278 (N_17278,N_16395,N_16067);
nor U17279 (N_17279,N_16160,N_16337);
nand U17280 (N_17280,N_16318,N_16383);
xnor U17281 (N_17281,N_16881,N_16182);
or U17282 (N_17282,N_16168,N_16681);
nand U17283 (N_17283,N_16279,N_16926);
nor U17284 (N_17284,N_16066,N_16972);
or U17285 (N_17285,N_16133,N_16009);
xor U17286 (N_17286,N_16561,N_16783);
xnor U17287 (N_17287,N_16378,N_16658);
nor U17288 (N_17288,N_16729,N_16401);
xor U17289 (N_17289,N_16101,N_16673);
xnor U17290 (N_17290,N_16237,N_16344);
xor U17291 (N_17291,N_16753,N_16249);
nor U17292 (N_17292,N_16719,N_16667);
or U17293 (N_17293,N_16637,N_16338);
or U17294 (N_17294,N_16058,N_16820);
or U17295 (N_17295,N_16495,N_16806);
nand U17296 (N_17296,N_16132,N_16412);
and U17297 (N_17297,N_16098,N_16711);
and U17298 (N_17298,N_16298,N_16215);
and U17299 (N_17299,N_16291,N_16975);
nand U17300 (N_17300,N_16439,N_16423);
nand U17301 (N_17301,N_16326,N_16019);
nand U17302 (N_17302,N_16935,N_16973);
nand U17303 (N_17303,N_16116,N_16678);
nand U17304 (N_17304,N_16193,N_16336);
xnor U17305 (N_17305,N_16349,N_16836);
or U17306 (N_17306,N_16235,N_16489);
xnor U17307 (N_17307,N_16330,N_16807);
or U17308 (N_17308,N_16226,N_16610);
and U17309 (N_17309,N_16484,N_16396);
xor U17310 (N_17310,N_16021,N_16450);
and U17311 (N_17311,N_16457,N_16432);
nor U17312 (N_17312,N_16166,N_16194);
nand U17313 (N_17313,N_16604,N_16579);
nor U17314 (N_17314,N_16560,N_16292);
and U17315 (N_17315,N_16062,N_16156);
and U17316 (N_17316,N_16722,N_16593);
and U17317 (N_17317,N_16191,N_16030);
or U17318 (N_17318,N_16863,N_16749);
nand U17319 (N_17319,N_16955,N_16715);
nor U17320 (N_17320,N_16790,N_16229);
nand U17321 (N_17321,N_16539,N_16208);
xor U17322 (N_17322,N_16516,N_16357);
or U17323 (N_17323,N_16599,N_16892);
xnor U17324 (N_17324,N_16454,N_16814);
nand U17325 (N_17325,N_16442,N_16609);
nand U17326 (N_17326,N_16026,N_16203);
nand U17327 (N_17327,N_16938,N_16726);
or U17328 (N_17328,N_16511,N_16995);
or U17329 (N_17329,N_16799,N_16497);
or U17330 (N_17330,N_16335,N_16617);
nor U17331 (N_17331,N_16157,N_16016);
nand U17332 (N_17332,N_16245,N_16117);
or U17333 (N_17333,N_16688,N_16761);
xnor U17334 (N_17334,N_16937,N_16102);
nand U17335 (N_17335,N_16402,N_16086);
nand U17336 (N_17336,N_16169,N_16135);
and U17337 (N_17337,N_16969,N_16443);
nor U17338 (N_17338,N_16339,N_16078);
and U17339 (N_17339,N_16730,N_16274);
nand U17340 (N_17340,N_16393,N_16988);
and U17341 (N_17341,N_16143,N_16565);
and U17342 (N_17342,N_16682,N_16387);
nand U17343 (N_17343,N_16174,N_16718);
nand U17344 (N_17344,N_16139,N_16051);
nor U17345 (N_17345,N_16659,N_16106);
and U17346 (N_17346,N_16216,N_16922);
xnor U17347 (N_17347,N_16574,N_16376);
nor U17348 (N_17348,N_16301,N_16507);
xor U17349 (N_17349,N_16964,N_16940);
xnor U17350 (N_17350,N_16348,N_16020);
and U17351 (N_17351,N_16923,N_16776);
or U17352 (N_17352,N_16693,N_16556);
and U17353 (N_17353,N_16343,N_16302);
nand U17354 (N_17354,N_16506,N_16239);
nor U17355 (N_17355,N_16601,N_16325);
xnor U17356 (N_17356,N_16110,N_16054);
nor U17357 (N_17357,N_16427,N_16675);
and U17358 (N_17358,N_16137,N_16771);
and U17359 (N_17359,N_16004,N_16181);
or U17360 (N_17360,N_16286,N_16250);
nand U17361 (N_17361,N_16258,N_16720);
nor U17362 (N_17362,N_16361,N_16104);
or U17363 (N_17363,N_16077,N_16027);
or U17364 (N_17364,N_16991,N_16630);
xor U17365 (N_17365,N_16449,N_16856);
or U17366 (N_17366,N_16538,N_16537);
xnor U17367 (N_17367,N_16575,N_16824);
and U17368 (N_17368,N_16755,N_16851);
or U17369 (N_17369,N_16162,N_16083);
and U17370 (N_17370,N_16703,N_16826);
nand U17371 (N_17371,N_16624,N_16300);
nand U17372 (N_17372,N_16684,N_16460);
xnor U17373 (N_17373,N_16927,N_16585);
xor U17374 (N_17374,N_16739,N_16097);
and U17375 (N_17375,N_16023,N_16392);
xor U17376 (N_17376,N_16813,N_16959);
nor U17377 (N_17377,N_16288,N_16503);
or U17378 (N_17378,N_16903,N_16154);
nand U17379 (N_17379,N_16910,N_16161);
nor U17380 (N_17380,N_16499,N_16440);
nand U17381 (N_17381,N_16417,N_16920);
or U17382 (N_17382,N_16858,N_16089);
nor U17383 (N_17383,N_16731,N_16323);
xor U17384 (N_17384,N_16744,N_16398);
nand U17385 (N_17385,N_16210,N_16308);
and U17386 (N_17386,N_16429,N_16752);
and U17387 (N_17387,N_16592,N_16462);
or U17388 (N_17388,N_16520,N_16642);
nand U17389 (N_17389,N_16173,N_16501);
nor U17390 (N_17390,N_16817,N_16888);
and U17391 (N_17391,N_16793,N_16939);
or U17392 (N_17392,N_16679,N_16997);
or U17393 (N_17393,N_16052,N_16379);
nor U17394 (N_17394,N_16333,N_16591);
nor U17395 (N_17395,N_16223,N_16146);
nor U17396 (N_17396,N_16849,N_16153);
or U17397 (N_17397,N_16844,N_16571);
or U17398 (N_17398,N_16530,N_16853);
xnor U17399 (N_17399,N_16303,N_16315);
nor U17400 (N_17400,N_16612,N_16870);
xor U17401 (N_17401,N_16000,N_16015);
nor U17402 (N_17402,N_16428,N_16149);
or U17403 (N_17403,N_16060,N_16525);
and U17404 (N_17404,N_16633,N_16476);
or U17405 (N_17405,N_16523,N_16649);
or U17406 (N_17406,N_16837,N_16698);
nand U17407 (N_17407,N_16380,N_16774);
or U17408 (N_17408,N_16481,N_16094);
nand U17409 (N_17409,N_16214,N_16759);
nand U17410 (N_17410,N_16307,N_16049);
nand U17411 (N_17411,N_16010,N_16987);
nor U17412 (N_17412,N_16057,N_16466);
nor U17413 (N_17413,N_16791,N_16885);
or U17414 (N_17414,N_16559,N_16390);
xor U17415 (N_17415,N_16540,N_16533);
nor U17416 (N_17416,N_16724,N_16238);
nor U17417 (N_17417,N_16763,N_16370);
nand U17418 (N_17418,N_16648,N_16779);
or U17419 (N_17419,N_16694,N_16808);
nand U17420 (N_17420,N_16690,N_16426);
nor U17421 (N_17421,N_16406,N_16990);
nor U17422 (N_17422,N_16354,N_16122);
xor U17423 (N_17423,N_16697,N_16871);
nand U17424 (N_17424,N_16846,N_16645);
nand U17425 (N_17425,N_16289,N_16409);
xor U17426 (N_17426,N_16366,N_16947);
or U17427 (N_17427,N_16140,N_16287);
and U17428 (N_17428,N_16452,N_16951);
nand U17429 (N_17429,N_16934,N_16056);
and U17430 (N_17430,N_16294,N_16570);
and U17431 (N_17431,N_16431,N_16350);
nand U17432 (N_17432,N_16605,N_16170);
nand U17433 (N_17433,N_16327,N_16653);
nand U17434 (N_17434,N_16603,N_16949);
xnor U17435 (N_17435,N_16582,N_16505);
nor U17436 (N_17436,N_16377,N_16583);
or U17437 (N_17437,N_16311,N_16721);
xor U17438 (N_17438,N_16465,N_16475);
and U17439 (N_17439,N_16996,N_16701);
xor U17440 (N_17440,N_16930,N_16696);
nor U17441 (N_17441,N_16897,N_16321);
and U17442 (N_17442,N_16524,N_16847);
nor U17443 (N_17443,N_16868,N_16451);
nand U17444 (N_17444,N_16404,N_16584);
and U17445 (N_17445,N_16260,N_16966);
or U17446 (N_17446,N_16998,N_16187);
nor U17447 (N_17447,N_16918,N_16418);
nand U17448 (N_17448,N_16728,N_16586);
nand U17449 (N_17449,N_16416,N_16184);
xnor U17450 (N_17450,N_16983,N_16105);
nor U17451 (N_17451,N_16115,N_16740);
nand U17452 (N_17452,N_16989,N_16087);
nor U17453 (N_17453,N_16919,N_16221);
xnor U17454 (N_17454,N_16036,N_16183);
nand U17455 (N_17455,N_16636,N_16825);
and U17456 (N_17456,N_16293,N_16717);
xnor U17457 (N_17457,N_16025,N_16231);
nand U17458 (N_17458,N_16950,N_16674);
and U17459 (N_17459,N_16974,N_16597);
nor U17460 (N_17460,N_16546,N_16830);
nand U17461 (N_17461,N_16388,N_16734);
and U17462 (N_17462,N_16515,N_16092);
xor U17463 (N_17463,N_16482,N_16775);
nor U17464 (N_17464,N_16686,N_16742);
nor U17465 (N_17465,N_16002,N_16399);
xnor U17466 (N_17466,N_16709,N_16118);
nand U17467 (N_17467,N_16558,N_16040);
or U17468 (N_17468,N_16929,N_16045);
nor U17469 (N_17469,N_16180,N_16108);
nor U17470 (N_17470,N_16261,N_16984);
and U17471 (N_17471,N_16611,N_16480);
nor U17472 (N_17472,N_16676,N_16620);
or U17473 (N_17473,N_16204,N_16131);
nand U17474 (N_17474,N_16789,N_16553);
or U17475 (N_17475,N_16522,N_16832);
and U17476 (N_17476,N_16488,N_16594);
nand U17477 (N_17477,N_16712,N_16264);
or U17478 (N_17478,N_16207,N_16784);
nor U17479 (N_17479,N_16305,N_16179);
nor U17480 (N_17480,N_16498,N_16050);
xor U17481 (N_17481,N_16978,N_16952);
or U17482 (N_17482,N_16479,N_16736);
nand U17483 (N_17483,N_16598,N_16165);
or U17484 (N_17484,N_16346,N_16875);
nand U17485 (N_17485,N_16386,N_16461);
nor U17486 (N_17486,N_16562,N_16345);
xor U17487 (N_17487,N_16320,N_16093);
or U17488 (N_17488,N_16757,N_16954);
nor U17489 (N_17489,N_16233,N_16351);
or U17490 (N_17490,N_16163,N_16317);
nor U17491 (N_17491,N_16541,N_16647);
and U17492 (N_17492,N_16079,N_16957);
and U17493 (N_17493,N_16171,N_16109);
xnor U17494 (N_17494,N_16683,N_16381);
nor U17495 (N_17495,N_16526,N_16804);
nor U17496 (N_17496,N_16928,N_16008);
nand U17497 (N_17497,N_16425,N_16596);
and U17498 (N_17498,N_16467,N_16967);
or U17499 (N_17499,N_16512,N_16551);
and U17500 (N_17500,N_16961,N_16788);
xor U17501 (N_17501,N_16066,N_16352);
nand U17502 (N_17502,N_16106,N_16257);
and U17503 (N_17503,N_16872,N_16893);
or U17504 (N_17504,N_16564,N_16112);
or U17505 (N_17505,N_16919,N_16971);
xnor U17506 (N_17506,N_16353,N_16024);
xor U17507 (N_17507,N_16814,N_16999);
nor U17508 (N_17508,N_16228,N_16446);
or U17509 (N_17509,N_16029,N_16704);
or U17510 (N_17510,N_16203,N_16837);
nand U17511 (N_17511,N_16505,N_16390);
nor U17512 (N_17512,N_16794,N_16990);
nor U17513 (N_17513,N_16904,N_16235);
nand U17514 (N_17514,N_16435,N_16960);
and U17515 (N_17515,N_16734,N_16357);
or U17516 (N_17516,N_16777,N_16768);
nand U17517 (N_17517,N_16375,N_16322);
or U17518 (N_17518,N_16810,N_16835);
nor U17519 (N_17519,N_16879,N_16097);
xor U17520 (N_17520,N_16871,N_16207);
nand U17521 (N_17521,N_16776,N_16231);
or U17522 (N_17522,N_16907,N_16821);
nand U17523 (N_17523,N_16988,N_16846);
and U17524 (N_17524,N_16899,N_16920);
and U17525 (N_17525,N_16753,N_16212);
nand U17526 (N_17526,N_16616,N_16300);
nand U17527 (N_17527,N_16611,N_16188);
or U17528 (N_17528,N_16098,N_16921);
nand U17529 (N_17529,N_16143,N_16219);
or U17530 (N_17530,N_16322,N_16335);
nor U17531 (N_17531,N_16267,N_16382);
nand U17532 (N_17532,N_16881,N_16628);
and U17533 (N_17533,N_16641,N_16145);
or U17534 (N_17534,N_16608,N_16766);
nand U17535 (N_17535,N_16632,N_16377);
or U17536 (N_17536,N_16703,N_16504);
and U17537 (N_17537,N_16110,N_16361);
nand U17538 (N_17538,N_16477,N_16001);
nor U17539 (N_17539,N_16660,N_16017);
or U17540 (N_17540,N_16130,N_16421);
or U17541 (N_17541,N_16025,N_16147);
xnor U17542 (N_17542,N_16789,N_16491);
nor U17543 (N_17543,N_16827,N_16831);
nand U17544 (N_17544,N_16232,N_16674);
xor U17545 (N_17545,N_16178,N_16029);
xnor U17546 (N_17546,N_16826,N_16742);
nor U17547 (N_17547,N_16994,N_16803);
xor U17548 (N_17548,N_16633,N_16674);
or U17549 (N_17549,N_16674,N_16494);
xnor U17550 (N_17550,N_16442,N_16196);
xor U17551 (N_17551,N_16424,N_16516);
nand U17552 (N_17552,N_16651,N_16732);
xnor U17553 (N_17553,N_16871,N_16773);
or U17554 (N_17554,N_16823,N_16030);
and U17555 (N_17555,N_16209,N_16235);
nand U17556 (N_17556,N_16140,N_16620);
xnor U17557 (N_17557,N_16279,N_16562);
nand U17558 (N_17558,N_16054,N_16349);
and U17559 (N_17559,N_16533,N_16899);
nand U17560 (N_17560,N_16850,N_16400);
xor U17561 (N_17561,N_16138,N_16128);
nand U17562 (N_17562,N_16080,N_16349);
or U17563 (N_17563,N_16821,N_16578);
nand U17564 (N_17564,N_16619,N_16277);
xor U17565 (N_17565,N_16370,N_16902);
xnor U17566 (N_17566,N_16527,N_16793);
or U17567 (N_17567,N_16462,N_16759);
nand U17568 (N_17568,N_16147,N_16238);
nor U17569 (N_17569,N_16525,N_16621);
and U17570 (N_17570,N_16436,N_16227);
or U17571 (N_17571,N_16928,N_16888);
and U17572 (N_17572,N_16074,N_16042);
and U17573 (N_17573,N_16551,N_16187);
or U17574 (N_17574,N_16196,N_16757);
and U17575 (N_17575,N_16795,N_16284);
nor U17576 (N_17576,N_16731,N_16928);
nor U17577 (N_17577,N_16917,N_16056);
nor U17578 (N_17578,N_16663,N_16149);
or U17579 (N_17579,N_16056,N_16189);
xor U17580 (N_17580,N_16457,N_16865);
nand U17581 (N_17581,N_16601,N_16026);
nand U17582 (N_17582,N_16842,N_16615);
nand U17583 (N_17583,N_16276,N_16597);
nor U17584 (N_17584,N_16738,N_16378);
xor U17585 (N_17585,N_16069,N_16138);
nor U17586 (N_17586,N_16485,N_16564);
xnor U17587 (N_17587,N_16682,N_16539);
and U17588 (N_17588,N_16840,N_16335);
nor U17589 (N_17589,N_16486,N_16015);
nor U17590 (N_17590,N_16925,N_16798);
nor U17591 (N_17591,N_16270,N_16664);
nor U17592 (N_17592,N_16607,N_16851);
and U17593 (N_17593,N_16998,N_16455);
or U17594 (N_17594,N_16272,N_16436);
xor U17595 (N_17595,N_16682,N_16103);
nand U17596 (N_17596,N_16421,N_16423);
nand U17597 (N_17597,N_16787,N_16511);
xor U17598 (N_17598,N_16876,N_16378);
or U17599 (N_17599,N_16060,N_16988);
nor U17600 (N_17600,N_16410,N_16512);
nand U17601 (N_17601,N_16659,N_16006);
xor U17602 (N_17602,N_16453,N_16008);
and U17603 (N_17603,N_16456,N_16900);
nor U17604 (N_17604,N_16155,N_16998);
or U17605 (N_17605,N_16246,N_16296);
xor U17606 (N_17606,N_16830,N_16960);
or U17607 (N_17607,N_16555,N_16574);
and U17608 (N_17608,N_16577,N_16451);
xnor U17609 (N_17609,N_16322,N_16516);
or U17610 (N_17610,N_16122,N_16538);
and U17611 (N_17611,N_16210,N_16868);
xnor U17612 (N_17612,N_16004,N_16339);
nand U17613 (N_17613,N_16860,N_16049);
and U17614 (N_17614,N_16946,N_16257);
nor U17615 (N_17615,N_16925,N_16636);
nor U17616 (N_17616,N_16647,N_16380);
nand U17617 (N_17617,N_16592,N_16020);
nand U17618 (N_17618,N_16342,N_16475);
and U17619 (N_17619,N_16105,N_16110);
nand U17620 (N_17620,N_16762,N_16598);
xor U17621 (N_17621,N_16772,N_16332);
or U17622 (N_17622,N_16683,N_16767);
nor U17623 (N_17623,N_16840,N_16220);
and U17624 (N_17624,N_16337,N_16262);
nand U17625 (N_17625,N_16770,N_16103);
and U17626 (N_17626,N_16745,N_16934);
nor U17627 (N_17627,N_16443,N_16820);
or U17628 (N_17628,N_16668,N_16663);
xor U17629 (N_17629,N_16263,N_16646);
nor U17630 (N_17630,N_16425,N_16627);
or U17631 (N_17631,N_16169,N_16487);
and U17632 (N_17632,N_16041,N_16609);
nor U17633 (N_17633,N_16366,N_16620);
xnor U17634 (N_17634,N_16641,N_16191);
and U17635 (N_17635,N_16412,N_16081);
nand U17636 (N_17636,N_16344,N_16055);
or U17637 (N_17637,N_16245,N_16233);
xnor U17638 (N_17638,N_16510,N_16215);
nor U17639 (N_17639,N_16942,N_16423);
nand U17640 (N_17640,N_16198,N_16727);
or U17641 (N_17641,N_16268,N_16545);
or U17642 (N_17642,N_16136,N_16636);
or U17643 (N_17643,N_16395,N_16794);
nand U17644 (N_17644,N_16795,N_16370);
and U17645 (N_17645,N_16360,N_16065);
and U17646 (N_17646,N_16309,N_16399);
and U17647 (N_17647,N_16331,N_16281);
and U17648 (N_17648,N_16327,N_16388);
and U17649 (N_17649,N_16684,N_16580);
xnor U17650 (N_17650,N_16490,N_16064);
or U17651 (N_17651,N_16253,N_16851);
or U17652 (N_17652,N_16337,N_16408);
and U17653 (N_17653,N_16478,N_16353);
xor U17654 (N_17654,N_16807,N_16356);
nand U17655 (N_17655,N_16631,N_16120);
and U17656 (N_17656,N_16640,N_16438);
xnor U17657 (N_17657,N_16335,N_16529);
nand U17658 (N_17658,N_16611,N_16893);
nor U17659 (N_17659,N_16749,N_16358);
and U17660 (N_17660,N_16711,N_16320);
nor U17661 (N_17661,N_16291,N_16054);
xor U17662 (N_17662,N_16034,N_16626);
nor U17663 (N_17663,N_16972,N_16853);
nand U17664 (N_17664,N_16969,N_16341);
and U17665 (N_17665,N_16772,N_16632);
or U17666 (N_17666,N_16960,N_16931);
or U17667 (N_17667,N_16383,N_16775);
and U17668 (N_17668,N_16232,N_16599);
nand U17669 (N_17669,N_16394,N_16048);
nand U17670 (N_17670,N_16363,N_16290);
nand U17671 (N_17671,N_16485,N_16858);
nand U17672 (N_17672,N_16158,N_16102);
and U17673 (N_17673,N_16773,N_16078);
nand U17674 (N_17674,N_16452,N_16475);
xor U17675 (N_17675,N_16822,N_16658);
and U17676 (N_17676,N_16756,N_16743);
nand U17677 (N_17677,N_16713,N_16926);
or U17678 (N_17678,N_16455,N_16473);
nor U17679 (N_17679,N_16924,N_16729);
or U17680 (N_17680,N_16554,N_16185);
nand U17681 (N_17681,N_16436,N_16171);
xnor U17682 (N_17682,N_16487,N_16591);
nand U17683 (N_17683,N_16711,N_16926);
nor U17684 (N_17684,N_16788,N_16326);
nand U17685 (N_17685,N_16115,N_16355);
and U17686 (N_17686,N_16332,N_16815);
nor U17687 (N_17687,N_16865,N_16906);
nor U17688 (N_17688,N_16833,N_16121);
nor U17689 (N_17689,N_16071,N_16651);
nand U17690 (N_17690,N_16086,N_16414);
and U17691 (N_17691,N_16828,N_16052);
nand U17692 (N_17692,N_16516,N_16954);
nand U17693 (N_17693,N_16865,N_16120);
xnor U17694 (N_17694,N_16043,N_16784);
nand U17695 (N_17695,N_16291,N_16855);
and U17696 (N_17696,N_16824,N_16172);
and U17697 (N_17697,N_16216,N_16946);
and U17698 (N_17698,N_16151,N_16330);
xnor U17699 (N_17699,N_16877,N_16002);
and U17700 (N_17700,N_16826,N_16265);
nor U17701 (N_17701,N_16003,N_16134);
xor U17702 (N_17702,N_16987,N_16013);
nand U17703 (N_17703,N_16053,N_16701);
nand U17704 (N_17704,N_16314,N_16628);
or U17705 (N_17705,N_16988,N_16733);
nand U17706 (N_17706,N_16315,N_16565);
and U17707 (N_17707,N_16471,N_16977);
nor U17708 (N_17708,N_16289,N_16990);
nor U17709 (N_17709,N_16778,N_16206);
nand U17710 (N_17710,N_16563,N_16070);
nor U17711 (N_17711,N_16515,N_16309);
or U17712 (N_17712,N_16287,N_16712);
nand U17713 (N_17713,N_16237,N_16646);
nor U17714 (N_17714,N_16052,N_16228);
or U17715 (N_17715,N_16966,N_16303);
or U17716 (N_17716,N_16334,N_16801);
xnor U17717 (N_17717,N_16924,N_16221);
nand U17718 (N_17718,N_16489,N_16212);
nor U17719 (N_17719,N_16350,N_16011);
xnor U17720 (N_17720,N_16635,N_16272);
or U17721 (N_17721,N_16962,N_16010);
nor U17722 (N_17722,N_16316,N_16141);
and U17723 (N_17723,N_16483,N_16746);
nand U17724 (N_17724,N_16924,N_16660);
xor U17725 (N_17725,N_16800,N_16518);
and U17726 (N_17726,N_16268,N_16802);
nor U17727 (N_17727,N_16597,N_16948);
nand U17728 (N_17728,N_16324,N_16197);
xnor U17729 (N_17729,N_16593,N_16060);
or U17730 (N_17730,N_16045,N_16902);
nor U17731 (N_17731,N_16055,N_16461);
nor U17732 (N_17732,N_16406,N_16287);
or U17733 (N_17733,N_16563,N_16832);
and U17734 (N_17734,N_16591,N_16024);
nand U17735 (N_17735,N_16875,N_16084);
nor U17736 (N_17736,N_16616,N_16720);
xnor U17737 (N_17737,N_16898,N_16400);
and U17738 (N_17738,N_16747,N_16328);
or U17739 (N_17739,N_16366,N_16044);
or U17740 (N_17740,N_16262,N_16021);
or U17741 (N_17741,N_16243,N_16716);
nand U17742 (N_17742,N_16309,N_16713);
xnor U17743 (N_17743,N_16781,N_16634);
and U17744 (N_17744,N_16291,N_16927);
or U17745 (N_17745,N_16297,N_16300);
xor U17746 (N_17746,N_16715,N_16636);
nand U17747 (N_17747,N_16549,N_16909);
xor U17748 (N_17748,N_16503,N_16774);
xor U17749 (N_17749,N_16431,N_16394);
and U17750 (N_17750,N_16299,N_16448);
nand U17751 (N_17751,N_16610,N_16867);
nand U17752 (N_17752,N_16894,N_16353);
nor U17753 (N_17753,N_16600,N_16874);
or U17754 (N_17754,N_16480,N_16203);
or U17755 (N_17755,N_16355,N_16459);
xor U17756 (N_17756,N_16318,N_16303);
or U17757 (N_17757,N_16049,N_16238);
nor U17758 (N_17758,N_16075,N_16279);
xor U17759 (N_17759,N_16484,N_16882);
and U17760 (N_17760,N_16966,N_16925);
nand U17761 (N_17761,N_16546,N_16656);
nand U17762 (N_17762,N_16428,N_16266);
and U17763 (N_17763,N_16683,N_16495);
nand U17764 (N_17764,N_16607,N_16763);
nand U17765 (N_17765,N_16543,N_16348);
xor U17766 (N_17766,N_16949,N_16053);
nor U17767 (N_17767,N_16202,N_16866);
or U17768 (N_17768,N_16601,N_16281);
xnor U17769 (N_17769,N_16338,N_16161);
or U17770 (N_17770,N_16119,N_16055);
and U17771 (N_17771,N_16898,N_16730);
xnor U17772 (N_17772,N_16384,N_16431);
and U17773 (N_17773,N_16789,N_16741);
xnor U17774 (N_17774,N_16739,N_16209);
nor U17775 (N_17775,N_16189,N_16395);
or U17776 (N_17776,N_16003,N_16557);
nand U17777 (N_17777,N_16386,N_16365);
or U17778 (N_17778,N_16538,N_16250);
nor U17779 (N_17779,N_16349,N_16492);
xor U17780 (N_17780,N_16249,N_16903);
nand U17781 (N_17781,N_16648,N_16346);
xor U17782 (N_17782,N_16531,N_16338);
and U17783 (N_17783,N_16548,N_16332);
and U17784 (N_17784,N_16672,N_16232);
or U17785 (N_17785,N_16169,N_16123);
nor U17786 (N_17786,N_16349,N_16451);
nor U17787 (N_17787,N_16166,N_16493);
xor U17788 (N_17788,N_16216,N_16211);
or U17789 (N_17789,N_16656,N_16708);
nand U17790 (N_17790,N_16936,N_16971);
nor U17791 (N_17791,N_16913,N_16235);
nor U17792 (N_17792,N_16178,N_16214);
nand U17793 (N_17793,N_16496,N_16917);
and U17794 (N_17794,N_16958,N_16912);
nand U17795 (N_17795,N_16602,N_16446);
nor U17796 (N_17796,N_16774,N_16518);
nor U17797 (N_17797,N_16060,N_16680);
nor U17798 (N_17798,N_16697,N_16576);
nor U17799 (N_17799,N_16334,N_16203);
xnor U17800 (N_17800,N_16334,N_16866);
nor U17801 (N_17801,N_16649,N_16165);
xor U17802 (N_17802,N_16277,N_16098);
nor U17803 (N_17803,N_16408,N_16309);
or U17804 (N_17804,N_16093,N_16756);
xnor U17805 (N_17805,N_16060,N_16362);
nor U17806 (N_17806,N_16654,N_16010);
and U17807 (N_17807,N_16407,N_16887);
xor U17808 (N_17808,N_16111,N_16397);
nor U17809 (N_17809,N_16479,N_16230);
or U17810 (N_17810,N_16254,N_16893);
and U17811 (N_17811,N_16536,N_16998);
or U17812 (N_17812,N_16315,N_16889);
nor U17813 (N_17813,N_16933,N_16590);
nand U17814 (N_17814,N_16428,N_16279);
nor U17815 (N_17815,N_16388,N_16307);
nand U17816 (N_17816,N_16302,N_16298);
nor U17817 (N_17817,N_16711,N_16284);
nor U17818 (N_17818,N_16459,N_16794);
nor U17819 (N_17819,N_16926,N_16795);
nor U17820 (N_17820,N_16230,N_16839);
and U17821 (N_17821,N_16561,N_16456);
xor U17822 (N_17822,N_16169,N_16471);
or U17823 (N_17823,N_16417,N_16024);
nand U17824 (N_17824,N_16267,N_16099);
xnor U17825 (N_17825,N_16206,N_16055);
xnor U17826 (N_17826,N_16114,N_16220);
or U17827 (N_17827,N_16537,N_16508);
nand U17828 (N_17828,N_16747,N_16503);
nor U17829 (N_17829,N_16254,N_16042);
nand U17830 (N_17830,N_16269,N_16564);
xor U17831 (N_17831,N_16473,N_16799);
or U17832 (N_17832,N_16139,N_16641);
nor U17833 (N_17833,N_16895,N_16819);
or U17834 (N_17834,N_16913,N_16857);
xnor U17835 (N_17835,N_16946,N_16516);
nor U17836 (N_17836,N_16119,N_16461);
xor U17837 (N_17837,N_16052,N_16813);
and U17838 (N_17838,N_16364,N_16361);
nor U17839 (N_17839,N_16608,N_16982);
and U17840 (N_17840,N_16788,N_16503);
nand U17841 (N_17841,N_16587,N_16873);
xnor U17842 (N_17842,N_16389,N_16769);
xor U17843 (N_17843,N_16349,N_16901);
xor U17844 (N_17844,N_16213,N_16845);
or U17845 (N_17845,N_16368,N_16036);
or U17846 (N_17846,N_16046,N_16591);
nor U17847 (N_17847,N_16548,N_16239);
nor U17848 (N_17848,N_16771,N_16913);
xor U17849 (N_17849,N_16098,N_16593);
nand U17850 (N_17850,N_16934,N_16145);
nor U17851 (N_17851,N_16711,N_16884);
or U17852 (N_17852,N_16299,N_16802);
xor U17853 (N_17853,N_16738,N_16190);
nand U17854 (N_17854,N_16061,N_16687);
nand U17855 (N_17855,N_16880,N_16302);
or U17856 (N_17856,N_16283,N_16671);
nand U17857 (N_17857,N_16823,N_16765);
or U17858 (N_17858,N_16421,N_16289);
and U17859 (N_17859,N_16341,N_16389);
nor U17860 (N_17860,N_16066,N_16978);
xnor U17861 (N_17861,N_16890,N_16270);
nand U17862 (N_17862,N_16324,N_16537);
nand U17863 (N_17863,N_16838,N_16678);
and U17864 (N_17864,N_16474,N_16231);
xor U17865 (N_17865,N_16616,N_16267);
xor U17866 (N_17866,N_16998,N_16722);
nand U17867 (N_17867,N_16380,N_16991);
nor U17868 (N_17868,N_16498,N_16432);
xor U17869 (N_17869,N_16908,N_16563);
and U17870 (N_17870,N_16231,N_16432);
and U17871 (N_17871,N_16151,N_16204);
xnor U17872 (N_17872,N_16992,N_16401);
nor U17873 (N_17873,N_16723,N_16264);
nand U17874 (N_17874,N_16413,N_16479);
nand U17875 (N_17875,N_16443,N_16627);
and U17876 (N_17876,N_16930,N_16518);
xnor U17877 (N_17877,N_16626,N_16016);
xor U17878 (N_17878,N_16843,N_16059);
and U17879 (N_17879,N_16430,N_16798);
and U17880 (N_17880,N_16899,N_16344);
xnor U17881 (N_17881,N_16265,N_16133);
and U17882 (N_17882,N_16433,N_16904);
xnor U17883 (N_17883,N_16685,N_16863);
nor U17884 (N_17884,N_16638,N_16871);
nor U17885 (N_17885,N_16822,N_16468);
and U17886 (N_17886,N_16175,N_16504);
xnor U17887 (N_17887,N_16807,N_16904);
xnor U17888 (N_17888,N_16318,N_16292);
nor U17889 (N_17889,N_16642,N_16877);
nand U17890 (N_17890,N_16425,N_16590);
or U17891 (N_17891,N_16128,N_16992);
nand U17892 (N_17892,N_16840,N_16876);
nand U17893 (N_17893,N_16428,N_16785);
nor U17894 (N_17894,N_16519,N_16481);
or U17895 (N_17895,N_16112,N_16582);
nor U17896 (N_17896,N_16943,N_16048);
nand U17897 (N_17897,N_16025,N_16259);
nand U17898 (N_17898,N_16800,N_16740);
or U17899 (N_17899,N_16326,N_16266);
nand U17900 (N_17900,N_16264,N_16866);
xnor U17901 (N_17901,N_16067,N_16594);
and U17902 (N_17902,N_16111,N_16628);
nor U17903 (N_17903,N_16875,N_16956);
nand U17904 (N_17904,N_16882,N_16288);
nand U17905 (N_17905,N_16182,N_16004);
and U17906 (N_17906,N_16984,N_16905);
nand U17907 (N_17907,N_16078,N_16724);
and U17908 (N_17908,N_16409,N_16536);
nand U17909 (N_17909,N_16076,N_16279);
and U17910 (N_17910,N_16893,N_16809);
nand U17911 (N_17911,N_16645,N_16152);
nand U17912 (N_17912,N_16163,N_16830);
xor U17913 (N_17913,N_16701,N_16040);
or U17914 (N_17914,N_16310,N_16683);
or U17915 (N_17915,N_16932,N_16257);
xor U17916 (N_17916,N_16454,N_16798);
and U17917 (N_17917,N_16260,N_16519);
nor U17918 (N_17918,N_16890,N_16182);
and U17919 (N_17919,N_16398,N_16125);
xor U17920 (N_17920,N_16932,N_16516);
nor U17921 (N_17921,N_16987,N_16966);
and U17922 (N_17922,N_16958,N_16539);
and U17923 (N_17923,N_16077,N_16128);
nor U17924 (N_17924,N_16309,N_16519);
or U17925 (N_17925,N_16785,N_16978);
and U17926 (N_17926,N_16803,N_16947);
xor U17927 (N_17927,N_16965,N_16916);
nor U17928 (N_17928,N_16476,N_16814);
nor U17929 (N_17929,N_16727,N_16916);
xnor U17930 (N_17930,N_16000,N_16226);
xor U17931 (N_17931,N_16051,N_16457);
xor U17932 (N_17932,N_16950,N_16976);
nand U17933 (N_17933,N_16301,N_16074);
or U17934 (N_17934,N_16046,N_16745);
nor U17935 (N_17935,N_16618,N_16358);
nand U17936 (N_17936,N_16323,N_16054);
nand U17937 (N_17937,N_16115,N_16137);
nand U17938 (N_17938,N_16851,N_16528);
nand U17939 (N_17939,N_16171,N_16671);
xnor U17940 (N_17940,N_16088,N_16627);
nand U17941 (N_17941,N_16960,N_16629);
nand U17942 (N_17942,N_16293,N_16104);
nand U17943 (N_17943,N_16664,N_16141);
nor U17944 (N_17944,N_16957,N_16962);
or U17945 (N_17945,N_16821,N_16510);
or U17946 (N_17946,N_16749,N_16680);
xor U17947 (N_17947,N_16008,N_16933);
nand U17948 (N_17948,N_16643,N_16695);
nor U17949 (N_17949,N_16400,N_16928);
and U17950 (N_17950,N_16640,N_16136);
or U17951 (N_17951,N_16502,N_16005);
and U17952 (N_17952,N_16912,N_16339);
nor U17953 (N_17953,N_16702,N_16156);
or U17954 (N_17954,N_16274,N_16253);
nor U17955 (N_17955,N_16511,N_16975);
nor U17956 (N_17956,N_16769,N_16018);
xor U17957 (N_17957,N_16736,N_16682);
or U17958 (N_17958,N_16501,N_16356);
nor U17959 (N_17959,N_16546,N_16453);
and U17960 (N_17960,N_16910,N_16299);
and U17961 (N_17961,N_16181,N_16054);
and U17962 (N_17962,N_16859,N_16242);
nor U17963 (N_17963,N_16306,N_16189);
nor U17964 (N_17964,N_16518,N_16982);
or U17965 (N_17965,N_16908,N_16121);
nand U17966 (N_17966,N_16646,N_16443);
or U17967 (N_17967,N_16595,N_16633);
or U17968 (N_17968,N_16145,N_16495);
nor U17969 (N_17969,N_16248,N_16412);
nor U17970 (N_17970,N_16250,N_16965);
and U17971 (N_17971,N_16767,N_16319);
nor U17972 (N_17972,N_16979,N_16781);
xnor U17973 (N_17973,N_16688,N_16459);
and U17974 (N_17974,N_16356,N_16919);
and U17975 (N_17975,N_16265,N_16875);
or U17976 (N_17976,N_16544,N_16295);
or U17977 (N_17977,N_16988,N_16658);
xnor U17978 (N_17978,N_16552,N_16737);
or U17979 (N_17979,N_16824,N_16061);
nand U17980 (N_17980,N_16119,N_16116);
nor U17981 (N_17981,N_16819,N_16623);
nor U17982 (N_17982,N_16597,N_16362);
nor U17983 (N_17983,N_16618,N_16353);
nand U17984 (N_17984,N_16725,N_16508);
nand U17985 (N_17985,N_16222,N_16062);
and U17986 (N_17986,N_16632,N_16265);
or U17987 (N_17987,N_16492,N_16721);
nor U17988 (N_17988,N_16594,N_16140);
or U17989 (N_17989,N_16590,N_16179);
or U17990 (N_17990,N_16246,N_16267);
nand U17991 (N_17991,N_16589,N_16723);
and U17992 (N_17992,N_16816,N_16487);
xnor U17993 (N_17993,N_16449,N_16476);
nand U17994 (N_17994,N_16076,N_16880);
or U17995 (N_17995,N_16056,N_16002);
and U17996 (N_17996,N_16998,N_16595);
nor U17997 (N_17997,N_16445,N_16120);
nand U17998 (N_17998,N_16930,N_16097);
nor U17999 (N_17999,N_16518,N_16322);
and U18000 (N_18000,N_17232,N_17165);
or U18001 (N_18001,N_17996,N_17277);
nor U18002 (N_18002,N_17004,N_17691);
and U18003 (N_18003,N_17158,N_17423);
nor U18004 (N_18004,N_17774,N_17023);
xnor U18005 (N_18005,N_17109,N_17933);
nand U18006 (N_18006,N_17212,N_17450);
and U18007 (N_18007,N_17640,N_17100);
and U18008 (N_18008,N_17539,N_17901);
nor U18009 (N_18009,N_17545,N_17818);
nand U18010 (N_18010,N_17571,N_17510);
or U18011 (N_18011,N_17718,N_17657);
and U18012 (N_18012,N_17059,N_17337);
nand U18013 (N_18013,N_17127,N_17446);
nor U18014 (N_18014,N_17819,N_17754);
or U18015 (N_18015,N_17010,N_17578);
or U18016 (N_18016,N_17550,N_17434);
xor U18017 (N_18017,N_17977,N_17912);
nor U18018 (N_18018,N_17359,N_17522);
nand U18019 (N_18019,N_17712,N_17982);
and U18020 (N_18020,N_17284,N_17231);
nand U18021 (N_18021,N_17855,N_17864);
or U18022 (N_18022,N_17590,N_17856);
nand U18023 (N_18023,N_17763,N_17064);
nand U18024 (N_18024,N_17796,N_17995);
xnor U18025 (N_18025,N_17611,N_17409);
xor U18026 (N_18026,N_17281,N_17719);
xor U18027 (N_18027,N_17119,N_17968);
nand U18028 (N_18028,N_17046,N_17956);
nor U18029 (N_18029,N_17765,N_17114);
or U18030 (N_18030,N_17490,N_17523);
or U18031 (N_18031,N_17186,N_17817);
nand U18032 (N_18032,N_17483,N_17683);
xor U18033 (N_18033,N_17316,N_17584);
and U18034 (N_18034,N_17549,N_17824);
or U18035 (N_18035,N_17932,N_17036);
nor U18036 (N_18036,N_17179,N_17356);
or U18037 (N_18037,N_17831,N_17069);
or U18038 (N_18038,N_17172,N_17162);
xor U18039 (N_18039,N_17641,N_17335);
nand U18040 (N_18040,N_17392,N_17779);
nor U18041 (N_18041,N_17776,N_17900);
or U18042 (N_18042,N_17676,N_17227);
nand U18043 (N_18043,N_17369,N_17123);
xor U18044 (N_18044,N_17040,N_17480);
xor U18045 (N_18045,N_17606,N_17519);
xor U18046 (N_18046,N_17031,N_17574);
or U18047 (N_18047,N_17960,N_17126);
nor U18048 (N_18048,N_17628,N_17426);
nor U18049 (N_18049,N_17035,N_17654);
nor U18050 (N_18050,N_17883,N_17703);
nand U18051 (N_18051,N_17467,N_17698);
xnor U18052 (N_18052,N_17219,N_17210);
or U18053 (N_18053,N_17319,N_17842);
nand U18054 (N_18054,N_17194,N_17854);
xnor U18055 (N_18055,N_17156,N_17500);
nand U18056 (N_18056,N_17680,N_17979);
or U18057 (N_18057,N_17800,N_17825);
and U18058 (N_18058,N_17432,N_17512);
xnor U18059 (N_18059,N_17853,N_17906);
or U18060 (N_18060,N_17192,N_17221);
xor U18061 (N_18061,N_17895,N_17844);
nand U18062 (N_18062,N_17273,N_17239);
nand U18063 (N_18063,N_17903,N_17990);
nor U18064 (N_18064,N_17575,N_17728);
xnor U18065 (N_18065,N_17044,N_17508);
or U18066 (N_18066,N_17799,N_17453);
xnor U18067 (N_18067,N_17645,N_17286);
nand U18068 (N_18068,N_17644,N_17345);
nand U18069 (N_18069,N_17967,N_17711);
or U18070 (N_18070,N_17878,N_17525);
or U18071 (N_18071,N_17976,N_17740);
nand U18072 (N_18072,N_17671,N_17601);
or U18073 (N_18073,N_17358,N_17433);
nor U18074 (N_18074,N_17049,N_17627);
nand U18075 (N_18075,N_17837,N_17940);
nor U18076 (N_18076,N_17764,N_17175);
nor U18077 (N_18077,N_17945,N_17177);
xor U18078 (N_18078,N_17889,N_17472);
or U18079 (N_18079,N_17843,N_17595);
xnor U18080 (N_18080,N_17669,N_17159);
xnor U18081 (N_18081,N_17516,N_17672);
or U18082 (N_18082,N_17767,N_17727);
or U18083 (N_18083,N_17737,N_17975);
nor U18084 (N_18084,N_17786,N_17447);
nand U18085 (N_18085,N_17095,N_17057);
xnor U18086 (N_18086,N_17350,N_17198);
nor U18087 (N_18087,N_17521,N_17213);
and U18088 (N_18088,N_17424,N_17581);
and U18089 (N_18089,N_17802,N_17759);
nand U18090 (N_18090,N_17464,N_17913);
or U18091 (N_18091,N_17739,N_17407);
nand U18092 (N_18092,N_17007,N_17371);
and U18093 (N_18093,N_17812,N_17093);
and U18094 (N_18094,N_17616,N_17043);
or U18095 (N_18095,N_17195,N_17448);
nor U18096 (N_18096,N_17478,N_17773);
xnor U18097 (N_18097,N_17931,N_17307);
or U18098 (N_18098,N_17005,N_17924);
and U18099 (N_18099,N_17013,N_17086);
nand U18100 (N_18100,N_17757,N_17816);
nor U18101 (N_18101,N_17230,N_17380);
xor U18102 (N_18102,N_17829,N_17922);
or U18103 (N_18103,N_17041,N_17804);
nor U18104 (N_18104,N_17164,N_17658);
and U18105 (N_18105,N_17839,N_17009);
and U18106 (N_18106,N_17511,N_17866);
or U18107 (N_18107,N_17139,N_17920);
nand U18108 (N_18108,N_17270,N_17425);
or U18109 (N_18109,N_17994,N_17451);
nand U18110 (N_18110,N_17257,N_17886);
or U18111 (N_18111,N_17012,N_17904);
or U18112 (N_18112,N_17325,N_17075);
nor U18113 (N_18113,N_17914,N_17459);
xnor U18114 (N_18114,N_17414,N_17838);
or U18115 (N_18115,N_17961,N_17813);
or U18116 (N_18116,N_17463,N_17921);
or U18117 (N_18117,N_17386,N_17531);
xor U18118 (N_18118,N_17437,N_17378);
and U18119 (N_18119,N_17555,N_17338);
xnor U18120 (N_18120,N_17300,N_17544);
and U18121 (N_18121,N_17588,N_17626);
nor U18122 (N_18122,N_17120,N_17428);
and U18123 (N_18123,N_17937,N_17241);
nand U18124 (N_18124,N_17798,N_17454);
or U18125 (N_18125,N_17534,N_17874);
nor U18126 (N_18126,N_17193,N_17305);
or U18127 (N_18127,N_17502,N_17706);
nor U18128 (N_18128,N_17214,N_17959);
xnor U18129 (N_18129,N_17520,N_17234);
or U18130 (N_18130,N_17998,N_17268);
and U18131 (N_18131,N_17220,N_17140);
xnor U18132 (N_18132,N_17117,N_17692);
and U18133 (N_18133,N_17686,N_17366);
xor U18134 (N_18134,N_17621,N_17872);
xor U18135 (N_18135,N_17456,N_17833);
and U18136 (N_18136,N_17289,N_17788);
nor U18137 (N_18137,N_17282,N_17943);
or U18138 (N_18138,N_17142,N_17184);
and U18139 (N_18139,N_17868,N_17202);
nand U18140 (N_18140,N_17431,N_17260);
and U18141 (N_18141,N_17176,N_17374);
and U18142 (N_18142,N_17527,N_17782);
nand U18143 (N_18143,N_17488,N_17361);
and U18144 (N_18144,N_17529,N_17614);
xnor U18145 (N_18145,N_17479,N_17935);
and U18146 (N_18146,N_17958,N_17503);
nor U18147 (N_18147,N_17694,N_17381);
nand U18148 (N_18148,N_17548,N_17551);
or U18149 (N_18149,N_17981,N_17188);
and U18150 (N_18150,N_17929,N_17665);
nor U18151 (N_18151,N_17097,N_17777);
and U18152 (N_18152,N_17725,N_17385);
nor U18153 (N_18153,N_17084,N_17707);
and U18154 (N_18154,N_17185,N_17072);
and U18155 (N_18155,N_17291,N_17887);
nand U18156 (N_18156,N_17587,N_17032);
nor U18157 (N_18157,N_17939,N_17331);
xor U18158 (N_18158,N_17318,N_17803);
or U18159 (N_18159,N_17417,N_17615);
nand U18160 (N_18160,N_17731,N_17546);
nor U18161 (N_18161,N_17293,N_17211);
nor U18162 (N_18162,N_17746,N_17443);
xor U18163 (N_18163,N_17476,N_17181);
and U18164 (N_18164,N_17577,N_17078);
xnor U18165 (N_18165,N_17966,N_17743);
and U18166 (N_18166,N_17849,N_17993);
or U18167 (N_18167,N_17659,N_17729);
and U18168 (N_18168,N_17637,N_17780);
xor U18169 (N_18169,N_17340,N_17000);
xnor U18170 (N_18170,N_17458,N_17905);
nand U18171 (N_18171,N_17047,N_17492);
nand U18172 (N_18172,N_17341,N_17149);
and U18173 (N_18173,N_17791,N_17760);
and U18174 (N_18174,N_17848,N_17267);
nor U18175 (N_18175,N_17630,N_17962);
or U18176 (N_18176,N_17021,N_17205);
and U18177 (N_18177,N_17222,N_17784);
or U18178 (N_18178,N_17794,N_17789);
xor U18179 (N_18179,N_17955,N_17438);
nand U18180 (N_18180,N_17643,N_17808);
or U18181 (N_18181,N_17190,N_17888);
nand U18182 (N_18182,N_17042,N_17399);
nand U18183 (N_18183,N_17363,N_17673);
nor U18184 (N_18184,N_17790,N_17554);
xor U18185 (N_18185,N_17594,N_17517);
or U18186 (N_18186,N_17295,N_17944);
or U18187 (N_18187,N_17250,N_17382);
nor U18188 (N_18188,N_17468,N_17070);
or U18189 (N_18189,N_17092,N_17001);
or U18190 (N_18190,N_17999,N_17034);
or U18191 (N_18191,N_17863,N_17173);
nand U18192 (N_18192,N_17543,N_17597);
and U18193 (N_18193,N_17607,N_17283);
nor U18194 (N_18194,N_17907,N_17721);
and U18195 (N_18195,N_17408,N_17208);
xor U18196 (N_18196,N_17207,N_17144);
and U18197 (N_18197,N_17766,N_17389);
xor U18198 (N_18198,N_17783,N_17357);
or U18199 (N_18199,N_17807,N_17376);
and U18200 (N_18200,N_17695,N_17327);
xor U18201 (N_18201,N_17169,N_17074);
or U18202 (N_18202,N_17246,N_17877);
xor U18203 (N_18203,N_17589,N_17237);
nor U18204 (N_18204,N_17952,N_17814);
or U18205 (N_18205,N_17401,N_17602);
nor U18206 (N_18206,N_17623,N_17751);
nand U18207 (N_18207,N_17992,N_17876);
nor U18208 (N_18208,N_17936,N_17068);
or U18209 (N_18209,N_17513,N_17847);
nand U18210 (N_18210,N_17017,N_17865);
or U18211 (N_18211,N_17138,N_17612);
nand U18212 (N_18212,N_17850,N_17836);
or U18213 (N_18213,N_17352,N_17562);
nand U18214 (N_18214,N_17247,N_17163);
nor U18215 (N_18215,N_17832,N_17244);
xor U18216 (N_18216,N_17094,N_17859);
or U18217 (N_18217,N_17226,N_17276);
and U18218 (N_18218,N_17153,N_17653);
nor U18219 (N_18219,N_17661,N_17349);
nor U18220 (N_18220,N_17598,N_17882);
nand U18221 (N_18221,N_17570,N_17430);
xnor U18222 (N_18222,N_17797,N_17398);
nand U18223 (N_18223,N_17403,N_17233);
or U18224 (N_18224,N_17506,N_17870);
and U18225 (N_18225,N_17178,N_17948);
nand U18226 (N_18226,N_17209,N_17274);
nor U18227 (N_18227,N_17667,N_17028);
or U18228 (N_18228,N_17465,N_17528);
and U18229 (N_18229,N_17620,N_17930);
and U18230 (N_18230,N_17189,N_17526);
nor U18231 (N_18231,N_17419,N_17280);
nand U18232 (N_18232,N_17333,N_17137);
nand U18233 (N_18233,N_17795,N_17862);
nor U18234 (N_18234,N_17923,N_17957);
or U18235 (N_18235,N_17204,N_17501);
nor U18236 (N_18236,N_17342,N_17772);
or U18237 (N_18237,N_17801,N_17826);
nand U18238 (N_18238,N_17805,N_17726);
nand U18239 (N_18239,N_17851,N_17778);
or U18240 (N_18240,N_17321,N_17604);
xor U18241 (N_18241,N_17312,N_17128);
and U18242 (N_18242,N_17063,N_17735);
and U18243 (N_18243,N_17006,N_17418);
nand U18244 (N_18244,N_17915,N_17600);
and U18245 (N_18245,N_17368,N_17015);
xnor U18246 (N_18246,N_17749,N_17593);
xnor U18247 (N_18247,N_17089,N_17422);
xor U18248 (N_18248,N_17974,N_17730);
or U18249 (N_18249,N_17633,N_17048);
and U18250 (N_18250,N_17540,N_17771);
nand U18251 (N_18251,N_17395,N_17987);
and U18252 (N_18252,N_17910,N_17390);
and U18253 (N_18253,N_17420,N_17224);
and U18254 (N_18254,N_17793,N_17055);
and U18255 (N_18255,N_17984,N_17107);
nor U18256 (N_18256,N_17411,N_17569);
xor U18257 (N_18257,N_17973,N_17689);
xor U18258 (N_18258,N_17662,N_17556);
or U18259 (N_18259,N_17256,N_17652);
or U18260 (N_18260,N_17634,N_17462);
and U18261 (N_18261,N_17037,N_17560);
nor U18262 (N_18262,N_17391,N_17457);
and U18263 (N_18263,N_17917,N_17756);
or U18264 (N_18264,N_17879,N_17925);
nand U18265 (N_18265,N_17442,N_17473);
nor U18266 (N_18266,N_17471,N_17716);
nand U18267 (N_18267,N_17532,N_17622);
or U18268 (N_18268,N_17646,N_17171);
nand U18269 (N_18269,N_17781,N_17474);
xor U18270 (N_18270,N_17576,N_17154);
xor U18271 (N_18271,N_17902,N_17505);
nor U18272 (N_18272,N_17991,N_17867);
or U18273 (N_18273,N_17322,N_17460);
nor U18274 (N_18274,N_17732,N_17315);
or U18275 (N_18275,N_17088,N_17263);
or U18276 (N_18276,N_17747,N_17083);
nand U18277 (N_18277,N_17236,N_17304);
nand U18278 (N_18278,N_17559,N_17493);
or U18279 (N_18279,N_17421,N_17235);
nand U18280 (N_18280,N_17741,N_17373);
nand U18281 (N_18281,N_17264,N_17722);
xor U18282 (N_18282,N_17191,N_17020);
nand U18283 (N_18283,N_17636,N_17497);
nor U18284 (N_18284,N_17477,N_17846);
or U18285 (N_18285,N_17537,N_17113);
xor U18286 (N_18286,N_17413,N_17161);
xor U18287 (N_18287,N_17563,N_17125);
nand U18288 (N_18288,N_17946,N_17384);
nor U18289 (N_18289,N_17324,N_17150);
xor U18290 (N_18290,N_17388,N_17610);
or U18291 (N_18291,N_17223,N_17452);
or U18292 (N_18292,N_17954,N_17104);
or U18293 (N_18293,N_17314,N_17926);
or U18294 (N_18294,N_17822,N_17033);
and U18295 (N_18295,N_17367,N_17174);
nor U18296 (N_18296,N_17152,N_17656);
and U18297 (N_18297,N_17196,N_17518);
nand U18298 (N_18298,N_17542,N_17266);
nand U18299 (N_18299,N_17690,N_17498);
nand U18300 (N_18300,N_17182,N_17168);
nor U18301 (N_18301,N_17909,N_17297);
or U18302 (N_18302,N_17538,N_17115);
xnor U18303 (N_18303,N_17348,N_17347);
nand U18304 (N_18304,N_17582,N_17255);
xnor U18305 (N_18305,N_17030,N_17484);
nor U18306 (N_18306,N_17670,N_17927);
and U18307 (N_18307,N_17820,N_17200);
nor U18308 (N_18308,N_17440,N_17141);
nor U18309 (N_18309,N_17339,N_17404);
nor U18310 (N_18310,N_17116,N_17899);
xnor U18311 (N_18311,N_17215,N_17827);
nand U18312 (N_18312,N_17775,N_17252);
and U18313 (N_18313,N_17061,N_17112);
nand U18314 (N_18314,N_17229,N_17353);
or U18315 (N_18315,N_17753,N_17320);
nor U18316 (N_18316,N_17714,N_17145);
and U18317 (N_18317,N_17253,N_17080);
nor U18318 (N_18318,N_17811,N_17285);
xor U18319 (N_18319,N_17087,N_17218);
and U18320 (N_18320,N_17110,N_17029);
or U18321 (N_18321,N_17343,N_17894);
or U18322 (N_18322,N_17122,N_17547);
xnor U18323 (N_18323,N_17770,N_17287);
xnor U18324 (N_18324,N_17713,N_17206);
nand U18325 (N_18325,N_17290,N_17259);
nand U18326 (N_18326,N_17891,N_17038);
nor U18327 (N_18327,N_17166,N_17199);
or U18328 (N_18328,N_17132,N_17393);
or U18329 (N_18329,N_17278,N_17596);
nand U18330 (N_18330,N_17011,N_17081);
xnor U18331 (N_18331,N_17989,N_17328);
or U18332 (N_18332,N_17697,N_17121);
and U18333 (N_18333,N_17858,N_17261);
and U18334 (N_18334,N_17752,N_17299);
and U18335 (N_18335,N_17288,N_17524);
nand U18336 (N_18336,N_17592,N_17014);
and U18337 (N_18337,N_17102,N_17701);
nand U18338 (N_18338,N_17918,N_17271);
or U18339 (N_18339,N_17823,N_17334);
nor U18340 (N_18340,N_17613,N_17370);
nor U18341 (N_18341,N_17648,N_17082);
and U18342 (N_18342,N_17830,N_17402);
xor U18343 (N_18343,N_17609,N_17496);
nand U18344 (N_18344,N_17580,N_17455);
or U18345 (N_18345,N_17362,N_17435);
xor U18346 (N_18346,N_17265,N_17301);
and U18347 (N_18347,N_17022,N_17101);
nand U18348 (N_18348,N_17769,N_17552);
nor U18349 (N_18349,N_17792,N_17618);
nor U18350 (N_18350,N_17916,N_17629);
nand U18351 (N_18351,N_17884,N_17514);
and U18352 (N_18352,N_17131,N_17225);
xor U18353 (N_18353,N_17262,N_17558);
and U18354 (N_18354,N_17568,N_17875);
or U18355 (N_18355,N_17449,N_17566);
xnor U18356 (N_18356,N_17852,N_17026);
xor U18357 (N_18357,N_17762,N_17396);
nor U18358 (N_18358,N_17986,N_17310);
and U18359 (N_18359,N_17509,N_17018);
nor U18360 (N_18360,N_17085,N_17561);
xnor U18361 (N_18361,N_17275,N_17696);
nand U18362 (N_18362,N_17016,N_17573);
nor U18363 (N_18363,N_17896,N_17638);
xnor U18364 (N_18364,N_17323,N_17311);
xnor U18365 (N_18365,N_17062,N_17723);
and U18366 (N_18366,N_17099,N_17655);
or U18367 (N_18367,N_17893,N_17679);
nand U18368 (N_18368,N_17167,N_17329);
xnor U18369 (N_18369,N_17885,N_17296);
or U18370 (N_18370,N_17203,N_17675);
and U18371 (N_18371,N_17605,N_17412);
or U18372 (N_18372,N_17845,N_17685);
xor U18373 (N_18373,N_17564,N_17201);
nor U18374 (N_18374,N_17745,N_17249);
nor U18375 (N_18375,N_17639,N_17332);
nor U18376 (N_18376,N_17079,N_17736);
xnor U18377 (N_18377,N_17585,N_17346);
xnor U18378 (N_18378,N_17649,N_17969);
xnor U18379 (N_18379,N_17942,N_17717);
and U18380 (N_18380,N_17130,N_17755);
nor U18381 (N_18381,N_17980,N_17330);
nand U18382 (N_18382,N_17197,N_17748);
xnor U18383 (N_18383,N_17365,N_17272);
xor U18384 (N_18384,N_17027,N_17687);
or U18385 (N_18385,N_17583,N_17668);
xnor U18386 (N_18386,N_17216,N_17688);
or U18387 (N_18387,N_17486,N_17003);
nand U18388 (N_18388,N_17090,N_17427);
nand U18389 (N_18389,N_17938,N_17586);
xnor U18390 (N_18390,N_17415,N_17351);
nand U18391 (N_18391,N_17445,N_17025);
or U18392 (N_18392,N_17060,N_17183);
nor U18393 (N_18393,N_17809,N_17377);
or U18394 (N_18394,N_17810,N_17572);
and U18395 (N_18395,N_17619,N_17024);
xnor U18396 (N_18396,N_17143,N_17002);
or U18397 (N_18397,N_17096,N_17344);
and U18398 (N_18398,N_17105,N_17983);
nor U18399 (N_18399,N_17058,N_17147);
xor U18400 (N_18400,N_17306,N_17504);
xor U18401 (N_18401,N_17785,N_17705);
xor U18402 (N_18402,N_17302,N_17245);
or U18403 (N_18403,N_17515,N_17146);
or U18404 (N_18404,N_17439,N_17397);
nand U18405 (N_18405,N_17536,N_17603);
and U18406 (N_18406,N_17317,N_17056);
nor U18407 (N_18407,N_17269,N_17313);
and U18408 (N_18408,N_17951,N_17469);
and U18409 (N_18409,N_17118,N_17066);
xnor U18410 (N_18410,N_17674,N_17405);
xnor U18411 (N_18411,N_17591,N_17880);
and U18412 (N_18412,N_17892,N_17298);
and U18413 (N_18413,N_17157,N_17180);
nand U18414 (N_18414,N_17632,N_17054);
xor U18415 (N_18415,N_17535,N_17077);
nand U18416 (N_18416,N_17869,N_17530);
nor U18417 (N_18417,N_17664,N_17360);
nor U18418 (N_18418,N_17111,N_17155);
and U18419 (N_18419,N_17985,N_17828);
nor U18420 (N_18420,N_17734,N_17941);
nand U18421 (N_18421,N_17466,N_17187);
and U18422 (N_18422,N_17103,N_17485);
xor U18423 (N_18423,N_17039,N_17553);
and U18424 (N_18424,N_17461,N_17702);
and U18425 (N_18425,N_17650,N_17170);
and U18426 (N_18426,N_17651,N_17821);
nand U18427 (N_18427,N_17890,N_17733);
xnor U18428 (N_18428,N_17949,N_17908);
nor U18429 (N_18429,N_17700,N_17254);
nor U18430 (N_18430,N_17708,N_17738);
xor U18431 (N_18431,N_17963,N_17787);
xnor U18432 (N_18432,N_17684,N_17965);
xnor U18433 (N_18433,N_17238,N_17815);
nor U18434 (N_18434,N_17475,N_17148);
nand U18435 (N_18435,N_17482,N_17608);
xor U18436 (N_18436,N_17091,N_17248);
or U18437 (N_18437,N_17898,N_17052);
and U18438 (N_18438,N_17950,N_17507);
nand U18439 (N_18439,N_17019,N_17383);
nand U18440 (N_18440,N_17067,N_17410);
or U18441 (N_18441,N_17860,N_17897);
and U18442 (N_18442,N_17861,N_17258);
or U18443 (N_18443,N_17677,N_17617);
or U18444 (N_18444,N_17136,N_17978);
xnor U18445 (N_18445,N_17567,N_17441);
nor U18446 (N_18446,N_17704,N_17071);
and U18447 (N_18447,N_17699,N_17354);
or U18448 (N_18448,N_17710,N_17750);
nor U18449 (N_18449,N_17294,N_17487);
nand U18450 (N_18450,N_17364,N_17709);
or U18451 (N_18451,N_17744,N_17124);
nand U18452 (N_18452,N_17768,N_17647);
or U18453 (N_18453,N_17631,N_17599);
xnor U18454 (N_18454,N_17133,N_17481);
and U18455 (N_18455,N_17565,N_17372);
xor U18456 (N_18456,N_17416,N_17579);
and U18457 (N_18457,N_17635,N_17303);
nand U18458 (N_18458,N_17715,N_17720);
or U18459 (N_18459,N_17494,N_17625);
xor U18460 (N_18460,N_17624,N_17911);
xnor U18461 (N_18461,N_17065,N_17988);
or U18462 (N_18462,N_17873,N_17151);
and U18463 (N_18463,N_17953,N_17928);
or U18464 (N_18464,N_17841,N_17073);
nand U18465 (N_18465,N_17436,N_17678);
nand U18466 (N_18466,N_17499,N_17919);
xor U18467 (N_18467,N_17533,N_17660);
nor U18468 (N_18468,N_17008,N_17135);
xnor U18469 (N_18469,N_17129,N_17106);
xnor U18470 (N_18470,N_17541,N_17682);
and U18471 (N_18471,N_17758,N_17681);
nand U18472 (N_18472,N_17693,N_17308);
or U18473 (N_18473,N_17076,N_17108);
nor U18474 (N_18474,N_17242,N_17964);
or U18475 (N_18475,N_17050,N_17495);
or U18476 (N_18476,N_17228,N_17871);
nand U18477 (N_18477,N_17834,N_17217);
xor U18478 (N_18478,N_17806,N_17663);
and U18479 (N_18479,N_17934,N_17970);
xor U18480 (N_18480,N_17279,N_17251);
or U18481 (N_18481,N_17666,N_17489);
xor U18482 (N_18482,N_17309,N_17406);
or U18483 (N_18483,N_17051,N_17387);
or U18484 (N_18484,N_17444,N_17243);
and U18485 (N_18485,N_17053,N_17947);
or U18486 (N_18486,N_17240,N_17724);
nand U18487 (N_18487,N_17742,N_17160);
nor U18488 (N_18488,N_17379,N_17098);
nand U18489 (N_18489,N_17761,N_17971);
nor U18490 (N_18490,N_17557,N_17429);
nand U18491 (N_18491,N_17470,N_17355);
and U18492 (N_18492,N_17326,N_17835);
nand U18493 (N_18493,N_17840,N_17045);
and U18494 (N_18494,N_17642,N_17336);
nand U18495 (N_18495,N_17292,N_17375);
or U18496 (N_18496,N_17134,N_17881);
nor U18497 (N_18497,N_17400,N_17857);
nor U18498 (N_18498,N_17972,N_17997);
nor U18499 (N_18499,N_17491,N_17394);
and U18500 (N_18500,N_17965,N_17890);
nand U18501 (N_18501,N_17073,N_17678);
or U18502 (N_18502,N_17602,N_17907);
xor U18503 (N_18503,N_17376,N_17494);
nand U18504 (N_18504,N_17327,N_17110);
xnor U18505 (N_18505,N_17161,N_17457);
nand U18506 (N_18506,N_17689,N_17176);
nor U18507 (N_18507,N_17026,N_17262);
xor U18508 (N_18508,N_17546,N_17161);
nand U18509 (N_18509,N_17752,N_17641);
nand U18510 (N_18510,N_17754,N_17156);
and U18511 (N_18511,N_17448,N_17245);
xnor U18512 (N_18512,N_17260,N_17158);
xnor U18513 (N_18513,N_17140,N_17271);
nand U18514 (N_18514,N_17071,N_17318);
nor U18515 (N_18515,N_17114,N_17379);
or U18516 (N_18516,N_17880,N_17308);
xnor U18517 (N_18517,N_17069,N_17663);
and U18518 (N_18518,N_17250,N_17967);
xnor U18519 (N_18519,N_17603,N_17947);
nor U18520 (N_18520,N_17704,N_17172);
nor U18521 (N_18521,N_17882,N_17317);
nor U18522 (N_18522,N_17440,N_17998);
and U18523 (N_18523,N_17722,N_17551);
and U18524 (N_18524,N_17963,N_17299);
nor U18525 (N_18525,N_17110,N_17958);
or U18526 (N_18526,N_17413,N_17181);
and U18527 (N_18527,N_17021,N_17321);
nand U18528 (N_18528,N_17402,N_17852);
nor U18529 (N_18529,N_17499,N_17173);
nand U18530 (N_18530,N_17674,N_17269);
nor U18531 (N_18531,N_17714,N_17446);
and U18532 (N_18532,N_17881,N_17808);
xor U18533 (N_18533,N_17234,N_17609);
nor U18534 (N_18534,N_17322,N_17850);
nor U18535 (N_18535,N_17313,N_17408);
nand U18536 (N_18536,N_17348,N_17822);
xor U18537 (N_18537,N_17763,N_17011);
xnor U18538 (N_18538,N_17660,N_17643);
xor U18539 (N_18539,N_17517,N_17270);
xor U18540 (N_18540,N_17741,N_17317);
and U18541 (N_18541,N_17304,N_17771);
xor U18542 (N_18542,N_17392,N_17521);
nand U18543 (N_18543,N_17271,N_17843);
or U18544 (N_18544,N_17741,N_17772);
nor U18545 (N_18545,N_17150,N_17805);
and U18546 (N_18546,N_17623,N_17933);
xnor U18547 (N_18547,N_17501,N_17390);
and U18548 (N_18548,N_17775,N_17096);
nor U18549 (N_18549,N_17667,N_17271);
nand U18550 (N_18550,N_17383,N_17608);
nand U18551 (N_18551,N_17517,N_17228);
nor U18552 (N_18552,N_17655,N_17241);
or U18553 (N_18553,N_17016,N_17395);
nand U18554 (N_18554,N_17931,N_17925);
and U18555 (N_18555,N_17370,N_17298);
nand U18556 (N_18556,N_17011,N_17581);
or U18557 (N_18557,N_17501,N_17705);
or U18558 (N_18558,N_17803,N_17602);
xnor U18559 (N_18559,N_17780,N_17534);
or U18560 (N_18560,N_17876,N_17469);
nand U18561 (N_18561,N_17995,N_17285);
xor U18562 (N_18562,N_17123,N_17470);
xnor U18563 (N_18563,N_17540,N_17159);
or U18564 (N_18564,N_17453,N_17849);
nand U18565 (N_18565,N_17701,N_17709);
xor U18566 (N_18566,N_17528,N_17496);
and U18567 (N_18567,N_17851,N_17326);
and U18568 (N_18568,N_17706,N_17246);
and U18569 (N_18569,N_17152,N_17125);
nor U18570 (N_18570,N_17495,N_17951);
nand U18571 (N_18571,N_17816,N_17609);
nor U18572 (N_18572,N_17858,N_17106);
nand U18573 (N_18573,N_17052,N_17612);
xnor U18574 (N_18574,N_17861,N_17054);
or U18575 (N_18575,N_17858,N_17220);
xnor U18576 (N_18576,N_17731,N_17195);
or U18577 (N_18577,N_17075,N_17032);
nand U18578 (N_18578,N_17350,N_17820);
or U18579 (N_18579,N_17553,N_17186);
xor U18580 (N_18580,N_17007,N_17432);
nand U18581 (N_18581,N_17249,N_17390);
or U18582 (N_18582,N_17821,N_17252);
and U18583 (N_18583,N_17022,N_17418);
or U18584 (N_18584,N_17233,N_17173);
nor U18585 (N_18585,N_17510,N_17316);
xor U18586 (N_18586,N_17198,N_17493);
and U18587 (N_18587,N_17535,N_17538);
nand U18588 (N_18588,N_17004,N_17768);
nand U18589 (N_18589,N_17900,N_17465);
nor U18590 (N_18590,N_17820,N_17613);
or U18591 (N_18591,N_17217,N_17720);
and U18592 (N_18592,N_17416,N_17982);
or U18593 (N_18593,N_17479,N_17918);
nand U18594 (N_18594,N_17485,N_17234);
nor U18595 (N_18595,N_17650,N_17528);
nor U18596 (N_18596,N_17113,N_17518);
nand U18597 (N_18597,N_17890,N_17083);
xor U18598 (N_18598,N_17260,N_17678);
xor U18599 (N_18599,N_17478,N_17531);
or U18600 (N_18600,N_17240,N_17116);
nor U18601 (N_18601,N_17232,N_17410);
and U18602 (N_18602,N_17080,N_17408);
xor U18603 (N_18603,N_17339,N_17096);
nand U18604 (N_18604,N_17532,N_17763);
or U18605 (N_18605,N_17855,N_17575);
or U18606 (N_18606,N_17537,N_17042);
nor U18607 (N_18607,N_17726,N_17022);
nor U18608 (N_18608,N_17562,N_17612);
nand U18609 (N_18609,N_17558,N_17101);
nor U18610 (N_18610,N_17101,N_17720);
and U18611 (N_18611,N_17328,N_17890);
and U18612 (N_18612,N_17907,N_17168);
nor U18613 (N_18613,N_17067,N_17178);
and U18614 (N_18614,N_17730,N_17300);
nor U18615 (N_18615,N_17137,N_17070);
or U18616 (N_18616,N_17738,N_17397);
xor U18617 (N_18617,N_17552,N_17194);
and U18618 (N_18618,N_17765,N_17410);
xnor U18619 (N_18619,N_17029,N_17535);
xnor U18620 (N_18620,N_17088,N_17218);
xnor U18621 (N_18621,N_17081,N_17907);
nor U18622 (N_18622,N_17236,N_17418);
and U18623 (N_18623,N_17173,N_17218);
nand U18624 (N_18624,N_17357,N_17079);
or U18625 (N_18625,N_17805,N_17385);
xnor U18626 (N_18626,N_17413,N_17036);
nor U18627 (N_18627,N_17536,N_17806);
nand U18628 (N_18628,N_17790,N_17683);
nor U18629 (N_18629,N_17300,N_17444);
and U18630 (N_18630,N_17124,N_17455);
or U18631 (N_18631,N_17043,N_17153);
or U18632 (N_18632,N_17975,N_17476);
nand U18633 (N_18633,N_17377,N_17957);
and U18634 (N_18634,N_17175,N_17248);
nor U18635 (N_18635,N_17308,N_17210);
or U18636 (N_18636,N_17695,N_17530);
nand U18637 (N_18637,N_17961,N_17156);
nor U18638 (N_18638,N_17553,N_17333);
and U18639 (N_18639,N_17311,N_17303);
nor U18640 (N_18640,N_17857,N_17428);
xor U18641 (N_18641,N_17771,N_17963);
xor U18642 (N_18642,N_17023,N_17094);
nor U18643 (N_18643,N_17181,N_17130);
nor U18644 (N_18644,N_17958,N_17504);
xor U18645 (N_18645,N_17935,N_17512);
and U18646 (N_18646,N_17840,N_17719);
and U18647 (N_18647,N_17002,N_17974);
nor U18648 (N_18648,N_17703,N_17773);
and U18649 (N_18649,N_17244,N_17530);
xnor U18650 (N_18650,N_17803,N_17458);
and U18651 (N_18651,N_17191,N_17275);
and U18652 (N_18652,N_17096,N_17099);
and U18653 (N_18653,N_17764,N_17279);
nor U18654 (N_18654,N_17254,N_17591);
and U18655 (N_18655,N_17708,N_17294);
nand U18656 (N_18656,N_17984,N_17717);
or U18657 (N_18657,N_17730,N_17581);
and U18658 (N_18658,N_17642,N_17537);
nand U18659 (N_18659,N_17987,N_17981);
xor U18660 (N_18660,N_17704,N_17228);
xor U18661 (N_18661,N_17639,N_17148);
and U18662 (N_18662,N_17406,N_17189);
or U18663 (N_18663,N_17687,N_17731);
or U18664 (N_18664,N_17964,N_17191);
and U18665 (N_18665,N_17094,N_17416);
and U18666 (N_18666,N_17288,N_17154);
or U18667 (N_18667,N_17801,N_17015);
and U18668 (N_18668,N_17637,N_17760);
or U18669 (N_18669,N_17229,N_17039);
or U18670 (N_18670,N_17423,N_17633);
nand U18671 (N_18671,N_17715,N_17311);
or U18672 (N_18672,N_17092,N_17337);
or U18673 (N_18673,N_17529,N_17994);
or U18674 (N_18674,N_17900,N_17712);
nor U18675 (N_18675,N_17850,N_17734);
nand U18676 (N_18676,N_17264,N_17451);
nand U18677 (N_18677,N_17065,N_17881);
nand U18678 (N_18678,N_17633,N_17865);
and U18679 (N_18679,N_17778,N_17456);
nor U18680 (N_18680,N_17533,N_17119);
nand U18681 (N_18681,N_17471,N_17074);
nor U18682 (N_18682,N_17379,N_17943);
xnor U18683 (N_18683,N_17931,N_17430);
xnor U18684 (N_18684,N_17452,N_17639);
and U18685 (N_18685,N_17210,N_17177);
nor U18686 (N_18686,N_17357,N_17477);
nor U18687 (N_18687,N_17061,N_17278);
nor U18688 (N_18688,N_17764,N_17214);
nand U18689 (N_18689,N_17059,N_17277);
or U18690 (N_18690,N_17739,N_17118);
xnor U18691 (N_18691,N_17021,N_17074);
nor U18692 (N_18692,N_17716,N_17068);
and U18693 (N_18693,N_17399,N_17171);
xnor U18694 (N_18694,N_17108,N_17299);
or U18695 (N_18695,N_17669,N_17053);
nor U18696 (N_18696,N_17575,N_17690);
xnor U18697 (N_18697,N_17520,N_17581);
or U18698 (N_18698,N_17787,N_17770);
xor U18699 (N_18699,N_17955,N_17302);
and U18700 (N_18700,N_17798,N_17916);
xnor U18701 (N_18701,N_17272,N_17933);
and U18702 (N_18702,N_17379,N_17743);
xor U18703 (N_18703,N_17499,N_17473);
or U18704 (N_18704,N_17099,N_17268);
xor U18705 (N_18705,N_17763,N_17431);
and U18706 (N_18706,N_17879,N_17579);
or U18707 (N_18707,N_17116,N_17357);
and U18708 (N_18708,N_17499,N_17608);
nor U18709 (N_18709,N_17683,N_17490);
nor U18710 (N_18710,N_17928,N_17576);
and U18711 (N_18711,N_17666,N_17370);
nand U18712 (N_18712,N_17967,N_17046);
nand U18713 (N_18713,N_17474,N_17087);
xor U18714 (N_18714,N_17458,N_17586);
or U18715 (N_18715,N_17626,N_17722);
nand U18716 (N_18716,N_17335,N_17563);
nor U18717 (N_18717,N_17595,N_17539);
xnor U18718 (N_18718,N_17403,N_17438);
nand U18719 (N_18719,N_17457,N_17618);
nand U18720 (N_18720,N_17602,N_17711);
and U18721 (N_18721,N_17677,N_17442);
nand U18722 (N_18722,N_17088,N_17469);
xor U18723 (N_18723,N_17980,N_17956);
xnor U18724 (N_18724,N_17753,N_17530);
nor U18725 (N_18725,N_17075,N_17724);
xnor U18726 (N_18726,N_17130,N_17714);
xor U18727 (N_18727,N_17991,N_17235);
nand U18728 (N_18728,N_17870,N_17651);
xor U18729 (N_18729,N_17637,N_17367);
xor U18730 (N_18730,N_17124,N_17532);
or U18731 (N_18731,N_17516,N_17085);
nor U18732 (N_18732,N_17803,N_17446);
xor U18733 (N_18733,N_17894,N_17397);
xor U18734 (N_18734,N_17209,N_17821);
or U18735 (N_18735,N_17407,N_17323);
nand U18736 (N_18736,N_17999,N_17634);
xnor U18737 (N_18737,N_17024,N_17319);
and U18738 (N_18738,N_17188,N_17039);
and U18739 (N_18739,N_17480,N_17855);
nor U18740 (N_18740,N_17384,N_17110);
nor U18741 (N_18741,N_17787,N_17037);
or U18742 (N_18742,N_17350,N_17568);
nor U18743 (N_18743,N_17282,N_17338);
nand U18744 (N_18744,N_17667,N_17968);
nor U18745 (N_18745,N_17599,N_17753);
nor U18746 (N_18746,N_17229,N_17278);
xnor U18747 (N_18747,N_17132,N_17300);
or U18748 (N_18748,N_17800,N_17829);
nor U18749 (N_18749,N_17298,N_17818);
nand U18750 (N_18750,N_17337,N_17840);
nand U18751 (N_18751,N_17837,N_17673);
or U18752 (N_18752,N_17816,N_17039);
and U18753 (N_18753,N_17782,N_17563);
nand U18754 (N_18754,N_17701,N_17218);
nor U18755 (N_18755,N_17560,N_17094);
xnor U18756 (N_18756,N_17218,N_17952);
and U18757 (N_18757,N_17561,N_17928);
and U18758 (N_18758,N_17416,N_17854);
nand U18759 (N_18759,N_17693,N_17045);
xor U18760 (N_18760,N_17625,N_17578);
or U18761 (N_18761,N_17883,N_17662);
nor U18762 (N_18762,N_17537,N_17555);
and U18763 (N_18763,N_17977,N_17217);
xnor U18764 (N_18764,N_17140,N_17018);
nor U18765 (N_18765,N_17437,N_17568);
nand U18766 (N_18766,N_17334,N_17933);
and U18767 (N_18767,N_17823,N_17353);
nand U18768 (N_18768,N_17704,N_17885);
and U18769 (N_18769,N_17737,N_17105);
nand U18770 (N_18770,N_17532,N_17992);
xor U18771 (N_18771,N_17764,N_17526);
and U18772 (N_18772,N_17501,N_17219);
and U18773 (N_18773,N_17748,N_17067);
xnor U18774 (N_18774,N_17061,N_17032);
or U18775 (N_18775,N_17353,N_17114);
nor U18776 (N_18776,N_17265,N_17707);
nand U18777 (N_18777,N_17013,N_17385);
nand U18778 (N_18778,N_17253,N_17643);
nor U18779 (N_18779,N_17594,N_17281);
nor U18780 (N_18780,N_17229,N_17239);
nand U18781 (N_18781,N_17808,N_17355);
or U18782 (N_18782,N_17393,N_17821);
nor U18783 (N_18783,N_17423,N_17665);
nor U18784 (N_18784,N_17798,N_17953);
nor U18785 (N_18785,N_17553,N_17661);
nor U18786 (N_18786,N_17689,N_17613);
xnor U18787 (N_18787,N_17062,N_17262);
and U18788 (N_18788,N_17258,N_17511);
nand U18789 (N_18789,N_17411,N_17875);
nand U18790 (N_18790,N_17708,N_17854);
xnor U18791 (N_18791,N_17164,N_17787);
xnor U18792 (N_18792,N_17718,N_17862);
or U18793 (N_18793,N_17221,N_17082);
or U18794 (N_18794,N_17961,N_17478);
xor U18795 (N_18795,N_17793,N_17065);
nor U18796 (N_18796,N_17547,N_17208);
nor U18797 (N_18797,N_17231,N_17472);
nor U18798 (N_18798,N_17365,N_17606);
nand U18799 (N_18799,N_17328,N_17525);
or U18800 (N_18800,N_17618,N_17565);
nand U18801 (N_18801,N_17838,N_17457);
and U18802 (N_18802,N_17117,N_17112);
or U18803 (N_18803,N_17433,N_17523);
nand U18804 (N_18804,N_17585,N_17760);
and U18805 (N_18805,N_17056,N_17694);
nand U18806 (N_18806,N_17948,N_17615);
nor U18807 (N_18807,N_17466,N_17569);
or U18808 (N_18808,N_17611,N_17748);
and U18809 (N_18809,N_17625,N_17071);
nor U18810 (N_18810,N_17617,N_17870);
and U18811 (N_18811,N_17847,N_17068);
nand U18812 (N_18812,N_17119,N_17509);
nor U18813 (N_18813,N_17683,N_17458);
xor U18814 (N_18814,N_17968,N_17244);
xnor U18815 (N_18815,N_17220,N_17461);
nor U18816 (N_18816,N_17791,N_17983);
or U18817 (N_18817,N_17427,N_17594);
or U18818 (N_18818,N_17349,N_17070);
nor U18819 (N_18819,N_17017,N_17449);
and U18820 (N_18820,N_17459,N_17009);
xor U18821 (N_18821,N_17584,N_17109);
nor U18822 (N_18822,N_17927,N_17636);
xnor U18823 (N_18823,N_17349,N_17049);
nand U18824 (N_18824,N_17361,N_17295);
nand U18825 (N_18825,N_17955,N_17039);
nor U18826 (N_18826,N_17967,N_17284);
xor U18827 (N_18827,N_17942,N_17222);
nand U18828 (N_18828,N_17084,N_17377);
xor U18829 (N_18829,N_17079,N_17007);
or U18830 (N_18830,N_17649,N_17517);
or U18831 (N_18831,N_17315,N_17247);
or U18832 (N_18832,N_17821,N_17459);
nor U18833 (N_18833,N_17972,N_17860);
and U18834 (N_18834,N_17385,N_17791);
nand U18835 (N_18835,N_17557,N_17311);
nand U18836 (N_18836,N_17655,N_17834);
or U18837 (N_18837,N_17367,N_17418);
nand U18838 (N_18838,N_17240,N_17941);
or U18839 (N_18839,N_17848,N_17407);
nor U18840 (N_18840,N_17860,N_17029);
and U18841 (N_18841,N_17583,N_17340);
or U18842 (N_18842,N_17246,N_17906);
and U18843 (N_18843,N_17211,N_17432);
nand U18844 (N_18844,N_17442,N_17499);
or U18845 (N_18845,N_17715,N_17299);
or U18846 (N_18846,N_17058,N_17386);
xnor U18847 (N_18847,N_17984,N_17173);
nor U18848 (N_18848,N_17628,N_17297);
nand U18849 (N_18849,N_17885,N_17087);
nor U18850 (N_18850,N_17864,N_17665);
or U18851 (N_18851,N_17651,N_17714);
nor U18852 (N_18852,N_17658,N_17487);
and U18853 (N_18853,N_17470,N_17356);
nor U18854 (N_18854,N_17667,N_17224);
nor U18855 (N_18855,N_17361,N_17704);
xor U18856 (N_18856,N_17538,N_17312);
and U18857 (N_18857,N_17240,N_17301);
nor U18858 (N_18858,N_17319,N_17996);
and U18859 (N_18859,N_17988,N_17765);
xor U18860 (N_18860,N_17419,N_17144);
and U18861 (N_18861,N_17112,N_17640);
or U18862 (N_18862,N_17614,N_17560);
xnor U18863 (N_18863,N_17499,N_17662);
nor U18864 (N_18864,N_17366,N_17030);
nand U18865 (N_18865,N_17737,N_17860);
or U18866 (N_18866,N_17784,N_17257);
or U18867 (N_18867,N_17591,N_17629);
or U18868 (N_18868,N_17876,N_17565);
nor U18869 (N_18869,N_17990,N_17052);
xnor U18870 (N_18870,N_17661,N_17563);
nand U18871 (N_18871,N_17256,N_17957);
and U18872 (N_18872,N_17245,N_17680);
nor U18873 (N_18873,N_17819,N_17866);
nor U18874 (N_18874,N_17880,N_17085);
nor U18875 (N_18875,N_17795,N_17884);
nand U18876 (N_18876,N_17385,N_17123);
xnor U18877 (N_18877,N_17841,N_17286);
and U18878 (N_18878,N_17140,N_17203);
xnor U18879 (N_18879,N_17365,N_17309);
or U18880 (N_18880,N_17733,N_17443);
nand U18881 (N_18881,N_17874,N_17128);
xor U18882 (N_18882,N_17651,N_17685);
nor U18883 (N_18883,N_17473,N_17552);
or U18884 (N_18884,N_17565,N_17101);
and U18885 (N_18885,N_17648,N_17079);
or U18886 (N_18886,N_17602,N_17244);
xor U18887 (N_18887,N_17141,N_17954);
nor U18888 (N_18888,N_17766,N_17282);
or U18889 (N_18889,N_17937,N_17415);
and U18890 (N_18890,N_17775,N_17112);
or U18891 (N_18891,N_17310,N_17286);
or U18892 (N_18892,N_17203,N_17033);
and U18893 (N_18893,N_17910,N_17215);
nand U18894 (N_18894,N_17484,N_17595);
xnor U18895 (N_18895,N_17166,N_17862);
nor U18896 (N_18896,N_17846,N_17252);
nor U18897 (N_18897,N_17820,N_17688);
nor U18898 (N_18898,N_17889,N_17217);
nand U18899 (N_18899,N_17082,N_17919);
or U18900 (N_18900,N_17079,N_17681);
nand U18901 (N_18901,N_17721,N_17583);
and U18902 (N_18902,N_17534,N_17433);
and U18903 (N_18903,N_17285,N_17295);
xnor U18904 (N_18904,N_17644,N_17697);
nor U18905 (N_18905,N_17515,N_17183);
or U18906 (N_18906,N_17528,N_17777);
or U18907 (N_18907,N_17208,N_17224);
xnor U18908 (N_18908,N_17187,N_17059);
nor U18909 (N_18909,N_17476,N_17223);
and U18910 (N_18910,N_17097,N_17737);
xnor U18911 (N_18911,N_17051,N_17196);
or U18912 (N_18912,N_17516,N_17730);
and U18913 (N_18913,N_17407,N_17113);
nor U18914 (N_18914,N_17909,N_17341);
or U18915 (N_18915,N_17037,N_17821);
xnor U18916 (N_18916,N_17927,N_17238);
or U18917 (N_18917,N_17693,N_17487);
nor U18918 (N_18918,N_17943,N_17779);
nand U18919 (N_18919,N_17984,N_17840);
or U18920 (N_18920,N_17676,N_17840);
nor U18921 (N_18921,N_17344,N_17030);
or U18922 (N_18922,N_17225,N_17301);
nand U18923 (N_18923,N_17730,N_17506);
xnor U18924 (N_18924,N_17747,N_17009);
nor U18925 (N_18925,N_17635,N_17432);
or U18926 (N_18926,N_17397,N_17517);
xnor U18927 (N_18927,N_17874,N_17049);
xor U18928 (N_18928,N_17805,N_17397);
xnor U18929 (N_18929,N_17058,N_17472);
and U18930 (N_18930,N_17198,N_17951);
nand U18931 (N_18931,N_17311,N_17226);
or U18932 (N_18932,N_17877,N_17122);
nor U18933 (N_18933,N_17105,N_17550);
and U18934 (N_18934,N_17258,N_17551);
nand U18935 (N_18935,N_17714,N_17260);
xnor U18936 (N_18936,N_17026,N_17870);
nor U18937 (N_18937,N_17329,N_17978);
xor U18938 (N_18938,N_17981,N_17757);
xor U18939 (N_18939,N_17406,N_17157);
and U18940 (N_18940,N_17592,N_17750);
nor U18941 (N_18941,N_17157,N_17910);
and U18942 (N_18942,N_17037,N_17025);
xor U18943 (N_18943,N_17489,N_17553);
xnor U18944 (N_18944,N_17692,N_17288);
xnor U18945 (N_18945,N_17891,N_17419);
and U18946 (N_18946,N_17634,N_17296);
or U18947 (N_18947,N_17394,N_17378);
nor U18948 (N_18948,N_17147,N_17380);
nand U18949 (N_18949,N_17963,N_17991);
nor U18950 (N_18950,N_17990,N_17831);
or U18951 (N_18951,N_17914,N_17024);
nand U18952 (N_18952,N_17831,N_17753);
and U18953 (N_18953,N_17269,N_17239);
nor U18954 (N_18954,N_17336,N_17984);
nand U18955 (N_18955,N_17926,N_17801);
nand U18956 (N_18956,N_17983,N_17566);
and U18957 (N_18957,N_17476,N_17382);
xor U18958 (N_18958,N_17749,N_17955);
xor U18959 (N_18959,N_17106,N_17616);
or U18960 (N_18960,N_17338,N_17334);
and U18961 (N_18961,N_17569,N_17826);
xnor U18962 (N_18962,N_17115,N_17498);
nand U18963 (N_18963,N_17182,N_17958);
nand U18964 (N_18964,N_17787,N_17658);
nor U18965 (N_18965,N_17330,N_17948);
and U18966 (N_18966,N_17173,N_17331);
and U18967 (N_18967,N_17752,N_17143);
and U18968 (N_18968,N_17385,N_17186);
nand U18969 (N_18969,N_17326,N_17594);
nor U18970 (N_18970,N_17895,N_17100);
or U18971 (N_18971,N_17351,N_17497);
xor U18972 (N_18972,N_17287,N_17430);
nand U18973 (N_18973,N_17193,N_17213);
or U18974 (N_18974,N_17640,N_17964);
nand U18975 (N_18975,N_17745,N_17293);
nor U18976 (N_18976,N_17175,N_17923);
nor U18977 (N_18977,N_17353,N_17028);
or U18978 (N_18978,N_17925,N_17854);
or U18979 (N_18979,N_17057,N_17761);
and U18980 (N_18980,N_17228,N_17172);
and U18981 (N_18981,N_17006,N_17757);
or U18982 (N_18982,N_17181,N_17361);
xnor U18983 (N_18983,N_17647,N_17421);
nand U18984 (N_18984,N_17067,N_17357);
nand U18985 (N_18985,N_17758,N_17780);
and U18986 (N_18986,N_17676,N_17724);
and U18987 (N_18987,N_17344,N_17259);
and U18988 (N_18988,N_17273,N_17222);
xnor U18989 (N_18989,N_17220,N_17023);
nor U18990 (N_18990,N_17849,N_17601);
xor U18991 (N_18991,N_17915,N_17278);
nand U18992 (N_18992,N_17196,N_17133);
and U18993 (N_18993,N_17905,N_17023);
xnor U18994 (N_18994,N_17820,N_17599);
nor U18995 (N_18995,N_17999,N_17187);
and U18996 (N_18996,N_17258,N_17161);
nand U18997 (N_18997,N_17008,N_17970);
nand U18998 (N_18998,N_17852,N_17667);
nor U18999 (N_18999,N_17854,N_17933);
xnor U19000 (N_19000,N_18022,N_18760);
nor U19001 (N_19001,N_18783,N_18954);
and U19002 (N_19002,N_18270,N_18267);
or U19003 (N_19003,N_18136,N_18466);
nand U19004 (N_19004,N_18587,N_18142);
xor U19005 (N_19005,N_18151,N_18492);
nor U19006 (N_19006,N_18771,N_18586);
and U19007 (N_19007,N_18279,N_18105);
and U19008 (N_19008,N_18986,N_18851);
xnor U19009 (N_19009,N_18835,N_18653);
nor U19010 (N_19010,N_18538,N_18591);
or U19011 (N_19011,N_18614,N_18915);
nand U19012 (N_19012,N_18581,N_18950);
and U19013 (N_19013,N_18768,N_18541);
or U19014 (N_19014,N_18332,N_18134);
or U19015 (N_19015,N_18819,N_18159);
or U19016 (N_19016,N_18124,N_18359);
nand U19017 (N_19017,N_18589,N_18679);
nand U19018 (N_19018,N_18969,N_18504);
nor U19019 (N_19019,N_18035,N_18329);
or U19020 (N_19020,N_18420,N_18817);
or U19021 (N_19021,N_18601,N_18340);
and U19022 (N_19022,N_18953,N_18394);
nand U19023 (N_19023,N_18863,N_18114);
and U19024 (N_19024,N_18223,N_18312);
or U19025 (N_19025,N_18836,N_18021);
or U19026 (N_19026,N_18827,N_18038);
and U19027 (N_19027,N_18200,N_18757);
and U19028 (N_19028,N_18291,N_18445);
nor U19029 (N_19029,N_18413,N_18714);
xnor U19030 (N_19030,N_18040,N_18424);
nand U19031 (N_19031,N_18456,N_18422);
and U19032 (N_19032,N_18683,N_18684);
xnor U19033 (N_19033,N_18885,N_18864);
xnor U19034 (N_19034,N_18091,N_18749);
nor U19035 (N_19035,N_18288,N_18352);
nor U19036 (N_19036,N_18410,N_18814);
nor U19037 (N_19037,N_18918,N_18143);
nand U19038 (N_19038,N_18774,N_18753);
or U19039 (N_19039,N_18370,N_18898);
nand U19040 (N_19040,N_18547,N_18009);
or U19041 (N_19041,N_18917,N_18371);
or U19042 (N_19042,N_18227,N_18772);
or U19043 (N_19043,N_18050,N_18901);
nor U19044 (N_19044,N_18841,N_18952);
and U19045 (N_19045,N_18500,N_18657);
xor U19046 (N_19046,N_18938,N_18391);
nor U19047 (N_19047,N_18387,N_18701);
or U19048 (N_19048,N_18483,N_18164);
xnor U19049 (N_19049,N_18717,N_18568);
or U19050 (N_19050,N_18770,N_18028);
and U19051 (N_19051,N_18567,N_18113);
xor U19052 (N_19052,N_18201,N_18230);
nand U19053 (N_19053,N_18577,N_18221);
and U19054 (N_19054,N_18059,N_18758);
or U19055 (N_19055,N_18847,N_18033);
nor U19056 (N_19056,N_18795,N_18607);
or U19057 (N_19057,N_18365,N_18588);
or U19058 (N_19058,N_18425,N_18545);
and U19059 (N_19059,N_18026,N_18297);
xor U19060 (N_19060,N_18542,N_18752);
xor U19061 (N_19061,N_18349,N_18180);
nor U19062 (N_19062,N_18574,N_18934);
and U19063 (N_19063,N_18535,N_18482);
nand U19064 (N_19064,N_18584,N_18030);
and U19065 (N_19065,N_18183,N_18775);
nor U19066 (N_19066,N_18912,N_18552);
nand U19067 (N_19067,N_18186,N_18649);
xor U19068 (N_19068,N_18914,N_18132);
xnor U19069 (N_19069,N_18673,N_18549);
nor U19070 (N_19070,N_18636,N_18472);
xnor U19071 (N_19071,N_18735,N_18037);
or U19072 (N_19072,N_18002,N_18295);
and U19073 (N_19073,N_18039,N_18285);
nor U19074 (N_19074,N_18364,N_18590);
or U19075 (N_19075,N_18519,N_18633);
and U19076 (N_19076,N_18304,N_18503);
and U19077 (N_19077,N_18497,N_18958);
xnor U19078 (N_19078,N_18991,N_18632);
xor U19079 (N_19079,N_18119,N_18678);
nor U19080 (N_19080,N_18237,N_18651);
and U19081 (N_19081,N_18762,N_18518);
nand U19082 (N_19082,N_18869,N_18536);
nand U19083 (N_19083,N_18027,N_18874);
xor U19084 (N_19084,N_18910,N_18184);
nor U19085 (N_19085,N_18619,N_18427);
and U19086 (N_19086,N_18540,N_18489);
nor U19087 (N_19087,N_18993,N_18647);
and U19088 (N_19088,N_18036,N_18524);
nand U19089 (N_19089,N_18621,N_18166);
nand U19090 (N_19090,N_18508,N_18506);
nand U19091 (N_19091,N_18511,N_18094);
nor U19092 (N_19092,N_18306,N_18389);
nand U19093 (N_19093,N_18487,N_18463);
nor U19094 (N_19094,N_18592,N_18362);
nor U19095 (N_19095,N_18579,N_18961);
xor U19096 (N_19096,N_18544,N_18996);
nand U19097 (N_19097,N_18974,N_18693);
nand U19098 (N_19098,N_18216,N_18404);
nor U19099 (N_19099,N_18913,N_18060);
or U19100 (N_19100,N_18942,N_18725);
xnor U19101 (N_19101,N_18686,N_18698);
and U19102 (N_19102,N_18010,N_18502);
nand U19103 (N_19103,N_18069,N_18606);
or U19104 (N_19104,N_18255,N_18431);
xor U19105 (N_19105,N_18555,N_18571);
nor U19106 (N_19106,N_18870,N_18242);
nor U19107 (N_19107,N_18397,N_18287);
nand U19108 (N_19108,N_18900,N_18711);
xnor U19109 (N_19109,N_18575,N_18042);
nor U19110 (N_19110,N_18104,N_18944);
or U19111 (N_19111,N_18298,N_18469);
or U19112 (N_19112,N_18258,N_18997);
nand U19113 (N_19113,N_18560,N_18945);
nand U19114 (N_19114,N_18564,N_18802);
and U19115 (N_19115,N_18246,N_18266);
and U19116 (N_19116,N_18602,N_18087);
xor U19117 (N_19117,N_18219,N_18943);
nor U19118 (N_19118,N_18350,N_18970);
xor U19119 (N_19119,N_18321,N_18562);
xor U19120 (N_19120,N_18994,N_18058);
and U19121 (N_19121,N_18973,N_18732);
xor U19122 (N_19122,N_18576,N_18401);
and U19123 (N_19123,N_18068,N_18737);
nand U19124 (N_19124,N_18680,N_18799);
nand U19125 (N_19125,N_18062,N_18889);
or U19126 (N_19126,N_18435,N_18800);
xnor U19127 (N_19127,N_18608,N_18721);
xnor U19128 (N_19128,N_18357,N_18224);
or U19129 (N_19129,N_18176,N_18729);
nor U19130 (N_19130,N_18556,N_18850);
nor U19131 (N_19131,N_18369,N_18065);
xor U19132 (N_19132,N_18667,N_18446);
nand U19133 (N_19133,N_18959,N_18668);
and U19134 (N_19134,N_18672,N_18139);
and U19135 (N_19135,N_18355,N_18655);
nor U19136 (N_19136,N_18890,N_18479);
xnor U19137 (N_19137,N_18470,N_18376);
nor U19138 (N_19138,N_18951,N_18380);
xor U19139 (N_19139,N_18292,N_18832);
and U19140 (N_19140,N_18498,N_18311);
or U19141 (N_19141,N_18894,N_18939);
and U19142 (N_19142,N_18765,N_18141);
or U19143 (N_19143,N_18326,N_18543);
nor U19144 (N_19144,N_18165,N_18043);
or U19145 (N_19145,N_18891,N_18353);
and U19146 (N_19146,N_18595,N_18766);
nor U19147 (N_19147,N_18083,N_18756);
xnor U19148 (N_19148,N_18175,N_18848);
nor U19149 (N_19149,N_18379,N_18190);
or U19150 (N_19150,N_18341,N_18310);
nor U19151 (N_19151,N_18513,N_18787);
and U19152 (N_19152,N_18599,N_18550);
xor U19153 (N_19153,N_18514,N_18532);
xnor U19154 (N_19154,N_18722,N_18031);
nand U19155 (N_19155,N_18642,N_18099);
nor U19156 (N_19156,N_18408,N_18229);
and U19157 (N_19157,N_18855,N_18853);
or U19158 (N_19158,N_18337,N_18813);
and U19159 (N_19159,N_18692,N_18648);
nor U19160 (N_19160,N_18277,N_18273);
or U19161 (N_19161,N_18989,N_18797);
or U19162 (N_19162,N_18925,N_18570);
nor U19163 (N_19163,N_18899,N_18073);
nand U19164 (N_19164,N_18202,N_18727);
nand U19165 (N_19165,N_18972,N_18041);
or U19166 (N_19166,N_18691,N_18730);
or U19167 (N_19167,N_18769,N_18845);
xor U19168 (N_19168,N_18309,N_18486);
and U19169 (N_19169,N_18481,N_18826);
nor U19170 (N_19170,N_18107,N_18919);
nand U19171 (N_19171,N_18409,N_18381);
or U19172 (N_19172,N_18613,N_18459);
nor U19173 (N_19173,N_18063,N_18904);
or U19174 (N_19174,N_18070,N_18325);
or U19175 (N_19175,N_18017,N_18286);
xnor U19176 (N_19176,N_18654,N_18145);
and U19177 (N_19177,N_18171,N_18215);
nand U19178 (N_19178,N_18331,N_18897);
xor U19179 (N_19179,N_18854,N_18212);
or U19180 (N_19180,N_18861,N_18748);
nor U19181 (N_19181,N_18004,N_18741);
and U19182 (N_19182,N_18324,N_18111);
and U19183 (N_19183,N_18363,N_18982);
or U19184 (N_19184,N_18308,N_18206);
nand U19185 (N_19185,N_18617,N_18024);
nor U19186 (N_19186,N_18108,N_18816);
nor U19187 (N_19187,N_18218,N_18034);
or U19188 (N_19188,N_18690,N_18429);
nand U19189 (N_19189,N_18937,N_18930);
nor U19190 (N_19190,N_18936,N_18128);
nand U19191 (N_19191,N_18534,N_18366);
nand U19192 (N_19192,N_18669,N_18208);
xor U19193 (N_19193,N_18493,N_18053);
and U19194 (N_19194,N_18434,N_18020);
xnor U19195 (N_19195,N_18232,N_18811);
xnor U19196 (N_19196,N_18097,N_18947);
nor U19197 (N_19197,N_18720,N_18101);
xnor U19198 (N_19198,N_18477,N_18174);
nor U19199 (N_19199,N_18763,N_18578);
nor U19200 (N_19200,N_18987,N_18923);
nand U19201 (N_19201,N_18249,N_18138);
and U19202 (N_19202,N_18345,N_18666);
or U19203 (N_19203,N_18928,N_18228);
nand U19204 (N_19204,N_18779,N_18383);
and U19205 (N_19205,N_18801,N_18551);
xor U19206 (N_19206,N_18728,N_18988);
or U19207 (N_19207,N_18054,N_18150);
or U19208 (N_19208,N_18857,N_18029);
or U19209 (N_19209,N_18344,N_18932);
and U19210 (N_19210,N_18005,N_18110);
nor U19211 (N_19211,N_18077,N_18135);
nand U19212 (N_19212,N_18018,N_18156);
nand U19213 (N_19213,N_18628,N_18985);
or U19214 (N_19214,N_18032,N_18315);
nand U19215 (N_19215,N_18072,N_18396);
nor U19216 (N_19216,N_18886,N_18259);
or U19217 (N_19217,N_18240,N_18265);
nor U19218 (N_19218,N_18565,N_18731);
nand U19219 (N_19219,N_18182,N_18906);
or U19220 (N_19220,N_18745,N_18983);
nand U19221 (N_19221,N_18011,N_18131);
xnor U19222 (N_19222,N_18301,N_18006);
nor U19223 (N_19223,N_18643,N_18903);
nand U19224 (N_19224,N_18168,N_18746);
and U19225 (N_19225,N_18630,N_18374);
nand U19226 (N_19226,N_18645,N_18457);
xor U19227 (N_19227,N_18251,N_18780);
nand U19228 (N_19228,N_18843,N_18755);
xnor U19229 (N_19229,N_18529,N_18708);
and U19230 (N_19230,N_18603,N_18622);
nand U19231 (N_19231,N_18276,N_18441);
nand U19232 (N_19232,N_18924,N_18220);
nand U19233 (N_19233,N_18406,N_18262);
nand U19234 (N_19234,N_18226,N_18979);
or U19235 (N_19235,N_18715,N_18467);
xor U19236 (N_19236,N_18172,N_18000);
or U19237 (N_19237,N_18257,N_18663);
or U19238 (N_19238,N_18407,N_18794);
nand U19239 (N_19239,N_18878,N_18393);
nor U19240 (N_19240,N_18554,N_18275);
or U19241 (N_19241,N_18382,N_18144);
xor U19242 (N_19242,N_18523,N_18754);
or U19243 (N_19243,N_18193,N_18594);
and U19244 (N_19244,N_18882,N_18573);
nor U19245 (N_19245,N_18507,N_18810);
nand U19246 (N_19246,N_18888,N_18759);
or U19247 (N_19247,N_18634,N_18675);
nand U19248 (N_19248,N_18335,N_18373);
nand U19249 (N_19249,N_18744,N_18834);
xnor U19250 (N_19250,N_18839,N_18207);
or U19251 (N_19251,N_18956,N_18596);
nor U19252 (N_19252,N_18883,N_18313);
or U19253 (N_19253,N_18557,N_18079);
xor U19254 (N_19254,N_18328,N_18076);
and U19255 (N_19255,N_18402,N_18471);
xor U19256 (N_19256,N_18405,N_18210);
xnor U19257 (N_19257,N_18868,N_18751);
xnor U19258 (N_19258,N_18147,N_18282);
or U19259 (N_19259,N_18008,N_18118);
or U19260 (N_19260,N_18490,N_18742);
or U19261 (N_19261,N_18616,N_18615);
or U19262 (N_19262,N_18347,N_18303);
or U19263 (N_19263,N_18048,N_18090);
and U19264 (N_19264,N_18222,N_18955);
or U19265 (N_19265,N_18239,N_18430);
xnor U19266 (N_19266,N_18305,N_18085);
xnor U19267 (N_19267,N_18170,N_18509);
nand U19268 (N_19268,N_18322,N_18788);
xnor U19269 (N_19269,N_18399,N_18887);
or U19270 (N_19270,N_18892,N_18895);
nor U19271 (N_19271,N_18314,N_18271);
nor U19272 (N_19272,N_18699,N_18248);
or U19273 (N_19273,N_18908,N_18747);
and U19274 (N_19274,N_18706,N_18450);
and U19275 (N_19275,N_18294,N_18921);
xnor U19276 (N_19276,N_18436,N_18244);
nand U19277 (N_19277,N_18044,N_18181);
or U19278 (N_19278,N_18962,N_18637);
and U19279 (N_19279,N_18558,N_18103);
nand U19280 (N_19280,N_18197,N_18999);
nand U19281 (N_19281,N_18515,N_18533);
nor U19282 (N_19282,N_18656,N_18019);
xnor U19283 (N_19283,N_18821,N_18474);
nand U19284 (N_19284,N_18454,N_18157);
xor U19285 (N_19285,N_18449,N_18652);
nor U19286 (N_19286,N_18149,N_18583);
and U19287 (N_19287,N_18437,N_18546);
and U19288 (N_19288,N_18612,N_18896);
xor U19289 (N_19289,N_18920,N_18278);
or U19290 (N_19290,N_18316,N_18968);
nand U19291 (N_19291,N_18078,N_18433);
and U19292 (N_19292,N_18859,N_18528);
nand U19293 (N_19293,N_18231,N_18569);
nand U19294 (N_19294,N_18750,N_18499);
nand U19295 (N_19295,N_18235,N_18724);
xor U19296 (N_19296,N_18225,N_18116);
nor U19297 (N_19297,N_18719,N_18163);
and U19298 (N_19298,N_18392,N_18179);
or U19299 (N_19299,N_18440,N_18833);
nand U19300 (N_19300,N_18452,N_18385);
nand U19301 (N_19301,N_18709,N_18274);
or U19302 (N_19302,N_18929,N_18842);
and U19303 (N_19303,N_18075,N_18354);
and U19304 (N_19304,N_18761,N_18453);
nor U19305 (N_19305,N_18548,N_18014);
xor U19306 (N_19306,N_18460,N_18488);
nor U19307 (N_19307,N_18395,N_18432);
or U19308 (N_19308,N_18782,N_18264);
and U19309 (N_19309,N_18290,N_18776);
and U19310 (N_19310,N_18377,N_18162);
or U19311 (N_19311,N_18773,N_18192);
or U19312 (N_19312,N_18798,N_18214);
or U19313 (N_19313,N_18803,N_18112);
nand U19314 (N_19314,N_18153,N_18705);
or U19315 (N_19315,N_18003,N_18967);
and U19316 (N_19316,N_18946,N_18473);
nand U19317 (N_19317,N_18080,N_18674);
nand U19318 (N_19318,N_18280,N_18137);
and U19319 (N_19319,N_18049,N_18926);
xnor U19320 (N_19320,N_18100,N_18444);
xor U19321 (N_19321,N_18209,N_18935);
or U19322 (N_19322,N_18261,N_18236);
or U19323 (N_19323,N_18458,N_18978);
or U19324 (N_19324,N_18815,N_18057);
xnor U19325 (N_19325,N_18629,N_18263);
and U19326 (N_19326,N_18609,N_18677);
or U19327 (N_19327,N_18023,N_18501);
nand U19328 (N_19328,N_18443,N_18611);
nor U19329 (N_19329,N_18188,N_18269);
nor U19330 (N_19330,N_18786,N_18696);
or U19331 (N_19331,N_18792,N_18013);
nor U19332 (N_19332,N_18793,N_18343);
or U19333 (N_19333,N_18922,N_18965);
and U19334 (N_19334,N_18293,N_18161);
or U19335 (N_19335,N_18241,N_18423);
nand U19336 (N_19336,N_18525,N_18082);
nand U19337 (N_19337,N_18644,N_18846);
nand U19338 (N_19338,N_18253,N_18909);
nor U19339 (N_19339,N_18734,N_18778);
xnor U19340 (N_19340,N_18860,N_18152);
xnor U19341 (N_19341,N_18957,N_18703);
nor U19342 (N_19342,N_18123,N_18484);
and U19343 (N_19343,N_18015,N_18169);
xor U19344 (N_19344,N_18320,N_18876);
and U19345 (N_19345,N_18877,N_18120);
nand U19346 (N_19346,N_18537,N_18398);
or U19347 (N_19347,N_18185,N_18372);
xnor U19348 (N_19348,N_18866,N_18055);
or U19349 (N_19349,N_18299,N_18710);
nor U19350 (N_19350,N_18415,N_18884);
nor U19351 (N_19351,N_18593,N_18966);
and U19352 (N_19352,N_18512,N_18805);
xnor U19353 (N_19353,N_18098,N_18386);
nand U19354 (N_19354,N_18976,N_18007);
or U19355 (N_19355,N_18739,N_18117);
xor U19356 (N_19356,N_18071,N_18155);
and U19357 (N_19357,N_18300,N_18659);
xor U19358 (N_19358,N_18808,N_18646);
xnor U19359 (N_19359,N_18238,N_18283);
xor U19360 (N_19360,N_18245,N_18442);
or U19361 (N_19361,N_18358,N_18167);
xor U19362 (N_19362,N_18317,N_18016);
and U19363 (N_19363,N_18384,N_18284);
or U19364 (N_19364,N_18960,N_18476);
nor U19365 (N_19365,N_18880,N_18624);
nor U19366 (N_19366,N_18940,N_18566);
and U19367 (N_19367,N_18045,N_18411);
xor U19368 (N_19368,N_18812,N_18893);
xor U19369 (N_19369,N_18682,N_18738);
or U19370 (N_19370,N_18820,N_18635);
nor U19371 (N_19371,N_18638,N_18256);
nor U19372 (N_19372,N_18559,N_18582);
xor U19373 (N_19373,N_18658,N_18639);
nand U19374 (N_19374,N_18995,N_18418);
or U19375 (N_19375,N_18640,N_18605);
or U19376 (N_19376,N_18133,N_18205);
xnor U19377 (N_19377,N_18378,N_18233);
and U19378 (N_19378,N_18074,N_18676);
xor U19379 (N_19379,N_18109,N_18234);
and U19380 (N_19380,N_18339,N_18419);
xnor U19381 (N_19381,N_18522,N_18585);
xor U19382 (N_19382,N_18828,N_18412);
and U19383 (N_19383,N_18189,N_18531);
and U19384 (N_19384,N_18849,N_18367);
or U19385 (N_19385,N_18281,N_18681);
nand U19386 (N_19386,N_18464,N_18822);
or U19387 (N_19387,N_18178,N_18081);
or U19388 (N_19388,N_18825,N_18650);
xnor U19389 (N_19389,N_18361,N_18356);
and U19390 (N_19390,N_18852,N_18390);
nor U19391 (N_19391,N_18796,N_18348);
and U19392 (N_19392,N_18302,N_18563);
and U19393 (N_19393,N_18689,N_18902);
and U19394 (N_19394,N_18623,N_18809);
nand U19395 (N_19395,N_18907,N_18338);
or U19396 (N_19396,N_18421,N_18056);
nand U19397 (N_19397,N_18086,N_18336);
or U19398 (N_19398,N_18992,N_18191);
nor U19399 (N_19399,N_18521,N_18610);
nor U19400 (N_19400,N_18671,N_18140);
and U19401 (N_19401,N_18767,N_18712);
xnor U19402 (N_19402,N_18046,N_18095);
xnor U19403 (N_19403,N_18704,N_18867);
or U19404 (N_19404,N_18084,N_18130);
nor U19405 (N_19405,N_18881,N_18478);
or U19406 (N_19406,N_18243,N_18831);
nor U19407 (N_19407,N_18451,N_18102);
xor U19408 (N_19408,N_18516,N_18187);
and U19409 (N_19409,N_18438,N_18426);
xor U19410 (N_19410,N_18334,N_18905);
and U19411 (N_19411,N_18873,N_18631);
or U19412 (N_19412,N_18495,N_18530);
nand U19413 (N_19413,N_18247,N_18428);
xnor U19414 (N_19414,N_18949,N_18790);
nor U19415 (N_19415,N_18252,N_18199);
nor U19416 (N_19416,N_18480,N_18777);
or U19417 (N_19417,N_18439,N_18665);
nand U19418 (N_19418,N_18620,N_18597);
nor U19419 (N_19419,N_18148,N_18700);
nor U19420 (N_19420,N_18447,N_18670);
nor U19421 (N_19421,N_18414,N_18333);
and U19422 (N_19422,N_18177,N_18475);
or U19423 (N_19423,N_18781,N_18468);
and U19424 (N_19424,N_18115,N_18198);
nor U19425 (N_19425,N_18088,N_18211);
or U19426 (N_19426,N_18598,N_18001);
nor U19427 (N_19427,N_18375,N_18448);
or U19428 (N_19428,N_18726,N_18526);
nand U19429 (N_19429,N_18051,N_18862);
and U19430 (N_19430,N_18695,N_18260);
nand U19431 (N_19431,N_18204,N_18342);
and U19432 (N_19432,N_18580,N_18911);
or U19433 (N_19433,N_18510,N_18461);
and U19434 (N_19434,N_18661,N_18688);
or U19435 (N_19435,N_18417,N_18064);
nand U19436 (N_19436,N_18254,N_18600);
xnor U19437 (N_19437,N_18804,N_18268);
xor U19438 (N_19438,N_18203,N_18660);
nor U19439 (N_19439,N_18685,N_18980);
xor U19440 (N_19440,N_18927,N_18289);
nor U19441 (N_19441,N_18830,N_18664);
xor U19442 (N_19442,N_18158,N_18733);
or U19443 (N_19443,N_18604,N_18694);
nor U19444 (N_19444,N_18572,N_18485);
nor U19445 (N_19445,N_18527,N_18807);
nand U19446 (N_19446,N_18879,N_18916);
and U19447 (N_19447,N_18875,N_18194);
and U19448 (N_19448,N_18403,N_18307);
or U19449 (N_19449,N_18723,N_18327);
or U19450 (N_19450,N_18092,N_18195);
or U19451 (N_19451,N_18626,N_18948);
or U19452 (N_19452,N_18618,N_18494);
or U19453 (N_19453,N_18840,N_18837);
and U19454 (N_19454,N_18963,N_18121);
and U19455 (N_19455,N_18561,N_18368);
or U19456 (N_19456,N_18089,N_18296);
xnor U19457 (N_19457,N_18641,N_18872);
nand U19458 (N_19458,N_18743,N_18196);
nand U19459 (N_19459,N_18146,N_18539);
or U19460 (N_19460,N_18697,N_18520);
nand U19461 (N_19461,N_18791,N_18818);
and U19462 (N_19462,N_18272,N_18217);
nor U19463 (N_19463,N_18122,N_18553);
xnor U19464 (N_19464,N_18971,N_18127);
nor U19465 (N_19465,N_18844,N_18129);
nor U19466 (N_19466,N_18096,N_18388);
nor U19467 (N_19467,N_18871,N_18707);
nor U19468 (N_19468,N_18455,N_18990);
or U19469 (N_19469,N_18465,N_18625);
or U19470 (N_19470,N_18318,N_18323);
nand U19471 (N_19471,N_18789,N_18856);
or U19472 (N_19472,N_18806,N_18319);
xor U19473 (N_19473,N_18662,N_18823);
xnor U19474 (N_19474,N_18931,N_18066);
or U19475 (N_19475,N_18824,N_18160);
or U19476 (N_19476,N_18462,N_18491);
nand U19477 (N_19477,N_18975,N_18067);
nand U19478 (N_19478,N_18829,N_18740);
nand U19479 (N_19479,N_18764,N_18346);
and U19480 (N_19480,N_18865,N_18173);
and U19481 (N_19481,N_18702,N_18998);
xnor U19482 (N_19482,N_18351,N_18784);
nor U19483 (N_19483,N_18416,N_18977);
or U19484 (N_19484,N_18106,N_18858);
nor U19485 (N_19485,N_18330,N_18517);
nor U19486 (N_19486,N_18047,N_18984);
and U19487 (N_19487,N_18941,N_18933);
nand U19488 (N_19488,N_18716,N_18838);
xnor U19489 (N_19489,N_18025,N_18213);
xnor U19490 (N_19490,N_18713,N_18718);
nor U19491 (N_19491,N_18360,N_18981);
and U19492 (N_19492,N_18400,N_18125);
xnor U19493 (N_19493,N_18627,N_18061);
xor U19494 (N_19494,N_18250,N_18736);
xor U19495 (N_19495,N_18505,N_18687);
or U19496 (N_19496,N_18052,N_18012);
xor U19497 (N_19497,N_18964,N_18154);
or U19498 (N_19498,N_18093,N_18785);
nor U19499 (N_19499,N_18496,N_18126);
nand U19500 (N_19500,N_18006,N_18286);
nand U19501 (N_19501,N_18307,N_18037);
nor U19502 (N_19502,N_18359,N_18295);
or U19503 (N_19503,N_18046,N_18197);
nand U19504 (N_19504,N_18512,N_18589);
or U19505 (N_19505,N_18666,N_18573);
xnor U19506 (N_19506,N_18175,N_18056);
and U19507 (N_19507,N_18768,N_18225);
nor U19508 (N_19508,N_18258,N_18292);
or U19509 (N_19509,N_18100,N_18077);
and U19510 (N_19510,N_18000,N_18047);
xnor U19511 (N_19511,N_18897,N_18286);
xor U19512 (N_19512,N_18524,N_18682);
or U19513 (N_19513,N_18005,N_18114);
nor U19514 (N_19514,N_18446,N_18764);
or U19515 (N_19515,N_18988,N_18080);
nor U19516 (N_19516,N_18708,N_18824);
or U19517 (N_19517,N_18335,N_18273);
nand U19518 (N_19518,N_18340,N_18878);
nand U19519 (N_19519,N_18671,N_18476);
nor U19520 (N_19520,N_18829,N_18887);
and U19521 (N_19521,N_18221,N_18761);
and U19522 (N_19522,N_18291,N_18223);
and U19523 (N_19523,N_18226,N_18738);
or U19524 (N_19524,N_18346,N_18062);
or U19525 (N_19525,N_18429,N_18906);
xor U19526 (N_19526,N_18645,N_18065);
nand U19527 (N_19527,N_18736,N_18310);
nand U19528 (N_19528,N_18964,N_18329);
nor U19529 (N_19529,N_18935,N_18433);
nand U19530 (N_19530,N_18337,N_18468);
nand U19531 (N_19531,N_18625,N_18440);
or U19532 (N_19532,N_18611,N_18809);
xor U19533 (N_19533,N_18618,N_18046);
and U19534 (N_19534,N_18805,N_18711);
xnor U19535 (N_19535,N_18954,N_18583);
or U19536 (N_19536,N_18959,N_18004);
or U19537 (N_19537,N_18427,N_18011);
xnor U19538 (N_19538,N_18930,N_18266);
and U19539 (N_19539,N_18116,N_18505);
nand U19540 (N_19540,N_18570,N_18066);
nand U19541 (N_19541,N_18579,N_18044);
nor U19542 (N_19542,N_18179,N_18317);
and U19543 (N_19543,N_18253,N_18823);
nand U19544 (N_19544,N_18422,N_18228);
or U19545 (N_19545,N_18265,N_18628);
and U19546 (N_19546,N_18509,N_18867);
or U19547 (N_19547,N_18545,N_18138);
xor U19548 (N_19548,N_18607,N_18126);
nor U19549 (N_19549,N_18494,N_18154);
nor U19550 (N_19550,N_18680,N_18727);
nand U19551 (N_19551,N_18559,N_18049);
xor U19552 (N_19552,N_18779,N_18359);
nand U19553 (N_19553,N_18318,N_18833);
and U19554 (N_19554,N_18496,N_18566);
or U19555 (N_19555,N_18105,N_18146);
and U19556 (N_19556,N_18306,N_18455);
nor U19557 (N_19557,N_18081,N_18330);
or U19558 (N_19558,N_18805,N_18027);
nor U19559 (N_19559,N_18620,N_18549);
or U19560 (N_19560,N_18570,N_18712);
nor U19561 (N_19561,N_18737,N_18809);
nand U19562 (N_19562,N_18638,N_18027);
xnor U19563 (N_19563,N_18690,N_18496);
nand U19564 (N_19564,N_18052,N_18907);
xnor U19565 (N_19565,N_18223,N_18533);
or U19566 (N_19566,N_18038,N_18133);
nor U19567 (N_19567,N_18321,N_18306);
nor U19568 (N_19568,N_18271,N_18741);
nor U19569 (N_19569,N_18391,N_18348);
or U19570 (N_19570,N_18898,N_18990);
nand U19571 (N_19571,N_18692,N_18946);
or U19572 (N_19572,N_18203,N_18475);
or U19573 (N_19573,N_18429,N_18126);
xnor U19574 (N_19574,N_18164,N_18871);
and U19575 (N_19575,N_18173,N_18524);
xnor U19576 (N_19576,N_18151,N_18400);
nand U19577 (N_19577,N_18483,N_18608);
or U19578 (N_19578,N_18705,N_18495);
nand U19579 (N_19579,N_18987,N_18476);
and U19580 (N_19580,N_18537,N_18676);
or U19581 (N_19581,N_18730,N_18624);
xor U19582 (N_19582,N_18592,N_18184);
or U19583 (N_19583,N_18382,N_18067);
and U19584 (N_19584,N_18137,N_18604);
nand U19585 (N_19585,N_18767,N_18454);
xnor U19586 (N_19586,N_18094,N_18075);
or U19587 (N_19587,N_18158,N_18026);
or U19588 (N_19588,N_18319,N_18428);
nand U19589 (N_19589,N_18489,N_18913);
xnor U19590 (N_19590,N_18073,N_18589);
xor U19591 (N_19591,N_18624,N_18248);
nor U19592 (N_19592,N_18395,N_18462);
nand U19593 (N_19593,N_18540,N_18754);
xor U19594 (N_19594,N_18823,N_18319);
nor U19595 (N_19595,N_18677,N_18807);
and U19596 (N_19596,N_18121,N_18896);
nor U19597 (N_19597,N_18036,N_18278);
nand U19598 (N_19598,N_18717,N_18948);
xnor U19599 (N_19599,N_18192,N_18523);
and U19600 (N_19600,N_18865,N_18127);
nor U19601 (N_19601,N_18885,N_18329);
nor U19602 (N_19602,N_18815,N_18547);
nor U19603 (N_19603,N_18080,N_18551);
or U19604 (N_19604,N_18823,N_18365);
nand U19605 (N_19605,N_18091,N_18146);
xor U19606 (N_19606,N_18406,N_18065);
nor U19607 (N_19607,N_18256,N_18143);
nor U19608 (N_19608,N_18569,N_18435);
xor U19609 (N_19609,N_18977,N_18187);
and U19610 (N_19610,N_18153,N_18337);
nand U19611 (N_19611,N_18985,N_18614);
nor U19612 (N_19612,N_18596,N_18120);
xor U19613 (N_19613,N_18031,N_18836);
or U19614 (N_19614,N_18762,N_18027);
nor U19615 (N_19615,N_18910,N_18070);
nor U19616 (N_19616,N_18842,N_18830);
nand U19617 (N_19617,N_18340,N_18921);
nand U19618 (N_19618,N_18860,N_18666);
and U19619 (N_19619,N_18919,N_18394);
nor U19620 (N_19620,N_18162,N_18303);
xnor U19621 (N_19621,N_18423,N_18704);
nand U19622 (N_19622,N_18654,N_18333);
nand U19623 (N_19623,N_18224,N_18251);
or U19624 (N_19624,N_18599,N_18184);
nor U19625 (N_19625,N_18391,N_18387);
nor U19626 (N_19626,N_18303,N_18170);
and U19627 (N_19627,N_18238,N_18368);
nor U19628 (N_19628,N_18673,N_18859);
xor U19629 (N_19629,N_18333,N_18556);
or U19630 (N_19630,N_18731,N_18222);
and U19631 (N_19631,N_18571,N_18077);
and U19632 (N_19632,N_18540,N_18938);
nor U19633 (N_19633,N_18692,N_18339);
xor U19634 (N_19634,N_18056,N_18128);
or U19635 (N_19635,N_18867,N_18841);
or U19636 (N_19636,N_18897,N_18204);
xor U19637 (N_19637,N_18743,N_18426);
nand U19638 (N_19638,N_18302,N_18623);
or U19639 (N_19639,N_18034,N_18287);
nor U19640 (N_19640,N_18248,N_18992);
nor U19641 (N_19641,N_18548,N_18407);
nor U19642 (N_19642,N_18586,N_18490);
and U19643 (N_19643,N_18539,N_18007);
and U19644 (N_19644,N_18711,N_18176);
nor U19645 (N_19645,N_18770,N_18855);
and U19646 (N_19646,N_18257,N_18291);
nand U19647 (N_19647,N_18448,N_18502);
or U19648 (N_19648,N_18125,N_18559);
nor U19649 (N_19649,N_18203,N_18854);
or U19650 (N_19650,N_18945,N_18368);
nand U19651 (N_19651,N_18051,N_18513);
nand U19652 (N_19652,N_18259,N_18906);
and U19653 (N_19653,N_18085,N_18096);
nor U19654 (N_19654,N_18139,N_18143);
xnor U19655 (N_19655,N_18119,N_18459);
and U19656 (N_19656,N_18669,N_18239);
nor U19657 (N_19657,N_18346,N_18160);
or U19658 (N_19658,N_18164,N_18213);
xor U19659 (N_19659,N_18285,N_18213);
nor U19660 (N_19660,N_18019,N_18295);
nor U19661 (N_19661,N_18937,N_18398);
and U19662 (N_19662,N_18151,N_18214);
and U19663 (N_19663,N_18931,N_18371);
nor U19664 (N_19664,N_18721,N_18088);
xor U19665 (N_19665,N_18056,N_18790);
and U19666 (N_19666,N_18636,N_18657);
or U19667 (N_19667,N_18490,N_18020);
or U19668 (N_19668,N_18736,N_18822);
or U19669 (N_19669,N_18447,N_18842);
or U19670 (N_19670,N_18740,N_18953);
nand U19671 (N_19671,N_18244,N_18441);
nand U19672 (N_19672,N_18981,N_18432);
nand U19673 (N_19673,N_18047,N_18645);
nand U19674 (N_19674,N_18925,N_18425);
or U19675 (N_19675,N_18743,N_18282);
xor U19676 (N_19676,N_18933,N_18151);
xnor U19677 (N_19677,N_18404,N_18068);
nand U19678 (N_19678,N_18006,N_18750);
and U19679 (N_19679,N_18247,N_18345);
xnor U19680 (N_19680,N_18396,N_18171);
xor U19681 (N_19681,N_18532,N_18245);
nor U19682 (N_19682,N_18316,N_18697);
nand U19683 (N_19683,N_18893,N_18972);
or U19684 (N_19684,N_18611,N_18297);
or U19685 (N_19685,N_18833,N_18087);
xor U19686 (N_19686,N_18661,N_18735);
and U19687 (N_19687,N_18130,N_18906);
xor U19688 (N_19688,N_18881,N_18295);
nor U19689 (N_19689,N_18476,N_18596);
nand U19690 (N_19690,N_18045,N_18829);
nand U19691 (N_19691,N_18201,N_18273);
or U19692 (N_19692,N_18904,N_18622);
xnor U19693 (N_19693,N_18059,N_18102);
xnor U19694 (N_19694,N_18824,N_18745);
xor U19695 (N_19695,N_18271,N_18454);
xnor U19696 (N_19696,N_18012,N_18992);
nor U19697 (N_19697,N_18145,N_18645);
and U19698 (N_19698,N_18290,N_18929);
nand U19699 (N_19699,N_18276,N_18246);
or U19700 (N_19700,N_18992,N_18051);
nor U19701 (N_19701,N_18272,N_18369);
nor U19702 (N_19702,N_18186,N_18578);
xor U19703 (N_19703,N_18646,N_18762);
or U19704 (N_19704,N_18675,N_18039);
and U19705 (N_19705,N_18164,N_18466);
or U19706 (N_19706,N_18744,N_18167);
or U19707 (N_19707,N_18695,N_18489);
nand U19708 (N_19708,N_18017,N_18714);
nand U19709 (N_19709,N_18882,N_18901);
nor U19710 (N_19710,N_18632,N_18198);
nand U19711 (N_19711,N_18927,N_18075);
or U19712 (N_19712,N_18271,N_18650);
nand U19713 (N_19713,N_18777,N_18679);
nand U19714 (N_19714,N_18779,N_18284);
nand U19715 (N_19715,N_18216,N_18864);
xor U19716 (N_19716,N_18413,N_18985);
or U19717 (N_19717,N_18057,N_18126);
or U19718 (N_19718,N_18370,N_18219);
or U19719 (N_19719,N_18076,N_18690);
nor U19720 (N_19720,N_18357,N_18660);
nand U19721 (N_19721,N_18148,N_18442);
nand U19722 (N_19722,N_18788,N_18844);
nor U19723 (N_19723,N_18788,N_18143);
xnor U19724 (N_19724,N_18990,N_18638);
nand U19725 (N_19725,N_18640,N_18912);
or U19726 (N_19726,N_18006,N_18100);
xnor U19727 (N_19727,N_18495,N_18243);
or U19728 (N_19728,N_18899,N_18488);
and U19729 (N_19729,N_18818,N_18594);
and U19730 (N_19730,N_18597,N_18133);
nor U19731 (N_19731,N_18383,N_18780);
nand U19732 (N_19732,N_18768,N_18461);
and U19733 (N_19733,N_18063,N_18754);
xor U19734 (N_19734,N_18925,N_18630);
or U19735 (N_19735,N_18392,N_18640);
xor U19736 (N_19736,N_18985,N_18566);
or U19737 (N_19737,N_18512,N_18280);
xnor U19738 (N_19738,N_18271,N_18871);
nand U19739 (N_19739,N_18293,N_18662);
nand U19740 (N_19740,N_18308,N_18878);
xor U19741 (N_19741,N_18239,N_18287);
nor U19742 (N_19742,N_18142,N_18654);
and U19743 (N_19743,N_18563,N_18419);
nand U19744 (N_19744,N_18438,N_18632);
nand U19745 (N_19745,N_18139,N_18298);
xnor U19746 (N_19746,N_18361,N_18801);
or U19747 (N_19747,N_18558,N_18310);
and U19748 (N_19748,N_18657,N_18206);
and U19749 (N_19749,N_18652,N_18452);
xnor U19750 (N_19750,N_18383,N_18454);
nand U19751 (N_19751,N_18818,N_18131);
nor U19752 (N_19752,N_18855,N_18299);
xnor U19753 (N_19753,N_18291,N_18020);
nand U19754 (N_19754,N_18953,N_18663);
and U19755 (N_19755,N_18203,N_18851);
or U19756 (N_19756,N_18667,N_18209);
xor U19757 (N_19757,N_18460,N_18699);
nand U19758 (N_19758,N_18003,N_18732);
and U19759 (N_19759,N_18951,N_18552);
nand U19760 (N_19760,N_18235,N_18336);
nand U19761 (N_19761,N_18577,N_18420);
nor U19762 (N_19762,N_18804,N_18633);
and U19763 (N_19763,N_18686,N_18349);
nor U19764 (N_19764,N_18003,N_18422);
nor U19765 (N_19765,N_18245,N_18222);
or U19766 (N_19766,N_18129,N_18727);
xnor U19767 (N_19767,N_18618,N_18286);
or U19768 (N_19768,N_18203,N_18811);
xnor U19769 (N_19769,N_18763,N_18729);
xor U19770 (N_19770,N_18797,N_18088);
and U19771 (N_19771,N_18625,N_18401);
xnor U19772 (N_19772,N_18799,N_18053);
nand U19773 (N_19773,N_18667,N_18436);
and U19774 (N_19774,N_18707,N_18838);
nor U19775 (N_19775,N_18412,N_18460);
and U19776 (N_19776,N_18584,N_18122);
and U19777 (N_19777,N_18651,N_18353);
or U19778 (N_19778,N_18021,N_18371);
and U19779 (N_19779,N_18469,N_18728);
nand U19780 (N_19780,N_18896,N_18773);
and U19781 (N_19781,N_18417,N_18034);
nor U19782 (N_19782,N_18861,N_18389);
or U19783 (N_19783,N_18247,N_18787);
nor U19784 (N_19784,N_18979,N_18782);
nand U19785 (N_19785,N_18129,N_18540);
nor U19786 (N_19786,N_18865,N_18050);
or U19787 (N_19787,N_18805,N_18011);
and U19788 (N_19788,N_18211,N_18970);
nor U19789 (N_19789,N_18594,N_18352);
nor U19790 (N_19790,N_18073,N_18420);
nor U19791 (N_19791,N_18927,N_18898);
nand U19792 (N_19792,N_18509,N_18167);
or U19793 (N_19793,N_18171,N_18855);
xnor U19794 (N_19794,N_18717,N_18964);
and U19795 (N_19795,N_18472,N_18009);
or U19796 (N_19796,N_18641,N_18228);
xor U19797 (N_19797,N_18562,N_18446);
and U19798 (N_19798,N_18598,N_18381);
nor U19799 (N_19799,N_18715,N_18071);
and U19800 (N_19800,N_18440,N_18237);
xor U19801 (N_19801,N_18026,N_18431);
nand U19802 (N_19802,N_18637,N_18237);
nor U19803 (N_19803,N_18422,N_18508);
nor U19804 (N_19804,N_18318,N_18775);
or U19805 (N_19805,N_18766,N_18001);
and U19806 (N_19806,N_18506,N_18162);
nor U19807 (N_19807,N_18672,N_18763);
nand U19808 (N_19808,N_18583,N_18316);
and U19809 (N_19809,N_18935,N_18597);
nand U19810 (N_19810,N_18370,N_18053);
and U19811 (N_19811,N_18263,N_18591);
or U19812 (N_19812,N_18640,N_18636);
xnor U19813 (N_19813,N_18145,N_18019);
nand U19814 (N_19814,N_18455,N_18634);
or U19815 (N_19815,N_18097,N_18738);
nor U19816 (N_19816,N_18154,N_18443);
xnor U19817 (N_19817,N_18446,N_18182);
or U19818 (N_19818,N_18529,N_18884);
or U19819 (N_19819,N_18998,N_18845);
nor U19820 (N_19820,N_18840,N_18183);
nor U19821 (N_19821,N_18500,N_18167);
xor U19822 (N_19822,N_18142,N_18959);
or U19823 (N_19823,N_18856,N_18314);
xnor U19824 (N_19824,N_18290,N_18195);
xor U19825 (N_19825,N_18110,N_18494);
or U19826 (N_19826,N_18883,N_18079);
nand U19827 (N_19827,N_18866,N_18491);
and U19828 (N_19828,N_18104,N_18921);
nor U19829 (N_19829,N_18127,N_18194);
nor U19830 (N_19830,N_18164,N_18432);
xnor U19831 (N_19831,N_18179,N_18240);
xnor U19832 (N_19832,N_18732,N_18276);
or U19833 (N_19833,N_18408,N_18916);
nor U19834 (N_19834,N_18479,N_18395);
or U19835 (N_19835,N_18217,N_18133);
and U19836 (N_19836,N_18554,N_18751);
or U19837 (N_19837,N_18981,N_18914);
and U19838 (N_19838,N_18537,N_18100);
nor U19839 (N_19839,N_18040,N_18085);
xnor U19840 (N_19840,N_18000,N_18431);
or U19841 (N_19841,N_18386,N_18400);
nor U19842 (N_19842,N_18984,N_18442);
or U19843 (N_19843,N_18202,N_18664);
and U19844 (N_19844,N_18470,N_18341);
and U19845 (N_19845,N_18008,N_18713);
and U19846 (N_19846,N_18197,N_18650);
xnor U19847 (N_19847,N_18067,N_18240);
xnor U19848 (N_19848,N_18249,N_18341);
xnor U19849 (N_19849,N_18789,N_18209);
nand U19850 (N_19850,N_18034,N_18442);
and U19851 (N_19851,N_18051,N_18745);
nor U19852 (N_19852,N_18869,N_18253);
and U19853 (N_19853,N_18559,N_18517);
xnor U19854 (N_19854,N_18479,N_18527);
nor U19855 (N_19855,N_18204,N_18843);
nor U19856 (N_19856,N_18297,N_18300);
nand U19857 (N_19857,N_18251,N_18450);
nand U19858 (N_19858,N_18271,N_18431);
nor U19859 (N_19859,N_18081,N_18162);
or U19860 (N_19860,N_18488,N_18267);
nand U19861 (N_19861,N_18711,N_18262);
nand U19862 (N_19862,N_18115,N_18879);
nand U19863 (N_19863,N_18772,N_18559);
and U19864 (N_19864,N_18225,N_18283);
nand U19865 (N_19865,N_18098,N_18419);
xor U19866 (N_19866,N_18205,N_18554);
or U19867 (N_19867,N_18777,N_18717);
xnor U19868 (N_19868,N_18935,N_18823);
or U19869 (N_19869,N_18278,N_18252);
or U19870 (N_19870,N_18712,N_18205);
nor U19871 (N_19871,N_18464,N_18940);
or U19872 (N_19872,N_18051,N_18502);
nor U19873 (N_19873,N_18128,N_18033);
and U19874 (N_19874,N_18505,N_18199);
and U19875 (N_19875,N_18101,N_18365);
xor U19876 (N_19876,N_18726,N_18688);
nand U19877 (N_19877,N_18013,N_18320);
nand U19878 (N_19878,N_18895,N_18914);
nor U19879 (N_19879,N_18701,N_18382);
and U19880 (N_19880,N_18158,N_18648);
nor U19881 (N_19881,N_18690,N_18839);
and U19882 (N_19882,N_18467,N_18336);
xor U19883 (N_19883,N_18671,N_18347);
nand U19884 (N_19884,N_18434,N_18259);
and U19885 (N_19885,N_18974,N_18696);
nand U19886 (N_19886,N_18920,N_18141);
and U19887 (N_19887,N_18304,N_18522);
or U19888 (N_19888,N_18726,N_18111);
nor U19889 (N_19889,N_18912,N_18900);
and U19890 (N_19890,N_18925,N_18068);
and U19891 (N_19891,N_18388,N_18053);
nor U19892 (N_19892,N_18992,N_18340);
or U19893 (N_19893,N_18462,N_18627);
nor U19894 (N_19894,N_18760,N_18360);
nand U19895 (N_19895,N_18397,N_18253);
and U19896 (N_19896,N_18138,N_18631);
nand U19897 (N_19897,N_18061,N_18340);
nand U19898 (N_19898,N_18066,N_18787);
nand U19899 (N_19899,N_18317,N_18893);
or U19900 (N_19900,N_18761,N_18922);
xor U19901 (N_19901,N_18806,N_18157);
or U19902 (N_19902,N_18027,N_18616);
or U19903 (N_19903,N_18406,N_18050);
nand U19904 (N_19904,N_18317,N_18819);
and U19905 (N_19905,N_18685,N_18462);
and U19906 (N_19906,N_18804,N_18784);
and U19907 (N_19907,N_18270,N_18605);
xor U19908 (N_19908,N_18346,N_18233);
nand U19909 (N_19909,N_18979,N_18018);
nor U19910 (N_19910,N_18242,N_18716);
nand U19911 (N_19911,N_18485,N_18738);
xnor U19912 (N_19912,N_18559,N_18892);
or U19913 (N_19913,N_18532,N_18777);
and U19914 (N_19914,N_18244,N_18051);
xor U19915 (N_19915,N_18990,N_18689);
and U19916 (N_19916,N_18494,N_18384);
and U19917 (N_19917,N_18996,N_18022);
nand U19918 (N_19918,N_18045,N_18513);
nand U19919 (N_19919,N_18667,N_18293);
nor U19920 (N_19920,N_18846,N_18159);
nor U19921 (N_19921,N_18605,N_18161);
nor U19922 (N_19922,N_18931,N_18520);
nor U19923 (N_19923,N_18836,N_18631);
nor U19924 (N_19924,N_18118,N_18318);
nor U19925 (N_19925,N_18103,N_18593);
xnor U19926 (N_19926,N_18137,N_18743);
nor U19927 (N_19927,N_18618,N_18925);
nand U19928 (N_19928,N_18955,N_18202);
nand U19929 (N_19929,N_18684,N_18043);
nor U19930 (N_19930,N_18704,N_18435);
nor U19931 (N_19931,N_18570,N_18852);
xor U19932 (N_19932,N_18779,N_18174);
or U19933 (N_19933,N_18388,N_18973);
xnor U19934 (N_19934,N_18448,N_18607);
nand U19935 (N_19935,N_18981,N_18118);
or U19936 (N_19936,N_18131,N_18365);
nor U19937 (N_19937,N_18482,N_18140);
nand U19938 (N_19938,N_18225,N_18114);
nand U19939 (N_19939,N_18670,N_18352);
nor U19940 (N_19940,N_18740,N_18814);
and U19941 (N_19941,N_18581,N_18686);
xnor U19942 (N_19942,N_18731,N_18459);
nand U19943 (N_19943,N_18520,N_18947);
xnor U19944 (N_19944,N_18048,N_18816);
nor U19945 (N_19945,N_18956,N_18327);
or U19946 (N_19946,N_18091,N_18563);
or U19947 (N_19947,N_18738,N_18079);
nor U19948 (N_19948,N_18714,N_18610);
and U19949 (N_19949,N_18901,N_18812);
nand U19950 (N_19950,N_18418,N_18686);
nor U19951 (N_19951,N_18262,N_18273);
and U19952 (N_19952,N_18493,N_18339);
or U19953 (N_19953,N_18244,N_18451);
nand U19954 (N_19954,N_18790,N_18611);
nand U19955 (N_19955,N_18681,N_18121);
and U19956 (N_19956,N_18692,N_18195);
nor U19957 (N_19957,N_18616,N_18973);
or U19958 (N_19958,N_18504,N_18238);
and U19959 (N_19959,N_18456,N_18164);
and U19960 (N_19960,N_18965,N_18529);
xnor U19961 (N_19961,N_18785,N_18052);
and U19962 (N_19962,N_18289,N_18972);
nor U19963 (N_19963,N_18740,N_18146);
nor U19964 (N_19964,N_18669,N_18406);
nand U19965 (N_19965,N_18388,N_18461);
nor U19966 (N_19966,N_18465,N_18384);
nand U19967 (N_19967,N_18787,N_18460);
xnor U19968 (N_19968,N_18951,N_18396);
nand U19969 (N_19969,N_18333,N_18652);
and U19970 (N_19970,N_18738,N_18053);
xor U19971 (N_19971,N_18135,N_18812);
nand U19972 (N_19972,N_18096,N_18371);
and U19973 (N_19973,N_18618,N_18490);
and U19974 (N_19974,N_18573,N_18521);
xor U19975 (N_19975,N_18658,N_18561);
xor U19976 (N_19976,N_18230,N_18000);
nand U19977 (N_19977,N_18833,N_18682);
and U19978 (N_19978,N_18667,N_18484);
nand U19979 (N_19979,N_18559,N_18023);
xnor U19980 (N_19980,N_18916,N_18457);
nand U19981 (N_19981,N_18089,N_18854);
nand U19982 (N_19982,N_18041,N_18538);
xnor U19983 (N_19983,N_18221,N_18280);
xor U19984 (N_19984,N_18419,N_18166);
or U19985 (N_19985,N_18225,N_18152);
nand U19986 (N_19986,N_18030,N_18775);
nor U19987 (N_19987,N_18249,N_18903);
or U19988 (N_19988,N_18927,N_18299);
nand U19989 (N_19989,N_18713,N_18894);
xnor U19990 (N_19990,N_18457,N_18482);
nor U19991 (N_19991,N_18639,N_18219);
nor U19992 (N_19992,N_18771,N_18479);
nand U19993 (N_19993,N_18502,N_18215);
xnor U19994 (N_19994,N_18496,N_18743);
xor U19995 (N_19995,N_18629,N_18389);
nor U19996 (N_19996,N_18613,N_18338);
nor U19997 (N_19997,N_18237,N_18066);
nand U19998 (N_19998,N_18277,N_18897);
xor U19999 (N_19999,N_18749,N_18841);
nand U20000 (N_20000,N_19471,N_19949);
or U20001 (N_20001,N_19518,N_19812);
nor U20002 (N_20002,N_19808,N_19843);
xnor U20003 (N_20003,N_19546,N_19063);
nand U20004 (N_20004,N_19517,N_19172);
or U20005 (N_20005,N_19775,N_19888);
and U20006 (N_20006,N_19248,N_19711);
xor U20007 (N_20007,N_19942,N_19866);
nand U20008 (N_20008,N_19487,N_19432);
nor U20009 (N_20009,N_19145,N_19270);
nand U20010 (N_20010,N_19175,N_19663);
and U20011 (N_20011,N_19390,N_19814);
xor U20012 (N_20012,N_19097,N_19996);
nand U20013 (N_20013,N_19096,N_19633);
xor U20014 (N_20014,N_19393,N_19596);
xnor U20015 (N_20015,N_19299,N_19014);
or U20016 (N_20016,N_19321,N_19740);
xor U20017 (N_20017,N_19274,N_19642);
and U20018 (N_20018,N_19442,N_19056);
nor U20019 (N_20019,N_19715,N_19406);
and U20020 (N_20020,N_19222,N_19915);
nand U20021 (N_20021,N_19832,N_19520);
xnor U20022 (N_20022,N_19875,N_19162);
nor U20023 (N_20023,N_19948,N_19408);
and U20024 (N_20024,N_19758,N_19603);
nand U20025 (N_20025,N_19804,N_19824);
and U20026 (N_20026,N_19239,N_19127);
nor U20027 (N_20027,N_19241,N_19320);
nand U20028 (N_20028,N_19375,N_19292);
nand U20029 (N_20029,N_19753,N_19280);
nor U20030 (N_20030,N_19577,N_19848);
nor U20031 (N_20031,N_19584,N_19331);
nand U20032 (N_20032,N_19865,N_19288);
and U20033 (N_20033,N_19041,N_19620);
nor U20034 (N_20034,N_19233,N_19240);
nand U20035 (N_20035,N_19896,N_19493);
and U20036 (N_20036,N_19975,N_19434);
nand U20037 (N_20037,N_19864,N_19606);
nand U20038 (N_20038,N_19821,N_19287);
nand U20039 (N_20039,N_19460,N_19857);
nand U20040 (N_20040,N_19858,N_19874);
and U20041 (N_20041,N_19319,N_19081);
nand U20042 (N_20042,N_19484,N_19072);
and U20043 (N_20043,N_19835,N_19541);
and U20044 (N_20044,N_19163,N_19730);
or U20045 (N_20045,N_19710,N_19469);
xor U20046 (N_20046,N_19568,N_19905);
nor U20047 (N_20047,N_19437,N_19306);
xor U20048 (N_20048,N_19261,N_19472);
and U20049 (N_20049,N_19787,N_19997);
nand U20050 (N_20050,N_19531,N_19677);
nand U20051 (N_20051,N_19533,N_19912);
or U20052 (N_20052,N_19330,N_19614);
nand U20053 (N_20053,N_19456,N_19553);
nand U20054 (N_20054,N_19149,N_19561);
nor U20055 (N_20055,N_19882,N_19772);
xor U20056 (N_20056,N_19994,N_19571);
or U20057 (N_20057,N_19588,N_19855);
or U20058 (N_20058,N_19295,N_19404);
xor U20059 (N_20059,N_19635,N_19687);
xor U20060 (N_20060,N_19226,N_19315);
nand U20061 (N_20061,N_19585,N_19567);
and U20062 (N_20062,N_19216,N_19581);
or U20063 (N_20063,N_19766,N_19329);
nor U20064 (N_20064,N_19387,N_19514);
xor U20065 (N_20065,N_19652,N_19177);
and U20066 (N_20066,N_19807,N_19282);
nand U20067 (N_20067,N_19968,N_19269);
and U20068 (N_20068,N_19289,N_19001);
xor U20069 (N_20069,N_19719,N_19862);
nor U20070 (N_20070,N_19675,N_19830);
nor U20071 (N_20071,N_19351,N_19921);
nand U20072 (N_20072,N_19077,N_19383);
and U20073 (N_20073,N_19872,N_19178);
nand U20074 (N_20074,N_19294,N_19300);
and U20075 (N_20075,N_19420,N_19703);
and U20076 (N_20076,N_19395,N_19630);
nor U20077 (N_20077,N_19119,N_19904);
and U20078 (N_20078,N_19970,N_19651);
nor U20079 (N_20079,N_19958,N_19445);
nand U20080 (N_20080,N_19556,N_19697);
xor U20081 (N_20081,N_19142,N_19025);
xor U20082 (N_20082,N_19680,N_19343);
and U20083 (N_20083,N_19078,N_19124);
or U20084 (N_20084,N_19622,N_19938);
nand U20085 (N_20085,N_19252,N_19380);
or U20086 (N_20086,N_19350,N_19899);
nor U20087 (N_20087,N_19168,N_19479);
nand U20088 (N_20088,N_19809,N_19369);
or U20089 (N_20089,N_19601,N_19881);
xnor U20090 (N_20090,N_19598,N_19190);
nor U20091 (N_20091,N_19424,N_19000);
xnor U20092 (N_20092,N_19061,N_19509);
nor U20093 (N_20093,N_19993,N_19324);
xnor U20094 (N_20094,N_19505,N_19754);
and U20095 (N_20095,N_19203,N_19842);
nand U20096 (N_20096,N_19731,N_19264);
or U20097 (N_20097,N_19782,N_19522);
nand U20098 (N_20098,N_19473,N_19370);
nand U20099 (N_20099,N_19026,N_19152);
or U20100 (N_20100,N_19836,N_19566);
nand U20101 (N_20101,N_19851,N_19759);
nand U20102 (N_20102,N_19853,N_19671);
nand U20103 (N_20103,N_19798,N_19047);
or U20104 (N_20104,N_19192,N_19694);
or U20105 (N_20105,N_19748,N_19786);
nor U20106 (N_20106,N_19037,N_19825);
and U20107 (N_20107,N_19764,N_19594);
nand U20108 (N_20108,N_19373,N_19173);
nand U20109 (N_20109,N_19455,N_19273);
nand U20110 (N_20110,N_19377,N_19805);
xor U20111 (N_20111,N_19305,N_19854);
nor U20112 (N_20112,N_19962,N_19547);
or U20113 (N_20113,N_19794,N_19504);
nand U20114 (N_20114,N_19323,N_19550);
xnor U20115 (N_20115,N_19636,N_19345);
and U20116 (N_20116,N_19342,N_19044);
or U20117 (N_20117,N_19511,N_19003);
and U20118 (N_20118,N_19111,N_19744);
and U20119 (N_20119,N_19153,N_19735);
nor U20120 (N_20120,N_19184,N_19777);
nand U20121 (N_20121,N_19684,N_19910);
xor U20122 (N_20122,N_19201,N_19086);
xor U20123 (N_20123,N_19823,N_19954);
and U20124 (N_20124,N_19562,N_19655);
or U20125 (N_20125,N_19117,N_19937);
or U20126 (N_20126,N_19451,N_19477);
xor U20127 (N_20127,N_19403,N_19946);
nor U20128 (N_20128,N_19412,N_19510);
or U20129 (N_20129,N_19422,N_19974);
and U20130 (N_20130,N_19980,N_19795);
nand U20131 (N_20131,N_19180,N_19413);
or U20132 (N_20132,N_19668,N_19291);
nand U20133 (N_20133,N_19641,N_19174);
and U20134 (N_20134,N_19712,N_19544);
xor U20135 (N_20135,N_19244,N_19618);
nand U20136 (N_20136,N_19771,N_19947);
and U20137 (N_20137,N_19347,N_19829);
and U20138 (N_20138,N_19046,N_19101);
xnor U20139 (N_20139,N_19931,N_19441);
nand U20140 (N_20140,N_19691,N_19893);
and U20141 (N_20141,N_19746,N_19155);
or U20142 (N_20142,N_19778,N_19672);
or U20143 (N_20143,N_19245,N_19191);
or U20144 (N_20144,N_19138,N_19376);
and U20145 (N_20145,N_19870,N_19978);
nor U20146 (N_20146,N_19845,N_19890);
and U20147 (N_20147,N_19067,N_19987);
nor U20148 (N_20148,N_19033,N_19426);
nor U20149 (N_20149,N_19924,N_19538);
and U20150 (N_20150,N_19116,N_19246);
nor U20151 (N_20151,N_19483,N_19353);
or U20152 (N_20152,N_19907,N_19869);
and U20153 (N_20153,N_19389,N_19834);
nor U20154 (N_20154,N_19335,N_19010);
nand U20155 (N_20155,N_19950,N_19963);
nor U20156 (N_20156,N_19030,N_19647);
nand U20157 (N_20157,N_19685,N_19151);
nand U20158 (N_20158,N_19590,N_19500);
nand U20159 (N_20159,N_19283,N_19150);
nor U20160 (N_20160,N_19727,N_19064);
and U20161 (N_20161,N_19070,N_19029);
and U20162 (N_20162,N_19849,N_19820);
or U20163 (N_20163,N_19513,N_19301);
nor U20164 (N_20164,N_19346,N_19976);
and U20165 (N_20165,N_19995,N_19999);
nand U20166 (N_20166,N_19444,N_19705);
or U20167 (N_20167,N_19654,N_19235);
and U20168 (N_20168,N_19723,N_19747);
and U20169 (N_20169,N_19068,N_19250);
or U20170 (N_20170,N_19113,N_19889);
nand U20171 (N_20171,N_19313,N_19088);
and U20172 (N_20172,N_19597,N_19815);
and U20173 (N_20173,N_19920,N_19625);
and U20174 (N_20174,N_19751,N_19491);
xnor U20175 (N_20175,N_19157,N_19349);
and U20176 (N_20176,N_19692,N_19414);
xnor U20177 (N_20177,N_19755,N_19580);
or U20178 (N_20178,N_19650,N_19645);
or U20179 (N_20179,N_19637,N_19411);
xor U20180 (N_20180,N_19489,N_19717);
or U20181 (N_20181,N_19956,N_19789);
xor U20182 (N_20182,N_19297,N_19200);
xnor U20183 (N_20183,N_19521,N_19091);
xor U20184 (N_20184,N_19108,N_19257);
or U20185 (N_20185,N_19498,N_19388);
or U20186 (N_20186,N_19016,N_19847);
xnor U20187 (N_20187,N_19761,N_19900);
and U20188 (N_20188,N_19262,N_19933);
nand U20189 (N_20189,N_19336,N_19219);
xnor U20190 (N_20190,N_19918,N_19932);
and U20191 (N_20191,N_19986,N_19617);
nand U20192 (N_20192,N_19176,N_19923);
and U20193 (N_20193,N_19573,N_19371);
or U20194 (N_20194,N_19217,N_19058);
and U20195 (N_20195,N_19673,N_19326);
and U20196 (N_20196,N_19199,N_19800);
and U20197 (N_20197,N_19419,N_19496);
xnor U20198 (N_20198,N_19548,N_19495);
nor U20199 (N_20199,N_19440,N_19130);
nand U20200 (N_20200,N_19154,N_19228);
xor U20201 (N_20201,N_19443,N_19578);
and U20202 (N_20202,N_19549,N_19208);
nor U20203 (N_20203,N_19732,N_19132);
nand U20204 (N_20204,N_19565,N_19340);
and U20205 (N_20205,N_19234,N_19075);
and U20206 (N_20206,N_19325,N_19988);
xnor U20207 (N_20207,N_19507,N_19019);
xor U20208 (N_20208,N_19856,N_19143);
or U20209 (N_20209,N_19537,N_19284);
nand U20210 (N_20210,N_19634,N_19470);
nor U20211 (N_20211,N_19608,N_19868);
nor U20212 (N_20212,N_19425,N_19629);
nand U20213 (N_20213,N_19318,N_19415);
xnor U20214 (N_20214,N_19038,N_19939);
xnor U20215 (N_20215,N_19605,N_19359);
and U20216 (N_20216,N_19121,N_19039);
xnor U20217 (N_20217,N_19073,N_19783);
xor U20218 (N_20218,N_19107,N_19666);
xor U20219 (N_20219,N_19913,N_19205);
nand U20220 (N_20220,N_19012,N_19187);
and U20221 (N_20221,N_19600,N_19861);
or U20222 (N_20222,N_19551,N_19526);
nand U20223 (N_20223,N_19658,N_19693);
nand U20224 (N_20224,N_19611,N_19409);
nand U20225 (N_20225,N_19136,N_19040);
and U20226 (N_20226,N_19678,N_19202);
or U20227 (N_20227,N_19819,N_19468);
nor U20228 (N_20228,N_19797,N_19362);
xnor U20229 (N_20229,N_19099,N_19344);
or U20230 (N_20230,N_19524,N_19066);
or U20231 (N_20231,N_19396,N_19700);
or U20232 (N_20232,N_19941,N_19756);
nor U20233 (N_20233,N_19196,N_19887);
nand U20234 (N_20234,N_19166,N_19131);
and U20235 (N_20235,N_19661,N_19035);
and U20236 (N_20236,N_19981,N_19171);
nor U20237 (N_20237,N_19427,N_19144);
nor U20238 (N_20238,N_19052,N_19276);
xor U20239 (N_20239,N_19583,N_19838);
and U20240 (N_20240,N_19643,N_19218);
or U20241 (N_20241,N_19281,N_19502);
xor U20242 (N_20242,N_19686,N_19007);
or U20243 (N_20243,N_19539,N_19615);
nand U20244 (N_20244,N_19574,N_19768);
xor U20245 (N_20245,N_19271,N_19267);
and U20246 (N_20246,N_19213,N_19901);
nand U20247 (N_20247,N_19708,N_19013);
and U20248 (N_20248,N_19702,N_19322);
or U20249 (N_20249,N_19765,N_19465);
or U20250 (N_20250,N_19895,N_19640);
or U20251 (N_20251,N_19841,N_19015);
nand U20252 (N_20252,N_19298,N_19207);
or U20253 (N_20253,N_19115,N_19743);
nor U20254 (N_20254,N_19688,N_19646);
xnor U20255 (N_20255,N_19259,N_19979);
nand U20256 (N_20256,N_19475,N_19619);
xor U20257 (N_20257,N_19185,N_19485);
nor U20258 (N_20258,N_19095,N_19368);
xnor U20259 (N_20259,N_19238,N_19911);
nand U20260 (N_20260,N_19966,N_19990);
xor U20261 (N_20261,N_19059,N_19796);
and U20262 (N_20262,N_19227,N_19198);
or U20263 (N_20263,N_19243,N_19828);
xor U20264 (N_20264,N_19360,N_19916);
nor U20265 (N_20265,N_19194,N_19555);
and U20266 (N_20266,N_19290,N_19811);
xor U20267 (N_20267,N_19022,N_19447);
nor U20268 (N_20268,N_19718,N_19628);
or U20269 (N_20269,N_19286,N_19927);
and U20270 (N_20270,N_19589,N_19112);
and U20271 (N_20271,N_19381,N_19639);
nand U20272 (N_20272,N_19716,N_19055);
xnor U20273 (N_20273,N_19348,N_19846);
nand U20274 (N_20274,N_19147,N_19497);
nand U20275 (N_20275,N_19255,N_19232);
and U20276 (N_20276,N_19860,N_19867);
nor U20277 (N_20277,N_19940,N_19114);
and U20278 (N_20278,N_19602,N_19833);
nor U20279 (N_20279,N_19372,N_19781);
or U20280 (N_20280,N_19231,N_19785);
xnor U20281 (N_20281,N_19429,N_19453);
nor U20282 (N_20282,N_19229,N_19126);
xor U20283 (N_20283,N_19023,N_19333);
nand U20284 (N_20284,N_19515,N_19363);
nand U20285 (N_20285,N_19586,N_19309);
or U20286 (N_20286,N_19110,N_19935);
and U20287 (N_20287,N_19263,N_19159);
nand U20288 (N_20288,N_19951,N_19822);
and U20289 (N_20289,N_19220,N_19891);
or U20290 (N_20290,N_19017,N_19384);
xor U20291 (N_20291,N_19579,N_19354);
or U20292 (N_20292,N_19183,N_19894);
nor U20293 (N_20293,N_19128,N_19928);
xnor U20294 (N_20294,N_19206,N_19466);
or U20295 (N_20295,N_19186,N_19738);
and U20296 (N_20296,N_19944,N_19418);
nand U20297 (N_20297,N_19382,N_19914);
and U20298 (N_20298,N_19791,N_19906);
and U20299 (N_20299,N_19474,N_19133);
nand U20300 (N_20300,N_19713,N_19105);
nor U20301 (N_20301,N_19595,N_19750);
nor U20302 (N_20302,N_19665,N_19612);
and U20303 (N_20303,N_19268,N_19050);
nand U20304 (N_20304,N_19402,N_19525);
xnor U20305 (N_20305,N_19311,N_19985);
nor U20306 (N_20306,N_19123,N_19506);
or U20307 (N_20307,N_19417,N_19767);
nor U20308 (N_20308,N_19083,N_19569);
nand U20309 (N_20309,N_19886,N_19043);
nor U20310 (N_20310,N_19535,N_19763);
nor U20311 (N_20311,N_19774,N_19967);
nand U20312 (N_20312,N_19929,N_19065);
or U20313 (N_20313,N_19793,N_19316);
or U20314 (N_20314,N_19314,N_19249);
nor U20315 (N_20315,N_19729,N_19728);
nor U20316 (N_20316,N_19071,N_19436);
and U20317 (N_20317,N_19883,N_19054);
nand U20318 (N_20318,N_19366,N_19638);
nand U20319 (N_20319,N_19850,N_19394);
nand U20320 (N_20320,N_19446,N_19745);
nand U20321 (N_20321,N_19837,N_19021);
nand U20322 (N_20322,N_19048,N_19140);
or U20323 (N_20323,N_19790,N_19532);
nand U20324 (N_20324,N_19272,N_19458);
nor U20325 (N_20325,N_19624,N_19439);
and U20326 (N_20326,N_19564,N_19873);
nor U20327 (N_20327,N_19512,N_19648);
nand U20328 (N_20328,N_19880,N_19662);
nor U20329 (N_20329,N_19356,N_19258);
and U20330 (N_20330,N_19438,N_19435);
nand U20331 (N_20331,N_19161,N_19167);
and U20332 (N_20332,N_19839,N_19757);
nor U20333 (N_20333,N_19179,N_19984);
or U20334 (N_20334,N_19508,N_19779);
nand U20335 (N_20335,N_19736,N_19523);
nor U20336 (N_20336,N_19977,N_19339);
or U20337 (N_20337,N_19752,N_19478);
xnor U20338 (N_20338,N_19042,N_19352);
xnor U20339 (N_20339,N_19604,N_19725);
xnor U20340 (N_20340,N_19223,N_19667);
xor U20341 (N_20341,N_19784,N_19361);
nand U20342 (N_20342,N_19934,N_19169);
nand U20343 (N_20343,N_19557,N_19328);
nand U20344 (N_20344,N_19773,N_19587);
xor U20345 (N_20345,N_19109,N_19279);
or U20346 (N_20346,N_19516,N_19897);
and U20347 (N_20347,N_19433,N_19092);
and U20348 (N_20348,N_19386,N_19733);
nor U20349 (N_20349,N_19462,N_19158);
xor U20350 (N_20350,N_19256,N_19749);
or U20351 (N_20351,N_19254,N_19737);
and U20352 (N_20352,N_19945,N_19265);
nor U20353 (N_20353,N_19660,N_19724);
or U20354 (N_20354,N_19721,N_19135);
nor U20355 (N_20355,N_19100,N_19069);
nand U20356 (N_20356,N_19399,N_19871);
nor U20357 (N_20357,N_19327,N_19308);
or U20358 (N_20358,N_19008,N_19631);
xnor U20359 (N_20359,N_19720,N_19476);
xnor U20360 (N_20360,N_19103,N_19307);
and U20361 (N_20361,N_19215,N_19627);
nand U20362 (N_20362,N_19285,N_19664);
or U20363 (N_20363,N_19407,N_19051);
and U20364 (N_20364,N_19379,N_19826);
and U20365 (N_20365,N_19714,N_19741);
nand U20366 (N_20366,N_19405,N_19090);
or U20367 (N_20367,N_19576,N_19401);
nand U20368 (N_20368,N_19397,N_19098);
and U20369 (N_20369,N_19844,N_19607);
or U20370 (N_20370,N_19011,N_19903);
nand U20371 (N_20371,N_19020,N_19801);
or U20372 (N_20372,N_19428,N_19006);
nand U20373 (N_20373,N_19189,N_19304);
and U20374 (N_20374,N_19225,N_19251);
xor U20375 (N_20375,N_19224,N_19852);
or U20376 (N_20376,N_19093,N_19957);
or U20377 (N_20377,N_19649,N_19696);
nor U20378 (N_20378,N_19094,N_19769);
and U20379 (N_20379,N_19034,N_19799);
nand U20380 (N_20380,N_19045,N_19181);
xnor U20381 (N_20381,N_19554,N_19334);
nor U20382 (N_20382,N_19572,N_19275);
and U20383 (N_20383,N_19613,N_19398);
and U20384 (N_20384,N_19087,N_19490);
or U20385 (N_20385,N_19210,N_19338);
nand U20386 (N_20386,N_19357,N_19813);
nor U20387 (N_20387,N_19623,N_19591);
nor U20388 (N_20388,N_19722,N_19632);
and U20389 (N_20389,N_19884,N_19626);
nor U20390 (N_20390,N_19141,N_19392);
xnor U20391 (N_20391,N_19818,N_19018);
nor U20392 (N_20392,N_19503,N_19670);
or U20393 (N_20393,N_19552,N_19193);
nand U20394 (N_20394,N_19961,N_19616);
and U20395 (N_20395,N_19780,N_19024);
nand U20396 (N_20396,N_19247,N_19971);
nor U20397 (N_20397,N_19709,N_19452);
nor U20398 (N_20398,N_19076,N_19317);
and U20399 (N_20399,N_19391,N_19104);
or U20400 (N_20400,N_19528,N_19480);
xor U20401 (N_20401,N_19592,N_19302);
nor U20402 (N_20402,N_19542,N_19488);
and U20403 (N_20403,N_19165,N_19296);
xor U20404 (N_20404,N_19558,N_19082);
and U20405 (N_20405,N_19028,N_19863);
nor U20406 (N_20406,N_19467,N_19085);
or U20407 (N_20407,N_19278,N_19908);
nand U20408 (N_20408,N_19621,N_19062);
nor U20409 (N_20409,N_19536,N_19965);
nor U20410 (N_20410,N_19683,N_19449);
nor U20411 (N_20411,N_19742,N_19005);
xnor U20412 (N_20412,N_19416,N_19337);
and U20413 (N_20413,N_19122,N_19204);
nor U20414 (N_20414,N_19690,N_19214);
or U20415 (N_20415,N_19461,N_19644);
nor U20416 (N_20416,N_19501,N_19817);
xor U20417 (N_20417,N_19534,N_19563);
nor U20418 (N_20418,N_19840,N_19423);
and U20419 (N_20419,N_19236,N_19410);
and U20420 (N_20420,N_19892,N_19653);
nand U20421 (N_20421,N_19679,N_19657);
xnor U20422 (N_20422,N_19464,N_19450);
and U20423 (N_20423,N_19955,N_19118);
nor U20424 (N_20424,N_19463,N_19230);
xor U20425 (N_20425,N_19027,N_19878);
nor U20426 (N_20426,N_19310,N_19898);
and U20427 (N_20427,N_19266,N_19919);
nand U20428 (N_20428,N_19374,N_19312);
nand U20429 (N_20429,N_19365,N_19698);
nor U20430 (N_20430,N_19953,N_19482);
xor U20431 (N_20431,N_19293,N_19943);
xor U20432 (N_20432,N_19926,N_19527);
nand U20433 (N_20433,N_19827,N_19879);
nor U20434 (N_20434,N_19770,N_19049);
xor U20435 (N_20435,N_19610,N_19164);
or U20436 (N_20436,N_19936,N_19582);
and U20437 (N_20437,N_19593,N_19969);
and U20438 (N_20438,N_19792,N_19499);
or U20439 (N_20439,N_19925,N_19982);
nor U20440 (N_20440,N_19053,N_19146);
or U20441 (N_20441,N_19358,N_19831);
and U20442 (N_20442,N_19734,N_19530);
nand U20443 (N_20443,N_19519,N_19211);
and U20444 (N_20444,N_19195,N_19120);
xnor U20445 (N_20445,N_19364,N_19002);
nand U20446 (N_20446,N_19960,N_19922);
and U20447 (N_20447,N_19991,N_19609);
nand U20448 (N_20448,N_19084,N_19959);
and U20449 (N_20449,N_19902,N_19156);
and U20450 (N_20450,N_19992,N_19776);
xor U20451 (N_20451,N_19909,N_19459);
xnor U20452 (N_20452,N_19102,N_19876);
nand U20453 (N_20453,N_19448,N_19430);
or U20454 (N_20454,N_19089,N_19964);
xor U20455 (N_20455,N_19400,N_19139);
xor U20456 (N_20456,N_19125,N_19332);
nand U20457 (N_20457,N_19930,N_19806);
and U20458 (N_20458,N_19560,N_19385);
nand U20459 (N_20459,N_19188,N_19803);
or U20460 (N_20460,N_19378,N_19137);
nor U20461 (N_20461,N_19303,N_19129);
nor U20462 (N_20462,N_19681,N_19057);
and U20463 (N_20463,N_19492,N_19656);
and U20464 (N_20464,N_19431,N_19704);
and U20465 (N_20465,N_19543,N_19036);
or U20466 (N_20466,N_19341,N_19009);
or U20467 (N_20467,N_19481,N_19080);
xor U20468 (N_20468,N_19454,N_19998);
xor U20469 (N_20469,N_19277,N_19032);
and U20470 (N_20470,N_19148,N_19659);
nor U20471 (N_20471,N_19726,N_19421);
nor U20472 (N_20472,N_19952,N_19197);
and U20473 (N_20473,N_19212,N_19060);
and U20474 (N_20474,N_19599,N_19816);
xnor U20475 (N_20475,N_19917,N_19367);
or U20476 (N_20476,N_19486,N_19209);
nand U20477 (N_20477,N_19182,N_19106);
or U20478 (N_20478,N_19253,N_19689);
and U20479 (N_20479,N_19699,N_19575);
or U20480 (N_20480,N_19529,N_19160);
xnor U20481 (N_20481,N_19031,N_19570);
xor U20482 (N_20482,N_19762,N_19242);
and U20483 (N_20483,N_19983,N_19669);
and U20484 (N_20484,N_19706,N_19674);
nand U20485 (N_20485,N_19760,N_19260);
nand U20486 (N_20486,N_19676,N_19810);
nor U20487 (N_20487,N_19802,N_19494);
nand U20488 (N_20488,N_19682,N_19707);
and U20489 (N_20489,N_19989,N_19559);
nand U20490 (N_20490,N_19170,N_19545);
xor U20491 (N_20491,N_19877,N_19972);
xnor U20492 (N_20492,N_19695,N_19355);
or U20493 (N_20493,N_19859,N_19739);
or U20494 (N_20494,N_19701,N_19788);
nand U20495 (N_20495,N_19237,N_19457);
nor U20496 (N_20496,N_19074,N_19004);
or U20497 (N_20497,N_19540,N_19973);
nor U20498 (N_20498,N_19221,N_19134);
xor U20499 (N_20499,N_19885,N_19079);
and U20500 (N_20500,N_19796,N_19056);
xnor U20501 (N_20501,N_19410,N_19164);
or U20502 (N_20502,N_19281,N_19617);
or U20503 (N_20503,N_19100,N_19356);
nor U20504 (N_20504,N_19937,N_19295);
or U20505 (N_20505,N_19844,N_19532);
nor U20506 (N_20506,N_19006,N_19424);
nand U20507 (N_20507,N_19752,N_19196);
xnor U20508 (N_20508,N_19738,N_19021);
xnor U20509 (N_20509,N_19364,N_19457);
xnor U20510 (N_20510,N_19560,N_19947);
or U20511 (N_20511,N_19842,N_19688);
nor U20512 (N_20512,N_19119,N_19219);
nor U20513 (N_20513,N_19188,N_19561);
or U20514 (N_20514,N_19445,N_19474);
nand U20515 (N_20515,N_19663,N_19731);
nor U20516 (N_20516,N_19091,N_19939);
or U20517 (N_20517,N_19652,N_19754);
or U20518 (N_20518,N_19088,N_19161);
nor U20519 (N_20519,N_19056,N_19435);
and U20520 (N_20520,N_19666,N_19185);
xnor U20521 (N_20521,N_19363,N_19693);
xnor U20522 (N_20522,N_19233,N_19294);
nor U20523 (N_20523,N_19857,N_19560);
nor U20524 (N_20524,N_19646,N_19954);
or U20525 (N_20525,N_19386,N_19384);
xor U20526 (N_20526,N_19944,N_19804);
nor U20527 (N_20527,N_19442,N_19438);
or U20528 (N_20528,N_19691,N_19661);
or U20529 (N_20529,N_19895,N_19564);
or U20530 (N_20530,N_19368,N_19342);
xor U20531 (N_20531,N_19433,N_19494);
or U20532 (N_20532,N_19420,N_19972);
nor U20533 (N_20533,N_19718,N_19769);
nand U20534 (N_20534,N_19035,N_19233);
xor U20535 (N_20535,N_19371,N_19404);
and U20536 (N_20536,N_19895,N_19507);
nand U20537 (N_20537,N_19695,N_19460);
and U20538 (N_20538,N_19908,N_19270);
and U20539 (N_20539,N_19613,N_19408);
or U20540 (N_20540,N_19031,N_19799);
xnor U20541 (N_20541,N_19158,N_19645);
or U20542 (N_20542,N_19658,N_19758);
or U20543 (N_20543,N_19218,N_19116);
nor U20544 (N_20544,N_19936,N_19678);
xor U20545 (N_20545,N_19401,N_19772);
and U20546 (N_20546,N_19989,N_19975);
or U20547 (N_20547,N_19890,N_19480);
nor U20548 (N_20548,N_19727,N_19032);
nor U20549 (N_20549,N_19164,N_19300);
nand U20550 (N_20550,N_19714,N_19043);
xnor U20551 (N_20551,N_19906,N_19249);
nor U20552 (N_20552,N_19750,N_19052);
nor U20553 (N_20553,N_19991,N_19426);
and U20554 (N_20554,N_19336,N_19817);
xnor U20555 (N_20555,N_19285,N_19882);
nand U20556 (N_20556,N_19534,N_19381);
and U20557 (N_20557,N_19601,N_19994);
nor U20558 (N_20558,N_19991,N_19904);
xor U20559 (N_20559,N_19612,N_19607);
nor U20560 (N_20560,N_19818,N_19747);
nor U20561 (N_20561,N_19583,N_19321);
and U20562 (N_20562,N_19384,N_19286);
nor U20563 (N_20563,N_19226,N_19875);
nor U20564 (N_20564,N_19504,N_19777);
and U20565 (N_20565,N_19459,N_19428);
xor U20566 (N_20566,N_19082,N_19993);
xor U20567 (N_20567,N_19754,N_19976);
or U20568 (N_20568,N_19120,N_19653);
nor U20569 (N_20569,N_19776,N_19672);
and U20570 (N_20570,N_19991,N_19400);
xor U20571 (N_20571,N_19483,N_19032);
or U20572 (N_20572,N_19647,N_19373);
or U20573 (N_20573,N_19676,N_19165);
and U20574 (N_20574,N_19698,N_19511);
nand U20575 (N_20575,N_19376,N_19212);
xor U20576 (N_20576,N_19776,N_19526);
or U20577 (N_20577,N_19228,N_19754);
xor U20578 (N_20578,N_19211,N_19122);
nor U20579 (N_20579,N_19067,N_19836);
nand U20580 (N_20580,N_19095,N_19395);
and U20581 (N_20581,N_19706,N_19550);
or U20582 (N_20582,N_19596,N_19285);
nand U20583 (N_20583,N_19501,N_19276);
xor U20584 (N_20584,N_19400,N_19600);
xnor U20585 (N_20585,N_19568,N_19129);
or U20586 (N_20586,N_19759,N_19983);
nand U20587 (N_20587,N_19061,N_19353);
nand U20588 (N_20588,N_19051,N_19532);
xnor U20589 (N_20589,N_19227,N_19041);
nand U20590 (N_20590,N_19873,N_19250);
xor U20591 (N_20591,N_19146,N_19745);
and U20592 (N_20592,N_19891,N_19480);
nor U20593 (N_20593,N_19318,N_19613);
xnor U20594 (N_20594,N_19090,N_19012);
xor U20595 (N_20595,N_19375,N_19883);
and U20596 (N_20596,N_19966,N_19938);
or U20597 (N_20597,N_19303,N_19740);
xor U20598 (N_20598,N_19572,N_19059);
nand U20599 (N_20599,N_19565,N_19346);
nor U20600 (N_20600,N_19888,N_19285);
and U20601 (N_20601,N_19834,N_19678);
xor U20602 (N_20602,N_19500,N_19878);
and U20603 (N_20603,N_19331,N_19850);
and U20604 (N_20604,N_19116,N_19147);
and U20605 (N_20605,N_19249,N_19156);
and U20606 (N_20606,N_19719,N_19747);
or U20607 (N_20607,N_19500,N_19561);
nor U20608 (N_20608,N_19553,N_19848);
and U20609 (N_20609,N_19063,N_19418);
or U20610 (N_20610,N_19303,N_19324);
xor U20611 (N_20611,N_19271,N_19032);
nor U20612 (N_20612,N_19477,N_19572);
nand U20613 (N_20613,N_19999,N_19298);
and U20614 (N_20614,N_19835,N_19596);
nand U20615 (N_20615,N_19282,N_19043);
nor U20616 (N_20616,N_19940,N_19167);
and U20617 (N_20617,N_19048,N_19035);
xnor U20618 (N_20618,N_19294,N_19766);
xor U20619 (N_20619,N_19986,N_19008);
and U20620 (N_20620,N_19935,N_19820);
and U20621 (N_20621,N_19660,N_19184);
nor U20622 (N_20622,N_19127,N_19524);
and U20623 (N_20623,N_19506,N_19646);
or U20624 (N_20624,N_19254,N_19752);
nand U20625 (N_20625,N_19217,N_19814);
and U20626 (N_20626,N_19683,N_19183);
xor U20627 (N_20627,N_19289,N_19784);
xnor U20628 (N_20628,N_19553,N_19291);
xnor U20629 (N_20629,N_19423,N_19024);
xnor U20630 (N_20630,N_19615,N_19747);
nor U20631 (N_20631,N_19786,N_19951);
nor U20632 (N_20632,N_19780,N_19546);
xor U20633 (N_20633,N_19533,N_19658);
nor U20634 (N_20634,N_19163,N_19166);
nor U20635 (N_20635,N_19814,N_19113);
nand U20636 (N_20636,N_19968,N_19020);
xor U20637 (N_20637,N_19783,N_19899);
nor U20638 (N_20638,N_19967,N_19093);
nand U20639 (N_20639,N_19624,N_19227);
xor U20640 (N_20640,N_19988,N_19306);
xor U20641 (N_20641,N_19857,N_19603);
or U20642 (N_20642,N_19569,N_19429);
and U20643 (N_20643,N_19339,N_19150);
or U20644 (N_20644,N_19214,N_19929);
nand U20645 (N_20645,N_19135,N_19762);
and U20646 (N_20646,N_19573,N_19498);
and U20647 (N_20647,N_19062,N_19382);
nor U20648 (N_20648,N_19379,N_19290);
and U20649 (N_20649,N_19359,N_19688);
nor U20650 (N_20650,N_19356,N_19593);
nand U20651 (N_20651,N_19757,N_19044);
and U20652 (N_20652,N_19144,N_19867);
and U20653 (N_20653,N_19035,N_19057);
nor U20654 (N_20654,N_19571,N_19619);
nor U20655 (N_20655,N_19349,N_19693);
nor U20656 (N_20656,N_19860,N_19394);
xnor U20657 (N_20657,N_19155,N_19542);
nand U20658 (N_20658,N_19753,N_19524);
nand U20659 (N_20659,N_19774,N_19542);
nor U20660 (N_20660,N_19837,N_19786);
nor U20661 (N_20661,N_19046,N_19606);
nor U20662 (N_20662,N_19006,N_19881);
nand U20663 (N_20663,N_19953,N_19866);
nor U20664 (N_20664,N_19163,N_19001);
and U20665 (N_20665,N_19249,N_19762);
and U20666 (N_20666,N_19385,N_19967);
nor U20667 (N_20667,N_19129,N_19959);
or U20668 (N_20668,N_19716,N_19912);
and U20669 (N_20669,N_19193,N_19194);
nor U20670 (N_20670,N_19501,N_19936);
nor U20671 (N_20671,N_19799,N_19782);
nand U20672 (N_20672,N_19061,N_19870);
xnor U20673 (N_20673,N_19269,N_19991);
or U20674 (N_20674,N_19542,N_19116);
nand U20675 (N_20675,N_19030,N_19660);
nand U20676 (N_20676,N_19467,N_19498);
or U20677 (N_20677,N_19673,N_19472);
xnor U20678 (N_20678,N_19532,N_19500);
nor U20679 (N_20679,N_19155,N_19004);
and U20680 (N_20680,N_19292,N_19206);
nand U20681 (N_20681,N_19650,N_19162);
and U20682 (N_20682,N_19628,N_19024);
xor U20683 (N_20683,N_19833,N_19415);
nand U20684 (N_20684,N_19697,N_19761);
or U20685 (N_20685,N_19679,N_19024);
or U20686 (N_20686,N_19755,N_19038);
nand U20687 (N_20687,N_19462,N_19166);
nor U20688 (N_20688,N_19403,N_19617);
or U20689 (N_20689,N_19916,N_19017);
and U20690 (N_20690,N_19015,N_19548);
nand U20691 (N_20691,N_19858,N_19516);
nor U20692 (N_20692,N_19345,N_19289);
and U20693 (N_20693,N_19794,N_19873);
or U20694 (N_20694,N_19883,N_19298);
or U20695 (N_20695,N_19781,N_19273);
and U20696 (N_20696,N_19545,N_19193);
or U20697 (N_20697,N_19580,N_19842);
nand U20698 (N_20698,N_19525,N_19197);
and U20699 (N_20699,N_19593,N_19577);
nand U20700 (N_20700,N_19369,N_19471);
nand U20701 (N_20701,N_19110,N_19687);
nand U20702 (N_20702,N_19775,N_19438);
xnor U20703 (N_20703,N_19592,N_19978);
and U20704 (N_20704,N_19682,N_19361);
nand U20705 (N_20705,N_19064,N_19751);
nor U20706 (N_20706,N_19595,N_19412);
nor U20707 (N_20707,N_19235,N_19842);
xor U20708 (N_20708,N_19687,N_19452);
nand U20709 (N_20709,N_19828,N_19241);
and U20710 (N_20710,N_19064,N_19689);
or U20711 (N_20711,N_19320,N_19395);
nor U20712 (N_20712,N_19297,N_19036);
and U20713 (N_20713,N_19597,N_19851);
and U20714 (N_20714,N_19273,N_19458);
xnor U20715 (N_20715,N_19597,N_19224);
and U20716 (N_20716,N_19371,N_19785);
and U20717 (N_20717,N_19592,N_19788);
or U20718 (N_20718,N_19997,N_19493);
and U20719 (N_20719,N_19277,N_19264);
nand U20720 (N_20720,N_19572,N_19282);
nand U20721 (N_20721,N_19162,N_19593);
xnor U20722 (N_20722,N_19071,N_19833);
nor U20723 (N_20723,N_19661,N_19395);
nor U20724 (N_20724,N_19690,N_19563);
nand U20725 (N_20725,N_19558,N_19486);
or U20726 (N_20726,N_19331,N_19751);
or U20727 (N_20727,N_19242,N_19570);
xor U20728 (N_20728,N_19660,N_19084);
xor U20729 (N_20729,N_19747,N_19168);
or U20730 (N_20730,N_19844,N_19286);
nor U20731 (N_20731,N_19509,N_19739);
nor U20732 (N_20732,N_19104,N_19059);
nor U20733 (N_20733,N_19266,N_19986);
nand U20734 (N_20734,N_19807,N_19025);
nand U20735 (N_20735,N_19617,N_19308);
nand U20736 (N_20736,N_19834,N_19100);
and U20737 (N_20737,N_19034,N_19365);
and U20738 (N_20738,N_19541,N_19188);
nor U20739 (N_20739,N_19666,N_19841);
and U20740 (N_20740,N_19010,N_19271);
nor U20741 (N_20741,N_19630,N_19625);
and U20742 (N_20742,N_19511,N_19604);
or U20743 (N_20743,N_19431,N_19509);
nand U20744 (N_20744,N_19829,N_19447);
and U20745 (N_20745,N_19037,N_19944);
nor U20746 (N_20746,N_19872,N_19036);
and U20747 (N_20747,N_19299,N_19301);
or U20748 (N_20748,N_19308,N_19556);
and U20749 (N_20749,N_19261,N_19501);
nand U20750 (N_20750,N_19264,N_19282);
nor U20751 (N_20751,N_19854,N_19349);
nor U20752 (N_20752,N_19757,N_19418);
xnor U20753 (N_20753,N_19267,N_19607);
or U20754 (N_20754,N_19382,N_19061);
nor U20755 (N_20755,N_19301,N_19627);
or U20756 (N_20756,N_19840,N_19981);
nor U20757 (N_20757,N_19482,N_19432);
xnor U20758 (N_20758,N_19959,N_19979);
or U20759 (N_20759,N_19334,N_19235);
xor U20760 (N_20760,N_19747,N_19286);
nor U20761 (N_20761,N_19987,N_19498);
and U20762 (N_20762,N_19927,N_19601);
nor U20763 (N_20763,N_19847,N_19580);
nand U20764 (N_20764,N_19746,N_19397);
and U20765 (N_20765,N_19043,N_19963);
nand U20766 (N_20766,N_19357,N_19748);
and U20767 (N_20767,N_19026,N_19671);
and U20768 (N_20768,N_19338,N_19711);
and U20769 (N_20769,N_19887,N_19855);
or U20770 (N_20770,N_19739,N_19734);
and U20771 (N_20771,N_19899,N_19542);
xnor U20772 (N_20772,N_19906,N_19557);
nand U20773 (N_20773,N_19354,N_19547);
and U20774 (N_20774,N_19147,N_19562);
xnor U20775 (N_20775,N_19341,N_19689);
or U20776 (N_20776,N_19423,N_19377);
xor U20777 (N_20777,N_19952,N_19826);
and U20778 (N_20778,N_19211,N_19135);
or U20779 (N_20779,N_19273,N_19787);
nor U20780 (N_20780,N_19256,N_19509);
nor U20781 (N_20781,N_19256,N_19602);
xnor U20782 (N_20782,N_19806,N_19172);
and U20783 (N_20783,N_19887,N_19648);
xnor U20784 (N_20784,N_19756,N_19008);
xor U20785 (N_20785,N_19945,N_19752);
nor U20786 (N_20786,N_19566,N_19492);
nor U20787 (N_20787,N_19193,N_19816);
nor U20788 (N_20788,N_19397,N_19800);
nor U20789 (N_20789,N_19343,N_19099);
or U20790 (N_20790,N_19042,N_19125);
and U20791 (N_20791,N_19619,N_19977);
nor U20792 (N_20792,N_19040,N_19597);
xnor U20793 (N_20793,N_19483,N_19235);
and U20794 (N_20794,N_19662,N_19663);
or U20795 (N_20795,N_19764,N_19299);
or U20796 (N_20796,N_19359,N_19085);
or U20797 (N_20797,N_19041,N_19854);
and U20798 (N_20798,N_19869,N_19167);
nor U20799 (N_20799,N_19275,N_19693);
nand U20800 (N_20800,N_19388,N_19531);
and U20801 (N_20801,N_19236,N_19785);
xnor U20802 (N_20802,N_19033,N_19334);
nor U20803 (N_20803,N_19351,N_19094);
or U20804 (N_20804,N_19258,N_19561);
nand U20805 (N_20805,N_19309,N_19024);
and U20806 (N_20806,N_19805,N_19191);
xor U20807 (N_20807,N_19663,N_19750);
nand U20808 (N_20808,N_19579,N_19045);
and U20809 (N_20809,N_19321,N_19752);
xor U20810 (N_20810,N_19962,N_19864);
nor U20811 (N_20811,N_19814,N_19787);
and U20812 (N_20812,N_19856,N_19096);
nor U20813 (N_20813,N_19933,N_19655);
and U20814 (N_20814,N_19377,N_19667);
and U20815 (N_20815,N_19830,N_19743);
xnor U20816 (N_20816,N_19262,N_19080);
or U20817 (N_20817,N_19735,N_19601);
xnor U20818 (N_20818,N_19821,N_19088);
nor U20819 (N_20819,N_19216,N_19521);
and U20820 (N_20820,N_19860,N_19777);
nand U20821 (N_20821,N_19785,N_19905);
nor U20822 (N_20822,N_19194,N_19246);
nor U20823 (N_20823,N_19096,N_19953);
nand U20824 (N_20824,N_19907,N_19659);
nand U20825 (N_20825,N_19755,N_19362);
nand U20826 (N_20826,N_19828,N_19913);
and U20827 (N_20827,N_19131,N_19930);
and U20828 (N_20828,N_19518,N_19599);
nor U20829 (N_20829,N_19881,N_19848);
or U20830 (N_20830,N_19430,N_19711);
or U20831 (N_20831,N_19678,N_19526);
xor U20832 (N_20832,N_19881,N_19205);
and U20833 (N_20833,N_19211,N_19341);
nor U20834 (N_20834,N_19711,N_19630);
nor U20835 (N_20835,N_19484,N_19248);
or U20836 (N_20836,N_19677,N_19332);
and U20837 (N_20837,N_19061,N_19430);
and U20838 (N_20838,N_19776,N_19651);
or U20839 (N_20839,N_19744,N_19168);
or U20840 (N_20840,N_19506,N_19492);
or U20841 (N_20841,N_19552,N_19151);
nand U20842 (N_20842,N_19102,N_19279);
or U20843 (N_20843,N_19339,N_19199);
xor U20844 (N_20844,N_19783,N_19146);
and U20845 (N_20845,N_19923,N_19170);
nor U20846 (N_20846,N_19651,N_19062);
or U20847 (N_20847,N_19269,N_19995);
nand U20848 (N_20848,N_19613,N_19943);
nor U20849 (N_20849,N_19439,N_19614);
and U20850 (N_20850,N_19649,N_19302);
and U20851 (N_20851,N_19272,N_19630);
and U20852 (N_20852,N_19872,N_19748);
nor U20853 (N_20853,N_19221,N_19406);
nor U20854 (N_20854,N_19957,N_19866);
and U20855 (N_20855,N_19937,N_19259);
xnor U20856 (N_20856,N_19334,N_19365);
nand U20857 (N_20857,N_19544,N_19174);
and U20858 (N_20858,N_19775,N_19309);
xor U20859 (N_20859,N_19753,N_19146);
and U20860 (N_20860,N_19687,N_19023);
nor U20861 (N_20861,N_19751,N_19897);
and U20862 (N_20862,N_19334,N_19896);
nand U20863 (N_20863,N_19768,N_19786);
xnor U20864 (N_20864,N_19681,N_19412);
nand U20865 (N_20865,N_19162,N_19124);
and U20866 (N_20866,N_19021,N_19651);
nor U20867 (N_20867,N_19579,N_19040);
nand U20868 (N_20868,N_19091,N_19321);
nor U20869 (N_20869,N_19445,N_19390);
xor U20870 (N_20870,N_19682,N_19241);
xor U20871 (N_20871,N_19706,N_19608);
and U20872 (N_20872,N_19158,N_19905);
nand U20873 (N_20873,N_19264,N_19939);
nor U20874 (N_20874,N_19422,N_19287);
nor U20875 (N_20875,N_19957,N_19152);
xnor U20876 (N_20876,N_19733,N_19673);
nor U20877 (N_20877,N_19442,N_19674);
and U20878 (N_20878,N_19816,N_19365);
and U20879 (N_20879,N_19427,N_19553);
nand U20880 (N_20880,N_19096,N_19937);
xor U20881 (N_20881,N_19132,N_19618);
or U20882 (N_20882,N_19014,N_19861);
nand U20883 (N_20883,N_19108,N_19320);
xor U20884 (N_20884,N_19809,N_19690);
xor U20885 (N_20885,N_19909,N_19001);
nor U20886 (N_20886,N_19896,N_19595);
nor U20887 (N_20887,N_19350,N_19599);
or U20888 (N_20888,N_19558,N_19409);
and U20889 (N_20889,N_19045,N_19705);
or U20890 (N_20890,N_19934,N_19408);
xnor U20891 (N_20891,N_19115,N_19357);
or U20892 (N_20892,N_19874,N_19825);
nand U20893 (N_20893,N_19694,N_19422);
or U20894 (N_20894,N_19820,N_19370);
nand U20895 (N_20895,N_19577,N_19295);
nand U20896 (N_20896,N_19931,N_19718);
xor U20897 (N_20897,N_19451,N_19024);
nor U20898 (N_20898,N_19018,N_19321);
nand U20899 (N_20899,N_19475,N_19714);
and U20900 (N_20900,N_19720,N_19540);
xnor U20901 (N_20901,N_19035,N_19087);
or U20902 (N_20902,N_19163,N_19255);
or U20903 (N_20903,N_19925,N_19800);
nor U20904 (N_20904,N_19827,N_19784);
xnor U20905 (N_20905,N_19005,N_19060);
and U20906 (N_20906,N_19094,N_19778);
xor U20907 (N_20907,N_19491,N_19497);
nor U20908 (N_20908,N_19420,N_19437);
nor U20909 (N_20909,N_19214,N_19082);
and U20910 (N_20910,N_19384,N_19425);
nand U20911 (N_20911,N_19315,N_19646);
xor U20912 (N_20912,N_19231,N_19607);
xnor U20913 (N_20913,N_19187,N_19632);
nor U20914 (N_20914,N_19582,N_19762);
xor U20915 (N_20915,N_19418,N_19863);
nor U20916 (N_20916,N_19258,N_19277);
nor U20917 (N_20917,N_19907,N_19628);
and U20918 (N_20918,N_19071,N_19463);
nand U20919 (N_20919,N_19795,N_19369);
and U20920 (N_20920,N_19735,N_19501);
or U20921 (N_20921,N_19082,N_19357);
xnor U20922 (N_20922,N_19126,N_19839);
xor U20923 (N_20923,N_19070,N_19775);
xor U20924 (N_20924,N_19879,N_19668);
and U20925 (N_20925,N_19405,N_19682);
and U20926 (N_20926,N_19149,N_19637);
nand U20927 (N_20927,N_19537,N_19556);
or U20928 (N_20928,N_19037,N_19651);
nor U20929 (N_20929,N_19346,N_19866);
nor U20930 (N_20930,N_19249,N_19124);
and U20931 (N_20931,N_19709,N_19538);
or U20932 (N_20932,N_19012,N_19394);
nand U20933 (N_20933,N_19209,N_19846);
nand U20934 (N_20934,N_19853,N_19580);
or U20935 (N_20935,N_19228,N_19476);
xnor U20936 (N_20936,N_19020,N_19587);
nand U20937 (N_20937,N_19428,N_19687);
nand U20938 (N_20938,N_19764,N_19671);
nand U20939 (N_20939,N_19837,N_19022);
nand U20940 (N_20940,N_19355,N_19420);
nand U20941 (N_20941,N_19870,N_19059);
nand U20942 (N_20942,N_19015,N_19116);
nand U20943 (N_20943,N_19226,N_19088);
or U20944 (N_20944,N_19968,N_19172);
or U20945 (N_20945,N_19401,N_19773);
xnor U20946 (N_20946,N_19830,N_19551);
nand U20947 (N_20947,N_19340,N_19196);
xor U20948 (N_20948,N_19530,N_19832);
xnor U20949 (N_20949,N_19736,N_19081);
and U20950 (N_20950,N_19808,N_19185);
and U20951 (N_20951,N_19764,N_19086);
nand U20952 (N_20952,N_19045,N_19772);
or U20953 (N_20953,N_19153,N_19211);
nor U20954 (N_20954,N_19979,N_19188);
nand U20955 (N_20955,N_19385,N_19496);
xnor U20956 (N_20956,N_19814,N_19466);
and U20957 (N_20957,N_19846,N_19974);
xor U20958 (N_20958,N_19713,N_19663);
xnor U20959 (N_20959,N_19035,N_19775);
nor U20960 (N_20960,N_19973,N_19908);
or U20961 (N_20961,N_19114,N_19287);
nor U20962 (N_20962,N_19824,N_19643);
and U20963 (N_20963,N_19816,N_19248);
or U20964 (N_20964,N_19311,N_19438);
and U20965 (N_20965,N_19470,N_19353);
nor U20966 (N_20966,N_19098,N_19831);
and U20967 (N_20967,N_19036,N_19955);
and U20968 (N_20968,N_19536,N_19642);
and U20969 (N_20969,N_19850,N_19877);
nor U20970 (N_20970,N_19484,N_19906);
xnor U20971 (N_20971,N_19721,N_19962);
nand U20972 (N_20972,N_19667,N_19821);
and U20973 (N_20973,N_19964,N_19766);
or U20974 (N_20974,N_19079,N_19256);
nand U20975 (N_20975,N_19352,N_19367);
xor U20976 (N_20976,N_19859,N_19058);
nor U20977 (N_20977,N_19623,N_19019);
or U20978 (N_20978,N_19712,N_19814);
nor U20979 (N_20979,N_19176,N_19011);
and U20980 (N_20980,N_19079,N_19193);
nand U20981 (N_20981,N_19843,N_19649);
xor U20982 (N_20982,N_19785,N_19362);
and U20983 (N_20983,N_19854,N_19122);
nand U20984 (N_20984,N_19339,N_19360);
nand U20985 (N_20985,N_19836,N_19478);
nand U20986 (N_20986,N_19672,N_19015);
nand U20987 (N_20987,N_19182,N_19123);
xnor U20988 (N_20988,N_19487,N_19799);
or U20989 (N_20989,N_19167,N_19665);
and U20990 (N_20990,N_19659,N_19678);
nor U20991 (N_20991,N_19139,N_19987);
or U20992 (N_20992,N_19137,N_19456);
xor U20993 (N_20993,N_19826,N_19682);
or U20994 (N_20994,N_19050,N_19393);
or U20995 (N_20995,N_19073,N_19758);
nor U20996 (N_20996,N_19528,N_19766);
or U20997 (N_20997,N_19977,N_19102);
xnor U20998 (N_20998,N_19844,N_19163);
nor U20999 (N_20999,N_19805,N_19433);
or U21000 (N_21000,N_20272,N_20798);
and U21001 (N_21001,N_20984,N_20691);
or U21002 (N_21002,N_20139,N_20213);
xnor U21003 (N_21003,N_20434,N_20048);
nor U21004 (N_21004,N_20853,N_20449);
and U21005 (N_21005,N_20134,N_20135);
nor U21006 (N_21006,N_20712,N_20929);
or U21007 (N_21007,N_20520,N_20343);
and U21008 (N_21008,N_20173,N_20211);
or U21009 (N_21009,N_20558,N_20465);
nand U21010 (N_21010,N_20540,N_20112);
nor U21011 (N_21011,N_20522,N_20001);
nor U21012 (N_21012,N_20000,N_20258);
or U21013 (N_21013,N_20072,N_20519);
xnor U21014 (N_21014,N_20829,N_20324);
nor U21015 (N_21015,N_20504,N_20336);
or U21016 (N_21016,N_20153,N_20689);
and U21017 (N_21017,N_20536,N_20709);
nor U21018 (N_21018,N_20468,N_20070);
nand U21019 (N_21019,N_20802,N_20813);
nand U21020 (N_21020,N_20163,N_20919);
nor U21021 (N_21021,N_20222,N_20552);
nor U21022 (N_21022,N_20470,N_20989);
or U21023 (N_21023,N_20482,N_20198);
and U21024 (N_21024,N_20484,N_20042);
nor U21025 (N_21025,N_20777,N_20553);
nand U21026 (N_21026,N_20035,N_20859);
or U21027 (N_21027,N_20964,N_20085);
or U21028 (N_21028,N_20566,N_20022);
and U21029 (N_21029,N_20227,N_20711);
or U21030 (N_21030,N_20422,N_20341);
or U21031 (N_21031,N_20843,N_20573);
and U21032 (N_21032,N_20684,N_20956);
nor U21033 (N_21033,N_20381,N_20763);
and U21034 (N_21034,N_20426,N_20122);
xor U21035 (N_21035,N_20062,N_20037);
nand U21036 (N_21036,N_20697,N_20026);
nand U21037 (N_21037,N_20496,N_20330);
or U21038 (N_21038,N_20963,N_20845);
nor U21039 (N_21039,N_20665,N_20832);
nor U21040 (N_21040,N_20148,N_20460);
or U21041 (N_21041,N_20841,N_20823);
and U21042 (N_21042,N_20888,N_20351);
and U21043 (N_21043,N_20701,N_20389);
nor U21044 (N_21044,N_20946,N_20523);
nor U21045 (N_21045,N_20215,N_20359);
nor U21046 (N_21046,N_20095,N_20912);
nor U21047 (N_21047,N_20957,N_20782);
xnor U21048 (N_21048,N_20795,N_20855);
xor U21049 (N_21049,N_20738,N_20725);
nand U21050 (N_21050,N_20203,N_20528);
and U21051 (N_21051,N_20995,N_20291);
and U21052 (N_21052,N_20113,N_20883);
nor U21053 (N_21053,N_20831,N_20298);
or U21054 (N_21054,N_20108,N_20694);
or U21055 (N_21055,N_20366,N_20078);
nand U21056 (N_21056,N_20145,N_20052);
xor U21057 (N_21057,N_20962,N_20115);
nand U21058 (N_21058,N_20388,N_20880);
nand U21059 (N_21059,N_20918,N_20350);
nand U21060 (N_21060,N_20539,N_20089);
xnor U21061 (N_21061,N_20983,N_20507);
and U21062 (N_21062,N_20877,N_20737);
xnor U21063 (N_21063,N_20819,N_20127);
and U21064 (N_21064,N_20043,N_20086);
xor U21065 (N_21065,N_20172,N_20270);
or U21066 (N_21066,N_20727,N_20276);
nand U21067 (N_21067,N_20615,N_20734);
or U21068 (N_21068,N_20164,N_20966);
nand U21069 (N_21069,N_20891,N_20401);
nor U21070 (N_21070,N_20597,N_20560);
or U21071 (N_21071,N_20892,N_20419);
and U21072 (N_21072,N_20921,N_20331);
nand U21073 (N_21073,N_20011,N_20472);
and U21074 (N_21074,N_20290,N_20809);
and U21075 (N_21075,N_20093,N_20194);
and U21076 (N_21076,N_20879,N_20865);
xor U21077 (N_21077,N_20474,N_20128);
or U21078 (N_21078,N_20099,N_20981);
or U21079 (N_21079,N_20774,N_20947);
and U21080 (N_21080,N_20352,N_20041);
xnor U21081 (N_21081,N_20609,N_20317);
nand U21082 (N_21082,N_20620,N_20284);
and U21083 (N_21083,N_20817,N_20903);
nand U21084 (N_21084,N_20444,N_20882);
or U21085 (N_21085,N_20543,N_20610);
nor U21086 (N_21086,N_20100,N_20742);
and U21087 (N_21087,N_20126,N_20902);
and U21088 (N_21088,N_20047,N_20618);
nand U21089 (N_21089,N_20844,N_20458);
nand U21090 (N_21090,N_20471,N_20051);
nand U21091 (N_21091,N_20822,N_20236);
xor U21092 (N_21092,N_20308,N_20762);
or U21093 (N_21093,N_20379,N_20658);
xor U21094 (N_21094,N_20239,N_20915);
and U21095 (N_21095,N_20028,N_20197);
nand U21096 (N_21096,N_20590,N_20629);
nor U21097 (N_21097,N_20327,N_20955);
nor U21098 (N_21098,N_20717,N_20600);
xnor U21099 (N_21099,N_20881,N_20268);
nor U21100 (N_21100,N_20116,N_20174);
or U21101 (N_21101,N_20289,N_20636);
xor U21102 (N_21102,N_20008,N_20369);
xor U21103 (N_21103,N_20740,N_20791);
and U21104 (N_21104,N_20716,N_20923);
and U21105 (N_21105,N_20110,N_20820);
and U21106 (N_21106,N_20541,N_20954);
nand U21107 (N_21107,N_20747,N_20598);
or U21108 (N_21108,N_20431,N_20358);
nor U21109 (N_21109,N_20514,N_20154);
and U21110 (N_21110,N_20617,N_20023);
nor U21111 (N_21111,N_20524,N_20733);
or U21112 (N_21112,N_20288,N_20337);
nor U21113 (N_21113,N_20825,N_20186);
and U21114 (N_21114,N_20538,N_20924);
nor U21115 (N_21115,N_20249,N_20643);
xnor U21116 (N_21116,N_20578,N_20776);
xor U21117 (N_21117,N_20207,N_20715);
nor U21118 (N_21118,N_20025,N_20094);
xnor U21119 (N_21119,N_20621,N_20703);
and U21120 (N_21120,N_20259,N_20926);
or U21121 (N_21121,N_20098,N_20155);
nor U21122 (N_21122,N_20058,N_20370);
nor U21123 (N_21123,N_20840,N_20282);
nor U21124 (N_21124,N_20296,N_20147);
and U21125 (N_21125,N_20015,N_20457);
nor U21126 (N_21126,N_20124,N_20220);
xor U21127 (N_21127,N_20107,N_20306);
xor U21128 (N_21128,N_20916,N_20205);
xnor U21129 (N_21129,N_20446,N_20392);
and U21130 (N_21130,N_20890,N_20430);
or U21131 (N_21131,N_20645,N_20451);
nor U21132 (N_21132,N_20726,N_20714);
or U21133 (N_21133,N_20068,N_20548);
or U21134 (N_21134,N_20050,N_20906);
xor U21135 (N_21135,N_20150,N_20669);
nor U21136 (N_21136,N_20624,N_20517);
or U21137 (N_21137,N_20410,N_20441);
xor U21138 (N_21138,N_20602,N_20167);
xnor U21139 (N_21139,N_20391,N_20861);
nor U21140 (N_21140,N_20132,N_20732);
nor U21141 (N_21141,N_20250,N_20547);
nor U21142 (N_21142,N_20265,N_20065);
nand U21143 (N_21143,N_20077,N_20469);
nor U21144 (N_21144,N_20481,N_20297);
or U21145 (N_21145,N_20644,N_20187);
nor U21146 (N_21146,N_20907,N_20349);
or U21147 (N_21147,N_20599,N_20530);
or U21148 (N_21148,N_20494,N_20261);
nor U21149 (N_21149,N_20944,N_20729);
nor U21150 (N_21150,N_20873,N_20666);
or U21151 (N_21151,N_20778,N_20661);
or U21152 (N_21152,N_20818,N_20588);
nor U21153 (N_21153,N_20679,N_20483);
and U21154 (N_21154,N_20235,N_20142);
and U21155 (N_21155,N_20651,N_20013);
xnor U21156 (N_21156,N_20057,N_20273);
nand U21157 (N_21157,N_20593,N_20529);
nand U21158 (N_21158,N_20020,N_20283);
nor U21159 (N_21159,N_20866,N_20997);
nor U21160 (N_21160,N_20695,N_20439);
nand U21161 (N_21161,N_20887,N_20503);
or U21162 (N_21162,N_20269,N_20302);
xor U21163 (N_21163,N_20869,N_20580);
nand U21164 (N_21164,N_20850,N_20626);
xor U21165 (N_21165,N_20931,N_20973);
nand U21166 (N_21166,N_20794,N_20678);
nand U21167 (N_21167,N_20189,N_20753);
nand U21168 (N_21168,N_20546,N_20648);
xor U21169 (N_21169,N_20980,N_20071);
xnor U21170 (N_21170,N_20839,N_20313);
nor U21171 (N_21171,N_20698,N_20429);
and U21172 (N_21172,N_20649,N_20216);
nor U21173 (N_21173,N_20511,N_20061);
and U21174 (N_21174,N_20664,N_20908);
nor U21175 (N_21175,N_20642,N_20165);
nand U21176 (N_21176,N_20413,N_20252);
and U21177 (N_21177,N_20886,N_20545);
xor U21178 (N_21178,N_20206,N_20638);
nand U21179 (N_21179,N_20510,N_20835);
and U21180 (N_21180,N_20316,N_20899);
xor U21181 (N_21181,N_20253,N_20033);
nor U21182 (N_21182,N_20385,N_20069);
nor U21183 (N_21183,N_20785,N_20526);
xor U21184 (N_21184,N_20575,N_20895);
or U21185 (N_21185,N_20491,N_20550);
nand U21186 (N_21186,N_20299,N_20828);
nor U21187 (N_21187,N_20783,N_20376);
and U21188 (N_21188,N_20506,N_20581);
or U21189 (N_21189,N_20192,N_20953);
or U21190 (N_21190,N_20990,N_20281);
and U21191 (N_21191,N_20579,N_20260);
xnor U21192 (N_21192,N_20927,N_20415);
nor U21193 (N_21193,N_20554,N_20394);
nand U21194 (N_21194,N_20488,N_20613);
nand U21195 (N_21195,N_20743,N_20685);
or U21196 (N_21196,N_20427,N_20897);
nand U21197 (N_21197,N_20606,N_20893);
and U21198 (N_21198,N_20007,N_20745);
or U21199 (N_21199,N_20706,N_20960);
nand U21200 (N_21200,N_20243,N_20119);
xor U21201 (N_21201,N_20162,N_20262);
or U21202 (N_21202,N_20278,N_20495);
nand U21203 (N_21203,N_20380,N_20399);
nor U21204 (N_21204,N_20979,N_20943);
or U21205 (N_21205,N_20190,N_20571);
nor U21206 (N_21206,N_20467,N_20386);
xor U21207 (N_21207,N_20994,N_20544);
nor U21208 (N_21208,N_20117,N_20219);
nand U21209 (N_21209,N_20237,N_20287);
and U21210 (N_21210,N_20871,N_20965);
nand U21211 (N_21211,N_20209,N_20567);
and U21212 (N_21212,N_20799,N_20251);
and U21213 (N_21213,N_20012,N_20787);
nor U21214 (N_21214,N_20789,N_20583);
nand U21215 (N_21215,N_20564,N_20502);
xor U21216 (N_21216,N_20464,N_20218);
xnor U21217 (N_21217,N_20801,N_20466);
and U21218 (N_21218,N_20286,N_20988);
nor U21219 (N_21219,N_20499,N_20238);
and U21220 (N_21220,N_20367,N_20682);
or U21221 (N_21221,N_20838,N_20807);
or U21222 (N_21222,N_20797,N_20130);
xor U21223 (N_21223,N_20310,N_20784);
nand U21224 (N_21224,N_20757,N_20687);
xnor U21225 (N_21225,N_20295,N_20992);
xnor U21226 (N_21226,N_20199,N_20515);
or U21227 (N_21227,N_20775,N_20677);
xnor U21228 (N_21228,N_20076,N_20404);
nor U21229 (N_21229,N_20447,N_20991);
nor U21230 (N_21230,N_20676,N_20241);
and U21231 (N_21231,N_20796,N_20834);
nor U21232 (N_21232,N_20372,N_20030);
nand U21233 (N_21233,N_20650,N_20329);
nor U21234 (N_21234,N_20565,N_20029);
or U21235 (N_21235,N_20229,N_20898);
xor U21236 (N_21236,N_20555,N_20166);
xor U21237 (N_21237,N_20326,N_20101);
xnor U21238 (N_21238,N_20300,N_20263);
nor U21239 (N_21239,N_20074,N_20905);
nor U21240 (N_21240,N_20371,N_20179);
nor U21241 (N_21241,N_20788,N_20088);
nor U21242 (N_21242,N_20445,N_20004);
nor U21243 (N_21243,N_20479,N_20563);
nor U21244 (N_21244,N_20138,N_20443);
nor U21245 (N_21245,N_20950,N_20040);
or U21246 (N_21246,N_20700,N_20756);
nand U21247 (N_21247,N_20357,N_20136);
or U21248 (N_21248,N_20945,N_20793);
and U21249 (N_21249,N_20630,N_20628);
and U21250 (N_21250,N_20623,N_20059);
or U21251 (N_21251,N_20005,N_20081);
nand U21252 (N_21252,N_20746,N_20006);
nand U21253 (N_21253,N_20605,N_20103);
nand U21254 (N_21254,N_20884,N_20417);
nand U21255 (N_21255,N_20156,N_20056);
or U21256 (N_21256,N_20513,N_20152);
nor U21257 (N_21257,N_20731,N_20346);
nor U21258 (N_21258,N_20083,N_20568);
nor U21259 (N_21259,N_20224,N_20201);
and U21260 (N_21260,N_20937,N_20455);
xor U21261 (N_21261,N_20333,N_20585);
xnor U21262 (N_21262,N_20724,N_20910);
and U21263 (N_21263,N_20305,N_20368);
nand U21264 (N_21264,N_20653,N_20312);
nand U21265 (N_21265,N_20266,N_20010);
xor U21266 (N_21266,N_20377,N_20752);
or U21267 (N_21267,N_20525,N_20728);
nor U21268 (N_21268,N_20200,N_20125);
and U21269 (N_21269,N_20473,N_20275);
nand U21270 (N_21270,N_20781,N_20292);
nand U21271 (N_21271,N_20332,N_20655);
nor U21272 (N_21272,N_20017,N_20255);
nor U21273 (N_21273,N_20181,N_20384);
xor U21274 (N_21274,N_20492,N_20812);
nor U21275 (N_21275,N_20111,N_20364);
nor U21276 (N_21276,N_20196,N_20137);
or U21277 (N_21277,N_20120,N_20815);
and U21278 (N_21278,N_20208,N_20378);
or U21279 (N_21279,N_20739,N_20987);
and U21280 (N_21280,N_20911,N_20003);
nand U21281 (N_21281,N_20978,N_20750);
nor U21282 (N_21282,N_20875,N_20018);
xnor U21283 (N_21283,N_20293,N_20240);
nor U21284 (N_21284,N_20395,N_20667);
nor U21285 (N_21285,N_20896,N_20972);
and U21286 (N_21286,N_20827,N_20044);
and U21287 (N_21287,N_20158,N_20505);
and U21288 (N_21288,N_20940,N_20195);
and U21289 (N_21289,N_20149,N_20039);
or U21290 (N_21290,N_20254,N_20758);
nor U21291 (N_21291,N_20748,N_20670);
nand U21292 (N_21292,N_20692,N_20055);
and U21293 (N_21293,N_20084,N_20486);
or U21294 (N_21294,N_20914,N_20870);
and U21295 (N_21295,N_20452,N_20212);
nor U21296 (N_21296,N_20542,N_20141);
xor U21297 (N_21297,N_20217,N_20177);
and U21298 (N_21298,N_20722,N_20414);
nand U21299 (N_21299,N_20450,N_20402);
and U21300 (N_21300,N_20334,N_20245);
nor U21301 (N_21301,N_20938,N_20968);
xnor U21302 (N_21302,N_20925,N_20398);
and U21303 (N_21303,N_20633,N_20425);
nor U21304 (N_21304,N_20230,N_20967);
nor U21305 (N_21305,N_20970,N_20002);
nor U21306 (N_21306,N_20675,N_20151);
and U21307 (N_21307,N_20267,N_20683);
nor U21308 (N_21308,N_20744,N_20982);
nor U21309 (N_21309,N_20647,N_20833);
and U21310 (N_21310,N_20348,N_20941);
or U21311 (N_21311,N_20713,N_20193);
nand U21312 (N_21312,N_20314,N_20779);
nor U21313 (N_21313,N_20347,N_20390);
or U21314 (N_21314,N_20080,N_20109);
nor U21315 (N_21315,N_20031,N_20920);
nand U21316 (N_21316,N_20885,N_20014);
xnor U21317 (N_21317,N_20027,N_20864);
xnor U21318 (N_21318,N_20420,N_20614);
and U21319 (N_21319,N_20512,N_20894);
or U21320 (N_21320,N_20418,N_20387);
xnor U21321 (N_21321,N_20688,N_20680);
nor U21322 (N_21322,N_20604,N_20256);
nand U21323 (N_21323,N_20355,N_20718);
and U21324 (N_21324,N_20274,N_20021);
nand U21325 (N_21325,N_20632,N_20285);
nor U21326 (N_21326,N_20416,N_20169);
xor U21327 (N_21327,N_20860,N_20131);
and U21328 (N_21328,N_20092,N_20456);
xnor U21329 (N_21329,N_20721,N_20303);
or U21330 (N_21330,N_20971,N_20674);
nand U21331 (N_21331,N_20900,N_20659);
nor U21332 (N_21332,N_20533,N_20400);
xor U21333 (N_21333,N_20765,N_20656);
and U21334 (N_21334,N_20475,N_20320);
nor U21335 (N_21335,N_20304,N_20323);
or U21336 (N_21336,N_20339,N_20766);
nor U21337 (N_21337,N_20639,N_20720);
or U21338 (N_21338,N_20576,N_20168);
and U21339 (N_21339,N_20657,N_20814);
nor U21340 (N_21340,N_20719,N_20360);
or U21341 (N_21341,N_20662,N_20143);
nand U21342 (N_21342,N_20868,N_20949);
xor U21343 (N_21343,N_20811,N_20928);
nor U21344 (N_21344,N_20338,N_20612);
xor U21345 (N_21345,N_20102,N_20437);
or U21346 (N_21346,N_20671,N_20448);
nand U21347 (N_21347,N_20397,N_20064);
nand U21348 (N_21348,N_20878,N_20476);
nand U21349 (N_21349,N_20363,N_20096);
nand U21350 (N_21350,N_20409,N_20403);
xnor U21351 (N_21351,N_20705,N_20374);
xor U21352 (N_21352,N_20279,N_20232);
xor U21353 (N_21353,N_20595,N_20749);
nand U21354 (N_21354,N_20591,N_20913);
nand U21355 (N_21355,N_20462,N_20412);
and U21356 (N_21356,N_20821,N_20951);
or U21357 (N_21357,N_20611,N_20231);
or U21358 (N_21358,N_20325,N_20764);
and U21359 (N_21359,N_20247,N_20375);
nand U21360 (N_21360,N_20534,N_20551);
xnor U21361 (N_21361,N_20640,N_20693);
nor U21362 (N_21362,N_20622,N_20559);
or U21363 (N_21363,N_20408,N_20652);
xnor U21364 (N_21364,N_20114,N_20681);
nor U21365 (N_21365,N_20161,N_20046);
nor U21366 (N_21366,N_20959,N_20301);
xnor U21367 (N_21367,N_20532,N_20406);
and U21368 (N_21368,N_20038,N_20735);
nand U21369 (N_21369,N_20271,N_20867);
xor U21370 (N_21370,N_20608,N_20019);
nand U21371 (N_21371,N_20311,N_20436);
and U21372 (N_21372,N_20660,N_20454);
nor U21373 (N_21373,N_20998,N_20075);
nand U21374 (N_21374,N_20922,N_20889);
nor U21375 (N_21375,N_20561,N_20294);
and U21376 (N_21376,N_20985,N_20383);
nand U21377 (N_21377,N_20699,N_20986);
nor U21378 (N_21378,N_20234,N_20405);
xor U21379 (N_21379,N_20751,N_20362);
or U21380 (N_21380,N_20354,N_20631);
or U21381 (N_21381,N_20257,N_20690);
nand U21382 (N_21382,N_20607,N_20790);
nand U21383 (N_21383,N_20625,N_20060);
nor U21384 (N_21384,N_20036,N_20862);
xor U21385 (N_21385,N_20121,N_20053);
or U21386 (N_21386,N_20948,N_20184);
nor U21387 (N_21387,N_20210,N_20993);
xnor U21388 (N_21388,N_20863,N_20569);
xnor U21389 (N_21389,N_20175,N_20182);
nor U21390 (N_21390,N_20668,N_20754);
or U21391 (N_21391,N_20577,N_20932);
nand U21392 (N_21392,N_20340,N_20857);
nand U21393 (N_21393,N_20936,N_20485);
xor U21394 (N_21394,N_20999,N_20616);
nand U21395 (N_21395,N_20328,N_20773);
and U21396 (N_21396,N_20854,N_20307);
and U21397 (N_21397,N_20342,N_20826);
xor U21398 (N_21398,N_20248,N_20091);
nor U21399 (N_21399,N_20942,N_20535);
xor U21400 (N_21400,N_20180,N_20803);
nor U21401 (N_21401,N_20702,N_20562);
xnor U21402 (N_21402,N_20453,N_20780);
and U21403 (N_21403,N_20244,N_20961);
nand U21404 (N_21404,N_20277,N_20759);
or U21405 (N_21405,N_20518,N_20601);
and U21406 (N_21406,N_20501,N_20202);
nand U21407 (N_21407,N_20584,N_20309);
xor U21408 (N_21408,N_20160,N_20438);
nand U21409 (N_21409,N_20423,N_20958);
xnor U21410 (N_21410,N_20901,N_20393);
xor U21411 (N_21411,N_20837,N_20373);
and U21412 (N_21412,N_20846,N_20847);
and U21413 (N_21413,N_20516,N_20531);
or U21414 (N_21414,N_20140,N_20586);
nand U21415 (N_21415,N_20767,N_20549);
or U21416 (N_21416,N_20769,N_20032);
nor U21417 (N_21417,N_20975,N_20170);
and U21418 (N_21418,N_20741,N_20952);
and U21419 (N_21419,N_20480,N_20365);
nor U21420 (N_21420,N_20489,N_20433);
nor U21421 (N_21421,N_20233,N_20396);
nor U21422 (N_21422,N_20498,N_20521);
nand U21423 (N_21423,N_20129,N_20428);
and U21424 (N_21424,N_20345,N_20223);
xor U21425 (N_21425,N_20185,N_20106);
and U21426 (N_21426,N_20707,N_20382);
or U21427 (N_21427,N_20090,N_20497);
xnor U21428 (N_21428,N_20315,N_20063);
and U21429 (N_21429,N_20634,N_20214);
or U21430 (N_21430,N_20808,N_20183);
nand U21431 (N_21431,N_20917,N_20939);
nand U21432 (N_21432,N_20073,N_20730);
and U21433 (N_21433,N_20146,N_20318);
and U21434 (N_21434,N_20572,N_20459);
xnor U21435 (N_21435,N_20874,N_20582);
xor U21436 (N_21436,N_20490,N_20344);
xnor U21437 (N_21437,N_20087,N_20105);
nor U21438 (N_21438,N_20704,N_20619);
nand U21439 (N_21439,N_20442,N_20144);
nand U21440 (N_21440,N_20188,N_20977);
nand U21441 (N_21441,N_20710,N_20356);
nor U21442 (N_21442,N_20641,N_20574);
nor U21443 (N_21443,N_20432,N_20935);
nor U21444 (N_21444,N_20596,N_20852);
nor U21445 (N_21445,N_20876,N_20934);
xnor U21446 (N_21446,N_20280,N_20104);
and U21447 (N_21447,N_20335,N_20673);
and U21448 (N_21448,N_20487,N_20755);
nand U21449 (N_21449,N_20570,N_20800);
nor U21450 (N_21450,N_20723,N_20556);
nor U21451 (N_21451,N_20176,N_20221);
or U21452 (N_21452,N_20016,N_20171);
nand U21453 (N_21453,N_20082,N_20696);
nand U21454 (N_21454,N_20191,N_20974);
nor U21455 (N_21455,N_20816,N_20440);
or U21456 (N_21456,N_20157,N_20830);
and U21457 (N_21457,N_20411,N_20909);
or U21458 (N_21458,N_20654,N_20225);
and U21459 (N_21459,N_20603,N_20435);
nand U21460 (N_21460,N_20461,N_20768);
nand U21461 (N_21461,N_20672,N_20204);
or U21462 (N_21462,N_20079,N_20933);
and U21463 (N_21463,N_20858,N_20594);
nor U21464 (N_21464,N_20477,N_20500);
nor U21465 (N_21465,N_20804,N_20627);
nand U21466 (N_21466,N_20592,N_20463);
xnor U21467 (N_21467,N_20049,N_20904);
or U21468 (N_21468,N_20322,N_20361);
and U21469 (N_21469,N_20848,N_20066);
xor U21470 (N_21470,N_20424,N_20509);
xor U21471 (N_21471,N_20242,N_20537);
nand U21472 (N_21472,N_20123,N_20319);
xor U21473 (N_21473,N_20637,N_20805);
nand U21474 (N_21474,N_20067,N_20824);
or U21475 (N_21475,N_20045,N_20508);
nand U21476 (N_21476,N_20527,N_20034);
and U21477 (N_21477,N_20407,N_20770);
nor U21478 (N_21478,N_20663,N_20024);
or U21479 (N_21479,N_20226,N_20589);
nor U21480 (N_21480,N_20761,N_20806);
xor U21481 (N_21481,N_20786,N_20493);
nand U21482 (N_21482,N_20930,N_20771);
or U21483 (N_21483,N_20842,N_20421);
nand U21484 (N_21484,N_20228,N_20054);
nand U21485 (N_21485,N_20264,N_20133);
and U21486 (N_21486,N_20760,N_20353);
nor U21487 (N_21487,N_20810,N_20478);
or U21488 (N_21488,N_20849,N_20686);
and U21489 (N_21489,N_20736,N_20557);
nand U21490 (N_21490,N_20321,N_20836);
or U21491 (N_21491,N_20996,N_20246);
nand U21492 (N_21492,N_20009,N_20969);
and U21493 (N_21493,N_20178,N_20851);
nand U21494 (N_21494,N_20635,N_20708);
or U21495 (N_21495,N_20856,N_20792);
nor U21496 (N_21496,N_20118,N_20097);
or U21497 (N_21497,N_20646,N_20587);
and U21498 (N_21498,N_20159,N_20772);
nand U21499 (N_21499,N_20872,N_20976);
and U21500 (N_21500,N_20257,N_20983);
nor U21501 (N_21501,N_20886,N_20646);
nand U21502 (N_21502,N_20105,N_20212);
or U21503 (N_21503,N_20103,N_20943);
nand U21504 (N_21504,N_20711,N_20878);
xnor U21505 (N_21505,N_20504,N_20056);
nor U21506 (N_21506,N_20728,N_20504);
or U21507 (N_21507,N_20774,N_20349);
nor U21508 (N_21508,N_20896,N_20019);
nor U21509 (N_21509,N_20465,N_20153);
nand U21510 (N_21510,N_20107,N_20211);
and U21511 (N_21511,N_20585,N_20578);
nor U21512 (N_21512,N_20777,N_20144);
and U21513 (N_21513,N_20429,N_20966);
nand U21514 (N_21514,N_20431,N_20623);
nand U21515 (N_21515,N_20900,N_20036);
nand U21516 (N_21516,N_20028,N_20256);
nand U21517 (N_21517,N_20578,N_20045);
nand U21518 (N_21518,N_20185,N_20391);
nor U21519 (N_21519,N_20165,N_20040);
xnor U21520 (N_21520,N_20326,N_20218);
or U21521 (N_21521,N_20370,N_20765);
and U21522 (N_21522,N_20830,N_20324);
or U21523 (N_21523,N_20746,N_20950);
nor U21524 (N_21524,N_20348,N_20328);
nand U21525 (N_21525,N_20222,N_20067);
or U21526 (N_21526,N_20534,N_20238);
xnor U21527 (N_21527,N_20321,N_20036);
or U21528 (N_21528,N_20519,N_20967);
nor U21529 (N_21529,N_20793,N_20042);
nand U21530 (N_21530,N_20738,N_20581);
and U21531 (N_21531,N_20952,N_20727);
nor U21532 (N_21532,N_20673,N_20731);
and U21533 (N_21533,N_20563,N_20927);
or U21534 (N_21534,N_20991,N_20019);
xnor U21535 (N_21535,N_20405,N_20866);
nand U21536 (N_21536,N_20561,N_20983);
xor U21537 (N_21537,N_20541,N_20314);
xor U21538 (N_21538,N_20004,N_20414);
or U21539 (N_21539,N_20055,N_20372);
nor U21540 (N_21540,N_20165,N_20896);
xnor U21541 (N_21541,N_20204,N_20382);
xor U21542 (N_21542,N_20776,N_20970);
xor U21543 (N_21543,N_20975,N_20384);
xor U21544 (N_21544,N_20386,N_20272);
nand U21545 (N_21545,N_20000,N_20346);
xor U21546 (N_21546,N_20707,N_20255);
and U21547 (N_21547,N_20240,N_20210);
or U21548 (N_21548,N_20280,N_20668);
nand U21549 (N_21549,N_20569,N_20488);
or U21550 (N_21550,N_20129,N_20044);
or U21551 (N_21551,N_20092,N_20564);
or U21552 (N_21552,N_20838,N_20540);
or U21553 (N_21553,N_20712,N_20273);
nor U21554 (N_21554,N_20386,N_20830);
and U21555 (N_21555,N_20127,N_20993);
xnor U21556 (N_21556,N_20858,N_20412);
nand U21557 (N_21557,N_20566,N_20594);
xnor U21558 (N_21558,N_20133,N_20010);
and U21559 (N_21559,N_20859,N_20220);
nor U21560 (N_21560,N_20302,N_20158);
nand U21561 (N_21561,N_20363,N_20920);
xnor U21562 (N_21562,N_20763,N_20891);
nand U21563 (N_21563,N_20834,N_20861);
nor U21564 (N_21564,N_20511,N_20360);
or U21565 (N_21565,N_20722,N_20845);
or U21566 (N_21566,N_20928,N_20750);
or U21567 (N_21567,N_20640,N_20524);
nand U21568 (N_21568,N_20751,N_20195);
xor U21569 (N_21569,N_20728,N_20045);
and U21570 (N_21570,N_20888,N_20145);
and U21571 (N_21571,N_20243,N_20236);
and U21572 (N_21572,N_20485,N_20835);
nor U21573 (N_21573,N_20580,N_20920);
and U21574 (N_21574,N_20338,N_20577);
xor U21575 (N_21575,N_20853,N_20426);
or U21576 (N_21576,N_20493,N_20018);
xnor U21577 (N_21577,N_20722,N_20274);
nand U21578 (N_21578,N_20257,N_20788);
xnor U21579 (N_21579,N_20621,N_20570);
nand U21580 (N_21580,N_20448,N_20213);
and U21581 (N_21581,N_20288,N_20595);
nand U21582 (N_21582,N_20700,N_20084);
and U21583 (N_21583,N_20556,N_20476);
or U21584 (N_21584,N_20432,N_20675);
or U21585 (N_21585,N_20461,N_20482);
or U21586 (N_21586,N_20417,N_20448);
nor U21587 (N_21587,N_20601,N_20066);
and U21588 (N_21588,N_20797,N_20329);
and U21589 (N_21589,N_20673,N_20000);
and U21590 (N_21590,N_20379,N_20603);
nand U21591 (N_21591,N_20656,N_20562);
nand U21592 (N_21592,N_20550,N_20982);
nand U21593 (N_21593,N_20202,N_20594);
nand U21594 (N_21594,N_20730,N_20462);
xnor U21595 (N_21595,N_20508,N_20689);
xor U21596 (N_21596,N_20901,N_20802);
nor U21597 (N_21597,N_20618,N_20919);
and U21598 (N_21598,N_20956,N_20524);
and U21599 (N_21599,N_20647,N_20531);
and U21600 (N_21600,N_20583,N_20623);
and U21601 (N_21601,N_20197,N_20317);
or U21602 (N_21602,N_20011,N_20959);
or U21603 (N_21603,N_20987,N_20151);
nand U21604 (N_21604,N_20190,N_20455);
nand U21605 (N_21605,N_20425,N_20314);
nor U21606 (N_21606,N_20656,N_20187);
nor U21607 (N_21607,N_20305,N_20341);
nand U21608 (N_21608,N_20324,N_20776);
nand U21609 (N_21609,N_20782,N_20666);
xor U21610 (N_21610,N_20544,N_20091);
and U21611 (N_21611,N_20462,N_20271);
nor U21612 (N_21612,N_20045,N_20521);
nor U21613 (N_21613,N_20970,N_20902);
xor U21614 (N_21614,N_20355,N_20600);
nand U21615 (N_21615,N_20421,N_20382);
xnor U21616 (N_21616,N_20554,N_20129);
nand U21617 (N_21617,N_20441,N_20575);
nand U21618 (N_21618,N_20060,N_20419);
and U21619 (N_21619,N_20978,N_20338);
xnor U21620 (N_21620,N_20124,N_20169);
xnor U21621 (N_21621,N_20982,N_20242);
nand U21622 (N_21622,N_20221,N_20555);
or U21623 (N_21623,N_20213,N_20806);
and U21624 (N_21624,N_20304,N_20060);
nand U21625 (N_21625,N_20420,N_20423);
and U21626 (N_21626,N_20541,N_20901);
nor U21627 (N_21627,N_20386,N_20828);
nor U21628 (N_21628,N_20062,N_20287);
or U21629 (N_21629,N_20253,N_20551);
nor U21630 (N_21630,N_20417,N_20453);
xor U21631 (N_21631,N_20544,N_20613);
and U21632 (N_21632,N_20765,N_20467);
nand U21633 (N_21633,N_20355,N_20578);
or U21634 (N_21634,N_20800,N_20083);
and U21635 (N_21635,N_20863,N_20123);
or U21636 (N_21636,N_20344,N_20392);
nand U21637 (N_21637,N_20942,N_20699);
and U21638 (N_21638,N_20501,N_20545);
nor U21639 (N_21639,N_20938,N_20907);
or U21640 (N_21640,N_20024,N_20613);
nor U21641 (N_21641,N_20444,N_20997);
or U21642 (N_21642,N_20835,N_20841);
nand U21643 (N_21643,N_20324,N_20862);
nor U21644 (N_21644,N_20769,N_20239);
xor U21645 (N_21645,N_20614,N_20899);
xor U21646 (N_21646,N_20137,N_20217);
nand U21647 (N_21647,N_20956,N_20207);
xor U21648 (N_21648,N_20214,N_20919);
and U21649 (N_21649,N_20530,N_20236);
nor U21650 (N_21650,N_20098,N_20265);
xnor U21651 (N_21651,N_20834,N_20428);
or U21652 (N_21652,N_20563,N_20348);
nand U21653 (N_21653,N_20420,N_20785);
nand U21654 (N_21654,N_20180,N_20231);
nand U21655 (N_21655,N_20509,N_20198);
and U21656 (N_21656,N_20838,N_20931);
nor U21657 (N_21657,N_20459,N_20186);
xnor U21658 (N_21658,N_20982,N_20545);
nand U21659 (N_21659,N_20058,N_20849);
nand U21660 (N_21660,N_20002,N_20800);
nand U21661 (N_21661,N_20505,N_20364);
and U21662 (N_21662,N_20617,N_20477);
or U21663 (N_21663,N_20699,N_20314);
xnor U21664 (N_21664,N_20823,N_20635);
nand U21665 (N_21665,N_20366,N_20789);
or U21666 (N_21666,N_20024,N_20625);
nor U21667 (N_21667,N_20471,N_20315);
nor U21668 (N_21668,N_20381,N_20599);
and U21669 (N_21669,N_20629,N_20803);
and U21670 (N_21670,N_20013,N_20718);
and U21671 (N_21671,N_20229,N_20698);
xor U21672 (N_21672,N_20004,N_20521);
nand U21673 (N_21673,N_20139,N_20337);
xor U21674 (N_21674,N_20815,N_20698);
and U21675 (N_21675,N_20703,N_20079);
nand U21676 (N_21676,N_20127,N_20597);
nand U21677 (N_21677,N_20567,N_20210);
and U21678 (N_21678,N_20569,N_20278);
xnor U21679 (N_21679,N_20879,N_20114);
or U21680 (N_21680,N_20694,N_20463);
or U21681 (N_21681,N_20466,N_20298);
xnor U21682 (N_21682,N_20448,N_20802);
and U21683 (N_21683,N_20094,N_20342);
nor U21684 (N_21684,N_20145,N_20705);
and U21685 (N_21685,N_20241,N_20534);
nor U21686 (N_21686,N_20128,N_20617);
nand U21687 (N_21687,N_20818,N_20486);
xor U21688 (N_21688,N_20498,N_20578);
and U21689 (N_21689,N_20289,N_20262);
nand U21690 (N_21690,N_20817,N_20180);
nor U21691 (N_21691,N_20287,N_20173);
xor U21692 (N_21692,N_20754,N_20348);
xor U21693 (N_21693,N_20295,N_20047);
xnor U21694 (N_21694,N_20421,N_20806);
and U21695 (N_21695,N_20863,N_20927);
or U21696 (N_21696,N_20011,N_20020);
or U21697 (N_21697,N_20822,N_20930);
nand U21698 (N_21698,N_20051,N_20994);
or U21699 (N_21699,N_20453,N_20615);
and U21700 (N_21700,N_20268,N_20511);
or U21701 (N_21701,N_20358,N_20195);
and U21702 (N_21702,N_20526,N_20728);
xor U21703 (N_21703,N_20297,N_20941);
nor U21704 (N_21704,N_20032,N_20085);
xor U21705 (N_21705,N_20846,N_20694);
or U21706 (N_21706,N_20775,N_20912);
or U21707 (N_21707,N_20953,N_20050);
and U21708 (N_21708,N_20252,N_20064);
nor U21709 (N_21709,N_20076,N_20373);
xor U21710 (N_21710,N_20149,N_20597);
and U21711 (N_21711,N_20743,N_20987);
nand U21712 (N_21712,N_20258,N_20201);
or U21713 (N_21713,N_20676,N_20478);
nand U21714 (N_21714,N_20229,N_20623);
xor U21715 (N_21715,N_20428,N_20762);
or U21716 (N_21716,N_20409,N_20097);
and U21717 (N_21717,N_20352,N_20990);
nor U21718 (N_21718,N_20698,N_20928);
and U21719 (N_21719,N_20334,N_20805);
or U21720 (N_21720,N_20517,N_20333);
nand U21721 (N_21721,N_20724,N_20671);
nand U21722 (N_21722,N_20309,N_20331);
or U21723 (N_21723,N_20442,N_20876);
nand U21724 (N_21724,N_20377,N_20059);
xnor U21725 (N_21725,N_20917,N_20220);
and U21726 (N_21726,N_20198,N_20179);
nor U21727 (N_21727,N_20067,N_20984);
or U21728 (N_21728,N_20947,N_20721);
xnor U21729 (N_21729,N_20258,N_20747);
and U21730 (N_21730,N_20942,N_20710);
xor U21731 (N_21731,N_20993,N_20677);
nor U21732 (N_21732,N_20060,N_20237);
nor U21733 (N_21733,N_20063,N_20020);
and U21734 (N_21734,N_20655,N_20166);
and U21735 (N_21735,N_20092,N_20968);
xnor U21736 (N_21736,N_20145,N_20698);
xnor U21737 (N_21737,N_20820,N_20690);
nor U21738 (N_21738,N_20635,N_20241);
nand U21739 (N_21739,N_20136,N_20436);
or U21740 (N_21740,N_20277,N_20274);
xnor U21741 (N_21741,N_20340,N_20084);
nand U21742 (N_21742,N_20556,N_20712);
xor U21743 (N_21743,N_20473,N_20210);
or U21744 (N_21744,N_20941,N_20940);
and U21745 (N_21745,N_20331,N_20659);
and U21746 (N_21746,N_20963,N_20415);
nand U21747 (N_21747,N_20435,N_20357);
nand U21748 (N_21748,N_20164,N_20193);
nand U21749 (N_21749,N_20246,N_20980);
xor U21750 (N_21750,N_20587,N_20019);
xor U21751 (N_21751,N_20586,N_20363);
nand U21752 (N_21752,N_20054,N_20870);
xor U21753 (N_21753,N_20203,N_20455);
nor U21754 (N_21754,N_20860,N_20253);
nand U21755 (N_21755,N_20944,N_20746);
or U21756 (N_21756,N_20166,N_20602);
and U21757 (N_21757,N_20370,N_20694);
nor U21758 (N_21758,N_20550,N_20689);
or U21759 (N_21759,N_20186,N_20751);
or U21760 (N_21760,N_20086,N_20734);
nand U21761 (N_21761,N_20979,N_20102);
nor U21762 (N_21762,N_20121,N_20671);
nand U21763 (N_21763,N_20526,N_20696);
and U21764 (N_21764,N_20508,N_20453);
and U21765 (N_21765,N_20530,N_20922);
nand U21766 (N_21766,N_20335,N_20888);
xnor U21767 (N_21767,N_20265,N_20380);
or U21768 (N_21768,N_20727,N_20845);
and U21769 (N_21769,N_20890,N_20877);
and U21770 (N_21770,N_20117,N_20414);
nor U21771 (N_21771,N_20782,N_20204);
xnor U21772 (N_21772,N_20960,N_20882);
or U21773 (N_21773,N_20088,N_20939);
xor U21774 (N_21774,N_20247,N_20154);
and U21775 (N_21775,N_20349,N_20686);
or U21776 (N_21776,N_20838,N_20969);
nand U21777 (N_21777,N_20017,N_20979);
nor U21778 (N_21778,N_20752,N_20204);
nor U21779 (N_21779,N_20986,N_20530);
and U21780 (N_21780,N_20675,N_20988);
nand U21781 (N_21781,N_20836,N_20726);
and U21782 (N_21782,N_20896,N_20231);
and U21783 (N_21783,N_20105,N_20354);
xnor U21784 (N_21784,N_20130,N_20703);
and U21785 (N_21785,N_20946,N_20011);
nand U21786 (N_21786,N_20682,N_20224);
or U21787 (N_21787,N_20713,N_20994);
xor U21788 (N_21788,N_20138,N_20182);
nor U21789 (N_21789,N_20013,N_20946);
nor U21790 (N_21790,N_20114,N_20004);
nor U21791 (N_21791,N_20647,N_20902);
nand U21792 (N_21792,N_20399,N_20521);
nand U21793 (N_21793,N_20089,N_20731);
and U21794 (N_21794,N_20414,N_20219);
nand U21795 (N_21795,N_20250,N_20194);
and U21796 (N_21796,N_20118,N_20084);
xnor U21797 (N_21797,N_20151,N_20464);
xnor U21798 (N_21798,N_20158,N_20127);
nor U21799 (N_21799,N_20088,N_20307);
and U21800 (N_21800,N_20681,N_20425);
and U21801 (N_21801,N_20177,N_20432);
nand U21802 (N_21802,N_20528,N_20255);
nand U21803 (N_21803,N_20731,N_20131);
xor U21804 (N_21804,N_20230,N_20386);
and U21805 (N_21805,N_20239,N_20214);
or U21806 (N_21806,N_20347,N_20887);
nand U21807 (N_21807,N_20026,N_20255);
and U21808 (N_21808,N_20333,N_20519);
nor U21809 (N_21809,N_20135,N_20698);
and U21810 (N_21810,N_20299,N_20570);
or U21811 (N_21811,N_20154,N_20599);
xnor U21812 (N_21812,N_20148,N_20513);
or U21813 (N_21813,N_20694,N_20607);
nand U21814 (N_21814,N_20789,N_20287);
nand U21815 (N_21815,N_20426,N_20647);
nand U21816 (N_21816,N_20470,N_20373);
and U21817 (N_21817,N_20110,N_20906);
xnor U21818 (N_21818,N_20876,N_20847);
nor U21819 (N_21819,N_20369,N_20048);
or U21820 (N_21820,N_20339,N_20788);
nand U21821 (N_21821,N_20799,N_20878);
nand U21822 (N_21822,N_20376,N_20196);
nand U21823 (N_21823,N_20411,N_20177);
xnor U21824 (N_21824,N_20330,N_20930);
xnor U21825 (N_21825,N_20506,N_20979);
nand U21826 (N_21826,N_20082,N_20840);
or U21827 (N_21827,N_20559,N_20399);
or U21828 (N_21828,N_20612,N_20618);
or U21829 (N_21829,N_20523,N_20391);
or U21830 (N_21830,N_20778,N_20877);
or U21831 (N_21831,N_20971,N_20330);
xor U21832 (N_21832,N_20333,N_20337);
or U21833 (N_21833,N_20348,N_20908);
nor U21834 (N_21834,N_20240,N_20292);
and U21835 (N_21835,N_20153,N_20342);
or U21836 (N_21836,N_20101,N_20128);
or U21837 (N_21837,N_20068,N_20651);
nand U21838 (N_21838,N_20731,N_20865);
nor U21839 (N_21839,N_20146,N_20914);
xor U21840 (N_21840,N_20589,N_20644);
nand U21841 (N_21841,N_20995,N_20634);
nor U21842 (N_21842,N_20470,N_20450);
and U21843 (N_21843,N_20075,N_20433);
nor U21844 (N_21844,N_20690,N_20702);
xor U21845 (N_21845,N_20244,N_20360);
and U21846 (N_21846,N_20631,N_20473);
xor U21847 (N_21847,N_20492,N_20087);
nor U21848 (N_21848,N_20859,N_20664);
nor U21849 (N_21849,N_20469,N_20181);
nor U21850 (N_21850,N_20000,N_20312);
xnor U21851 (N_21851,N_20532,N_20776);
and U21852 (N_21852,N_20151,N_20855);
nand U21853 (N_21853,N_20345,N_20096);
or U21854 (N_21854,N_20620,N_20280);
and U21855 (N_21855,N_20761,N_20007);
or U21856 (N_21856,N_20049,N_20161);
nand U21857 (N_21857,N_20015,N_20180);
or U21858 (N_21858,N_20778,N_20832);
or U21859 (N_21859,N_20868,N_20098);
xnor U21860 (N_21860,N_20172,N_20788);
or U21861 (N_21861,N_20884,N_20546);
nor U21862 (N_21862,N_20812,N_20814);
xor U21863 (N_21863,N_20468,N_20444);
nand U21864 (N_21864,N_20959,N_20659);
nand U21865 (N_21865,N_20963,N_20139);
xor U21866 (N_21866,N_20570,N_20416);
xor U21867 (N_21867,N_20568,N_20486);
nor U21868 (N_21868,N_20568,N_20132);
nand U21869 (N_21869,N_20166,N_20451);
nand U21870 (N_21870,N_20203,N_20408);
nor U21871 (N_21871,N_20982,N_20704);
and U21872 (N_21872,N_20344,N_20947);
and U21873 (N_21873,N_20894,N_20619);
nor U21874 (N_21874,N_20314,N_20386);
or U21875 (N_21875,N_20819,N_20094);
xnor U21876 (N_21876,N_20057,N_20823);
nand U21877 (N_21877,N_20976,N_20171);
and U21878 (N_21878,N_20444,N_20030);
nand U21879 (N_21879,N_20588,N_20198);
or U21880 (N_21880,N_20629,N_20256);
nor U21881 (N_21881,N_20204,N_20573);
nand U21882 (N_21882,N_20690,N_20737);
nand U21883 (N_21883,N_20703,N_20384);
xnor U21884 (N_21884,N_20881,N_20051);
nor U21885 (N_21885,N_20272,N_20218);
nand U21886 (N_21886,N_20535,N_20832);
nor U21887 (N_21887,N_20221,N_20534);
nor U21888 (N_21888,N_20278,N_20822);
or U21889 (N_21889,N_20382,N_20375);
nand U21890 (N_21890,N_20031,N_20640);
nor U21891 (N_21891,N_20077,N_20984);
nand U21892 (N_21892,N_20802,N_20656);
nor U21893 (N_21893,N_20399,N_20957);
nand U21894 (N_21894,N_20105,N_20877);
or U21895 (N_21895,N_20867,N_20999);
or U21896 (N_21896,N_20426,N_20435);
and U21897 (N_21897,N_20910,N_20236);
xor U21898 (N_21898,N_20437,N_20436);
and U21899 (N_21899,N_20077,N_20443);
nand U21900 (N_21900,N_20617,N_20603);
and U21901 (N_21901,N_20024,N_20650);
xor U21902 (N_21902,N_20801,N_20407);
xor U21903 (N_21903,N_20714,N_20708);
xnor U21904 (N_21904,N_20211,N_20464);
nand U21905 (N_21905,N_20082,N_20076);
xor U21906 (N_21906,N_20912,N_20235);
or U21907 (N_21907,N_20738,N_20121);
xor U21908 (N_21908,N_20825,N_20407);
and U21909 (N_21909,N_20620,N_20512);
nand U21910 (N_21910,N_20137,N_20534);
nand U21911 (N_21911,N_20940,N_20244);
xnor U21912 (N_21912,N_20864,N_20147);
nand U21913 (N_21913,N_20748,N_20202);
xnor U21914 (N_21914,N_20839,N_20179);
nor U21915 (N_21915,N_20587,N_20282);
nand U21916 (N_21916,N_20979,N_20773);
or U21917 (N_21917,N_20213,N_20552);
nor U21918 (N_21918,N_20233,N_20003);
nor U21919 (N_21919,N_20156,N_20009);
nor U21920 (N_21920,N_20327,N_20642);
and U21921 (N_21921,N_20423,N_20346);
xnor U21922 (N_21922,N_20466,N_20002);
xor U21923 (N_21923,N_20086,N_20808);
xor U21924 (N_21924,N_20506,N_20509);
or U21925 (N_21925,N_20708,N_20606);
nor U21926 (N_21926,N_20669,N_20846);
or U21927 (N_21927,N_20112,N_20795);
xnor U21928 (N_21928,N_20608,N_20697);
xnor U21929 (N_21929,N_20345,N_20685);
nand U21930 (N_21930,N_20696,N_20703);
and U21931 (N_21931,N_20072,N_20224);
xor U21932 (N_21932,N_20813,N_20194);
and U21933 (N_21933,N_20428,N_20071);
or U21934 (N_21934,N_20599,N_20099);
nand U21935 (N_21935,N_20460,N_20971);
or U21936 (N_21936,N_20761,N_20080);
nor U21937 (N_21937,N_20793,N_20411);
nor U21938 (N_21938,N_20910,N_20981);
nor U21939 (N_21939,N_20346,N_20415);
and U21940 (N_21940,N_20973,N_20400);
and U21941 (N_21941,N_20117,N_20702);
nand U21942 (N_21942,N_20685,N_20842);
and U21943 (N_21943,N_20453,N_20438);
xor U21944 (N_21944,N_20545,N_20383);
xnor U21945 (N_21945,N_20396,N_20755);
xor U21946 (N_21946,N_20712,N_20843);
and U21947 (N_21947,N_20279,N_20335);
and U21948 (N_21948,N_20114,N_20403);
and U21949 (N_21949,N_20135,N_20736);
nor U21950 (N_21950,N_20281,N_20414);
nor U21951 (N_21951,N_20603,N_20216);
nand U21952 (N_21952,N_20617,N_20830);
and U21953 (N_21953,N_20585,N_20416);
nor U21954 (N_21954,N_20322,N_20236);
and U21955 (N_21955,N_20158,N_20494);
or U21956 (N_21956,N_20515,N_20215);
xor U21957 (N_21957,N_20484,N_20166);
nor U21958 (N_21958,N_20164,N_20674);
or U21959 (N_21959,N_20459,N_20371);
and U21960 (N_21960,N_20832,N_20741);
nor U21961 (N_21961,N_20708,N_20689);
xor U21962 (N_21962,N_20976,N_20188);
or U21963 (N_21963,N_20533,N_20439);
or U21964 (N_21964,N_20001,N_20053);
nor U21965 (N_21965,N_20234,N_20731);
or U21966 (N_21966,N_20390,N_20565);
nand U21967 (N_21967,N_20484,N_20293);
and U21968 (N_21968,N_20686,N_20371);
xnor U21969 (N_21969,N_20631,N_20750);
or U21970 (N_21970,N_20069,N_20902);
nor U21971 (N_21971,N_20480,N_20821);
or U21972 (N_21972,N_20399,N_20897);
xnor U21973 (N_21973,N_20654,N_20757);
and U21974 (N_21974,N_20345,N_20089);
xor U21975 (N_21975,N_20937,N_20944);
xnor U21976 (N_21976,N_20310,N_20910);
or U21977 (N_21977,N_20062,N_20895);
and U21978 (N_21978,N_20813,N_20129);
xnor U21979 (N_21979,N_20683,N_20005);
nor U21980 (N_21980,N_20810,N_20750);
or U21981 (N_21981,N_20031,N_20421);
nor U21982 (N_21982,N_20534,N_20042);
and U21983 (N_21983,N_20199,N_20331);
nand U21984 (N_21984,N_20834,N_20752);
nor U21985 (N_21985,N_20151,N_20760);
xnor U21986 (N_21986,N_20419,N_20062);
or U21987 (N_21987,N_20686,N_20210);
nor U21988 (N_21988,N_20455,N_20368);
or U21989 (N_21989,N_20387,N_20324);
or U21990 (N_21990,N_20649,N_20903);
nand U21991 (N_21991,N_20284,N_20137);
nor U21992 (N_21992,N_20988,N_20009);
nor U21993 (N_21993,N_20600,N_20076);
and U21994 (N_21994,N_20181,N_20542);
xor U21995 (N_21995,N_20929,N_20988);
xor U21996 (N_21996,N_20030,N_20088);
nor U21997 (N_21997,N_20516,N_20650);
nor U21998 (N_21998,N_20629,N_20282);
or U21999 (N_21999,N_20795,N_20917);
and U22000 (N_22000,N_21545,N_21343);
nor U22001 (N_22001,N_21188,N_21586);
and U22002 (N_22002,N_21975,N_21938);
or U22003 (N_22003,N_21385,N_21052);
and U22004 (N_22004,N_21452,N_21147);
or U22005 (N_22005,N_21522,N_21762);
and U22006 (N_22006,N_21799,N_21252);
and U22007 (N_22007,N_21443,N_21595);
nor U22008 (N_22008,N_21139,N_21968);
nand U22009 (N_22009,N_21940,N_21227);
or U22010 (N_22010,N_21064,N_21041);
and U22011 (N_22011,N_21539,N_21246);
xor U22012 (N_22012,N_21202,N_21901);
nor U22013 (N_22013,N_21504,N_21319);
nand U22014 (N_22014,N_21137,N_21196);
xnor U22015 (N_22015,N_21836,N_21873);
or U22016 (N_22016,N_21007,N_21379);
and U22017 (N_22017,N_21008,N_21301);
and U22018 (N_22018,N_21528,N_21014);
xor U22019 (N_22019,N_21791,N_21328);
xor U22020 (N_22020,N_21541,N_21006);
and U22021 (N_22021,N_21620,N_21814);
xnor U22022 (N_22022,N_21375,N_21792);
nand U22023 (N_22023,N_21451,N_21396);
and U22024 (N_22024,N_21412,N_21480);
nand U22025 (N_22025,N_21662,N_21200);
nor U22026 (N_22026,N_21436,N_21768);
or U22027 (N_22027,N_21894,N_21497);
nand U22028 (N_22028,N_21341,N_21135);
or U22029 (N_22029,N_21761,N_21323);
and U22030 (N_22030,N_21760,N_21141);
nand U22031 (N_22031,N_21566,N_21399);
nor U22032 (N_22032,N_21699,N_21066);
nand U22033 (N_22033,N_21616,N_21228);
or U22034 (N_22034,N_21303,N_21548);
nor U22035 (N_22035,N_21454,N_21963);
and U22036 (N_22036,N_21384,N_21287);
nand U22037 (N_22037,N_21868,N_21306);
xnor U22038 (N_22038,N_21839,N_21780);
or U22039 (N_22039,N_21476,N_21063);
nand U22040 (N_22040,N_21523,N_21819);
nor U22041 (N_22041,N_21872,N_21828);
or U22042 (N_22042,N_21101,N_21832);
or U22043 (N_22043,N_21980,N_21646);
and U22044 (N_22044,N_21499,N_21992);
and U22045 (N_22045,N_21989,N_21233);
and U22046 (N_22046,N_21296,N_21648);
or U22047 (N_22047,N_21182,N_21720);
xor U22048 (N_22048,N_21298,N_21735);
xor U22049 (N_22049,N_21218,N_21338);
or U22050 (N_22050,N_21840,N_21517);
nor U22051 (N_22051,N_21487,N_21891);
xnor U22052 (N_22052,N_21515,N_21494);
nor U22053 (N_22053,N_21903,N_21425);
or U22054 (N_22054,N_21837,N_21361);
nand U22055 (N_22055,N_21352,N_21171);
nand U22056 (N_22056,N_21689,N_21194);
nand U22057 (N_22057,N_21776,N_21278);
xor U22058 (N_22058,N_21823,N_21329);
nand U22059 (N_22059,N_21160,N_21580);
and U22060 (N_22060,N_21048,N_21906);
nand U22061 (N_22061,N_21897,N_21677);
or U22062 (N_22062,N_21815,N_21559);
and U22063 (N_22063,N_21473,N_21021);
xnor U22064 (N_22064,N_21433,N_21603);
and U22065 (N_22065,N_21082,N_21702);
nand U22066 (N_22066,N_21056,N_21138);
nand U22067 (N_22067,N_21697,N_21337);
nand U22068 (N_22068,N_21299,N_21125);
xnor U22069 (N_22069,N_21964,N_21054);
nor U22070 (N_22070,N_21513,N_21681);
nand U22071 (N_22071,N_21250,N_21251);
xor U22072 (N_22072,N_21459,N_21393);
nand U22073 (N_22073,N_21816,N_21865);
nand U22074 (N_22074,N_21952,N_21929);
nor U22075 (N_22075,N_21093,N_21498);
nand U22076 (N_22076,N_21569,N_21464);
xor U22077 (N_22077,N_21033,N_21954);
and U22078 (N_22078,N_21059,N_21268);
and U22079 (N_22079,N_21267,N_21055);
xor U22080 (N_22080,N_21178,N_21594);
or U22081 (N_22081,N_21684,N_21009);
or U22082 (N_22082,N_21564,N_21700);
or U22083 (N_22083,N_21547,N_21416);
nand U22084 (N_22084,N_21358,N_21560);
and U22085 (N_22085,N_21982,N_21411);
nor U22086 (N_22086,N_21856,N_21095);
nor U22087 (N_22087,N_21265,N_21822);
nand U22088 (N_22088,N_21479,N_21482);
or U22089 (N_22089,N_21167,N_21225);
and U22090 (N_22090,N_21809,N_21861);
nand U22091 (N_22091,N_21496,N_21575);
nand U22092 (N_22092,N_21849,N_21979);
nand U22093 (N_22093,N_21049,N_21269);
nor U22094 (N_22094,N_21474,N_21893);
nor U22095 (N_22095,N_21653,N_21552);
nand U22096 (N_22096,N_21585,N_21676);
nand U22097 (N_22097,N_21530,N_21026);
nand U22098 (N_22098,N_21829,N_21945);
xor U22099 (N_22099,N_21333,N_21180);
nand U22100 (N_22100,N_21773,N_21161);
nand U22101 (N_22101,N_21036,N_21288);
and U22102 (N_22102,N_21405,N_21234);
and U22103 (N_22103,N_21775,N_21902);
xnor U22104 (N_22104,N_21395,N_21132);
nor U22105 (N_22105,N_21781,N_21350);
or U22106 (N_22106,N_21942,N_21658);
or U22107 (N_22107,N_21119,N_21624);
xor U22108 (N_22108,N_21802,N_21495);
nand U22109 (N_22109,N_21285,N_21181);
xnor U22110 (N_22110,N_21738,N_21165);
or U22111 (N_22111,N_21198,N_21308);
and U22112 (N_22112,N_21630,N_21596);
nor U22113 (N_22113,N_21568,N_21870);
xnor U22114 (N_22114,N_21788,N_21953);
nand U22115 (N_22115,N_21888,N_21882);
and U22116 (N_22116,N_21898,N_21919);
nand U22117 (N_22117,N_21877,N_21549);
nor U22118 (N_22118,N_21998,N_21294);
nand U22119 (N_22119,N_21001,N_21824);
or U22120 (N_22120,N_21544,N_21766);
xnor U22121 (N_22121,N_21205,N_21310);
or U22122 (N_22122,N_21053,N_21020);
nand U22123 (N_22123,N_21555,N_21364);
or U22124 (N_22124,N_21332,N_21561);
nand U22125 (N_22125,N_21032,N_21626);
nor U22126 (N_22126,N_21440,N_21483);
and U22127 (N_22127,N_21857,N_21912);
xnor U22128 (N_22128,N_21793,N_21346);
xnor U22129 (N_22129,N_21633,N_21214);
nor U22130 (N_22130,N_21850,N_21907);
or U22131 (N_22131,N_21543,N_21531);
nor U22132 (N_22132,N_21605,N_21074);
or U22133 (N_22133,N_21261,N_21068);
nor U22134 (N_22134,N_21157,N_21121);
nand U22135 (N_22135,N_21537,N_21102);
nand U22136 (N_22136,N_21509,N_21748);
nand U22137 (N_22137,N_21712,N_21086);
nand U22138 (N_22138,N_21974,N_21862);
and U22139 (N_22139,N_21217,N_21719);
or U22140 (N_22140,N_21330,N_21737);
or U22141 (N_22141,N_21471,N_21270);
nand U22142 (N_22142,N_21682,N_21441);
and U22143 (N_22143,N_21711,N_21804);
and U22144 (N_22144,N_21300,N_21223);
or U22145 (N_22145,N_21229,N_21935);
and U22146 (N_22146,N_21327,N_21576);
nand U22147 (N_22147,N_21211,N_21191);
or U22148 (N_22148,N_21415,N_21455);
nand U22149 (N_22149,N_21149,N_21623);
and U22150 (N_22150,N_21860,N_21869);
xor U22151 (N_22151,N_21800,N_21029);
nand U22152 (N_22152,N_21978,N_21146);
or U22153 (N_22153,N_21371,N_21625);
nor U22154 (N_22154,N_21686,N_21256);
nand U22155 (N_22155,N_21209,N_21127);
nor U22156 (N_22156,N_21602,N_21820);
nor U22157 (N_22157,N_21988,N_21004);
or U22158 (N_22158,N_21790,N_21264);
or U22159 (N_22159,N_21615,N_21900);
or U22160 (N_22160,N_21619,N_21947);
or U22161 (N_22161,N_21599,N_21842);
xnor U22162 (N_22162,N_21279,N_21739);
and U22163 (N_22163,N_21601,N_21273);
and U22164 (N_22164,N_21282,N_21673);
nor U22165 (N_22165,N_21466,N_21959);
xor U22166 (N_22166,N_21750,N_21812);
nand U22167 (N_22167,N_21520,N_21117);
xor U22168 (N_22168,N_21172,N_21481);
xnor U22169 (N_22169,N_21290,N_21448);
nor U22170 (N_22170,N_21166,N_21846);
nor U22171 (N_22171,N_21920,N_21022);
nand U22172 (N_22172,N_21113,N_21116);
and U22173 (N_22173,N_21084,N_21948);
and U22174 (N_22174,N_21755,N_21219);
or U22175 (N_22175,N_21707,N_21307);
xor U22176 (N_22176,N_21075,N_21694);
xor U22177 (N_22177,N_21216,N_21174);
nand U22178 (N_22178,N_21195,N_21691);
xor U22179 (N_22179,N_21142,N_21011);
and U22180 (N_22180,N_21969,N_21749);
and U22181 (N_22181,N_21933,N_21756);
nor U22182 (N_22182,N_21374,N_21176);
xnor U22183 (N_22183,N_21394,N_21248);
xnor U22184 (N_22184,N_21345,N_21035);
or U22185 (N_22185,N_21321,N_21342);
nor U22186 (N_22186,N_21960,N_21999);
nand U22187 (N_22187,N_21771,N_21003);
nand U22188 (N_22188,N_21263,N_21987);
xor U22189 (N_22189,N_21642,N_21631);
or U22190 (N_22190,N_21058,N_21918);
or U22191 (N_22191,N_21883,N_21511);
nor U22192 (N_22192,N_21302,N_21462);
or U22193 (N_22193,N_21449,N_21659);
and U22194 (N_22194,N_21597,N_21221);
nand U22195 (N_22195,N_21796,N_21500);
nor U22196 (N_22196,N_21914,N_21984);
or U22197 (N_22197,N_21478,N_21420);
and U22198 (N_22198,N_21372,N_21851);
or U22199 (N_22199,N_21281,N_21240);
nor U22200 (N_22200,N_21028,N_21885);
nor U22201 (N_22201,N_21716,N_21928);
or U22202 (N_22202,N_21986,N_21734);
xnor U22203 (N_22203,N_21508,N_21104);
xor U22204 (N_22204,N_21810,N_21667);
and U22205 (N_22205,N_21752,N_21617);
nor U22206 (N_22206,N_21985,N_21419);
or U22207 (N_22207,N_21946,N_21365);
nand U22208 (N_22208,N_21746,N_21961);
nand U22209 (N_22209,N_21852,N_21593);
or U22210 (N_22210,N_21542,N_21239);
xor U22211 (N_22211,N_21930,N_21878);
xnor U22212 (N_22212,N_21859,N_21271);
nand U22213 (N_22213,N_21778,N_21971);
nor U22214 (N_22214,N_21108,N_21962);
nand U22215 (N_22215,N_21051,N_21636);
or U22216 (N_22216,N_21997,N_21613);
nor U22217 (N_22217,N_21817,N_21787);
xnor U22218 (N_22218,N_21621,N_21030);
and U22219 (N_22219,N_21351,N_21944);
nand U22220 (N_22220,N_21638,N_21785);
nand U22221 (N_22221,N_21806,N_21422);
xor U22222 (N_22222,N_21512,N_21406);
xnor U22223 (N_22223,N_21841,N_21732);
xor U22224 (N_22224,N_21484,N_21789);
nand U22225 (N_22225,N_21805,N_21465);
and U22226 (N_22226,N_21100,N_21743);
or U22227 (N_22227,N_21794,N_21879);
or U22228 (N_22228,N_21591,N_21316);
nand U22229 (N_22229,N_21115,N_21320);
or U22230 (N_22230,N_21254,N_21450);
and U22231 (N_22231,N_21916,N_21641);
and U22232 (N_22232,N_21204,N_21129);
or U22233 (N_22233,N_21931,N_21589);
or U22234 (N_22234,N_21065,N_21460);
and U22235 (N_22235,N_21297,N_21925);
and U22236 (N_22236,N_21243,N_21939);
or U22237 (N_22237,N_21016,N_21486);
nand U22238 (N_22238,N_21803,N_21808);
nand U22239 (N_22239,N_21884,N_21220);
or U22240 (N_22240,N_21098,N_21164);
nor U22241 (N_22241,N_21610,N_21527);
nor U22242 (N_22242,N_21255,N_21538);
and U22243 (N_22243,N_21380,N_21991);
and U22244 (N_22244,N_21490,N_21833);
nor U22245 (N_22245,N_21249,N_21366);
nor U22246 (N_22246,N_21259,N_21057);
or U22247 (N_22247,N_21190,N_21876);
nand U22248 (N_22248,N_21091,N_21661);
nand U22249 (N_22249,N_21344,N_21177);
nor U22250 (N_22250,N_21525,N_21072);
xor U22251 (N_22251,N_21736,N_21587);
nand U22252 (N_22252,N_21370,N_21578);
nand U22253 (N_22253,N_21040,N_21764);
nand U22254 (N_22254,N_21854,N_21050);
and U22255 (N_22255,N_21604,N_21671);
xor U22256 (N_22256,N_21521,N_21210);
nor U22257 (N_22257,N_21280,N_21044);
nor U22258 (N_22258,N_21077,N_21286);
nand U22259 (N_22259,N_21643,N_21080);
or U22260 (N_22260,N_21242,N_21253);
nand U22261 (N_22261,N_21418,N_21145);
nand U22262 (N_22262,N_21027,N_21453);
nor U22263 (N_22263,N_21292,N_21845);
nor U22264 (N_22264,N_21083,N_21213);
xnor U22265 (N_22265,N_21070,N_21696);
and U22266 (N_22266,N_21688,N_21073);
xnor U22267 (N_22267,N_21915,N_21314);
nor U22268 (N_22268,N_21170,N_21786);
nand U22269 (N_22269,N_21231,N_21598);
nand U22270 (N_22270,N_21921,N_21359);
nand U22271 (N_22271,N_21046,N_21990);
nand U22272 (N_22272,N_21956,N_21038);
xnor U22273 (N_22273,N_21703,N_21488);
or U22274 (N_22274,N_21154,N_21363);
nand U22275 (N_22275,N_21524,N_21047);
nand U22276 (N_22276,N_21133,N_21535);
or U22277 (N_22277,N_21144,N_21612);
nor U22278 (N_22278,N_21042,N_21391);
nor U22279 (N_22279,N_21304,N_21197);
and U22280 (N_22280,N_21140,N_21967);
nor U22281 (N_22281,N_21556,N_21112);
nand U22282 (N_22282,N_21740,N_21401);
and U22283 (N_22283,N_21501,N_21326);
and U22284 (N_22284,N_21582,N_21122);
nand U22285 (N_22285,N_21187,N_21774);
or U22286 (N_22286,N_21710,N_21431);
and U22287 (N_22287,N_21571,N_21890);
or U22288 (N_22288,N_21291,N_21693);
and U22289 (N_22289,N_21018,N_21715);
nor U22290 (N_22290,N_21034,N_21163);
nand U22291 (N_22291,N_21640,N_21238);
nor U22292 (N_22292,N_21927,N_21705);
or U22293 (N_22293,N_21503,N_21784);
nor U22294 (N_22294,N_21446,N_21674);
and U22295 (N_22295,N_21650,N_21472);
nand U22296 (N_22296,N_21505,N_21934);
nor U22297 (N_22297,N_21099,N_21444);
nor U22298 (N_22298,N_21002,N_21169);
nor U22299 (N_22299,N_21305,N_21972);
and U22300 (N_22300,N_21722,N_21708);
and U22301 (N_22301,N_21655,N_21754);
nand U22302 (N_22302,N_21728,N_21356);
nor U22303 (N_22303,N_21324,N_21461);
or U22304 (N_22304,N_21844,N_21120);
or U22305 (N_22305,N_21097,N_21657);
nor U22306 (N_22306,N_21423,N_21043);
and U22307 (N_22307,N_21143,N_21647);
nand U22308 (N_22308,N_21367,N_21215);
or U22309 (N_22309,N_21409,N_21895);
nor U22310 (N_22310,N_21000,N_21212);
nand U22311 (N_22311,N_21434,N_21069);
nor U22312 (N_22312,N_21519,N_21562);
and U22313 (N_22313,N_21362,N_21574);
xor U22314 (N_22314,N_21744,N_21880);
nor U22315 (N_22315,N_21896,N_21089);
and U22316 (N_22316,N_21622,N_21039);
or U22317 (N_22317,N_21996,N_21680);
nor U22318 (N_22318,N_21311,N_21349);
nor U22319 (N_22319,N_21600,N_21772);
nand U22320 (N_22320,N_21148,N_21309);
and U22321 (N_22321,N_21645,N_21668);
and U22322 (N_22322,N_21798,N_21695);
nand U22323 (N_22323,N_21357,N_21553);
nor U22324 (N_22324,N_21570,N_21763);
or U22325 (N_22325,N_21635,N_21951);
nor U22326 (N_22326,N_21173,N_21607);
nand U22327 (N_22327,N_21741,N_21821);
or U22328 (N_22328,N_21757,N_21106);
xnor U22329 (N_22329,N_21134,N_21672);
nand U22330 (N_22330,N_21489,N_21887);
and U22331 (N_22331,N_21546,N_21404);
xnor U22332 (N_22332,N_21886,N_21855);
or U22333 (N_22333,N_21150,N_21414);
or U22334 (N_22334,N_21110,N_21639);
nand U22335 (N_22335,N_21704,N_21811);
or U22336 (N_22336,N_21533,N_21966);
nor U22337 (N_22337,N_21729,N_21312);
or U22338 (N_22338,N_21258,N_21567);
xnor U22339 (N_22339,N_21958,N_21588);
and U22340 (N_22340,N_21128,N_21666);
xor U22341 (N_22341,N_21368,N_21848);
xor U22342 (N_22342,N_21275,N_21557);
nor U22343 (N_22343,N_21369,N_21813);
or U22344 (N_22344,N_21827,N_21664);
xnor U22345 (N_22345,N_21230,N_21071);
and U22346 (N_22346,N_21005,N_21670);
xnor U22347 (N_22347,N_21685,N_21076);
nor U22348 (N_22348,N_21970,N_21383);
nand U22349 (N_22349,N_21731,N_21207);
and U22350 (N_22350,N_21573,N_21995);
and U22351 (N_22351,N_21224,N_21654);
and U22352 (N_22352,N_21062,N_21922);
or U22353 (N_22353,N_21060,N_21376);
or U22354 (N_22354,N_21386,N_21665);
xnor U22355 (N_22355,N_21532,N_21241);
xnor U22356 (N_22356,N_21325,N_21417);
nand U22357 (N_22357,N_21107,N_21426);
nor U22358 (N_22358,N_21186,N_21818);
or U22359 (N_22359,N_21551,N_21184);
nor U22360 (N_22360,N_21105,N_21260);
or U22361 (N_22361,N_21579,N_21118);
nand U22362 (N_22362,N_21159,N_21632);
nand U22363 (N_22363,N_21717,N_21909);
and U22364 (N_22364,N_21936,N_21733);
nand U22365 (N_22365,N_21013,N_21467);
or U22366 (N_22366,N_21977,N_21085);
or U22367 (N_22367,N_21400,N_21826);
nand U22368 (N_22368,N_21724,N_21427);
xnor U22369 (N_22369,N_21067,N_21583);
or U22370 (N_22370,N_21644,N_21313);
xor U22371 (N_22371,N_21831,N_21382);
or U22372 (N_22372,N_21335,N_21943);
xnor U22373 (N_22373,N_21061,N_21558);
nand U22374 (N_22374,N_21608,N_21581);
nor U22375 (N_22375,N_21795,N_21277);
nand U22376 (N_22376,N_21023,N_21529);
nor U22377 (N_22377,N_21257,N_21387);
nor U22378 (N_22378,N_21834,N_21429);
nor U22379 (N_22379,N_21010,N_21683);
or U22380 (N_22380,N_21858,N_21019);
nor U22381 (N_22381,N_21272,N_21096);
and U22382 (N_22382,N_21516,N_21899);
nor U22383 (N_22383,N_21905,N_21199);
xor U22384 (N_22384,N_21540,N_21770);
xor U22385 (N_22385,N_21130,N_21126);
xnor U22386 (N_22386,N_21295,N_21206);
nand U22387 (N_22387,N_21284,N_21331);
xnor U22388 (N_22388,N_21208,N_21510);
or U22389 (N_22389,N_21955,N_21266);
or U22390 (N_22390,N_21407,N_21153);
xor U22391 (N_22391,N_21192,N_21526);
nand U22392 (N_22392,N_21874,N_21435);
nor U22393 (N_22393,N_21917,N_21663);
or U22394 (N_22394,N_21475,N_21355);
and U22395 (N_22395,N_21024,N_21782);
xnor U22396 (N_22396,N_21892,N_21618);
nand U22397 (N_22397,N_21315,N_21226);
xor U22398 (N_22398,N_21276,N_21079);
nor U22399 (N_22399,N_21506,N_21183);
nor U22400 (N_22400,N_21424,N_21611);
nor U22401 (N_22401,N_21572,N_21322);
and U22402 (N_22402,N_21536,N_21765);
nand U22403 (N_22403,N_21155,N_21373);
nor U22404 (N_22404,N_21692,N_21124);
nand U22405 (N_22405,N_21244,N_21838);
nor U22406 (N_22406,N_21769,N_21911);
nand U22407 (N_22407,N_21428,N_21777);
and U22408 (N_22408,N_21678,N_21726);
nand U22409 (N_22409,N_21193,N_21477);
xnor U22410 (N_22410,N_21871,N_21468);
nand U22411 (N_22411,N_21957,N_21637);
or U22412 (N_22412,N_21976,N_21565);
and U22413 (N_22413,N_21442,N_21293);
or U22414 (N_22414,N_21031,N_21687);
xor U22415 (N_22415,N_21701,N_21797);
and U22416 (N_22416,N_21863,N_21012);
nor U22417 (N_22417,N_21973,N_21179);
xnor U22418 (N_22418,N_21432,N_21924);
xnor U22419 (N_22419,N_21445,N_21398);
nor U22420 (N_22420,N_21392,N_21354);
nand U22421 (N_22421,N_21377,N_21590);
nand U22422 (N_22422,N_21721,N_21438);
nor U22423 (N_22423,N_21923,N_21908);
nand U22424 (N_22424,N_21103,N_21904);
or U22425 (N_22425,N_21045,N_21725);
nor U22426 (N_22426,N_21390,N_21318);
and U22427 (N_22427,N_21807,N_21402);
nor U22428 (N_22428,N_21336,N_21713);
nand U22429 (N_22429,N_21675,N_21245);
and U22430 (N_22430,N_21965,N_21825);
and U22431 (N_22431,N_21439,N_21388);
xnor U22432 (N_22432,N_21758,N_21554);
nor U22433 (N_22433,N_21162,N_21514);
and U22434 (N_22434,N_21485,N_21759);
nand U22435 (N_22435,N_21201,N_21235);
or U22436 (N_22436,N_21941,N_21723);
or U22437 (N_22437,N_21993,N_21679);
xnor U22438 (N_22438,N_21088,N_21087);
xor U22439 (N_22439,N_21136,N_21463);
nor U22440 (N_22440,N_21262,N_21751);
nand U22441 (N_22441,N_21983,N_21563);
and U22442 (N_22442,N_21584,N_21017);
or U22443 (N_22443,N_21507,N_21843);
nor U22444 (N_22444,N_21081,N_21926);
nand U22445 (N_22445,N_21730,N_21881);
nor U22446 (N_22446,N_21151,N_21727);
and U22447 (N_22447,N_21801,N_21994);
nand U22448 (N_22448,N_21430,N_21718);
xor U22449 (N_22449,N_21493,N_21981);
nand U22450 (N_22450,N_21203,N_21492);
and U22451 (N_22451,N_21742,N_21469);
nand U22452 (N_22452,N_21949,N_21847);
and U22453 (N_22453,N_21709,N_21706);
xor U22454 (N_22454,N_21247,N_21932);
or U22455 (N_22455,N_21025,N_21783);
nor U22456 (N_22456,N_21348,N_21090);
and U22457 (N_22457,N_21094,N_21168);
or U22458 (N_22458,N_21491,N_21408);
nor U22459 (N_22459,N_21421,N_21649);
and U22460 (N_22460,N_21156,N_21037);
xor U22461 (N_22461,N_21334,N_21669);
xnor U22462 (N_22462,N_21592,N_21779);
or U22463 (N_22463,N_21232,N_21185);
and U22464 (N_22464,N_21652,N_21114);
and U22465 (N_22465,N_21456,N_21389);
nor U22466 (N_22466,N_21634,N_21078);
and U22467 (N_22467,N_21457,N_21698);
nand U22468 (N_22468,N_21092,N_21189);
and U22469 (N_22469,N_21397,N_21378);
nand U22470 (N_22470,N_21937,N_21222);
and U22471 (N_22471,N_21747,N_21353);
nor U22472 (N_22472,N_21651,N_21656);
and U22473 (N_22473,N_21866,N_21913);
nand U22474 (N_22474,N_21714,N_21606);
or U22475 (N_22475,N_21767,N_21274);
or U22476 (N_22476,N_21236,N_21745);
and U22477 (N_22477,N_21835,N_21458);
nor U22478 (N_22478,N_21910,N_21470);
nand U22479 (N_22479,N_21629,N_21609);
or U22480 (N_22480,N_21534,N_21347);
nor U22481 (N_22481,N_21889,N_21403);
nand U22482 (N_22482,N_21753,N_21109);
and U22483 (N_22483,N_21317,N_21853);
nand U22484 (N_22484,N_21158,N_21410);
or U22485 (N_22485,N_21340,N_21550);
nand U22486 (N_22486,N_21283,N_21437);
nand U22487 (N_22487,N_21123,N_21875);
nor U22488 (N_22488,N_21867,N_21660);
nand U22489 (N_22489,N_21628,N_21950);
and U22490 (N_22490,N_21518,N_21175);
xnor U22491 (N_22491,N_21502,N_21131);
or U22492 (N_22492,N_21339,N_21381);
and U22493 (N_22493,N_21864,N_21152);
nor U22494 (N_22494,N_21614,N_21237);
or U22495 (N_22495,N_21627,N_21447);
nor U22496 (N_22496,N_21690,N_21015);
nand U22497 (N_22497,N_21111,N_21360);
and U22498 (N_22498,N_21413,N_21577);
or U22499 (N_22499,N_21289,N_21830);
nand U22500 (N_22500,N_21600,N_21862);
xnor U22501 (N_22501,N_21925,N_21466);
nand U22502 (N_22502,N_21034,N_21864);
or U22503 (N_22503,N_21893,N_21958);
and U22504 (N_22504,N_21639,N_21636);
xor U22505 (N_22505,N_21467,N_21441);
xnor U22506 (N_22506,N_21091,N_21736);
or U22507 (N_22507,N_21634,N_21053);
nand U22508 (N_22508,N_21468,N_21498);
xnor U22509 (N_22509,N_21856,N_21413);
xor U22510 (N_22510,N_21936,N_21432);
or U22511 (N_22511,N_21394,N_21717);
and U22512 (N_22512,N_21168,N_21350);
nor U22513 (N_22513,N_21264,N_21469);
and U22514 (N_22514,N_21515,N_21416);
and U22515 (N_22515,N_21502,N_21414);
nand U22516 (N_22516,N_21981,N_21204);
xor U22517 (N_22517,N_21683,N_21881);
and U22518 (N_22518,N_21937,N_21554);
nor U22519 (N_22519,N_21114,N_21956);
or U22520 (N_22520,N_21850,N_21834);
nand U22521 (N_22521,N_21387,N_21690);
xor U22522 (N_22522,N_21453,N_21240);
nand U22523 (N_22523,N_21082,N_21638);
and U22524 (N_22524,N_21858,N_21254);
or U22525 (N_22525,N_21569,N_21074);
and U22526 (N_22526,N_21123,N_21348);
xnor U22527 (N_22527,N_21270,N_21298);
or U22528 (N_22528,N_21390,N_21156);
nand U22529 (N_22529,N_21044,N_21692);
nand U22530 (N_22530,N_21931,N_21451);
xnor U22531 (N_22531,N_21017,N_21336);
nor U22532 (N_22532,N_21591,N_21790);
nor U22533 (N_22533,N_21919,N_21177);
nand U22534 (N_22534,N_21499,N_21138);
or U22535 (N_22535,N_21871,N_21362);
nand U22536 (N_22536,N_21456,N_21311);
nand U22537 (N_22537,N_21379,N_21250);
or U22538 (N_22538,N_21005,N_21449);
xnor U22539 (N_22539,N_21225,N_21460);
nand U22540 (N_22540,N_21956,N_21815);
or U22541 (N_22541,N_21359,N_21424);
xnor U22542 (N_22542,N_21120,N_21132);
nand U22543 (N_22543,N_21751,N_21523);
nand U22544 (N_22544,N_21082,N_21183);
nor U22545 (N_22545,N_21863,N_21130);
nor U22546 (N_22546,N_21813,N_21845);
or U22547 (N_22547,N_21978,N_21751);
nor U22548 (N_22548,N_21037,N_21761);
nand U22549 (N_22549,N_21960,N_21175);
or U22550 (N_22550,N_21512,N_21465);
and U22551 (N_22551,N_21738,N_21531);
and U22552 (N_22552,N_21920,N_21059);
xor U22553 (N_22553,N_21932,N_21299);
or U22554 (N_22554,N_21944,N_21010);
or U22555 (N_22555,N_21845,N_21653);
and U22556 (N_22556,N_21181,N_21504);
xnor U22557 (N_22557,N_21048,N_21281);
nand U22558 (N_22558,N_21630,N_21865);
nand U22559 (N_22559,N_21473,N_21537);
and U22560 (N_22560,N_21241,N_21037);
nand U22561 (N_22561,N_21121,N_21668);
or U22562 (N_22562,N_21204,N_21150);
nand U22563 (N_22563,N_21111,N_21131);
and U22564 (N_22564,N_21850,N_21749);
nand U22565 (N_22565,N_21502,N_21739);
nand U22566 (N_22566,N_21760,N_21647);
or U22567 (N_22567,N_21710,N_21055);
nand U22568 (N_22568,N_21348,N_21739);
nand U22569 (N_22569,N_21186,N_21808);
nor U22570 (N_22570,N_21908,N_21678);
xnor U22571 (N_22571,N_21844,N_21432);
nand U22572 (N_22572,N_21348,N_21487);
xnor U22573 (N_22573,N_21180,N_21643);
nor U22574 (N_22574,N_21262,N_21733);
nand U22575 (N_22575,N_21429,N_21274);
and U22576 (N_22576,N_21893,N_21435);
and U22577 (N_22577,N_21914,N_21286);
nand U22578 (N_22578,N_21561,N_21489);
or U22579 (N_22579,N_21486,N_21163);
and U22580 (N_22580,N_21564,N_21139);
or U22581 (N_22581,N_21525,N_21460);
and U22582 (N_22582,N_21161,N_21512);
or U22583 (N_22583,N_21151,N_21112);
or U22584 (N_22584,N_21509,N_21445);
or U22585 (N_22585,N_21001,N_21266);
nor U22586 (N_22586,N_21483,N_21295);
nor U22587 (N_22587,N_21457,N_21245);
xnor U22588 (N_22588,N_21927,N_21078);
or U22589 (N_22589,N_21538,N_21341);
xnor U22590 (N_22590,N_21832,N_21481);
or U22591 (N_22591,N_21617,N_21262);
or U22592 (N_22592,N_21006,N_21179);
or U22593 (N_22593,N_21815,N_21270);
xor U22594 (N_22594,N_21417,N_21092);
nor U22595 (N_22595,N_21315,N_21673);
nand U22596 (N_22596,N_21504,N_21609);
nor U22597 (N_22597,N_21874,N_21886);
nand U22598 (N_22598,N_21549,N_21905);
and U22599 (N_22599,N_21026,N_21668);
and U22600 (N_22600,N_21648,N_21440);
or U22601 (N_22601,N_21265,N_21031);
and U22602 (N_22602,N_21602,N_21915);
xnor U22603 (N_22603,N_21399,N_21366);
nand U22604 (N_22604,N_21307,N_21872);
and U22605 (N_22605,N_21191,N_21154);
and U22606 (N_22606,N_21406,N_21107);
nor U22607 (N_22607,N_21154,N_21933);
nor U22608 (N_22608,N_21672,N_21754);
or U22609 (N_22609,N_21505,N_21346);
nor U22610 (N_22610,N_21531,N_21576);
nor U22611 (N_22611,N_21812,N_21480);
xor U22612 (N_22612,N_21823,N_21211);
and U22613 (N_22613,N_21153,N_21251);
nor U22614 (N_22614,N_21094,N_21086);
and U22615 (N_22615,N_21762,N_21509);
and U22616 (N_22616,N_21530,N_21478);
xor U22617 (N_22617,N_21384,N_21308);
or U22618 (N_22618,N_21703,N_21760);
xnor U22619 (N_22619,N_21295,N_21546);
nor U22620 (N_22620,N_21098,N_21237);
xor U22621 (N_22621,N_21568,N_21850);
nand U22622 (N_22622,N_21821,N_21183);
xor U22623 (N_22623,N_21145,N_21403);
nand U22624 (N_22624,N_21503,N_21933);
nor U22625 (N_22625,N_21803,N_21992);
xnor U22626 (N_22626,N_21933,N_21390);
or U22627 (N_22627,N_21553,N_21607);
and U22628 (N_22628,N_21480,N_21210);
and U22629 (N_22629,N_21769,N_21611);
or U22630 (N_22630,N_21139,N_21752);
nor U22631 (N_22631,N_21845,N_21523);
or U22632 (N_22632,N_21250,N_21577);
or U22633 (N_22633,N_21860,N_21055);
nand U22634 (N_22634,N_21360,N_21270);
nand U22635 (N_22635,N_21219,N_21652);
or U22636 (N_22636,N_21710,N_21226);
and U22637 (N_22637,N_21197,N_21518);
xnor U22638 (N_22638,N_21792,N_21013);
xnor U22639 (N_22639,N_21538,N_21990);
nand U22640 (N_22640,N_21324,N_21927);
or U22641 (N_22641,N_21525,N_21975);
xor U22642 (N_22642,N_21010,N_21221);
nand U22643 (N_22643,N_21488,N_21998);
nand U22644 (N_22644,N_21838,N_21787);
nand U22645 (N_22645,N_21663,N_21522);
xnor U22646 (N_22646,N_21509,N_21488);
xnor U22647 (N_22647,N_21947,N_21401);
or U22648 (N_22648,N_21481,N_21976);
and U22649 (N_22649,N_21430,N_21572);
and U22650 (N_22650,N_21053,N_21533);
nand U22651 (N_22651,N_21433,N_21120);
nor U22652 (N_22652,N_21260,N_21344);
and U22653 (N_22653,N_21777,N_21961);
nand U22654 (N_22654,N_21756,N_21285);
and U22655 (N_22655,N_21937,N_21969);
and U22656 (N_22656,N_21804,N_21300);
nor U22657 (N_22657,N_21317,N_21040);
xnor U22658 (N_22658,N_21875,N_21087);
and U22659 (N_22659,N_21469,N_21554);
and U22660 (N_22660,N_21304,N_21438);
or U22661 (N_22661,N_21589,N_21940);
nand U22662 (N_22662,N_21890,N_21862);
xnor U22663 (N_22663,N_21000,N_21988);
and U22664 (N_22664,N_21744,N_21515);
and U22665 (N_22665,N_21936,N_21483);
and U22666 (N_22666,N_21703,N_21649);
and U22667 (N_22667,N_21921,N_21956);
or U22668 (N_22668,N_21160,N_21648);
nor U22669 (N_22669,N_21874,N_21881);
nor U22670 (N_22670,N_21884,N_21174);
nand U22671 (N_22671,N_21060,N_21898);
xnor U22672 (N_22672,N_21265,N_21870);
xor U22673 (N_22673,N_21286,N_21466);
nand U22674 (N_22674,N_21822,N_21643);
xor U22675 (N_22675,N_21296,N_21530);
and U22676 (N_22676,N_21012,N_21339);
xnor U22677 (N_22677,N_21900,N_21629);
and U22678 (N_22678,N_21161,N_21118);
nor U22679 (N_22679,N_21452,N_21388);
xnor U22680 (N_22680,N_21298,N_21496);
xor U22681 (N_22681,N_21995,N_21074);
nand U22682 (N_22682,N_21019,N_21260);
xor U22683 (N_22683,N_21547,N_21813);
xor U22684 (N_22684,N_21738,N_21764);
and U22685 (N_22685,N_21727,N_21291);
nor U22686 (N_22686,N_21301,N_21830);
and U22687 (N_22687,N_21965,N_21500);
nor U22688 (N_22688,N_21280,N_21396);
nor U22689 (N_22689,N_21685,N_21915);
or U22690 (N_22690,N_21924,N_21875);
and U22691 (N_22691,N_21950,N_21425);
nor U22692 (N_22692,N_21629,N_21551);
nand U22693 (N_22693,N_21918,N_21789);
nor U22694 (N_22694,N_21836,N_21148);
xnor U22695 (N_22695,N_21381,N_21829);
or U22696 (N_22696,N_21022,N_21497);
nor U22697 (N_22697,N_21715,N_21533);
nor U22698 (N_22698,N_21063,N_21738);
nor U22699 (N_22699,N_21734,N_21118);
nand U22700 (N_22700,N_21430,N_21840);
nor U22701 (N_22701,N_21824,N_21543);
nor U22702 (N_22702,N_21119,N_21456);
nor U22703 (N_22703,N_21071,N_21944);
nor U22704 (N_22704,N_21929,N_21158);
xnor U22705 (N_22705,N_21018,N_21063);
and U22706 (N_22706,N_21520,N_21496);
xor U22707 (N_22707,N_21320,N_21859);
or U22708 (N_22708,N_21707,N_21886);
xnor U22709 (N_22709,N_21064,N_21192);
and U22710 (N_22710,N_21785,N_21411);
nand U22711 (N_22711,N_21602,N_21585);
nor U22712 (N_22712,N_21870,N_21030);
and U22713 (N_22713,N_21548,N_21052);
nor U22714 (N_22714,N_21255,N_21031);
or U22715 (N_22715,N_21202,N_21600);
xnor U22716 (N_22716,N_21223,N_21075);
nand U22717 (N_22717,N_21112,N_21984);
and U22718 (N_22718,N_21563,N_21691);
or U22719 (N_22719,N_21164,N_21709);
or U22720 (N_22720,N_21304,N_21809);
or U22721 (N_22721,N_21475,N_21654);
nor U22722 (N_22722,N_21818,N_21083);
xor U22723 (N_22723,N_21823,N_21557);
and U22724 (N_22724,N_21355,N_21018);
nor U22725 (N_22725,N_21740,N_21862);
nor U22726 (N_22726,N_21189,N_21728);
xnor U22727 (N_22727,N_21219,N_21978);
and U22728 (N_22728,N_21523,N_21317);
xor U22729 (N_22729,N_21595,N_21946);
nor U22730 (N_22730,N_21438,N_21774);
xnor U22731 (N_22731,N_21749,N_21760);
or U22732 (N_22732,N_21025,N_21175);
nand U22733 (N_22733,N_21552,N_21631);
or U22734 (N_22734,N_21435,N_21896);
and U22735 (N_22735,N_21660,N_21215);
xor U22736 (N_22736,N_21712,N_21365);
nor U22737 (N_22737,N_21391,N_21547);
xnor U22738 (N_22738,N_21311,N_21407);
and U22739 (N_22739,N_21983,N_21603);
nand U22740 (N_22740,N_21466,N_21855);
and U22741 (N_22741,N_21000,N_21637);
or U22742 (N_22742,N_21536,N_21106);
nor U22743 (N_22743,N_21207,N_21468);
nand U22744 (N_22744,N_21121,N_21267);
xnor U22745 (N_22745,N_21900,N_21199);
nand U22746 (N_22746,N_21921,N_21079);
or U22747 (N_22747,N_21622,N_21216);
nand U22748 (N_22748,N_21389,N_21573);
xnor U22749 (N_22749,N_21510,N_21728);
nand U22750 (N_22750,N_21538,N_21607);
xnor U22751 (N_22751,N_21885,N_21113);
xnor U22752 (N_22752,N_21335,N_21193);
and U22753 (N_22753,N_21069,N_21131);
and U22754 (N_22754,N_21322,N_21919);
nor U22755 (N_22755,N_21158,N_21213);
or U22756 (N_22756,N_21647,N_21155);
nand U22757 (N_22757,N_21079,N_21536);
nor U22758 (N_22758,N_21714,N_21567);
or U22759 (N_22759,N_21862,N_21629);
or U22760 (N_22760,N_21525,N_21712);
xnor U22761 (N_22761,N_21849,N_21485);
nor U22762 (N_22762,N_21761,N_21470);
nand U22763 (N_22763,N_21123,N_21839);
and U22764 (N_22764,N_21577,N_21791);
and U22765 (N_22765,N_21822,N_21349);
and U22766 (N_22766,N_21932,N_21126);
and U22767 (N_22767,N_21220,N_21854);
and U22768 (N_22768,N_21222,N_21243);
nor U22769 (N_22769,N_21584,N_21116);
xor U22770 (N_22770,N_21691,N_21900);
nand U22771 (N_22771,N_21943,N_21003);
or U22772 (N_22772,N_21242,N_21090);
and U22773 (N_22773,N_21963,N_21347);
xnor U22774 (N_22774,N_21752,N_21636);
and U22775 (N_22775,N_21689,N_21404);
nand U22776 (N_22776,N_21735,N_21599);
or U22777 (N_22777,N_21383,N_21976);
nor U22778 (N_22778,N_21920,N_21184);
xor U22779 (N_22779,N_21250,N_21225);
nor U22780 (N_22780,N_21017,N_21066);
and U22781 (N_22781,N_21482,N_21351);
and U22782 (N_22782,N_21784,N_21616);
or U22783 (N_22783,N_21748,N_21093);
or U22784 (N_22784,N_21253,N_21475);
and U22785 (N_22785,N_21225,N_21493);
nand U22786 (N_22786,N_21506,N_21970);
xnor U22787 (N_22787,N_21556,N_21069);
and U22788 (N_22788,N_21744,N_21022);
or U22789 (N_22789,N_21525,N_21170);
and U22790 (N_22790,N_21229,N_21582);
nand U22791 (N_22791,N_21199,N_21479);
nor U22792 (N_22792,N_21746,N_21504);
and U22793 (N_22793,N_21224,N_21856);
xor U22794 (N_22794,N_21635,N_21174);
nand U22795 (N_22795,N_21556,N_21255);
nand U22796 (N_22796,N_21391,N_21530);
nand U22797 (N_22797,N_21346,N_21784);
or U22798 (N_22798,N_21080,N_21177);
nor U22799 (N_22799,N_21972,N_21031);
and U22800 (N_22800,N_21947,N_21734);
or U22801 (N_22801,N_21700,N_21458);
or U22802 (N_22802,N_21076,N_21058);
and U22803 (N_22803,N_21772,N_21092);
and U22804 (N_22804,N_21346,N_21181);
xor U22805 (N_22805,N_21281,N_21659);
and U22806 (N_22806,N_21361,N_21993);
xnor U22807 (N_22807,N_21206,N_21495);
xnor U22808 (N_22808,N_21746,N_21563);
nor U22809 (N_22809,N_21655,N_21923);
nand U22810 (N_22810,N_21165,N_21972);
xnor U22811 (N_22811,N_21776,N_21494);
nor U22812 (N_22812,N_21194,N_21918);
and U22813 (N_22813,N_21249,N_21676);
and U22814 (N_22814,N_21526,N_21985);
xor U22815 (N_22815,N_21791,N_21985);
nor U22816 (N_22816,N_21153,N_21511);
nor U22817 (N_22817,N_21451,N_21930);
nor U22818 (N_22818,N_21337,N_21738);
xnor U22819 (N_22819,N_21668,N_21159);
xnor U22820 (N_22820,N_21746,N_21938);
xor U22821 (N_22821,N_21990,N_21460);
or U22822 (N_22822,N_21229,N_21496);
xor U22823 (N_22823,N_21445,N_21470);
nand U22824 (N_22824,N_21688,N_21402);
and U22825 (N_22825,N_21638,N_21972);
nor U22826 (N_22826,N_21102,N_21223);
or U22827 (N_22827,N_21399,N_21675);
xnor U22828 (N_22828,N_21923,N_21631);
nand U22829 (N_22829,N_21808,N_21636);
xnor U22830 (N_22830,N_21134,N_21329);
nand U22831 (N_22831,N_21565,N_21581);
xor U22832 (N_22832,N_21711,N_21985);
xor U22833 (N_22833,N_21115,N_21496);
nor U22834 (N_22834,N_21156,N_21102);
xor U22835 (N_22835,N_21346,N_21007);
and U22836 (N_22836,N_21770,N_21027);
xnor U22837 (N_22837,N_21052,N_21725);
nor U22838 (N_22838,N_21829,N_21185);
xor U22839 (N_22839,N_21218,N_21824);
nor U22840 (N_22840,N_21581,N_21661);
and U22841 (N_22841,N_21458,N_21931);
xor U22842 (N_22842,N_21477,N_21026);
nand U22843 (N_22843,N_21560,N_21899);
and U22844 (N_22844,N_21297,N_21207);
nor U22845 (N_22845,N_21128,N_21113);
xnor U22846 (N_22846,N_21856,N_21479);
nand U22847 (N_22847,N_21174,N_21891);
nor U22848 (N_22848,N_21206,N_21706);
xnor U22849 (N_22849,N_21066,N_21250);
nand U22850 (N_22850,N_21622,N_21751);
or U22851 (N_22851,N_21859,N_21341);
nor U22852 (N_22852,N_21962,N_21225);
or U22853 (N_22853,N_21281,N_21720);
nor U22854 (N_22854,N_21916,N_21276);
xor U22855 (N_22855,N_21561,N_21590);
nor U22856 (N_22856,N_21356,N_21017);
xor U22857 (N_22857,N_21373,N_21142);
or U22858 (N_22858,N_21101,N_21450);
xnor U22859 (N_22859,N_21552,N_21788);
nand U22860 (N_22860,N_21594,N_21729);
nor U22861 (N_22861,N_21642,N_21436);
or U22862 (N_22862,N_21254,N_21348);
nor U22863 (N_22863,N_21164,N_21065);
xor U22864 (N_22864,N_21916,N_21561);
nor U22865 (N_22865,N_21191,N_21441);
xor U22866 (N_22866,N_21296,N_21852);
and U22867 (N_22867,N_21195,N_21096);
and U22868 (N_22868,N_21886,N_21438);
or U22869 (N_22869,N_21924,N_21520);
nand U22870 (N_22870,N_21169,N_21408);
xor U22871 (N_22871,N_21890,N_21717);
xor U22872 (N_22872,N_21623,N_21974);
nor U22873 (N_22873,N_21358,N_21415);
and U22874 (N_22874,N_21787,N_21661);
nor U22875 (N_22875,N_21116,N_21403);
or U22876 (N_22876,N_21572,N_21816);
and U22877 (N_22877,N_21498,N_21616);
or U22878 (N_22878,N_21953,N_21525);
or U22879 (N_22879,N_21922,N_21705);
or U22880 (N_22880,N_21327,N_21932);
and U22881 (N_22881,N_21699,N_21914);
xnor U22882 (N_22882,N_21810,N_21872);
xnor U22883 (N_22883,N_21379,N_21903);
nand U22884 (N_22884,N_21505,N_21550);
and U22885 (N_22885,N_21822,N_21534);
and U22886 (N_22886,N_21182,N_21129);
nor U22887 (N_22887,N_21885,N_21689);
or U22888 (N_22888,N_21700,N_21461);
nor U22889 (N_22889,N_21887,N_21378);
nor U22890 (N_22890,N_21971,N_21333);
and U22891 (N_22891,N_21853,N_21765);
nand U22892 (N_22892,N_21096,N_21897);
or U22893 (N_22893,N_21438,N_21454);
and U22894 (N_22894,N_21112,N_21166);
nand U22895 (N_22895,N_21369,N_21754);
or U22896 (N_22896,N_21691,N_21599);
or U22897 (N_22897,N_21541,N_21686);
or U22898 (N_22898,N_21047,N_21756);
xnor U22899 (N_22899,N_21560,N_21533);
xnor U22900 (N_22900,N_21582,N_21811);
xor U22901 (N_22901,N_21695,N_21725);
and U22902 (N_22902,N_21839,N_21735);
nor U22903 (N_22903,N_21456,N_21435);
or U22904 (N_22904,N_21463,N_21007);
and U22905 (N_22905,N_21620,N_21148);
and U22906 (N_22906,N_21859,N_21843);
nand U22907 (N_22907,N_21656,N_21772);
nand U22908 (N_22908,N_21077,N_21334);
nor U22909 (N_22909,N_21669,N_21788);
nand U22910 (N_22910,N_21371,N_21288);
and U22911 (N_22911,N_21531,N_21571);
or U22912 (N_22912,N_21269,N_21844);
nand U22913 (N_22913,N_21898,N_21145);
and U22914 (N_22914,N_21892,N_21259);
nor U22915 (N_22915,N_21528,N_21743);
xnor U22916 (N_22916,N_21707,N_21148);
xor U22917 (N_22917,N_21183,N_21924);
nor U22918 (N_22918,N_21400,N_21762);
xnor U22919 (N_22919,N_21971,N_21120);
or U22920 (N_22920,N_21110,N_21280);
nand U22921 (N_22921,N_21804,N_21380);
and U22922 (N_22922,N_21609,N_21998);
xnor U22923 (N_22923,N_21466,N_21803);
nand U22924 (N_22924,N_21225,N_21973);
nor U22925 (N_22925,N_21899,N_21472);
xnor U22926 (N_22926,N_21716,N_21192);
or U22927 (N_22927,N_21835,N_21151);
and U22928 (N_22928,N_21966,N_21099);
xor U22929 (N_22929,N_21348,N_21396);
nand U22930 (N_22930,N_21959,N_21648);
or U22931 (N_22931,N_21405,N_21383);
and U22932 (N_22932,N_21178,N_21138);
nor U22933 (N_22933,N_21497,N_21304);
and U22934 (N_22934,N_21394,N_21737);
xnor U22935 (N_22935,N_21540,N_21302);
nand U22936 (N_22936,N_21388,N_21525);
or U22937 (N_22937,N_21545,N_21963);
and U22938 (N_22938,N_21119,N_21235);
and U22939 (N_22939,N_21868,N_21959);
nor U22940 (N_22940,N_21058,N_21501);
xor U22941 (N_22941,N_21743,N_21476);
and U22942 (N_22942,N_21898,N_21759);
nand U22943 (N_22943,N_21881,N_21939);
xnor U22944 (N_22944,N_21381,N_21360);
xor U22945 (N_22945,N_21211,N_21331);
nand U22946 (N_22946,N_21253,N_21768);
or U22947 (N_22947,N_21857,N_21449);
xnor U22948 (N_22948,N_21237,N_21231);
nand U22949 (N_22949,N_21455,N_21013);
and U22950 (N_22950,N_21316,N_21737);
and U22951 (N_22951,N_21390,N_21373);
nand U22952 (N_22952,N_21865,N_21493);
and U22953 (N_22953,N_21625,N_21589);
and U22954 (N_22954,N_21803,N_21501);
and U22955 (N_22955,N_21705,N_21486);
xor U22956 (N_22956,N_21991,N_21574);
and U22957 (N_22957,N_21937,N_21702);
nand U22958 (N_22958,N_21676,N_21957);
xor U22959 (N_22959,N_21954,N_21691);
nand U22960 (N_22960,N_21661,N_21297);
nor U22961 (N_22961,N_21194,N_21137);
nand U22962 (N_22962,N_21421,N_21209);
nor U22963 (N_22963,N_21582,N_21100);
and U22964 (N_22964,N_21060,N_21439);
xor U22965 (N_22965,N_21768,N_21908);
or U22966 (N_22966,N_21385,N_21784);
and U22967 (N_22967,N_21867,N_21360);
nand U22968 (N_22968,N_21332,N_21284);
and U22969 (N_22969,N_21314,N_21239);
xnor U22970 (N_22970,N_21514,N_21297);
or U22971 (N_22971,N_21039,N_21959);
nand U22972 (N_22972,N_21144,N_21106);
and U22973 (N_22973,N_21569,N_21541);
nor U22974 (N_22974,N_21502,N_21456);
and U22975 (N_22975,N_21967,N_21230);
or U22976 (N_22976,N_21970,N_21823);
xor U22977 (N_22977,N_21990,N_21195);
nor U22978 (N_22978,N_21052,N_21159);
or U22979 (N_22979,N_21235,N_21178);
nand U22980 (N_22980,N_21299,N_21930);
xnor U22981 (N_22981,N_21471,N_21814);
or U22982 (N_22982,N_21203,N_21765);
nor U22983 (N_22983,N_21578,N_21131);
and U22984 (N_22984,N_21627,N_21688);
nor U22985 (N_22985,N_21883,N_21985);
nand U22986 (N_22986,N_21802,N_21858);
nand U22987 (N_22987,N_21071,N_21836);
xnor U22988 (N_22988,N_21871,N_21397);
xor U22989 (N_22989,N_21067,N_21267);
nand U22990 (N_22990,N_21035,N_21718);
nor U22991 (N_22991,N_21636,N_21115);
nand U22992 (N_22992,N_21489,N_21420);
xnor U22993 (N_22993,N_21274,N_21509);
xor U22994 (N_22994,N_21351,N_21025);
xnor U22995 (N_22995,N_21921,N_21787);
and U22996 (N_22996,N_21434,N_21688);
or U22997 (N_22997,N_21922,N_21985);
nand U22998 (N_22998,N_21828,N_21878);
or U22999 (N_22999,N_21879,N_21683);
or U23000 (N_23000,N_22151,N_22582);
xor U23001 (N_23001,N_22036,N_22828);
or U23002 (N_23002,N_22784,N_22860);
nand U23003 (N_23003,N_22906,N_22969);
nand U23004 (N_23004,N_22685,N_22696);
or U23005 (N_23005,N_22429,N_22074);
nor U23006 (N_23006,N_22686,N_22426);
nand U23007 (N_23007,N_22076,N_22260);
nand U23008 (N_23008,N_22902,N_22681);
nor U23009 (N_23009,N_22812,N_22659);
nand U23010 (N_23010,N_22952,N_22556);
and U23011 (N_23011,N_22214,N_22626);
nor U23012 (N_23012,N_22719,N_22810);
xor U23013 (N_23013,N_22738,N_22264);
and U23014 (N_23014,N_22372,N_22829);
nor U23015 (N_23015,N_22342,N_22639);
nor U23016 (N_23016,N_22033,N_22647);
or U23017 (N_23017,N_22682,N_22565);
nand U23018 (N_23018,N_22588,N_22974);
or U23019 (N_23019,N_22722,N_22936);
nor U23020 (N_23020,N_22535,N_22634);
xnor U23021 (N_23021,N_22825,N_22038);
nor U23022 (N_23022,N_22774,N_22017);
xor U23023 (N_23023,N_22912,N_22631);
nor U23024 (N_23024,N_22942,N_22472);
or U23025 (N_23025,N_22951,N_22893);
and U23026 (N_23026,N_22619,N_22311);
nor U23027 (N_23027,N_22579,N_22813);
xnor U23028 (N_23028,N_22628,N_22736);
or U23029 (N_23029,N_22744,N_22019);
xor U23030 (N_23030,N_22028,N_22894);
or U23031 (N_23031,N_22760,N_22694);
or U23032 (N_23032,N_22529,N_22649);
and U23033 (N_23033,N_22559,N_22864);
and U23034 (N_23034,N_22504,N_22469);
and U23035 (N_23035,N_22710,N_22403);
and U23036 (N_23036,N_22612,N_22586);
and U23037 (N_23037,N_22416,N_22175);
and U23038 (N_23038,N_22616,N_22240);
xor U23039 (N_23039,N_22709,N_22259);
nor U23040 (N_23040,N_22961,N_22419);
or U23041 (N_23041,N_22176,N_22415);
or U23042 (N_23042,N_22518,N_22883);
nand U23043 (N_23043,N_22304,N_22247);
nand U23044 (N_23044,N_22560,N_22135);
xnor U23045 (N_23045,N_22862,N_22528);
xnor U23046 (N_23046,N_22370,N_22935);
nand U23047 (N_23047,N_22910,N_22023);
nor U23048 (N_23048,N_22436,N_22932);
xor U23049 (N_23049,N_22439,N_22119);
nand U23050 (N_23050,N_22078,N_22000);
nand U23051 (N_23051,N_22684,N_22997);
nand U23052 (N_23052,N_22059,N_22716);
and U23053 (N_23053,N_22369,N_22352);
or U23054 (N_23054,N_22447,N_22377);
nand U23055 (N_23055,N_22053,N_22088);
xnor U23056 (N_23056,N_22795,N_22975);
or U23057 (N_23057,N_22152,N_22930);
xnor U23058 (N_23058,N_22082,N_22394);
nor U23059 (N_23059,N_22671,N_22618);
nand U23060 (N_23060,N_22237,N_22479);
nor U23061 (N_23061,N_22102,N_22536);
xor U23062 (N_23062,N_22547,N_22968);
or U23063 (N_23063,N_22374,N_22139);
nor U23064 (N_23064,N_22690,N_22021);
xnor U23065 (N_23065,N_22454,N_22723);
nand U23066 (N_23066,N_22324,N_22672);
xor U23067 (N_23067,N_22727,N_22406);
or U23068 (N_23068,N_22138,N_22923);
nor U23069 (N_23069,N_22087,N_22045);
nor U23070 (N_23070,N_22830,N_22758);
xor U23071 (N_23071,N_22804,N_22858);
and U23072 (N_23072,N_22113,N_22850);
or U23073 (N_23073,N_22411,N_22363);
nor U23074 (N_23074,N_22283,N_22305);
and U23075 (N_23075,N_22978,N_22458);
nand U23076 (N_23076,N_22487,N_22446);
xnor U23077 (N_23077,N_22897,N_22115);
nor U23078 (N_23078,N_22590,N_22869);
nor U23079 (N_23079,N_22180,N_22674);
and U23080 (N_23080,N_22382,N_22186);
and U23081 (N_23081,N_22605,N_22246);
or U23082 (N_23082,N_22269,N_22707);
nor U23083 (N_23083,N_22482,N_22293);
nor U23084 (N_23084,N_22179,N_22800);
or U23085 (N_23085,N_22958,N_22622);
and U23086 (N_23086,N_22405,N_22357);
or U23087 (N_23087,N_22770,N_22717);
or U23088 (N_23088,N_22281,N_22356);
xnor U23089 (N_23089,N_22809,N_22903);
nand U23090 (N_23090,N_22383,N_22300);
nand U23091 (N_23091,N_22623,N_22303);
nor U23092 (N_23092,N_22703,N_22235);
nand U23093 (N_23093,N_22753,N_22699);
and U23094 (N_23094,N_22348,N_22194);
nand U23095 (N_23095,N_22483,N_22270);
and U23096 (N_23096,N_22614,N_22927);
xnor U23097 (N_23097,N_22325,N_22276);
or U23098 (N_23098,N_22944,N_22554);
or U23099 (N_23099,N_22286,N_22987);
or U23100 (N_23100,N_22338,N_22872);
nand U23101 (N_23101,N_22852,N_22039);
nor U23102 (N_23102,N_22851,N_22277);
xnor U23103 (N_23103,N_22054,N_22089);
and U23104 (N_23104,N_22667,N_22938);
and U23105 (N_23105,N_22972,N_22947);
xor U23106 (N_23106,N_22513,N_22787);
and U23107 (N_23107,N_22500,N_22531);
nor U23108 (N_23108,N_22189,N_22721);
nand U23109 (N_23109,N_22937,N_22421);
or U23110 (N_23110,N_22607,N_22391);
or U23111 (N_23111,N_22549,N_22174);
nand U23112 (N_23112,N_22470,N_22637);
and U23113 (N_23113,N_22512,N_22929);
nor U23114 (N_23114,N_22498,N_22648);
and U23115 (N_23115,N_22256,N_22199);
nor U23116 (N_23116,N_22025,N_22700);
xnor U23117 (N_23117,N_22066,N_22558);
or U23118 (N_23118,N_22012,N_22859);
or U23119 (N_23119,N_22577,N_22833);
nor U23120 (N_23120,N_22640,N_22835);
or U23121 (N_23121,N_22677,N_22125);
or U23122 (N_23122,N_22735,N_22473);
or U23123 (N_23123,N_22546,N_22654);
or U23124 (N_23124,N_22344,N_22629);
nor U23125 (N_23125,N_22730,N_22386);
nand U23126 (N_23126,N_22678,N_22171);
and U23127 (N_23127,N_22056,N_22704);
xnor U23128 (N_23128,N_22361,N_22123);
xnor U23129 (N_23129,N_22339,N_22250);
and U23130 (N_23130,N_22853,N_22495);
xor U23131 (N_23131,N_22491,N_22211);
and U23132 (N_23132,N_22408,N_22219);
nand U23133 (N_23133,N_22816,N_22514);
nand U23134 (N_23134,N_22266,N_22210);
nor U23135 (N_23135,N_22899,N_22541);
nand U23136 (N_23136,N_22392,N_22687);
nor U23137 (N_23137,N_22578,N_22192);
xnor U23138 (N_23138,N_22802,N_22380);
and U23139 (N_23139,N_22085,N_22551);
xor U23140 (N_23140,N_22731,N_22844);
xor U23141 (N_23141,N_22279,N_22014);
nor U23142 (N_23142,N_22561,N_22569);
or U23143 (N_23143,N_22042,N_22061);
nand U23144 (N_23144,N_22073,N_22966);
xor U23145 (N_23145,N_22327,N_22353);
nand U23146 (N_23146,N_22335,N_22763);
nand U23147 (N_23147,N_22794,N_22101);
xnor U23148 (N_23148,N_22431,N_22792);
nand U23149 (N_23149,N_22530,N_22395);
xor U23150 (N_23150,N_22861,N_22052);
or U23151 (N_23151,N_22777,N_22563);
or U23152 (N_23152,N_22432,N_22093);
nor U23153 (N_23153,N_22414,N_22789);
nand U23154 (N_23154,N_22609,N_22440);
or U23155 (N_23155,N_22463,N_22740);
nand U23156 (N_23156,N_22100,N_22438);
xor U23157 (N_23157,N_22627,N_22516);
xnor U23158 (N_23158,N_22575,N_22956);
nor U23159 (N_23159,N_22092,N_22567);
nand U23160 (N_23160,N_22752,N_22769);
nor U23161 (N_23161,N_22583,N_22287);
nor U23162 (N_23162,N_22332,N_22520);
nor U23163 (N_23163,N_22739,N_22691);
or U23164 (N_23164,N_22594,N_22302);
nor U23165 (N_23165,N_22477,N_22030);
nor U23166 (N_23166,N_22288,N_22815);
nand U23167 (N_23167,N_22116,N_22570);
and U23168 (N_23168,N_22350,N_22244);
or U23169 (N_23169,N_22765,N_22867);
or U23170 (N_23170,N_22708,N_22026);
nor U23171 (N_23171,N_22697,N_22824);
nor U23172 (N_23172,N_22226,N_22959);
xnor U23173 (N_23173,N_22946,N_22320);
nand U23174 (N_23174,N_22509,N_22013);
or U23175 (N_23175,N_22020,N_22613);
or U23176 (N_23176,N_22257,N_22163);
nand U23177 (N_23177,N_22878,N_22148);
or U23178 (N_23178,N_22010,N_22705);
or U23179 (N_23179,N_22114,N_22295);
or U23180 (N_23180,N_22775,N_22451);
or U23181 (N_23181,N_22349,N_22538);
or U23182 (N_23182,N_22204,N_22050);
nor U23183 (N_23183,N_22232,N_22404);
or U23184 (N_23184,N_22786,N_22423);
xor U23185 (N_23185,N_22328,N_22918);
nand U23186 (N_23186,N_22664,N_22086);
or U23187 (N_23187,N_22358,N_22006);
xor U23188 (N_23188,N_22109,N_22355);
nand U23189 (N_23189,N_22949,N_22243);
and U23190 (N_23190,N_22007,N_22212);
xor U23191 (N_23191,N_22838,N_22268);
and U23192 (N_23192,N_22166,N_22132);
or U23193 (N_23193,N_22203,N_22315);
nor U23194 (N_23194,N_22106,N_22475);
or U23195 (N_23195,N_22149,N_22943);
xnor U23196 (N_23196,N_22826,N_22728);
or U23197 (N_23197,N_22761,N_22022);
or U23198 (N_23198,N_22955,N_22371);
or U23199 (N_23199,N_22772,N_22322);
or U23200 (N_23200,N_22108,N_22510);
or U23201 (N_23201,N_22720,N_22112);
and U23202 (N_23202,N_22005,N_22611);
or U23203 (N_23203,N_22091,N_22597);
or U23204 (N_23204,N_22187,N_22016);
xnor U23205 (N_23205,N_22190,N_22759);
nand U23206 (N_23206,N_22522,N_22928);
nand U23207 (N_23207,N_22865,N_22982);
nor U23208 (N_23208,N_22988,N_22953);
and U23209 (N_23209,N_22048,N_22027);
and U23210 (N_23210,N_22107,N_22499);
nand U23211 (N_23211,N_22445,N_22553);
or U23212 (N_23212,N_22562,N_22688);
xor U23213 (N_23213,N_22231,N_22127);
xnor U23214 (N_23214,N_22548,N_22990);
xor U23215 (N_23215,N_22907,N_22989);
or U23216 (N_23216,N_22400,N_22651);
nand U23217 (N_23217,N_22837,N_22275);
and U23218 (N_23218,N_22433,N_22417);
nor U23219 (N_23219,N_22222,N_22343);
xnor U23220 (N_23220,N_22347,N_22185);
or U23221 (N_23221,N_22849,N_22539);
nand U23222 (N_23222,N_22455,N_22037);
nor U23223 (N_23223,N_22873,N_22669);
and U23224 (N_23224,N_22496,N_22584);
or U23225 (N_23225,N_22313,N_22653);
or U23226 (N_23226,N_22202,N_22230);
xor U23227 (N_23227,N_22435,N_22225);
or U23228 (N_23228,N_22146,N_22517);
nor U23229 (N_23229,N_22791,N_22796);
nand U23230 (N_23230,N_22248,N_22821);
or U23231 (N_23231,N_22398,N_22044);
nor U23232 (N_23232,N_22459,N_22750);
nand U23233 (N_23233,N_22261,N_22729);
or U23234 (N_23234,N_22814,N_22993);
and U23235 (N_23235,N_22909,N_22181);
and U23236 (N_23236,N_22603,N_22841);
nand U23237 (N_23237,N_22031,N_22373);
xor U23238 (N_23238,N_22124,N_22920);
nor U23239 (N_23239,N_22284,N_22839);
or U23240 (N_23240,N_22533,N_22168);
and U23241 (N_23241,N_22967,N_22798);
nor U23242 (N_23242,N_22318,N_22505);
nand U23243 (N_23243,N_22480,N_22188);
xnor U23244 (N_23244,N_22657,N_22581);
nor U23245 (N_23245,N_22725,N_22515);
or U23246 (N_23246,N_22099,N_22715);
nand U23247 (N_23247,N_22863,N_22818);
nor U23248 (N_23248,N_22788,N_22675);
or U23249 (N_23249,N_22790,N_22797);
nor U23250 (N_23250,N_22104,N_22167);
nor U23251 (N_23251,N_22901,N_22840);
nand U23252 (N_23252,N_22360,N_22995);
nand U23253 (N_23253,N_22018,N_22573);
nand U23254 (N_23254,N_22580,N_22144);
or U23255 (N_23255,N_22337,N_22385);
or U23256 (N_23256,N_22117,N_22488);
or U23257 (N_23257,N_22393,N_22610);
nand U23258 (N_23258,N_22916,N_22881);
and U23259 (N_23259,N_22768,N_22985);
xnor U23260 (N_23260,N_22537,N_22766);
xor U23261 (N_23261,N_22658,N_22817);
xor U23262 (N_23262,N_22399,N_22478);
xnor U23263 (N_23263,N_22645,N_22885);
and U23264 (N_23264,N_22615,N_22698);
and U23265 (N_23265,N_22857,N_22291);
nand U23266 (N_23266,N_22819,N_22868);
nor U23267 (N_23267,N_22655,N_22776);
or U23268 (N_23268,N_22223,N_22600);
or U23269 (N_23269,N_22574,N_22663);
nor U23270 (N_23270,N_22413,N_22680);
xor U23271 (N_23271,N_22822,N_22384);
xnor U23272 (N_23272,N_22258,N_22743);
xnor U23273 (N_23273,N_22272,N_22094);
nand U23274 (N_23274,N_22141,N_22633);
or U23275 (N_23275,N_22806,N_22757);
or U23276 (N_23276,N_22236,N_22641);
or U23277 (N_23277,N_22737,N_22206);
or U23278 (N_23278,N_22397,N_22205);
or U23279 (N_23279,N_22887,N_22781);
nand U23280 (N_23280,N_22177,N_22122);
nand U23281 (N_23281,N_22120,N_22058);
nand U23282 (N_23282,N_22506,N_22754);
or U23283 (N_23283,N_22378,N_22252);
xnor U23284 (N_23284,N_22301,N_22096);
nor U23285 (N_23285,N_22443,N_22874);
nor U23286 (N_23286,N_22646,N_22057);
or U23287 (N_23287,N_22051,N_22388);
and U23288 (N_23288,N_22711,N_22136);
xnor U23289 (N_23289,N_22599,N_22345);
or U23290 (N_23290,N_22501,N_22326);
nor U23291 (N_23291,N_22024,N_22292);
xnor U23292 (N_23292,N_22870,N_22207);
and U23293 (N_23293,N_22278,N_22742);
nor U23294 (N_23294,N_22164,N_22733);
or U23295 (N_23295,N_22689,N_22845);
nand U23296 (N_23296,N_22241,N_22793);
nor U23297 (N_23297,N_22466,N_22983);
nor U23298 (N_23298,N_22552,N_22069);
and U23299 (N_23299,N_22090,N_22424);
nand U23300 (N_23300,N_22726,N_22457);
xnor U23301 (N_23301,N_22055,N_22888);
xnor U23302 (N_23302,N_22389,N_22081);
nor U23303 (N_23303,N_22508,N_22129);
xor U23304 (N_23304,N_22065,N_22854);
xor U23305 (N_23305,N_22608,N_22808);
xnor U23306 (N_23306,N_22029,N_22330);
nor U23307 (N_23307,N_22035,N_22493);
nand U23308 (N_23308,N_22110,N_22103);
nand U23309 (N_23309,N_22919,N_22756);
nor U23310 (N_23310,N_22805,N_22449);
or U23311 (N_23311,N_22980,N_22251);
nand U23312 (N_23312,N_22062,N_22941);
and U23313 (N_23313,N_22939,N_22882);
nand U23314 (N_23314,N_22604,N_22229);
and U23315 (N_23315,N_22156,N_22820);
nor U23316 (N_23316,N_22665,N_22595);
nand U23317 (N_23317,N_22150,N_22049);
or U23318 (N_23318,N_22410,N_22234);
nand U23319 (N_23319,N_22566,N_22336);
nor U23320 (N_23320,N_22067,N_22191);
nor U23321 (N_23321,N_22002,N_22497);
and U23322 (N_23322,N_22273,N_22323);
nand U23323 (N_23323,N_22034,N_22592);
nand U23324 (N_23324,N_22262,N_22991);
nor U23325 (N_23325,N_22157,N_22444);
and U23326 (N_23326,N_22456,N_22494);
nand U23327 (N_23327,N_22856,N_22585);
and U23328 (N_23328,N_22783,N_22153);
nand U23329 (N_23329,N_22714,N_22282);
xnor U23330 (N_23330,N_22218,N_22137);
nor U23331 (N_23331,N_22911,N_22986);
or U23332 (N_23332,N_22242,N_22351);
nand U23333 (N_23333,N_22368,N_22077);
xor U23334 (N_23334,N_22354,N_22746);
nand U23335 (N_23335,N_22316,N_22503);
xnor U23336 (N_23336,N_22255,N_22779);
and U23337 (N_23337,N_22162,N_22544);
or U23338 (N_23338,N_22312,N_22962);
nand U23339 (N_23339,N_22884,N_22617);
or U23340 (N_23340,N_22803,N_22523);
xnor U23341 (N_23341,N_22886,N_22527);
or U23342 (N_23342,N_22834,N_22926);
nand U23343 (N_23343,N_22507,N_22263);
and U23344 (N_23344,N_22172,N_22591);
and U23345 (N_23345,N_22173,N_22462);
and U23346 (N_23346,N_22183,N_22306);
xnor U23347 (N_23347,N_22064,N_22948);
or U23348 (N_23348,N_22158,N_22200);
nor U23349 (N_23349,N_22409,N_22133);
nor U23350 (N_23350,N_22245,N_22976);
nor U23351 (N_23351,N_22428,N_22249);
nand U23352 (N_23352,N_22159,N_22238);
or U23353 (N_23353,N_22001,N_22823);
nor U23354 (N_23354,N_22572,N_22450);
or U23355 (N_23355,N_22362,N_22917);
nand U23356 (N_23356,N_22964,N_22145);
or U23357 (N_23357,N_22576,N_22996);
and U23358 (N_23358,N_22407,N_22892);
xnor U23359 (N_23359,N_22492,N_22847);
xnor U23360 (N_23360,N_22913,N_22143);
and U23361 (N_23361,N_22084,N_22239);
nand U23362 (N_23362,N_22442,N_22811);
and U23363 (N_23363,N_22525,N_22047);
nor U23364 (N_23364,N_22196,N_22606);
and U23365 (N_23365,N_22642,N_22785);
and U23366 (N_23366,N_22540,N_22521);
nand U23367 (N_23367,N_22542,N_22490);
or U23368 (N_23368,N_22265,N_22340);
and U23369 (N_23369,N_22254,N_22656);
nand U23370 (N_23370,N_22430,N_22638);
or U23371 (N_23371,N_22915,N_22448);
nand U23372 (N_23372,N_22217,N_22846);
nor U23373 (N_23373,N_22895,N_22732);
and U23374 (N_23374,N_22161,N_22807);
or U23375 (N_23375,N_22904,N_22998);
and U23376 (N_23376,N_22224,N_22402);
and U23377 (N_23377,N_22474,N_22644);
nand U23378 (N_23378,N_22587,N_22063);
nand U23379 (N_23379,N_22624,N_22364);
xor U23380 (N_23380,N_22670,N_22679);
or U23381 (N_23381,N_22693,N_22486);
nor U23382 (N_23382,N_22543,N_22111);
nor U23383 (N_23383,N_22940,N_22041);
xor U23384 (N_23384,N_22040,N_22412);
or U23385 (N_23385,N_22147,N_22130);
nor U23386 (N_23386,N_22121,N_22836);
nand U23387 (N_23387,N_22914,N_22875);
nor U23388 (N_23388,N_22706,N_22227);
xnor U23389 (N_23389,N_22650,N_22891);
and U23390 (N_23390,N_22992,N_22718);
nand U23391 (N_23391,N_22799,N_22984);
xor U23392 (N_23392,N_22079,N_22890);
or U23393 (N_23393,N_22748,N_22009);
and U23394 (N_23394,N_22134,N_22317);
xor U23395 (N_23395,N_22905,N_22105);
nor U23396 (N_23396,N_22749,N_22755);
nand U23397 (N_23397,N_22201,N_22341);
and U23398 (N_23398,N_22954,N_22602);
xor U23399 (N_23399,N_22198,N_22668);
xor U23400 (N_23400,N_22285,N_22712);
xor U23401 (N_23401,N_22519,N_22702);
nand U23402 (N_23402,N_22751,N_22564);
nor U23403 (N_23403,N_22309,N_22060);
nand U23404 (N_23404,N_22142,N_22557);
or U23405 (N_23405,N_22464,N_22801);
nand U23406 (N_23406,N_22128,N_22843);
or U23407 (N_23407,N_22971,N_22734);
and U23408 (N_23408,N_22925,N_22346);
nand U23409 (N_23409,N_22924,N_22933);
xnor U23410 (N_23410,N_22950,N_22922);
nor U23411 (N_23411,N_22842,N_22880);
nor U23412 (N_23412,N_22233,N_22095);
nand U23413 (N_23413,N_22876,N_22465);
nand U23414 (N_23414,N_22550,N_22908);
nor U23415 (N_23415,N_22661,N_22228);
xnor U23416 (N_23416,N_22097,N_22334);
nand U23417 (N_23417,N_22420,N_22692);
and U23418 (N_23418,N_22379,N_22195);
or U23419 (N_23419,N_22832,N_22294);
and U23420 (N_23420,N_22762,N_22871);
xor U23421 (N_23421,N_22154,N_22741);
xnor U23422 (N_23422,N_22931,N_22945);
nor U23423 (N_23423,N_22003,N_22182);
xor U23424 (N_23424,N_22072,N_22589);
nor U23425 (N_23425,N_22376,N_22960);
and U23426 (N_23426,N_22724,N_22596);
nor U23427 (N_23427,N_22484,N_22418);
nand U23428 (N_23428,N_22220,N_22461);
nor U23429 (N_23429,N_22193,N_22630);
or U23430 (N_23430,N_22216,N_22329);
and U23431 (N_23431,N_22660,N_22848);
xor U23432 (N_23432,N_22178,N_22877);
nand U23433 (N_23433,N_22331,N_22131);
and U23434 (N_23434,N_22215,N_22299);
nor U23435 (N_23435,N_22098,N_22401);
or U23436 (N_23436,N_22452,N_22643);
xnor U23437 (N_23437,N_22314,N_22427);
xnor U23438 (N_23438,N_22683,N_22625);
xnor U23439 (N_23439,N_22896,N_22032);
xnor U23440 (N_23440,N_22855,N_22545);
nor U23441 (N_23441,N_22297,N_22534);
nand U23442 (N_23442,N_22367,N_22441);
and U23443 (N_23443,N_22568,N_22701);
nand U23444 (N_23444,N_22898,N_22011);
xnor U23445 (N_23445,N_22771,N_22080);
nand U23446 (N_23446,N_22140,N_22068);
nand U23447 (N_23447,N_22170,N_22511);
nand U23448 (N_23448,N_22476,N_22965);
or U23449 (N_23449,N_22999,N_22662);
xor U23450 (N_23450,N_22425,N_22071);
nor U23451 (N_23451,N_22453,N_22747);
and U23452 (N_23452,N_22434,N_22310);
nand U23453 (N_23453,N_22831,N_22184);
xnor U23454 (N_23454,N_22267,N_22981);
and U23455 (N_23455,N_22481,N_22934);
xnor U23456 (N_23456,N_22970,N_22008);
xnor U23457 (N_23457,N_22489,N_22155);
nor U23458 (N_23458,N_22160,N_22197);
nor U23459 (N_23459,N_22046,N_22307);
xnor U23460 (N_23460,N_22767,N_22666);
and U23461 (N_23461,N_22994,N_22365);
nand U23462 (N_23462,N_22695,N_22979);
or U23463 (N_23463,N_22598,N_22676);
and U23464 (N_23464,N_22621,N_22387);
or U23465 (N_23465,N_22208,N_22015);
nor U23466 (N_23466,N_22526,N_22366);
nand U23467 (N_23467,N_22532,N_22601);
xor U23468 (N_23468,N_22126,N_22390);
nor U23469 (N_23469,N_22375,N_22900);
xor U23470 (N_23470,N_22280,N_22319);
nor U23471 (N_23471,N_22879,N_22296);
or U23472 (N_23472,N_22289,N_22485);
nand U23473 (N_23473,N_22620,N_22221);
xor U23474 (N_23474,N_22977,N_22963);
nand U23475 (N_23475,N_22921,N_22083);
or U23476 (N_23476,N_22213,N_22043);
or U23477 (N_23477,N_22780,N_22274);
nor U23478 (N_23478,N_22467,N_22422);
nand U23479 (N_23479,N_22713,N_22889);
or U23480 (N_23480,N_22437,N_22636);
nand U23481 (N_23481,N_22745,N_22635);
nand U23482 (N_23482,N_22298,N_22973);
nor U23483 (N_23483,N_22070,N_22381);
xnor U23484 (N_23484,N_22782,N_22502);
or U23485 (N_23485,N_22773,N_22764);
xnor U23486 (N_23486,N_22253,N_22308);
nor U23487 (N_23487,N_22593,N_22271);
and U23488 (N_23488,N_22290,N_22827);
and U23489 (N_23489,N_22471,N_22075);
nor U23490 (N_23490,N_22165,N_22396);
nor U23491 (N_23491,N_22866,N_22333);
nand U23492 (N_23492,N_22957,N_22004);
nand U23493 (N_23493,N_22571,N_22524);
xor U23494 (N_23494,N_22460,N_22118);
or U23495 (N_23495,N_22555,N_22652);
nand U23496 (N_23496,N_22673,N_22321);
and U23497 (N_23497,N_22359,N_22169);
nand U23498 (N_23498,N_22778,N_22209);
or U23499 (N_23499,N_22468,N_22632);
xor U23500 (N_23500,N_22523,N_22858);
or U23501 (N_23501,N_22943,N_22819);
and U23502 (N_23502,N_22523,N_22647);
xnor U23503 (N_23503,N_22710,N_22124);
nand U23504 (N_23504,N_22553,N_22495);
nor U23505 (N_23505,N_22035,N_22430);
or U23506 (N_23506,N_22935,N_22812);
nor U23507 (N_23507,N_22934,N_22885);
and U23508 (N_23508,N_22121,N_22609);
xnor U23509 (N_23509,N_22147,N_22279);
xor U23510 (N_23510,N_22176,N_22903);
nor U23511 (N_23511,N_22966,N_22277);
or U23512 (N_23512,N_22721,N_22504);
and U23513 (N_23513,N_22754,N_22383);
nand U23514 (N_23514,N_22353,N_22188);
xor U23515 (N_23515,N_22443,N_22027);
nand U23516 (N_23516,N_22279,N_22927);
or U23517 (N_23517,N_22390,N_22432);
xnor U23518 (N_23518,N_22743,N_22467);
xnor U23519 (N_23519,N_22975,N_22982);
and U23520 (N_23520,N_22656,N_22888);
xor U23521 (N_23521,N_22292,N_22917);
nand U23522 (N_23522,N_22063,N_22887);
and U23523 (N_23523,N_22641,N_22343);
or U23524 (N_23524,N_22440,N_22617);
nor U23525 (N_23525,N_22358,N_22144);
nor U23526 (N_23526,N_22409,N_22172);
nor U23527 (N_23527,N_22240,N_22418);
nor U23528 (N_23528,N_22588,N_22352);
nand U23529 (N_23529,N_22986,N_22487);
nor U23530 (N_23530,N_22822,N_22543);
nand U23531 (N_23531,N_22146,N_22856);
xnor U23532 (N_23532,N_22586,N_22995);
nor U23533 (N_23533,N_22556,N_22836);
xnor U23534 (N_23534,N_22513,N_22329);
nor U23535 (N_23535,N_22016,N_22096);
nand U23536 (N_23536,N_22481,N_22807);
nor U23537 (N_23537,N_22436,N_22806);
and U23538 (N_23538,N_22161,N_22239);
nand U23539 (N_23539,N_22409,N_22106);
and U23540 (N_23540,N_22851,N_22284);
xnor U23541 (N_23541,N_22688,N_22601);
nor U23542 (N_23542,N_22307,N_22781);
nor U23543 (N_23543,N_22535,N_22042);
xor U23544 (N_23544,N_22664,N_22385);
nand U23545 (N_23545,N_22000,N_22134);
nor U23546 (N_23546,N_22632,N_22578);
nor U23547 (N_23547,N_22841,N_22349);
nor U23548 (N_23548,N_22623,N_22147);
and U23549 (N_23549,N_22818,N_22963);
xor U23550 (N_23550,N_22377,N_22708);
nand U23551 (N_23551,N_22296,N_22851);
nor U23552 (N_23552,N_22342,N_22779);
nor U23553 (N_23553,N_22537,N_22034);
nand U23554 (N_23554,N_22033,N_22426);
xor U23555 (N_23555,N_22530,N_22509);
nand U23556 (N_23556,N_22589,N_22413);
or U23557 (N_23557,N_22378,N_22808);
nor U23558 (N_23558,N_22645,N_22015);
xnor U23559 (N_23559,N_22407,N_22951);
and U23560 (N_23560,N_22913,N_22447);
xor U23561 (N_23561,N_22421,N_22417);
nor U23562 (N_23562,N_22231,N_22729);
or U23563 (N_23563,N_22095,N_22487);
or U23564 (N_23564,N_22413,N_22844);
nor U23565 (N_23565,N_22391,N_22918);
xor U23566 (N_23566,N_22443,N_22545);
nand U23567 (N_23567,N_22611,N_22231);
nand U23568 (N_23568,N_22777,N_22215);
nor U23569 (N_23569,N_22224,N_22689);
or U23570 (N_23570,N_22383,N_22781);
nand U23571 (N_23571,N_22580,N_22907);
nand U23572 (N_23572,N_22286,N_22863);
and U23573 (N_23573,N_22192,N_22699);
nor U23574 (N_23574,N_22260,N_22498);
nor U23575 (N_23575,N_22149,N_22439);
nor U23576 (N_23576,N_22090,N_22862);
or U23577 (N_23577,N_22086,N_22479);
nor U23578 (N_23578,N_22186,N_22841);
or U23579 (N_23579,N_22841,N_22013);
or U23580 (N_23580,N_22230,N_22329);
nand U23581 (N_23581,N_22080,N_22315);
xor U23582 (N_23582,N_22055,N_22722);
nand U23583 (N_23583,N_22163,N_22071);
xnor U23584 (N_23584,N_22864,N_22419);
nand U23585 (N_23585,N_22501,N_22583);
or U23586 (N_23586,N_22086,N_22435);
or U23587 (N_23587,N_22693,N_22561);
or U23588 (N_23588,N_22788,N_22100);
nand U23589 (N_23589,N_22570,N_22858);
xnor U23590 (N_23590,N_22698,N_22476);
xnor U23591 (N_23591,N_22159,N_22488);
xnor U23592 (N_23592,N_22509,N_22740);
nand U23593 (N_23593,N_22683,N_22133);
nand U23594 (N_23594,N_22712,N_22384);
or U23595 (N_23595,N_22996,N_22970);
or U23596 (N_23596,N_22345,N_22251);
or U23597 (N_23597,N_22759,N_22726);
xor U23598 (N_23598,N_22955,N_22416);
xor U23599 (N_23599,N_22461,N_22489);
nand U23600 (N_23600,N_22652,N_22946);
and U23601 (N_23601,N_22482,N_22883);
nand U23602 (N_23602,N_22796,N_22864);
and U23603 (N_23603,N_22371,N_22989);
nand U23604 (N_23604,N_22326,N_22624);
nor U23605 (N_23605,N_22700,N_22414);
xor U23606 (N_23606,N_22015,N_22575);
and U23607 (N_23607,N_22682,N_22908);
nand U23608 (N_23608,N_22306,N_22685);
nor U23609 (N_23609,N_22040,N_22962);
nand U23610 (N_23610,N_22198,N_22320);
xnor U23611 (N_23611,N_22882,N_22636);
nand U23612 (N_23612,N_22162,N_22238);
xnor U23613 (N_23613,N_22522,N_22129);
nand U23614 (N_23614,N_22371,N_22857);
or U23615 (N_23615,N_22291,N_22189);
nor U23616 (N_23616,N_22321,N_22697);
xnor U23617 (N_23617,N_22275,N_22059);
nand U23618 (N_23618,N_22974,N_22613);
or U23619 (N_23619,N_22116,N_22811);
xnor U23620 (N_23620,N_22531,N_22757);
and U23621 (N_23621,N_22939,N_22274);
or U23622 (N_23622,N_22210,N_22442);
nand U23623 (N_23623,N_22393,N_22354);
nor U23624 (N_23624,N_22593,N_22397);
or U23625 (N_23625,N_22711,N_22399);
xnor U23626 (N_23626,N_22319,N_22681);
nor U23627 (N_23627,N_22460,N_22073);
nand U23628 (N_23628,N_22744,N_22654);
or U23629 (N_23629,N_22244,N_22660);
or U23630 (N_23630,N_22605,N_22369);
nand U23631 (N_23631,N_22224,N_22904);
nor U23632 (N_23632,N_22143,N_22734);
and U23633 (N_23633,N_22375,N_22239);
and U23634 (N_23634,N_22614,N_22397);
nand U23635 (N_23635,N_22766,N_22916);
and U23636 (N_23636,N_22496,N_22868);
or U23637 (N_23637,N_22106,N_22344);
nor U23638 (N_23638,N_22442,N_22541);
xnor U23639 (N_23639,N_22747,N_22471);
nand U23640 (N_23640,N_22951,N_22674);
or U23641 (N_23641,N_22290,N_22255);
nand U23642 (N_23642,N_22860,N_22430);
or U23643 (N_23643,N_22833,N_22426);
and U23644 (N_23644,N_22095,N_22352);
nor U23645 (N_23645,N_22286,N_22829);
nand U23646 (N_23646,N_22604,N_22702);
and U23647 (N_23647,N_22651,N_22359);
nor U23648 (N_23648,N_22880,N_22371);
nand U23649 (N_23649,N_22415,N_22913);
or U23650 (N_23650,N_22496,N_22748);
nor U23651 (N_23651,N_22939,N_22443);
or U23652 (N_23652,N_22721,N_22963);
xor U23653 (N_23653,N_22166,N_22951);
xnor U23654 (N_23654,N_22283,N_22268);
xnor U23655 (N_23655,N_22476,N_22709);
nor U23656 (N_23656,N_22726,N_22233);
nand U23657 (N_23657,N_22490,N_22981);
nand U23658 (N_23658,N_22437,N_22204);
and U23659 (N_23659,N_22588,N_22721);
and U23660 (N_23660,N_22840,N_22833);
or U23661 (N_23661,N_22457,N_22462);
nor U23662 (N_23662,N_22436,N_22977);
or U23663 (N_23663,N_22149,N_22353);
nor U23664 (N_23664,N_22567,N_22873);
and U23665 (N_23665,N_22853,N_22033);
xnor U23666 (N_23666,N_22485,N_22438);
xnor U23667 (N_23667,N_22506,N_22953);
or U23668 (N_23668,N_22468,N_22720);
xnor U23669 (N_23669,N_22399,N_22811);
nand U23670 (N_23670,N_22237,N_22593);
or U23671 (N_23671,N_22384,N_22587);
nand U23672 (N_23672,N_22477,N_22989);
or U23673 (N_23673,N_22835,N_22823);
or U23674 (N_23674,N_22727,N_22852);
or U23675 (N_23675,N_22165,N_22208);
nor U23676 (N_23676,N_22762,N_22054);
or U23677 (N_23677,N_22569,N_22302);
xnor U23678 (N_23678,N_22656,N_22878);
and U23679 (N_23679,N_22307,N_22869);
and U23680 (N_23680,N_22904,N_22993);
xnor U23681 (N_23681,N_22531,N_22292);
nor U23682 (N_23682,N_22193,N_22673);
or U23683 (N_23683,N_22941,N_22348);
nor U23684 (N_23684,N_22428,N_22972);
and U23685 (N_23685,N_22826,N_22081);
and U23686 (N_23686,N_22680,N_22948);
nand U23687 (N_23687,N_22514,N_22668);
or U23688 (N_23688,N_22217,N_22019);
nor U23689 (N_23689,N_22422,N_22237);
or U23690 (N_23690,N_22494,N_22245);
nor U23691 (N_23691,N_22729,N_22976);
or U23692 (N_23692,N_22551,N_22071);
and U23693 (N_23693,N_22689,N_22104);
or U23694 (N_23694,N_22892,N_22399);
nand U23695 (N_23695,N_22312,N_22122);
and U23696 (N_23696,N_22967,N_22707);
or U23697 (N_23697,N_22055,N_22209);
or U23698 (N_23698,N_22327,N_22461);
xnor U23699 (N_23699,N_22621,N_22637);
or U23700 (N_23700,N_22599,N_22866);
or U23701 (N_23701,N_22733,N_22041);
and U23702 (N_23702,N_22122,N_22093);
nor U23703 (N_23703,N_22952,N_22706);
nand U23704 (N_23704,N_22323,N_22961);
xor U23705 (N_23705,N_22567,N_22944);
or U23706 (N_23706,N_22518,N_22596);
xor U23707 (N_23707,N_22536,N_22938);
and U23708 (N_23708,N_22749,N_22801);
nand U23709 (N_23709,N_22257,N_22477);
and U23710 (N_23710,N_22716,N_22367);
nor U23711 (N_23711,N_22097,N_22760);
nor U23712 (N_23712,N_22111,N_22199);
nand U23713 (N_23713,N_22090,N_22070);
xnor U23714 (N_23714,N_22506,N_22489);
or U23715 (N_23715,N_22297,N_22601);
and U23716 (N_23716,N_22707,N_22629);
nand U23717 (N_23717,N_22777,N_22095);
nor U23718 (N_23718,N_22108,N_22417);
xor U23719 (N_23719,N_22766,N_22056);
nand U23720 (N_23720,N_22814,N_22185);
xnor U23721 (N_23721,N_22729,N_22504);
or U23722 (N_23722,N_22655,N_22893);
nand U23723 (N_23723,N_22493,N_22012);
nor U23724 (N_23724,N_22059,N_22630);
or U23725 (N_23725,N_22168,N_22120);
and U23726 (N_23726,N_22570,N_22300);
nor U23727 (N_23727,N_22885,N_22202);
xnor U23728 (N_23728,N_22490,N_22262);
and U23729 (N_23729,N_22791,N_22091);
and U23730 (N_23730,N_22252,N_22144);
xor U23731 (N_23731,N_22750,N_22043);
xor U23732 (N_23732,N_22330,N_22262);
xor U23733 (N_23733,N_22822,N_22425);
or U23734 (N_23734,N_22848,N_22800);
and U23735 (N_23735,N_22965,N_22939);
nor U23736 (N_23736,N_22064,N_22495);
or U23737 (N_23737,N_22469,N_22246);
xnor U23738 (N_23738,N_22430,N_22720);
and U23739 (N_23739,N_22665,N_22154);
and U23740 (N_23740,N_22909,N_22492);
and U23741 (N_23741,N_22753,N_22720);
nor U23742 (N_23742,N_22441,N_22705);
xnor U23743 (N_23743,N_22888,N_22155);
nor U23744 (N_23744,N_22332,N_22225);
or U23745 (N_23745,N_22398,N_22994);
or U23746 (N_23746,N_22355,N_22331);
nor U23747 (N_23747,N_22952,N_22904);
or U23748 (N_23748,N_22827,N_22356);
or U23749 (N_23749,N_22013,N_22484);
nand U23750 (N_23750,N_22330,N_22479);
nand U23751 (N_23751,N_22259,N_22378);
or U23752 (N_23752,N_22490,N_22319);
nor U23753 (N_23753,N_22830,N_22717);
nor U23754 (N_23754,N_22185,N_22253);
and U23755 (N_23755,N_22053,N_22985);
or U23756 (N_23756,N_22154,N_22579);
nor U23757 (N_23757,N_22742,N_22195);
nor U23758 (N_23758,N_22084,N_22295);
xor U23759 (N_23759,N_22987,N_22774);
nand U23760 (N_23760,N_22853,N_22420);
and U23761 (N_23761,N_22283,N_22345);
and U23762 (N_23762,N_22873,N_22988);
nand U23763 (N_23763,N_22469,N_22500);
or U23764 (N_23764,N_22082,N_22276);
or U23765 (N_23765,N_22458,N_22768);
nor U23766 (N_23766,N_22900,N_22930);
or U23767 (N_23767,N_22254,N_22354);
nand U23768 (N_23768,N_22502,N_22645);
nor U23769 (N_23769,N_22045,N_22816);
or U23770 (N_23770,N_22962,N_22388);
xor U23771 (N_23771,N_22359,N_22084);
nor U23772 (N_23772,N_22129,N_22293);
nand U23773 (N_23773,N_22348,N_22987);
and U23774 (N_23774,N_22264,N_22709);
xor U23775 (N_23775,N_22240,N_22049);
or U23776 (N_23776,N_22237,N_22412);
nor U23777 (N_23777,N_22982,N_22918);
xor U23778 (N_23778,N_22194,N_22277);
nand U23779 (N_23779,N_22834,N_22095);
nor U23780 (N_23780,N_22172,N_22157);
nand U23781 (N_23781,N_22424,N_22047);
nand U23782 (N_23782,N_22934,N_22960);
xor U23783 (N_23783,N_22987,N_22682);
and U23784 (N_23784,N_22452,N_22627);
xnor U23785 (N_23785,N_22480,N_22950);
or U23786 (N_23786,N_22739,N_22433);
and U23787 (N_23787,N_22503,N_22895);
nand U23788 (N_23788,N_22340,N_22803);
nor U23789 (N_23789,N_22513,N_22376);
and U23790 (N_23790,N_22984,N_22967);
xnor U23791 (N_23791,N_22949,N_22221);
xor U23792 (N_23792,N_22582,N_22004);
and U23793 (N_23793,N_22176,N_22223);
xnor U23794 (N_23794,N_22603,N_22599);
xor U23795 (N_23795,N_22663,N_22367);
or U23796 (N_23796,N_22456,N_22851);
and U23797 (N_23797,N_22889,N_22904);
xor U23798 (N_23798,N_22097,N_22252);
nor U23799 (N_23799,N_22243,N_22151);
and U23800 (N_23800,N_22093,N_22748);
nor U23801 (N_23801,N_22461,N_22242);
nand U23802 (N_23802,N_22295,N_22169);
or U23803 (N_23803,N_22807,N_22305);
xor U23804 (N_23804,N_22971,N_22537);
and U23805 (N_23805,N_22027,N_22767);
nor U23806 (N_23806,N_22351,N_22352);
or U23807 (N_23807,N_22273,N_22647);
and U23808 (N_23808,N_22667,N_22912);
xor U23809 (N_23809,N_22328,N_22628);
or U23810 (N_23810,N_22669,N_22548);
nand U23811 (N_23811,N_22070,N_22541);
nand U23812 (N_23812,N_22572,N_22585);
xnor U23813 (N_23813,N_22689,N_22405);
xor U23814 (N_23814,N_22999,N_22733);
nor U23815 (N_23815,N_22089,N_22644);
and U23816 (N_23816,N_22912,N_22366);
nand U23817 (N_23817,N_22621,N_22983);
nand U23818 (N_23818,N_22243,N_22024);
nand U23819 (N_23819,N_22317,N_22497);
and U23820 (N_23820,N_22258,N_22752);
xnor U23821 (N_23821,N_22044,N_22270);
and U23822 (N_23822,N_22488,N_22118);
and U23823 (N_23823,N_22320,N_22896);
xor U23824 (N_23824,N_22640,N_22923);
xor U23825 (N_23825,N_22976,N_22785);
and U23826 (N_23826,N_22108,N_22924);
nand U23827 (N_23827,N_22428,N_22815);
or U23828 (N_23828,N_22656,N_22979);
and U23829 (N_23829,N_22416,N_22269);
nor U23830 (N_23830,N_22397,N_22525);
or U23831 (N_23831,N_22552,N_22766);
nor U23832 (N_23832,N_22328,N_22092);
and U23833 (N_23833,N_22798,N_22192);
and U23834 (N_23834,N_22194,N_22247);
and U23835 (N_23835,N_22487,N_22838);
and U23836 (N_23836,N_22569,N_22487);
and U23837 (N_23837,N_22270,N_22211);
nor U23838 (N_23838,N_22925,N_22910);
and U23839 (N_23839,N_22019,N_22747);
xor U23840 (N_23840,N_22304,N_22408);
nand U23841 (N_23841,N_22687,N_22699);
nand U23842 (N_23842,N_22624,N_22023);
xnor U23843 (N_23843,N_22866,N_22831);
or U23844 (N_23844,N_22252,N_22361);
or U23845 (N_23845,N_22713,N_22784);
xor U23846 (N_23846,N_22712,N_22434);
and U23847 (N_23847,N_22336,N_22632);
and U23848 (N_23848,N_22905,N_22762);
nand U23849 (N_23849,N_22115,N_22458);
and U23850 (N_23850,N_22135,N_22613);
and U23851 (N_23851,N_22125,N_22937);
xnor U23852 (N_23852,N_22291,N_22373);
xor U23853 (N_23853,N_22925,N_22612);
nor U23854 (N_23854,N_22222,N_22249);
nor U23855 (N_23855,N_22434,N_22868);
and U23856 (N_23856,N_22212,N_22022);
and U23857 (N_23857,N_22477,N_22627);
xnor U23858 (N_23858,N_22794,N_22217);
nor U23859 (N_23859,N_22777,N_22201);
xnor U23860 (N_23860,N_22792,N_22998);
nor U23861 (N_23861,N_22941,N_22034);
nor U23862 (N_23862,N_22329,N_22198);
or U23863 (N_23863,N_22949,N_22986);
nand U23864 (N_23864,N_22830,N_22067);
nor U23865 (N_23865,N_22920,N_22364);
nor U23866 (N_23866,N_22700,N_22841);
nand U23867 (N_23867,N_22900,N_22578);
xnor U23868 (N_23868,N_22633,N_22801);
and U23869 (N_23869,N_22644,N_22616);
nor U23870 (N_23870,N_22115,N_22983);
or U23871 (N_23871,N_22056,N_22166);
and U23872 (N_23872,N_22340,N_22810);
or U23873 (N_23873,N_22014,N_22900);
and U23874 (N_23874,N_22717,N_22769);
nand U23875 (N_23875,N_22353,N_22064);
and U23876 (N_23876,N_22577,N_22561);
nand U23877 (N_23877,N_22554,N_22464);
nor U23878 (N_23878,N_22014,N_22874);
or U23879 (N_23879,N_22206,N_22900);
or U23880 (N_23880,N_22610,N_22749);
and U23881 (N_23881,N_22463,N_22805);
xor U23882 (N_23882,N_22396,N_22139);
xnor U23883 (N_23883,N_22596,N_22981);
xor U23884 (N_23884,N_22155,N_22457);
nor U23885 (N_23885,N_22689,N_22612);
or U23886 (N_23886,N_22814,N_22756);
nor U23887 (N_23887,N_22474,N_22252);
or U23888 (N_23888,N_22301,N_22365);
nor U23889 (N_23889,N_22025,N_22236);
and U23890 (N_23890,N_22053,N_22203);
nand U23891 (N_23891,N_22542,N_22132);
xnor U23892 (N_23892,N_22105,N_22658);
xnor U23893 (N_23893,N_22539,N_22936);
xor U23894 (N_23894,N_22222,N_22615);
and U23895 (N_23895,N_22844,N_22900);
nand U23896 (N_23896,N_22929,N_22253);
or U23897 (N_23897,N_22396,N_22374);
nand U23898 (N_23898,N_22002,N_22523);
nand U23899 (N_23899,N_22526,N_22903);
nor U23900 (N_23900,N_22832,N_22018);
or U23901 (N_23901,N_22139,N_22076);
nand U23902 (N_23902,N_22653,N_22719);
nand U23903 (N_23903,N_22176,N_22339);
xnor U23904 (N_23904,N_22007,N_22595);
nor U23905 (N_23905,N_22676,N_22047);
and U23906 (N_23906,N_22467,N_22219);
xnor U23907 (N_23907,N_22446,N_22961);
xnor U23908 (N_23908,N_22505,N_22638);
nor U23909 (N_23909,N_22815,N_22570);
or U23910 (N_23910,N_22475,N_22685);
xor U23911 (N_23911,N_22692,N_22975);
nor U23912 (N_23912,N_22411,N_22410);
nand U23913 (N_23913,N_22394,N_22724);
nand U23914 (N_23914,N_22293,N_22327);
or U23915 (N_23915,N_22718,N_22985);
and U23916 (N_23916,N_22721,N_22047);
nand U23917 (N_23917,N_22026,N_22573);
or U23918 (N_23918,N_22762,N_22397);
nor U23919 (N_23919,N_22737,N_22142);
or U23920 (N_23920,N_22517,N_22528);
nor U23921 (N_23921,N_22993,N_22439);
or U23922 (N_23922,N_22768,N_22797);
xor U23923 (N_23923,N_22226,N_22954);
nand U23924 (N_23924,N_22254,N_22683);
or U23925 (N_23925,N_22555,N_22552);
xnor U23926 (N_23926,N_22375,N_22494);
nor U23927 (N_23927,N_22028,N_22923);
nor U23928 (N_23928,N_22749,N_22144);
nor U23929 (N_23929,N_22126,N_22173);
xor U23930 (N_23930,N_22564,N_22019);
and U23931 (N_23931,N_22519,N_22555);
or U23932 (N_23932,N_22926,N_22458);
nand U23933 (N_23933,N_22829,N_22489);
and U23934 (N_23934,N_22084,N_22303);
nor U23935 (N_23935,N_22881,N_22555);
xnor U23936 (N_23936,N_22653,N_22381);
or U23937 (N_23937,N_22582,N_22542);
nor U23938 (N_23938,N_22011,N_22219);
nor U23939 (N_23939,N_22721,N_22366);
nor U23940 (N_23940,N_22323,N_22243);
nand U23941 (N_23941,N_22004,N_22670);
and U23942 (N_23942,N_22489,N_22599);
xor U23943 (N_23943,N_22209,N_22902);
and U23944 (N_23944,N_22343,N_22589);
nor U23945 (N_23945,N_22822,N_22775);
nor U23946 (N_23946,N_22061,N_22510);
and U23947 (N_23947,N_22111,N_22979);
nand U23948 (N_23948,N_22314,N_22135);
or U23949 (N_23949,N_22618,N_22759);
xor U23950 (N_23950,N_22944,N_22153);
or U23951 (N_23951,N_22105,N_22237);
and U23952 (N_23952,N_22529,N_22237);
nor U23953 (N_23953,N_22754,N_22304);
nand U23954 (N_23954,N_22824,N_22900);
and U23955 (N_23955,N_22542,N_22368);
and U23956 (N_23956,N_22651,N_22820);
xnor U23957 (N_23957,N_22463,N_22629);
xor U23958 (N_23958,N_22576,N_22137);
and U23959 (N_23959,N_22779,N_22301);
nor U23960 (N_23960,N_22387,N_22335);
and U23961 (N_23961,N_22259,N_22352);
xnor U23962 (N_23962,N_22107,N_22204);
nor U23963 (N_23963,N_22329,N_22316);
or U23964 (N_23964,N_22310,N_22823);
nand U23965 (N_23965,N_22903,N_22227);
nand U23966 (N_23966,N_22743,N_22222);
or U23967 (N_23967,N_22825,N_22096);
and U23968 (N_23968,N_22548,N_22235);
nand U23969 (N_23969,N_22331,N_22169);
and U23970 (N_23970,N_22860,N_22990);
nor U23971 (N_23971,N_22978,N_22524);
or U23972 (N_23972,N_22921,N_22816);
nand U23973 (N_23973,N_22602,N_22938);
nand U23974 (N_23974,N_22665,N_22589);
nand U23975 (N_23975,N_22261,N_22185);
and U23976 (N_23976,N_22424,N_22820);
nand U23977 (N_23977,N_22792,N_22098);
nor U23978 (N_23978,N_22320,N_22981);
or U23979 (N_23979,N_22320,N_22495);
xnor U23980 (N_23980,N_22324,N_22794);
nor U23981 (N_23981,N_22851,N_22776);
nand U23982 (N_23982,N_22281,N_22788);
or U23983 (N_23983,N_22933,N_22176);
nor U23984 (N_23984,N_22283,N_22002);
nor U23985 (N_23985,N_22183,N_22732);
nand U23986 (N_23986,N_22019,N_22039);
and U23987 (N_23987,N_22437,N_22008);
xnor U23988 (N_23988,N_22417,N_22539);
nand U23989 (N_23989,N_22031,N_22346);
nor U23990 (N_23990,N_22460,N_22583);
nor U23991 (N_23991,N_22770,N_22326);
and U23992 (N_23992,N_22040,N_22178);
and U23993 (N_23993,N_22257,N_22997);
and U23994 (N_23994,N_22926,N_22756);
xnor U23995 (N_23995,N_22436,N_22696);
and U23996 (N_23996,N_22725,N_22143);
xor U23997 (N_23997,N_22839,N_22930);
and U23998 (N_23998,N_22114,N_22218);
nor U23999 (N_23999,N_22412,N_22340);
nand U24000 (N_24000,N_23525,N_23513);
nand U24001 (N_24001,N_23278,N_23779);
nand U24002 (N_24002,N_23687,N_23579);
and U24003 (N_24003,N_23068,N_23038);
xnor U24004 (N_24004,N_23137,N_23328);
nor U24005 (N_24005,N_23797,N_23150);
or U24006 (N_24006,N_23645,N_23059);
nand U24007 (N_24007,N_23171,N_23776);
or U24008 (N_24008,N_23417,N_23808);
xor U24009 (N_24009,N_23860,N_23652);
or U24010 (N_24010,N_23330,N_23706);
nand U24011 (N_24011,N_23932,N_23662);
xnor U24012 (N_24012,N_23156,N_23358);
nand U24013 (N_24013,N_23405,N_23683);
xnor U24014 (N_24014,N_23173,N_23206);
and U24015 (N_24015,N_23461,N_23226);
or U24016 (N_24016,N_23654,N_23664);
xor U24017 (N_24017,N_23164,N_23750);
or U24018 (N_24018,N_23688,N_23462);
nor U24019 (N_24019,N_23876,N_23445);
nor U24020 (N_24020,N_23300,N_23239);
and U24021 (N_24021,N_23773,N_23718);
nor U24022 (N_24022,N_23653,N_23188);
xnor U24023 (N_24023,N_23637,N_23472);
nor U24024 (N_24024,N_23191,N_23460);
nand U24025 (N_24025,N_23064,N_23276);
nor U24026 (N_24026,N_23177,N_23163);
or U24027 (N_24027,N_23247,N_23283);
and U24028 (N_24028,N_23279,N_23946);
xor U24029 (N_24029,N_23108,N_23784);
and U24030 (N_24030,N_23160,N_23744);
nor U24031 (N_24031,N_23721,N_23891);
nand U24032 (N_24032,N_23404,N_23319);
nand U24033 (N_24033,N_23923,N_23015);
or U24034 (N_24034,N_23062,N_23293);
or U24035 (N_24035,N_23117,N_23303);
nand U24036 (N_24036,N_23848,N_23692);
nor U24037 (N_24037,N_23847,N_23408);
nor U24038 (N_24038,N_23092,N_23909);
xnor U24039 (N_24039,N_23730,N_23903);
or U24040 (N_24040,N_23524,N_23954);
nand U24041 (N_24041,N_23597,N_23185);
xnor U24042 (N_24042,N_23864,N_23559);
nand U24043 (N_24043,N_23898,N_23257);
nor U24044 (N_24044,N_23421,N_23798);
nand U24045 (N_24045,N_23021,N_23512);
nor U24046 (N_24046,N_23691,N_23456);
or U24047 (N_24047,N_23708,N_23577);
or U24048 (N_24048,N_23621,N_23235);
or U24049 (N_24049,N_23424,N_23429);
nor U24050 (N_24050,N_23819,N_23938);
xor U24051 (N_24051,N_23782,N_23071);
nor U24052 (N_24052,N_23479,N_23097);
or U24053 (N_24053,N_23605,N_23237);
xor U24054 (N_24054,N_23942,N_23659);
or U24055 (N_24055,N_23740,N_23897);
and U24056 (N_24056,N_23965,N_23961);
xor U24057 (N_24057,N_23990,N_23478);
or U24058 (N_24058,N_23701,N_23075);
nand U24059 (N_24059,N_23355,N_23553);
nor U24060 (N_24060,N_23363,N_23918);
and U24061 (N_24061,N_23305,N_23713);
and U24062 (N_24062,N_23366,N_23100);
and U24063 (N_24063,N_23049,N_23018);
or U24064 (N_24064,N_23787,N_23403);
and U24065 (N_24065,N_23801,N_23480);
and U24066 (N_24066,N_23045,N_23501);
nor U24067 (N_24067,N_23988,N_23302);
nor U24068 (N_24068,N_23287,N_23763);
or U24069 (N_24069,N_23452,N_23994);
or U24070 (N_24070,N_23896,N_23707);
xnor U24071 (N_24071,N_23837,N_23865);
nor U24072 (N_24072,N_23074,N_23322);
or U24073 (N_24073,N_23552,N_23246);
nand U24074 (N_24074,N_23975,N_23192);
nor U24075 (N_24075,N_23518,N_23116);
xnor U24076 (N_24076,N_23600,N_23202);
nand U24077 (N_24077,N_23588,N_23667);
or U24078 (N_24078,N_23436,N_23207);
xnor U24079 (N_24079,N_23581,N_23218);
and U24080 (N_24080,N_23810,N_23323);
nor U24081 (N_24081,N_23894,N_23329);
or U24082 (N_24082,N_23282,N_23829);
nand U24083 (N_24083,N_23504,N_23020);
and U24084 (N_24084,N_23011,N_23873);
or U24085 (N_24085,N_23034,N_23746);
or U24086 (N_24086,N_23105,N_23422);
or U24087 (N_24087,N_23446,N_23966);
nand U24088 (N_24088,N_23517,N_23854);
nor U24089 (N_24089,N_23542,N_23989);
and U24090 (N_24090,N_23168,N_23385);
and U24091 (N_24091,N_23359,N_23384);
or U24092 (N_24092,N_23943,N_23892);
and U24093 (N_24093,N_23863,N_23466);
or U24094 (N_24094,N_23426,N_23904);
nand U24095 (N_24095,N_23743,N_23227);
or U24096 (N_24096,N_23986,N_23759);
nor U24097 (N_24097,N_23599,N_23981);
nand U24098 (N_24098,N_23199,N_23624);
xnor U24099 (N_24099,N_23415,N_23113);
nor U24100 (N_24100,N_23031,N_23560);
or U24101 (N_24101,N_23925,N_23170);
nor U24102 (N_24102,N_23842,N_23545);
and U24103 (N_24103,N_23009,N_23371);
and U24104 (N_24104,N_23657,N_23976);
nor U24105 (N_24105,N_23522,N_23809);
nor U24106 (N_24106,N_23843,N_23134);
and U24107 (N_24107,N_23194,N_23209);
or U24108 (N_24108,N_23094,N_23115);
nand U24109 (N_24109,N_23334,N_23564);
nand U24110 (N_24110,N_23233,N_23789);
or U24111 (N_24111,N_23310,N_23221);
xnor U24112 (N_24112,N_23070,N_23146);
nand U24113 (N_24113,N_23214,N_23136);
nand U24114 (N_24114,N_23252,N_23814);
nand U24115 (N_24115,N_23447,N_23546);
or U24116 (N_24116,N_23855,N_23258);
nand U24117 (N_24117,N_23344,N_23827);
or U24118 (N_24118,N_23576,N_23399);
nor U24119 (N_24119,N_23660,N_23338);
or U24120 (N_24120,N_23601,N_23915);
xnor U24121 (N_24121,N_23457,N_23430);
xnor U24122 (N_24122,N_23748,N_23617);
nor U24123 (N_24123,N_23933,N_23535);
nor U24124 (N_24124,N_23742,N_23704);
or U24125 (N_24125,N_23416,N_23845);
or U24126 (N_24126,N_23783,N_23222);
or U24127 (N_24127,N_23042,N_23130);
nand U24128 (N_24128,N_23902,N_23548);
nor U24129 (N_24129,N_23592,N_23555);
and U24130 (N_24130,N_23857,N_23261);
nor U24131 (N_24131,N_23353,N_23443);
nor U24132 (N_24132,N_23423,N_23294);
and U24133 (N_24133,N_23931,N_23412);
and U24134 (N_24134,N_23387,N_23341);
nand U24135 (N_24135,N_23037,N_23318);
or U24136 (N_24136,N_23488,N_23534);
or U24137 (N_24137,N_23493,N_23913);
or U24138 (N_24138,N_23474,N_23272);
nor U24139 (N_24139,N_23066,N_23839);
nand U24140 (N_24140,N_23851,N_23309);
xor U24141 (N_24141,N_23292,N_23505);
xor U24142 (N_24142,N_23811,N_23957);
xnor U24143 (N_24143,N_23129,N_23032);
nand U24144 (N_24144,N_23515,N_23425);
xnor U24145 (N_24145,N_23536,N_23469);
or U24146 (N_24146,N_23270,N_23095);
and U24147 (N_24147,N_23566,N_23141);
nor U24148 (N_24148,N_23835,N_23234);
nand U24149 (N_24149,N_23537,N_23354);
or U24150 (N_24150,N_23777,N_23131);
xnor U24151 (N_24151,N_23398,N_23312);
and U24152 (N_24152,N_23228,N_23022);
nand U24153 (N_24153,N_23219,N_23658);
nand U24154 (N_24154,N_23065,N_23816);
xnor U24155 (N_24155,N_23427,N_23080);
xnor U24156 (N_24156,N_23076,N_23268);
and U24157 (N_24157,N_23884,N_23912);
nand U24158 (N_24158,N_23771,N_23967);
nor U24159 (N_24159,N_23602,N_23333);
and U24160 (N_24160,N_23331,N_23383);
xnor U24161 (N_24161,N_23054,N_23167);
or U24162 (N_24162,N_23574,N_23541);
or U24163 (N_24163,N_23400,N_23551);
or U24164 (N_24164,N_23241,N_23732);
and U24165 (N_24165,N_23804,N_23491);
nand U24166 (N_24166,N_23217,N_23340);
nand U24167 (N_24167,N_23264,N_23005);
nand U24168 (N_24168,N_23477,N_23475);
and U24169 (N_24169,N_23802,N_23378);
xnor U24170 (N_24170,N_23569,N_23148);
or U24171 (N_24171,N_23767,N_23490);
nor U24172 (N_24172,N_23367,N_23500);
and U24173 (N_24173,N_23905,N_23317);
or U24174 (N_24174,N_23959,N_23822);
nand U24175 (N_24175,N_23179,N_23775);
nor U24176 (N_24176,N_23396,N_23585);
and U24177 (N_24177,N_23544,N_23960);
nor U24178 (N_24178,N_23610,N_23788);
xnor U24179 (N_24179,N_23663,N_23041);
xnor U24180 (N_24180,N_23785,N_23147);
or U24181 (N_24181,N_23640,N_23000);
and U24182 (N_24182,N_23858,N_23924);
nor U24183 (N_24183,N_23539,N_23275);
or U24184 (N_24184,N_23459,N_23502);
or U24185 (N_24185,N_23248,N_23995);
nor U24186 (N_24186,N_23296,N_23869);
or U24187 (N_24187,N_23067,N_23004);
or U24188 (N_24188,N_23244,N_23947);
and U24189 (N_24189,N_23286,N_23882);
nand U24190 (N_24190,N_23971,N_23514);
and U24191 (N_24191,N_23166,N_23696);
or U24192 (N_24192,N_23265,N_23381);
nor U24193 (N_24193,N_23372,N_23757);
nand U24194 (N_24194,N_23817,N_23030);
xor U24195 (N_24195,N_23313,N_23060);
nand U24196 (N_24196,N_23705,N_23729);
nor U24197 (N_24197,N_23911,N_23240);
xor U24198 (N_24198,N_23928,N_23674);
nand U24199 (N_24199,N_23772,N_23291);
and U24200 (N_24200,N_23435,N_23304);
and U24201 (N_24201,N_23453,N_23665);
xor U24202 (N_24202,N_23008,N_23528);
or U24203 (N_24203,N_23752,N_23583);
or U24204 (N_24204,N_23917,N_23118);
nor U24205 (N_24205,N_23135,N_23812);
xor U24206 (N_24206,N_23343,N_23119);
nand U24207 (N_24207,N_23320,N_23326);
xor U24208 (N_24208,N_23273,N_23028);
or U24209 (N_24209,N_23582,N_23499);
xnor U24210 (N_24210,N_23571,N_23970);
nand U24211 (N_24211,N_23103,N_23053);
or U24212 (N_24212,N_23288,N_23057);
or U24213 (N_24213,N_23106,N_23428);
nor U24214 (N_24214,N_23133,N_23349);
nor U24215 (N_24215,N_23375,N_23991);
xnor U24216 (N_24216,N_23944,N_23158);
and U24217 (N_24217,N_23382,N_23332);
and U24218 (N_24218,N_23468,N_23538);
nand U24219 (N_24219,N_23764,N_23088);
nand U24220 (N_24220,N_23212,N_23232);
xnor U24221 (N_24221,N_23509,N_23082);
and U24222 (N_24222,N_23591,N_23710);
nand U24223 (N_24223,N_23781,N_23521);
and U24224 (N_24224,N_23321,N_23449);
nand U24225 (N_24225,N_23295,N_23737);
xor U24226 (N_24226,N_23977,N_23736);
xnor U24227 (N_24227,N_23051,N_23124);
or U24228 (N_24228,N_23339,N_23128);
and U24229 (N_24229,N_23554,N_23675);
or U24230 (N_24230,N_23671,N_23724);
xnor U24231 (N_24231,N_23531,N_23872);
xor U24232 (N_24232,N_23984,N_23336);
nand U24233 (N_24233,N_23717,N_23877);
and U24234 (N_24234,N_23670,N_23953);
xor U24235 (N_24235,N_23281,N_23983);
or U24236 (N_24236,N_23609,N_23867);
nor U24237 (N_24237,N_23254,N_23039);
and U24238 (N_24238,N_23840,N_23697);
nand U24239 (N_24239,N_23464,N_23012);
and U24240 (N_24240,N_23910,N_23935);
or U24241 (N_24241,N_23586,N_23723);
and U24242 (N_24242,N_23165,N_23603);
or U24243 (N_24243,N_23745,N_23616);
nor U24244 (N_24244,N_23655,N_23418);
or U24245 (N_24245,N_23871,N_23019);
nor U24246 (N_24246,N_23044,N_23629);
nor U24247 (N_24247,N_23888,N_23369);
nand U24248 (N_24248,N_23993,N_23997);
or U24249 (N_24249,N_23486,N_23467);
or U24250 (N_24250,N_23825,N_23803);
nor U24251 (N_24251,N_23392,N_23438);
or U24252 (N_24252,N_23895,N_23394);
and U24253 (N_24253,N_23619,N_23831);
nor U24254 (N_24254,N_23887,N_23138);
and U24255 (N_24255,N_23454,N_23906);
xor U24256 (N_24256,N_23143,N_23596);
xor U24257 (N_24257,N_23210,N_23434);
nor U24258 (N_24258,N_23875,N_23711);
xor U24259 (N_24259,N_23722,N_23361);
xor U24260 (N_24260,N_23140,N_23727);
and U24261 (N_24261,N_23881,N_23155);
nand U24262 (N_24262,N_23828,N_23852);
or U24263 (N_24263,N_23731,N_23325);
nor U24264 (N_24264,N_23186,N_23393);
nand U24265 (N_24265,N_23673,N_23805);
nor U24266 (N_24266,N_23978,N_23519);
xor U24267 (N_24267,N_23225,N_23195);
nand U24268 (N_24268,N_23243,N_23735);
xnor U24269 (N_24269,N_23125,N_23738);
or U24270 (N_24270,N_23216,N_23087);
xor U24271 (N_24271,N_23963,N_23823);
xnor U24272 (N_24272,N_23002,N_23590);
or U24273 (N_24273,N_23589,N_23029);
nor U24274 (N_24274,N_23681,N_23362);
xor U24275 (N_24275,N_23420,N_23914);
nor U24276 (N_24276,N_23496,N_23807);
and U24277 (N_24277,N_23725,N_23149);
nor U24278 (N_24278,N_23980,N_23678);
and U24279 (N_24279,N_23650,N_23250);
xor U24280 (N_24280,N_23639,N_23685);
and U24281 (N_24281,N_23052,N_23284);
nand U24282 (N_24282,N_23187,N_23256);
or U24283 (N_24283,N_23255,N_23813);
or U24284 (N_24284,N_23091,N_23547);
or U24285 (N_24285,N_23390,N_23679);
nand U24286 (N_24286,N_23543,N_23793);
xnor U24287 (N_24287,N_23335,N_23862);
nor U24288 (N_24288,N_23523,N_23719);
xor U24289 (N_24289,N_23267,N_23506);
nor U24290 (N_24290,N_23540,N_23846);
nor U24291 (N_24291,N_23575,N_23102);
or U24292 (N_24292,N_23765,N_23373);
or U24293 (N_24293,N_23922,N_23850);
nor U24294 (N_24294,N_23684,N_23703);
nand U24295 (N_24295,N_23529,N_23756);
xnor U24296 (N_24296,N_23716,N_23162);
and U24297 (N_24297,N_23370,N_23992);
and U24298 (N_24298,N_23886,N_23532);
xnor U24299 (N_24299,N_23072,N_23883);
and U24300 (N_24300,N_23451,N_23614);
or U24301 (N_24301,N_23955,N_23142);
nor U24302 (N_24302,N_23768,N_23680);
nand U24303 (N_24303,N_23643,N_23013);
or U24304 (N_24304,N_23401,N_23494);
and U24305 (N_24305,N_23766,N_23379);
and U24306 (N_24306,N_23458,N_23608);
nand U24307 (N_24307,N_23958,N_23612);
nand U24308 (N_24308,N_23180,N_23441);
or U24309 (N_24309,N_23920,N_23927);
xor U24310 (N_24310,N_23594,N_23123);
or U24311 (N_24311,N_23290,N_23040);
and U24312 (N_24312,N_23093,N_23567);
or U24313 (N_24313,N_23236,N_23127);
xnor U24314 (N_24314,N_23414,N_23263);
nand U24315 (N_24315,N_23649,N_23587);
or U24316 (N_24316,N_23826,N_23190);
and U24317 (N_24317,N_23482,N_23838);
or U24318 (N_24318,N_23623,N_23791);
nor U24319 (N_24319,N_23121,N_23712);
nor U24320 (N_24320,N_23376,N_23189);
and U24321 (N_24321,N_23634,N_23778);
or U24322 (N_24322,N_23593,N_23078);
or U24323 (N_24323,N_23646,N_23213);
nor U24324 (N_24324,N_23820,N_23700);
xnor U24325 (N_24325,N_23666,N_23604);
xnor U24326 (N_24326,N_23016,N_23606);
and U24327 (N_24327,N_23557,N_23699);
xor U24328 (N_24328,N_23205,N_23901);
nor U24329 (N_24329,N_23999,N_23471);
xor U24330 (N_24330,N_23485,N_23157);
or U24331 (N_24331,N_23899,N_23998);
xnor U24332 (N_24332,N_23308,N_23169);
nand U24333 (N_24333,N_23492,N_23689);
or U24334 (N_24334,N_23948,N_23949);
nor U24335 (N_24335,N_23741,N_23686);
nor U24336 (N_24336,N_23562,N_23503);
or U24337 (N_24337,N_23647,N_23316);
nand U24338 (N_24338,N_23739,N_23985);
and U24339 (N_24339,N_23058,N_23861);
and U24340 (N_24340,N_23676,N_23668);
and U24341 (N_24341,N_23790,N_23274);
nor U24342 (N_24342,N_23715,N_23346);
nor U24343 (N_24343,N_23386,N_23628);
and U24344 (N_24344,N_23510,N_23556);
nand U24345 (N_24345,N_23644,N_23025);
and U24346 (N_24346,N_23419,N_23196);
nor U24347 (N_24347,N_23878,N_23465);
nor U24348 (N_24348,N_23132,N_23900);
xnor U24349 (N_24349,N_23533,N_23511);
nor U24350 (N_24350,N_23890,N_23607);
nor U24351 (N_24351,N_23161,N_23356);
nand U24352 (N_24352,N_23348,N_23007);
nand U24353 (N_24353,N_23260,N_23198);
or U24354 (N_24354,N_23111,N_23620);
nand U24355 (N_24355,N_23230,N_23003);
or U24356 (N_24356,N_23301,N_23017);
xnor U24357 (N_24357,N_23968,N_23444);
xor U24358 (N_24358,N_23656,N_23047);
nor U24359 (N_24359,N_23433,N_23174);
and U24360 (N_24360,N_23497,N_23154);
or U24361 (N_24361,N_23758,N_23859);
nand U24362 (N_24362,N_23096,N_23720);
or U24363 (N_24363,N_23830,N_23632);
xnor U24364 (N_24364,N_23856,N_23406);
nand U24365 (N_24365,N_23974,N_23800);
nor U24366 (N_24366,N_23110,N_23470);
nand U24367 (N_24367,N_23622,N_23578);
nand U24368 (N_24368,N_23939,N_23661);
nor U24369 (N_24369,N_23262,N_23249);
nand U24370 (N_24370,N_23972,N_23099);
xnor U24371 (N_24371,N_23324,N_23437);
nor U24372 (N_24372,N_23682,N_23342);
or U24373 (N_24373,N_23432,N_23570);
nand U24374 (N_24374,N_23853,N_23941);
xor U24375 (N_24375,N_23495,N_23033);
nor U24376 (N_24376,N_23048,N_23806);
and U24377 (N_24377,N_23774,N_23014);
nor U24378 (N_24378,N_23081,N_23613);
and U24379 (N_24379,N_23215,N_23786);
and U24380 (N_24380,N_23979,N_23109);
xnor U24381 (N_24381,N_23907,N_23734);
nand U24382 (N_24382,N_23498,N_23733);
nor U24383 (N_24383,N_23694,N_23693);
and U24384 (N_24384,N_23175,N_23821);
nor U24385 (N_24385,N_23450,N_23751);
nand U24386 (N_24386,N_23483,N_23229);
and U24387 (N_24387,N_23345,N_23549);
xnor U24388 (N_24388,N_23084,N_23755);
xor U24389 (N_24389,N_23027,N_23299);
nand U24390 (N_24390,N_23061,N_23937);
and U24391 (N_24391,N_23749,N_23982);
nand U24392 (N_24392,N_23580,N_23368);
nor U24393 (N_24393,N_23360,N_23409);
and U24394 (N_24394,N_23635,N_23908);
nand U24395 (N_24395,N_23391,N_23507);
nand U24396 (N_24396,N_23558,N_23940);
and U24397 (N_24397,N_23389,N_23176);
nand U24398 (N_24398,N_23598,N_23996);
nand U24399 (N_24399,N_23046,N_23584);
or U24400 (N_24400,N_23868,N_23006);
and U24401 (N_24401,N_23231,N_23834);
or U24402 (N_24402,N_23266,N_23481);
and U24403 (N_24403,N_23431,N_23043);
nor U24404 (N_24404,N_23035,N_23377);
or U24405 (N_24405,N_23159,N_23120);
or U24406 (N_24406,N_23351,N_23259);
xnor U24407 (N_24407,N_23615,N_23145);
nor U24408 (N_24408,N_23402,N_23153);
nor U24409 (N_24409,N_23484,N_23642);
xnor U24410 (N_24410,N_23024,N_23473);
xnor U24411 (N_24411,N_23380,N_23879);
xnor U24412 (N_24412,N_23930,N_23698);
and U24413 (N_24413,N_23626,N_23950);
nand U24414 (N_24414,N_23618,N_23595);
nand U24415 (N_24415,N_23726,N_23844);
nand U24416 (N_24416,N_23926,N_23780);
or U24417 (N_24417,N_23085,N_23122);
nor U24418 (N_24418,N_23126,N_23669);
nand U24419 (N_24419,N_23184,N_23253);
and U24420 (N_24420,N_23832,N_23144);
and U24421 (N_24421,N_23568,N_23516);
or U24422 (N_24422,N_23956,N_23337);
nand U24423 (N_24423,N_23762,N_23747);
nand U24424 (N_24424,N_23089,N_23280);
nor U24425 (N_24425,N_23530,N_23573);
or U24426 (N_24426,N_23315,N_23841);
or U24427 (N_24427,N_23307,N_23936);
xor U24428 (N_24428,N_23357,N_23885);
and U24429 (N_24429,N_23695,N_23672);
nor U24430 (N_24430,N_23083,N_23242);
xnor U24431 (N_24431,N_23714,N_23709);
or U24432 (N_24432,N_23440,N_23489);
xnor U24433 (N_24433,N_23572,N_23090);
xor U24434 (N_24434,N_23023,N_23754);
nand U24435 (N_24435,N_23036,N_23919);
and U24436 (N_24436,N_23327,N_23636);
nand U24437 (N_24437,N_23001,N_23794);
xnor U24438 (N_24438,N_23631,N_23311);
nor U24439 (N_24439,N_23824,N_23104);
and U24440 (N_24440,N_23448,N_23056);
xnor U24441 (N_24441,N_23374,N_23880);
xor U24442 (N_24442,N_23350,N_23388);
xnor U24443 (N_24443,N_23760,N_23197);
and U24444 (N_24444,N_23410,N_23487);
nor U24445 (N_24445,N_23364,N_23770);
or U24446 (N_24446,N_23476,N_23563);
or U24447 (N_24447,N_23934,N_23753);
xnor U24448 (N_24448,N_23114,N_23289);
and U24449 (N_24449,N_23208,N_23050);
nor U24450 (N_24450,N_23139,N_23413);
nor U24451 (N_24451,N_23520,N_23352);
or U24452 (N_24452,N_23365,N_23347);
nor U24453 (N_24453,N_23945,N_23026);
and U24454 (N_24454,N_23463,N_23152);
nand U24455 (N_24455,N_23439,N_23182);
or U24456 (N_24456,N_23285,N_23916);
nor U24457 (N_24457,N_23112,N_23193);
nand U24458 (N_24458,N_23277,N_23690);
and U24459 (N_24459,N_23098,N_23172);
nand U24460 (N_24460,N_23298,N_23211);
nand U24461 (N_24461,N_23455,N_23677);
and U24462 (N_24462,N_23889,N_23651);
and U24463 (N_24463,N_23565,N_23201);
or U24464 (N_24464,N_23893,N_23183);
and U24465 (N_24465,N_23397,N_23921);
nand U24466 (N_24466,N_23611,N_23874);
xor U24467 (N_24467,N_23055,N_23245);
and U24468 (N_24468,N_23962,N_23799);
nor U24469 (N_24469,N_23866,N_23200);
or U24470 (N_24470,N_23411,N_23633);
and U24471 (N_24471,N_23086,N_23836);
and U24472 (N_24472,N_23969,N_23630);
or U24473 (N_24473,N_23627,N_23063);
and U24474 (N_24474,N_23269,N_23010);
nand U24475 (N_24475,N_23407,N_23833);
or U24476 (N_24476,N_23761,N_23204);
nor U24477 (N_24477,N_23815,N_23203);
and U24478 (N_24478,N_23795,N_23251);
nor U24479 (N_24479,N_23297,N_23849);
and U24480 (N_24480,N_23306,N_23625);
nand U24481 (N_24481,N_23641,N_23178);
nor U24482 (N_24482,N_23561,N_23929);
nand U24483 (N_24483,N_23728,N_23224);
nor U24484 (N_24484,N_23526,N_23964);
and U24485 (N_24485,N_23951,N_23314);
nor U24486 (N_24486,N_23702,N_23952);
or U24487 (N_24487,N_23073,N_23508);
nand U24488 (N_24488,N_23181,N_23101);
xnor U24489 (N_24489,N_23442,N_23223);
xor U24490 (N_24490,N_23796,N_23769);
nor U24491 (N_24491,N_23818,N_23069);
or U24492 (N_24492,N_23220,N_23870);
nor U24493 (N_24493,N_23107,N_23648);
nor U24494 (N_24494,N_23792,N_23973);
nand U24495 (N_24495,N_23987,N_23638);
or U24496 (N_24496,N_23151,N_23238);
xor U24497 (N_24497,N_23271,N_23527);
and U24498 (N_24498,N_23395,N_23077);
nand U24499 (N_24499,N_23550,N_23079);
or U24500 (N_24500,N_23839,N_23128);
nand U24501 (N_24501,N_23925,N_23958);
xnor U24502 (N_24502,N_23771,N_23144);
xor U24503 (N_24503,N_23949,N_23207);
or U24504 (N_24504,N_23490,N_23435);
xnor U24505 (N_24505,N_23744,N_23262);
nand U24506 (N_24506,N_23165,N_23539);
nor U24507 (N_24507,N_23505,N_23841);
or U24508 (N_24508,N_23774,N_23464);
nor U24509 (N_24509,N_23529,N_23311);
and U24510 (N_24510,N_23156,N_23588);
nand U24511 (N_24511,N_23565,N_23881);
nand U24512 (N_24512,N_23996,N_23929);
nand U24513 (N_24513,N_23643,N_23291);
xnor U24514 (N_24514,N_23166,N_23169);
nor U24515 (N_24515,N_23934,N_23579);
nor U24516 (N_24516,N_23191,N_23396);
and U24517 (N_24517,N_23258,N_23490);
and U24518 (N_24518,N_23380,N_23167);
and U24519 (N_24519,N_23335,N_23076);
and U24520 (N_24520,N_23213,N_23552);
xnor U24521 (N_24521,N_23530,N_23761);
nor U24522 (N_24522,N_23696,N_23612);
nand U24523 (N_24523,N_23005,N_23373);
or U24524 (N_24524,N_23294,N_23386);
nor U24525 (N_24525,N_23179,N_23778);
and U24526 (N_24526,N_23439,N_23113);
nand U24527 (N_24527,N_23452,N_23098);
xor U24528 (N_24528,N_23050,N_23021);
or U24529 (N_24529,N_23826,N_23875);
nor U24530 (N_24530,N_23275,N_23873);
and U24531 (N_24531,N_23514,N_23893);
or U24532 (N_24532,N_23595,N_23730);
nor U24533 (N_24533,N_23971,N_23867);
or U24534 (N_24534,N_23309,N_23520);
xnor U24535 (N_24535,N_23748,N_23891);
or U24536 (N_24536,N_23341,N_23332);
xor U24537 (N_24537,N_23363,N_23850);
xor U24538 (N_24538,N_23794,N_23866);
nor U24539 (N_24539,N_23403,N_23037);
or U24540 (N_24540,N_23434,N_23863);
nand U24541 (N_24541,N_23931,N_23544);
xor U24542 (N_24542,N_23501,N_23120);
or U24543 (N_24543,N_23655,N_23280);
nand U24544 (N_24544,N_23092,N_23861);
or U24545 (N_24545,N_23953,N_23088);
nand U24546 (N_24546,N_23028,N_23607);
and U24547 (N_24547,N_23698,N_23057);
nand U24548 (N_24548,N_23199,N_23939);
xor U24549 (N_24549,N_23019,N_23129);
and U24550 (N_24550,N_23119,N_23583);
nand U24551 (N_24551,N_23615,N_23620);
nor U24552 (N_24552,N_23448,N_23682);
or U24553 (N_24553,N_23611,N_23663);
or U24554 (N_24554,N_23009,N_23253);
and U24555 (N_24555,N_23833,N_23278);
nand U24556 (N_24556,N_23608,N_23015);
or U24557 (N_24557,N_23430,N_23547);
and U24558 (N_24558,N_23444,N_23290);
nand U24559 (N_24559,N_23291,N_23900);
nor U24560 (N_24560,N_23162,N_23387);
nand U24561 (N_24561,N_23464,N_23982);
xnor U24562 (N_24562,N_23729,N_23451);
or U24563 (N_24563,N_23746,N_23340);
or U24564 (N_24564,N_23542,N_23555);
nor U24565 (N_24565,N_23398,N_23132);
nand U24566 (N_24566,N_23960,N_23639);
xor U24567 (N_24567,N_23814,N_23226);
or U24568 (N_24568,N_23962,N_23886);
nand U24569 (N_24569,N_23661,N_23297);
and U24570 (N_24570,N_23065,N_23797);
or U24571 (N_24571,N_23744,N_23201);
and U24572 (N_24572,N_23536,N_23859);
nand U24573 (N_24573,N_23461,N_23078);
and U24574 (N_24574,N_23881,N_23709);
and U24575 (N_24575,N_23783,N_23777);
or U24576 (N_24576,N_23447,N_23019);
nor U24577 (N_24577,N_23138,N_23190);
and U24578 (N_24578,N_23112,N_23870);
and U24579 (N_24579,N_23059,N_23046);
or U24580 (N_24580,N_23849,N_23782);
nand U24581 (N_24581,N_23923,N_23975);
and U24582 (N_24582,N_23250,N_23115);
and U24583 (N_24583,N_23360,N_23567);
and U24584 (N_24584,N_23087,N_23487);
nand U24585 (N_24585,N_23203,N_23373);
and U24586 (N_24586,N_23011,N_23744);
xor U24587 (N_24587,N_23221,N_23645);
nand U24588 (N_24588,N_23357,N_23851);
xor U24589 (N_24589,N_23793,N_23952);
or U24590 (N_24590,N_23451,N_23746);
or U24591 (N_24591,N_23009,N_23701);
nand U24592 (N_24592,N_23604,N_23539);
xnor U24593 (N_24593,N_23526,N_23535);
xnor U24594 (N_24594,N_23735,N_23132);
xor U24595 (N_24595,N_23235,N_23509);
xor U24596 (N_24596,N_23176,N_23781);
or U24597 (N_24597,N_23547,N_23788);
xnor U24598 (N_24598,N_23378,N_23883);
and U24599 (N_24599,N_23625,N_23616);
nand U24600 (N_24600,N_23633,N_23817);
and U24601 (N_24601,N_23120,N_23781);
and U24602 (N_24602,N_23422,N_23535);
xor U24603 (N_24603,N_23987,N_23424);
nor U24604 (N_24604,N_23694,N_23259);
and U24605 (N_24605,N_23450,N_23108);
xnor U24606 (N_24606,N_23442,N_23936);
nand U24607 (N_24607,N_23407,N_23487);
and U24608 (N_24608,N_23789,N_23321);
xor U24609 (N_24609,N_23118,N_23704);
nor U24610 (N_24610,N_23499,N_23104);
and U24611 (N_24611,N_23141,N_23023);
nor U24612 (N_24612,N_23863,N_23138);
and U24613 (N_24613,N_23776,N_23623);
nor U24614 (N_24614,N_23198,N_23314);
nand U24615 (N_24615,N_23736,N_23557);
or U24616 (N_24616,N_23888,N_23225);
and U24617 (N_24617,N_23059,N_23278);
nand U24618 (N_24618,N_23233,N_23699);
nand U24619 (N_24619,N_23060,N_23721);
and U24620 (N_24620,N_23451,N_23970);
xnor U24621 (N_24621,N_23053,N_23537);
xor U24622 (N_24622,N_23648,N_23993);
and U24623 (N_24623,N_23773,N_23606);
nor U24624 (N_24624,N_23898,N_23319);
or U24625 (N_24625,N_23699,N_23556);
nand U24626 (N_24626,N_23800,N_23134);
or U24627 (N_24627,N_23311,N_23445);
xor U24628 (N_24628,N_23360,N_23267);
xor U24629 (N_24629,N_23183,N_23400);
xor U24630 (N_24630,N_23289,N_23635);
and U24631 (N_24631,N_23681,N_23764);
nor U24632 (N_24632,N_23493,N_23827);
xor U24633 (N_24633,N_23346,N_23102);
nor U24634 (N_24634,N_23908,N_23751);
nand U24635 (N_24635,N_23025,N_23867);
and U24636 (N_24636,N_23835,N_23542);
and U24637 (N_24637,N_23969,N_23823);
and U24638 (N_24638,N_23287,N_23505);
or U24639 (N_24639,N_23740,N_23714);
nand U24640 (N_24640,N_23033,N_23806);
xnor U24641 (N_24641,N_23773,N_23673);
nor U24642 (N_24642,N_23653,N_23108);
xor U24643 (N_24643,N_23282,N_23745);
or U24644 (N_24644,N_23480,N_23219);
nand U24645 (N_24645,N_23526,N_23722);
nand U24646 (N_24646,N_23881,N_23808);
xnor U24647 (N_24647,N_23734,N_23832);
nand U24648 (N_24648,N_23987,N_23890);
nor U24649 (N_24649,N_23990,N_23399);
and U24650 (N_24650,N_23169,N_23593);
and U24651 (N_24651,N_23687,N_23673);
nand U24652 (N_24652,N_23970,N_23173);
and U24653 (N_24653,N_23414,N_23131);
xor U24654 (N_24654,N_23486,N_23758);
nand U24655 (N_24655,N_23466,N_23502);
nor U24656 (N_24656,N_23805,N_23210);
nand U24657 (N_24657,N_23964,N_23120);
and U24658 (N_24658,N_23255,N_23235);
and U24659 (N_24659,N_23969,N_23900);
or U24660 (N_24660,N_23322,N_23123);
nor U24661 (N_24661,N_23524,N_23850);
xor U24662 (N_24662,N_23248,N_23976);
or U24663 (N_24663,N_23343,N_23175);
xor U24664 (N_24664,N_23786,N_23261);
and U24665 (N_24665,N_23083,N_23757);
nor U24666 (N_24666,N_23759,N_23065);
xor U24667 (N_24667,N_23975,N_23711);
and U24668 (N_24668,N_23800,N_23879);
or U24669 (N_24669,N_23239,N_23493);
nor U24670 (N_24670,N_23500,N_23967);
xnor U24671 (N_24671,N_23563,N_23379);
or U24672 (N_24672,N_23416,N_23660);
xor U24673 (N_24673,N_23553,N_23947);
nand U24674 (N_24674,N_23463,N_23265);
nand U24675 (N_24675,N_23069,N_23889);
or U24676 (N_24676,N_23781,N_23893);
and U24677 (N_24677,N_23454,N_23246);
nand U24678 (N_24678,N_23086,N_23960);
xnor U24679 (N_24679,N_23099,N_23208);
nor U24680 (N_24680,N_23992,N_23494);
and U24681 (N_24681,N_23175,N_23878);
and U24682 (N_24682,N_23421,N_23264);
nand U24683 (N_24683,N_23970,N_23107);
and U24684 (N_24684,N_23591,N_23845);
or U24685 (N_24685,N_23717,N_23895);
nand U24686 (N_24686,N_23403,N_23133);
nand U24687 (N_24687,N_23385,N_23346);
nor U24688 (N_24688,N_23336,N_23472);
nor U24689 (N_24689,N_23595,N_23914);
xnor U24690 (N_24690,N_23795,N_23423);
and U24691 (N_24691,N_23259,N_23751);
nand U24692 (N_24692,N_23648,N_23409);
nor U24693 (N_24693,N_23969,N_23766);
nand U24694 (N_24694,N_23080,N_23356);
xnor U24695 (N_24695,N_23742,N_23229);
and U24696 (N_24696,N_23954,N_23181);
or U24697 (N_24697,N_23475,N_23493);
xor U24698 (N_24698,N_23511,N_23318);
and U24699 (N_24699,N_23345,N_23693);
or U24700 (N_24700,N_23409,N_23547);
xnor U24701 (N_24701,N_23911,N_23626);
nor U24702 (N_24702,N_23650,N_23135);
xor U24703 (N_24703,N_23581,N_23337);
nor U24704 (N_24704,N_23735,N_23860);
and U24705 (N_24705,N_23203,N_23127);
nor U24706 (N_24706,N_23882,N_23208);
or U24707 (N_24707,N_23193,N_23480);
and U24708 (N_24708,N_23834,N_23254);
nand U24709 (N_24709,N_23623,N_23278);
or U24710 (N_24710,N_23948,N_23362);
xor U24711 (N_24711,N_23929,N_23491);
nand U24712 (N_24712,N_23960,N_23489);
and U24713 (N_24713,N_23571,N_23666);
xnor U24714 (N_24714,N_23582,N_23389);
xnor U24715 (N_24715,N_23466,N_23013);
nor U24716 (N_24716,N_23787,N_23393);
xnor U24717 (N_24717,N_23335,N_23837);
nand U24718 (N_24718,N_23192,N_23432);
nand U24719 (N_24719,N_23166,N_23290);
and U24720 (N_24720,N_23627,N_23820);
xnor U24721 (N_24721,N_23897,N_23392);
and U24722 (N_24722,N_23792,N_23984);
nand U24723 (N_24723,N_23849,N_23982);
nor U24724 (N_24724,N_23833,N_23100);
or U24725 (N_24725,N_23645,N_23303);
and U24726 (N_24726,N_23644,N_23018);
xnor U24727 (N_24727,N_23844,N_23567);
xor U24728 (N_24728,N_23235,N_23117);
nand U24729 (N_24729,N_23275,N_23795);
and U24730 (N_24730,N_23058,N_23845);
and U24731 (N_24731,N_23495,N_23065);
or U24732 (N_24732,N_23562,N_23852);
and U24733 (N_24733,N_23933,N_23229);
or U24734 (N_24734,N_23851,N_23227);
xor U24735 (N_24735,N_23683,N_23449);
xnor U24736 (N_24736,N_23068,N_23474);
or U24737 (N_24737,N_23514,N_23858);
and U24738 (N_24738,N_23603,N_23881);
and U24739 (N_24739,N_23019,N_23990);
nor U24740 (N_24740,N_23071,N_23203);
xor U24741 (N_24741,N_23214,N_23636);
or U24742 (N_24742,N_23622,N_23071);
xor U24743 (N_24743,N_23943,N_23019);
and U24744 (N_24744,N_23255,N_23849);
nor U24745 (N_24745,N_23233,N_23531);
nand U24746 (N_24746,N_23626,N_23293);
and U24747 (N_24747,N_23761,N_23297);
nand U24748 (N_24748,N_23227,N_23582);
nand U24749 (N_24749,N_23819,N_23883);
nand U24750 (N_24750,N_23154,N_23554);
xnor U24751 (N_24751,N_23209,N_23596);
and U24752 (N_24752,N_23844,N_23392);
nor U24753 (N_24753,N_23272,N_23319);
and U24754 (N_24754,N_23960,N_23574);
nor U24755 (N_24755,N_23385,N_23642);
xnor U24756 (N_24756,N_23498,N_23776);
xor U24757 (N_24757,N_23374,N_23007);
nand U24758 (N_24758,N_23163,N_23226);
nand U24759 (N_24759,N_23720,N_23186);
and U24760 (N_24760,N_23892,N_23357);
nor U24761 (N_24761,N_23044,N_23967);
xnor U24762 (N_24762,N_23826,N_23709);
nand U24763 (N_24763,N_23755,N_23302);
xor U24764 (N_24764,N_23424,N_23348);
nand U24765 (N_24765,N_23000,N_23597);
xnor U24766 (N_24766,N_23037,N_23366);
nor U24767 (N_24767,N_23718,N_23264);
or U24768 (N_24768,N_23060,N_23137);
nor U24769 (N_24769,N_23325,N_23740);
nand U24770 (N_24770,N_23819,N_23115);
nand U24771 (N_24771,N_23098,N_23844);
nor U24772 (N_24772,N_23969,N_23469);
nand U24773 (N_24773,N_23043,N_23949);
xor U24774 (N_24774,N_23806,N_23152);
nor U24775 (N_24775,N_23839,N_23453);
nor U24776 (N_24776,N_23969,N_23887);
nor U24777 (N_24777,N_23329,N_23604);
nor U24778 (N_24778,N_23368,N_23287);
and U24779 (N_24779,N_23129,N_23961);
and U24780 (N_24780,N_23131,N_23434);
nor U24781 (N_24781,N_23742,N_23036);
or U24782 (N_24782,N_23023,N_23276);
or U24783 (N_24783,N_23361,N_23488);
xor U24784 (N_24784,N_23494,N_23029);
or U24785 (N_24785,N_23517,N_23354);
nand U24786 (N_24786,N_23970,N_23139);
and U24787 (N_24787,N_23625,N_23733);
nor U24788 (N_24788,N_23387,N_23142);
nor U24789 (N_24789,N_23948,N_23912);
or U24790 (N_24790,N_23708,N_23535);
or U24791 (N_24791,N_23110,N_23973);
nor U24792 (N_24792,N_23510,N_23523);
and U24793 (N_24793,N_23938,N_23388);
nor U24794 (N_24794,N_23434,N_23935);
and U24795 (N_24795,N_23148,N_23380);
and U24796 (N_24796,N_23718,N_23143);
or U24797 (N_24797,N_23724,N_23142);
nand U24798 (N_24798,N_23894,N_23754);
and U24799 (N_24799,N_23916,N_23680);
xnor U24800 (N_24800,N_23195,N_23790);
or U24801 (N_24801,N_23630,N_23265);
xnor U24802 (N_24802,N_23184,N_23753);
or U24803 (N_24803,N_23125,N_23498);
and U24804 (N_24804,N_23201,N_23824);
nor U24805 (N_24805,N_23983,N_23145);
or U24806 (N_24806,N_23159,N_23371);
or U24807 (N_24807,N_23681,N_23380);
nand U24808 (N_24808,N_23014,N_23284);
xnor U24809 (N_24809,N_23768,N_23607);
and U24810 (N_24810,N_23844,N_23635);
or U24811 (N_24811,N_23004,N_23684);
and U24812 (N_24812,N_23706,N_23640);
nand U24813 (N_24813,N_23540,N_23861);
nand U24814 (N_24814,N_23650,N_23484);
and U24815 (N_24815,N_23221,N_23053);
xnor U24816 (N_24816,N_23352,N_23047);
and U24817 (N_24817,N_23089,N_23596);
and U24818 (N_24818,N_23751,N_23962);
and U24819 (N_24819,N_23994,N_23297);
and U24820 (N_24820,N_23205,N_23014);
and U24821 (N_24821,N_23939,N_23937);
or U24822 (N_24822,N_23111,N_23955);
xnor U24823 (N_24823,N_23274,N_23249);
or U24824 (N_24824,N_23710,N_23357);
and U24825 (N_24825,N_23056,N_23794);
and U24826 (N_24826,N_23413,N_23204);
and U24827 (N_24827,N_23821,N_23833);
and U24828 (N_24828,N_23214,N_23278);
nor U24829 (N_24829,N_23765,N_23361);
nor U24830 (N_24830,N_23279,N_23160);
or U24831 (N_24831,N_23110,N_23258);
or U24832 (N_24832,N_23288,N_23654);
nor U24833 (N_24833,N_23599,N_23998);
and U24834 (N_24834,N_23458,N_23586);
nor U24835 (N_24835,N_23154,N_23080);
xor U24836 (N_24836,N_23842,N_23541);
and U24837 (N_24837,N_23544,N_23809);
and U24838 (N_24838,N_23497,N_23816);
xnor U24839 (N_24839,N_23888,N_23073);
xor U24840 (N_24840,N_23069,N_23718);
and U24841 (N_24841,N_23281,N_23192);
or U24842 (N_24842,N_23926,N_23773);
xnor U24843 (N_24843,N_23723,N_23595);
xnor U24844 (N_24844,N_23562,N_23242);
and U24845 (N_24845,N_23237,N_23776);
xnor U24846 (N_24846,N_23837,N_23127);
xnor U24847 (N_24847,N_23993,N_23139);
xor U24848 (N_24848,N_23182,N_23228);
nor U24849 (N_24849,N_23758,N_23029);
nor U24850 (N_24850,N_23074,N_23906);
nand U24851 (N_24851,N_23932,N_23448);
nor U24852 (N_24852,N_23508,N_23119);
nor U24853 (N_24853,N_23939,N_23029);
nor U24854 (N_24854,N_23045,N_23270);
or U24855 (N_24855,N_23498,N_23079);
xor U24856 (N_24856,N_23349,N_23842);
xor U24857 (N_24857,N_23490,N_23198);
and U24858 (N_24858,N_23605,N_23448);
nor U24859 (N_24859,N_23663,N_23568);
xnor U24860 (N_24860,N_23154,N_23294);
nand U24861 (N_24861,N_23495,N_23688);
nor U24862 (N_24862,N_23545,N_23197);
or U24863 (N_24863,N_23705,N_23894);
and U24864 (N_24864,N_23897,N_23158);
or U24865 (N_24865,N_23581,N_23531);
and U24866 (N_24866,N_23324,N_23660);
nor U24867 (N_24867,N_23373,N_23485);
nand U24868 (N_24868,N_23722,N_23808);
nor U24869 (N_24869,N_23212,N_23957);
nand U24870 (N_24870,N_23526,N_23659);
nor U24871 (N_24871,N_23100,N_23682);
nand U24872 (N_24872,N_23768,N_23666);
nor U24873 (N_24873,N_23518,N_23246);
or U24874 (N_24874,N_23669,N_23493);
nand U24875 (N_24875,N_23419,N_23594);
and U24876 (N_24876,N_23946,N_23211);
or U24877 (N_24877,N_23423,N_23719);
xor U24878 (N_24878,N_23126,N_23529);
and U24879 (N_24879,N_23025,N_23258);
nand U24880 (N_24880,N_23221,N_23231);
nand U24881 (N_24881,N_23417,N_23518);
nand U24882 (N_24882,N_23091,N_23172);
nor U24883 (N_24883,N_23803,N_23760);
xnor U24884 (N_24884,N_23967,N_23486);
nand U24885 (N_24885,N_23231,N_23909);
nor U24886 (N_24886,N_23318,N_23708);
nand U24887 (N_24887,N_23034,N_23446);
xnor U24888 (N_24888,N_23251,N_23543);
xnor U24889 (N_24889,N_23069,N_23241);
and U24890 (N_24890,N_23686,N_23316);
or U24891 (N_24891,N_23642,N_23997);
xor U24892 (N_24892,N_23233,N_23287);
and U24893 (N_24893,N_23913,N_23109);
xor U24894 (N_24894,N_23040,N_23957);
nand U24895 (N_24895,N_23731,N_23737);
nor U24896 (N_24896,N_23586,N_23211);
xnor U24897 (N_24897,N_23376,N_23775);
and U24898 (N_24898,N_23948,N_23636);
or U24899 (N_24899,N_23126,N_23524);
nand U24900 (N_24900,N_23571,N_23901);
nand U24901 (N_24901,N_23418,N_23952);
and U24902 (N_24902,N_23388,N_23023);
or U24903 (N_24903,N_23786,N_23961);
nor U24904 (N_24904,N_23341,N_23486);
xnor U24905 (N_24905,N_23837,N_23862);
nor U24906 (N_24906,N_23468,N_23063);
xnor U24907 (N_24907,N_23767,N_23780);
or U24908 (N_24908,N_23229,N_23762);
xor U24909 (N_24909,N_23171,N_23230);
and U24910 (N_24910,N_23668,N_23678);
nand U24911 (N_24911,N_23477,N_23515);
or U24912 (N_24912,N_23600,N_23156);
xor U24913 (N_24913,N_23790,N_23836);
xor U24914 (N_24914,N_23102,N_23300);
and U24915 (N_24915,N_23948,N_23495);
nor U24916 (N_24916,N_23588,N_23183);
nand U24917 (N_24917,N_23405,N_23074);
nand U24918 (N_24918,N_23535,N_23625);
or U24919 (N_24919,N_23090,N_23759);
nand U24920 (N_24920,N_23221,N_23235);
nor U24921 (N_24921,N_23060,N_23612);
and U24922 (N_24922,N_23408,N_23869);
xnor U24923 (N_24923,N_23880,N_23355);
and U24924 (N_24924,N_23920,N_23803);
and U24925 (N_24925,N_23839,N_23682);
xor U24926 (N_24926,N_23044,N_23595);
nand U24927 (N_24927,N_23668,N_23357);
nor U24928 (N_24928,N_23671,N_23397);
or U24929 (N_24929,N_23945,N_23054);
or U24930 (N_24930,N_23004,N_23476);
nand U24931 (N_24931,N_23810,N_23756);
xnor U24932 (N_24932,N_23187,N_23536);
or U24933 (N_24933,N_23776,N_23200);
nand U24934 (N_24934,N_23184,N_23982);
nand U24935 (N_24935,N_23686,N_23708);
or U24936 (N_24936,N_23578,N_23302);
and U24937 (N_24937,N_23899,N_23190);
nand U24938 (N_24938,N_23686,N_23607);
and U24939 (N_24939,N_23139,N_23090);
or U24940 (N_24940,N_23441,N_23101);
or U24941 (N_24941,N_23593,N_23544);
and U24942 (N_24942,N_23194,N_23258);
and U24943 (N_24943,N_23059,N_23657);
nor U24944 (N_24944,N_23605,N_23299);
and U24945 (N_24945,N_23005,N_23191);
nor U24946 (N_24946,N_23253,N_23811);
nor U24947 (N_24947,N_23299,N_23026);
or U24948 (N_24948,N_23449,N_23110);
or U24949 (N_24949,N_23053,N_23363);
nor U24950 (N_24950,N_23640,N_23939);
nor U24951 (N_24951,N_23016,N_23446);
and U24952 (N_24952,N_23205,N_23589);
nor U24953 (N_24953,N_23853,N_23498);
nor U24954 (N_24954,N_23969,N_23680);
nor U24955 (N_24955,N_23492,N_23312);
nor U24956 (N_24956,N_23850,N_23068);
nand U24957 (N_24957,N_23059,N_23967);
nor U24958 (N_24958,N_23077,N_23219);
xor U24959 (N_24959,N_23157,N_23903);
nor U24960 (N_24960,N_23026,N_23855);
and U24961 (N_24961,N_23923,N_23962);
xor U24962 (N_24962,N_23002,N_23935);
nand U24963 (N_24963,N_23068,N_23307);
nand U24964 (N_24964,N_23805,N_23348);
nand U24965 (N_24965,N_23215,N_23659);
and U24966 (N_24966,N_23369,N_23097);
nand U24967 (N_24967,N_23749,N_23958);
nor U24968 (N_24968,N_23212,N_23306);
and U24969 (N_24969,N_23883,N_23131);
or U24970 (N_24970,N_23485,N_23502);
xor U24971 (N_24971,N_23680,N_23862);
nand U24972 (N_24972,N_23265,N_23840);
or U24973 (N_24973,N_23831,N_23295);
nor U24974 (N_24974,N_23128,N_23930);
or U24975 (N_24975,N_23397,N_23611);
and U24976 (N_24976,N_23758,N_23440);
nor U24977 (N_24977,N_23909,N_23304);
or U24978 (N_24978,N_23700,N_23718);
nand U24979 (N_24979,N_23041,N_23686);
xnor U24980 (N_24980,N_23977,N_23825);
or U24981 (N_24981,N_23638,N_23664);
or U24982 (N_24982,N_23567,N_23939);
nor U24983 (N_24983,N_23636,N_23404);
and U24984 (N_24984,N_23363,N_23655);
nor U24985 (N_24985,N_23931,N_23071);
nor U24986 (N_24986,N_23202,N_23975);
nor U24987 (N_24987,N_23317,N_23275);
xor U24988 (N_24988,N_23452,N_23976);
or U24989 (N_24989,N_23922,N_23209);
nor U24990 (N_24990,N_23085,N_23713);
or U24991 (N_24991,N_23307,N_23540);
and U24992 (N_24992,N_23701,N_23233);
nand U24993 (N_24993,N_23422,N_23540);
xor U24994 (N_24994,N_23585,N_23419);
nand U24995 (N_24995,N_23469,N_23324);
or U24996 (N_24996,N_23466,N_23077);
or U24997 (N_24997,N_23099,N_23567);
xor U24998 (N_24998,N_23414,N_23776);
xor U24999 (N_24999,N_23226,N_23706);
or U25000 (N_25000,N_24495,N_24230);
or U25001 (N_25001,N_24265,N_24754);
xnor U25002 (N_25002,N_24090,N_24907);
xnor U25003 (N_25003,N_24177,N_24087);
or U25004 (N_25004,N_24527,N_24570);
and U25005 (N_25005,N_24212,N_24328);
xnor U25006 (N_25006,N_24530,N_24523);
nand U25007 (N_25007,N_24613,N_24716);
nand U25008 (N_25008,N_24232,N_24884);
nor U25009 (N_25009,N_24057,N_24650);
nand U25010 (N_25010,N_24713,N_24569);
xor U25011 (N_25011,N_24467,N_24364);
nand U25012 (N_25012,N_24120,N_24429);
nand U25013 (N_25013,N_24701,N_24099);
xnor U25014 (N_25014,N_24235,N_24741);
nor U25015 (N_25015,N_24266,N_24590);
and U25016 (N_25016,N_24589,N_24399);
nor U25017 (N_25017,N_24392,N_24359);
or U25018 (N_25018,N_24791,N_24211);
nor U25019 (N_25019,N_24019,N_24047);
or U25020 (N_25020,N_24167,N_24101);
nor U25021 (N_25021,N_24353,N_24053);
xnor U25022 (N_25022,N_24144,N_24281);
nor U25023 (N_25023,N_24011,N_24448);
xnor U25024 (N_25024,N_24318,N_24420);
nor U25025 (N_25025,N_24348,N_24288);
or U25026 (N_25026,N_24383,N_24479);
nor U25027 (N_25027,N_24185,N_24830);
nand U25028 (N_25028,N_24943,N_24885);
or U25029 (N_25029,N_24588,N_24894);
or U25030 (N_25030,N_24749,N_24492);
and U25031 (N_25031,N_24093,N_24654);
nor U25032 (N_25032,N_24639,N_24610);
xor U25033 (N_25033,N_24108,N_24055);
and U25034 (N_25034,N_24842,N_24450);
nor U25035 (N_25035,N_24476,N_24107);
or U25036 (N_25036,N_24059,N_24028);
and U25037 (N_25037,N_24603,N_24234);
xnor U25038 (N_25038,N_24665,N_24637);
xnor U25039 (N_25039,N_24256,N_24298);
nor U25040 (N_25040,N_24465,N_24784);
nand U25041 (N_25041,N_24435,N_24483);
xor U25042 (N_25042,N_24086,N_24748);
or U25043 (N_25043,N_24294,N_24634);
xnor U25044 (N_25044,N_24797,N_24506);
nor U25045 (N_25045,N_24829,N_24195);
xnor U25046 (N_25046,N_24264,N_24568);
or U25047 (N_25047,N_24729,N_24471);
xor U25048 (N_25048,N_24083,N_24586);
or U25049 (N_25049,N_24719,N_24157);
and U25050 (N_25050,N_24076,N_24947);
or U25051 (N_25051,N_24773,N_24389);
nor U25052 (N_25052,N_24272,N_24980);
or U25053 (N_25053,N_24540,N_24934);
or U25054 (N_25054,N_24463,N_24440);
and U25055 (N_25055,N_24605,N_24519);
nand U25056 (N_25056,N_24507,N_24788);
or U25057 (N_25057,N_24812,N_24106);
or U25058 (N_25058,N_24329,N_24037);
nor U25059 (N_25059,N_24398,N_24814);
nand U25060 (N_25060,N_24950,N_24869);
and U25061 (N_25061,N_24684,N_24405);
nand U25062 (N_25062,N_24453,N_24113);
xnor U25063 (N_25063,N_24501,N_24370);
nor U25064 (N_25064,N_24189,N_24133);
xor U25065 (N_25065,N_24706,N_24341);
xnor U25066 (N_25066,N_24160,N_24388);
nand U25067 (N_25067,N_24813,N_24752);
nand U25068 (N_25068,N_24430,N_24614);
and U25069 (N_25069,N_24960,N_24514);
xnor U25070 (N_25070,N_24488,N_24198);
xor U25071 (N_25071,N_24895,N_24269);
nand U25072 (N_25072,N_24132,N_24216);
and U25073 (N_25073,N_24284,N_24493);
nor U25074 (N_25074,N_24686,N_24599);
xor U25075 (N_25075,N_24871,N_24222);
xor U25076 (N_25076,N_24914,N_24640);
and U25077 (N_25077,N_24844,N_24792);
and U25078 (N_25078,N_24623,N_24202);
or U25079 (N_25079,N_24809,N_24764);
or U25080 (N_25080,N_24832,N_24699);
nor U25081 (N_25081,N_24877,N_24626);
nor U25082 (N_25082,N_24659,N_24508);
nor U25083 (N_25083,N_24477,N_24025);
xor U25084 (N_25084,N_24485,N_24441);
and U25085 (N_25085,N_24197,N_24986);
or U25086 (N_25086,N_24546,N_24282);
nor U25087 (N_25087,N_24557,N_24179);
or U25088 (N_25088,N_24491,N_24336);
nor U25089 (N_25089,N_24065,N_24021);
and U25090 (N_25090,N_24816,N_24163);
nand U25091 (N_25091,N_24733,N_24368);
xor U25092 (N_25092,N_24852,N_24662);
nand U25093 (N_25093,N_24742,N_24793);
nor U25094 (N_25094,N_24680,N_24082);
and U25095 (N_25095,N_24854,N_24154);
xnor U25096 (N_25096,N_24751,N_24574);
and U25097 (N_25097,N_24757,N_24989);
nand U25098 (N_25098,N_24903,N_24690);
nand U25099 (N_25099,N_24602,N_24461);
nor U25100 (N_25100,N_24660,N_24984);
nand U25101 (N_25101,N_24587,N_24941);
and U25102 (N_25102,N_24343,N_24924);
xor U25103 (N_25103,N_24990,N_24290);
and U25104 (N_25104,N_24831,N_24124);
or U25105 (N_25105,N_24102,N_24513);
and U25106 (N_25106,N_24755,N_24425);
nor U25107 (N_25107,N_24002,N_24456);
and U25108 (N_25108,N_24436,N_24434);
or U25109 (N_25109,N_24088,N_24423);
and U25110 (N_25110,N_24270,N_24421);
or U25111 (N_25111,N_24330,N_24607);
xor U25112 (N_25112,N_24029,N_24581);
nor U25113 (N_25113,N_24332,N_24882);
nand U25114 (N_25114,N_24072,N_24302);
nor U25115 (N_25115,N_24118,N_24122);
nand U25116 (N_25116,N_24126,N_24847);
xnor U25117 (N_25117,N_24003,N_24502);
and U25118 (N_25118,N_24473,N_24172);
nand U25119 (N_25119,N_24666,N_24181);
or U25120 (N_25120,N_24223,N_24097);
nor U25121 (N_25121,N_24412,N_24503);
xnor U25122 (N_25122,N_24168,N_24394);
and U25123 (N_25123,N_24679,N_24825);
nand U25124 (N_25124,N_24201,N_24112);
nor U25125 (N_25125,N_24048,N_24904);
nor U25126 (N_25126,N_24677,N_24678);
and U25127 (N_25127,N_24459,N_24732);
nor U25128 (N_25128,N_24942,N_24015);
or U25129 (N_25129,N_24247,N_24656);
nand U25130 (N_25130,N_24182,N_24811);
nor U25131 (N_25131,N_24860,N_24210);
nor U25132 (N_25132,N_24580,N_24549);
nand U25133 (N_25133,N_24948,N_24458);
or U25134 (N_25134,N_24965,N_24200);
xnor U25135 (N_25135,N_24305,N_24886);
nand U25136 (N_25136,N_24609,N_24049);
or U25137 (N_25137,N_24881,N_24236);
nand U25138 (N_25138,N_24078,N_24416);
nand U25139 (N_25139,N_24379,N_24770);
or U25140 (N_25140,N_24422,N_24710);
or U25141 (N_25141,N_24846,N_24820);
nand U25142 (N_25142,N_24096,N_24967);
nand U25143 (N_25143,N_24912,N_24129);
and U25144 (N_25144,N_24567,N_24455);
xnor U25145 (N_25145,N_24808,N_24462);
nand U25146 (N_25146,N_24487,N_24839);
and U25147 (N_25147,N_24556,N_24897);
nor U25148 (N_25148,N_24277,N_24511);
nor U25149 (N_25149,N_24311,N_24248);
nor U25150 (N_25150,N_24199,N_24066);
nand U25151 (N_25151,N_24104,N_24873);
nand U25152 (N_25152,N_24880,N_24105);
and U25153 (N_25153,N_24286,N_24073);
xnor U25154 (N_25154,N_24632,N_24402);
and U25155 (N_25155,N_24625,N_24718);
xor U25156 (N_25156,N_24123,N_24743);
nor U25157 (N_25157,N_24531,N_24464);
and U25158 (N_25158,N_24692,N_24522);
and U25159 (N_25159,N_24396,N_24601);
nor U25160 (N_25160,N_24356,N_24628);
xor U25161 (N_25161,N_24447,N_24085);
xnor U25162 (N_25162,N_24469,N_24111);
xnor U25163 (N_25163,N_24619,N_24382);
nand U25164 (N_25164,N_24786,N_24648);
nand U25165 (N_25165,N_24801,N_24481);
nor U25166 (N_25166,N_24314,N_24803);
nor U25167 (N_25167,N_24584,N_24593);
and U25168 (N_25168,N_24631,N_24417);
or U25169 (N_25169,N_24604,N_24572);
xnor U25170 (N_25170,N_24283,N_24357);
nand U25171 (N_25171,N_24176,N_24013);
xor U25172 (N_25172,N_24034,N_24611);
xnor U25173 (N_25173,N_24320,N_24923);
nor U25174 (N_25174,N_24896,N_24415);
and U25175 (N_25175,N_24433,N_24951);
nand U25176 (N_25176,N_24616,N_24432);
nand U25177 (N_25177,N_24276,N_24213);
nor U25178 (N_25178,N_24615,N_24279);
xnor U25179 (N_25179,N_24386,N_24375);
and U25180 (N_25180,N_24804,N_24252);
xor U25181 (N_25181,N_24915,N_24390);
xor U25182 (N_25182,N_24064,N_24703);
and U25183 (N_25183,N_24007,N_24977);
nor U25184 (N_25184,N_24532,N_24358);
nand U25185 (N_25185,N_24309,N_24633);
nor U25186 (N_25186,N_24795,N_24856);
xor U25187 (N_25187,N_24419,N_24018);
and U25188 (N_25188,N_24670,N_24683);
or U25189 (N_25189,N_24413,N_24303);
and U25190 (N_25190,N_24494,N_24169);
or U25191 (N_25191,N_24945,N_24334);
xnor U25192 (N_25192,N_24141,N_24164);
xor U25193 (N_25193,N_24414,N_24009);
or U25194 (N_25194,N_24110,N_24250);
xor U25195 (N_25195,N_24152,N_24393);
xor U25196 (N_25196,N_24001,N_24178);
or U25197 (N_25197,N_24555,N_24851);
or U25198 (N_25198,N_24621,N_24667);
or U25199 (N_25199,N_24515,N_24292);
nor U25200 (N_25200,N_24249,N_24996);
xor U25201 (N_25201,N_24765,N_24962);
xnor U25202 (N_25202,N_24997,N_24240);
nand U25203 (N_25203,N_24987,N_24868);
or U25204 (N_25204,N_24963,N_24777);
nor U25205 (N_25205,N_24418,N_24478);
or U25206 (N_25206,N_24901,N_24208);
xor U25207 (N_25207,N_24925,N_24509);
or U25208 (N_25208,N_24153,N_24134);
nor U25209 (N_25209,N_24597,N_24685);
and U25210 (N_25210,N_24327,N_24084);
or U25211 (N_25211,N_24909,N_24004);
xnor U25212 (N_25212,N_24117,N_24917);
or U25213 (N_25213,N_24058,N_24406);
and U25214 (N_25214,N_24595,N_24952);
or U25215 (N_25215,N_24241,N_24746);
nand U25216 (N_25216,N_24608,N_24794);
xnor U25217 (N_25217,N_24403,N_24306);
or U25218 (N_25218,N_24378,N_24166);
nor U25219 (N_25219,N_24561,N_24135);
and U25220 (N_25220,N_24038,N_24278);
and U25221 (N_25221,N_24271,N_24349);
or U25222 (N_25222,N_24778,N_24982);
and U25223 (N_25223,N_24898,N_24939);
xor U25224 (N_25224,N_24983,N_24280);
xor U25225 (N_25225,N_24720,N_24673);
and U25226 (N_25226,N_24867,N_24700);
and U25227 (N_25227,N_24079,N_24528);
nor U25228 (N_25228,N_24850,N_24369);
and U25229 (N_25229,N_24675,N_24779);
nand U25230 (N_25230,N_24438,N_24664);
and U25231 (N_25231,N_24260,N_24428);
xnor U25232 (N_25232,N_24726,N_24864);
or U25233 (N_25233,N_24554,N_24890);
or U25234 (N_25234,N_24674,N_24571);
or U25235 (N_25235,N_24437,N_24734);
or U25236 (N_25236,N_24022,N_24974);
and U25237 (N_25237,N_24326,N_24151);
and U25238 (N_25238,N_24138,N_24756);
or U25239 (N_25239,N_24142,N_24838);
or U25240 (N_25240,N_24612,N_24910);
xor U25241 (N_25241,N_24771,N_24253);
and U25242 (N_25242,N_24565,N_24259);
and U25243 (N_25243,N_24920,N_24194);
nand U25244 (N_25244,N_24069,N_24295);
xor U25245 (N_25245,N_24036,N_24537);
nor U25246 (N_25246,N_24317,N_24310);
or U25247 (N_25247,N_24693,N_24985);
and U25248 (N_25248,N_24347,N_24559);
or U25249 (N_25249,N_24709,N_24342);
nor U25250 (N_25250,N_24730,N_24759);
nor U25251 (N_25251,N_24374,N_24312);
xor U25252 (N_25252,N_24297,N_24702);
and U25253 (N_25253,N_24857,N_24165);
nor U25254 (N_25254,N_24636,N_24629);
xor U25255 (N_25255,N_24694,N_24156);
xor U25256 (N_25256,N_24999,N_24750);
xor U25257 (N_25257,N_24174,N_24642);
and U25258 (N_25258,N_24217,N_24472);
nand U25259 (N_25259,N_24395,N_24242);
nand U25260 (N_25260,N_24443,N_24548);
and U25261 (N_25261,N_24397,N_24772);
nand U25262 (N_25262,N_24582,N_24878);
or U25263 (N_25263,N_24641,N_24780);
and U25264 (N_25264,N_24712,N_24040);
xor U25265 (N_25265,N_24063,N_24762);
or U25266 (N_25266,N_24539,N_24188);
and U25267 (N_25267,N_24100,N_24352);
xnor U25268 (N_25268,N_24535,N_24354);
nor U25269 (N_25269,N_24563,N_24361);
and U25270 (N_25270,N_24221,N_24681);
and U25271 (N_25271,N_24457,N_24927);
xnor U25272 (N_25272,N_24553,N_24930);
and U25273 (N_25273,N_24400,N_24377);
and U25274 (N_25274,N_24769,N_24024);
xor U25275 (N_25275,N_24689,N_24475);
and U25276 (N_25276,N_24731,N_24688);
and U25277 (N_25277,N_24544,N_24979);
nor U25278 (N_25278,N_24331,N_24293);
and U25279 (N_25279,N_24103,N_24866);
nand U25280 (N_25280,N_24973,N_24845);
nand U25281 (N_25281,N_24442,N_24121);
nor U25282 (N_25282,N_24970,N_24722);
nor U25283 (N_25283,N_24171,N_24954);
nand U25284 (N_25284,N_24131,N_24870);
and U25285 (N_25285,N_24824,N_24991);
or U25286 (N_25286,N_24949,N_24928);
nand U25287 (N_25287,N_24052,N_24969);
and U25288 (N_25288,N_24843,N_24682);
xnor U25289 (N_25289,N_24094,N_24366);
nor U25290 (N_25290,N_24575,N_24075);
xnor U25291 (N_25291,N_24490,N_24499);
xor U25292 (N_25292,N_24340,N_24466);
nand U25293 (N_25293,N_24192,N_24091);
nor U25294 (N_25294,N_24835,N_24385);
xnor U25295 (N_25295,N_24033,N_24841);
xor U25296 (N_25296,N_24872,N_24191);
nor U25297 (N_25297,N_24285,N_24550);
and U25298 (N_25298,N_24335,N_24020);
nor U25299 (N_25299,N_24562,N_24606);
nor U25300 (N_25300,N_24600,N_24944);
nand U25301 (N_25301,N_24000,N_24802);
and U25302 (N_25302,N_24043,N_24325);
nand U25303 (N_25303,N_24541,N_24411);
or U25304 (N_25304,N_24728,N_24671);
xor U25305 (N_25305,N_24698,N_24672);
xnor U25306 (N_25306,N_24552,N_24827);
nand U25307 (N_25307,N_24139,N_24060);
or U25308 (N_25308,N_24697,N_24818);
or U25309 (N_25309,N_24206,N_24220);
nand U25310 (N_25310,N_24787,N_24577);
nor U25311 (N_25311,N_24031,N_24598);
nand U25312 (N_25312,N_24401,N_24339);
xnor U25313 (N_25313,N_24207,N_24579);
xnor U25314 (N_25314,N_24908,N_24891);
or U25315 (N_25315,N_24721,N_24926);
or U25316 (N_25316,N_24972,N_24922);
xnor U25317 (N_25317,N_24480,N_24140);
and U25318 (N_25318,N_24258,N_24653);
xnor U25319 (N_25319,N_24127,N_24714);
xor U25320 (N_25320,N_24173,N_24267);
or U25321 (N_25321,N_24861,N_24865);
xnor U25322 (N_25322,N_24529,N_24184);
xor U25323 (N_25323,N_24815,N_24807);
xnor U25324 (N_25324,N_24921,N_24130);
or U25325 (N_25325,N_24218,N_24929);
and U25326 (N_25326,N_24887,N_24900);
and U25327 (N_25327,N_24345,N_24992);
or U25328 (N_25328,N_24360,N_24739);
nor U25329 (N_25329,N_24035,N_24763);
or U25330 (N_25330,N_24074,N_24030);
and U25331 (N_25331,N_24578,N_24961);
nand U25332 (N_25332,N_24251,N_24255);
or U25333 (N_25333,N_24798,N_24149);
or U25334 (N_25334,N_24039,N_24454);
nor U25335 (N_25335,N_24964,N_24876);
and U25336 (N_25336,N_24026,N_24077);
and U25337 (N_25337,N_24145,N_24239);
and U25338 (N_25338,N_24724,N_24879);
nand U25339 (N_25339,N_24109,N_24148);
nor U25340 (N_25340,N_24573,N_24781);
and U25341 (N_25341,N_24268,N_24445);
xnor U25342 (N_25342,N_24547,N_24014);
nor U25343 (N_25343,N_24214,N_24116);
xnor U25344 (N_25344,N_24257,N_24193);
xnor U25345 (N_25345,N_24012,N_24933);
or U25346 (N_25346,N_24067,N_24446);
or U25347 (N_25347,N_24505,N_24658);
xor U25348 (N_25348,N_24913,N_24758);
nand U25349 (N_25349,N_24518,N_24451);
and U25350 (N_25350,N_24668,N_24596);
and U25351 (N_25351,N_24452,N_24875);
or U25352 (N_25352,N_24744,N_24966);
or U25353 (N_25353,N_24054,N_24551);
or U25354 (N_25354,N_24833,N_24051);
and U25355 (N_25355,N_24050,N_24766);
and U25356 (N_25356,N_24424,N_24564);
nand U25357 (N_25357,N_24916,N_24380);
nand U25358 (N_25358,N_24289,N_24262);
nand U25359 (N_25359,N_24322,N_24439);
and U25360 (N_25360,N_24959,N_24905);
nor U25361 (N_25361,N_24526,N_24470);
and U25362 (N_25362,N_24071,N_24204);
xor U25363 (N_25363,N_24081,N_24005);
xor U25364 (N_25364,N_24315,N_24027);
xor U25365 (N_25365,N_24498,N_24367);
nand U25366 (N_25366,N_24800,N_24016);
or U25367 (N_25367,N_24183,N_24224);
and U25368 (N_25368,N_24638,N_24828);
nand U25369 (N_25369,N_24953,N_24957);
or U25370 (N_25370,N_24321,N_24727);
nand U25371 (N_25371,N_24711,N_24657);
xnor U25372 (N_25372,N_24125,N_24520);
nor U25373 (N_25373,N_24849,N_24525);
nand U25374 (N_25374,N_24299,N_24008);
and U25375 (N_25375,N_24404,N_24010);
nor U25376 (N_25376,N_24524,N_24715);
xor U25377 (N_25377,N_24978,N_24649);
or U25378 (N_25378,N_24776,N_24371);
or U25379 (N_25379,N_24161,N_24696);
nand U25380 (N_25380,N_24521,N_24316);
and U25381 (N_25381,N_24823,N_24170);
nor U25382 (N_25382,N_24484,N_24363);
or U25383 (N_25383,N_24796,N_24645);
nand U25384 (N_25384,N_24837,N_24517);
or U25385 (N_25385,N_24237,N_24243);
and U25386 (N_25386,N_24785,N_24245);
or U25387 (N_25387,N_24238,N_24187);
nand U25388 (N_25388,N_24061,N_24410);
xnor U25389 (N_25389,N_24032,N_24676);
and U25390 (N_25390,N_24936,N_24560);
nand U25391 (N_25391,N_24669,N_24046);
nand U25392 (N_25392,N_24583,N_24128);
xnor U25393 (N_25393,N_24227,N_24209);
and U25394 (N_25394,N_24203,N_24162);
nand U25395 (N_25395,N_24147,N_24215);
or U25396 (N_25396,N_24355,N_24301);
xor U25397 (N_25397,N_24307,N_24576);
or U25398 (N_25398,N_24275,N_24098);
xnor U25399 (N_25399,N_24760,N_24017);
or U25400 (N_25400,N_24545,N_24175);
nand U25401 (N_25401,N_24810,N_24994);
xor U25402 (N_25402,N_24993,N_24747);
nand U25403 (N_25403,N_24226,N_24707);
xnor U25404 (N_25404,N_24337,N_24042);
and U25405 (N_25405,N_24630,N_24889);
nor U25406 (N_25406,N_24976,N_24543);
and U25407 (N_25407,N_24918,N_24643);
nor U25408 (N_25408,N_24858,N_24635);
nor U25409 (N_25409,N_24460,N_24585);
xnor U25410 (N_25410,N_24114,N_24822);
xnor U25411 (N_25411,N_24231,N_24119);
or U25412 (N_25412,N_24044,N_24687);
xnor U25413 (N_25413,N_24995,N_24542);
nor U25414 (N_25414,N_24691,N_24883);
nand U25415 (N_25415,N_24534,N_24180);
nand U25416 (N_25416,N_24313,N_24955);
and U25417 (N_25417,N_24935,N_24273);
or U25418 (N_25418,N_24627,N_24474);
nand U25419 (N_25419,N_24190,N_24753);
or U25420 (N_25420,N_24735,N_24855);
nand U25421 (N_25421,N_24919,N_24504);
and U25422 (N_25422,N_24362,N_24817);
and U25423 (N_25423,N_24940,N_24427);
nor U25424 (N_25424,N_24806,N_24496);
nor U25425 (N_25425,N_24449,N_24387);
or U25426 (N_25426,N_24946,N_24848);
nand U25427 (N_25427,N_24431,N_24196);
or U25428 (N_25428,N_24767,N_24651);
xnor U25429 (N_25429,N_24931,N_24874);
nor U25430 (N_25430,N_24391,N_24409);
and U25431 (N_25431,N_24761,N_24350);
and U25432 (N_25432,N_24407,N_24782);
nand U25433 (N_25433,N_24620,N_24594);
and U25434 (N_25434,N_24932,N_24489);
xor U25435 (N_25435,N_24045,N_24115);
nor U25436 (N_25436,N_24911,N_24346);
or U25437 (N_25437,N_24647,N_24186);
or U25438 (N_25438,N_24225,N_24774);
and U25439 (N_25439,N_24333,N_24263);
xnor U25440 (N_25440,N_24956,N_24975);
or U25441 (N_25441,N_24988,N_24261);
nor U25442 (N_25442,N_24233,N_24906);
and U25443 (N_25443,N_24644,N_24538);
nor U25444 (N_25444,N_24646,N_24708);
or U25445 (N_25445,N_24723,N_24591);
nor U25446 (N_25446,N_24622,N_24783);
nor U25447 (N_25447,N_24338,N_24902);
or U25448 (N_25448,N_24408,N_24862);
nor U25449 (N_25449,N_24137,N_24738);
nand U25450 (N_25450,N_24618,N_24080);
nor U25451 (N_25451,N_24937,N_24655);
and U25452 (N_25452,N_24836,N_24516);
or U25453 (N_25453,N_24274,N_24095);
and U25454 (N_25454,N_24789,N_24958);
nand U25455 (N_25455,N_24468,N_24893);
nand U25456 (N_25456,N_24041,N_24444);
nor U25457 (N_25457,N_24150,N_24089);
or U25458 (N_25458,N_24291,N_24892);
xor U25459 (N_25459,N_24486,N_24205);
nor U25460 (N_25460,N_24287,N_24373);
or U25461 (N_25461,N_24652,N_24737);
nand U25462 (N_25462,N_24790,N_24323);
xor U25463 (N_25463,N_24859,N_24246);
nand U25464 (N_25464,N_24799,N_24899);
nor U25465 (N_25465,N_24717,N_24745);
and U25466 (N_25466,N_24705,N_24775);
xnor U25467 (N_25467,N_24146,N_24888);
or U25468 (N_25468,N_24482,N_24136);
nor U25469 (N_25469,N_24998,N_24092);
or U25470 (N_25470,N_24023,N_24840);
nor U25471 (N_25471,N_24229,N_24938);
nand U25472 (N_25472,N_24500,N_24968);
xor U25473 (N_25473,N_24296,N_24155);
nor U25474 (N_25474,N_24617,N_24372);
xnor U25475 (N_25475,N_24981,N_24158);
nand U25476 (N_25476,N_24254,N_24308);
and U25477 (N_25477,N_24566,N_24512);
nor U25478 (N_25478,N_24663,N_24740);
nor U25479 (N_25479,N_24159,N_24592);
nor U25480 (N_25480,N_24624,N_24143);
or U25481 (N_25481,N_24304,N_24344);
xnor U25482 (N_25482,N_24661,N_24319);
xor U25483 (N_25483,N_24768,N_24070);
xor U25484 (N_25484,N_24365,N_24376);
nand U25485 (N_25485,N_24863,N_24826);
nor U25486 (N_25486,N_24056,N_24853);
and U25487 (N_25487,N_24351,N_24228);
xor U25488 (N_25488,N_24819,N_24725);
nor U25489 (N_25489,N_24219,N_24384);
xor U25490 (N_25490,N_24426,N_24736);
nor U25491 (N_25491,N_24805,N_24510);
and U25492 (N_25492,N_24244,N_24704);
nor U25493 (N_25493,N_24533,N_24971);
xor U25494 (N_25494,N_24536,N_24834);
or U25495 (N_25495,N_24558,N_24324);
and U25496 (N_25496,N_24497,N_24062);
xnor U25497 (N_25497,N_24381,N_24068);
and U25498 (N_25498,N_24821,N_24006);
nand U25499 (N_25499,N_24695,N_24300);
or U25500 (N_25500,N_24317,N_24197);
or U25501 (N_25501,N_24446,N_24998);
nor U25502 (N_25502,N_24092,N_24039);
or U25503 (N_25503,N_24915,N_24644);
and U25504 (N_25504,N_24679,N_24894);
xnor U25505 (N_25505,N_24244,N_24749);
or U25506 (N_25506,N_24963,N_24935);
or U25507 (N_25507,N_24342,N_24320);
and U25508 (N_25508,N_24766,N_24793);
and U25509 (N_25509,N_24745,N_24769);
nor U25510 (N_25510,N_24085,N_24787);
xor U25511 (N_25511,N_24241,N_24306);
xnor U25512 (N_25512,N_24969,N_24137);
nand U25513 (N_25513,N_24828,N_24709);
nor U25514 (N_25514,N_24108,N_24005);
or U25515 (N_25515,N_24792,N_24509);
xor U25516 (N_25516,N_24229,N_24887);
nor U25517 (N_25517,N_24570,N_24000);
nor U25518 (N_25518,N_24707,N_24593);
and U25519 (N_25519,N_24860,N_24629);
or U25520 (N_25520,N_24779,N_24043);
nor U25521 (N_25521,N_24882,N_24805);
nor U25522 (N_25522,N_24746,N_24833);
xor U25523 (N_25523,N_24305,N_24630);
or U25524 (N_25524,N_24740,N_24353);
nand U25525 (N_25525,N_24041,N_24937);
nand U25526 (N_25526,N_24193,N_24638);
nor U25527 (N_25527,N_24206,N_24108);
nand U25528 (N_25528,N_24907,N_24865);
or U25529 (N_25529,N_24507,N_24643);
nor U25530 (N_25530,N_24704,N_24105);
or U25531 (N_25531,N_24379,N_24030);
or U25532 (N_25532,N_24934,N_24127);
and U25533 (N_25533,N_24341,N_24475);
nand U25534 (N_25534,N_24822,N_24066);
or U25535 (N_25535,N_24668,N_24462);
nand U25536 (N_25536,N_24834,N_24422);
and U25537 (N_25537,N_24376,N_24438);
and U25538 (N_25538,N_24914,N_24308);
nor U25539 (N_25539,N_24976,N_24722);
nor U25540 (N_25540,N_24089,N_24031);
and U25541 (N_25541,N_24125,N_24945);
nand U25542 (N_25542,N_24904,N_24525);
and U25543 (N_25543,N_24945,N_24059);
and U25544 (N_25544,N_24895,N_24964);
and U25545 (N_25545,N_24941,N_24002);
and U25546 (N_25546,N_24753,N_24759);
nand U25547 (N_25547,N_24922,N_24924);
xor U25548 (N_25548,N_24500,N_24267);
or U25549 (N_25549,N_24136,N_24632);
or U25550 (N_25550,N_24409,N_24368);
or U25551 (N_25551,N_24079,N_24227);
or U25552 (N_25552,N_24250,N_24313);
xor U25553 (N_25553,N_24390,N_24221);
xnor U25554 (N_25554,N_24986,N_24670);
xnor U25555 (N_25555,N_24455,N_24067);
and U25556 (N_25556,N_24530,N_24543);
and U25557 (N_25557,N_24735,N_24501);
or U25558 (N_25558,N_24825,N_24236);
xnor U25559 (N_25559,N_24631,N_24865);
nand U25560 (N_25560,N_24268,N_24573);
and U25561 (N_25561,N_24738,N_24586);
nor U25562 (N_25562,N_24830,N_24889);
and U25563 (N_25563,N_24024,N_24829);
or U25564 (N_25564,N_24622,N_24087);
xor U25565 (N_25565,N_24979,N_24361);
or U25566 (N_25566,N_24352,N_24844);
or U25567 (N_25567,N_24756,N_24290);
and U25568 (N_25568,N_24044,N_24402);
nor U25569 (N_25569,N_24292,N_24665);
nor U25570 (N_25570,N_24811,N_24039);
nor U25571 (N_25571,N_24771,N_24523);
or U25572 (N_25572,N_24495,N_24190);
and U25573 (N_25573,N_24120,N_24864);
nand U25574 (N_25574,N_24262,N_24402);
nor U25575 (N_25575,N_24803,N_24491);
nor U25576 (N_25576,N_24453,N_24951);
or U25577 (N_25577,N_24345,N_24516);
nor U25578 (N_25578,N_24322,N_24251);
xor U25579 (N_25579,N_24840,N_24379);
nor U25580 (N_25580,N_24624,N_24289);
xnor U25581 (N_25581,N_24715,N_24517);
and U25582 (N_25582,N_24217,N_24083);
nand U25583 (N_25583,N_24155,N_24283);
nand U25584 (N_25584,N_24431,N_24895);
nand U25585 (N_25585,N_24677,N_24219);
nand U25586 (N_25586,N_24029,N_24558);
nor U25587 (N_25587,N_24962,N_24389);
nand U25588 (N_25588,N_24177,N_24007);
and U25589 (N_25589,N_24640,N_24772);
or U25590 (N_25590,N_24822,N_24674);
nand U25591 (N_25591,N_24800,N_24421);
and U25592 (N_25592,N_24357,N_24393);
xor U25593 (N_25593,N_24820,N_24049);
nand U25594 (N_25594,N_24322,N_24547);
nand U25595 (N_25595,N_24868,N_24194);
xnor U25596 (N_25596,N_24918,N_24396);
or U25597 (N_25597,N_24110,N_24173);
or U25598 (N_25598,N_24800,N_24953);
or U25599 (N_25599,N_24625,N_24223);
nor U25600 (N_25600,N_24381,N_24482);
and U25601 (N_25601,N_24154,N_24296);
and U25602 (N_25602,N_24262,N_24129);
nand U25603 (N_25603,N_24390,N_24148);
nand U25604 (N_25604,N_24562,N_24137);
nor U25605 (N_25605,N_24041,N_24741);
xnor U25606 (N_25606,N_24656,N_24878);
xnor U25607 (N_25607,N_24095,N_24726);
or U25608 (N_25608,N_24428,N_24564);
or U25609 (N_25609,N_24764,N_24531);
xnor U25610 (N_25610,N_24066,N_24671);
or U25611 (N_25611,N_24496,N_24303);
and U25612 (N_25612,N_24788,N_24101);
and U25613 (N_25613,N_24097,N_24421);
xor U25614 (N_25614,N_24510,N_24374);
or U25615 (N_25615,N_24734,N_24228);
or U25616 (N_25616,N_24331,N_24675);
and U25617 (N_25617,N_24129,N_24363);
nand U25618 (N_25618,N_24826,N_24039);
xor U25619 (N_25619,N_24651,N_24451);
or U25620 (N_25620,N_24068,N_24354);
and U25621 (N_25621,N_24393,N_24598);
and U25622 (N_25622,N_24114,N_24723);
xnor U25623 (N_25623,N_24779,N_24240);
nor U25624 (N_25624,N_24956,N_24933);
or U25625 (N_25625,N_24523,N_24764);
nand U25626 (N_25626,N_24005,N_24884);
and U25627 (N_25627,N_24639,N_24285);
xnor U25628 (N_25628,N_24427,N_24801);
xnor U25629 (N_25629,N_24146,N_24206);
xnor U25630 (N_25630,N_24750,N_24713);
or U25631 (N_25631,N_24990,N_24718);
nand U25632 (N_25632,N_24516,N_24244);
or U25633 (N_25633,N_24367,N_24318);
or U25634 (N_25634,N_24913,N_24971);
or U25635 (N_25635,N_24901,N_24320);
nand U25636 (N_25636,N_24531,N_24449);
xnor U25637 (N_25637,N_24369,N_24091);
nor U25638 (N_25638,N_24752,N_24190);
nand U25639 (N_25639,N_24336,N_24685);
xnor U25640 (N_25640,N_24288,N_24424);
and U25641 (N_25641,N_24754,N_24601);
xnor U25642 (N_25642,N_24374,N_24222);
xnor U25643 (N_25643,N_24364,N_24997);
or U25644 (N_25644,N_24218,N_24287);
and U25645 (N_25645,N_24177,N_24290);
or U25646 (N_25646,N_24908,N_24608);
and U25647 (N_25647,N_24115,N_24961);
nor U25648 (N_25648,N_24144,N_24860);
xor U25649 (N_25649,N_24800,N_24641);
xor U25650 (N_25650,N_24166,N_24513);
or U25651 (N_25651,N_24801,N_24001);
or U25652 (N_25652,N_24985,N_24584);
xnor U25653 (N_25653,N_24909,N_24603);
or U25654 (N_25654,N_24138,N_24936);
or U25655 (N_25655,N_24479,N_24104);
or U25656 (N_25656,N_24018,N_24927);
xor U25657 (N_25657,N_24282,N_24193);
nand U25658 (N_25658,N_24820,N_24116);
xor U25659 (N_25659,N_24497,N_24569);
nand U25660 (N_25660,N_24015,N_24388);
and U25661 (N_25661,N_24827,N_24838);
and U25662 (N_25662,N_24912,N_24335);
xor U25663 (N_25663,N_24840,N_24450);
xnor U25664 (N_25664,N_24234,N_24193);
nor U25665 (N_25665,N_24757,N_24760);
nand U25666 (N_25666,N_24889,N_24902);
and U25667 (N_25667,N_24596,N_24224);
and U25668 (N_25668,N_24129,N_24014);
or U25669 (N_25669,N_24060,N_24550);
nor U25670 (N_25670,N_24585,N_24512);
nor U25671 (N_25671,N_24383,N_24314);
nor U25672 (N_25672,N_24457,N_24768);
and U25673 (N_25673,N_24767,N_24531);
and U25674 (N_25674,N_24346,N_24871);
xnor U25675 (N_25675,N_24793,N_24500);
nand U25676 (N_25676,N_24071,N_24567);
nand U25677 (N_25677,N_24973,N_24693);
or U25678 (N_25678,N_24348,N_24825);
nand U25679 (N_25679,N_24583,N_24094);
and U25680 (N_25680,N_24825,N_24046);
and U25681 (N_25681,N_24225,N_24289);
nor U25682 (N_25682,N_24321,N_24856);
xnor U25683 (N_25683,N_24929,N_24064);
nand U25684 (N_25684,N_24770,N_24580);
or U25685 (N_25685,N_24520,N_24242);
nand U25686 (N_25686,N_24107,N_24253);
xnor U25687 (N_25687,N_24531,N_24845);
nand U25688 (N_25688,N_24789,N_24923);
and U25689 (N_25689,N_24104,N_24901);
nor U25690 (N_25690,N_24587,N_24229);
and U25691 (N_25691,N_24340,N_24478);
or U25692 (N_25692,N_24222,N_24830);
and U25693 (N_25693,N_24121,N_24554);
nor U25694 (N_25694,N_24686,N_24671);
nor U25695 (N_25695,N_24006,N_24658);
nand U25696 (N_25696,N_24200,N_24982);
and U25697 (N_25697,N_24694,N_24773);
or U25698 (N_25698,N_24256,N_24916);
or U25699 (N_25699,N_24492,N_24568);
nand U25700 (N_25700,N_24590,N_24119);
nand U25701 (N_25701,N_24240,N_24933);
nand U25702 (N_25702,N_24203,N_24580);
nand U25703 (N_25703,N_24757,N_24410);
or U25704 (N_25704,N_24259,N_24724);
nor U25705 (N_25705,N_24650,N_24032);
or U25706 (N_25706,N_24513,N_24935);
or U25707 (N_25707,N_24071,N_24608);
nor U25708 (N_25708,N_24630,N_24923);
and U25709 (N_25709,N_24327,N_24048);
or U25710 (N_25710,N_24842,N_24559);
and U25711 (N_25711,N_24910,N_24209);
nor U25712 (N_25712,N_24929,N_24376);
xor U25713 (N_25713,N_24600,N_24381);
nand U25714 (N_25714,N_24062,N_24771);
or U25715 (N_25715,N_24075,N_24332);
nand U25716 (N_25716,N_24551,N_24396);
or U25717 (N_25717,N_24520,N_24462);
nand U25718 (N_25718,N_24851,N_24929);
nor U25719 (N_25719,N_24773,N_24990);
and U25720 (N_25720,N_24041,N_24664);
nand U25721 (N_25721,N_24498,N_24381);
and U25722 (N_25722,N_24924,N_24050);
xnor U25723 (N_25723,N_24498,N_24511);
and U25724 (N_25724,N_24876,N_24505);
xnor U25725 (N_25725,N_24586,N_24835);
and U25726 (N_25726,N_24278,N_24321);
xnor U25727 (N_25727,N_24738,N_24652);
nand U25728 (N_25728,N_24291,N_24121);
and U25729 (N_25729,N_24509,N_24707);
and U25730 (N_25730,N_24615,N_24322);
and U25731 (N_25731,N_24712,N_24318);
nor U25732 (N_25732,N_24080,N_24338);
or U25733 (N_25733,N_24765,N_24687);
nor U25734 (N_25734,N_24761,N_24264);
or U25735 (N_25735,N_24791,N_24562);
and U25736 (N_25736,N_24712,N_24224);
or U25737 (N_25737,N_24721,N_24394);
nor U25738 (N_25738,N_24237,N_24722);
and U25739 (N_25739,N_24793,N_24454);
xor U25740 (N_25740,N_24398,N_24300);
xnor U25741 (N_25741,N_24238,N_24620);
or U25742 (N_25742,N_24583,N_24301);
nand U25743 (N_25743,N_24977,N_24226);
nor U25744 (N_25744,N_24639,N_24560);
and U25745 (N_25745,N_24385,N_24899);
nor U25746 (N_25746,N_24490,N_24905);
nor U25747 (N_25747,N_24275,N_24051);
or U25748 (N_25748,N_24202,N_24697);
xor U25749 (N_25749,N_24863,N_24308);
and U25750 (N_25750,N_24779,N_24323);
nor U25751 (N_25751,N_24231,N_24168);
and U25752 (N_25752,N_24427,N_24209);
nand U25753 (N_25753,N_24102,N_24811);
xnor U25754 (N_25754,N_24413,N_24511);
or U25755 (N_25755,N_24423,N_24180);
xnor U25756 (N_25756,N_24288,N_24054);
or U25757 (N_25757,N_24725,N_24822);
and U25758 (N_25758,N_24248,N_24665);
and U25759 (N_25759,N_24600,N_24734);
nor U25760 (N_25760,N_24162,N_24933);
nor U25761 (N_25761,N_24156,N_24423);
nand U25762 (N_25762,N_24703,N_24732);
or U25763 (N_25763,N_24549,N_24959);
nand U25764 (N_25764,N_24216,N_24030);
nor U25765 (N_25765,N_24155,N_24842);
or U25766 (N_25766,N_24111,N_24201);
xnor U25767 (N_25767,N_24672,N_24626);
nor U25768 (N_25768,N_24937,N_24237);
nor U25769 (N_25769,N_24236,N_24647);
nand U25770 (N_25770,N_24540,N_24449);
nand U25771 (N_25771,N_24738,N_24209);
xor U25772 (N_25772,N_24939,N_24824);
xor U25773 (N_25773,N_24259,N_24991);
or U25774 (N_25774,N_24785,N_24522);
and U25775 (N_25775,N_24425,N_24141);
and U25776 (N_25776,N_24606,N_24341);
nand U25777 (N_25777,N_24524,N_24879);
and U25778 (N_25778,N_24522,N_24713);
nand U25779 (N_25779,N_24426,N_24260);
and U25780 (N_25780,N_24473,N_24389);
nor U25781 (N_25781,N_24009,N_24159);
or U25782 (N_25782,N_24545,N_24832);
xor U25783 (N_25783,N_24671,N_24062);
xnor U25784 (N_25784,N_24530,N_24320);
xor U25785 (N_25785,N_24886,N_24911);
or U25786 (N_25786,N_24625,N_24207);
and U25787 (N_25787,N_24847,N_24789);
xnor U25788 (N_25788,N_24001,N_24021);
or U25789 (N_25789,N_24445,N_24899);
xnor U25790 (N_25790,N_24629,N_24760);
and U25791 (N_25791,N_24966,N_24945);
nor U25792 (N_25792,N_24959,N_24968);
nor U25793 (N_25793,N_24988,N_24433);
or U25794 (N_25794,N_24392,N_24959);
and U25795 (N_25795,N_24587,N_24381);
nor U25796 (N_25796,N_24631,N_24581);
and U25797 (N_25797,N_24457,N_24853);
nand U25798 (N_25798,N_24957,N_24114);
xnor U25799 (N_25799,N_24683,N_24378);
or U25800 (N_25800,N_24773,N_24346);
nand U25801 (N_25801,N_24435,N_24109);
and U25802 (N_25802,N_24335,N_24373);
xor U25803 (N_25803,N_24448,N_24935);
nor U25804 (N_25804,N_24171,N_24384);
nand U25805 (N_25805,N_24253,N_24886);
or U25806 (N_25806,N_24373,N_24938);
or U25807 (N_25807,N_24590,N_24781);
nor U25808 (N_25808,N_24599,N_24093);
and U25809 (N_25809,N_24543,N_24967);
or U25810 (N_25810,N_24486,N_24649);
nor U25811 (N_25811,N_24332,N_24815);
nor U25812 (N_25812,N_24235,N_24378);
or U25813 (N_25813,N_24436,N_24126);
and U25814 (N_25814,N_24585,N_24262);
nor U25815 (N_25815,N_24293,N_24567);
nand U25816 (N_25816,N_24627,N_24493);
xor U25817 (N_25817,N_24782,N_24507);
and U25818 (N_25818,N_24560,N_24337);
nand U25819 (N_25819,N_24097,N_24759);
and U25820 (N_25820,N_24948,N_24650);
nor U25821 (N_25821,N_24208,N_24036);
or U25822 (N_25822,N_24275,N_24285);
nand U25823 (N_25823,N_24846,N_24732);
nor U25824 (N_25824,N_24589,N_24948);
or U25825 (N_25825,N_24207,N_24551);
and U25826 (N_25826,N_24454,N_24148);
xor U25827 (N_25827,N_24113,N_24495);
or U25828 (N_25828,N_24520,N_24268);
nor U25829 (N_25829,N_24746,N_24941);
and U25830 (N_25830,N_24527,N_24721);
or U25831 (N_25831,N_24724,N_24063);
and U25832 (N_25832,N_24441,N_24184);
and U25833 (N_25833,N_24966,N_24515);
and U25834 (N_25834,N_24002,N_24194);
nand U25835 (N_25835,N_24631,N_24048);
nor U25836 (N_25836,N_24368,N_24566);
and U25837 (N_25837,N_24469,N_24561);
xnor U25838 (N_25838,N_24787,N_24115);
xor U25839 (N_25839,N_24714,N_24984);
and U25840 (N_25840,N_24175,N_24550);
and U25841 (N_25841,N_24553,N_24349);
nor U25842 (N_25842,N_24828,N_24115);
or U25843 (N_25843,N_24549,N_24023);
nand U25844 (N_25844,N_24478,N_24837);
nor U25845 (N_25845,N_24866,N_24365);
nor U25846 (N_25846,N_24482,N_24048);
nor U25847 (N_25847,N_24039,N_24755);
xnor U25848 (N_25848,N_24028,N_24372);
or U25849 (N_25849,N_24744,N_24043);
nor U25850 (N_25850,N_24728,N_24767);
and U25851 (N_25851,N_24308,N_24871);
xnor U25852 (N_25852,N_24859,N_24625);
nand U25853 (N_25853,N_24446,N_24181);
nor U25854 (N_25854,N_24108,N_24371);
xnor U25855 (N_25855,N_24144,N_24570);
nor U25856 (N_25856,N_24218,N_24798);
or U25857 (N_25857,N_24412,N_24422);
nand U25858 (N_25858,N_24925,N_24106);
nor U25859 (N_25859,N_24062,N_24400);
nor U25860 (N_25860,N_24728,N_24724);
nand U25861 (N_25861,N_24390,N_24614);
xnor U25862 (N_25862,N_24712,N_24270);
nor U25863 (N_25863,N_24822,N_24807);
or U25864 (N_25864,N_24864,N_24685);
xor U25865 (N_25865,N_24806,N_24467);
and U25866 (N_25866,N_24726,N_24938);
nand U25867 (N_25867,N_24005,N_24426);
or U25868 (N_25868,N_24990,N_24686);
nor U25869 (N_25869,N_24612,N_24890);
or U25870 (N_25870,N_24974,N_24212);
nor U25871 (N_25871,N_24930,N_24829);
or U25872 (N_25872,N_24781,N_24061);
xor U25873 (N_25873,N_24883,N_24578);
and U25874 (N_25874,N_24964,N_24856);
xnor U25875 (N_25875,N_24896,N_24925);
or U25876 (N_25876,N_24314,N_24883);
nor U25877 (N_25877,N_24741,N_24972);
nor U25878 (N_25878,N_24239,N_24654);
nor U25879 (N_25879,N_24922,N_24110);
nand U25880 (N_25880,N_24075,N_24537);
nor U25881 (N_25881,N_24731,N_24253);
and U25882 (N_25882,N_24152,N_24459);
and U25883 (N_25883,N_24908,N_24478);
or U25884 (N_25884,N_24208,N_24770);
nand U25885 (N_25885,N_24906,N_24895);
nand U25886 (N_25886,N_24654,N_24858);
nor U25887 (N_25887,N_24001,N_24331);
nand U25888 (N_25888,N_24819,N_24923);
or U25889 (N_25889,N_24931,N_24126);
xnor U25890 (N_25890,N_24177,N_24097);
xor U25891 (N_25891,N_24264,N_24028);
xor U25892 (N_25892,N_24126,N_24228);
and U25893 (N_25893,N_24361,N_24713);
nor U25894 (N_25894,N_24530,N_24649);
or U25895 (N_25895,N_24045,N_24814);
nand U25896 (N_25896,N_24359,N_24363);
nand U25897 (N_25897,N_24183,N_24265);
nand U25898 (N_25898,N_24718,N_24783);
nand U25899 (N_25899,N_24033,N_24967);
xnor U25900 (N_25900,N_24805,N_24765);
nand U25901 (N_25901,N_24630,N_24767);
xnor U25902 (N_25902,N_24937,N_24722);
and U25903 (N_25903,N_24811,N_24078);
xnor U25904 (N_25904,N_24321,N_24896);
nand U25905 (N_25905,N_24501,N_24039);
nor U25906 (N_25906,N_24752,N_24811);
or U25907 (N_25907,N_24125,N_24338);
nand U25908 (N_25908,N_24140,N_24717);
and U25909 (N_25909,N_24583,N_24352);
nand U25910 (N_25910,N_24117,N_24925);
or U25911 (N_25911,N_24363,N_24277);
xor U25912 (N_25912,N_24320,N_24112);
nand U25913 (N_25913,N_24252,N_24182);
xor U25914 (N_25914,N_24411,N_24274);
nor U25915 (N_25915,N_24765,N_24832);
or U25916 (N_25916,N_24417,N_24403);
nand U25917 (N_25917,N_24068,N_24165);
xor U25918 (N_25918,N_24456,N_24060);
and U25919 (N_25919,N_24334,N_24621);
nor U25920 (N_25920,N_24064,N_24554);
or U25921 (N_25921,N_24846,N_24226);
xor U25922 (N_25922,N_24498,N_24858);
and U25923 (N_25923,N_24667,N_24486);
nand U25924 (N_25924,N_24354,N_24912);
nand U25925 (N_25925,N_24551,N_24530);
nor U25926 (N_25926,N_24914,N_24487);
nor U25927 (N_25927,N_24869,N_24254);
nand U25928 (N_25928,N_24835,N_24766);
and U25929 (N_25929,N_24254,N_24078);
xor U25930 (N_25930,N_24057,N_24094);
xor U25931 (N_25931,N_24134,N_24453);
or U25932 (N_25932,N_24829,N_24984);
nand U25933 (N_25933,N_24949,N_24287);
xnor U25934 (N_25934,N_24076,N_24282);
or U25935 (N_25935,N_24256,N_24226);
nor U25936 (N_25936,N_24676,N_24090);
or U25937 (N_25937,N_24727,N_24866);
xnor U25938 (N_25938,N_24195,N_24652);
and U25939 (N_25939,N_24151,N_24456);
xnor U25940 (N_25940,N_24382,N_24374);
xor U25941 (N_25941,N_24645,N_24409);
or U25942 (N_25942,N_24831,N_24776);
nor U25943 (N_25943,N_24938,N_24448);
and U25944 (N_25944,N_24691,N_24765);
nand U25945 (N_25945,N_24505,N_24935);
xor U25946 (N_25946,N_24536,N_24546);
and U25947 (N_25947,N_24021,N_24433);
xor U25948 (N_25948,N_24276,N_24443);
nor U25949 (N_25949,N_24276,N_24335);
nand U25950 (N_25950,N_24223,N_24803);
nand U25951 (N_25951,N_24827,N_24419);
or U25952 (N_25952,N_24992,N_24289);
nor U25953 (N_25953,N_24500,N_24744);
nand U25954 (N_25954,N_24260,N_24571);
nand U25955 (N_25955,N_24631,N_24516);
xor U25956 (N_25956,N_24279,N_24159);
xnor U25957 (N_25957,N_24181,N_24159);
or U25958 (N_25958,N_24002,N_24660);
nor U25959 (N_25959,N_24705,N_24583);
xnor U25960 (N_25960,N_24410,N_24146);
or U25961 (N_25961,N_24733,N_24436);
xor U25962 (N_25962,N_24970,N_24521);
and U25963 (N_25963,N_24047,N_24150);
nor U25964 (N_25964,N_24100,N_24456);
or U25965 (N_25965,N_24309,N_24137);
nor U25966 (N_25966,N_24532,N_24548);
or U25967 (N_25967,N_24143,N_24766);
nand U25968 (N_25968,N_24920,N_24579);
nand U25969 (N_25969,N_24707,N_24193);
xor U25970 (N_25970,N_24283,N_24450);
xor U25971 (N_25971,N_24184,N_24501);
and U25972 (N_25972,N_24204,N_24774);
xor U25973 (N_25973,N_24846,N_24937);
and U25974 (N_25974,N_24757,N_24388);
nor U25975 (N_25975,N_24391,N_24846);
xnor U25976 (N_25976,N_24352,N_24772);
and U25977 (N_25977,N_24924,N_24120);
nand U25978 (N_25978,N_24868,N_24300);
nand U25979 (N_25979,N_24960,N_24555);
and U25980 (N_25980,N_24247,N_24676);
xnor U25981 (N_25981,N_24534,N_24985);
and U25982 (N_25982,N_24986,N_24852);
nand U25983 (N_25983,N_24192,N_24685);
or U25984 (N_25984,N_24900,N_24263);
or U25985 (N_25985,N_24315,N_24901);
nand U25986 (N_25986,N_24560,N_24583);
and U25987 (N_25987,N_24808,N_24300);
xnor U25988 (N_25988,N_24801,N_24665);
nand U25989 (N_25989,N_24065,N_24806);
nand U25990 (N_25990,N_24041,N_24735);
nor U25991 (N_25991,N_24183,N_24825);
nand U25992 (N_25992,N_24468,N_24218);
nand U25993 (N_25993,N_24187,N_24098);
nor U25994 (N_25994,N_24017,N_24605);
xnor U25995 (N_25995,N_24856,N_24597);
nand U25996 (N_25996,N_24966,N_24925);
or U25997 (N_25997,N_24972,N_24721);
or U25998 (N_25998,N_24279,N_24614);
and U25999 (N_25999,N_24501,N_24587);
nand U26000 (N_26000,N_25235,N_25458);
nor U26001 (N_26001,N_25054,N_25699);
xnor U26002 (N_26002,N_25871,N_25150);
nor U26003 (N_26003,N_25934,N_25250);
nor U26004 (N_26004,N_25507,N_25634);
xor U26005 (N_26005,N_25378,N_25554);
nor U26006 (N_26006,N_25876,N_25140);
xor U26007 (N_26007,N_25447,N_25337);
nand U26008 (N_26008,N_25761,N_25468);
nand U26009 (N_26009,N_25676,N_25174);
nand U26010 (N_26010,N_25947,N_25521);
xor U26011 (N_26011,N_25734,N_25846);
nor U26012 (N_26012,N_25342,N_25954);
or U26013 (N_26013,N_25248,N_25939);
nand U26014 (N_26014,N_25074,N_25598);
nand U26015 (N_26015,N_25192,N_25181);
or U26016 (N_26016,N_25773,N_25249);
and U26017 (N_26017,N_25223,N_25182);
and U26018 (N_26018,N_25066,N_25286);
xnor U26019 (N_26019,N_25523,N_25115);
xor U26020 (N_26020,N_25518,N_25352);
nand U26021 (N_26021,N_25845,N_25608);
xnor U26022 (N_26022,N_25719,N_25051);
nand U26023 (N_26023,N_25321,N_25813);
nor U26024 (N_26024,N_25515,N_25664);
nand U26025 (N_26025,N_25013,N_25918);
nand U26026 (N_26026,N_25156,N_25986);
nor U26027 (N_26027,N_25126,N_25470);
xor U26028 (N_26028,N_25217,N_25258);
and U26029 (N_26029,N_25298,N_25390);
or U26030 (N_26030,N_25087,N_25604);
nor U26031 (N_26031,N_25536,N_25693);
and U26032 (N_26032,N_25474,N_25927);
xor U26033 (N_26033,N_25964,N_25567);
xnor U26034 (N_26034,N_25748,N_25508);
and U26035 (N_26035,N_25798,N_25835);
and U26036 (N_26036,N_25269,N_25456);
xnor U26037 (N_26037,N_25696,N_25362);
or U26038 (N_26038,N_25862,N_25102);
or U26039 (N_26039,N_25389,N_25722);
or U26040 (N_26040,N_25328,N_25014);
nor U26041 (N_26041,N_25672,N_25267);
and U26042 (N_26042,N_25842,N_25797);
or U26043 (N_26043,N_25443,N_25714);
nand U26044 (N_26044,N_25800,N_25422);
nand U26045 (N_26045,N_25516,N_25068);
nand U26046 (N_26046,N_25828,N_25301);
or U26047 (N_26047,N_25173,N_25692);
xor U26048 (N_26048,N_25681,N_25886);
and U26049 (N_26049,N_25000,N_25906);
and U26050 (N_26050,N_25732,N_25711);
and U26051 (N_26051,N_25225,N_25715);
nor U26052 (N_26052,N_25643,N_25185);
xnor U26053 (N_26053,N_25988,N_25650);
xor U26054 (N_26054,N_25602,N_25877);
or U26055 (N_26055,N_25038,N_25170);
nor U26056 (N_26056,N_25485,N_25666);
nand U26057 (N_26057,N_25701,N_25981);
nor U26058 (N_26058,N_25600,N_25319);
nand U26059 (N_26059,N_25762,N_25308);
nor U26060 (N_26060,N_25289,N_25280);
nor U26061 (N_26061,N_25429,N_25582);
or U26062 (N_26062,N_25403,N_25492);
nand U26063 (N_26063,N_25622,N_25164);
xor U26064 (N_26064,N_25490,N_25537);
or U26065 (N_26065,N_25198,N_25579);
or U26066 (N_26066,N_25256,N_25767);
nand U26067 (N_26067,N_25294,N_25398);
or U26068 (N_26068,N_25254,N_25242);
or U26069 (N_26069,N_25989,N_25824);
or U26070 (N_26070,N_25427,N_25766);
xnor U26071 (N_26071,N_25478,N_25619);
and U26072 (N_26072,N_25453,N_25612);
nor U26073 (N_26073,N_25647,N_25826);
xnor U26074 (N_26074,N_25610,N_25099);
or U26075 (N_26075,N_25060,N_25010);
xnor U26076 (N_26076,N_25159,N_25117);
or U26077 (N_26077,N_25417,N_25071);
xnor U26078 (N_26078,N_25116,N_25740);
nand U26079 (N_26079,N_25314,N_25659);
and U26080 (N_26080,N_25348,N_25146);
nor U26081 (N_26081,N_25555,N_25177);
nand U26082 (N_26082,N_25607,N_25787);
or U26083 (N_26083,N_25034,N_25752);
nand U26084 (N_26084,N_25645,N_25171);
or U26085 (N_26085,N_25464,N_25112);
or U26086 (N_26086,N_25902,N_25450);
nor U26087 (N_26087,N_25510,N_25107);
xor U26088 (N_26088,N_25799,N_25895);
nor U26089 (N_26089,N_25420,N_25239);
nor U26090 (N_26090,N_25475,N_25165);
and U26091 (N_26091,N_25514,N_25631);
xnor U26092 (N_26092,N_25392,N_25015);
nor U26093 (N_26093,N_25397,N_25993);
nand U26094 (N_26094,N_25245,N_25724);
nor U26095 (N_26095,N_25416,N_25093);
xor U26096 (N_26096,N_25519,N_25935);
or U26097 (N_26097,N_25572,N_25090);
and U26098 (N_26098,N_25794,N_25288);
or U26099 (N_26099,N_25705,N_25590);
nor U26100 (N_26100,N_25266,N_25749);
or U26101 (N_26101,N_25941,N_25606);
and U26102 (N_26102,N_25825,N_25589);
or U26103 (N_26103,N_25530,N_25931);
or U26104 (N_26104,N_25305,N_25372);
and U26105 (N_26105,N_25866,N_25229);
nand U26106 (N_26106,N_25023,N_25889);
or U26107 (N_26107,N_25671,N_25996);
or U26108 (N_26108,N_25728,N_25162);
nand U26109 (N_26109,N_25428,N_25216);
nor U26110 (N_26110,N_25349,N_25587);
nor U26111 (N_26111,N_25404,N_25039);
xor U26112 (N_26112,N_25960,N_25419);
nand U26113 (N_26113,N_25304,N_25737);
xnor U26114 (N_26114,N_25393,N_25501);
nor U26115 (N_26115,N_25230,N_25292);
nor U26116 (N_26116,N_25400,N_25726);
or U26117 (N_26117,N_25978,N_25418);
or U26118 (N_26118,N_25157,N_25955);
nand U26119 (N_26119,N_25409,N_25768);
or U26120 (N_26120,N_25599,N_25609);
and U26121 (N_26121,N_25236,N_25709);
and U26122 (N_26122,N_25985,N_25970);
nand U26123 (N_26123,N_25287,N_25961);
xnor U26124 (N_26124,N_25035,N_25439);
nand U26125 (N_26125,N_25459,N_25855);
nand U26126 (N_26126,N_25496,N_25415);
xnor U26127 (N_26127,N_25574,N_25710);
or U26128 (N_26128,N_25476,N_25884);
nor U26129 (N_26129,N_25208,N_25333);
nor U26130 (N_26130,N_25736,N_25682);
nand U26131 (N_26131,N_25114,N_25702);
xnor U26132 (N_26132,N_25848,N_25499);
and U26133 (N_26133,N_25983,N_25820);
nand U26134 (N_26134,N_25317,N_25808);
or U26135 (N_26135,N_25706,N_25780);
nand U26136 (N_26136,N_25406,N_25481);
or U26137 (N_26137,N_25119,N_25534);
or U26138 (N_26138,N_25279,N_25462);
nor U26139 (N_26139,N_25457,N_25691);
nor U26140 (N_26140,N_25641,N_25100);
nand U26141 (N_26141,N_25195,N_25479);
xnor U26142 (N_26142,N_25270,N_25153);
and U26143 (N_26143,N_25818,N_25907);
or U26144 (N_26144,N_25882,N_25080);
nand U26145 (N_26145,N_25541,N_25336);
and U26146 (N_26146,N_25027,N_25653);
nand U26147 (N_26147,N_25727,N_25327);
nor U26148 (N_26148,N_25796,N_25169);
xnor U26149 (N_26149,N_25967,N_25055);
or U26150 (N_26150,N_25984,N_25781);
nand U26151 (N_26151,N_25668,N_25442);
and U26152 (N_26152,N_25227,N_25512);
nor U26153 (N_26153,N_25841,N_25637);
and U26154 (N_26154,N_25004,N_25571);
and U26155 (N_26155,N_25956,N_25725);
nand U26156 (N_26156,N_25058,N_25811);
and U26157 (N_26157,N_25703,N_25913);
and U26158 (N_26158,N_25802,N_25969);
xnor U26159 (N_26159,N_25048,N_25391);
nand U26160 (N_26160,N_25313,N_25677);
or U26161 (N_26161,N_25311,N_25987);
and U26162 (N_26162,N_25678,N_25477);
or U26163 (N_26163,N_25777,N_25361);
nand U26164 (N_26164,N_25595,N_25751);
nand U26165 (N_26165,N_25340,N_25290);
and U26166 (N_26166,N_25898,N_25001);
and U26167 (N_26167,N_25547,N_25375);
or U26168 (N_26168,N_25148,N_25088);
nor U26169 (N_26169,N_25030,N_25928);
or U26170 (N_26170,N_25972,N_25592);
or U26171 (N_26171,N_25020,N_25371);
or U26172 (N_26172,N_25944,N_25531);
nor U26173 (N_26173,N_25872,N_25293);
nand U26174 (N_26174,N_25747,N_25809);
nor U26175 (N_26175,N_25346,N_25839);
and U26176 (N_26176,N_25785,N_25190);
nor U26177 (N_26177,N_25441,N_25366);
xor U26178 (N_26178,N_25910,N_25394);
nand U26179 (N_26179,N_25444,N_25929);
xor U26180 (N_26180,N_25847,N_25538);
nor U26181 (N_26181,N_25585,N_25557);
xnor U26182 (N_26182,N_25905,N_25203);
xor U26183 (N_26183,N_25662,N_25994);
and U26184 (N_26184,N_25132,N_25938);
and U26185 (N_26185,N_25936,N_25196);
or U26186 (N_26186,N_25665,N_25957);
or U26187 (N_26187,N_25296,N_25325);
nand U26188 (N_26188,N_25187,N_25801);
xnor U26189 (N_26189,N_25999,N_25188);
nor U26190 (N_26190,N_25613,N_25899);
nor U26191 (N_26191,N_25125,N_25383);
nand U26192 (N_26192,N_25551,N_25810);
and U26193 (N_26193,N_25875,N_25310);
or U26194 (N_26194,N_25471,N_25863);
nand U26195 (N_26195,N_25565,N_25224);
nand U26196 (N_26196,N_25903,N_25656);
or U26197 (N_26197,N_25002,N_25489);
nand U26198 (N_26198,N_25651,N_25660);
nand U26199 (N_26199,N_25275,N_25505);
nor U26200 (N_26200,N_25033,N_25306);
nor U26201 (N_26201,N_25916,N_25282);
nor U26202 (N_26202,N_25491,N_25025);
or U26203 (N_26203,N_25219,N_25106);
nand U26204 (N_26204,N_25779,N_25532);
and U26205 (N_26205,N_25615,N_25888);
nand U26206 (N_26206,N_25784,N_25617);
xor U26207 (N_26207,N_25577,N_25494);
and U26208 (N_26208,N_25949,N_25858);
xor U26209 (N_26209,N_25368,N_25979);
nor U26210 (N_26210,N_25260,N_25804);
nor U26211 (N_26211,N_25384,N_25374);
nand U26212 (N_26212,N_25614,N_25550);
or U26213 (N_26213,N_25951,N_25240);
or U26214 (N_26214,N_25118,N_25277);
nand U26215 (N_26215,N_25921,N_25483);
nor U26216 (N_26216,N_25022,N_25019);
or U26217 (N_26217,N_25620,N_25881);
nor U26218 (N_26218,N_25821,N_25454);
and U26219 (N_26219,N_25973,N_25948);
or U26220 (N_26220,N_25226,N_25109);
xnor U26221 (N_26221,N_25200,N_25209);
xnor U26222 (N_26222,N_25549,N_25220);
or U26223 (N_26223,N_25834,N_25852);
nor U26224 (N_26224,N_25199,N_25933);
xor U26225 (N_26225,N_25312,N_25497);
xnor U26226 (N_26226,N_25950,N_25210);
and U26227 (N_26227,N_25963,N_25160);
and U26228 (N_26228,N_25679,N_25104);
nor U26229 (N_26229,N_25110,N_25360);
and U26230 (N_26230,N_25894,N_25204);
and U26231 (N_26231,N_25197,N_25642);
nand U26232 (N_26232,N_25975,N_25830);
xor U26233 (N_26233,N_25237,N_25255);
or U26234 (N_26234,N_25924,N_25601);
or U26235 (N_26235,N_25867,N_25893);
nand U26236 (N_26236,N_25044,N_25186);
nor U26237 (N_26237,N_25564,N_25576);
xor U26238 (N_26238,N_25654,N_25271);
or U26239 (N_26239,N_25430,N_25111);
xor U26240 (N_26240,N_25860,N_25584);
xnor U26241 (N_26241,N_25303,N_25733);
or U26242 (N_26242,N_25755,N_25261);
or U26243 (N_26243,N_25569,N_25509);
nand U26244 (N_26244,N_25062,N_25854);
nand U26245 (N_26245,N_25788,N_25524);
or U26246 (N_26246,N_25285,N_25661);
nor U26247 (N_26247,N_25466,N_25688);
or U26248 (N_26248,N_25302,N_25221);
xnor U26249 (N_26249,N_25700,N_25029);
nor U26250 (N_26250,N_25320,N_25233);
or U26251 (N_26251,N_25018,N_25684);
nor U26252 (N_26252,N_25874,N_25201);
xnor U26253 (N_26253,N_25307,N_25021);
xnor U26254 (N_26254,N_25925,N_25354);
and U26255 (N_26255,N_25667,N_25624);
or U26256 (N_26256,N_25206,N_25982);
and U26257 (N_26257,N_25919,N_25669);
xnor U26258 (N_26258,N_25488,N_25341);
xnor U26259 (N_26259,N_25640,N_25857);
nand U26260 (N_26260,N_25425,N_25016);
xnor U26261 (N_26261,N_25032,N_25091);
or U26262 (N_26262,N_25094,N_25380);
nor U26263 (N_26263,N_25542,N_25544);
and U26264 (N_26264,N_25347,N_25228);
or U26265 (N_26265,N_25440,N_25853);
xor U26266 (N_26266,N_25382,N_25883);
xor U26267 (N_26267,N_25469,N_25353);
xnor U26268 (N_26268,N_25072,N_25364);
or U26269 (N_26269,N_25059,N_25713);
and U26270 (N_26270,N_25358,N_25851);
nor U26271 (N_26271,N_25890,N_25323);
and U26272 (N_26272,N_25695,N_25369);
nor U26273 (N_26273,N_25730,N_25652);
xor U26274 (N_26274,N_25007,N_25124);
nand U26275 (N_26275,N_25373,N_25596);
nor U26276 (N_26276,N_25388,N_25817);
or U26277 (N_26277,N_25795,N_25081);
and U26278 (N_26278,N_25411,N_25178);
nor U26279 (N_26279,N_25774,N_25128);
xnor U26280 (N_26280,N_25952,N_25526);
nor U26281 (N_26281,N_25892,N_25775);
nand U26282 (N_26282,N_25528,N_25827);
and U26283 (N_26283,N_25139,N_25721);
nand U26284 (N_26284,N_25522,N_25076);
or U26285 (N_26285,N_25593,N_25792);
or U26286 (N_26286,N_25142,N_25559);
or U26287 (N_26287,N_25067,N_25437);
or U26288 (N_26288,N_25832,N_25562);
nand U26289 (N_26289,N_25451,N_25089);
and U26290 (N_26290,N_25591,N_25042);
nor U26291 (N_26291,N_25135,N_25756);
xor U26292 (N_26292,N_25942,N_25553);
xnor U26293 (N_26293,N_25234,N_25945);
xor U26294 (N_26294,N_25739,N_25151);
xnor U26295 (N_26295,N_25920,N_25663);
xor U26296 (N_26296,N_25129,N_25829);
nand U26297 (N_26297,N_25793,N_25473);
nor U26298 (N_26298,N_25923,N_25690);
or U26299 (N_26299,N_25718,N_25145);
nor U26300 (N_26300,N_25815,N_25603);
or U26301 (N_26301,N_25356,N_25535);
xnor U26302 (N_26302,N_25729,N_25720);
xnor U26303 (N_26303,N_25315,N_25658);
nor U26304 (N_26304,N_25120,N_25446);
xor U26305 (N_26305,N_25434,N_25465);
nand U26306 (N_26306,N_25687,N_25268);
nor U26307 (N_26307,N_25316,N_25175);
xnor U26308 (N_26308,N_25697,N_25694);
nand U26309 (N_26309,N_25098,N_25791);
or U26310 (N_26310,N_25561,N_25517);
nand U26311 (N_26311,N_25363,N_25152);
or U26312 (N_26312,N_25636,N_25460);
xor U26313 (N_26313,N_25069,N_25511);
and U26314 (N_26314,N_25548,N_25163);
nor U26315 (N_26315,N_25050,N_25257);
and U26316 (N_26316,N_25545,N_25410);
or U26317 (N_26317,N_25168,N_25241);
xnor U26318 (N_26318,N_25189,N_25822);
nor U26319 (N_26319,N_25716,N_25539);
and U26320 (N_26320,N_25133,N_25786);
and U26321 (N_26321,N_25097,N_25402);
xnor U26322 (N_26322,N_25052,N_25626);
xnor U26323 (N_26323,N_25741,N_25966);
or U26324 (N_26324,N_25082,N_25202);
and U26325 (N_26325,N_25359,N_25588);
or U26326 (N_26326,N_25864,N_25502);
xor U26327 (N_26327,N_25379,N_25003);
and U26328 (N_26328,N_25686,N_25167);
xnor U26329 (N_26329,N_25309,N_25061);
nor U26330 (N_26330,N_25273,N_25041);
or U26331 (N_26331,N_25101,N_25213);
nand U26332 (N_26332,N_25017,N_25037);
and U26333 (N_26333,N_25904,N_25011);
xnor U26334 (N_26334,N_25130,N_25646);
and U26335 (N_26335,N_25597,N_25543);
nor U26336 (N_26336,N_25959,N_25707);
xor U26337 (N_26337,N_25759,N_25105);
xor U26338 (N_26338,N_25008,N_25231);
or U26339 (N_26339,N_25487,N_25085);
nor U26340 (N_26340,N_25330,N_25627);
and U26341 (N_26341,N_25395,N_25991);
and U26342 (N_26342,N_25436,N_25968);
nand U26343 (N_26343,N_25758,N_25908);
nand U26344 (N_26344,N_25435,N_25318);
nor U26345 (N_26345,N_25583,N_25036);
and U26346 (N_26346,N_25616,N_25789);
and U26347 (N_26347,N_25805,N_25806);
xor U26348 (N_26348,N_25424,N_25043);
and U26349 (N_26349,N_25423,N_25618);
nand U26350 (N_26350,N_25426,N_25265);
nand U26351 (N_26351,N_25776,N_25926);
or U26352 (N_26352,N_25772,N_25770);
nand U26353 (N_26353,N_25901,N_25922);
and U26354 (N_26354,N_25449,N_25965);
xor U26355 (N_26355,N_25191,N_25324);
or U26356 (N_26356,N_25765,N_25742);
nor U26357 (N_26357,N_25399,N_25078);
nand U26358 (N_26358,N_25744,N_25870);
and U26359 (N_26359,N_25141,N_25568);
xor U26360 (N_26360,N_25484,N_25504);
and U26361 (N_26361,N_25915,N_25276);
nand U26362 (N_26362,N_25743,N_25005);
nor U26363 (N_26363,N_25909,N_25370);
or U26364 (N_26364,N_25272,N_25322);
or U26365 (N_26365,N_25621,N_25685);
xnor U26366 (N_26366,N_25079,N_25251);
xnor U26367 (N_26367,N_25264,N_25482);
or U26368 (N_26368,N_25056,N_25012);
or U26369 (N_26369,N_25134,N_25812);
nor U26370 (N_26370,N_25529,N_25218);
nor U26371 (N_26371,N_25207,N_25083);
xor U26372 (N_26372,N_25075,N_25205);
nand U26373 (N_26373,N_25006,N_25856);
or U26374 (N_26374,N_25500,N_25556);
or U26375 (N_26375,N_25147,N_25746);
nand U26376 (N_26376,N_25026,N_25149);
or U26377 (N_26377,N_25084,N_25731);
nor U26378 (N_26378,N_25843,N_25648);
nor U26379 (N_26379,N_25448,N_25351);
xor U26380 (N_26380,N_25831,N_25253);
and U26381 (N_26381,N_25339,N_25031);
and U26382 (N_26382,N_25405,N_25558);
or U26383 (N_26383,N_25580,N_25738);
xnor U26384 (N_26384,N_25611,N_25525);
and U26385 (N_26385,N_25009,N_25252);
xnor U26386 (N_26386,N_25176,N_25452);
nor U26387 (N_26387,N_25977,N_25407);
or U26388 (N_26388,N_25086,N_25844);
xor U26389 (N_26389,N_25885,N_25381);
xnor U26390 (N_26390,N_25657,N_25334);
or U26391 (N_26391,N_25896,N_25262);
or U26392 (N_26392,N_25878,N_25345);
nor U26393 (N_26393,N_25172,N_25865);
or U26394 (N_26394,N_25143,N_25480);
nand U26395 (N_26395,N_25166,N_25520);
and U26396 (N_26396,N_25683,N_25344);
nand U26397 (N_26397,N_25533,N_25586);
and U26398 (N_26398,N_25632,N_25673);
xnor U26399 (N_26399,N_25486,N_25958);
nand U26400 (N_26400,N_25122,N_25232);
and U26401 (N_26401,N_25432,N_25343);
and U26402 (N_26402,N_25763,N_25639);
nand U26403 (N_26403,N_25943,N_25063);
nor U26404 (N_26404,N_25698,N_25995);
nand U26405 (N_26405,N_25386,N_25912);
or U26406 (N_26406,N_25623,N_25689);
nor U26407 (N_26407,N_25046,N_25814);
or U26408 (N_26408,N_25891,N_25717);
nand U26409 (N_26409,N_25385,N_25546);
or U26410 (N_26410,N_25708,N_25629);
xnor U26411 (N_26411,N_25680,N_25365);
xor U26412 (N_26412,N_25940,N_25914);
and U26413 (N_26413,N_25764,N_25295);
nand U26414 (N_26414,N_25329,N_25625);
or U26415 (N_26415,N_25495,N_25144);
and U26416 (N_26416,N_25838,N_25376);
xnor U26417 (N_26417,N_25655,N_25263);
and U26418 (N_26418,N_25723,N_25869);
or U26419 (N_26419,N_25911,N_25712);
nand U26420 (N_26420,N_25823,N_25513);
nor U26421 (N_26421,N_25527,N_25463);
or U26422 (N_26422,N_25121,N_25992);
and U26423 (N_26423,N_25753,N_25184);
nor U26424 (N_26424,N_25946,N_25045);
xor U26425 (N_26425,N_25215,N_25998);
or U26426 (N_26426,N_25879,N_25070);
or U26427 (N_26427,N_25897,N_25976);
xnor U26428 (N_26428,N_25136,N_25900);
nor U26429 (N_26429,N_25816,N_25438);
or U26430 (N_26430,N_25638,N_25335);
xor U26431 (N_26431,N_25154,N_25493);
xnor U26432 (N_26432,N_25735,N_25849);
nor U26433 (N_26433,N_25837,N_25594);
and U26434 (N_26434,N_25840,N_25243);
nor U26435 (N_26435,N_25782,N_25861);
or U26436 (N_26436,N_25297,N_25790);
nor U26437 (N_26437,N_25644,N_25754);
nand U26438 (N_26438,N_25974,N_25971);
nand U26439 (N_26439,N_25675,N_25183);
nand U26440 (N_26440,N_25778,N_25563);
nor U26441 (N_26441,N_25868,N_25445);
or U26442 (N_26442,N_25131,N_25413);
nand U26443 (N_26443,N_25506,N_25421);
xor U26444 (N_26444,N_25073,N_25807);
xnor U26445 (N_26445,N_25573,N_25750);
xor U26446 (N_26446,N_25578,N_25244);
xor U26447 (N_26447,N_25350,N_25819);
or U26448 (N_26448,N_25367,N_25455);
or U26449 (N_26449,N_25997,N_25540);
or U26450 (N_26450,N_25331,N_25222);
nor U26451 (N_26451,N_25932,N_25990);
or U26452 (N_26452,N_25096,N_25123);
xnor U26453 (N_26453,N_25850,N_25064);
or U26454 (N_26454,N_25566,N_25472);
and U26455 (N_26455,N_25357,N_25575);
and U26456 (N_26456,N_25238,N_25401);
nor U26457 (N_26457,N_25635,N_25745);
and U26458 (N_26458,N_25259,N_25103);
xnor U26459 (N_26459,N_25408,N_25560);
nand U26460 (N_26460,N_25461,N_25247);
xor U26461 (N_26461,N_25387,N_25769);
or U26462 (N_26462,N_25605,N_25284);
or U26463 (N_26463,N_25771,N_25332);
or U26464 (N_26464,N_25503,N_25278);
nor U26465 (N_26465,N_25630,N_25193);
nor U26466 (N_26466,N_25937,N_25552);
or U26467 (N_26467,N_25783,N_25953);
xnor U26468 (N_26468,N_25024,N_25833);
nand U26469 (N_26469,N_25246,N_25138);
xor U26470 (N_26470,N_25649,N_25179);
xnor U26471 (N_26471,N_25092,N_25930);
and U26472 (N_26472,N_25300,N_25028);
or U26473 (N_26473,N_25057,N_25628);
xor U26474 (N_26474,N_25467,N_25194);
or U26475 (N_26475,N_25498,N_25670);
xnor U26476 (N_26476,N_25053,N_25859);
and U26477 (N_26477,N_25214,N_25283);
nand U26478 (N_26478,N_25180,N_25077);
and U26479 (N_26479,N_25414,N_25355);
or U26480 (N_26480,N_25155,N_25570);
nand U26481 (N_26481,N_25127,N_25281);
nand U26482 (N_26482,N_25158,N_25291);
xor U26483 (N_26483,N_25980,N_25757);
and U26484 (N_26484,N_25917,N_25880);
or U26485 (N_26485,N_25674,N_25412);
or U26486 (N_26486,N_25431,N_25047);
or U26487 (N_26487,N_25873,N_25962);
nand U26488 (N_26488,N_25887,N_25299);
xor U26489 (N_26489,N_25803,N_25161);
or U26490 (N_26490,N_25113,N_25377);
or U26491 (N_26491,N_25212,N_25326);
nor U26492 (N_26492,N_25396,N_25338);
and U26493 (N_26493,N_25049,N_25095);
or U26494 (N_26494,N_25065,N_25433);
or U26495 (N_26495,N_25633,N_25040);
xnor U26496 (N_26496,N_25274,N_25704);
or U26497 (N_26497,N_25108,N_25836);
nor U26498 (N_26498,N_25760,N_25137);
nor U26499 (N_26499,N_25211,N_25581);
nor U26500 (N_26500,N_25181,N_25225);
nand U26501 (N_26501,N_25234,N_25508);
or U26502 (N_26502,N_25430,N_25008);
nand U26503 (N_26503,N_25382,N_25032);
nand U26504 (N_26504,N_25475,N_25905);
or U26505 (N_26505,N_25901,N_25935);
nor U26506 (N_26506,N_25102,N_25185);
xnor U26507 (N_26507,N_25410,N_25430);
nor U26508 (N_26508,N_25294,N_25396);
or U26509 (N_26509,N_25244,N_25079);
nand U26510 (N_26510,N_25003,N_25163);
nand U26511 (N_26511,N_25872,N_25976);
nand U26512 (N_26512,N_25206,N_25300);
and U26513 (N_26513,N_25391,N_25499);
xor U26514 (N_26514,N_25669,N_25316);
nor U26515 (N_26515,N_25305,N_25687);
and U26516 (N_26516,N_25364,N_25007);
xor U26517 (N_26517,N_25730,N_25100);
xor U26518 (N_26518,N_25399,N_25862);
nand U26519 (N_26519,N_25699,N_25311);
or U26520 (N_26520,N_25726,N_25207);
and U26521 (N_26521,N_25856,N_25341);
and U26522 (N_26522,N_25610,N_25317);
nor U26523 (N_26523,N_25978,N_25742);
or U26524 (N_26524,N_25574,N_25377);
or U26525 (N_26525,N_25221,N_25313);
or U26526 (N_26526,N_25941,N_25345);
nor U26527 (N_26527,N_25347,N_25708);
xnor U26528 (N_26528,N_25041,N_25448);
nor U26529 (N_26529,N_25708,N_25381);
and U26530 (N_26530,N_25886,N_25684);
and U26531 (N_26531,N_25892,N_25367);
and U26532 (N_26532,N_25101,N_25294);
nor U26533 (N_26533,N_25388,N_25891);
or U26534 (N_26534,N_25369,N_25419);
or U26535 (N_26535,N_25005,N_25622);
xnor U26536 (N_26536,N_25366,N_25088);
nand U26537 (N_26537,N_25018,N_25221);
nor U26538 (N_26538,N_25354,N_25709);
and U26539 (N_26539,N_25931,N_25802);
nor U26540 (N_26540,N_25750,N_25849);
nor U26541 (N_26541,N_25396,N_25768);
nand U26542 (N_26542,N_25577,N_25317);
nor U26543 (N_26543,N_25858,N_25007);
xnor U26544 (N_26544,N_25924,N_25433);
and U26545 (N_26545,N_25260,N_25515);
nand U26546 (N_26546,N_25192,N_25683);
xnor U26547 (N_26547,N_25257,N_25488);
xor U26548 (N_26548,N_25762,N_25637);
nor U26549 (N_26549,N_25054,N_25637);
nand U26550 (N_26550,N_25915,N_25389);
nor U26551 (N_26551,N_25181,N_25661);
and U26552 (N_26552,N_25055,N_25194);
or U26553 (N_26553,N_25952,N_25125);
nand U26554 (N_26554,N_25496,N_25484);
nand U26555 (N_26555,N_25429,N_25008);
xnor U26556 (N_26556,N_25583,N_25730);
or U26557 (N_26557,N_25598,N_25389);
nor U26558 (N_26558,N_25136,N_25923);
or U26559 (N_26559,N_25100,N_25375);
xor U26560 (N_26560,N_25429,N_25390);
nand U26561 (N_26561,N_25197,N_25375);
or U26562 (N_26562,N_25656,N_25972);
xnor U26563 (N_26563,N_25570,N_25970);
xor U26564 (N_26564,N_25599,N_25967);
and U26565 (N_26565,N_25622,N_25384);
nor U26566 (N_26566,N_25141,N_25039);
or U26567 (N_26567,N_25430,N_25306);
nand U26568 (N_26568,N_25780,N_25769);
xnor U26569 (N_26569,N_25184,N_25820);
nand U26570 (N_26570,N_25904,N_25281);
xnor U26571 (N_26571,N_25317,N_25917);
or U26572 (N_26572,N_25159,N_25094);
and U26573 (N_26573,N_25859,N_25535);
or U26574 (N_26574,N_25893,N_25317);
nand U26575 (N_26575,N_25623,N_25190);
nor U26576 (N_26576,N_25494,N_25927);
nand U26577 (N_26577,N_25541,N_25233);
xnor U26578 (N_26578,N_25325,N_25494);
xnor U26579 (N_26579,N_25286,N_25082);
xor U26580 (N_26580,N_25639,N_25172);
nand U26581 (N_26581,N_25498,N_25852);
or U26582 (N_26582,N_25814,N_25612);
nand U26583 (N_26583,N_25499,N_25230);
nand U26584 (N_26584,N_25620,N_25696);
nand U26585 (N_26585,N_25102,N_25384);
and U26586 (N_26586,N_25481,N_25455);
or U26587 (N_26587,N_25475,N_25404);
nor U26588 (N_26588,N_25515,N_25490);
xor U26589 (N_26589,N_25858,N_25419);
nor U26590 (N_26590,N_25843,N_25523);
xnor U26591 (N_26591,N_25192,N_25413);
or U26592 (N_26592,N_25319,N_25589);
nor U26593 (N_26593,N_25558,N_25260);
nor U26594 (N_26594,N_25587,N_25477);
and U26595 (N_26595,N_25952,N_25429);
nand U26596 (N_26596,N_25389,N_25541);
or U26597 (N_26597,N_25287,N_25843);
xor U26598 (N_26598,N_25586,N_25504);
and U26599 (N_26599,N_25935,N_25468);
or U26600 (N_26600,N_25941,N_25879);
xnor U26601 (N_26601,N_25754,N_25520);
or U26602 (N_26602,N_25489,N_25127);
nor U26603 (N_26603,N_25676,N_25268);
or U26604 (N_26604,N_25247,N_25858);
nor U26605 (N_26605,N_25768,N_25322);
or U26606 (N_26606,N_25137,N_25115);
nor U26607 (N_26607,N_25240,N_25123);
or U26608 (N_26608,N_25839,N_25597);
xor U26609 (N_26609,N_25385,N_25627);
or U26610 (N_26610,N_25160,N_25570);
and U26611 (N_26611,N_25973,N_25798);
or U26612 (N_26612,N_25426,N_25627);
or U26613 (N_26613,N_25962,N_25928);
or U26614 (N_26614,N_25773,N_25644);
nand U26615 (N_26615,N_25442,N_25229);
nand U26616 (N_26616,N_25840,N_25506);
xnor U26617 (N_26617,N_25363,N_25456);
or U26618 (N_26618,N_25007,N_25548);
xor U26619 (N_26619,N_25677,N_25819);
xnor U26620 (N_26620,N_25519,N_25186);
or U26621 (N_26621,N_25516,N_25553);
and U26622 (N_26622,N_25562,N_25839);
nor U26623 (N_26623,N_25387,N_25232);
xor U26624 (N_26624,N_25505,N_25169);
nor U26625 (N_26625,N_25327,N_25522);
and U26626 (N_26626,N_25426,N_25903);
nand U26627 (N_26627,N_25773,N_25778);
or U26628 (N_26628,N_25517,N_25125);
or U26629 (N_26629,N_25365,N_25603);
or U26630 (N_26630,N_25854,N_25809);
xor U26631 (N_26631,N_25813,N_25311);
nor U26632 (N_26632,N_25326,N_25424);
nor U26633 (N_26633,N_25307,N_25270);
and U26634 (N_26634,N_25231,N_25363);
or U26635 (N_26635,N_25228,N_25983);
and U26636 (N_26636,N_25177,N_25450);
nand U26637 (N_26637,N_25936,N_25200);
nor U26638 (N_26638,N_25284,N_25325);
nand U26639 (N_26639,N_25643,N_25711);
or U26640 (N_26640,N_25885,N_25189);
nand U26641 (N_26641,N_25214,N_25614);
nor U26642 (N_26642,N_25925,N_25465);
and U26643 (N_26643,N_25727,N_25570);
nand U26644 (N_26644,N_25594,N_25156);
nand U26645 (N_26645,N_25340,N_25894);
and U26646 (N_26646,N_25816,N_25249);
xor U26647 (N_26647,N_25052,N_25744);
or U26648 (N_26648,N_25506,N_25258);
nand U26649 (N_26649,N_25006,N_25813);
xnor U26650 (N_26650,N_25360,N_25277);
and U26651 (N_26651,N_25320,N_25355);
xnor U26652 (N_26652,N_25229,N_25437);
and U26653 (N_26653,N_25845,N_25918);
and U26654 (N_26654,N_25145,N_25398);
nand U26655 (N_26655,N_25206,N_25922);
and U26656 (N_26656,N_25548,N_25087);
and U26657 (N_26657,N_25609,N_25938);
or U26658 (N_26658,N_25542,N_25766);
and U26659 (N_26659,N_25413,N_25455);
xnor U26660 (N_26660,N_25346,N_25613);
nor U26661 (N_26661,N_25962,N_25540);
or U26662 (N_26662,N_25446,N_25783);
nor U26663 (N_26663,N_25708,N_25550);
nor U26664 (N_26664,N_25306,N_25959);
and U26665 (N_26665,N_25663,N_25329);
nand U26666 (N_26666,N_25732,N_25988);
xor U26667 (N_26667,N_25164,N_25223);
xor U26668 (N_26668,N_25403,N_25177);
nor U26669 (N_26669,N_25000,N_25538);
nand U26670 (N_26670,N_25717,N_25727);
nand U26671 (N_26671,N_25334,N_25278);
or U26672 (N_26672,N_25173,N_25013);
xnor U26673 (N_26673,N_25590,N_25951);
xor U26674 (N_26674,N_25500,N_25090);
nand U26675 (N_26675,N_25570,N_25629);
nor U26676 (N_26676,N_25602,N_25223);
nand U26677 (N_26677,N_25034,N_25928);
nand U26678 (N_26678,N_25939,N_25838);
and U26679 (N_26679,N_25639,N_25585);
xnor U26680 (N_26680,N_25412,N_25614);
nand U26681 (N_26681,N_25778,N_25380);
xor U26682 (N_26682,N_25328,N_25750);
xor U26683 (N_26683,N_25130,N_25207);
xnor U26684 (N_26684,N_25525,N_25349);
or U26685 (N_26685,N_25568,N_25331);
nor U26686 (N_26686,N_25420,N_25043);
nor U26687 (N_26687,N_25342,N_25843);
xor U26688 (N_26688,N_25127,N_25852);
nand U26689 (N_26689,N_25927,N_25666);
nor U26690 (N_26690,N_25703,N_25878);
nor U26691 (N_26691,N_25345,N_25513);
xor U26692 (N_26692,N_25069,N_25991);
nor U26693 (N_26693,N_25374,N_25126);
xnor U26694 (N_26694,N_25944,N_25450);
nor U26695 (N_26695,N_25031,N_25803);
and U26696 (N_26696,N_25700,N_25179);
and U26697 (N_26697,N_25380,N_25594);
and U26698 (N_26698,N_25923,N_25233);
and U26699 (N_26699,N_25710,N_25163);
or U26700 (N_26700,N_25708,N_25765);
and U26701 (N_26701,N_25302,N_25268);
nand U26702 (N_26702,N_25564,N_25026);
xnor U26703 (N_26703,N_25593,N_25415);
xnor U26704 (N_26704,N_25738,N_25260);
xor U26705 (N_26705,N_25804,N_25873);
xor U26706 (N_26706,N_25591,N_25079);
or U26707 (N_26707,N_25358,N_25946);
and U26708 (N_26708,N_25535,N_25896);
xnor U26709 (N_26709,N_25239,N_25426);
nor U26710 (N_26710,N_25100,N_25153);
or U26711 (N_26711,N_25250,N_25176);
or U26712 (N_26712,N_25769,N_25821);
or U26713 (N_26713,N_25890,N_25052);
nand U26714 (N_26714,N_25175,N_25689);
nand U26715 (N_26715,N_25704,N_25296);
nor U26716 (N_26716,N_25922,N_25952);
or U26717 (N_26717,N_25403,N_25282);
and U26718 (N_26718,N_25525,N_25116);
or U26719 (N_26719,N_25040,N_25374);
and U26720 (N_26720,N_25954,N_25365);
nand U26721 (N_26721,N_25772,N_25358);
xor U26722 (N_26722,N_25864,N_25327);
nand U26723 (N_26723,N_25469,N_25239);
nor U26724 (N_26724,N_25109,N_25182);
and U26725 (N_26725,N_25598,N_25243);
xor U26726 (N_26726,N_25451,N_25185);
nand U26727 (N_26727,N_25167,N_25050);
xnor U26728 (N_26728,N_25877,N_25612);
nand U26729 (N_26729,N_25605,N_25287);
nor U26730 (N_26730,N_25554,N_25091);
and U26731 (N_26731,N_25902,N_25892);
or U26732 (N_26732,N_25386,N_25857);
or U26733 (N_26733,N_25586,N_25958);
and U26734 (N_26734,N_25747,N_25999);
xor U26735 (N_26735,N_25082,N_25066);
xor U26736 (N_26736,N_25358,N_25293);
nand U26737 (N_26737,N_25494,N_25697);
xnor U26738 (N_26738,N_25345,N_25726);
xor U26739 (N_26739,N_25609,N_25239);
and U26740 (N_26740,N_25153,N_25765);
nand U26741 (N_26741,N_25375,N_25540);
or U26742 (N_26742,N_25254,N_25469);
or U26743 (N_26743,N_25547,N_25728);
nand U26744 (N_26744,N_25293,N_25706);
and U26745 (N_26745,N_25861,N_25396);
nor U26746 (N_26746,N_25650,N_25653);
nand U26747 (N_26747,N_25601,N_25778);
nor U26748 (N_26748,N_25720,N_25234);
xor U26749 (N_26749,N_25516,N_25770);
or U26750 (N_26750,N_25522,N_25211);
nor U26751 (N_26751,N_25474,N_25085);
and U26752 (N_26752,N_25203,N_25955);
nor U26753 (N_26753,N_25128,N_25824);
and U26754 (N_26754,N_25639,N_25091);
or U26755 (N_26755,N_25725,N_25710);
nand U26756 (N_26756,N_25443,N_25859);
and U26757 (N_26757,N_25281,N_25585);
nand U26758 (N_26758,N_25714,N_25250);
or U26759 (N_26759,N_25692,N_25332);
or U26760 (N_26760,N_25832,N_25014);
nand U26761 (N_26761,N_25036,N_25645);
and U26762 (N_26762,N_25849,N_25694);
nor U26763 (N_26763,N_25679,N_25255);
and U26764 (N_26764,N_25090,N_25569);
nor U26765 (N_26765,N_25617,N_25179);
xnor U26766 (N_26766,N_25869,N_25454);
or U26767 (N_26767,N_25077,N_25330);
nand U26768 (N_26768,N_25827,N_25862);
or U26769 (N_26769,N_25101,N_25830);
nor U26770 (N_26770,N_25809,N_25757);
nand U26771 (N_26771,N_25259,N_25386);
nor U26772 (N_26772,N_25614,N_25021);
and U26773 (N_26773,N_25786,N_25119);
nand U26774 (N_26774,N_25720,N_25294);
xor U26775 (N_26775,N_25502,N_25015);
nor U26776 (N_26776,N_25624,N_25292);
and U26777 (N_26777,N_25625,N_25870);
and U26778 (N_26778,N_25572,N_25604);
and U26779 (N_26779,N_25871,N_25881);
xnor U26780 (N_26780,N_25783,N_25514);
xnor U26781 (N_26781,N_25730,N_25276);
nand U26782 (N_26782,N_25639,N_25237);
xor U26783 (N_26783,N_25204,N_25424);
and U26784 (N_26784,N_25955,N_25082);
xnor U26785 (N_26785,N_25545,N_25031);
xnor U26786 (N_26786,N_25188,N_25717);
nand U26787 (N_26787,N_25308,N_25192);
and U26788 (N_26788,N_25322,N_25090);
and U26789 (N_26789,N_25556,N_25224);
nand U26790 (N_26790,N_25385,N_25261);
or U26791 (N_26791,N_25657,N_25712);
nand U26792 (N_26792,N_25441,N_25425);
nand U26793 (N_26793,N_25112,N_25400);
nand U26794 (N_26794,N_25670,N_25058);
nor U26795 (N_26795,N_25280,N_25224);
nand U26796 (N_26796,N_25595,N_25140);
nor U26797 (N_26797,N_25591,N_25332);
nor U26798 (N_26798,N_25051,N_25795);
nor U26799 (N_26799,N_25467,N_25558);
nor U26800 (N_26800,N_25137,N_25679);
nor U26801 (N_26801,N_25491,N_25049);
nor U26802 (N_26802,N_25049,N_25035);
and U26803 (N_26803,N_25037,N_25671);
and U26804 (N_26804,N_25309,N_25517);
nor U26805 (N_26805,N_25173,N_25904);
nor U26806 (N_26806,N_25215,N_25247);
xor U26807 (N_26807,N_25928,N_25663);
nand U26808 (N_26808,N_25205,N_25238);
nor U26809 (N_26809,N_25712,N_25954);
nand U26810 (N_26810,N_25105,N_25749);
nor U26811 (N_26811,N_25819,N_25075);
nor U26812 (N_26812,N_25983,N_25771);
nand U26813 (N_26813,N_25724,N_25263);
xor U26814 (N_26814,N_25133,N_25746);
nand U26815 (N_26815,N_25547,N_25403);
xor U26816 (N_26816,N_25026,N_25188);
and U26817 (N_26817,N_25149,N_25199);
xnor U26818 (N_26818,N_25953,N_25212);
nor U26819 (N_26819,N_25357,N_25935);
and U26820 (N_26820,N_25146,N_25992);
nor U26821 (N_26821,N_25410,N_25864);
and U26822 (N_26822,N_25660,N_25418);
and U26823 (N_26823,N_25057,N_25524);
nand U26824 (N_26824,N_25997,N_25516);
xnor U26825 (N_26825,N_25174,N_25417);
nor U26826 (N_26826,N_25472,N_25361);
nand U26827 (N_26827,N_25637,N_25902);
xor U26828 (N_26828,N_25499,N_25367);
xor U26829 (N_26829,N_25653,N_25376);
or U26830 (N_26830,N_25089,N_25389);
or U26831 (N_26831,N_25151,N_25421);
nor U26832 (N_26832,N_25653,N_25623);
and U26833 (N_26833,N_25318,N_25953);
or U26834 (N_26834,N_25888,N_25629);
xor U26835 (N_26835,N_25429,N_25697);
nand U26836 (N_26836,N_25782,N_25886);
xnor U26837 (N_26837,N_25707,N_25154);
nand U26838 (N_26838,N_25455,N_25201);
or U26839 (N_26839,N_25008,N_25216);
nand U26840 (N_26840,N_25913,N_25024);
and U26841 (N_26841,N_25230,N_25071);
or U26842 (N_26842,N_25788,N_25938);
or U26843 (N_26843,N_25147,N_25640);
xor U26844 (N_26844,N_25015,N_25570);
nor U26845 (N_26845,N_25234,N_25351);
xnor U26846 (N_26846,N_25592,N_25580);
or U26847 (N_26847,N_25519,N_25358);
nor U26848 (N_26848,N_25372,N_25523);
xnor U26849 (N_26849,N_25435,N_25918);
and U26850 (N_26850,N_25371,N_25861);
or U26851 (N_26851,N_25957,N_25180);
or U26852 (N_26852,N_25355,N_25075);
xnor U26853 (N_26853,N_25445,N_25426);
xor U26854 (N_26854,N_25056,N_25113);
nor U26855 (N_26855,N_25501,N_25068);
nor U26856 (N_26856,N_25160,N_25254);
or U26857 (N_26857,N_25435,N_25319);
nand U26858 (N_26858,N_25132,N_25037);
xnor U26859 (N_26859,N_25650,N_25283);
nor U26860 (N_26860,N_25384,N_25351);
and U26861 (N_26861,N_25840,N_25682);
or U26862 (N_26862,N_25392,N_25602);
and U26863 (N_26863,N_25289,N_25407);
xor U26864 (N_26864,N_25160,N_25740);
xor U26865 (N_26865,N_25984,N_25686);
xnor U26866 (N_26866,N_25982,N_25335);
nand U26867 (N_26867,N_25237,N_25176);
nand U26868 (N_26868,N_25069,N_25103);
nand U26869 (N_26869,N_25261,N_25909);
nor U26870 (N_26870,N_25923,N_25664);
nand U26871 (N_26871,N_25940,N_25743);
nand U26872 (N_26872,N_25218,N_25378);
or U26873 (N_26873,N_25852,N_25876);
and U26874 (N_26874,N_25986,N_25599);
xnor U26875 (N_26875,N_25535,N_25089);
or U26876 (N_26876,N_25926,N_25551);
nand U26877 (N_26877,N_25435,N_25617);
xor U26878 (N_26878,N_25406,N_25619);
or U26879 (N_26879,N_25258,N_25208);
xor U26880 (N_26880,N_25876,N_25257);
and U26881 (N_26881,N_25521,N_25362);
nor U26882 (N_26882,N_25972,N_25444);
or U26883 (N_26883,N_25296,N_25316);
or U26884 (N_26884,N_25125,N_25087);
nand U26885 (N_26885,N_25558,N_25042);
and U26886 (N_26886,N_25960,N_25462);
nand U26887 (N_26887,N_25643,N_25993);
xor U26888 (N_26888,N_25706,N_25726);
nor U26889 (N_26889,N_25239,N_25895);
and U26890 (N_26890,N_25329,N_25654);
or U26891 (N_26891,N_25822,N_25755);
and U26892 (N_26892,N_25751,N_25192);
nor U26893 (N_26893,N_25546,N_25991);
nor U26894 (N_26894,N_25704,N_25298);
or U26895 (N_26895,N_25707,N_25096);
nand U26896 (N_26896,N_25822,N_25531);
nand U26897 (N_26897,N_25092,N_25908);
and U26898 (N_26898,N_25538,N_25003);
xor U26899 (N_26899,N_25683,N_25576);
nor U26900 (N_26900,N_25347,N_25952);
nor U26901 (N_26901,N_25248,N_25278);
or U26902 (N_26902,N_25524,N_25178);
and U26903 (N_26903,N_25542,N_25283);
xnor U26904 (N_26904,N_25405,N_25499);
or U26905 (N_26905,N_25846,N_25632);
and U26906 (N_26906,N_25400,N_25091);
nor U26907 (N_26907,N_25990,N_25258);
nor U26908 (N_26908,N_25531,N_25950);
and U26909 (N_26909,N_25852,N_25288);
and U26910 (N_26910,N_25824,N_25041);
and U26911 (N_26911,N_25790,N_25045);
or U26912 (N_26912,N_25520,N_25251);
or U26913 (N_26913,N_25029,N_25686);
xnor U26914 (N_26914,N_25963,N_25182);
and U26915 (N_26915,N_25363,N_25716);
and U26916 (N_26916,N_25906,N_25580);
nand U26917 (N_26917,N_25511,N_25185);
and U26918 (N_26918,N_25231,N_25403);
or U26919 (N_26919,N_25645,N_25732);
xor U26920 (N_26920,N_25012,N_25830);
and U26921 (N_26921,N_25134,N_25558);
nor U26922 (N_26922,N_25533,N_25282);
nor U26923 (N_26923,N_25259,N_25039);
or U26924 (N_26924,N_25843,N_25286);
nor U26925 (N_26925,N_25404,N_25732);
xor U26926 (N_26926,N_25147,N_25717);
or U26927 (N_26927,N_25213,N_25409);
or U26928 (N_26928,N_25383,N_25572);
nor U26929 (N_26929,N_25112,N_25608);
or U26930 (N_26930,N_25341,N_25570);
xor U26931 (N_26931,N_25915,N_25975);
nand U26932 (N_26932,N_25425,N_25965);
xor U26933 (N_26933,N_25136,N_25805);
nor U26934 (N_26934,N_25797,N_25176);
xnor U26935 (N_26935,N_25893,N_25838);
xnor U26936 (N_26936,N_25990,N_25425);
nor U26937 (N_26937,N_25605,N_25936);
xnor U26938 (N_26938,N_25831,N_25893);
and U26939 (N_26939,N_25856,N_25039);
and U26940 (N_26940,N_25355,N_25098);
and U26941 (N_26941,N_25835,N_25987);
nand U26942 (N_26942,N_25034,N_25040);
and U26943 (N_26943,N_25024,N_25635);
nand U26944 (N_26944,N_25493,N_25990);
nor U26945 (N_26945,N_25412,N_25697);
xor U26946 (N_26946,N_25421,N_25429);
nor U26947 (N_26947,N_25081,N_25585);
or U26948 (N_26948,N_25270,N_25018);
nor U26949 (N_26949,N_25591,N_25741);
xnor U26950 (N_26950,N_25382,N_25929);
or U26951 (N_26951,N_25790,N_25307);
nand U26952 (N_26952,N_25224,N_25756);
nor U26953 (N_26953,N_25322,N_25605);
and U26954 (N_26954,N_25181,N_25651);
nand U26955 (N_26955,N_25152,N_25425);
nor U26956 (N_26956,N_25622,N_25817);
nor U26957 (N_26957,N_25983,N_25855);
or U26958 (N_26958,N_25458,N_25782);
or U26959 (N_26959,N_25540,N_25206);
and U26960 (N_26960,N_25624,N_25858);
xnor U26961 (N_26961,N_25855,N_25375);
or U26962 (N_26962,N_25372,N_25371);
nor U26963 (N_26963,N_25009,N_25883);
and U26964 (N_26964,N_25830,N_25289);
xor U26965 (N_26965,N_25261,N_25752);
nand U26966 (N_26966,N_25114,N_25538);
and U26967 (N_26967,N_25424,N_25580);
and U26968 (N_26968,N_25766,N_25344);
and U26969 (N_26969,N_25786,N_25454);
and U26970 (N_26970,N_25455,N_25505);
or U26971 (N_26971,N_25970,N_25396);
nor U26972 (N_26972,N_25424,N_25747);
xor U26973 (N_26973,N_25576,N_25327);
nand U26974 (N_26974,N_25212,N_25883);
nand U26975 (N_26975,N_25924,N_25287);
xor U26976 (N_26976,N_25189,N_25989);
or U26977 (N_26977,N_25995,N_25159);
or U26978 (N_26978,N_25096,N_25404);
xnor U26979 (N_26979,N_25747,N_25648);
xnor U26980 (N_26980,N_25223,N_25584);
or U26981 (N_26981,N_25139,N_25006);
or U26982 (N_26982,N_25755,N_25359);
xnor U26983 (N_26983,N_25063,N_25252);
and U26984 (N_26984,N_25862,N_25929);
or U26985 (N_26985,N_25642,N_25822);
nor U26986 (N_26986,N_25808,N_25162);
xnor U26987 (N_26987,N_25595,N_25570);
xor U26988 (N_26988,N_25729,N_25119);
and U26989 (N_26989,N_25808,N_25453);
and U26990 (N_26990,N_25496,N_25110);
and U26991 (N_26991,N_25400,N_25218);
and U26992 (N_26992,N_25193,N_25111);
nor U26993 (N_26993,N_25955,N_25629);
xor U26994 (N_26994,N_25382,N_25208);
or U26995 (N_26995,N_25826,N_25751);
or U26996 (N_26996,N_25604,N_25099);
or U26997 (N_26997,N_25124,N_25430);
xnor U26998 (N_26998,N_25544,N_25036);
or U26999 (N_26999,N_25422,N_25501);
xor U27000 (N_27000,N_26541,N_26296);
or U27001 (N_27001,N_26225,N_26482);
and U27002 (N_27002,N_26236,N_26895);
nand U27003 (N_27003,N_26184,N_26919);
or U27004 (N_27004,N_26268,N_26618);
and U27005 (N_27005,N_26059,N_26954);
nor U27006 (N_27006,N_26497,N_26393);
xor U27007 (N_27007,N_26190,N_26921);
and U27008 (N_27008,N_26906,N_26454);
or U27009 (N_27009,N_26446,N_26480);
or U27010 (N_27010,N_26743,N_26503);
xnor U27011 (N_27011,N_26256,N_26474);
or U27012 (N_27012,N_26732,N_26460);
or U27013 (N_27013,N_26778,N_26198);
or U27014 (N_27014,N_26109,N_26404);
and U27015 (N_27015,N_26138,N_26661);
nand U27016 (N_27016,N_26733,N_26413);
xor U27017 (N_27017,N_26143,N_26420);
nor U27018 (N_27018,N_26053,N_26311);
xor U27019 (N_27019,N_26683,N_26527);
nand U27020 (N_27020,N_26013,N_26955);
nand U27021 (N_27021,N_26471,N_26858);
or U27022 (N_27022,N_26774,N_26470);
nor U27023 (N_27023,N_26985,N_26362);
or U27024 (N_27024,N_26800,N_26081);
and U27025 (N_27025,N_26004,N_26770);
and U27026 (N_27026,N_26974,N_26376);
nor U27027 (N_27027,N_26408,N_26044);
nand U27028 (N_27028,N_26119,N_26685);
nand U27029 (N_27029,N_26307,N_26623);
or U27030 (N_27030,N_26982,N_26567);
xor U27031 (N_27031,N_26852,N_26656);
and U27032 (N_27032,N_26836,N_26434);
nand U27033 (N_27033,N_26767,N_26084);
and U27034 (N_27034,N_26910,N_26556);
nand U27035 (N_27035,N_26325,N_26018);
nand U27036 (N_27036,N_26811,N_26933);
nand U27037 (N_27037,N_26837,N_26019);
nor U27038 (N_27038,N_26030,N_26739);
and U27039 (N_27039,N_26417,N_26638);
nand U27040 (N_27040,N_26813,N_26211);
nor U27041 (N_27041,N_26189,N_26622);
and U27042 (N_27042,N_26841,N_26022);
or U27043 (N_27043,N_26007,N_26601);
xnor U27044 (N_27044,N_26602,N_26883);
nand U27045 (N_27045,N_26114,N_26331);
nand U27046 (N_27046,N_26864,N_26402);
nand U27047 (N_27047,N_26032,N_26709);
and U27048 (N_27048,N_26534,N_26243);
nor U27049 (N_27049,N_26006,N_26970);
nand U27050 (N_27050,N_26549,N_26241);
xor U27051 (N_27051,N_26036,N_26346);
nor U27052 (N_27052,N_26350,N_26106);
nor U27053 (N_27053,N_26940,N_26870);
nor U27054 (N_27054,N_26320,N_26738);
xnor U27055 (N_27055,N_26810,N_26688);
xnor U27056 (N_27056,N_26768,N_26449);
xnor U27057 (N_27057,N_26303,N_26597);
nor U27058 (N_27058,N_26917,N_26334);
and U27059 (N_27059,N_26377,N_26294);
xnor U27060 (N_27060,N_26002,N_26188);
or U27061 (N_27061,N_26835,N_26866);
and U27062 (N_27062,N_26664,N_26140);
or U27063 (N_27063,N_26719,N_26900);
or U27064 (N_27064,N_26599,N_26505);
or U27065 (N_27065,N_26832,N_26913);
nor U27066 (N_27066,N_26660,N_26698);
xnor U27067 (N_27067,N_26686,N_26088);
nor U27068 (N_27068,N_26441,N_26983);
xor U27069 (N_27069,N_26113,N_26747);
nor U27070 (N_27070,N_26563,N_26815);
and U27071 (N_27071,N_26422,N_26519);
and U27072 (N_27072,N_26579,N_26077);
and U27073 (N_27073,N_26516,N_26266);
or U27074 (N_27074,N_26699,N_26416);
and U27075 (N_27075,N_26082,N_26526);
nand U27076 (N_27076,N_26989,N_26171);
nor U27077 (N_27077,N_26472,N_26158);
and U27078 (N_27078,N_26169,N_26343);
and U27079 (N_27079,N_26561,N_26339);
or U27080 (N_27080,N_26639,N_26857);
or U27081 (N_27081,N_26001,N_26730);
or U27082 (N_27082,N_26851,N_26994);
nor U27083 (N_27083,N_26382,N_26406);
and U27084 (N_27084,N_26244,N_26528);
or U27085 (N_27085,N_26263,N_26340);
xnor U27086 (N_27086,N_26634,N_26038);
and U27087 (N_27087,N_26609,N_26667);
xor U27088 (N_27088,N_26378,N_26095);
or U27089 (N_27089,N_26000,N_26742);
or U27090 (N_27090,N_26112,N_26961);
nand U27091 (N_27091,N_26199,N_26876);
nor U27092 (N_27092,N_26123,N_26819);
nand U27093 (N_27093,N_26297,N_26222);
nand U27094 (N_27094,N_26783,N_26966);
nor U27095 (N_27095,N_26553,N_26170);
nand U27096 (N_27096,N_26555,N_26267);
xor U27097 (N_27097,N_26489,N_26375);
nand U27098 (N_27098,N_26322,N_26093);
or U27099 (N_27099,N_26010,N_26435);
nor U27100 (N_27100,N_26461,N_26094);
nand U27101 (N_27101,N_26429,N_26157);
and U27102 (N_27102,N_26751,N_26050);
nand U27103 (N_27103,N_26120,N_26057);
and U27104 (N_27104,N_26695,N_26293);
nand U27105 (N_27105,N_26364,N_26485);
nor U27106 (N_27106,N_26554,N_26711);
nand U27107 (N_27107,N_26672,N_26752);
nand U27108 (N_27108,N_26098,N_26260);
and U27109 (N_27109,N_26818,N_26275);
and U27110 (N_27110,N_26279,N_26637);
nand U27111 (N_27111,N_26701,N_26306);
nor U27112 (N_27112,N_26755,N_26995);
nor U27113 (N_27113,N_26608,N_26353);
or U27114 (N_27114,N_26079,N_26669);
nor U27115 (N_27115,N_26287,N_26005);
and U27116 (N_27116,N_26042,N_26809);
nand U27117 (N_27117,N_26734,N_26369);
nor U27118 (N_27118,N_26465,N_26808);
xor U27119 (N_27119,N_26744,N_26593);
nor U27120 (N_27120,N_26682,N_26504);
nand U27121 (N_27121,N_26178,N_26028);
nor U27122 (N_27122,N_26590,N_26905);
or U27123 (N_27123,N_26415,N_26899);
nand U27124 (N_27124,N_26749,N_26312);
xor U27125 (N_27125,N_26814,N_26806);
and U27126 (N_27126,N_26037,N_26075);
xor U27127 (N_27127,N_26107,N_26160);
or U27128 (N_27128,N_26721,N_26360);
or U27129 (N_27129,N_26203,N_26115);
and U27130 (N_27130,N_26889,N_26969);
and U27131 (N_27131,N_26099,N_26668);
and U27132 (N_27132,N_26365,N_26938);
nand U27133 (N_27133,N_26904,N_26968);
nand U27134 (N_27134,N_26183,N_26017);
xor U27135 (N_27135,N_26912,N_26391);
nor U27136 (N_27136,N_26574,N_26344);
nor U27137 (N_27137,N_26746,N_26568);
nor U27138 (N_27138,N_26546,N_26722);
and U27139 (N_27139,N_26849,N_26024);
or U27140 (N_27140,N_26349,N_26911);
nor U27141 (N_27141,N_26610,N_26789);
and U27142 (N_27142,N_26923,N_26598);
or U27143 (N_27143,N_26591,N_26164);
nand U27144 (N_27144,N_26736,N_26765);
xor U27145 (N_27145,N_26918,N_26569);
or U27146 (N_27146,N_26657,N_26323);
nor U27147 (N_27147,N_26288,N_26963);
nor U27148 (N_27148,N_26512,N_26802);
xnor U27149 (N_27149,N_26511,N_26562);
and U27150 (N_27150,N_26473,N_26674);
and U27151 (N_27151,N_26706,N_26759);
or U27152 (N_27152,N_26803,N_26620);
xor U27153 (N_27153,N_26552,N_26619);
xnor U27154 (N_27154,N_26934,N_26833);
xor U27155 (N_27155,N_26187,N_26087);
xor U27156 (N_27156,N_26197,N_26272);
or U27157 (N_27157,N_26831,N_26874);
nand U27158 (N_27158,N_26444,N_26853);
xor U27159 (N_27159,N_26723,N_26101);
or U27160 (N_27160,N_26863,N_26436);
nor U27161 (N_27161,N_26979,N_26621);
nand U27162 (N_27162,N_26882,N_26048);
or U27163 (N_27163,N_26679,N_26838);
xor U27164 (N_27164,N_26229,N_26418);
nor U27165 (N_27165,N_26425,N_26993);
xor U27166 (N_27166,N_26176,N_26300);
xor U27167 (N_27167,N_26697,N_26206);
xor U27168 (N_27168,N_26745,N_26606);
or U27169 (N_27169,N_26223,N_26144);
and U27170 (N_27170,N_26131,N_26359);
and U27171 (N_27171,N_26873,N_26351);
nand U27172 (N_27172,N_26582,N_26047);
nand U27173 (N_27173,N_26174,N_26467);
or U27174 (N_27174,N_26128,N_26595);
or U27175 (N_27175,N_26705,N_26948);
nand U27176 (N_27176,N_26495,N_26756);
nor U27177 (N_27177,N_26145,N_26490);
and U27178 (N_27178,N_26321,N_26137);
and U27179 (N_27179,N_26855,N_26400);
nor U27180 (N_27180,N_26161,N_26588);
and U27181 (N_27181,N_26121,N_26166);
nand U27182 (N_27182,N_26255,N_26642);
or U27183 (N_27183,N_26310,N_26513);
nand U27184 (N_27184,N_26367,N_26927);
or U27185 (N_27185,N_26845,N_26515);
xor U27186 (N_27186,N_26020,N_26283);
and U27187 (N_27187,N_26731,N_26259);
nor U27188 (N_27188,N_26068,N_26978);
or U27189 (N_27189,N_26871,N_26635);
xor U27190 (N_27190,N_26726,N_26146);
nor U27191 (N_27191,N_26510,N_26548);
xor U27192 (N_27192,N_26884,N_26647);
xor U27193 (N_27193,N_26676,N_26142);
nor U27194 (N_27194,N_26846,N_26027);
nand U27195 (N_27195,N_26600,N_26537);
xnor U27196 (N_27196,N_26403,N_26572);
and U27197 (N_27197,N_26455,N_26551);
nand U27198 (N_27198,N_26118,N_26894);
and U27199 (N_27199,N_26865,N_26580);
xnor U27200 (N_27200,N_26015,N_26258);
and U27201 (N_27201,N_26034,N_26366);
xnor U27202 (N_27202,N_26784,N_26061);
or U27203 (N_27203,N_26014,N_26265);
or U27204 (N_27204,N_26887,N_26867);
nor U27205 (N_27205,N_26085,N_26335);
xor U27206 (N_27206,N_26401,N_26076);
xnor U27207 (N_27207,N_26397,N_26735);
nand U27208 (N_27208,N_26280,N_26058);
or U27209 (N_27209,N_26196,N_26847);
and U27210 (N_27210,N_26565,N_26456);
xor U27211 (N_27211,N_26285,N_26067);
or U27212 (N_27212,N_26775,N_26453);
nor U27213 (N_27213,N_26702,N_26926);
or U27214 (N_27214,N_26330,N_26916);
and U27215 (N_27215,N_26824,N_26257);
xnor U27216 (N_27216,N_26439,N_26486);
and U27217 (N_27217,N_26689,N_26135);
nand U27218 (N_27218,N_26134,N_26844);
or U27219 (N_27219,N_26080,N_26617);
or U27220 (N_27220,N_26469,N_26932);
nor U27221 (N_27221,N_26943,N_26102);
or U27222 (N_27222,N_26771,N_26165);
nand U27223 (N_27223,N_26707,N_26720);
nor U27224 (N_27224,N_26725,N_26653);
xor U27225 (N_27225,N_26052,N_26522);
and U27226 (N_27226,N_26372,N_26336);
nor U27227 (N_27227,N_26830,N_26286);
nor U27228 (N_27228,N_26941,N_26407);
or U27229 (N_27229,N_26564,N_26097);
and U27230 (N_27230,N_26459,N_26741);
and U27231 (N_27231,N_26421,N_26262);
nand U27232 (N_27232,N_26728,N_26398);
or U27233 (N_27233,N_26517,N_26633);
or U27234 (N_27234,N_26690,N_26281);
and U27235 (N_27235,N_26754,N_26152);
xnor U27236 (N_27236,N_26298,N_26445);
nand U27237 (N_27237,N_26958,N_26999);
and U27238 (N_27238,N_26662,N_26615);
and U27239 (N_27239,N_26315,N_26319);
and U27240 (N_27240,N_26959,N_26980);
and U27241 (N_27241,N_26869,N_26484);
nor U27242 (N_27242,N_26525,N_26273);
or U27243 (N_27243,N_26877,N_26629);
xor U27244 (N_27244,N_26448,N_26305);
nor U27245 (N_27245,N_26859,N_26646);
xnor U27246 (N_27246,N_26399,N_26626);
xnor U27247 (N_27247,N_26915,N_26613);
nand U27248 (N_27248,N_26766,N_26826);
nand U27249 (N_27249,N_26872,N_26762);
nand U27250 (N_27250,N_26361,N_26089);
nand U27251 (N_27251,N_26862,N_26008);
xor U27252 (N_27252,N_26337,N_26922);
or U27253 (N_27253,N_26840,N_26231);
nor U27254 (N_27254,N_26892,N_26781);
nor U27255 (N_27255,N_26544,N_26072);
xnor U27256 (N_27256,N_26405,N_26409);
nor U27257 (N_27257,N_26172,N_26536);
nand U27258 (N_27258,N_26062,N_26828);
xnor U27259 (N_27259,N_26996,N_26960);
xnor U27260 (N_27260,N_26508,N_26247);
nor U27261 (N_27261,N_26463,N_26506);
xnor U27262 (N_27262,N_26185,N_26691);
nand U27263 (N_27263,N_26431,N_26825);
nand U27264 (N_27264,N_26854,N_26724);
nand U27265 (N_27265,N_26239,N_26096);
nand U27266 (N_27266,N_26971,N_26428);
nand U27267 (N_27267,N_26779,N_26973);
xor U27268 (N_27268,N_26217,N_26105);
or U27269 (N_27269,N_26326,N_26897);
and U27270 (N_27270,N_26909,N_26530);
xor U27271 (N_27271,N_26308,N_26205);
or U27272 (N_27272,N_26821,N_26386);
nand U27273 (N_27273,N_26631,N_26440);
and U27274 (N_27274,N_26712,N_26104);
or U27275 (N_27275,N_26925,N_26786);
nand U27276 (N_27276,N_26003,N_26529);
or U27277 (N_27277,N_26545,N_26773);
nor U27278 (N_27278,N_26603,N_26514);
nor U27279 (N_27279,N_26843,N_26476);
nand U27280 (N_27280,N_26991,N_26594);
or U27281 (N_27281,N_26487,N_26232);
xnor U27282 (N_27282,N_26521,N_26383);
nand U27283 (N_27283,N_26065,N_26498);
or U27284 (N_27284,N_26207,N_26295);
nand U27285 (N_27285,N_26538,N_26316);
nand U27286 (N_27286,N_26758,N_26499);
or U27287 (N_27287,N_26878,N_26410);
xor U27288 (N_27288,N_26776,N_26764);
xor U27289 (N_27289,N_26318,N_26289);
xnor U27290 (N_27290,N_26753,N_26043);
nor U27291 (N_27291,N_26539,N_26678);
xnor U27292 (N_27292,N_26625,N_26162);
and U27293 (N_27293,N_26136,N_26012);
or U27294 (N_27294,N_26798,N_26447);
and U27295 (N_27295,N_26981,N_26886);
xnor U27296 (N_27296,N_26129,N_26163);
nand U27297 (N_27297,N_26083,N_26788);
xnor U27298 (N_27298,N_26451,N_26956);
and U27299 (N_27299,N_26761,N_26957);
or U27300 (N_27300,N_26896,N_26936);
nand U27301 (N_27301,N_26893,N_26793);
and U27302 (N_27302,N_26898,N_26357);
nand U27303 (N_27303,N_26794,N_26108);
xor U27304 (N_27304,N_26939,N_26727);
nor U27305 (N_27305,N_26299,N_26122);
or U27306 (N_27306,N_26560,N_26975);
and U27307 (N_27307,N_26237,N_26195);
xnor U27308 (N_27308,N_26063,N_26924);
nor U27309 (N_27309,N_26861,N_26226);
xor U27310 (N_27310,N_26769,N_26935);
xnor U27311 (N_27311,N_26791,N_26253);
xor U27312 (N_27312,N_26665,N_26071);
xor U27313 (N_27313,N_26713,N_26997);
nand U27314 (N_27314,N_26799,N_26245);
xnor U27315 (N_27315,N_26204,N_26443);
or U27316 (N_27316,N_26433,N_26596);
xnor U27317 (N_27317,N_26558,N_26907);
or U27318 (N_27318,N_26117,N_26233);
and U27319 (N_27319,N_26384,N_26585);
xnor U27320 (N_27320,N_26209,N_26494);
or U27321 (N_27321,N_26414,N_26860);
nand U27322 (N_27322,N_26394,N_26827);
nor U27323 (N_27323,N_26009,N_26592);
and U27324 (N_27324,N_26354,N_26478);
nor U27325 (N_27325,N_26292,N_26891);
xnor U27326 (N_27326,N_26130,N_26442);
and U27327 (N_27327,N_26518,N_26450);
nor U27328 (N_27328,N_26483,N_26250);
xnor U27329 (N_27329,N_26868,N_26332);
nor U27330 (N_27330,N_26557,N_26202);
or U27331 (N_27331,N_26931,N_26575);
nor U27332 (N_27332,N_26612,N_26666);
nand U27333 (N_27333,N_26566,N_26908);
or U27334 (N_27334,N_26092,N_26796);
xnor U27335 (N_27335,N_26605,N_26944);
xnor U27336 (N_27336,N_26249,N_26070);
or U27337 (N_27337,N_26452,N_26133);
nand U27338 (N_27338,N_26842,N_26021);
and U27339 (N_27339,N_26227,N_26324);
nand U27340 (N_27340,N_26718,N_26920);
and U27341 (N_27341,N_26496,N_26385);
and U27342 (N_27342,N_26839,N_26348);
or U27343 (N_27343,N_26951,N_26126);
nand U27344 (N_27344,N_26524,N_26714);
and U27345 (N_27345,N_26795,N_26046);
xnor U27346 (N_27346,N_26193,N_26424);
nor U27347 (N_27347,N_26757,N_26578);
nand U27348 (N_27348,N_26073,N_26304);
or U27349 (N_27349,N_26984,N_26125);
and U27350 (N_27350,N_26500,N_26040);
nand U27351 (N_27351,N_26964,N_26329);
and U27352 (N_27352,N_26477,N_26381);
nor U27353 (N_27353,N_26438,N_26501);
and U27354 (N_27354,N_26468,N_26930);
nor U27355 (N_27355,N_26977,N_26380);
nor U27356 (N_27356,N_26587,N_26167);
nor U27357 (N_27357,N_26696,N_26992);
or U27358 (N_27358,N_26154,N_26212);
nand U27359 (N_27359,N_26186,N_26141);
or U27360 (N_27360,N_26327,N_26693);
nand U27361 (N_27361,N_26412,N_26139);
or U27362 (N_27362,N_26586,N_26708);
or U27363 (N_27363,N_26492,N_26277);
and U27364 (N_27364,N_26238,N_26986);
nor U27365 (N_27365,N_26988,N_26807);
xnor U27366 (N_27366,N_26248,N_26888);
xor U27367 (N_27367,N_26902,N_26547);
xnor U27368 (N_27368,N_26663,N_26023);
nand U27369 (N_27369,N_26645,N_26801);
nor U27370 (N_27370,N_26937,N_26159);
or U27371 (N_27371,N_26254,N_26822);
nand U27372 (N_27372,N_26432,N_26729);
xor U27373 (N_27373,N_26147,N_26488);
and U27374 (N_27374,N_26509,N_26103);
nand U27375 (N_27375,N_26234,N_26651);
nand U27376 (N_27376,N_26387,N_26031);
or U27377 (N_27377,N_26149,N_26589);
or U27378 (N_27378,N_26604,N_26881);
nor U27379 (N_27379,N_26156,N_26270);
and U27380 (N_27380,N_26390,N_26636);
nand U27381 (N_27381,N_26704,N_26879);
nand U27382 (N_27382,N_26388,N_26230);
or U27383 (N_27383,N_26535,N_26314);
xnor U27384 (N_27384,N_26987,N_26641);
or U27385 (N_27385,N_26716,N_26692);
nor U27386 (N_27386,N_26655,N_26054);
and U27387 (N_27387,N_26356,N_26033);
nor U27388 (N_27388,N_26627,N_26074);
or U27389 (N_27389,N_26584,N_26650);
nand U27390 (N_27390,N_26652,N_26278);
nor U27391 (N_27391,N_26829,N_26218);
nand U27392 (N_27392,N_26182,N_26928);
nand U27393 (N_27393,N_26942,N_26805);
xnor U27394 (N_27394,N_26155,N_26025);
nor U27395 (N_27395,N_26214,N_26252);
xor U27396 (N_27396,N_26559,N_26466);
or U27397 (N_27397,N_26675,N_26191);
or U27398 (N_27398,N_26532,N_26347);
and U27399 (N_27399,N_26903,N_26116);
nand U27400 (N_27400,N_26373,N_26782);
nor U27401 (N_27401,N_26520,N_26224);
and U27402 (N_27402,N_26111,N_26777);
nand U27403 (N_27403,N_26389,N_26370);
nor U27404 (N_27404,N_26965,N_26313);
nor U27405 (N_27405,N_26055,N_26150);
xor U27406 (N_27406,N_26901,N_26251);
xor U27407 (N_27407,N_26419,N_26817);
xnor U27408 (N_27408,N_26220,N_26570);
nand U27409 (N_27409,N_26953,N_26649);
or U27410 (N_27410,N_26531,N_26264);
nor U27411 (N_27411,N_26069,N_26790);
nand U27412 (N_27412,N_26640,N_26426);
nor U27413 (N_27413,N_26998,N_26430);
xor U27414 (N_27414,N_26885,N_26914);
and U27415 (N_27415,N_26890,N_26100);
nor U27416 (N_27416,N_26880,N_26213);
and U27417 (N_27417,N_26066,N_26309);
or U27418 (N_27418,N_26345,N_26246);
or U27419 (N_27419,N_26523,N_26792);
xnor U27420 (N_27420,N_26717,N_26284);
and U27421 (N_27421,N_26302,N_26816);
xnor U27422 (N_27422,N_26715,N_26875);
xor U27423 (N_27423,N_26671,N_26060);
and U27424 (N_27424,N_26290,N_26972);
nand U27425 (N_27425,N_26533,N_26614);
xnor U27426 (N_27426,N_26475,N_26396);
or U27427 (N_27427,N_26328,N_26291);
xnor U27428 (N_27428,N_26550,N_26947);
or U27429 (N_27429,N_26628,N_26703);
xor U27430 (N_27430,N_26481,N_26064);
or U27431 (N_27431,N_26820,N_26464);
or U27432 (N_27432,N_26049,N_26045);
nor U27433 (N_27433,N_26039,N_26571);
and U27434 (N_27434,N_26201,N_26659);
and U27435 (N_27435,N_26078,N_26670);
nor U27436 (N_27436,N_26946,N_26684);
or U27437 (N_27437,N_26427,N_26374);
and U27438 (N_27438,N_26760,N_26235);
and U27439 (N_27439,N_26379,N_26624);
nor U27440 (N_27440,N_26945,N_26240);
or U27441 (N_27441,N_26437,N_26180);
nor U27442 (N_27442,N_26127,N_26834);
and U27443 (N_27443,N_26269,N_26215);
xnor U27444 (N_27444,N_26210,N_26687);
nor U27445 (N_27445,N_26363,N_26276);
or U27446 (N_27446,N_26644,N_26700);
nor U27447 (N_27447,N_26502,N_26179);
xor U27448 (N_27448,N_26261,N_26677);
or U27449 (N_27449,N_26355,N_26763);
nor U27450 (N_27450,N_26110,N_26168);
nor U27451 (N_27451,N_26962,N_26457);
xnor U27452 (N_27452,N_26216,N_26194);
nand U27453 (N_27453,N_26173,N_26797);
nor U27454 (N_27454,N_26648,N_26630);
nand U27455 (N_27455,N_26395,N_26658);
xor U27456 (N_27456,N_26411,N_26576);
nor U27457 (N_27457,N_26352,N_26056);
nand U27458 (N_27458,N_26577,N_26581);
nand U27459 (N_27459,N_26342,N_26848);
xor U27460 (N_27460,N_26673,N_26750);
or U27461 (N_27461,N_26148,N_26772);
and U27462 (N_27462,N_26200,N_26132);
nor U27463 (N_27463,N_26804,N_26694);
nor U27464 (N_27464,N_26011,N_26242);
nor U27465 (N_27465,N_26090,N_26680);
xor U27466 (N_27466,N_26181,N_26317);
xnor U27467 (N_27467,N_26274,N_26228);
or U27468 (N_27468,N_26643,N_26542);
xnor U27469 (N_27469,N_26990,N_26823);
or U27470 (N_27470,N_26041,N_26026);
nand U27471 (N_27471,N_26737,N_26812);
xor U27472 (N_27472,N_26479,N_26301);
nor U27473 (N_27473,N_26151,N_26175);
xor U27474 (N_27474,N_26856,N_26035);
xor U27475 (N_27475,N_26462,N_26710);
xnor U27476 (N_27476,N_26221,N_26458);
nand U27477 (N_27477,N_26338,N_26632);
nor U27478 (N_27478,N_26967,N_26219);
and U27479 (N_27479,N_26607,N_26681);
and U27480 (N_27480,N_26785,N_26333);
xnor U27481 (N_27481,N_26787,N_26341);
nand U27482 (N_27482,N_26392,N_26493);
or U27483 (N_27483,N_26540,N_26091);
xor U27484 (N_27484,N_26371,N_26029);
nor U27485 (N_27485,N_26368,N_26780);
nand U27486 (N_27486,N_26543,N_26423);
and U27487 (N_27487,N_26748,N_26491);
xnor U27488 (N_27488,N_26192,N_26271);
and U27489 (N_27489,N_26051,N_26952);
nand U27490 (N_27490,N_26850,N_26616);
and U27491 (N_27491,N_26740,N_26282);
xor U27492 (N_27492,N_26950,N_26153);
nor U27493 (N_27493,N_26611,N_26358);
nand U27494 (N_27494,N_26086,N_26507);
or U27495 (N_27495,N_26177,N_26124);
nand U27496 (N_27496,N_26573,N_26949);
xnor U27497 (N_27497,N_26654,N_26016);
and U27498 (N_27498,N_26583,N_26976);
and U27499 (N_27499,N_26929,N_26208);
nand U27500 (N_27500,N_26094,N_26675);
nand U27501 (N_27501,N_26964,N_26723);
nor U27502 (N_27502,N_26888,N_26932);
or U27503 (N_27503,N_26492,N_26980);
xnor U27504 (N_27504,N_26760,N_26939);
nor U27505 (N_27505,N_26159,N_26783);
or U27506 (N_27506,N_26920,N_26329);
and U27507 (N_27507,N_26676,N_26802);
and U27508 (N_27508,N_26087,N_26320);
and U27509 (N_27509,N_26022,N_26794);
and U27510 (N_27510,N_26440,N_26452);
nand U27511 (N_27511,N_26956,N_26600);
nor U27512 (N_27512,N_26947,N_26564);
or U27513 (N_27513,N_26292,N_26100);
or U27514 (N_27514,N_26917,N_26801);
nand U27515 (N_27515,N_26380,N_26390);
and U27516 (N_27516,N_26319,N_26945);
nand U27517 (N_27517,N_26495,N_26414);
nor U27518 (N_27518,N_26697,N_26289);
nand U27519 (N_27519,N_26788,N_26811);
nor U27520 (N_27520,N_26833,N_26913);
and U27521 (N_27521,N_26174,N_26418);
nor U27522 (N_27522,N_26506,N_26616);
nand U27523 (N_27523,N_26172,N_26311);
xnor U27524 (N_27524,N_26661,N_26031);
nand U27525 (N_27525,N_26050,N_26026);
or U27526 (N_27526,N_26554,N_26355);
or U27527 (N_27527,N_26163,N_26412);
or U27528 (N_27528,N_26901,N_26292);
nor U27529 (N_27529,N_26101,N_26316);
nor U27530 (N_27530,N_26530,N_26484);
nand U27531 (N_27531,N_26987,N_26978);
and U27532 (N_27532,N_26498,N_26053);
nor U27533 (N_27533,N_26687,N_26497);
nor U27534 (N_27534,N_26810,N_26545);
nor U27535 (N_27535,N_26480,N_26643);
nor U27536 (N_27536,N_26678,N_26915);
nand U27537 (N_27537,N_26578,N_26873);
nand U27538 (N_27538,N_26991,N_26653);
and U27539 (N_27539,N_26232,N_26331);
and U27540 (N_27540,N_26692,N_26678);
nand U27541 (N_27541,N_26828,N_26830);
xor U27542 (N_27542,N_26183,N_26864);
nor U27543 (N_27543,N_26094,N_26393);
nor U27544 (N_27544,N_26097,N_26658);
and U27545 (N_27545,N_26156,N_26549);
xor U27546 (N_27546,N_26399,N_26780);
nand U27547 (N_27547,N_26565,N_26320);
or U27548 (N_27548,N_26839,N_26661);
or U27549 (N_27549,N_26914,N_26213);
nor U27550 (N_27550,N_26516,N_26199);
or U27551 (N_27551,N_26592,N_26799);
nor U27552 (N_27552,N_26510,N_26565);
nor U27553 (N_27553,N_26511,N_26113);
and U27554 (N_27554,N_26605,N_26902);
nand U27555 (N_27555,N_26594,N_26665);
and U27556 (N_27556,N_26784,N_26436);
or U27557 (N_27557,N_26707,N_26329);
nor U27558 (N_27558,N_26720,N_26563);
nand U27559 (N_27559,N_26980,N_26495);
nand U27560 (N_27560,N_26333,N_26420);
nand U27561 (N_27561,N_26539,N_26392);
or U27562 (N_27562,N_26058,N_26288);
or U27563 (N_27563,N_26123,N_26549);
and U27564 (N_27564,N_26025,N_26900);
or U27565 (N_27565,N_26011,N_26536);
or U27566 (N_27566,N_26686,N_26271);
or U27567 (N_27567,N_26339,N_26994);
or U27568 (N_27568,N_26870,N_26597);
and U27569 (N_27569,N_26526,N_26863);
nand U27570 (N_27570,N_26338,N_26544);
and U27571 (N_27571,N_26698,N_26462);
and U27572 (N_27572,N_26433,N_26328);
and U27573 (N_27573,N_26566,N_26856);
xnor U27574 (N_27574,N_26998,N_26638);
or U27575 (N_27575,N_26222,N_26651);
nor U27576 (N_27576,N_26338,N_26060);
xor U27577 (N_27577,N_26904,N_26501);
and U27578 (N_27578,N_26142,N_26975);
nor U27579 (N_27579,N_26871,N_26031);
nor U27580 (N_27580,N_26398,N_26420);
nand U27581 (N_27581,N_26167,N_26225);
and U27582 (N_27582,N_26549,N_26229);
nor U27583 (N_27583,N_26953,N_26760);
and U27584 (N_27584,N_26668,N_26244);
or U27585 (N_27585,N_26217,N_26721);
nand U27586 (N_27586,N_26348,N_26167);
nand U27587 (N_27587,N_26651,N_26624);
nor U27588 (N_27588,N_26873,N_26387);
xnor U27589 (N_27589,N_26435,N_26271);
nand U27590 (N_27590,N_26035,N_26157);
nor U27591 (N_27591,N_26752,N_26235);
nor U27592 (N_27592,N_26185,N_26970);
and U27593 (N_27593,N_26001,N_26241);
or U27594 (N_27594,N_26465,N_26671);
or U27595 (N_27595,N_26990,N_26912);
xnor U27596 (N_27596,N_26995,N_26599);
xnor U27597 (N_27597,N_26854,N_26909);
or U27598 (N_27598,N_26533,N_26280);
xnor U27599 (N_27599,N_26984,N_26263);
nand U27600 (N_27600,N_26762,N_26431);
xnor U27601 (N_27601,N_26040,N_26652);
or U27602 (N_27602,N_26503,N_26972);
nand U27603 (N_27603,N_26142,N_26175);
xor U27604 (N_27604,N_26266,N_26117);
xor U27605 (N_27605,N_26691,N_26095);
xnor U27606 (N_27606,N_26275,N_26836);
or U27607 (N_27607,N_26585,N_26129);
nor U27608 (N_27608,N_26677,N_26329);
nand U27609 (N_27609,N_26975,N_26232);
or U27610 (N_27610,N_26879,N_26558);
and U27611 (N_27611,N_26691,N_26029);
nand U27612 (N_27612,N_26942,N_26773);
xor U27613 (N_27613,N_26336,N_26437);
nor U27614 (N_27614,N_26868,N_26226);
and U27615 (N_27615,N_26211,N_26545);
xnor U27616 (N_27616,N_26446,N_26303);
and U27617 (N_27617,N_26926,N_26646);
nand U27618 (N_27618,N_26046,N_26758);
and U27619 (N_27619,N_26618,N_26584);
and U27620 (N_27620,N_26062,N_26263);
nand U27621 (N_27621,N_26947,N_26178);
and U27622 (N_27622,N_26589,N_26465);
or U27623 (N_27623,N_26908,N_26523);
and U27624 (N_27624,N_26251,N_26153);
and U27625 (N_27625,N_26552,N_26642);
and U27626 (N_27626,N_26444,N_26994);
nand U27627 (N_27627,N_26935,N_26387);
nand U27628 (N_27628,N_26428,N_26363);
or U27629 (N_27629,N_26815,N_26595);
xnor U27630 (N_27630,N_26588,N_26229);
xnor U27631 (N_27631,N_26430,N_26424);
and U27632 (N_27632,N_26517,N_26091);
nor U27633 (N_27633,N_26728,N_26075);
xor U27634 (N_27634,N_26781,N_26221);
or U27635 (N_27635,N_26788,N_26139);
nand U27636 (N_27636,N_26793,N_26164);
or U27637 (N_27637,N_26993,N_26469);
nand U27638 (N_27638,N_26069,N_26589);
nand U27639 (N_27639,N_26228,N_26983);
nor U27640 (N_27640,N_26079,N_26176);
or U27641 (N_27641,N_26981,N_26894);
or U27642 (N_27642,N_26803,N_26192);
and U27643 (N_27643,N_26893,N_26154);
nor U27644 (N_27644,N_26662,N_26189);
nand U27645 (N_27645,N_26390,N_26409);
nor U27646 (N_27646,N_26635,N_26880);
nand U27647 (N_27647,N_26334,N_26251);
nor U27648 (N_27648,N_26529,N_26309);
xnor U27649 (N_27649,N_26335,N_26616);
nand U27650 (N_27650,N_26199,N_26157);
and U27651 (N_27651,N_26437,N_26365);
or U27652 (N_27652,N_26092,N_26874);
xnor U27653 (N_27653,N_26236,N_26527);
nand U27654 (N_27654,N_26582,N_26188);
or U27655 (N_27655,N_26418,N_26009);
and U27656 (N_27656,N_26748,N_26822);
and U27657 (N_27657,N_26661,N_26693);
xor U27658 (N_27658,N_26200,N_26728);
nand U27659 (N_27659,N_26330,N_26026);
nor U27660 (N_27660,N_26835,N_26761);
xnor U27661 (N_27661,N_26260,N_26320);
or U27662 (N_27662,N_26010,N_26501);
xnor U27663 (N_27663,N_26306,N_26062);
nor U27664 (N_27664,N_26806,N_26755);
nor U27665 (N_27665,N_26664,N_26268);
or U27666 (N_27666,N_26185,N_26149);
and U27667 (N_27667,N_26679,N_26050);
xnor U27668 (N_27668,N_26368,N_26256);
xor U27669 (N_27669,N_26290,N_26412);
or U27670 (N_27670,N_26367,N_26256);
xnor U27671 (N_27671,N_26540,N_26393);
or U27672 (N_27672,N_26837,N_26054);
nand U27673 (N_27673,N_26475,N_26043);
nor U27674 (N_27674,N_26795,N_26630);
xor U27675 (N_27675,N_26023,N_26826);
xor U27676 (N_27676,N_26926,N_26324);
xnor U27677 (N_27677,N_26232,N_26653);
or U27678 (N_27678,N_26691,N_26993);
nor U27679 (N_27679,N_26000,N_26790);
nand U27680 (N_27680,N_26390,N_26039);
nand U27681 (N_27681,N_26076,N_26087);
nor U27682 (N_27682,N_26204,N_26035);
or U27683 (N_27683,N_26980,N_26001);
or U27684 (N_27684,N_26642,N_26628);
or U27685 (N_27685,N_26236,N_26286);
nor U27686 (N_27686,N_26608,N_26792);
nand U27687 (N_27687,N_26826,N_26836);
or U27688 (N_27688,N_26742,N_26937);
or U27689 (N_27689,N_26872,N_26035);
xor U27690 (N_27690,N_26797,N_26542);
nor U27691 (N_27691,N_26517,N_26562);
nand U27692 (N_27692,N_26269,N_26095);
xnor U27693 (N_27693,N_26698,N_26362);
or U27694 (N_27694,N_26138,N_26976);
nor U27695 (N_27695,N_26231,N_26683);
or U27696 (N_27696,N_26047,N_26117);
or U27697 (N_27697,N_26111,N_26289);
or U27698 (N_27698,N_26379,N_26317);
or U27699 (N_27699,N_26301,N_26596);
nand U27700 (N_27700,N_26762,N_26456);
nand U27701 (N_27701,N_26340,N_26120);
or U27702 (N_27702,N_26043,N_26444);
and U27703 (N_27703,N_26305,N_26283);
xor U27704 (N_27704,N_26646,N_26397);
or U27705 (N_27705,N_26692,N_26192);
xor U27706 (N_27706,N_26221,N_26193);
xor U27707 (N_27707,N_26228,N_26190);
xor U27708 (N_27708,N_26237,N_26108);
nor U27709 (N_27709,N_26870,N_26016);
and U27710 (N_27710,N_26288,N_26455);
or U27711 (N_27711,N_26237,N_26806);
nor U27712 (N_27712,N_26498,N_26078);
xnor U27713 (N_27713,N_26731,N_26081);
and U27714 (N_27714,N_26428,N_26544);
or U27715 (N_27715,N_26427,N_26326);
nor U27716 (N_27716,N_26517,N_26964);
nor U27717 (N_27717,N_26515,N_26197);
and U27718 (N_27718,N_26254,N_26767);
nor U27719 (N_27719,N_26893,N_26982);
nor U27720 (N_27720,N_26082,N_26254);
nand U27721 (N_27721,N_26023,N_26338);
or U27722 (N_27722,N_26370,N_26964);
nor U27723 (N_27723,N_26594,N_26899);
nand U27724 (N_27724,N_26447,N_26888);
nand U27725 (N_27725,N_26449,N_26576);
xnor U27726 (N_27726,N_26482,N_26715);
nor U27727 (N_27727,N_26488,N_26762);
or U27728 (N_27728,N_26096,N_26608);
nand U27729 (N_27729,N_26180,N_26367);
xor U27730 (N_27730,N_26976,N_26661);
nor U27731 (N_27731,N_26627,N_26783);
or U27732 (N_27732,N_26270,N_26474);
xor U27733 (N_27733,N_26689,N_26209);
xnor U27734 (N_27734,N_26600,N_26556);
or U27735 (N_27735,N_26437,N_26030);
or U27736 (N_27736,N_26292,N_26589);
or U27737 (N_27737,N_26032,N_26488);
nor U27738 (N_27738,N_26375,N_26604);
nand U27739 (N_27739,N_26066,N_26576);
xnor U27740 (N_27740,N_26679,N_26512);
xnor U27741 (N_27741,N_26943,N_26225);
nor U27742 (N_27742,N_26453,N_26110);
xor U27743 (N_27743,N_26081,N_26417);
xor U27744 (N_27744,N_26955,N_26700);
or U27745 (N_27745,N_26297,N_26537);
nor U27746 (N_27746,N_26355,N_26680);
nor U27747 (N_27747,N_26171,N_26747);
and U27748 (N_27748,N_26198,N_26752);
and U27749 (N_27749,N_26194,N_26992);
nand U27750 (N_27750,N_26607,N_26715);
nand U27751 (N_27751,N_26770,N_26154);
or U27752 (N_27752,N_26143,N_26788);
xor U27753 (N_27753,N_26543,N_26003);
xnor U27754 (N_27754,N_26564,N_26633);
nor U27755 (N_27755,N_26020,N_26594);
xnor U27756 (N_27756,N_26557,N_26234);
nor U27757 (N_27757,N_26443,N_26219);
or U27758 (N_27758,N_26540,N_26389);
nor U27759 (N_27759,N_26852,N_26082);
or U27760 (N_27760,N_26234,N_26197);
and U27761 (N_27761,N_26110,N_26857);
nor U27762 (N_27762,N_26582,N_26333);
or U27763 (N_27763,N_26642,N_26970);
xor U27764 (N_27764,N_26217,N_26990);
or U27765 (N_27765,N_26928,N_26531);
nor U27766 (N_27766,N_26433,N_26626);
xnor U27767 (N_27767,N_26526,N_26212);
xor U27768 (N_27768,N_26651,N_26174);
xor U27769 (N_27769,N_26859,N_26021);
nand U27770 (N_27770,N_26766,N_26015);
nand U27771 (N_27771,N_26109,N_26389);
or U27772 (N_27772,N_26191,N_26616);
nand U27773 (N_27773,N_26090,N_26745);
nor U27774 (N_27774,N_26650,N_26505);
nor U27775 (N_27775,N_26523,N_26865);
or U27776 (N_27776,N_26647,N_26116);
nor U27777 (N_27777,N_26287,N_26931);
nor U27778 (N_27778,N_26646,N_26296);
xor U27779 (N_27779,N_26641,N_26735);
nand U27780 (N_27780,N_26771,N_26431);
or U27781 (N_27781,N_26850,N_26153);
nand U27782 (N_27782,N_26691,N_26406);
and U27783 (N_27783,N_26421,N_26939);
xnor U27784 (N_27784,N_26416,N_26439);
and U27785 (N_27785,N_26782,N_26078);
nand U27786 (N_27786,N_26429,N_26524);
xor U27787 (N_27787,N_26447,N_26757);
xnor U27788 (N_27788,N_26870,N_26784);
nor U27789 (N_27789,N_26843,N_26019);
xnor U27790 (N_27790,N_26145,N_26734);
or U27791 (N_27791,N_26461,N_26829);
xnor U27792 (N_27792,N_26746,N_26734);
or U27793 (N_27793,N_26281,N_26154);
or U27794 (N_27794,N_26619,N_26787);
nor U27795 (N_27795,N_26040,N_26014);
xnor U27796 (N_27796,N_26528,N_26423);
or U27797 (N_27797,N_26589,N_26857);
nand U27798 (N_27798,N_26773,N_26487);
or U27799 (N_27799,N_26039,N_26905);
or U27800 (N_27800,N_26838,N_26385);
xor U27801 (N_27801,N_26319,N_26588);
xor U27802 (N_27802,N_26244,N_26123);
nand U27803 (N_27803,N_26123,N_26729);
xnor U27804 (N_27804,N_26111,N_26893);
xor U27805 (N_27805,N_26064,N_26398);
xor U27806 (N_27806,N_26356,N_26405);
and U27807 (N_27807,N_26172,N_26794);
nor U27808 (N_27808,N_26771,N_26681);
or U27809 (N_27809,N_26917,N_26996);
nor U27810 (N_27810,N_26717,N_26188);
nor U27811 (N_27811,N_26634,N_26937);
nand U27812 (N_27812,N_26839,N_26786);
nor U27813 (N_27813,N_26877,N_26029);
xor U27814 (N_27814,N_26712,N_26060);
xnor U27815 (N_27815,N_26099,N_26746);
and U27816 (N_27816,N_26509,N_26604);
nand U27817 (N_27817,N_26214,N_26584);
or U27818 (N_27818,N_26078,N_26281);
nand U27819 (N_27819,N_26346,N_26682);
nand U27820 (N_27820,N_26482,N_26372);
xnor U27821 (N_27821,N_26546,N_26738);
or U27822 (N_27822,N_26204,N_26873);
and U27823 (N_27823,N_26685,N_26496);
or U27824 (N_27824,N_26469,N_26023);
nor U27825 (N_27825,N_26257,N_26767);
or U27826 (N_27826,N_26917,N_26418);
nor U27827 (N_27827,N_26086,N_26184);
or U27828 (N_27828,N_26866,N_26181);
nor U27829 (N_27829,N_26761,N_26632);
xnor U27830 (N_27830,N_26360,N_26369);
xor U27831 (N_27831,N_26206,N_26861);
or U27832 (N_27832,N_26012,N_26609);
xor U27833 (N_27833,N_26101,N_26483);
xor U27834 (N_27834,N_26052,N_26559);
and U27835 (N_27835,N_26055,N_26426);
nor U27836 (N_27836,N_26744,N_26506);
and U27837 (N_27837,N_26761,N_26444);
or U27838 (N_27838,N_26310,N_26803);
nor U27839 (N_27839,N_26773,N_26842);
xnor U27840 (N_27840,N_26220,N_26824);
nor U27841 (N_27841,N_26131,N_26567);
or U27842 (N_27842,N_26140,N_26734);
nand U27843 (N_27843,N_26413,N_26037);
or U27844 (N_27844,N_26212,N_26516);
xnor U27845 (N_27845,N_26206,N_26958);
or U27846 (N_27846,N_26829,N_26630);
and U27847 (N_27847,N_26390,N_26534);
or U27848 (N_27848,N_26248,N_26136);
or U27849 (N_27849,N_26997,N_26153);
nor U27850 (N_27850,N_26939,N_26423);
nand U27851 (N_27851,N_26606,N_26216);
or U27852 (N_27852,N_26808,N_26648);
and U27853 (N_27853,N_26053,N_26276);
nand U27854 (N_27854,N_26931,N_26167);
and U27855 (N_27855,N_26906,N_26224);
nand U27856 (N_27856,N_26827,N_26449);
nand U27857 (N_27857,N_26923,N_26296);
and U27858 (N_27858,N_26796,N_26917);
xnor U27859 (N_27859,N_26848,N_26818);
xnor U27860 (N_27860,N_26706,N_26727);
nand U27861 (N_27861,N_26861,N_26919);
and U27862 (N_27862,N_26157,N_26240);
nand U27863 (N_27863,N_26700,N_26566);
nor U27864 (N_27864,N_26752,N_26706);
nor U27865 (N_27865,N_26189,N_26212);
or U27866 (N_27866,N_26793,N_26721);
and U27867 (N_27867,N_26176,N_26247);
xor U27868 (N_27868,N_26260,N_26553);
or U27869 (N_27869,N_26372,N_26594);
nor U27870 (N_27870,N_26575,N_26682);
xnor U27871 (N_27871,N_26288,N_26561);
xnor U27872 (N_27872,N_26229,N_26940);
or U27873 (N_27873,N_26090,N_26442);
nor U27874 (N_27874,N_26302,N_26065);
or U27875 (N_27875,N_26972,N_26427);
and U27876 (N_27876,N_26125,N_26869);
or U27877 (N_27877,N_26621,N_26600);
and U27878 (N_27878,N_26003,N_26376);
nor U27879 (N_27879,N_26656,N_26800);
and U27880 (N_27880,N_26286,N_26745);
nand U27881 (N_27881,N_26702,N_26378);
and U27882 (N_27882,N_26687,N_26051);
or U27883 (N_27883,N_26628,N_26283);
or U27884 (N_27884,N_26970,N_26615);
and U27885 (N_27885,N_26118,N_26875);
and U27886 (N_27886,N_26269,N_26176);
xor U27887 (N_27887,N_26627,N_26118);
nor U27888 (N_27888,N_26713,N_26616);
xor U27889 (N_27889,N_26028,N_26122);
nor U27890 (N_27890,N_26825,N_26659);
or U27891 (N_27891,N_26141,N_26453);
xnor U27892 (N_27892,N_26177,N_26964);
xor U27893 (N_27893,N_26223,N_26927);
nor U27894 (N_27894,N_26365,N_26179);
xor U27895 (N_27895,N_26592,N_26645);
and U27896 (N_27896,N_26716,N_26725);
nand U27897 (N_27897,N_26867,N_26173);
and U27898 (N_27898,N_26848,N_26797);
and U27899 (N_27899,N_26070,N_26051);
nand U27900 (N_27900,N_26844,N_26765);
or U27901 (N_27901,N_26484,N_26258);
nand U27902 (N_27902,N_26649,N_26985);
or U27903 (N_27903,N_26364,N_26851);
xor U27904 (N_27904,N_26058,N_26467);
nand U27905 (N_27905,N_26219,N_26684);
nor U27906 (N_27906,N_26351,N_26068);
nand U27907 (N_27907,N_26241,N_26757);
nand U27908 (N_27908,N_26990,N_26526);
nor U27909 (N_27909,N_26936,N_26460);
xnor U27910 (N_27910,N_26363,N_26471);
or U27911 (N_27911,N_26834,N_26278);
xor U27912 (N_27912,N_26928,N_26279);
nor U27913 (N_27913,N_26308,N_26368);
and U27914 (N_27914,N_26709,N_26859);
and U27915 (N_27915,N_26284,N_26375);
nor U27916 (N_27916,N_26603,N_26411);
nand U27917 (N_27917,N_26491,N_26833);
nand U27918 (N_27918,N_26087,N_26210);
and U27919 (N_27919,N_26203,N_26511);
and U27920 (N_27920,N_26566,N_26544);
nand U27921 (N_27921,N_26268,N_26365);
and U27922 (N_27922,N_26727,N_26646);
xor U27923 (N_27923,N_26177,N_26000);
xnor U27924 (N_27924,N_26382,N_26786);
nor U27925 (N_27925,N_26865,N_26539);
or U27926 (N_27926,N_26122,N_26757);
and U27927 (N_27927,N_26853,N_26272);
nor U27928 (N_27928,N_26641,N_26007);
nand U27929 (N_27929,N_26364,N_26402);
and U27930 (N_27930,N_26087,N_26495);
and U27931 (N_27931,N_26899,N_26663);
nand U27932 (N_27932,N_26986,N_26072);
and U27933 (N_27933,N_26830,N_26817);
nand U27934 (N_27934,N_26618,N_26021);
xnor U27935 (N_27935,N_26389,N_26892);
nor U27936 (N_27936,N_26462,N_26510);
nand U27937 (N_27937,N_26302,N_26664);
nor U27938 (N_27938,N_26041,N_26606);
and U27939 (N_27939,N_26074,N_26138);
xor U27940 (N_27940,N_26218,N_26759);
or U27941 (N_27941,N_26136,N_26298);
and U27942 (N_27942,N_26269,N_26924);
and U27943 (N_27943,N_26158,N_26245);
xor U27944 (N_27944,N_26127,N_26880);
nor U27945 (N_27945,N_26535,N_26131);
and U27946 (N_27946,N_26137,N_26684);
nand U27947 (N_27947,N_26479,N_26191);
nor U27948 (N_27948,N_26922,N_26057);
nor U27949 (N_27949,N_26218,N_26612);
xnor U27950 (N_27950,N_26096,N_26809);
and U27951 (N_27951,N_26530,N_26356);
xor U27952 (N_27952,N_26832,N_26987);
xnor U27953 (N_27953,N_26946,N_26006);
xnor U27954 (N_27954,N_26015,N_26051);
and U27955 (N_27955,N_26802,N_26539);
and U27956 (N_27956,N_26891,N_26538);
xnor U27957 (N_27957,N_26734,N_26203);
and U27958 (N_27958,N_26991,N_26237);
nor U27959 (N_27959,N_26396,N_26691);
nand U27960 (N_27960,N_26188,N_26057);
or U27961 (N_27961,N_26712,N_26716);
or U27962 (N_27962,N_26618,N_26344);
nand U27963 (N_27963,N_26051,N_26708);
and U27964 (N_27964,N_26317,N_26162);
xnor U27965 (N_27965,N_26785,N_26520);
and U27966 (N_27966,N_26446,N_26295);
xor U27967 (N_27967,N_26428,N_26946);
xnor U27968 (N_27968,N_26815,N_26650);
and U27969 (N_27969,N_26995,N_26309);
nand U27970 (N_27970,N_26630,N_26924);
xnor U27971 (N_27971,N_26477,N_26964);
xor U27972 (N_27972,N_26273,N_26359);
and U27973 (N_27973,N_26541,N_26984);
or U27974 (N_27974,N_26385,N_26895);
xnor U27975 (N_27975,N_26426,N_26907);
nand U27976 (N_27976,N_26100,N_26943);
and U27977 (N_27977,N_26870,N_26041);
xnor U27978 (N_27978,N_26814,N_26280);
nand U27979 (N_27979,N_26640,N_26826);
or U27980 (N_27980,N_26753,N_26425);
or U27981 (N_27981,N_26981,N_26696);
and U27982 (N_27982,N_26927,N_26456);
xnor U27983 (N_27983,N_26480,N_26393);
xor U27984 (N_27984,N_26682,N_26859);
and U27985 (N_27985,N_26167,N_26681);
and U27986 (N_27986,N_26712,N_26776);
xnor U27987 (N_27987,N_26300,N_26341);
nand U27988 (N_27988,N_26771,N_26875);
nand U27989 (N_27989,N_26259,N_26003);
xnor U27990 (N_27990,N_26483,N_26968);
and U27991 (N_27991,N_26546,N_26906);
or U27992 (N_27992,N_26143,N_26306);
or U27993 (N_27993,N_26415,N_26956);
nor U27994 (N_27994,N_26598,N_26069);
nor U27995 (N_27995,N_26239,N_26695);
and U27996 (N_27996,N_26110,N_26044);
nor U27997 (N_27997,N_26895,N_26001);
and U27998 (N_27998,N_26440,N_26405);
xor U27999 (N_27999,N_26938,N_26766);
and U28000 (N_28000,N_27672,N_27057);
and U28001 (N_28001,N_27684,N_27938);
nand U28002 (N_28002,N_27438,N_27676);
nand U28003 (N_28003,N_27584,N_27119);
or U28004 (N_28004,N_27709,N_27964);
nor U28005 (N_28005,N_27960,N_27050);
nor U28006 (N_28006,N_27562,N_27995);
or U28007 (N_28007,N_27434,N_27303);
xor U28008 (N_28008,N_27895,N_27178);
nor U28009 (N_28009,N_27332,N_27358);
nand U28010 (N_28010,N_27070,N_27167);
xor U28011 (N_28011,N_27716,N_27413);
nor U28012 (N_28012,N_27124,N_27678);
xnor U28013 (N_28013,N_27444,N_27028);
nand U28014 (N_28014,N_27707,N_27309);
or U28015 (N_28015,N_27915,N_27181);
or U28016 (N_28016,N_27592,N_27018);
or U28017 (N_28017,N_27862,N_27816);
or U28018 (N_28018,N_27474,N_27525);
and U28019 (N_28019,N_27841,N_27172);
nor U28020 (N_28020,N_27488,N_27962);
or U28021 (N_28021,N_27887,N_27865);
xor U28022 (N_28022,N_27643,N_27593);
and U28023 (N_28023,N_27763,N_27105);
nor U28024 (N_28024,N_27086,N_27958);
nor U28025 (N_28025,N_27100,N_27576);
or U28026 (N_28026,N_27904,N_27701);
and U28027 (N_28027,N_27024,N_27943);
nor U28028 (N_28028,N_27538,N_27829);
xnor U28029 (N_28029,N_27273,N_27751);
and U28030 (N_28030,N_27374,N_27547);
or U28031 (N_28031,N_27598,N_27099);
nor U28032 (N_28032,N_27612,N_27885);
and U28033 (N_28033,N_27421,N_27809);
nand U28034 (N_28034,N_27839,N_27311);
nor U28035 (N_28035,N_27649,N_27361);
xnor U28036 (N_28036,N_27875,N_27770);
xor U28037 (N_28037,N_27208,N_27138);
nand U28038 (N_28038,N_27985,N_27692);
and U28039 (N_28039,N_27949,N_27133);
nor U28040 (N_28040,N_27121,N_27994);
and U28041 (N_28041,N_27876,N_27450);
or U28042 (N_28042,N_27320,N_27858);
or U28043 (N_28043,N_27927,N_27842);
and U28044 (N_28044,N_27458,N_27477);
and U28045 (N_28045,N_27834,N_27799);
and U28046 (N_28046,N_27624,N_27803);
nand U28047 (N_28047,N_27398,N_27744);
xnor U28048 (N_28048,N_27338,N_27517);
xnor U28049 (N_28049,N_27503,N_27725);
xor U28050 (N_28050,N_27571,N_27023);
xnor U28051 (N_28051,N_27778,N_27369);
nand U28052 (N_28052,N_27628,N_27342);
and U28053 (N_28053,N_27227,N_27804);
nor U28054 (N_28054,N_27674,N_27510);
xnor U28055 (N_28055,N_27671,N_27791);
nand U28056 (N_28056,N_27840,N_27681);
xnor U28057 (N_28057,N_27917,N_27360);
nor U28058 (N_28058,N_27722,N_27104);
nand U28059 (N_28059,N_27148,N_27341);
nand U28060 (N_28060,N_27171,N_27093);
and U28061 (N_28061,N_27176,N_27288);
nor U28062 (N_28062,N_27245,N_27997);
or U28063 (N_28063,N_27587,N_27020);
and U28064 (N_28064,N_27255,N_27122);
or U28065 (N_28065,N_27185,N_27063);
or U28066 (N_28066,N_27098,N_27597);
or U28067 (N_28067,N_27975,N_27578);
nor U28068 (N_28068,N_27388,N_27696);
nand U28069 (N_28069,N_27500,N_27715);
or U28070 (N_28070,N_27989,N_27430);
or U28071 (N_28071,N_27198,N_27683);
nor U28072 (N_28072,N_27627,N_27354);
nor U28073 (N_28073,N_27765,N_27297);
and U28074 (N_28074,N_27053,N_27397);
nand U28075 (N_28075,N_27077,N_27864);
xor U28076 (N_28076,N_27455,N_27760);
or U28077 (N_28077,N_27195,N_27505);
nand U28078 (N_28078,N_27193,N_27449);
nand U28079 (N_28079,N_27118,N_27890);
and U28080 (N_28080,N_27512,N_27331);
and U28081 (N_28081,N_27016,N_27293);
and U28082 (N_28082,N_27164,N_27036);
xor U28083 (N_28083,N_27226,N_27559);
nand U28084 (N_28084,N_27797,N_27409);
xor U28085 (N_28085,N_27441,N_27033);
nor U28086 (N_28086,N_27615,N_27254);
xnor U28087 (N_28087,N_27758,N_27629);
nand U28088 (N_28088,N_27321,N_27012);
nor U28089 (N_28089,N_27131,N_27898);
or U28090 (N_28090,N_27846,N_27375);
and U28091 (N_28091,N_27498,N_27201);
or U28092 (N_28092,N_27111,N_27998);
and U28093 (N_28093,N_27468,N_27249);
nand U28094 (N_28094,N_27655,N_27196);
xor U28095 (N_28095,N_27463,N_27056);
and U28096 (N_28096,N_27340,N_27811);
xor U28097 (N_28097,N_27225,N_27912);
xor U28098 (N_28098,N_27079,N_27608);
and U28099 (N_28099,N_27596,N_27714);
and U28100 (N_28100,N_27609,N_27824);
nand U28101 (N_28101,N_27194,N_27749);
or U28102 (N_28102,N_27435,N_27262);
nand U28103 (N_28103,N_27395,N_27981);
nand U28104 (N_28104,N_27886,N_27582);
nand U28105 (N_28105,N_27212,N_27078);
or U28106 (N_28106,N_27832,N_27518);
nand U28107 (N_28107,N_27881,N_27563);
nor U28108 (N_28108,N_27359,N_27507);
nor U28109 (N_28109,N_27591,N_27837);
xor U28110 (N_28110,N_27800,N_27236);
and U28111 (N_28111,N_27919,N_27580);
and U28112 (N_28112,N_27290,N_27626);
and U28113 (N_28113,N_27738,N_27776);
xor U28114 (N_28114,N_27200,N_27418);
xnor U28115 (N_28115,N_27367,N_27669);
nand U28116 (N_28116,N_27848,N_27555);
nor U28117 (N_28117,N_27852,N_27183);
xnor U28118 (N_28118,N_27777,N_27909);
or U28119 (N_28119,N_27601,N_27386);
xor U28120 (N_28120,N_27940,N_27143);
xor U28121 (N_28121,N_27215,N_27038);
nor U28122 (N_28122,N_27810,N_27007);
xnor U28123 (N_28123,N_27537,N_27316);
and U28124 (N_28124,N_27990,N_27853);
and U28125 (N_28125,N_27731,N_27656);
and U28126 (N_28126,N_27873,N_27126);
nand U28127 (N_28127,N_27527,N_27049);
nand U28128 (N_28128,N_27257,N_27412);
nor U28129 (N_28129,N_27424,N_27581);
nand U28130 (N_28130,N_27792,N_27353);
nand U28131 (N_28131,N_27606,N_27149);
xnor U28132 (N_28132,N_27123,N_27246);
nor U28133 (N_28133,N_27452,N_27357);
or U28134 (N_28134,N_27888,N_27796);
xnor U28135 (N_28135,N_27602,N_27337);
or U28136 (N_28136,N_27611,N_27892);
and U28137 (N_28137,N_27823,N_27607);
and U28138 (N_28138,N_27153,N_27097);
or U28139 (N_28139,N_27160,N_27698);
and U28140 (N_28140,N_27771,N_27190);
xor U28141 (N_28141,N_27906,N_27788);
and U28142 (N_28142,N_27729,N_27774);
nand U28143 (N_28143,N_27821,N_27156);
nor U28144 (N_28144,N_27174,N_27936);
or U28145 (N_28145,N_27222,N_27937);
or U28146 (N_28146,N_27453,N_27429);
nand U28147 (N_28147,N_27289,N_27334);
and U28148 (N_28148,N_27762,N_27380);
nand U28149 (N_28149,N_27266,N_27849);
and U28150 (N_28150,N_27433,N_27805);
xnor U28151 (N_28151,N_27577,N_27673);
nor U28152 (N_28152,N_27371,N_27022);
nand U28153 (N_28153,N_27594,N_27759);
nand U28154 (N_28154,N_27646,N_27182);
nand U28155 (N_28155,N_27166,N_27180);
and U28156 (N_28156,N_27860,N_27532);
or U28157 (N_28157,N_27158,N_27793);
nand U28158 (N_28158,N_27318,N_27206);
and U28159 (N_28159,N_27735,N_27475);
and U28160 (N_28160,N_27769,N_27946);
xnor U28161 (N_28161,N_27017,N_27252);
nand U28162 (N_28162,N_27281,N_27702);
nand U28163 (N_28163,N_27218,N_27426);
nand U28164 (N_28164,N_27263,N_27447);
and U28165 (N_28165,N_27700,N_27941);
nand U28166 (N_28166,N_27711,N_27746);
nand U28167 (N_28167,N_27719,N_27569);
or U28168 (N_28168,N_27736,N_27085);
and U28169 (N_28169,N_27043,N_27491);
xnor U28170 (N_28170,N_27566,N_27819);
xnor U28171 (N_28171,N_27728,N_27460);
nor U28172 (N_28172,N_27094,N_27713);
or U28173 (N_28173,N_27389,N_27726);
xnor U28174 (N_28174,N_27071,N_27457);
nand U28175 (N_28175,N_27640,N_27410);
or U28176 (N_28176,N_27396,N_27233);
nand U28177 (N_28177,N_27349,N_27934);
nor U28178 (N_28178,N_27925,N_27499);
nor U28179 (N_28179,N_27516,N_27031);
nor U28180 (N_28180,N_27818,N_27355);
nand U28181 (N_28181,N_27586,N_27567);
nor U28182 (N_28182,N_27366,N_27270);
or U28183 (N_28183,N_27259,N_27723);
nand U28184 (N_28184,N_27436,N_27061);
nand U28185 (N_28185,N_27670,N_27838);
nand U28186 (N_28186,N_27784,N_27871);
nand U28187 (N_28187,N_27058,N_27220);
xor U28188 (N_28188,N_27961,N_27115);
and U28189 (N_28189,N_27037,N_27029);
and U28190 (N_28190,N_27199,N_27391);
nand U28191 (N_28191,N_27689,N_27637);
or U28192 (N_28192,N_27451,N_27327);
xnor U28193 (N_28193,N_27635,N_27269);
xor U28194 (N_28194,N_27550,N_27323);
nand U28195 (N_28195,N_27945,N_27390);
xnor U28196 (N_28196,N_27630,N_27668);
nand U28197 (N_28197,N_27542,N_27419);
and U28198 (N_28198,N_27084,N_27704);
or U28199 (N_28199,N_27456,N_27991);
and U28200 (N_28200,N_27494,N_27169);
and U28201 (N_28201,N_27055,N_27526);
or U28202 (N_28202,N_27425,N_27423);
xor U28203 (N_28203,N_27652,N_27688);
nor U28204 (N_28204,N_27779,N_27431);
or U28205 (N_28205,N_27277,N_27046);
and U28206 (N_28206,N_27015,N_27387);
and U28207 (N_28207,N_27267,N_27411);
nor U28208 (N_28208,N_27207,N_27151);
xor U28209 (N_28209,N_27090,N_27365);
xnor U28210 (N_28210,N_27968,N_27383);
or U28211 (N_28211,N_27062,N_27059);
and U28212 (N_28212,N_27908,N_27276);
nor U28213 (N_28213,N_27928,N_27644);
or U28214 (N_28214,N_27712,N_27533);
or U28215 (N_28215,N_27248,N_27000);
xnor U28216 (N_28216,N_27659,N_27150);
xor U28217 (N_28217,N_27025,N_27953);
nor U28218 (N_28218,N_27492,N_27756);
xor U28219 (N_28219,N_27787,N_27284);
or U28220 (N_28220,N_27159,N_27872);
xor U28221 (N_28221,N_27978,N_27951);
nor U28222 (N_28222,N_27544,N_27192);
or U28223 (N_28223,N_27127,N_27521);
xor U28224 (N_28224,N_27219,N_27914);
or U28225 (N_28225,N_27610,N_27027);
and U28226 (N_28226,N_27552,N_27761);
xnor U28227 (N_28227,N_27616,N_27146);
or U28228 (N_28228,N_27041,N_27911);
and U28229 (N_28229,N_27685,N_27221);
or U28230 (N_28230,N_27330,N_27278);
xnor U28231 (N_28231,N_27733,N_27891);
nand U28232 (N_28232,N_27579,N_27379);
xnor U28233 (N_28233,N_27144,N_27481);
and U28234 (N_28234,N_27753,N_27750);
or U28235 (N_28235,N_27939,N_27047);
xor U28236 (N_28236,N_27370,N_27496);
nor U28237 (N_28237,N_27165,N_27346);
nand U28238 (N_28238,N_27699,N_27446);
and U28239 (N_28239,N_27623,N_27096);
nand U28240 (N_28240,N_27161,N_27243);
or U28241 (N_28241,N_27322,N_27480);
xnor U28242 (N_28242,N_27617,N_27866);
xor U28243 (N_28243,N_27781,N_27382);
nand U28244 (N_28244,N_27663,N_27910);
nand U28245 (N_28245,N_27343,N_27622);
and U28246 (N_28246,N_27372,N_27798);
nand U28247 (N_28247,N_27665,N_27926);
xnor U28248 (N_28248,N_27922,N_27137);
xnor U28249 (N_28249,N_27405,N_27717);
nor U28250 (N_28250,N_27442,N_27001);
or U28251 (N_28251,N_27690,N_27825);
and U28252 (N_28252,N_27479,N_27209);
nor U28253 (N_28253,N_27013,N_27666);
nand U28254 (N_28254,N_27724,N_27693);
xor U28255 (N_28255,N_27088,N_27109);
nor U28256 (N_28256,N_27264,N_27406);
or U28257 (N_28257,N_27972,N_27965);
and U28258 (N_28258,N_27280,N_27680);
xnor U28259 (N_28259,N_27040,N_27613);
or U28260 (N_28260,N_27009,N_27963);
xnor U28261 (N_28261,N_27184,N_27954);
and U28262 (N_28262,N_27801,N_27984);
nand U28263 (N_28263,N_27850,N_27545);
xnor U28264 (N_28264,N_27145,N_27484);
and U28265 (N_28265,N_27068,N_27363);
or U28266 (N_28266,N_27339,N_27114);
xor U28267 (N_28267,N_27741,N_27708);
and U28268 (N_28268,N_27642,N_27974);
xor U28269 (N_28269,N_27443,N_27268);
xor U28270 (N_28270,N_27006,N_27948);
or U28271 (N_28271,N_27393,N_27234);
nor U28272 (N_28272,N_27979,N_27599);
nor U28273 (N_28273,N_27575,N_27064);
xor U28274 (N_28274,N_27286,N_27345);
or U28275 (N_28275,N_27502,N_27554);
or U28276 (N_28276,N_27999,N_27721);
and U28277 (N_28277,N_27588,N_27335);
or U28278 (N_28278,N_27427,N_27877);
nand U28279 (N_28279,N_27996,N_27661);
nor U28280 (N_28280,N_27767,N_27298);
nor U28281 (N_28281,N_27859,N_27570);
and U28282 (N_28282,N_27147,N_27734);
or U28283 (N_28283,N_27415,N_27732);
xnor U28284 (N_28284,N_27112,N_27328);
nand U28285 (N_28285,N_27506,N_27253);
nor U28286 (N_28286,N_27140,N_27324);
or U28287 (N_28287,N_27154,N_27556);
and U28288 (N_28288,N_27814,N_27101);
xor U28289 (N_28289,N_27224,N_27534);
xor U28290 (N_28290,N_27305,N_27175);
and U28291 (N_28291,N_27439,N_27141);
nand U28292 (N_28292,N_27706,N_27844);
and U28293 (N_28293,N_27639,N_27894);
or U28294 (N_28294,N_27271,N_27966);
nor U28295 (N_28295,N_27074,N_27485);
nand U28296 (N_28296,N_27081,N_27679);
or U28297 (N_28297,N_27030,N_27903);
or U28298 (N_28298,N_27239,N_27210);
and U28299 (N_28299,N_27827,N_27718);
and U28300 (N_28300,N_27362,N_27136);
or U28301 (N_28301,N_27319,N_27907);
nand U28302 (N_28302,N_27102,N_27470);
nand U28303 (N_28303,N_27667,N_27614);
or U28304 (N_28304,N_27634,N_27296);
xnor U28305 (N_28305,N_27603,N_27117);
and U28306 (N_28306,N_27993,N_27476);
nor U28307 (N_28307,N_27631,N_27251);
nor U28308 (N_28308,N_27205,N_27952);
xnor U28309 (N_28309,N_27931,N_27310);
nand U28310 (N_28310,N_27564,N_27132);
and U28311 (N_28311,N_27187,N_27549);
or U28312 (N_28312,N_27560,N_27420);
xor U28313 (N_28313,N_27513,N_27574);
nor U28314 (N_28314,N_27188,N_27923);
and U28315 (N_28315,N_27459,N_27658);
nand U28316 (N_28316,N_27918,N_27287);
or U28317 (N_28317,N_27950,N_27466);
nand U28318 (N_28318,N_27247,N_27710);
xnor U28319 (N_28319,N_27955,N_27794);
nor U28320 (N_28320,N_27947,N_27432);
nand U28321 (N_28321,N_27835,N_27535);
or U28322 (N_28322,N_27490,N_27113);
xnor U28323 (N_28323,N_27867,N_27944);
nor U28324 (N_28324,N_27052,N_27072);
nor U28325 (N_28325,N_27032,N_27959);
and U28326 (N_28326,N_27830,N_27897);
nor U28327 (N_28327,N_27857,N_27775);
or U28328 (N_28328,N_27103,N_27536);
and U28329 (N_28329,N_27807,N_27983);
nand U28330 (N_28330,N_27238,N_27854);
or U28331 (N_28331,N_27282,N_27351);
nor U28332 (N_28332,N_27987,N_27461);
nand U28333 (N_28333,N_27971,N_27314);
or U28334 (N_28334,N_27660,N_27752);
nand U28335 (N_28335,N_27497,N_27478);
or U28336 (N_28336,N_27605,N_27069);
xnor U28337 (N_28337,N_27285,N_27065);
nand U28338 (N_28338,N_27299,N_27815);
nand U28339 (N_28339,N_27394,N_27845);
nor U28340 (N_28340,N_27932,N_27336);
nor U28341 (N_28341,N_27657,N_27590);
and U28342 (N_28342,N_27501,N_27977);
nand U28343 (N_28343,N_27011,N_27551);
and U28344 (N_28344,N_27802,N_27026);
and U28345 (N_28345,N_27408,N_27163);
xor U28346 (N_28346,N_27157,N_27045);
xor U28347 (N_28347,N_27933,N_27847);
and U28348 (N_28348,N_27235,N_27373);
xor U28349 (N_28349,N_27471,N_27524);
or U28350 (N_28350,N_27530,N_27080);
xnor U28351 (N_28351,N_27633,N_27073);
xnor U28352 (N_28352,N_27529,N_27486);
and U28353 (N_28353,N_27697,N_27986);
and U28354 (N_28354,N_27110,N_27691);
and U28355 (N_28355,N_27817,N_27350);
nand U28356 (N_28356,N_27618,N_27469);
or U28357 (N_28357,N_27745,N_27091);
and U28358 (N_28358,N_27186,N_27116);
nand U28359 (N_28359,N_27976,N_27956);
or U28360 (N_28360,N_27924,N_27014);
nand U28361 (N_28361,N_27356,N_27326);
and U28362 (N_28362,N_27044,N_27988);
xnor U28363 (N_28363,N_27921,N_27177);
xor U28364 (N_28364,N_27295,N_27901);
xor U28365 (N_28365,N_27782,N_27211);
nand U28366 (N_28366,N_27325,N_27511);
nor U28367 (N_28367,N_27399,N_27883);
xnor U28368 (N_28368,N_27035,N_27645);
nand U28369 (N_28369,N_27258,N_27508);
nor U28370 (N_28370,N_27543,N_27294);
and U28371 (N_28371,N_27005,N_27315);
xnor U28372 (N_28372,N_27216,N_27313);
or U28373 (N_28373,N_27317,N_27764);
xnor U28374 (N_28374,N_27806,N_27089);
nor U28375 (N_28375,N_27755,N_27135);
and U28376 (N_28376,N_27076,N_27002);
nor U28377 (N_28377,N_27067,N_27768);
xor U28378 (N_28378,N_27573,N_27256);
xnor U28379 (N_28379,N_27152,N_27565);
or U28380 (N_28380,N_27381,N_27348);
or U28381 (N_28381,N_27308,N_27487);
or U28382 (N_28382,N_27651,N_27473);
xor U28383 (N_28383,N_27275,N_27230);
nand U28384 (N_28384,N_27333,N_27329);
and U28385 (N_28385,N_27523,N_27650);
nand U28386 (N_28386,N_27274,N_27561);
or U28387 (N_28387,N_27539,N_27757);
or U28388 (N_28388,N_27856,N_27377);
xnor U28389 (N_28389,N_27232,N_27139);
and U28390 (N_28390,N_27428,N_27493);
or U28391 (N_28391,N_27019,N_27142);
or U28392 (N_28392,N_27528,N_27982);
nor U28393 (N_28393,N_27705,N_27638);
xnor U28394 (N_28394,N_27870,N_27307);
nand U28395 (N_28395,N_27522,N_27747);
and U28396 (N_28396,N_27812,N_27973);
nand U28397 (N_28397,N_27636,N_27213);
xor U28398 (N_28398,N_27170,N_27283);
and U28399 (N_28399,N_27869,N_27541);
or U28400 (N_28400,N_27107,N_27703);
or U28401 (N_28401,N_27942,N_27272);
and U28402 (N_28402,N_27730,N_27240);
nor U28403 (N_28403,N_27748,N_27843);
or U28404 (N_28404,N_27483,N_27595);
xor U28405 (N_28405,N_27054,N_27831);
nor U28406 (N_28406,N_27244,N_27376);
nor U28407 (N_28407,N_27677,N_27967);
or U28408 (N_28408,N_27740,N_27155);
or U28409 (N_28409,N_27168,N_27861);
nand U28410 (N_28410,N_27401,N_27416);
xnor U28411 (N_28411,N_27664,N_27197);
xor U28412 (N_28412,N_27051,N_27772);
and U28413 (N_28413,N_27509,N_27836);
nor U28414 (N_28414,N_27620,N_27833);
and U28415 (N_28415,N_27515,N_27520);
nand U28416 (N_28416,N_27173,N_27695);
and U28417 (N_28417,N_27417,N_27900);
xor U28418 (N_28418,N_27082,N_27727);
nor U28419 (N_28419,N_27905,N_27407);
and U28420 (N_28420,N_27514,N_27010);
and U28421 (N_28421,N_27879,N_27902);
and U28422 (N_28422,N_27422,N_27414);
nand U28423 (N_28423,N_27223,N_27042);
nor U28424 (N_28424,N_27179,N_27739);
or U28425 (N_28425,N_27495,N_27694);
nor U28426 (N_28426,N_27504,N_27851);
and U28427 (N_28427,N_27548,N_27347);
xnor U28428 (N_28428,N_27773,N_27392);
and U28429 (N_28429,N_27465,N_27930);
or U28430 (N_28430,N_27632,N_27662);
or U28431 (N_28431,N_27312,N_27378);
nand U28432 (N_28432,N_27589,N_27682);
or U28433 (N_28433,N_27822,N_27783);
nor U28434 (N_28434,N_27130,N_27304);
or U28435 (N_28435,N_27820,N_27929);
nand U28436 (N_28436,N_27403,N_27619);
or U28437 (N_28437,N_27265,N_27204);
nand U28438 (N_28438,N_27826,N_27048);
and U28439 (N_28439,N_27095,N_27687);
xnor U28440 (N_28440,N_27231,N_27352);
or U28441 (N_28441,N_27203,N_27789);
nand U28442 (N_28442,N_27106,N_27546);
and U28443 (N_28443,N_27120,N_27531);
nand U28444 (N_28444,N_27553,N_27790);
xor U28445 (N_28445,N_27134,N_27060);
xnor U28446 (N_28446,N_27884,N_27558);
xnor U28447 (N_28447,N_27880,N_27980);
and U28448 (N_28448,N_27291,N_27128);
and U28449 (N_28449,N_27472,N_27039);
or U28450 (N_28450,N_27402,N_27868);
nand U28451 (N_28451,N_27874,N_27675);
or U28452 (N_28452,N_27214,N_27743);
nand U28453 (N_28453,N_27034,N_27242);
nor U28454 (N_28454,N_27557,N_27654);
and U28455 (N_28455,N_27129,N_27992);
or U28456 (N_28456,N_27786,N_27828);
nor U28457 (N_28457,N_27021,N_27087);
or U28458 (N_28458,N_27957,N_27813);
and U28459 (N_28459,N_27489,N_27250);
and U28460 (N_28460,N_27686,N_27467);
nand U28461 (N_28461,N_27648,N_27437);
nand U28462 (N_28462,N_27899,N_27766);
nor U28463 (N_28463,N_27237,N_27780);
nand U28464 (N_28464,N_27162,N_27385);
xnor U28465 (N_28465,N_27241,N_27785);
or U28466 (N_28466,N_27125,N_27066);
xnor U28467 (N_28467,N_27261,N_27625);
nand U28468 (N_28468,N_27969,N_27464);
xnor U28469 (N_28469,N_27344,N_27916);
nor U28470 (N_28470,N_27600,N_27641);
nor U28471 (N_28471,N_27653,N_27092);
nor U28472 (N_28472,N_27448,N_27279);
nand U28473 (N_28473,N_27202,N_27519);
or U28474 (N_28474,N_27896,N_27808);
nor U28475 (N_28475,N_27302,N_27075);
or U28476 (N_28476,N_27191,N_27003);
xor U28477 (N_28477,N_27568,N_27572);
nor U28478 (N_28478,N_27855,N_27260);
nor U28479 (N_28479,N_27882,N_27292);
and U28480 (N_28480,N_27889,N_27621);
nor U28481 (N_28481,N_27217,N_27583);
nor U28482 (N_28482,N_27108,N_27368);
xnor U28483 (N_28483,N_27008,N_27300);
and U28484 (N_28484,N_27301,N_27970);
and U28485 (N_28485,N_27454,N_27440);
nand U28486 (N_28486,N_27913,N_27742);
nand U28487 (N_28487,N_27604,N_27647);
or U28488 (N_28488,N_27482,N_27893);
and U28489 (N_28489,N_27935,N_27404);
or U28490 (N_28490,N_27878,N_27720);
xor U28491 (N_28491,N_27229,N_27384);
xor U28492 (N_28492,N_27400,N_27920);
or U28493 (N_28493,N_27228,N_27737);
xnor U28494 (N_28494,N_27306,N_27863);
xor U28495 (N_28495,N_27795,N_27083);
nor U28496 (N_28496,N_27445,N_27189);
or U28497 (N_28497,N_27462,N_27540);
xnor U28498 (N_28498,N_27364,N_27754);
and U28499 (N_28499,N_27004,N_27585);
nor U28500 (N_28500,N_27110,N_27137);
nor U28501 (N_28501,N_27748,N_27061);
and U28502 (N_28502,N_27018,N_27670);
or U28503 (N_28503,N_27613,N_27811);
nand U28504 (N_28504,N_27578,N_27661);
and U28505 (N_28505,N_27558,N_27098);
or U28506 (N_28506,N_27820,N_27337);
or U28507 (N_28507,N_27969,N_27210);
and U28508 (N_28508,N_27639,N_27863);
nor U28509 (N_28509,N_27102,N_27953);
nand U28510 (N_28510,N_27716,N_27990);
or U28511 (N_28511,N_27246,N_27181);
xnor U28512 (N_28512,N_27294,N_27364);
or U28513 (N_28513,N_27636,N_27221);
nor U28514 (N_28514,N_27078,N_27379);
and U28515 (N_28515,N_27112,N_27896);
nor U28516 (N_28516,N_27188,N_27568);
nand U28517 (N_28517,N_27180,N_27514);
and U28518 (N_28518,N_27486,N_27824);
nor U28519 (N_28519,N_27248,N_27402);
and U28520 (N_28520,N_27318,N_27604);
nand U28521 (N_28521,N_27046,N_27478);
or U28522 (N_28522,N_27652,N_27935);
nor U28523 (N_28523,N_27914,N_27208);
nand U28524 (N_28524,N_27955,N_27222);
or U28525 (N_28525,N_27071,N_27418);
nor U28526 (N_28526,N_27135,N_27842);
and U28527 (N_28527,N_27642,N_27288);
xnor U28528 (N_28528,N_27321,N_27740);
and U28529 (N_28529,N_27410,N_27605);
nor U28530 (N_28530,N_27854,N_27249);
xnor U28531 (N_28531,N_27980,N_27158);
xnor U28532 (N_28532,N_27669,N_27985);
nor U28533 (N_28533,N_27760,N_27370);
xor U28534 (N_28534,N_27652,N_27675);
or U28535 (N_28535,N_27312,N_27540);
and U28536 (N_28536,N_27245,N_27585);
xnor U28537 (N_28537,N_27064,N_27411);
xor U28538 (N_28538,N_27025,N_27671);
and U28539 (N_28539,N_27859,N_27280);
or U28540 (N_28540,N_27533,N_27339);
and U28541 (N_28541,N_27531,N_27263);
nand U28542 (N_28542,N_27725,N_27567);
nor U28543 (N_28543,N_27397,N_27147);
nor U28544 (N_28544,N_27830,N_27505);
nor U28545 (N_28545,N_27506,N_27062);
xnor U28546 (N_28546,N_27223,N_27312);
nand U28547 (N_28547,N_27988,N_27030);
or U28548 (N_28548,N_27121,N_27009);
or U28549 (N_28549,N_27860,N_27775);
nor U28550 (N_28550,N_27250,N_27219);
and U28551 (N_28551,N_27247,N_27578);
xnor U28552 (N_28552,N_27457,N_27124);
or U28553 (N_28553,N_27865,N_27262);
and U28554 (N_28554,N_27431,N_27714);
xor U28555 (N_28555,N_27072,N_27561);
nand U28556 (N_28556,N_27304,N_27455);
nand U28557 (N_28557,N_27457,N_27770);
and U28558 (N_28558,N_27250,N_27187);
and U28559 (N_28559,N_27834,N_27505);
nand U28560 (N_28560,N_27172,N_27681);
xnor U28561 (N_28561,N_27521,N_27993);
nor U28562 (N_28562,N_27915,N_27960);
nor U28563 (N_28563,N_27170,N_27131);
and U28564 (N_28564,N_27025,N_27850);
and U28565 (N_28565,N_27213,N_27890);
nor U28566 (N_28566,N_27528,N_27728);
nand U28567 (N_28567,N_27211,N_27486);
and U28568 (N_28568,N_27117,N_27225);
nand U28569 (N_28569,N_27017,N_27244);
xor U28570 (N_28570,N_27869,N_27163);
and U28571 (N_28571,N_27737,N_27515);
xor U28572 (N_28572,N_27252,N_27343);
nor U28573 (N_28573,N_27836,N_27414);
or U28574 (N_28574,N_27756,N_27942);
nand U28575 (N_28575,N_27066,N_27081);
xor U28576 (N_28576,N_27657,N_27358);
or U28577 (N_28577,N_27915,N_27283);
nor U28578 (N_28578,N_27803,N_27725);
xnor U28579 (N_28579,N_27350,N_27696);
or U28580 (N_28580,N_27855,N_27651);
and U28581 (N_28581,N_27279,N_27610);
and U28582 (N_28582,N_27424,N_27743);
nand U28583 (N_28583,N_27132,N_27593);
xor U28584 (N_28584,N_27750,N_27604);
nor U28585 (N_28585,N_27387,N_27294);
nand U28586 (N_28586,N_27536,N_27960);
and U28587 (N_28587,N_27926,N_27140);
or U28588 (N_28588,N_27691,N_27338);
nor U28589 (N_28589,N_27318,N_27117);
xor U28590 (N_28590,N_27167,N_27275);
xnor U28591 (N_28591,N_27596,N_27099);
or U28592 (N_28592,N_27907,N_27378);
xor U28593 (N_28593,N_27597,N_27840);
or U28594 (N_28594,N_27966,N_27290);
and U28595 (N_28595,N_27393,N_27968);
xor U28596 (N_28596,N_27716,N_27015);
nor U28597 (N_28597,N_27908,N_27845);
xnor U28598 (N_28598,N_27320,N_27692);
nand U28599 (N_28599,N_27139,N_27072);
nor U28600 (N_28600,N_27506,N_27364);
and U28601 (N_28601,N_27634,N_27287);
nand U28602 (N_28602,N_27455,N_27600);
and U28603 (N_28603,N_27144,N_27838);
nand U28604 (N_28604,N_27598,N_27621);
xor U28605 (N_28605,N_27376,N_27642);
xor U28606 (N_28606,N_27615,N_27589);
or U28607 (N_28607,N_27815,N_27327);
nand U28608 (N_28608,N_27367,N_27162);
nor U28609 (N_28609,N_27268,N_27791);
or U28610 (N_28610,N_27901,N_27151);
nor U28611 (N_28611,N_27742,N_27044);
or U28612 (N_28612,N_27842,N_27332);
nand U28613 (N_28613,N_27532,N_27189);
xnor U28614 (N_28614,N_27744,N_27863);
nor U28615 (N_28615,N_27853,N_27522);
or U28616 (N_28616,N_27620,N_27087);
and U28617 (N_28617,N_27534,N_27908);
nand U28618 (N_28618,N_27456,N_27451);
xor U28619 (N_28619,N_27260,N_27750);
or U28620 (N_28620,N_27819,N_27375);
nand U28621 (N_28621,N_27747,N_27686);
nand U28622 (N_28622,N_27709,N_27486);
nor U28623 (N_28623,N_27747,N_27511);
or U28624 (N_28624,N_27271,N_27096);
and U28625 (N_28625,N_27594,N_27481);
nor U28626 (N_28626,N_27788,N_27568);
xor U28627 (N_28627,N_27227,N_27749);
nor U28628 (N_28628,N_27234,N_27485);
nand U28629 (N_28629,N_27750,N_27439);
or U28630 (N_28630,N_27734,N_27213);
nand U28631 (N_28631,N_27393,N_27240);
nor U28632 (N_28632,N_27242,N_27318);
nand U28633 (N_28633,N_27443,N_27840);
or U28634 (N_28634,N_27433,N_27749);
nor U28635 (N_28635,N_27716,N_27327);
xnor U28636 (N_28636,N_27501,N_27076);
xor U28637 (N_28637,N_27555,N_27085);
xor U28638 (N_28638,N_27389,N_27197);
or U28639 (N_28639,N_27645,N_27979);
xor U28640 (N_28640,N_27294,N_27185);
nor U28641 (N_28641,N_27161,N_27963);
and U28642 (N_28642,N_27472,N_27217);
nor U28643 (N_28643,N_27354,N_27678);
or U28644 (N_28644,N_27325,N_27436);
nand U28645 (N_28645,N_27964,N_27298);
xnor U28646 (N_28646,N_27483,N_27405);
nand U28647 (N_28647,N_27051,N_27674);
or U28648 (N_28648,N_27318,N_27625);
xor U28649 (N_28649,N_27750,N_27896);
nor U28650 (N_28650,N_27717,N_27957);
nor U28651 (N_28651,N_27426,N_27521);
nor U28652 (N_28652,N_27458,N_27528);
nor U28653 (N_28653,N_27372,N_27318);
or U28654 (N_28654,N_27891,N_27087);
xnor U28655 (N_28655,N_27930,N_27252);
nor U28656 (N_28656,N_27627,N_27969);
nor U28657 (N_28657,N_27026,N_27279);
and U28658 (N_28658,N_27191,N_27341);
nand U28659 (N_28659,N_27926,N_27458);
or U28660 (N_28660,N_27286,N_27357);
xnor U28661 (N_28661,N_27568,N_27928);
nand U28662 (N_28662,N_27274,N_27225);
nor U28663 (N_28663,N_27096,N_27491);
or U28664 (N_28664,N_27387,N_27883);
or U28665 (N_28665,N_27650,N_27570);
and U28666 (N_28666,N_27142,N_27335);
or U28667 (N_28667,N_27880,N_27989);
xor U28668 (N_28668,N_27284,N_27426);
or U28669 (N_28669,N_27075,N_27594);
and U28670 (N_28670,N_27140,N_27418);
and U28671 (N_28671,N_27817,N_27139);
nor U28672 (N_28672,N_27296,N_27452);
or U28673 (N_28673,N_27139,N_27399);
or U28674 (N_28674,N_27951,N_27191);
nor U28675 (N_28675,N_27644,N_27473);
nand U28676 (N_28676,N_27116,N_27795);
and U28677 (N_28677,N_27176,N_27370);
or U28678 (N_28678,N_27851,N_27953);
or U28679 (N_28679,N_27964,N_27500);
xor U28680 (N_28680,N_27036,N_27342);
nor U28681 (N_28681,N_27212,N_27187);
xnor U28682 (N_28682,N_27563,N_27759);
xnor U28683 (N_28683,N_27374,N_27283);
and U28684 (N_28684,N_27994,N_27428);
or U28685 (N_28685,N_27071,N_27795);
xnor U28686 (N_28686,N_27295,N_27068);
nand U28687 (N_28687,N_27361,N_27518);
nor U28688 (N_28688,N_27912,N_27430);
or U28689 (N_28689,N_27723,N_27667);
and U28690 (N_28690,N_27379,N_27562);
or U28691 (N_28691,N_27664,N_27413);
nor U28692 (N_28692,N_27375,N_27029);
xor U28693 (N_28693,N_27536,N_27582);
nand U28694 (N_28694,N_27473,N_27953);
or U28695 (N_28695,N_27558,N_27615);
and U28696 (N_28696,N_27708,N_27218);
xnor U28697 (N_28697,N_27469,N_27737);
and U28698 (N_28698,N_27588,N_27843);
and U28699 (N_28699,N_27196,N_27039);
nand U28700 (N_28700,N_27947,N_27004);
nor U28701 (N_28701,N_27743,N_27115);
nand U28702 (N_28702,N_27378,N_27059);
and U28703 (N_28703,N_27160,N_27947);
and U28704 (N_28704,N_27675,N_27846);
nand U28705 (N_28705,N_27184,N_27743);
xor U28706 (N_28706,N_27487,N_27322);
nor U28707 (N_28707,N_27444,N_27678);
nand U28708 (N_28708,N_27537,N_27298);
nand U28709 (N_28709,N_27510,N_27640);
or U28710 (N_28710,N_27718,N_27276);
xnor U28711 (N_28711,N_27028,N_27763);
and U28712 (N_28712,N_27469,N_27727);
or U28713 (N_28713,N_27932,N_27142);
and U28714 (N_28714,N_27904,N_27486);
xnor U28715 (N_28715,N_27060,N_27532);
xnor U28716 (N_28716,N_27949,N_27116);
nand U28717 (N_28717,N_27812,N_27728);
nand U28718 (N_28718,N_27779,N_27650);
nor U28719 (N_28719,N_27446,N_27238);
xor U28720 (N_28720,N_27865,N_27683);
nor U28721 (N_28721,N_27512,N_27349);
xnor U28722 (N_28722,N_27508,N_27504);
nand U28723 (N_28723,N_27017,N_27079);
nand U28724 (N_28724,N_27331,N_27809);
nand U28725 (N_28725,N_27175,N_27493);
nand U28726 (N_28726,N_27733,N_27493);
nand U28727 (N_28727,N_27734,N_27874);
nor U28728 (N_28728,N_27615,N_27238);
and U28729 (N_28729,N_27834,N_27984);
xor U28730 (N_28730,N_27218,N_27990);
or U28731 (N_28731,N_27822,N_27336);
or U28732 (N_28732,N_27155,N_27581);
and U28733 (N_28733,N_27058,N_27069);
and U28734 (N_28734,N_27968,N_27651);
or U28735 (N_28735,N_27799,N_27863);
xor U28736 (N_28736,N_27858,N_27887);
xor U28737 (N_28737,N_27071,N_27232);
nor U28738 (N_28738,N_27936,N_27034);
nand U28739 (N_28739,N_27494,N_27789);
and U28740 (N_28740,N_27942,N_27904);
nor U28741 (N_28741,N_27148,N_27458);
xor U28742 (N_28742,N_27087,N_27267);
and U28743 (N_28743,N_27393,N_27659);
or U28744 (N_28744,N_27297,N_27743);
or U28745 (N_28745,N_27049,N_27867);
and U28746 (N_28746,N_27895,N_27319);
nand U28747 (N_28747,N_27802,N_27662);
and U28748 (N_28748,N_27762,N_27856);
or U28749 (N_28749,N_27192,N_27160);
nor U28750 (N_28750,N_27222,N_27881);
nand U28751 (N_28751,N_27197,N_27041);
nand U28752 (N_28752,N_27233,N_27828);
nand U28753 (N_28753,N_27324,N_27188);
and U28754 (N_28754,N_27854,N_27446);
xor U28755 (N_28755,N_27291,N_27058);
nand U28756 (N_28756,N_27914,N_27989);
and U28757 (N_28757,N_27417,N_27293);
xor U28758 (N_28758,N_27425,N_27900);
or U28759 (N_28759,N_27770,N_27110);
xnor U28760 (N_28760,N_27414,N_27951);
or U28761 (N_28761,N_27332,N_27771);
xnor U28762 (N_28762,N_27300,N_27053);
nand U28763 (N_28763,N_27406,N_27408);
nand U28764 (N_28764,N_27769,N_27223);
or U28765 (N_28765,N_27442,N_27709);
nand U28766 (N_28766,N_27155,N_27230);
nand U28767 (N_28767,N_27697,N_27173);
nor U28768 (N_28768,N_27643,N_27455);
nand U28769 (N_28769,N_27137,N_27937);
nand U28770 (N_28770,N_27901,N_27919);
or U28771 (N_28771,N_27565,N_27059);
and U28772 (N_28772,N_27259,N_27100);
xor U28773 (N_28773,N_27092,N_27042);
nand U28774 (N_28774,N_27066,N_27965);
and U28775 (N_28775,N_27550,N_27666);
and U28776 (N_28776,N_27216,N_27179);
or U28777 (N_28777,N_27927,N_27311);
and U28778 (N_28778,N_27379,N_27805);
nand U28779 (N_28779,N_27888,N_27934);
or U28780 (N_28780,N_27612,N_27180);
and U28781 (N_28781,N_27795,N_27017);
and U28782 (N_28782,N_27792,N_27653);
and U28783 (N_28783,N_27387,N_27921);
nor U28784 (N_28784,N_27882,N_27197);
nand U28785 (N_28785,N_27994,N_27617);
and U28786 (N_28786,N_27112,N_27606);
and U28787 (N_28787,N_27705,N_27451);
and U28788 (N_28788,N_27325,N_27215);
xor U28789 (N_28789,N_27397,N_27701);
xor U28790 (N_28790,N_27899,N_27297);
xor U28791 (N_28791,N_27214,N_27229);
xor U28792 (N_28792,N_27189,N_27188);
and U28793 (N_28793,N_27945,N_27930);
nor U28794 (N_28794,N_27979,N_27232);
nor U28795 (N_28795,N_27515,N_27070);
and U28796 (N_28796,N_27050,N_27633);
and U28797 (N_28797,N_27963,N_27929);
or U28798 (N_28798,N_27625,N_27057);
or U28799 (N_28799,N_27818,N_27844);
and U28800 (N_28800,N_27696,N_27126);
xor U28801 (N_28801,N_27866,N_27678);
and U28802 (N_28802,N_27949,N_27279);
xnor U28803 (N_28803,N_27343,N_27171);
or U28804 (N_28804,N_27405,N_27370);
and U28805 (N_28805,N_27495,N_27898);
and U28806 (N_28806,N_27489,N_27665);
nand U28807 (N_28807,N_27373,N_27245);
and U28808 (N_28808,N_27128,N_27398);
nand U28809 (N_28809,N_27389,N_27908);
and U28810 (N_28810,N_27974,N_27915);
nor U28811 (N_28811,N_27324,N_27167);
or U28812 (N_28812,N_27459,N_27362);
or U28813 (N_28813,N_27524,N_27883);
xnor U28814 (N_28814,N_27613,N_27662);
nand U28815 (N_28815,N_27331,N_27439);
xnor U28816 (N_28816,N_27697,N_27912);
nand U28817 (N_28817,N_27012,N_27237);
xnor U28818 (N_28818,N_27996,N_27858);
and U28819 (N_28819,N_27266,N_27416);
nand U28820 (N_28820,N_27780,N_27268);
and U28821 (N_28821,N_27134,N_27767);
nor U28822 (N_28822,N_27570,N_27008);
xor U28823 (N_28823,N_27589,N_27371);
nand U28824 (N_28824,N_27048,N_27439);
nor U28825 (N_28825,N_27203,N_27195);
or U28826 (N_28826,N_27066,N_27121);
xnor U28827 (N_28827,N_27480,N_27368);
and U28828 (N_28828,N_27650,N_27008);
nor U28829 (N_28829,N_27735,N_27089);
and U28830 (N_28830,N_27241,N_27603);
and U28831 (N_28831,N_27769,N_27607);
xnor U28832 (N_28832,N_27750,N_27319);
and U28833 (N_28833,N_27745,N_27592);
and U28834 (N_28834,N_27019,N_27689);
and U28835 (N_28835,N_27770,N_27950);
nor U28836 (N_28836,N_27525,N_27139);
nor U28837 (N_28837,N_27994,N_27047);
or U28838 (N_28838,N_27097,N_27662);
nand U28839 (N_28839,N_27171,N_27966);
nor U28840 (N_28840,N_27112,N_27462);
xor U28841 (N_28841,N_27052,N_27029);
nor U28842 (N_28842,N_27994,N_27747);
or U28843 (N_28843,N_27152,N_27487);
or U28844 (N_28844,N_27864,N_27330);
nand U28845 (N_28845,N_27049,N_27209);
xnor U28846 (N_28846,N_27911,N_27352);
or U28847 (N_28847,N_27058,N_27518);
nand U28848 (N_28848,N_27064,N_27256);
nor U28849 (N_28849,N_27946,N_27953);
xnor U28850 (N_28850,N_27650,N_27614);
nor U28851 (N_28851,N_27445,N_27317);
or U28852 (N_28852,N_27156,N_27394);
or U28853 (N_28853,N_27101,N_27588);
or U28854 (N_28854,N_27381,N_27869);
xnor U28855 (N_28855,N_27578,N_27603);
or U28856 (N_28856,N_27970,N_27791);
nand U28857 (N_28857,N_27912,N_27778);
and U28858 (N_28858,N_27595,N_27633);
nor U28859 (N_28859,N_27565,N_27204);
or U28860 (N_28860,N_27939,N_27172);
xor U28861 (N_28861,N_27632,N_27986);
nor U28862 (N_28862,N_27912,N_27203);
nor U28863 (N_28863,N_27447,N_27664);
xnor U28864 (N_28864,N_27090,N_27476);
nand U28865 (N_28865,N_27534,N_27199);
nand U28866 (N_28866,N_27121,N_27473);
or U28867 (N_28867,N_27638,N_27510);
xnor U28868 (N_28868,N_27609,N_27092);
nor U28869 (N_28869,N_27848,N_27652);
nand U28870 (N_28870,N_27415,N_27986);
and U28871 (N_28871,N_27824,N_27755);
or U28872 (N_28872,N_27566,N_27754);
or U28873 (N_28873,N_27682,N_27571);
nand U28874 (N_28874,N_27924,N_27115);
xor U28875 (N_28875,N_27102,N_27370);
nor U28876 (N_28876,N_27336,N_27694);
and U28877 (N_28877,N_27675,N_27765);
nor U28878 (N_28878,N_27294,N_27127);
nor U28879 (N_28879,N_27883,N_27158);
xnor U28880 (N_28880,N_27197,N_27829);
nor U28881 (N_28881,N_27304,N_27430);
nor U28882 (N_28882,N_27556,N_27026);
or U28883 (N_28883,N_27365,N_27531);
xor U28884 (N_28884,N_27960,N_27105);
or U28885 (N_28885,N_27249,N_27166);
and U28886 (N_28886,N_27612,N_27301);
and U28887 (N_28887,N_27896,N_27693);
nand U28888 (N_28888,N_27671,N_27836);
xnor U28889 (N_28889,N_27160,N_27057);
nor U28890 (N_28890,N_27305,N_27955);
or U28891 (N_28891,N_27494,N_27629);
xnor U28892 (N_28892,N_27164,N_27037);
nor U28893 (N_28893,N_27633,N_27724);
nand U28894 (N_28894,N_27407,N_27115);
and U28895 (N_28895,N_27848,N_27720);
nand U28896 (N_28896,N_27284,N_27950);
nand U28897 (N_28897,N_27994,N_27533);
nand U28898 (N_28898,N_27007,N_27958);
or U28899 (N_28899,N_27102,N_27561);
and U28900 (N_28900,N_27819,N_27926);
or U28901 (N_28901,N_27417,N_27749);
and U28902 (N_28902,N_27821,N_27839);
xnor U28903 (N_28903,N_27528,N_27182);
or U28904 (N_28904,N_27369,N_27606);
nor U28905 (N_28905,N_27319,N_27006);
or U28906 (N_28906,N_27308,N_27146);
and U28907 (N_28907,N_27757,N_27035);
and U28908 (N_28908,N_27450,N_27088);
or U28909 (N_28909,N_27138,N_27357);
or U28910 (N_28910,N_27657,N_27317);
nor U28911 (N_28911,N_27687,N_27789);
and U28912 (N_28912,N_27490,N_27469);
or U28913 (N_28913,N_27522,N_27294);
or U28914 (N_28914,N_27484,N_27766);
and U28915 (N_28915,N_27453,N_27169);
nand U28916 (N_28916,N_27691,N_27856);
or U28917 (N_28917,N_27610,N_27776);
nand U28918 (N_28918,N_27239,N_27056);
xnor U28919 (N_28919,N_27179,N_27933);
or U28920 (N_28920,N_27007,N_27086);
xor U28921 (N_28921,N_27282,N_27808);
or U28922 (N_28922,N_27935,N_27266);
nand U28923 (N_28923,N_27185,N_27688);
xor U28924 (N_28924,N_27454,N_27390);
or U28925 (N_28925,N_27375,N_27847);
xnor U28926 (N_28926,N_27858,N_27580);
nand U28927 (N_28927,N_27509,N_27847);
nor U28928 (N_28928,N_27537,N_27437);
or U28929 (N_28929,N_27315,N_27712);
and U28930 (N_28930,N_27492,N_27277);
and U28931 (N_28931,N_27378,N_27938);
nor U28932 (N_28932,N_27796,N_27503);
or U28933 (N_28933,N_27063,N_27406);
or U28934 (N_28934,N_27214,N_27641);
xor U28935 (N_28935,N_27178,N_27409);
nand U28936 (N_28936,N_27594,N_27341);
xnor U28937 (N_28937,N_27960,N_27734);
nand U28938 (N_28938,N_27236,N_27595);
xor U28939 (N_28939,N_27816,N_27645);
xor U28940 (N_28940,N_27383,N_27354);
nor U28941 (N_28941,N_27343,N_27958);
nor U28942 (N_28942,N_27718,N_27485);
or U28943 (N_28943,N_27368,N_27349);
nor U28944 (N_28944,N_27633,N_27042);
or U28945 (N_28945,N_27490,N_27270);
and U28946 (N_28946,N_27032,N_27035);
xnor U28947 (N_28947,N_27144,N_27737);
nor U28948 (N_28948,N_27676,N_27990);
nor U28949 (N_28949,N_27459,N_27869);
or U28950 (N_28950,N_27455,N_27589);
nor U28951 (N_28951,N_27787,N_27719);
or U28952 (N_28952,N_27439,N_27590);
nand U28953 (N_28953,N_27786,N_27097);
nor U28954 (N_28954,N_27022,N_27100);
xor U28955 (N_28955,N_27280,N_27061);
and U28956 (N_28956,N_27258,N_27037);
nand U28957 (N_28957,N_27397,N_27539);
nand U28958 (N_28958,N_27298,N_27468);
and U28959 (N_28959,N_27311,N_27598);
or U28960 (N_28960,N_27403,N_27570);
and U28961 (N_28961,N_27061,N_27959);
nor U28962 (N_28962,N_27290,N_27300);
nor U28963 (N_28963,N_27499,N_27600);
nand U28964 (N_28964,N_27530,N_27147);
or U28965 (N_28965,N_27282,N_27625);
and U28966 (N_28966,N_27462,N_27429);
nand U28967 (N_28967,N_27886,N_27774);
xor U28968 (N_28968,N_27113,N_27806);
nor U28969 (N_28969,N_27972,N_27268);
nor U28970 (N_28970,N_27861,N_27850);
and U28971 (N_28971,N_27760,N_27068);
nand U28972 (N_28972,N_27085,N_27702);
nor U28973 (N_28973,N_27450,N_27172);
xor U28974 (N_28974,N_27814,N_27632);
nor U28975 (N_28975,N_27013,N_27782);
and U28976 (N_28976,N_27616,N_27990);
or U28977 (N_28977,N_27561,N_27658);
nand U28978 (N_28978,N_27335,N_27482);
nand U28979 (N_28979,N_27630,N_27411);
xor U28980 (N_28980,N_27381,N_27866);
nand U28981 (N_28981,N_27493,N_27967);
nor U28982 (N_28982,N_27894,N_27945);
and U28983 (N_28983,N_27874,N_27610);
and U28984 (N_28984,N_27842,N_27513);
or U28985 (N_28985,N_27042,N_27239);
xor U28986 (N_28986,N_27736,N_27320);
or U28987 (N_28987,N_27700,N_27263);
nor U28988 (N_28988,N_27585,N_27587);
and U28989 (N_28989,N_27337,N_27063);
and U28990 (N_28990,N_27040,N_27992);
nor U28991 (N_28991,N_27151,N_27992);
xnor U28992 (N_28992,N_27051,N_27531);
nand U28993 (N_28993,N_27263,N_27115);
or U28994 (N_28994,N_27916,N_27438);
nand U28995 (N_28995,N_27897,N_27697);
nand U28996 (N_28996,N_27046,N_27496);
nor U28997 (N_28997,N_27761,N_27852);
and U28998 (N_28998,N_27801,N_27720);
or U28999 (N_28999,N_27126,N_27667);
nor U29000 (N_29000,N_28398,N_28781);
and U29001 (N_29001,N_28024,N_28451);
nor U29002 (N_29002,N_28165,N_28225);
and U29003 (N_29003,N_28906,N_28306);
or U29004 (N_29004,N_28933,N_28517);
nand U29005 (N_29005,N_28394,N_28077);
nand U29006 (N_29006,N_28673,N_28229);
xor U29007 (N_29007,N_28195,N_28094);
and U29008 (N_29008,N_28827,N_28824);
nand U29009 (N_29009,N_28053,N_28025);
nor U29010 (N_29010,N_28262,N_28426);
nor U29011 (N_29011,N_28898,N_28360);
nor U29012 (N_29012,N_28457,N_28694);
and U29013 (N_29013,N_28779,N_28632);
xor U29014 (N_29014,N_28159,N_28459);
nor U29015 (N_29015,N_28331,N_28812);
xor U29016 (N_29016,N_28819,N_28961);
nor U29017 (N_29017,N_28402,N_28874);
and U29018 (N_29018,N_28114,N_28136);
nor U29019 (N_29019,N_28616,N_28832);
nor U29020 (N_29020,N_28263,N_28298);
nand U29021 (N_29021,N_28974,N_28629);
nand U29022 (N_29022,N_28559,N_28671);
nor U29023 (N_29023,N_28943,N_28344);
nor U29024 (N_29024,N_28351,N_28003);
nand U29025 (N_29025,N_28654,N_28279);
or U29026 (N_29026,N_28889,N_28293);
xor U29027 (N_29027,N_28826,N_28822);
nand U29028 (N_29028,N_28986,N_28504);
nor U29029 (N_29029,N_28625,N_28439);
or U29030 (N_29030,N_28729,N_28541);
xnor U29031 (N_29031,N_28390,N_28818);
nor U29032 (N_29032,N_28998,N_28330);
xnor U29033 (N_29033,N_28442,N_28295);
and U29034 (N_29034,N_28901,N_28923);
or U29035 (N_29035,N_28609,N_28947);
nand U29036 (N_29036,N_28709,N_28621);
and U29037 (N_29037,N_28783,N_28042);
and U29038 (N_29038,N_28406,N_28760);
and U29039 (N_29039,N_28059,N_28039);
nor U29040 (N_29040,N_28046,N_28335);
xnor U29041 (N_29041,N_28886,N_28768);
xor U29042 (N_29042,N_28190,N_28318);
nand U29043 (N_29043,N_28372,N_28867);
or U29044 (N_29044,N_28757,N_28339);
or U29045 (N_29045,N_28092,N_28524);
nor U29046 (N_29046,N_28536,N_28622);
and U29047 (N_29047,N_28181,N_28510);
or U29048 (N_29048,N_28422,N_28154);
xor U29049 (N_29049,N_28036,N_28037);
xor U29050 (N_29050,N_28844,N_28991);
or U29051 (N_29051,N_28034,N_28883);
and U29052 (N_29052,N_28932,N_28786);
nor U29053 (N_29053,N_28137,N_28474);
or U29054 (N_29054,N_28382,N_28070);
and U29055 (N_29055,N_28206,N_28311);
nand U29056 (N_29056,N_28728,N_28948);
xnor U29057 (N_29057,N_28276,N_28065);
xor U29058 (N_29058,N_28496,N_28023);
nor U29059 (N_29059,N_28926,N_28585);
and U29060 (N_29060,N_28499,N_28458);
or U29061 (N_29061,N_28550,N_28209);
or U29062 (N_29062,N_28610,N_28535);
nor U29063 (N_29063,N_28951,N_28858);
and U29064 (N_29064,N_28139,N_28838);
xnor U29065 (N_29065,N_28870,N_28424);
and U29066 (N_29066,N_28678,N_28075);
nor U29067 (N_29067,N_28085,N_28526);
xnor U29068 (N_29068,N_28656,N_28096);
nand U29069 (N_29069,N_28753,N_28196);
xnor U29070 (N_29070,N_28102,N_28375);
nand U29071 (N_29071,N_28916,N_28189);
nor U29072 (N_29072,N_28871,N_28975);
xnor U29073 (N_29073,N_28589,N_28359);
and U29074 (N_29074,N_28650,N_28796);
or U29075 (N_29075,N_28099,N_28745);
nor U29076 (N_29076,N_28565,N_28670);
nor U29077 (N_29077,N_28962,N_28447);
nand U29078 (N_29078,N_28333,N_28133);
xor U29079 (N_29079,N_28661,N_28291);
nand U29080 (N_29080,N_28855,N_28058);
nor U29081 (N_29081,N_28104,N_28437);
nand U29082 (N_29082,N_28055,N_28149);
nand U29083 (N_29083,N_28806,N_28516);
nor U29084 (N_29084,N_28505,N_28681);
nor U29085 (N_29085,N_28934,N_28441);
nor U29086 (N_29086,N_28007,N_28476);
nor U29087 (N_29087,N_28045,N_28749);
nor U29088 (N_29088,N_28854,N_28322);
or U29089 (N_29089,N_28266,N_28035);
nor U29090 (N_29090,N_28186,N_28241);
or U29091 (N_29091,N_28172,N_28155);
xnor U29092 (N_29092,N_28759,N_28506);
nand U29093 (N_29093,N_28723,N_28989);
nand U29094 (N_29094,N_28044,N_28269);
nor U29095 (N_29095,N_28066,N_28959);
nor U29096 (N_29096,N_28350,N_28529);
or U29097 (N_29097,N_28325,N_28686);
xnor U29098 (N_29098,N_28987,N_28081);
or U29099 (N_29099,N_28721,N_28471);
nor U29100 (N_29100,N_28762,N_28261);
or U29101 (N_29101,N_28392,N_28970);
or U29102 (N_29102,N_28573,N_28275);
xnor U29103 (N_29103,N_28810,N_28117);
or U29104 (N_29104,N_28539,N_28346);
or U29105 (N_29105,N_28988,N_28869);
and U29106 (N_29106,N_28198,N_28579);
xor U29107 (N_29107,N_28316,N_28775);
nor U29108 (N_29108,N_28255,N_28483);
and U29109 (N_29109,N_28135,N_28495);
nor U29110 (N_29110,N_28792,N_28342);
nand U29111 (N_29111,N_28166,N_28720);
and U29112 (N_29112,N_28863,N_28326);
xnor U29113 (N_29113,N_28690,N_28202);
nand U29114 (N_29114,N_28481,N_28780);
or U29115 (N_29115,N_28493,N_28737);
and U29116 (N_29116,N_28141,N_28057);
nor U29117 (N_29117,N_28002,N_28501);
nor U29118 (N_29118,N_28450,N_28001);
nand U29119 (N_29119,N_28646,N_28286);
or U29120 (N_29120,N_28093,N_28368);
nand U29121 (N_29121,N_28265,N_28126);
nand U29122 (N_29122,N_28887,N_28929);
xor U29123 (N_29123,N_28105,N_28774);
nand U29124 (N_29124,N_28803,N_28937);
or U29125 (N_29125,N_28436,N_28252);
nand U29126 (N_29126,N_28688,N_28902);
xor U29127 (N_29127,N_28453,N_28772);
or U29128 (N_29128,N_28233,N_28310);
nor U29129 (N_29129,N_28598,N_28809);
nor U29130 (N_29130,N_28733,N_28460);
nand U29131 (N_29131,N_28121,N_28672);
and U29132 (N_29132,N_28373,N_28395);
and U29133 (N_29133,N_28313,N_28866);
and U29134 (N_29134,N_28531,N_28801);
or U29135 (N_29135,N_28755,N_28486);
and U29136 (N_29136,N_28289,N_28304);
nor U29137 (N_29137,N_28773,N_28861);
xnor U29138 (N_29138,N_28732,N_28743);
xor U29139 (N_29139,N_28319,N_28845);
xor U29140 (N_29140,N_28634,N_28240);
nor U29141 (N_29141,N_28689,N_28581);
xor U29142 (N_29142,N_28715,N_28973);
xor U29143 (N_29143,N_28389,N_28257);
xnor U29144 (N_29144,N_28226,N_28317);
or U29145 (N_29145,N_28894,N_28846);
or U29146 (N_29146,N_28795,N_28778);
or U29147 (N_29147,N_28659,N_28340);
nor U29148 (N_29148,N_28477,N_28630);
or U29149 (N_29149,N_28494,N_28599);
nand U29150 (N_29150,N_28216,N_28387);
or U29151 (N_29151,N_28299,N_28015);
xnor U29152 (N_29152,N_28183,N_28177);
nor U29153 (N_29153,N_28830,N_28677);
and U29154 (N_29154,N_28520,N_28909);
nor U29155 (N_29155,N_28692,N_28582);
xor U29156 (N_29156,N_28853,N_28983);
nor U29157 (N_29157,N_28079,N_28563);
or U29158 (N_29158,N_28461,N_28256);
nor U29159 (N_29159,N_28586,N_28764);
nor U29160 (N_29160,N_28738,N_28560);
nor U29161 (N_29161,N_28297,N_28356);
nor U29162 (N_29162,N_28555,N_28676);
nand U29163 (N_29163,N_28419,N_28511);
xor U29164 (N_29164,N_28074,N_28719);
nor U29165 (N_29165,N_28605,N_28651);
xor U29166 (N_29166,N_28432,N_28400);
nand U29167 (N_29167,N_28124,N_28712);
or U29168 (N_29168,N_28321,N_28590);
or U29169 (N_29169,N_28146,N_28821);
nor U29170 (N_29170,N_28403,N_28982);
or U29171 (N_29171,N_28110,N_28355);
nor U29172 (N_29172,N_28469,N_28132);
xnor U29173 (N_29173,N_28928,N_28788);
nand U29174 (N_29174,N_28296,N_28487);
and U29175 (N_29175,N_28770,N_28143);
xnor U29176 (N_29176,N_28100,N_28706);
or U29177 (N_29177,N_28969,N_28736);
and U29178 (N_29178,N_28281,N_28848);
or U29179 (N_29179,N_28060,N_28575);
xor U29180 (N_29180,N_28184,N_28163);
xnor U29181 (N_29181,N_28153,N_28636);
nor U29182 (N_29182,N_28769,N_28613);
and U29183 (N_29183,N_28258,N_28120);
xnor U29184 (N_29184,N_28679,N_28466);
xor U29185 (N_29185,N_28073,N_28594);
nor U29186 (N_29186,N_28927,N_28602);
nand U29187 (N_29187,N_28080,N_28160);
xor U29188 (N_29188,N_28203,N_28776);
or U29189 (N_29189,N_28016,N_28725);
or U29190 (N_29190,N_28608,N_28842);
nor U29191 (N_29191,N_28884,N_28680);
nor U29192 (N_29192,N_28649,N_28250);
xor U29193 (N_29193,N_28445,N_28940);
or U29194 (N_29194,N_28239,N_28816);
and U29195 (N_29195,N_28569,N_28668);
or U29196 (N_29196,N_28349,N_28833);
nand U29197 (N_29197,N_28164,N_28664);
nor U29198 (N_29198,N_28882,N_28361);
or U29199 (N_29199,N_28981,N_28307);
or U29200 (N_29200,N_28031,N_28591);
xor U29201 (N_29201,N_28013,N_28717);
and U29202 (N_29202,N_28048,N_28470);
or U29203 (N_29203,N_28829,N_28026);
or U29204 (N_29204,N_28302,N_28949);
xor U29205 (N_29205,N_28823,N_28374);
nor U29206 (N_29206,N_28534,N_28794);
xor U29207 (N_29207,N_28614,N_28305);
nand U29208 (N_29208,N_28147,N_28038);
nand U29209 (N_29209,N_28956,N_28207);
or U29210 (N_29210,N_28404,N_28260);
or U29211 (N_29211,N_28264,N_28918);
nand U29212 (N_29212,N_28027,N_28201);
or U29213 (N_29213,N_28101,N_28623);
or U29214 (N_29214,N_28587,N_28808);
and U29215 (N_29215,N_28817,N_28831);
or U29216 (N_29216,N_28378,N_28008);
nand U29217 (N_29217,N_28702,N_28532);
or U29218 (N_29218,N_28953,N_28489);
and U29219 (N_29219,N_28980,N_28642);
and U29220 (N_29220,N_28353,N_28379);
nand U29221 (N_29221,N_28345,N_28028);
xnor U29222 (N_29222,N_28811,N_28872);
or U29223 (N_29223,N_28414,N_28718);
and U29224 (N_29224,N_28767,N_28309);
xor U29225 (N_29225,N_28456,N_28662);
xor U29226 (N_29226,N_28278,N_28512);
nor U29227 (N_29227,N_28628,N_28421);
nor U29228 (N_29228,N_28367,N_28014);
xnor U29229 (N_29229,N_28643,N_28549);
and U29230 (N_29230,N_28711,N_28840);
and U29231 (N_29231,N_28547,N_28005);
xor U29232 (N_29232,N_28924,N_28019);
xnor U29233 (N_29233,N_28750,N_28362);
nand U29234 (N_29234,N_28371,N_28968);
xor U29235 (N_29235,N_28592,N_28967);
nor U29236 (N_29236,N_28548,N_28793);
xor U29237 (N_29237,N_28851,N_28523);
and U29238 (N_29238,N_28624,N_28354);
and U29239 (N_29239,N_28399,N_28259);
or U29240 (N_29240,N_28468,N_28997);
or U29241 (N_29241,N_28554,N_28984);
or U29242 (N_29242,N_28220,N_28455);
nand U29243 (N_29243,N_28544,N_28268);
or U29244 (N_29244,N_28875,N_28785);
nand U29245 (N_29245,N_28566,N_28498);
or U29246 (N_29246,N_28935,N_28612);
nand U29247 (N_29247,N_28423,N_28029);
and U29248 (N_29248,N_28211,N_28485);
or U29249 (N_29249,N_28248,N_28868);
nor U29250 (N_29250,N_28742,N_28430);
xnor U29251 (N_29251,N_28782,N_28542);
xor U29252 (N_29252,N_28519,N_28696);
xnor U29253 (N_29253,N_28683,N_28665);
and U29254 (N_29254,N_28915,N_28283);
xnor U29255 (N_29255,N_28618,N_28675);
or U29256 (N_29256,N_28140,N_28763);
nand U29257 (N_29257,N_28417,N_28352);
nand U29258 (N_29258,N_28347,N_28401);
xor U29259 (N_29259,N_28507,N_28807);
or U29260 (N_29260,N_28218,N_28011);
nor U29261 (N_29261,N_28601,N_28653);
nor U29262 (N_29262,N_28513,N_28580);
xnor U29263 (N_29263,N_28734,N_28950);
and U29264 (N_29264,N_28115,N_28619);
or U29265 (N_29265,N_28508,N_28064);
xnor U29266 (N_29266,N_28145,N_28267);
or U29267 (N_29267,N_28254,N_28864);
or U29268 (N_29268,N_28285,N_28062);
or U29269 (N_29269,N_28393,N_28633);
or U29270 (N_29270,N_28205,N_28328);
and U29271 (N_29271,N_28332,N_28448);
and U29272 (N_29272,N_28658,N_28213);
nand U29273 (N_29273,N_28879,N_28941);
nand U29274 (N_29274,N_28540,N_28859);
or U29275 (N_29275,N_28288,N_28052);
xor U29276 (N_29276,N_28179,N_28597);
or U29277 (N_29277,N_28251,N_28976);
nand U29278 (N_29278,N_28323,N_28896);
nand U29279 (N_29279,N_28123,N_28237);
and U29280 (N_29280,N_28385,N_28522);
or U29281 (N_29281,N_28054,N_28161);
nand U29282 (N_29282,N_28880,N_28480);
and U29283 (N_29283,N_28682,N_28113);
xnor U29284 (N_29284,N_28193,N_28428);
xor U29285 (N_29285,N_28227,N_28553);
nor U29286 (N_29286,N_28647,N_28551);
and U29287 (N_29287,N_28805,N_28944);
nor U29288 (N_29288,N_28097,N_28804);
or U29289 (N_29289,N_28771,N_28936);
and U29290 (N_29290,N_28000,N_28134);
and U29291 (N_29291,N_28273,N_28971);
xnor U29292 (N_29292,N_28475,N_28050);
nor U29293 (N_29293,N_28068,N_28129);
and U29294 (N_29294,N_28109,N_28314);
nand U29295 (N_29295,N_28178,N_28040);
xor U29296 (N_29296,N_28942,N_28169);
and U29297 (N_29297,N_28041,N_28790);
or U29298 (N_29298,N_28952,N_28663);
and U29299 (N_29299,N_28063,N_28088);
xnor U29300 (N_29300,N_28525,N_28912);
and U29301 (N_29301,N_28922,N_28391);
nand U29302 (N_29302,N_28568,N_28452);
or U29303 (N_29303,N_28862,N_28825);
nand U29304 (N_29304,N_28090,N_28082);
nand U29305 (N_29305,N_28890,N_28584);
xor U29306 (N_29306,N_28638,N_28488);
or U29307 (N_29307,N_28364,N_28021);
or U29308 (N_29308,N_28231,N_28637);
xnor U29309 (N_29309,N_28684,N_28300);
or U29310 (N_29310,N_28600,N_28130);
or U29311 (N_29311,N_28731,N_28383);
or U29312 (N_29312,N_28722,N_28187);
nand U29313 (N_29313,N_28687,N_28413);
nand U29314 (N_29314,N_28892,N_28815);
xnor U29315 (N_29315,N_28545,N_28235);
xor U29316 (N_29316,N_28223,N_28841);
nand U29317 (N_29317,N_28168,N_28434);
nand U29318 (N_29318,N_28552,N_28282);
nand U29319 (N_29319,N_28271,N_28217);
nor U29320 (N_29320,N_28604,N_28502);
nor U29321 (N_29321,N_28707,N_28192);
nor U29322 (N_29322,N_28290,N_28337);
and U29323 (N_29323,N_28365,N_28946);
or U29324 (N_29324,N_28188,N_28979);
nand U29325 (N_29325,N_28197,N_28860);
and U29326 (N_29326,N_28171,N_28107);
nand U29327 (N_29327,N_28693,N_28873);
and U29328 (N_29328,N_28641,N_28324);
and U29329 (N_29329,N_28999,N_28410);
nand U29330 (N_29330,N_28022,N_28479);
and U29331 (N_29331,N_28899,N_28444);
nor U29332 (N_29332,N_28484,N_28242);
nand U29333 (N_29333,N_28577,N_28409);
nor U29334 (N_29334,N_28343,N_28144);
or U29335 (N_29335,N_28537,N_28384);
and U29336 (N_29336,N_28595,N_28897);
nor U29337 (N_29337,N_28463,N_28639);
xnor U29338 (N_29338,N_28657,N_28162);
nor U29339 (N_29339,N_28972,N_28877);
nor U29340 (N_29340,N_28176,N_28813);
nand U29341 (N_29341,N_28708,N_28405);
or U29342 (N_29342,N_28703,N_28357);
or U29343 (N_29343,N_28945,N_28334);
nor U29344 (N_29344,N_28215,N_28546);
nand U29345 (N_29345,N_28095,N_28234);
nor U29346 (N_29346,N_28348,N_28797);
nand U29347 (N_29347,N_28704,N_28528);
xor U29348 (N_29348,N_28397,N_28607);
or U29349 (N_29349,N_28128,N_28067);
and U29350 (N_29350,N_28412,N_28515);
nor U29351 (N_29351,N_28086,N_28834);
or U29352 (N_29352,N_28992,N_28930);
nand U29353 (N_29353,N_28284,N_28977);
xor U29354 (N_29354,N_28533,N_28931);
and U29355 (N_29355,N_28802,N_28900);
nand U29356 (N_29356,N_28847,N_28411);
or U29357 (N_29357,N_28611,N_28212);
or U29358 (N_29358,N_28701,N_28740);
xor U29359 (N_29359,N_28174,N_28363);
nor U29360 (N_29360,N_28878,N_28669);
nand U29361 (N_29361,N_28030,N_28210);
nor U29362 (N_29362,N_28645,N_28925);
nand U29363 (N_29363,N_28230,N_28713);
nor U29364 (N_29364,N_28849,N_28514);
or U29365 (N_29365,N_28119,N_28440);
xnor U29366 (N_29366,N_28049,N_28416);
nor U29367 (N_29367,N_28503,N_28150);
or U29368 (N_29368,N_28754,N_28561);
or U29369 (N_29369,N_28908,N_28530);
or U29370 (N_29370,N_28170,N_28881);
nand U29371 (N_29371,N_28004,N_28814);
and U29372 (N_29372,N_28726,N_28472);
and U29373 (N_29373,N_28103,N_28500);
nand U29374 (N_29374,N_28955,N_28572);
nor U29375 (N_29375,N_28996,N_28888);
and U29376 (N_29376,N_28963,N_28018);
or U29377 (N_29377,N_28061,N_28857);
nor U29378 (N_29378,N_28157,N_28244);
xnor U29379 (N_29379,N_28938,N_28843);
or U29380 (N_29380,N_28521,N_28377);
xnor U29381 (N_29381,N_28995,N_28051);
or U29382 (N_29382,N_28329,N_28564);
and U29383 (N_29383,N_28185,N_28603);
nand U29384 (N_29384,N_28799,N_28960);
xnor U29385 (N_29385,N_28228,N_28751);
or U29386 (N_29386,N_28911,N_28308);
nor U29387 (N_29387,N_28238,N_28538);
nor U29388 (N_29388,N_28084,N_28415);
nor U29389 (N_29389,N_28756,N_28583);
or U29390 (N_29390,N_28913,N_28232);
and U29391 (N_29391,N_28697,N_28852);
or U29392 (N_29392,N_28509,N_28012);
or U29393 (N_29393,N_28017,N_28358);
nor U29394 (N_29394,N_28735,N_28236);
and U29395 (N_29395,N_28571,N_28490);
nand U29396 (N_29396,N_28666,N_28606);
xor U29397 (N_29397,N_28667,N_28777);
nor U29398 (N_29398,N_28567,N_28069);
nor U29399 (N_29399,N_28388,N_28072);
nand U29400 (N_29400,N_28116,N_28800);
xor U29401 (N_29401,N_28784,N_28253);
xor U29402 (N_29402,N_28965,N_28089);
xnor U29403 (N_29403,N_28173,N_28214);
nand U29404 (N_29404,N_28798,N_28699);
nor U29405 (N_29405,N_28910,N_28462);
nor U29406 (N_29406,N_28626,N_28446);
nor U29407 (N_29407,N_28994,N_28705);
xor U29408 (N_29408,N_28766,N_28246);
and U29409 (N_29409,N_28557,N_28917);
nand U29410 (N_29410,N_28903,N_28836);
nand U29411 (N_29411,N_28978,N_28839);
nor U29412 (N_29412,N_28820,N_28370);
nand U29413 (N_29413,N_28741,N_28631);
nor U29414 (N_29414,N_28301,N_28744);
and U29415 (N_29415,N_28182,N_28791);
xnor U29416 (N_29416,N_28369,N_28224);
xor U29417 (N_29417,N_28433,N_28674);
and U29418 (N_29418,N_28527,N_28118);
and U29419 (N_29419,N_28009,N_28876);
nor U29420 (N_29420,N_28127,N_28076);
or U29421 (N_29421,N_28386,N_28338);
nor U29422 (N_29422,N_28287,N_28245);
nor U29423 (N_29423,N_28274,N_28427);
xor U29424 (N_29424,N_28006,N_28985);
nand U29425 (N_29425,N_28247,N_28914);
nand U29426 (N_29426,N_28966,N_28835);
or U29427 (N_29427,N_28710,N_28122);
or U29428 (N_29428,N_28765,N_28431);
nand U29429 (N_29429,N_28083,N_28222);
or U29430 (N_29430,N_28964,N_28620);
or U29431 (N_29431,N_28907,N_28071);
xor U29432 (N_29432,N_28714,N_28435);
or U29433 (N_29433,N_28396,N_28142);
nor U29434 (N_29434,N_28315,N_28954);
and U29435 (N_29435,N_28655,N_28652);
nand U29436 (N_29436,N_28243,N_28125);
xor U29437 (N_29437,N_28556,N_28408);
nand U29438 (N_29438,N_28648,N_28558);
and U29439 (N_29439,N_28131,N_28336);
nand U29440 (N_29440,N_28716,N_28615);
nand U29441 (N_29441,N_28921,N_28518);
nor U29442 (N_29442,N_28492,N_28588);
and U29443 (N_29443,N_28112,N_28761);
nor U29444 (N_29444,N_28429,N_28312);
xor U29445 (N_29445,N_28543,N_28294);
xor U29446 (N_29446,N_28151,N_28219);
xor U29447 (N_29447,N_28108,N_28644);
and U29448 (N_29448,N_28491,N_28056);
xnor U29449 (N_29449,N_28691,N_28837);
or U29450 (N_29450,N_28380,N_28175);
xor U29451 (N_29451,N_28199,N_28482);
and U29452 (N_29452,N_28895,N_28919);
and U29453 (N_29453,N_28904,N_28752);
nand U29454 (N_29454,N_28789,N_28562);
or U29455 (N_29455,N_28156,N_28746);
nor U29456 (N_29456,N_28856,N_28640);
nor U29457 (N_29457,N_28087,N_28576);
nand U29458 (N_29458,N_28033,N_28497);
nand U29459 (N_29459,N_28574,N_28194);
and U29460 (N_29460,N_28449,N_28047);
nor U29461 (N_29461,N_28727,N_28221);
xor U29462 (N_29462,N_28700,N_28724);
xnor U29463 (N_29463,N_28578,N_28292);
and U29464 (N_29464,N_28593,N_28376);
xnor U29465 (N_29465,N_28152,N_28420);
nand U29466 (N_29466,N_28032,N_28366);
nor U29467 (N_29467,N_28191,N_28465);
and U29468 (N_29468,N_28957,N_28280);
and U29469 (N_29469,N_28180,N_28891);
nor U29470 (N_29470,N_28478,N_28464);
nand U29471 (N_29471,N_28596,N_28320);
nand U29472 (N_29472,N_28249,N_28148);
and U29473 (N_29473,N_28905,N_28270);
and U29474 (N_29474,N_28381,N_28885);
or U29475 (N_29475,N_28739,N_28200);
or U29476 (N_29476,N_28454,N_28303);
or U29477 (N_29477,N_28418,N_28106);
nor U29478 (N_29478,N_28167,N_28865);
and U29479 (N_29479,N_28341,N_28043);
nand U29480 (N_29480,N_28098,N_28939);
and U29481 (N_29481,N_28893,N_28138);
nand U29482 (N_29482,N_28698,N_28660);
xor U29483 (N_29483,N_28010,N_28443);
or U29484 (N_29484,N_28407,N_28208);
nand U29485 (N_29485,N_28748,N_28920);
or U29486 (N_29486,N_28158,N_28627);
nor U29487 (N_29487,N_28078,N_28438);
xnor U29488 (N_29488,N_28990,N_28570);
nand U29489 (N_29489,N_28020,N_28425);
or U29490 (N_29490,N_28111,N_28091);
xor U29491 (N_29491,N_28747,N_28204);
xor U29492 (N_29492,N_28958,N_28277);
xnor U29493 (N_29493,N_28467,N_28730);
nor U29494 (N_29494,N_28850,N_28617);
and U29495 (N_29495,N_28685,N_28473);
xor U29496 (N_29496,N_28828,N_28758);
and U29497 (N_29497,N_28993,N_28327);
or U29498 (N_29498,N_28272,N_28635);
xnor U29499 (N_29499,N_28787,N_28695);
or U29500 (N_29500,N_28730,N_28139);
and U29501 (N_29501,N_28658,N_28110);
nor U29502 (N_29502,N_28814,N_28404);
xnor U29503 (N_29503,N_28236,N_28614);
nand U29504 (N_29504,N_28156,N_28413);
nand U29505 (N_29505,N_28336,N_28694);
xnor U29506 (N_29506,N_28602,N_28162);
xor U29507 (N_29507,N_28276,N_28893);
xnor U29508 (N_29508,N_28792,N_28636);
xnor U29509 (N_29509,N_28184,N_28656);
or U29510 (N_29510,N_28286,N_28662);
nor U29511 (N_29511,N_28435,N_28396);
nand U29512 (N_29512,N_28386,N_28956);
or U29513 (N_29513,N_28254,N_28827);
and U29514 (N_29514,N_28076,N_28811);
nand U29515 (N_29515,N_28285,N_28277);
xor U29516 (N_29516,N_28455,N_28929);
nand U29517 (N_29517,N_28916,N_28295);
or U29518 (N_29518,N_28621,N_28448);
and U29519 (N_29519,N_28517,N_28897);
nand U29520 (N_29520,N_28418,N_28513);
or U29521 (N_29521,N_28164,N_28047);
and U29522 (N_29522,N_28154,N_28354);
nor U29523 (N_29523,N_28093,N_28798);
and U29524 (N_29524,N_28909,N_28290);
xor U29525 (N_29525,N_28170,N_28435);
xnor U29526 (N_29526,N_28907,N_28617);
nor U29527 (N_29527,N_28461,N_28852);
or U29528 (N_29528,N_28513,N_28862);
nand U29529 (N_29529,N_28879,N_28228);
xnor U29530 (N_29530,N_28147,N_28800);
nor U29531 (N_29531,N_28422,N_28746);
and U29532 (N_29532,N_28220,N_28399);
nor U29533 (N_29533,N_28213,N_28921);
or U29534 (N_29534,N_28048,N_28030);
and U29535 (N_29535,N_28950,N_28503);
nand U29536 (N_29536,N_28282,N_28674);
nor U29537 (N_29537,N_28403,N_28988);
or U29538 (N_29538,N_28126,N_28845);
or U29539 (N_29539,N_28717,N_28636);
xor U29540 (N_29540,N_28637,N_28729);
or U29541 (N_29541,N_28699,N_28919);
nand U29542 (N_29542,N_28309,N_28256);
and U29543 (N_29543,N_28793,N_28544);
xor U29544 (N_29544,N_28743,N_28521);
or U29545 (N_29545,N_28758,N_28915);
or U29546 (N_29546,N_28165,N_28368);
or U29547 (N_29547,N_28433,N_28217);
or U29548 (N_29548,N_28218,N_28697);
xor U29549 (N_29549,N_28761,N_28596);
and U29550 (N_29550,N_28063,N_28710);
nand U29551 (N_29551,N_28783,N_28023);
or U29552 (N_29552,N_28277,N_28898);
and U29553 (N_29553,N_28477,N_28097);
nor U29554 (N_29554,N_28899,N_28969);
and U29555 (N_29555,N_28527,N_28442);
nor U29556 (N_29556,N_28335,N_28953);
and U29557 (N_29557,N_28064,N_28007);
or U29558 (N_29558,N_28872,N_28891);
nand U29559 (N_29559,N_28457,N_28732);
or U29560 (N_29560,N_28658,N_28252);
and U29561 (N_29561,N_28354,N_28762);
nor U29562 (N_29562,N_28151,N_28420);
nand U29563 (N_29563,N_28928,N_28676);
nor U29564 (N_29564,N_28196,N_28672);
and U29565 (N_29565,N_28924,N_28057);
or U29566 (N_29566,N_28610,N_28924);
and U29567 (N_29567,N_28006,N_28884);
or U29568 (N_29568,N_28456,N_28941);
and U29569 (N_29569,N_28930,N_28489);
xor U29570 (N_29570,N_28264,N_28738);
or U29571 (N_29571,N_28442,N_28543);
nor U29572 (N_29572,N_28543,N_28819);
nor U29573 (N_29573,N_28869,N_28859);
nand U29574 (N_29574,N_28802,N_28363);
nand U29575 (N_29575,N_28349,N_28747);
nand U29576 (N_29576,N_28572,N_28115);
and U29577 (N_29577,N_28573,N_28185);
or U29578 (N_29578,N_28455,N_28668);
nor U29579 (N_29579,N_28955,N_28742);
xor U29580 (N_29580,N_28360,N_28582);
xor U29581 (N_29581,N_28937,N_28778);
nor U29582 (N_29582,N_28482,N_28213);
xnor U29583 (N_29583,N_28783,N_28316);
xor U29584 (N_29584,N_28357,N_28885);
and U29585 (N_29585,N_28551,N_28405);
xnor U29586 (N_29586,N_28894,N_28612);
nor U29587 (N_29587,N_28230,N_28637);
nor U29588 (N_29588,N_28309,N_28738);
nor U29589 (N_29589,N_28487,N_28101);
nor U29590 (N_29590,N_28727,N_28536);
nand U29591 (N_29591,N_28574,N_28565);
nand U29592 (N_29592,N_28521,N_28168);
xnor U29593 (N_29593,N_28152,N_28948);
or U29594 (N_29594,N_28962,N_28274);
or U29595 (N_29595,N_28146,N_28251);
nand U29596 (N_29596,N_28100,N_28451);
xor U29597 (N_29597,N_28081,N_28960);
nand U29598 (N_29598,N_28770,N_28786);
or U29599 (N_29599,N_28457,N_28593);
xnor U29600 (N_29600,N_28134,N_28699);
or U29601 (N_29601,N_28969,N_28020);
nand U29602 (N_29602,N_28199,N_28441);
nand U29603 (N_29603,N_28132,N_28473);
nor U29604 (N_29604,N_28213,N_28784);
or U29605 (N_29605,N_28251,N_28380);
and U29606 (N_29606,N_28212,N_28344);
nor U29607 (N_29607,N_28862,N_28138);
xnor U29608 (N_29608,N_28874,N_28309);
and U29609 (N_29609,N_28930,N_28104);
nand U29610 (N_29610,N_28602,N_28976);
or U29611 (N_29611,N_28473,N_28048);
nor U29612 (N_29612,N_28514,N_28268);
xnor U29613 (N_29613,N_28337,N_28646);
xor U29614 (N_29614,N_28825,N_28284);
xor U29615 (N_29615,N_28610,N_28494);
nand U29616 (N_29616,N_28351,N_28789);
xor U29617 (N_29617,N_28170,N_28809);
nor U29618 (N_29618,N_28333,N_28885);
or U29619 (N_29619,N_28252,N_28894);
xor U29620 (N_29620,N_28586,N_28601);
or U29621 (N_29621,N_28297,N_28246);
xnor U29622 (N_29622,N_28993,N_28347);
and U29623 (N_29623,N_28217,N_28314);
xnor U29624 (N_29624,N_28288,N_28696);
or U29625 (N_29625,N_28013,N_28220);
xor U29626 (N_29626,N_28833,N_28121);
nor U29627 (N_29627,N_28769,N_28932);
or U29628 (N_29628,N_28767,N_28105);
and U29629 (N_29629,N_28503,N_28755);
nand U29630 (N_29630,N_28916,N_28483);
or U29631 (N_29631,N_28023,N_28310);
nand U29632 (N_29632,N_28722,N_28493);
and U29633 (N_29633,N_28193,N_28088);
or U29634 (N_29634,N_28398,N_28130);
or U29635 (N_29635,N_28451,N_28933);
and U29636 (N_29636,N_28490,N_28185);
xor U29637 (N_29637,N_28299,N_28838);
and U29638 (N_29638,N_28879,N_28461);
nand U29639 (N_29639,N_28403,N_28022);
and U29640 (N_29640,N_28074,N_28683);
or U29641 (N_29641,N_28969,N_28902);
xor U29642 (N_29642,N_28098,N_28297);
xor U29643 (N_29643,N_28687,N_28782);
nor U29644 (N_29644,N_28227,N_28752);
or U29645 (N_29645,N_28146,N_28526);
or U29646 (N_29646,N_28647,N_28583);
nand U29647 (N_29647,N_28176,N_28674);
nor U29648 (N_29648,N_28819,N_28571);
nor U29649 (N_29649,N_28781,N_28648);
and U29650 (N_29650,N_28365,N_28444);
nor U29651 (N_29651,N_28801,N_28633);
xnor U29652 (N_29652,N_28664,N_28561);
nand U29653 (N_29653,N_28269,N_28836);
xor U29654 (N_29654,N_28014,N_28178);
nor U29655 (N_29655,N_28773,N_28750);
nor U29656 (N_29656,N_28814,N_28499);
and U29657 (N_29657,N_28097,N_28829);
or U29658 (N_29658,N_28476,N_28209);
xor U29659 (N_29659,N_28436,N_28537);
xnor U29660 (N_29660,N_28062,N_28254);
and U29661 (N_29661,N_28044,N_28900);
xor U29662 (N_29662,N_28655,N_28575);
or U29663 (N_29663,N_28420,N_28999);
xnor U29664 (N_29664,N_28124,N_28080);
nor U29665 (N_29665,N_28718,N_28847);
or U29666 (N_29666,N_28100,N_28397);
and U29667 (N_29667,N_28884,N_28212);
nand U29668 (N_29668,N_28717,N_28172);
or U29669 (N_29669,N_28594,N_28384);
xor U29670 (N_29670,N_28599,N_28055);
and U29671 (N_29671,N_28886,N_28715);
xor U29672 (N_29672,N_28703,N_28389);
xor U29673 (N_29673,N_28953,N_28843);
and U29674 (N_29674,N_28275,N_28048);
and U29675 (N_29675,N_28854,N_28578);
nor U29676 (N_29676,N_28539,N_28339);
xnor U29677 (N_29677,N_28821,N_28303);
and U29678 (N_29678,N_28760,N_28855);
xnor U29679 (N_29679,N_28092,N_28174);
nand U29680 (N_29680,N_28135,N_28986);
or U29681 (N_29681,N_28062,N_28856);
xnor U29682 (N_29682,N_28919,N_28276);
or U29683 (N_29683,N_28234,N_28097);
and U29684 (N_29684,N_28309,N_28266);
nor U29685 (N_29685,N_28036,N_28839);
nand U29686 (N_29686,N_28689,N_28364);
xor U29687 (N_29687,N_28964,N_28490);
xnor U29688 (N_29688,N_28236,N_28752);
or U29689 (N_29689,N_28576,N_28779);
and U29690 (N_29690,N_28974,N_28038);
nand U29691 (N_29691,N_28526,N_28893);
nand U29692 (N_29692,N_28972,N_28835);
nand U29693 (N_29693,N_28104,N_28248);
nor U29694 (N_29694,N_28436,N_28684);
nand U29695 (N_29695,N_28336,N_28289);
nand U29696 (N_29696,N_28010,N_28544);
xnor U29697 (N_29697,N_28029,N_28841);
xnor U29698 (N_29698,N_28824,N_28723);
and U29699 (N_29699,N_28589,N_28986);
nand U29700 (N_29700,N_28188,N_28680);
nor U29701 (N_29701,N_28489,N_28878);
nand U29702 (N_29702,N_28976,N_28311);
nor U29703 (N_29703,N_28663,N_28738);
xor U29704 (N_29704,N_28184,N_28393);
nand U29705 (N_29705,N_28201,N_28567);
and U29706 (N_29706,N_28590,N_28685);
and U29707 (N_29707,N_28635,N_28695);
nor U29708 (N_29708,N_28063,N_28873);
and U29709 (N_29709,N_28862,N_28609);
or U29710 (N_29710,N_28981,N_28853);
and U29711 (N_29711,N_28827,N_28219);
xor U29712 (N_29712,N_28210,N_28671);
xor U29713 (N_29713,N_28495,N_28700);
or U29714 (N_29714,N_28457,N_28858);
or U29715 (N_29715,N_28467,N_28301);
nor U29716 (N_29716,N_28898,N_28698);
nand U29717 (N_29717,N_28580,N_28401);
nand U29718 (N_29718,N_28356,N_28661);
and U29719 (N_29719,N_28678,N_28386);
nand U29720 (N_29720,N_28721,N_28168);
or U29721 (N_29721,N_28026,N_28781);
and U29722 (N_29722,N_28577,N_28587);
or U29723 (N_29723,N_28082,N_28128);
and U29724 (N_29724,N_28070,N_28549);
xnor U29725 (N_29725,N_28134,N_28338);
and U29726 (N_29726,N_28397,N_28317);
and U29727 (N_29727,N_28304,N_28430);
nor U29728 (N_29728,N_28550,N_28629);
xor U29729 (N_29729,N_28144,N_28358);
nor U29730 (N_29730,N_28259,N_28555);
or U29731 (N_29731,N_28676,N_28527);
and U29732 (N_29732,N_28772,N_28312);
or U29733 (N_29733,N_28616,N_28595);
or U29734 (N_29734,N_28707,N_28580);
xor U29735 (N_29735,N_28999,N_28770);
or U29736 (N_29736,N_28218,N_28108);
nor U29737 (N_29737,N_28310,N_28500);
or U29738 (N_29738,N_28907,N_28919);
or U29739 (N_29739,N_28802,N_28951);
nand U29740 (N_29740,N_28220,N_28809);
and U29741 (N_29741,N_28766,N_28950);
or U29742 (N_29742,N_28553,N_28116);
xor U29743 (N_29743,N_28376,N_28377);
nor U29744 (N_29744,N_28412,N_28106);
or U29745 (N_29745,N_28417,N_28786);
nand U29746 (N_29746,N_28291,N_28636);
or U29747 (N_29747,N_28179,N_28811);
nor U29748 (N_29748,N_28061,N_28392);
or U29749 (N_29749,N_28616,N_28135);
and U29750 (N_29750,N_28320,N_28094);
or U29751 (N_29751,N_28866,N_28381);
nor U29752 (N_29752,N_28559,N_28644);
and U29753 (N_29753,N_28554,N_28945);
xnor U29754 (N_29754,N_28649,N_28721);
or U29755 (N_29755,N_28461,N_28822);
nor U29756 (N_29756,N_28656,N_28897);
nor U29757 (N_29757,N_28521,N_28753);
nand U29758 (N_29758,N_28110,N_28354);
nor U29759 (N_29759,N_28140,N_28001);
and U29760 (N_29760,N_28965,N_28773);
and U29761 (N_29761,N_28097,N_28215);
xor U29762 (N_29762,N_28167,N_28091);
and U29763 (N_29763,N_28558,N_28151);
or U29764 (N_29764,N_28410,N_28269);
nand U29765 (N_29765,N_28817,N_28177);
xnor U29766 (N_29766,N_28036,N_28335);
nor U29767 (N_29767,N_28873,N_28332);
xor U29768 (N_29768,N_28509,N_28990);
nand U29769 (N_29769,N_28701,N_28781);
and U29770 (N_29770,N_28226,N_28669);
nor U29771 (N_29771,N_28573,N_28873);
nor U29772 (N_29772,N_28037,N_28734);
or U29773 (N_29773,N_28442,N_28165);
or U29774 (N_29774,N_28041,N_28017);
nand U29775 (N_29775,N_28994,N_28721);
and U29776 (N_29776,N_28080,N_28854);
xor U29777 (N_29777,N_28979,N_28563);
and U29778 (N_29778,N_28707,N_28215);
or U29779 (N_29779,N_28536,N_28869);
and U29780 (N_29780,N_28230,N_28561);
nor U29781 (N_29781,N_28085,N_28994);
xor U29782 (N_29782,N_28361,N_28199);
nand U29783 (N_29783,N_28733,N_28688);
or U29784 (N_29784,N_28773,N_28307);
and U29785 (N_29785,N_28149,N_28244);
nor U29786 (N_29786,N_28500,N_28196);
xor U29787 (N_29787,N_28136,N_28579);
or U29788 (N_29788,N_28179,N_28482);
or U29789 (N_29789,N_28873,N_28077);
or U29790 (N_29790,N_28364,N_28943);
nor U29791 (N_29791,N_28736,N_28933);
nand U29792 (N_29792,N_28698,N_28796);
nand U29793 (N_29793,N_28758,N_28659);
or U29794 (N_29794,N_28093,N_28495);
nand U29795 (N_29795,N_28569,N_28331);
and U29796 (N_29796,N_28258,N_28524);
nand U29797 (N_29797,N_28278,N_28499);
or U29798 (N_29798,N_28666,N_28421);
xnor U29799 (N_29799,N_28250,N_28562);
nand U29800 (N_29800,N_28302,N_28497);
xor U29801 (N_29801,N_28850,N_28229);
nor U29802 (N_29802,N_28757,N_28064);
or U29803 (N_29803,N_28589,N_28004);
xor U29804 (N_29804,N_28201,N_28495);
xnor U29805 (N_29805,N_28088,N_28342);
nor U29806 (N_29806,N_28961,N_28270);
nor U29807 (N_29807,N_28039,N_28621);
and U29808 (N_29808,N_28692,N_28849);
nand U29809 (N_29809,N_28024,N_28719);
xnor U29810 (N_29810,N_28971,N_28649);
xor U29811 (N_29811,N_28236,N_28209);
xor U29812 (N_29812,N_28367,N_28868);
xor U29813 (N_29813,N_28718,N_28649);
nor U29814 (N_29814,N_28099,N_28449);
xor U29815 (N_29815,N_28385,N_28924);
or U29816 (N_29816,N_28009,N_28787);
xor U29817 (N_29817,N_28186,N_28708);
xor U29818 (N_29818,N_28347,N_28961);
nor U29819 (N_29819,N_28735,N_28451);
nand U29820 (N_29820,N_28901,N_28889);
xnor U29821 (N_29821,N_28938,N_28663);
and U29822 (N_29822,N_28285,N_28425);
nor U29823 (N_29823,N_28488,N_28753);
nor U29824 (N_29824,N_28181,N_28454);
or U29825 (N_29825,N_28134,N_28051);
nand U29826 (N_29826,N_28905,N_28927);
xor U29827 (N_29827,N_28003,N_28779);
or U29828 (N_29828,N_28070,N_28189);
xor U29829 (N_29829,N_28313,N_28013);
or U29830 (N_29830,N_28204,N_28403);
xnor U29831 (N_29831,N_28553,N_28544);
or U29832 (N_29832,N_28388,N_28469);
or U29833 (N_29833,N_28475,N_28438);
and U29834 (N_29834,N_28024,N_28946);
nor U29835 (N_29835,N_28598,N_28985);
xnor U29836 (N_29836,N_28375,N_28135);
and U29837 (N_29837,N_28375,N_28794);
xor U29838 (N_29838,N_28307,N_28868);
nand U29839 (N_29839,N_28811,N_28531);
xnor U29840 (N_29840,N_28608,N_28857);
nor U29841 (N_29841,N_28218,N_28237);
nor U29842 (N_29842,N_28778,N_28193);
or U29843 (N_29843,N_28549,N_28142);
nand U29844 (N_29844,N_28325,N_28882);
and U29845 (N_29845,N_28437,N_28111);
xor U29846 (N_29846,N_28408,N_28153);
and U29847 (N_29847,N_28177,N_28504);
and U29848 (N_29848,N_28260,N_28125);
or U29849 (N_29849,N_28309,N_28216);
nor U29850 (N_29850,N_28105,N_28315);
nor U29851 (N_29851,N_28283,N_28734);
nand U29852 (N_29852,N_28075,N_28513);
and U29853 (N_29853,N_28627,N_28388);
nor U29854 (N_29854,N_28908,N_28489);
and U29855 (N_29855,N_28937,N_28336);
xor U29856 (N_29856,N_28992,N_28984);
nor U29857 (N_29857,N_28621,N_28336);
nor U29858 (N_29858,N_28182,N_28997);
nor U29859 (N_29859,N_28852,N_28971);
or U29860 (N_29860,N_28778,N_28798);
or U29861 (N_29861,N_28223,N_28207);
or U29862 (N_29862,N_28165,N_28502);
or U29863 (N_29863,N_28263,N_28775);
nand U29864 (N_29864,N_28657,N_28025);
and U29865 (N_29865,N_28461,N_28632);
nand U29866 (N_29866,N_28575,N_28763);
nor U29867 (N_29867,N_28718,N_28416);
and U29868 (N_29868,N_28217,N_28189);
or U29869 (N_29869,N_28743,N_28464);
nor U29870 (N_29870,N_28113,N_28953);
xnor U29871 (N_29871,N_28218,N_28418);
nor U29872 (N_29872,N_28646,N_28413);
xnor U29873 (N_29873,N_28203,N_28820);
nand U29874 (N_29874,N_28906,N_28367);
or U29875 (N_29875,N_28628,N_28670);
nand U29876 (N_29876,N_28561,N_28365);
or U29877 (N_29877,N_28287,N_28481);
or U29878 (N_29878,N_28787,N_28575);
xor U29879 (N_29879,N_28913,N_28764);
nand U29880 (N_29880,N_28004,N_28723);
xor U29881 (N_29881,N_28667,N_28755);
xnor U29882 (N_29882,N_28531,N_28090);
xnor U29883 (N_29883,N_28504,N_28982);
nand U29884 (N_29884,N_28907,N_28160);
xor U29885 (N_29885,N_28787,N_28357);
nor U29886 (N_29886,N_28142,N_28835);
nor U29887 (N_29887,N_28720,N_28577);
nor U29888 (N_29888,N_28202,N_28815);
and U29889 (N_29889,N_28703,N_28784);
xor U29890 (N_29890,N_28878,N_28013);
nor U29891 (N_29891,N_28980,N_28414);
nor U29892 (N_29892,N_28558,N_28992);
nor U29893 (N_29893,N_28305,N_28398);
nor U29894 (N_29894,N_28298,N_28558);
nor U29895 (N_29895,N_28924,N_28946);
or U29896 (N_29896,N_28216,N_28543);
nand U29897 (N_29897,N_28636,N_28337);
xnor U29898 (N_29898,N_28446,N_28380);
or U29899 (N_29899,N_28904,N_28800);
xor U29900 (N_29900,N_28050,N_28443);
xor U29901 (N_29901,N_28924,N_28350);
nand U29902 (N_29902,N_28553,N_28905);
nor U29903 (N_29903,N_28593,N_28213);
xnor U29904 (N_29904,N_28508,N_28911);
or U29905 (N_29905,N_28159,N_28327);
xor U29906 (N_29906,N_28526,N_28517);
nor U29907 (N_29907,N_28521,N_28372);
or U29908 (N_29908,N_28788,N_28756);
and U29909 (N_29909,N_28763,N_28577);
nor U29910 (N_29910,N_28238,N_28982);
and U29911 (N_29911,N_28901,N_28315);
nand U29912 (N_29912,N_28618,N_28824);
and U29913 (N_29913,N_28903,N_28740);
and U29914 (N_29914,N_28833,N_28027);
and U29915 (N_29915,N_28860,N_28159);
or U29916 (N_29916,N_28349,N_28300);
nand U29917 (N_29917,N_28007,N_28396);
nor U29918 (N_29918,N_28227,N_28613);
xor U29919 (N_29919,N_28864,N_28307);
or U29920 (N_29920,N_28618,N_28661);
nand U29921 (N_29921,N_28914,N_28280);
nand U29922 (N_29922,N_28682,N_28883);
nor U29923 (N_29923,N_28634,N_28530);
or U29924 (N_29924,N_28199,N_28325);
or U29925 (N_29925,N_28636,N_28987);
or U29926 (N_29926,N_28504,N_28922);
and U29927 (N_29927,N_28295,N_28495);
xor U29928 (N_29928,N_28465,N_28851);
xor U29929 (N_29929,N_28166,N_28699);
and U29930 (N_29930,N_28419,N_28141);
xor U29931 (N_29931,N_28749,N_28823);
nor U29932 (N_29932,N_28433,N_28093);
or U29933 (N_29933,N_28236,N_28684);
nand U29934 (N_29934,N_28074,N_28226);
xor U29935 (N_29935,N_28083,N_28912);
nor U29936 (N_29936,N_28655,N_28574);
xor U29937 (N_29937,N_28051,N_28942);
xor U29938 (N_29938,N_28451,N_28002);
or U29939 (N_29939,N_28722,N_28989);
nand U29940 (N_29940,N_28411,N_28177);
nand U29941 (N_29941,N_28039,N_28455);
nor U29942 (N_29942,N_28526,N_28408);
xor U29943 (N_29943,N_28255,N_28425);
nand U29944 (N_29944,N_28638,N_28730);
or U29945 (N_29945,N_28456,N_28576);
or U29946 (N_29946,N_28175,N_28065);
or U29947 (N_29947,N_28222,N_28555);
or U29948 (N_29948,N_28404,N_28908);
nor U29949 (N_29949,N_28224,N_28915);
and U29950 (N_29950,N_28852,N_28165);
nor U29951 (N_29951,N_28671,N_28681);
nand U29952 (N_29952,N_28335,N_28242);
nand U29953 (N_29953,N_28868,N_28303);
nor U29954 (N_29954,N_28777,N_28090);
nor U29955 (N_29955,N_28675,N_28542);
and U29956 (N_29956,N_28130,N_28516);
nand U29957 (N_29957,N_28068,N_28497);
or U29958 (N_29958,N_28019,N_28675);
nand U29959 (N_29959,N_28038,N_28753);
nor U29960 (N_29960,N_28324,N_28490);
nand U29961 (N_29961,N_28229,N_28181);
or U29962 (N_29962,N_28795,N_28096);
or U29963 (N_29963,N_28895,N_28606);
nor U29964 (N_29964,N_28122,N_28706);
nand U29965 (N_29965,N_28068,N_28366);
or U29966 (N_29966,N_28157,N_28821);
and U29967 (N_29967,N_28324,N_28871);
and U29968 (N_29968,N_28867,N_28140);
xnor U29969 (N_29969,N_28583,N_28322);
xor U29970 (N_29970,N_28747,N_28309);
nor U29971 (N_29971,N_28854,N_28065);
nand U29972 (N_29972,N_28587,N_28492);
and U29973 (N_29973,N_28114,N_28748);
or U29974 (N_29974,N_28333,N_28422);
nor U29975 (N_29975,N_28080,N_28925);
xnor U29976 (N_29976,N_28849,N_28595);
nor U29977 (N_29977,N_28990,N_28736);
nand U29978 (N_29978,N_28538,N_28469);
and U29979 (N_29979,N_28283,N_28426);
and U29980 (N_29980,N_28289,N_28409);
nor U29981 (N_29981,N_28874,N_28480);
nand U29982 (N_29982,N_28364,N_28120);
or U29983 (N_29983,N_28616,N_28877);
and U29984 (N_29984,N_28305,N_28237);
nand U29985 (N_29985,N_28110,N_28333);
or U29986 (N_29986,N_28164,N_28807);
and U29987 (N_29987,N_28024,N_28690);
xnor U29988 (N_29988,N_28077,N_28935);
or U29989 (N_29989,N_28077,N_28335);
nor U29990 (N_29990,N_28701,N_28132);
nor U29991 (N_29991,N_28387,N_28352);
nor U29992 (N_29992,N_28039,N_28294);
xnor U29993 (N_29993,N_28049,N_28592);
xor U29994 (N_29994,N_28521,N_28660);
nor U29995 (N_29995,N_28260,N_28547);
xor U29996 (N_29996,N_28319,N_28117);
xnor U29997 (N_29997,N_28278,N_28397);
or U29998 (N_29998,N_28184,N_28462);
nor U29999 (N_29999,N_28030,N_28639);
or UO_0 (O_0,N_29844,N_29818);
and UO_1 (O_1,N_29593,N_29392);
nor UO_2 (O_2,N_29707,N_29098);
or UO_3 (O_3,N_29631,N_29495);
nor UO_4 (O_4,N_29718,N_29850);
or UO_5 (O_5,N_29244,N_29548);
xor UO_6 (O_6,N_29658,N_29117);
or UO_7 (O_7,N_29561,N_29231);
xor UO_8 (O_8,N_29408,N_29185);
nor UO_9 (O_9,N_29123,N_29960);
nand UO_10 (O_10,N_29876,N_29405);
nor UO_11 (O_11,N_29459,N_29996);
and UO_12 (O_12,N_29926,N_29653);
nor UO_13 (O_13,N_29949,N_29167);
nor UO_14 (O_14,N_29272,N_29282);
and UO_15 (O_15,N_29087,N_29596);
and UO_16 (O_16,N_29204,N_29440);
nor UO_17 (O_17,N_29727,N_29371);
or UO_18 (O_18,N_29964,N_29385);
or UO_19 (O_19,N_29635,N_29309);
and UO_20 (O_20,N_29175,N_29080);
nor UO_21 (O_21,N_29894,N_29293);
or UO_22 (O_22,N_29796,N_29815);
and UO_23 (O_23,N_29798,N_29530);
xor UO_24 (O_24,N_29461,N_29633);
and UO_25 (O_25,N_29366,N_29835);
or UO_26 (O_26,N_29952,N_29017);
or UO_27 (O_27,N_29959,N_29501);
nand UO_28 (O_28,N_29662,N_29875);
nor UO_29 (O_29,N_29337,N_29715);
or UO_30 (O_30,N_29755,N_29620);
and UO_31 (O_31,N_29702,N_29383);
and UO_32 (O_32,N_29567,N_29216);
or UO_33 (O_33,N_29479,N_29699);
and UO_34 (O_34,N_29121,N_29586);
xnor UO_35 (O_35,N_29981,N_29521);
nand UO_36 (O_36,N_29068,N_29011);
or UO_37 (O_37,N_29616,N_29673);
and UO_38 (O_38,N_29628,N_29783);
and UO_39 (O_39,N_29667,N_29790);
nor UO_40 (O_40,N_29895,N_29097);
nor UO_41 (O_41,N_29523,N_29536);
and UO_42 (O_42,N_29693,N_29859);
or UO_43 (O_43,N_29529,N_29012);
or UO_44 (O_44,N_29075,N_29809);
or UO_45 (O_45,N_29283,N_29073);
nor UO_46 (O_46,N_29430,N_29558);
or UO_47 (O_47,N_29056,N_29050);
or UO_48 (O_48,N_29607,N_29574);
nor UO_49 (O_49,N_29769,N_29608);
and UO_50 (O_50,N_29497,N_29448);
and UO_51 (O_51,N_29191,N_29575);
and UO_52 (O_52,N_29065,N_29297);
nor UO_53 (O_53,N_29901,N_29524);
or UO_54 (O_54,N_29453,N_29552);
nor UO_55 (O_55,N_29989,N_29443);
xor UO_56 (O_56,N_29668,N_29014);
nor UO_57 (O_57,N_29236,N_29277);
xnor UO_58 (O_58,N_29577,N_29200);
and UO_59 (O_59,N_29039,N_29004);
and UO_60 (O_60,N_29446,N_29510);
nand UO_61 (O_61,N_29909,N_29108);
and UO_62 (O_62,N_29275,N_29889);
or UO_63 (O_63,N_29795,N_29849);
nor UO_64 (O_64,N_29131,N_29760);
or UO_65 (O_65,N_29793,N_29998);
nand UO_66 (O_66,N_29923,N_29520);
and UO_67 (O_67,N_29339,N_29058);
or UO_68 (O_68,N_29963,N_29541);
xnor UO_69 (O_69,N_29265,N_29001);
and UO_70 (O_70,N_29736,N_29797);
nor UO_71 (O_71,N_29462,N_29566);
nor UO_72 (O_72,N_29100,N_29109);
or UO_73 (O_73,N_29090,N_29215);
xor UO_74 (O_74,N_29550,N_29456);
and UO_75 (O_75,N_29880,N_29776);
nand UO_76 (O_76,N_29027,N_29999);
and UO_77 (O_77,N_29929,N_29931);
nor UO_78 (O_78,N_29554,N_29871);
or UO_79 (O_79,N_29762,N_29868);
nand UO_80 (O_80,N_29295,N_29799);
nor UO_81 (O_81,N_29500,N_29209);
nand UO_82 (O_82,N_29221,N_29840);
nor UO_83 (O_83,N_29107,N_29201);
nand UO_84 (O_84,N_29910,N_29086);
nor UO_85 (O_85,N_29245,N_29413);
nor UO_86 (O_86,N_29825,N_29143);
xnor UO_87 (O_87,N_29890,N_29691);
nor UO_88 (O_88,N_29846,N_29176);
xor UO_89 (O_89,N_29370,N_29393);
and UO_90 (O_90,N_29525,N_29274);
or UO_91 (O_91,N_29396,N_29344);
nand UO_92 (O_92,N_29332,N_29280);
or UO_93 (O_93,N_29938,N_29284);
nand UO_94 (O_94,N_29847,N_29390);
nand UO_95 (O_95,N_29626,N_29819);
xnor UO_96 (O_96,N_29331,N_29303);
or UO_97 (O_97,N_29737,N_29739);
and UO_98 (O_98,N_29007,N_29124);
and UO_99 (O_99,N_29666,N_29580);
nand UO_100 (O_100,N_29278,N_29489);
or UO_101 (O_101,N_29042,N_29873);
nor UO_102 (O_102,N_29092,N_29933);
nor UO_103 (O_103,N_29387,N_29672);
or UO_104 (O_104,N_29036,N_29758);
nand UO_105 (O_105,N_29692,N_29454);
or UO_106 (O_106,N_29881,N_29382);
or UO_107 (O_107,N_29624,N_29407);
nand UO_108 (O_108,N_29374,N_29937);
nand UO_109 (O_109,N_29634,N_29404);
nand UO_110 (O_110,N_29146,N_29917);
nand UO_111 (O_111,N_29709,N_29024);
or UO_112 (O_112,N_29202,N_29941);
and UO_113 (O_113,N_29333,N_29531);
and UO_114 (O_114,N_29887,N_29922);
and UO_115 (O_115,N_29855,N_29246);
and UO_116 (O_116,N_29677,N_29301);
nor UO_117 (O_117,N_29255,N_29350);
and UO_118 (O_118,N_29805,N_29439);
and UO_119 (O_119,N_29263,N_29152);
or UO_120 (O_120,N_29587,N_29729);
nand UO_121 (O_121,N_29779,N_29701);
and UO_122 (O_122,N_29903,N_29502);
xnor UO_123 (O_123,N_29877,N_29359);
and UO_124 (O_124,N_29507,N_29982);
nand UO_125 (O_125,N_29165,N_29064);
nand UO_126 (O_126,N_29576,N_29617);
or UO_127 (O_127,N_29071,N_29285);
or UO_128 (O_128,N_29774,N_29410);
xor UO_129 (O_129,N_29319,N_29182);
nand UO_130 (O_130,N_29091,N_29994);
nand UO_131 (O_131,N_29735,N_29082);
xor UO_132 (O_132,N_29426,N_29435);
nand UO_133 (O_133,N_29589,N_29351);
nand UO_134 (O_134,N_29179,N_29652);
nor UO_135 (O_135,N_29939,N_29979);
nand UO_136 (O_136,N_29025,N_29015);
xor UO_137 (O_137,N_29806,N_29824);
xnor UO_138 (O_138,N_29766,N_29708);
or UO_139 (O_139,N_29432,N_29487);
xnor UO_140 (O_140,N_29357,N_29679);
xnor UO_141 (O_141,N_29427,N_29096);
nor UO_142 (O_142,N_29338,N_29801);
nand UO_143 (O_143,N_29545,N_29988);
nand UO_144 (O_144,N_29271,N_29967);
nor UO_145 (O_145,N_29111,N_29335);
nand UO_146 (O_146,N_29786,N_29623);
and UO_147 (O_147,N_29643,N_29311);
nand UO_148 (O_148,N_29638,N_29680);
nand UO_149 (O_149,N_29112,N_29972);
or UO_150 (O_150,N_29640,N_29557);
or UO_151 (O_151,N_29342,N_29033);
or UO_152 (O_152,N_29389,N_29040);
or UO_153 (O_153,N_29993,N_29913);
or UO_154 (O_154,N_29379,N_29522);
or UO_155 (O_155,N_29914,N_29180);
nor UO_156 (O_156,N_29581,N_29018);
and UO_157 (O_157,N_29464,N_29340);
and UO_158 (O_158,N_29136,N_29060);
and UO_159 (O_159,N_29118,N_29892);
nand UO_160 (O_160,N_29526,N_29232);
nand UO_161 (O_161,N_29153,N_29714);
nand UO_162 (O_162,N_29141,N_29711);
xnor UO_163 (O_163,N_29838,N_29916);
or UO_164 (O_164,N_29388,N_29326);
or UO_165 (O_165,N_29544,N_29037);
nor UO_166 (O_166,N_29978,N_29261);
or UO_167 (O_167,N_29023,N_29005);
nand UO_168 (O_168,N_29866,N_29619);
and UO_169 (O_169,N_29578,N_29281);
or UO_170 (O_170,N_29764,N_29368);
nor UO_171 (O_171,N_29987,N_29885);
or UO_172 (O_172,N_29535,N_29647);
nor UO_173 (O_173,N_29116,N_29279);
or UO_174 (O_174,N_29605,N_29980);
xnor UO_175 (O_175,N_29163,N_29854);
nand UO_176 (O_176,N_29352,N_29227);
nand UO_177 (O_177,N_29807,N_29196);
or UO_178 (O_178,N_29595,N_29481);
or UO_179 (O_179,N_29782,N_29599);
nor UO_180 (O_180,N_29069,N_29564);
and UO_181 (O_181,N_29600,N_29676);
and UO_182 (O_182,N_29642,N_29241);
nand UO_183 (O_183,N_29164,N_29156);
nor UO_184 (O_184,N_29083,N_29513);
or UO_185 (O_185,N_29419,N_29114);
or UO_186 (O_186,N_29476,N_29334);
xnor UO_187 (O_187,N_29812,N_29899);
or UO_188 (O_188,N_29906,N_29035);
nand UO_189 (O_189,N_29170,N_29028);
nand UO_190 (O_190,N_29816,N_29716);
nor UO_191 (O_191,N_29829,N_29808);
nand UO_192 (O_192,N_29137,N_29920);
nor UO_193 (O_193,N_29690,N_29681);
and UO_194 (O_194,N_29898,N_29486);
or UO_195 (O_195,N_29444,N_29710);
and UO_196 (O_196,N_29474,N_29678);
and UO_197 (O_197,N_29343,N_29059);
nor UO_198 (O_198,N_29833,N_29328);
xnor UO_199 (O_199,N_29239,N_29294);
nor UO_200 (O_200,N_29115,N_29173);
and UO_201 (O_201,N_29395,N_29740);
and UO_202 (O_202,N_29252,N_29290);
xnor UO_203 (O_203,N_29752,N_29936);
and UO_204 (O_204,N_29992,N_29423);
xor UO_205 (O_205,N_29965,N_29912);
xor UO_206 (O_206,N_29433,N_29742);
nand UO_207 (O_207,N_29171,N_29450);
and UO_208 (O_208,N_29970,N_29306);
nand UO_209 (O_209,N_29579,N_29703);
xnor UO_210 (O_210,N_29921,N_29817);
or UO_211 (O_211,N_29416,N_29656);
and UO_212 (O_212,N_29957,N_29078);
xnor UO_213 (O_213,N_29897,N_29904);
xnor UO_214 (O_214,N_29128,N_29190);
and UO_215 (O_215,N_29251,N_29700);
xnor UO_216 (O_216,N_29494,N_29315);
nor UO_217 (O_217,N_29602,N_29590);
nor UO_218 (O_218,N_29573,N_29519);
and UO_219 (O_219,N_29373,N_29313);
and UO_220 (O_220,N_29414,N_29571);
xnor UO_221 (O_221,N_29888,N_29105);
nor UO_222 (O_222,N_29601,N_29365);
or UO_223 (O_223,N_29534,N_29951);
nand UO_224 (O_224,N_29103,N_29197);
xnor UO_225 (O_225,N_29650,N_29367);
xor UO_226 (O_226,N_29377,N_29355);
and UO_227 (O_227,N_29420,N_29759);
or UO_228 (O_228,N_29229,N_29858);
nand UO_229 (O_229,N_29428,N_29663);
and UO_230 (O_230,N_29768,N_29287);
xnor UO_231 (O_231,N_29654,N_29961);
nand UO_232 (O_232,N_29750,N_29498);
xnor UO_233 (O_233,N_29113,N_29145);
or UO_234 (O_234,N_29611,N_29482);
nor UO_235 (O_235,N_29689,N_29300);
nor UO_236 (O_236,N_29346,N_29496);
or UO_237 (O_237,N_29588,N_29276);
xnor UO_238 (O_238,N_29101,N_29353);
nand UO_239 (O_239,N_29259,N_29364);
or UO_240 (O_240,N_29598,N_29253);
nor UO_241 (O_241,N_29148,N_29956);
nand UO_242 (O_242,N_29597,N_29447);
xor UO_243 (O_243,N_29659,N_29771);
xnor UO_244 (O_244,N_29738,N_29528);
or UO_245 (O_245,N_29054,N_29562);
or UO_246 (O_246,N_29983,N_29509);
nand UO_247 (O_247,N_29038,N_29618);
xnor UO_248 (O_248,N_29424,N_29843);
xor UO_249 (O_249,N_29316,N_29325);
nor UO_250 (O_250,N_29770,N_29199);
or UO_251 (O_251,N_29804,N_29256);
nand UO_252 (O_252,N_29968,N_29748);
nand UO_253 (O_253,N_29286,N_29719);
nor UO_254 (O_254,N_29211,N_29845);
nand UO_255 (O_255,N_29052,N_29186);
nor UO_256 (O_256,N_29472,N_29264);
and UO_257 (O_257,N_29238,N_29606);
xor UO_258 (O_258,N_29363,N_29369);
nor UO_259 (O_259,N_29205,N_29753);
nor UO_260 (O_260,N_29403,N_29911);
or UO_261 (O_261,N_29347,N_29161);
nor UO_262 (O_262,N_29184,N_29220);
nand UO_263 (O_263,N_29198,N_29480);
nor UO_264 (O_264,N_29572,N_29627);
nor UO_265 (O_265,N_29234,N_29984);
and UO_266 (O_266,N_29225,N_29865);
and UO_267 (O_267,N_29094,N_29019);
nand UO_268 (O_268,N_29135,N_29088);
or UO_269 (O_269,N_29927,N_29953);
or UO_270 (O_270,N_29803,N_29151);
or UO_271 (O_271,N_29675,N_29948);
xnor UO_272 (O_272,N_29686,N_29749);
xor UO_273 (O_273,N_29954,N_29207);
nor UO_274 (O_274,N_29969,N_29731);
nand UO_275 (O_275,N_29990,N_29079);
nand UO_276 (O_276,N_29883,N_29418);
nor UO_277 (O_277,N_29412,N_29745);
nand UO_278 (O_278,N_29950,N_29734);
nor UO_279 (O_279,N_29049,N_29041);
or UO_280 (O_280,N_29537,N_29930);
nand UO_281 (O_281,N_29886,N_29026);
or UO_282 (O_282,N_29250,N_29884);
nand UO_283 (O_283,N_29584,N_29555);
xnor UO_284 (O_284,N_29072,N_29228);
nand UO_285 (O_285,N_29613,N_29077);
and UO_286 (O_286,N_29324,N_29104);
and UO_287 (O_287,N_29240,N_29070);
xor UO_288 (O_288,N_29178,N_29076);
nor UO_289 (O_289,N_29661,N_29000);
xor UO_290 (O_290,N_29973,N_29905);
xor UO_291 (O_291,N_29823,N_29784);
xor UO_292 (O_292,N_29591,N_29696);
nand UO_293 (O_293,N_29349,N_29637);
xnor UO_294 (O_294,N_29262,N_29051);
or UO_295 (O_295,N_29995,N_29682);
nand UO_296 (O_296,N_29378,N_29110);
nor UO_297 (O_297,N_29166,N_29030);
and UO_298 (O_298,N_29308,N_29991);
nor UO_299 (O_299,N_29943,N_29125);
xnor UO_300 (O_300,N_29106,N_29133);
xnor UO_301 (O_301,N_29438,N_29781);
xor UO_302 (O_302,N_29384,N_29460);
xor UO_303 (O_303,N_29397,N_29158);
and UO_304 (O_304,N_29095,N_29008);
nand UO_305 (O_305,N_29822,N_29401);
nor UO_306 (O_306,N_29465,N_29746);
nand UO_307 (O_307,N_29451,N_29399);
nor UO_308 (O_308,N_29836,N_29506);
or UO_309 (O_309,N_29830,N_29546);
nor UO_310 (O_310,N_29174,N_29757);
or UO_311 (O_311,N_29516,N_29569);
nor UO_312 (O_312,N_29664,N_29473);
and UO_313 (O_313,N_29067,N_29192);
and UO_314 (O_314,N_29788,N_29126);
and UO_315 (O_315,N_29687,N_29724);
nor UO_316 (O_316,N_29348,N_29674);
and UO_317 (O_317,N_29733,N_29499);
xor UO_318 (O_318,N_29168,N_29706);
or UO_319 (O_319,N_29458,N_29935);
or UO_320 (O_320,N_29955,N_29445);
nor UO_321 (O_321,N_29188,N_29794);
xnor UO_322 (O_322,N_29243,N_29778);
nor UO_323 (O_323,N_29312,N_29547);
nand UO_324 (O_324,N_29908,N_29518);
or UO_325 (O_325,N_29560,N_29467);
xor UO_326 (O_326,N_29155,N_29085);
xnor UO_327 (O_327,N_29213,N_29183);
or UO_328 (O_328,N_29940,N_29538);
nor UO_329 (O_329,N_29013,N_29400);
nor UO_330 (O_330,N_29341,N_29649);
xor UO_331 (O_331,N_29415,N_29360);
and UO_332 (O_332,N_29132,N_29127);
nor UO_333 (O_333,N_29744,N_29919);
nor UO_334 (O_334,N_29792,N_29612);
or UO_335 (O_335,N_29493,N_29632);
nor UO_336 (O_336,N_29032,N_29469);
xor UO_337 (O_337,N_29218,N_29775);
and UO_338 (O_338,N_29491,N_29977);
and UO_339 (O_339,N_29629,N_29247);
xor UO_340 (O_340,N_29470,N_29372);
or UO_341 (O_341,N_29206,N_29345);
xor UO_342 (O_342,N_29874,N_29842);
nand UO_343 (O_343,N_29485,N_29302);
or UO_344 (O_344,N_29697,N_29878);
nor UO_345 (O_345,N_29832,N_29140);
nand UO_346 (O_346,N_29305,N_29237);
xnor UO_347 (O_347,N_29645,N_29242);
nand UO_348 (O_348,N_29327,N_29532);
nor UO_349 (O_349,N_29648,N_29289);
and UO_350 (O_350,N_29893,N_29398);
or UO_351 (O_351,N_29828,N_29515);
or UO_352 (O_352,N_29665,N_29260);
and UO_353 (O_353,N_29021,N_29622);
xnor UO_354 (O_354,N_29743,N_29651);
nand UO_355 (O_355,N_29615,N_29639);
nor UO_356 (O_356,N_29570,N_29002);
nor UO_357 (O_357,N_29867,N_29046);
nor UO_358 (O_358,N_29483,N_29266);
and UO_359 (O_359,N_29636,N_29861);
nor UO_360 (O_360,N_29756,N_29212);
xor UO_361 (O_361,N_29820,N_29230);
or UO_362 (O_362,N_29031,N_29853);
nand UO_363 (O_363,N_29870,N_29655);
or UO_364 (O_364,N_29505,N_29226);
and UO_365 (O_365,N_29821,N_29120);
nor UO_366 (O_366,N_29958,N_29705);
or UO_367 (O_367,N_29291,N_29375);
nand UO_368 (O_368,N_29273,N_29542);
xor UO_369 (O_369,N_29789,N_29010);
nand UO_370 (O_370,N_29354,N_29203);
nor UO_371 (O_371,N_29975,N_29827);
nand UO_372 (O_372,N_29045,N_29857);
xnor UO_373 (O_373,N_29568,N_29869);
or UO_374 (O_374,N_29583,N_29685);
nand UO_375 (O_375,N_29436,N_29800);
or UO_376 (O_376,N_29997,N_29802);
xor UO_377 (O_377,N_29061,N_29891);
nand UO_378 (O_378,N_29763,N_29773);
nand UO_379 (O_379,N_29380,N_29863);
or UO_380 (O_380,N_29044,N_29925);
and UO_381 (O_381,N_29503,N_29310);
nor UO_382 (O_382,N_29296,N_29722);
and UO_383 (O_383,N_29455,N_29466);
and UO_384 (O_384,N_29814,N_29434);
xnor UO_385 (O_385,N_29376,N_29932);
xnor UO_386 (O_386,N_29093,N_29129);
nor UO_387 (O_387,N_29660,N_29694);
or UO_388 (O_388,N_29504,N_29723);
xnor UO_389 (O_389,N_29947,N_29712);
nand UO_390 (O_390,N_29195,N_29053);
nor UO_391 (O_391,N_29540,N_29900);
nor UO_392 (O_392,N_29066,N_29902);
xnor UO_393 (O_393,N_29646,N_29478);
and UO_394 (O_394,N_29726,N_29767);
or UO_395 (O_395,N_29425,N_29402);
or UO_396 (O_396,N_29217,N_29625);
or UO_397 (O_397,N_29329,N_29527);
nor UO_398 (O_398,N_29945,N_29813);
and UO_399 (O_399,N_29747,N_29918);
xor UO_400 (O_400,N_29644,N_29463);
nor UO_401 (O_401,N_29442,N_29475);
xor UO_402 (O_402,N_29150,N_29421);
nor UO_403 (O_403,N_29669,N_29971);
or UO_404 (O_404,N_29222,N_29429);
or UO_405 (O_405,N_29856,N_29394);
or UO_406 (O_406,N_29304,N_29728);
nand UO_407 (O_407,N_29417,N_29490);
xnor UO_408 (O_408,N_29089,N_29826);
nand UO_409 (O_409,N_29754,N_29139);
or UO_410 (O_410,N_29683,N_29254);
xor UO_411 (O_411,N_29055,N_29288);
or UO_412 (O_412,N_29449,N_29047);
nor UO_413 (O_413,N_29057,N_29553);
xnor UO_414 (O_414,N_29730,N_29322);
nor UO_415 (O_415,N_29603,N_29269);
xnor UO_416 (O_416,N_29621,N_29549);
nand UO_417 (O_417,N_29177,N_29468);
and UO_418 (O_418,N_29138,N_29944);
and UO_419 (O_419,N_29585,N_29698);
nor UO_420 (O_420,N_29543,N_29223);
or UO_421 (O_421,N_29864,N_29020);
nor UO_422 (O_422,N_29062,N_29713);
or UO_423 (O_423,N_29181,N_29249);
xnor UO_424 (O_424,N_29122,N_29172);
xnor UO_425 (O_425,N_29457,N_29048);
or UO_426 (O_426,N_29134,N_29193);
nand UO_427 (O_427,N_29362,N_29942);
xor UO_428 (O_428,N_29684,N_29811);
xor UO_429 (O_429,N_29081,N_29307);
nand UO_430 (O_430,N_29533,N_29986);
xnor UO_431 (O_431,N_29063,N_29386);
or UO_432 (O_432,N_29777,N_29022);
and UO_433 (O_433,N_29928,N_29610);
and UO_434 (O_434,N_29321,N_29556);
and UO_435 (O_435,N_29704,N_29772);
and UO_436 (O_436,N_29422,N_29144);
or UO_437 (O_437,N_29488,N_29946);
and UO_438 (O_438,N_29406,N_29671);
or UO_439 (O_439,N_29508,N_29219);
or UO_440 (O_440,N_29517,N_29976);
and UO_441 (O_441,N_29839,N_29851);
nor UO_442 (O_442,N_29741,N_29514);
nand UO_443 (O_443,N_29162,N_29119);
or UO_444 (O_444,N_29471,N_29224);
nor UO_445 (O_445,N_29160,N_29299);
and UO_446 (O_446,N_29159,N_29761);
or UO_447 (O_447,N_29582,N_29785);
xnor UO_448 (O_448,N_29604,N_29323);
xor UO_449 (O_449,N_29592,N_29765);
or UO_450 (O_450,N_29214,N_29102);
xnor UO_451 (O_451,N_29559,N_29431);
and UO_452 (O_452,N_29551,N_29985);
xor UO_453 (O_453,N_29872,N_29511);
xor UO_454 (O_454,N_29381,N_29248);
and UO_455 (O_455,N_29336,N_29477);
or UO_456 (O_456,N_29154,N_29670);
and UO_457 (O_457,N_29034,N_29029);
and UO_458 (O_458,N_29565,N_29043);
nor UO_459 (O_459,N_29356,N_29609);
or UO_460 (O_460,N_29441,N_29268);
nand UO_461 (O_461,N_29330,N_29657);
or UO_462 (O_462,N_29896,N_29147);
and UO_463 (O_463,N_29594,N_29512);
or UO_464 (O_464,N_29235,N_29966);
xor UO_465 (O_465,N_29934,N_29009);
nor UO_466 (O_466,N_29732,N_29907);
nand UO_467 (O_467,N_29142,N_29267);
nor UO_468 (O_468,N_29084,N_29317);
nor UO_469 (O_469,N_29492,N_29016);
or UO_470 (O_470,N_29539,N_29194);
xnor UO_471 (O_471,N_29852,N_29641);
nand UO_472 (O_472,N_29099,N_29862);
and UO_473 (O_473,N_29484,N_29292);
xnor UO_474 (O_474,N_29717,N_29721);
nand UO_475 (O_475,N_29725,N_29320);
nand UO_476 (O_476,N_29787,N_29006);
nor UO_477 (O_477,N_29860,N_29879);
nor UO_478 (O_478,N_29257,N_29361);
and UO_479 (O_479,N_29169,N_29962);
nand UO_480 (O_480,N_29074,N_29974);
nand UO_481 (O_481,N_29437,N_29149);
or UO_482 (O_482,N_29314,N_29831);
or UO_483 (O_483,N_29210,N_29882);
xnor UO_484 (O_484,N_29270,N_29810);
and UO_485 (O_485,N_29187,N_29208);
nand UO_486 (O_486,N_29003,N_29924);
or UO_487 (O_487,N_29452,N_29915);
nor UO_488 (O_488,N_29695,N_29298);
nor UO_489 (O_489,N_29358,N_29391);
and UO_490 (O_490,N_29614,N_29837);
nor UO_491 (O_491,N_29780,N_29841);
nor UO_492 (O_492,N_29409,N_29130);
xnor UO_493 (O_493,N_29318,N_29791);
nor UO_494 (O_494,N_29751,N_29157);
nand UO_495 (O_495,N_29563,N_29189);
and UO_496 (O_496,N_29233,N_29848);
or UO_497 (O_497,N_29258,N_29630);
or UO_498 (O_498,N_29411,N_29688);
nor UO_499 (O_499,N_29720,N_29834);
nand UO_500 (O_500,N_29745,N_29510);
xor UO_501 (O_501,N_29290,N_29748);
nand UO_502 (O_502,N_29090,N_29521);
and UO_503 (O_503,N_29377,N_29917);
nand UO_504 (O_504,N_29192,N_29178);
nand UO_505 (O_505,N_29986,N_29532);
nor UO_506 (O_506,N_29998,N_29365);
or UO_507 (O_507,N_29542,N_29310);
and UO_508 (O_508,N_29781,N_29638);
nor UO_509 (O_509,N_29661,N_29971);
and UO_510 (O_510,N_29117,N_29343);
nand UO_511 (O_511,N_29004,N_29205);
or UO_512 (O_512,N_29365,N_29559);
nor UO_513 (O_513,N_29409,N_29356);
and UO_514 (O_514,N_29341,N_29732);
nand UO_515 (O_515,N_29481,N_29148);
or UO_516 (O_516,N_29616,N_29315);
and UO_517 (O_517,N_29708,N_29877);
and UO_518 (O_518,N_29793,N_29865);
or UO_519 (O_519,N_29241,N_29189);
xor UO_520 (O_520,N_29545,N_29270);
xor UO_521 (O_521,N_29714,N_29098);
nand UO_522 (O_522,N_29312,N_29154);
nor UO_523 (O_523,N_29075,N_29342);
and UO_524 (O_524,N_29284,N_29017);
nand UO_525 (O_525,N_29338,N_29523);
nor UO_526 (O_526,N_29749,N_29254);
and UO_527 (O_527,N_29974,N_29523);
nand UO_528 (O_528,N_29038,N_29856);
xnor UO_529 (O_529,N_29670,N_29363);
nand UO_530 (O_530,N_29822,N_29738);
or UO_531 (O_531,N_29963,N_29544);
xnor UO_532 (O_532,N_29573,N_29740);
and UO_533 (O_533,N_29692,N_29278);
xor UO_534 (O_534,N_29358,N_29326);
and UO_535 (O_535,N_29816,N_29430);
or UO_536 (O_536,N_29731,N_29074);
xor UO_537 (O_537,N_29243,N_29714);
and UO_538 (O_538,N_29706,N_29128);
nor UO_539 (O_539,N_29637,N_29224);
nor UO_540 (O_540,N_29985,N_29949);
nor UO_541 (O_541,N_29967,N_29496);
and UO_542 (O_542,N_29204,N_29120);
nand UO_543 (O_543,N_29869,N_29852);
xnor UO_544 (O_544,N_29941,N_29427);
xor UO_545 (O_545,N_29464,N_29876);
nor UO_546 (O_546,N_29901,N_29990);
nand UO_547 (O_547,N_29351,N_29103);
or UO_548 (O_548,N_29489,N_29843);
nand UO_549 (O_549,N_29724,N_29031);
xor UO_550 (O_550,N_29865,N_29677);
and UO_551 (O_551,N_29744,N_29419);
nor UO_552 (O_552,N_29185,N_29568);
nand UO_553 (O_553,N_29088,N_29888);
nor UO_554 (O_554,N_29784,N_29710);
nor UO_555 (O_555,N_29211,N_29646);
xnor UO_556 (O_556,N_29862,N_29126);
xor UO_557 (O_557,N_29338,N_29443);
xor UO_558 (O_558,N_29758,N_29302);
xor UO_559 (O_559,N_29178,N_29092);
or UO_560 (O_560,N_29966,N_29560);
and UO_561 (O_561,N_29395,N_29058);
xnor UO_562 (O_562,N_29569,N_29404);
nor UO_563 (O_563,N_29136,N_29290);
nor UO_564 (O_564,N_29129,N_29775);
nand UO_565 (O_565,N_29068,N_29071);
xnor UO_566 (O_566,N_29568,N_29741);
and UO_567 (O_567,N_29516,N_29875);
xor UO_568 (O_568,N_29313,N_29868);
xnor UO_569 (O_569,N_29388,N_29992);
and UO_570 (O_570,N_29554,N_29210);
or UO_571 (O_571,N_29273,N_29289);
nand UO_572 (O_572,N_29081,N_29087);
nor UO_573 (O_573,N_29718,N_29288);
and UO_574 (O_574,N_29536,N_29410);
xor UO_575 (O_575,N_29694,N_29320);
nor UO_576 (O_576,N_29705,N_29093);
or UO_577 (O_577,N_29303,N_29759);
nor UO_578 (O_578,N_29606,N_29787);
or UO_579 (O_579,N_29415,N_29840);
or UO_580 (O_580,N_29738,N_29656);
xnor UO_581 (O_581,N_29427,N_29269);
or UO_582 (O_582,N_29942,N_29886);
nand UO_583 (O_583,N_29718,N_29737);
and UO_584 (O_584,N_29721,N_29456);
nor UO_585 (O_585,N_29844,N_29590);
nand UO_586 (O_586,N_29119,N_29989);
and UO_587 (O_587,N_29078,N_29996);
xor UO_588 (O_588,N_29211,N_29629);
nand UO_589 (O_589,N_29593,N_29355);
nand UO_590 (O_590,N_29401,N_29450);
nand UO_591 (O_591,N_29204,N_29751);
nand UO_592 (O_592,N_29388,N_29276);
or UO_593 (O_593,N_29257,N_29457);
and UO_594 (O_594,N_29809,N_29948);
nor UO_595 (O_595,N_29102,N_29543);
xor UO_596 (O_596,N_29261,N_29424);
nand UO_597 (O_597,N_29706,N_29032);
xor UO_598 (O_598,N_29882,N_29588);
or UO_599 (O_599,N_29265,N_29178);
nor UO_600 (O_600,N_29847,N_29168);
nor UO_601 (O_601,N_29368,N_29738);
nand UO_602 (O_602,N_29824,N_29657);
xnor UO_603 (O_603,N_29105,N_29083);
and UO_604 (O_604,N_29276,N_29189);
nand UO_605 (O_605,N_29024,N_29386);
xnor UO_606 (O_606,N_29516,N_29328);
and UO_607 (O_607,N_29499,N_29466);
or UO_608 (O_608,N_29622,N_29129);
xor UO_609 (O_609,N_29075,N_29336);
or UO_610 (O_610,N_29327,N_29959);
nor UO_611 (O_611,N_29673,N_29833);
nor UO_612 (O_612,N_29908,N_29183);
nand UO_613 (O_613,N_29830,N_29880);
or UO_614 (O_614,N_29698,N_29159);
or UO_615 (O_615,N_29680,N_29001);
or UO_616 (O_616,N_29890,N_29199);
nand UO_617 (O_617,N_29168,N_29534);
nor UO_618 (O_618,N_29299,N_29719);
xnor UO_619 (O_619,N_29181,N_29106);
and UO_620 (O_620,N_29733,N_29747);
or UO_621 (O_621,N_29045,N_29140);
nor UO_622 (O_622,N_29791,N_29565);
and UO_623 (O_623,N_29031,N_29658);
nor UO_624 (O_624,N_29262,N_29611);
or UO_625 (O_625,N_29174,N_29906);
and UO_626 (O_626,N_29110,N_29824);
nand UO_627 (O_627,N_29052,N_29909);
nor UO_628 (O_628,N_29445,N_29626);
nand UO_629 (O_629,N_29683,N_29253);
xor UO_630 (O_630,N_29096,N_29497);
and UO_631 (O_631,N_29024,N_29057);
and UO_632 (O_632,N_29835,N_29828);
xnor UO_633 (O_633,N_29556,N_29133);
nor UO_634 (O_634,N_29607,N_29844);
and UO_635 (O_635,N_29382,N_29921);
xor UO_636 (O_636,N_29258,N_29145);
nor UO_637 (O_637,N_29409,N_29437);
or UO_638 (O_638,N_29030,N_29298);
or UO_639 (O_639,N_29252,N_29258);
and UO_640 (O_640,N_29811,N_29049);
and UO_641 (O_641,N_29184,N_29559);
and UO_642 (O_642,N_29499,N_29314);
xnor UO_643 (O_643,N_29871,N_29169);
nand UO_644 (O_644,N_29675,N_29784);
and UO_645 (O_645,N_29226,N_29282);
nand UO_646 (O_646,N_29745,N_29193);
nand UO_647 (O_647,N_29529,N_29442);
and UO_648 (O_648,N_29880,N_29651);
nand UO_649 (O_649,N_29009,N_29345);
nor UO_650 (O_650,N_29988,N_29903);
nand UO_651 (O_651,N_29267,N_29588);
xor UO_652 (O_652,N_29291,N_29706);
nor UO_653 (O_653,N_29405,N_29074);
xor UO_654 (O_654,N_29563,N_29433);
xor UO_655 (O_655,N_29073,N_29426);
nor UO_656 (O_656,N_29486,N_29458);
or UO_657 (O_657,N_29089,N_29385);
xnor UO_658 (O_658,N_29786,N_29080);
nand UO_659 (O_659,N_29386,N_29219);
and UO_660 (O_660,N_29470,N_29960);
or UO_661 (O_661,N_29990,N_29406);
and UO_662 (O_662,N_29012,N_29779);
or UO_663 (O_663,N_29120,N_29504);
and UO_664 (O_664,N_29662,N_29846);
xor UO_665 (O_665,N_29546,N_29601);
nor UO_666 (O_666,N_29571,N_29897);
xnor UO_667 (O_667,N_29356,N_29242);
xor UO_668 (O_668,N_29922,N_29724);
xor UO_669 (O_669,N_29856,N_29769);
or UO_670 (O_670,N_29106,N_29620);
or UO_671 (O_671,N_29685,N_29455);
nor UO_672 (O_672,N_29485,N_29171);
nand UO_673 (O_673,N_29037,N_29175);
nand UO_674 (O_674,N_29018,N_29612);
nor UO_675 (O_675,N_29913,N_29710);
or UO_676 (O_676,N_29760,N_29896);
nor UO_677 (O_677,N_29434,N_29428);
and UO_678 (O_678,N_29829,N_29173);
xnor UO_679 (O_679,N_29585,N_29319);
or UO_680 (O_680,N_29169,N_29020);
xnor UO_681 (O_681,N_29922,N_29016);
nand UO_682 (O_682,N_29256,N_29879);
nand UO_683 (O_683,N_29208,N_29755);
nor UO_684 (O_684,N_29761,N_29415);
or UO_685 (O_685,N_29475,N_29722);
and UO_686 (O_686,N_29292,N_29750);
nor UO_687 (O_687,N_29560,N_29161);
nor UO_688 (O_688,N_29487,N_29874);
or UO_689 (O_689,N_29318,N_29307);
xor UO_690 (O_690,N_29903,N_29331);
nor UO_691 (O_691,N_29372,N_29373);
and UO_692 (O_692,N_29263,N_29236);
nor UO_693 (O_693,N_29770,N_29648);
xnor UO_694 (O_694,N_29072,N_29775);
nand UO_695 (O_695,N_29945,N_29733);
and UO_696 (O_696,N_29265,N_29617);
nor UO_697 (O_697,N_29547,N_29187);
or UO_698 (O_698,N_29823,N_29561);
or UO_699 (O_699,N_29253,N_29884);
xnor UO_700 (O_700,N_29776,N_29487);
nor UO_701 (O_701,N_29979,N_29632);
nor UO_702 (O_702,N_29041,N_29762);
or UO_703 (O_703,N_29211,N_29336);
or UO_704 (O_704,N_29957,N_29383);
xor UO_705 (O_705,N_29514,N_29415);
nand UO_706 (O_706,N_29798,N_29845);
or UO_707 (O_707,N_29260,N_29859);
and UO_708 (O_708,N_29109,N_29111);
xor UO_709 (O_709,N_29194,N_29355);
and UO_710 (O_710,N_29855,N_29485);
xnor UO_711 (O_711,N_29205,N_29134);
nand UO_712 (O_712,N_29488,N_29402);
or UO_713 (O_713,N_29471,N_29127);
and UO_714 (O_714,N_29188,N_29732);
nand UO_715 (O_715,N_29716,N_29108);
xor UO_716 (O_716,N_29877,N_29320);
nand UO_717 (O_717,N_29999,N_29148);
nor UO_718 (O_718,N_29789,N_29414);
nand UO_719 (O_719,N_29716,N_29663);
and UO_720 (O_720,N_29636,N_29614);
and UO_721 (O_721,N_29706,N_29571);
or UO_722 (O_722,N_29882,N_29796);
and UO_723 (O_723,N_29153,N_29402);
or UO_724 (O_724,N_29802,N_29331);
xor UO_725 (O_725,N_29568,N_29205);
nor UO_726 (O_726,N_29613,N_29522);
nand UO_727 (O_727,N_29035,N_29149);
nor UO_728 (O_728,N_29564,N_29872);
and UO_729 (O_729,N_29239,N_29002);
nand UO_730 (O_730,N_29011,N_29450);
or UO_731 (O_731,N_29622,N_29641);
or UO_732 (O_732,N_29806,N_29895);
and UO_733 (O_733,N_29250,N_29878);
nor UO_734 (O_734,N_29238,N_29472);
nand UO_735 (O_735,N_29840,N_29772);
xnor UO_736 (O_736,N_29081,N_29703);
or UO_737 (O_737,N_29681,N_29190);
nor UO_738 (O_738,N_29154,N_29217);
or UO_739 (O_739,N_29351,N_29979);
xnor UO_740 (O_740,N_29013,N_29607);
or UO_741 (O_741,N_29874,N_29212);
xnor UO_742 (O_742,N_29997,N_29827);
nor UO_743 (O_743,N_29478,N_29684);
nand UO_744 (O_744,N_29910,N_29567);
nor UO_745 (O_745,N_29362,N_29974);
and UO_746 (O_746,N_29760,N_29977);
or UO_747 (O_747,N_29653,N_29408);
and UO_748 (O_748,N_29832,N_29379);
nor UO_749 (O_749,N_29796,N_29051);
nor UO_750 (O_750,N_29032,N_29432);
and UO_751 (O_751,N_29284,N_29662);
and UO_752 (O_752,N_29978,N_29546);
nand UO_753 (O_753,N_29525,N_29658);
nor UO_754 (O_754,N_29328,N_29980);
xnor UO_755 (O_755,N_29528,N_29560);
or UO_756 (O_756,N_29535,N_29511);
or UO_757 (O_757,N_29941,N_29195);
and UO_758 (O_758,N_29511,N_29884);
nor UO_759 (O_759,N_29738,N_29852);
nor UO_760 (O_760,N_29263,N_29644);
nor UO_761 (O_761,N_29826,N_29489);
xnor UO_762 (O_762,N_29400,N_29466);
nand UO_763 (O_763,N_29421,N_29899);
xor UO_764 (O_764,N_29722,N_29487);
xor UO_765 (O_765,N_29154,N_29643);
or UO_766 (O_766,N_29835,N_29203);
and UO_767 (O_767,N_29035,N_29322);
nand UO_768 (O_768,N_29191,N_29555);
and UO_769 (O_769,N_29697,N_29574);
xnor UO_770 (O_770,N_29754,N_29844);
nand UO_771 (O_771,N_29280,N_29700);
and UO_772 (O_772,N_29172,N_29979);
or UO_773 (O_773,N_29948,N_29658);
nand UO_774 (O_774,N_29438,N_29617);
xnor UO_775 (O_775,N_29832,N_29718);
nand UO_776 (O_776,N_29961,N_29450);
or UO_777 (O_777,N_29242,N_29561);
or UO_778 (O_778,N_29180,N_29258);
or UO_779 (O_779,N_29051,N_29982);
nand UO_780 (O_780,N_29951,N_29877);
or UO_781 (O_781,N_29742,N_29973);
xnor UO_782 (O_782,N_29649,N_29017);
nor UO_783 (O_783,N_29953,N_29946);
and UO_784 (O_784,N_29487,N_29129);
and UO_785 (O_785,N_29246,N_29527);
nor UO_786 (O_786,N_29255,N_29312);
nor UO_787 (O_787,N_29649,N_29222);
xnor UO_788 (O_788,N_29012,N_29971);
or UO_789 (O_789,N_29642,N_29542);
and UO_790 (O_790,N_29852,N_29793);
nor UO_791 (O_791,N_29038,N_29360);
or UO_792 (O_792,N_29297,N_29598);
nor UO_793 (O_793,N_29016,N_29788);
and UO_794 (O_794,N_29047,N_29786);
nor UO_795 (O_795,N_29905,N_29960);
xor UO_796 (O_796,N_29073,N_29965);
nor UO_797 (O_797,N_29375,N_29475);
xor UO_798 (O_798,N_29810,N_29848);
nor UO_799 (O_799,N_29358,N_29206);
nand UO_800 (O_800,N_29891,N_29932);
xnor UO_801 (O_801,N_29054,N_29159);
nand UO_802 (O_802,N_29018,N_29163);
and UO_803 (O_803,N_29033,N_29471);
and UO_804 (O_804,N_29878,N_29486);
and UO_805 (O_805,N_29055,N_29534);
nand UO_806 (O_806,N_29891,N_29375);
nand UO_807 (O_807,N_29053,N_29641);
xnor UO_808 (O_808,N_29610,N_29401);
nor UO_809 (O_809,N_29489,N_29378);
nand UO_810 (O_810,N_29323,N_29706);
and UO_811 (O_811,N_29793,N_29476);
nand UO_812 (O_812,N_29519,N_29185);
or UO_813 (O_813,N_29366,N_29948);
or UO_814 (O_814,N_29142,N_29055);
xnor UO_815 (O_815,N_29277,N_29164);
and UO_816 (O_816,N_29000,N_29858);
nand UO_817 (O_817,N_29258,N_29916);
nand UO_818 (O_818,N_29393,N_29034);
and UO_819 (O_819,N_29355,N_29343);
nor UO_820 (O_820,N_29118,N_29256);
or UO_821 (O_821,N_29643,N_29529);
or UO_822 (O_822,N_29511,N_29413);
nand UO_823 (O_823,N_29584,N_29755);
and UO_824 (O_824,N_29338,N_29327);
nand UO_825 (O_825,N_29945,N_29428);
nand UO_826 (O_826,N_29731,N_29955);
or UO_827 (O_827,N_29949,N_29882);
nand UO_828 (O_828,N_29902,N_29007);
or UO_829 (O_829,N_29324,N_29224);
and UO_830 (O_830,N_29192,N_29334);
nand UO_831 (O_831,N_29132,N_29211);
and UO_832 (O_832,N_29816,N_29066);
or UO_833 (O_833,N_29732,N_29037);
xor UO_834 (O_834,N_29861,N_29342);
nand UO_835 (O_835,N_29086,N_29860);
xor UO_836 (O_836,N_29283,N_29724);
nor UO_837 (O_837,N_29867,N_29622);
or UO_838 (O_838,N_29626,N_29993);
or UO_839 (O_839,N_29840,N_29271);
nand UO_840 (O_840,N_29320,N_29160);
and UO_841 (O_841,N_29404,N_29352);
xor UO_842 (O_842,N_29611,N_29160);
nand UO_843 (O_843,N_29809,N_29153);
and UO_844 (O_844,N_29207,N_29604);
nor UO_845 (O_845,N_29617,N_29340);
xnor UO_846 (O_846,N_29035,N_29064);
or UO_847 (O_847,N_29397,N_29912);
xor UO_848 (O_848,N_29704,N_29857);
or UO_849 (O_849,N_29703,N_29050);
or UO_850 (O_850,N_29584,N_29760);
and UO_851 (O_851,N_29563,N_29017);
or UO_852 (O_852,N_29114,N_29403);
or UO_853 (O_853,N_29182,N_29451);
nor UO_854 (O_854,N_29923,N_29158);
or UO_855 (O_855,N_29801,N_29027);
nor UO_856 (O_856,N_29989,N_29381);
xor UO_857 (O_857,N_29732,N_29168);
nand UO_858 (O_858,N_29677,N_29148);
and UO_859 (O_859,N_29168,N_29910);
xnor UO_860 (O_860,N_29022,N_29140);
nor UO_861 (O_861,N_29909,N_29195);
or UO_862 (O_862,N_29160,N_29325);
xnor UO_863 (O_863,N_29307,N_29717);
and UO_864 (O_864,N_29178,N_29544);
nand UO_865 (O_865,N_29675,N_29707);
nand UO_866 (O_866,N_29039,N_29656);
and UO_867 (O_867,N_29901,N_29462);
xor UO_868 (O_868,N_29689,N_29667);
and UO_869 (O_869,N_29263,N_29807);
and UO_870 (O_870,N_29348,N_29840);
and UO_871 (O_871,N_29804,N_29747);
xor UO_872 (O_872,N_29397,N_29241);
or UO_873 (O_873,N_29431,N_29151);
nand UO_874 (O_874,N_29030,N_29319);
or UO_875 (O_875,N_29720,N_29468);
and UO_876 (O_876,N_29041,N_29799);
or UO_877 (O_877,N_29370,N_29290);
nor UO_878 (O_878,N_29501,N_29495);
xnor UO_879 (O_879,N_29846,N_29167);
xnor UO_880 (O_880,N_29096,N_29500);
nand UO_881 (O_881,N_29976,N_29027);
nand UO_882 (O_882,N_29875,N_29746);
and UO_883 (O_883,N_29187,N_29270);
nor UO_884 (O_884,N_29077,N_29710);
nor UO_885 (O_885,N_29722,N_29549);
and UO_886 (O_886,N_29064,N_29646);
nand UO_887 (O_887,N_29708,N_29761);
nand UO_888 (O_888,N_29717,N_29874);
nor UO_889 (O_889,N_29584,N_29744);
xnor UO_890 (O_890,N_29047,N_29520);
nor UO_891 (O_891,N_29122,N_29885);
and UO_892 (O_892,N_29618,N_29970);
nand UO_893 (O_893,N_29091,N_29397);
xor UO_894 (O_894,N_29655,N_29565);
and UO_895 (O_895,N_29204,N_29334);
nor UO_896 (O_896,N_29498,N_29608);
nand UO_897 (O_897,N_29395,N_29640);
nand UO_898 (O_898,N_29024,N_29264);
and UO_899 (O_899,N_29417,N_29966);
or UO_900 (O_900,N_29375,N_29316);
and UO_901 (O_901,N_29565,N_29889);
xnor UO_902 (O_902,N_29275,N_29370);
xnor UO_903 (O_903,N_29365,N_29862);
nor UO_904 (O_904,N_29283,N_29922);
xor UO_905 (O_905,N_29338,N_29571);
nor UO_906 (O_906,N_29251,N_29487);
and UO_907 (O_907,N_29712,N_29147);
xor UO_908 (O_908,N_29928,N_29600);
and UO_909 (O_909,N_29332,N_29800);
or UO_910 (O_910,N_29744,N_29504);
nor UO_911 (O_911,N_29167,N_29910);
nor UO_912 (O_912,N_29781,N_29579);
nor UO_913 (O_913,N_29488,N_29033);
xnor UO_914 (O_914,N_29202,N_29103);
xnor UO_915 (O_915,N_29049,N_29788);
and UO_916 (O_916,N_29384,N_29598);
and UO_917 (O_917,N_29591,N_29619);
nand UO_918 (O_918,N_29393,N_29837);
xnor UO_919 (O_919,N_29227,N_29031);
nor UO_920 (O_920,N_29657,N_29015);
nor UO_921 (O_921,N_29067,N_29802);
or UO_922 (O_922,N_29701,N_29824);
or UO_923 (O_923,N_29489,N_29148);
or UO_924 (O_924,N_29990,N_29118);
nand UO_925 (O_925,N_29920,N_29131);
and UO_926 (O_926,N_29835,N_29967);
nand UO_927 (O_927,N_29441,N_29458);
or UO_928 (O_928,N_29244,N_29906);
and UO_929 (O_929,N_29145,N_29856);
xor UO_930 (O_930,N_29073,N_29252);
or UO_931 (O_931,N_29925,N_29196);
and UO_932 (O_932,N_29082,N_29460);
xor UO_933 (O_933,N_29194,N_29516);
nand UO_934 (O_934,N_29403,N_29179);
and UO_935 (O_935,N_29962,N_29990);
or UO_936 (O_936,N_29771,N_29070);
nor UO_937 (O_937,N_29783,N_29076);
nor UO_938 (O_938,N_29404,N_29691);
and UO_939 (O_939,N_29254,N_29611);
and UO_940 (O_940,N_29452,N_29360);
and UO_941 (O_941,N_29780,N_29971);
nor UO_942 (O_942,N_29323,N_29852);
nand UO_943 (O_943,N_29779,N_29741);
nand UO_944 (O_944,N_29907,N_29727);
or UO_945 (O_945,N_29385,N_29778);
nor UO_946 (O_946,N_29271,N_29399);
nor UO_947 (O_947,N_29832,N_29914);
nor UO_948 (O_948,N_29899,N_29953);
nor UO_949 (O_949,N_29021,N_29369);
xnor UO_950 (O_950,N_29746,N_29893);
and UO_951 (O_951,N_29178,N_29429);
or UO_952 (O_952,N_29498,N_29278);
and UO_953 (O_953,N_29583,N_29491);
nor UO_954 (O_954,N_29237,N_29116);
or UO_955 (O_955,N_29379,N_29535);
xnor UO_956 (O_956,N_29319,N_29552);
or UO_957 (O_957,N_29972,N_29798);
and UO_958 (O_958,N_29333,N_29612);
xnor UO_959 (O_959,N_29747,N_29485);
nand UO_960 (O_960,N_29709,N_29573);
and UO_961 (O_961,N_29670,N_29163);
nor UO_962 (O_962,N_29747,N_29588);
nor UO_963 (O_963,N_29510,N_29811);
and UO_964 (O_964,N_29113,N_29426);
nor UO_965 (O_965,N_29948,N_29872);
and UO_966 (O_966,N_29920,N_29727);
and UO_967 (O_967,N_29137,N_29810);
nand UO_968 (O_968,N_29859,N_29004);
xnor UO_969 (O_969,N_29011,N_29445);
nor UO_970 (O_970,N_29254,N_29692);
xor UO_971 (O_971,N_29084,N_29686);
nand UO_972 (O_972,N_29246,N_29866);
nand UO_973 (O_973,N_29572,N_29176);
nor UO_974 (O_974,N_29947,N_29312);
xor UO_975 (O_975,N_29274,N_29996);
nor UO_976 (O_976,N_29735,N_29343);
xnor UO_977 (O_977,N_29539,N_29435);
or UO_978 (O_978,N_29312,N_29591);
and UO_979 (O_979,N_29473,N_29076);
nand UO_980 (O_980,N_29061,N_29763);
and UO_981 (O_981,N_29425,N_29426);
nor UO_982 (O_982,N_29962,N_29590);
or UO_983 (O_983,N_29563,N_29072);
nor UO_984 (O_984,N_29529,N_29120);
nor UO_985 (O_985,N_29279,N_29873);
and UO_986 (O_986,N_29542,N_29335);
nor UO_987 (O_987,N_29978,N_29312);
or UO_988 (O_988,N_29798,N_29840);
xor UO_989 (O_989,N_29628,N_29620);
nor UO_990 (O_990,N_29520,N_29523);
nand UO_991 (O_991,N_29656,N_29672);
or UO_992 (O_992,N_29497,N_29211);
nand UO_993 (O_993,N_29523,N_29145);
xor UO_994 (O_994,N_29827,N_29429);
and UO_995 (O_995,N_29461,N_29805);
or UO_996 (O_996,N_29293,N_29463);
or UO_997 (O_997,N_29272,N_29293);
and UO_998 (O_998,N_29812,N_29243);
and UO_999 (O_999,N_29914,N_29922);
or UO_1000 (O_1000,N_29692,N_29562);
xor UO_1001 (O_1001,N_29767,N_29801);
nand UO_1002 (O_1002,N_29018,N_29002);
nor UO_1003 (O_1003,N_29458,N_29693);
xnor UO_1004 (O_1004,N_29730,N_29996);
or UO_1005 (O_1005,N_29106,N_29395);
or UO_1006 (O_1006,N_29675,N_29267);
xnor UO_1007 (O_1007,N_29970,N_29984);
nand UO_1008 (O_1008,N_29991,N_29542);
nor UO_1009 (O_1009,N_29090,N_29459);
xnor UO_1010 (O_1010,N_29639,N_29486);
or UO_1011 (O_1011,N_29552,N_29858);
or UO_1012 (O_1012,N_29012,N_29369);
xnor UO_1013 (O_1013,N_29397,N_29538);
xor UO_1014 (O_1014,N_29833,N_29894);
xor UO_1015 (O_1015,N_29052,N_29614);
nand UO_1016 (O_1016,N_29532,N_29580);
and UO_1017 (O_1017,N_29835,N_29025);
xnor UO_1018 (O_1018,N_29922,N_29846);
or UO_1019 (O_1019,N_29372,N_29931);
nand UO_1020 (O_1020,N_29205,N_29337);
nor UO_1021 (O_1021,N_29440,N_29117);
xor UO_1022 (O_1022,N_29314,N_29072);
and UO_1023 (O_1023,N_29157,N_29290);
xnor UO_1024 (O_1024,N_29383,N_29182);
or UO_1025 (O_1025,N_29816,N_29116);
or UO_1026 (O_1026,N_29785,N_29200);
or UO_1027 (O_1027,N_29521,N_29769);
nor UO_1028 (O_1028,N_29034,N_29989);
xor UO_1029 (O_1029,N_29510,N_29260);
nand UO_1030 (O_1030,N_29994,N_29035);
and UO_1031 (O_1031,N_29465,N_29722);
xor UO_1032 (O_1032,N_29607,N_29913);
nor UO_1033 (O_1033,N_29846,N_29245);
nand UO_1034 (O_1034,N_29310,N_29274);
nand UO_1035 (O_1035,N_29657,N_29728);
and UO_1036 (O_1036,N_29996,N_29309);
xor UO_1037 (O_1037,N_29703,N_29362);
or UO_1038 (O_1038,N_29795,N_29049);
nor UO_1039 (O_1039,N_29680,N_29456);
or UO_1040 (O_1040,N_29930,N_29119);
xnor UO_1041 (O_1041,N_29679,N_29069);
xnor UO_1042 (O_1042,N_29068,N_29934);
xnor UO_1043 (O_1043,N_29741,N_29431);
nand UO_1044 (O_1044,N_29139,N_29239);
and UO_1045 (O_1045,N_29622,N_29887);
or UO_1046 (O_1046,N_29210,N_29020);
nand UO_1047 (O_1047,N_29621,N_29569);
xor UO_1048 (O_1048,N_29011,N_29805);
nand UO_1049 (O_1049,N_29682,N_29771);
or UO_1050 (O_1050,N_29474,N_29211);
or UO_1051 (O_1051,N_29277,N_29786);
and UO_1052 (O_1052,N_29764,N_29693);
nor UO_1053 (O_1053,N_29296,N_29733);
xor UO_1054 (O_1054,N_29327,N_29994);
xor UO_1055 (O_1055,N_29944,N_29049);
xnor UO_1056 (O_1056,N_29227,N_29070);
xnor UO_1057 (O_1057,N_29935,N_29387);
xor UO_1058 (O_1058,N_29632,N_29672);
xnor UO_1059 (O_1059,N_29506,N_29330);
and UO_1060 (O_1060,N_29186,N_29042);
xor UO_1061 (O_1061,N_29353,N_29515);
nor UO_1062 (O_1062,N_29369,N_29415);
and UO_1063 (O_1063,N_29270,N_29863);
or UO_1064 (O_1064,N_29044,N_29884);
nor UO_1065 (O_1065,N_29883,N_29797);
nand UO_1066 (O_1066,N_29270,N_29883);
nor UO_1067 (O_1067,N_29535,N_29616);
nor UO_1068 (O_1068,N_29634,N_29745);
nand UO_1069 (O_1069,N_29227,N_29606);
nor UO_1070 (O_1070,N_29201,N_29865);
nand UO_1071 (O_1071,N_29253,N_29174);
xnor UO_1072 (O_1072,N_29453,N_29499);
nand UO_1073 (O_1073,N_29598,N_29968);
or UO_1074 (O_1074,N_29850,N_29178);
xnor UO_1075 (O_1075,N_29647,N_29714);
xnor UO_1076 (O_1076,N_29464,N_29428);
nand UO_1077 (O_1077,N_29921,N_29154);
xnor UO_1078 (O_1078,N_29528,N_29593);
or UO_1079 (O_1079,N_29648,N_29288);
nor UO_1080 (O_1080,N_29571,N_29531);
and UO_1081 (O_1081,N_29969,N_29963);
xor UO_1082 (O_1082,N_29203,N_29914);
nor UO_1083 (O_1083,N_29528,N_29215);
or UO_1084 (O_1084,N_29118,N_29665);
nor UO_1085 (O_1085,N_29329,N_29624);
nand UO_1086 (O_1086,N_29871,N_29997);
nor UO_1087 (O_1087,N_29874,N_29265);
and UO_1088 (O_1088,N_29218,N_29064);
nor UO_1089 (O_1089,N_29008,N_29753);
nor UO_1090 (O_1090,N_29458,N_29508);
nor UO_1091 (O_1091,N_29855,N_29969);
or UO_1092 (O_1092,N_29426,N_29938);
nor UO_1093 (O_1093,N_29154,N_29280);
nand UO_1094 (O_1094,N_29498,N_29010);
nor UO_1095 (O_1095,N_29353,N_29390);
and UO_1096 (O_1096,N_29101,N_29210);
or UO_1097 (O_1097,N_29131,N_29909);
and UO_1098 (O_1098,N_29858,N_29966);
or UO_1099 (O_1099,N_29486,N_29215);
nor UO_1100 (O_1100,N_29560,N_29832);
xnor UO_1101 (O_1101,N_29836,N_29592);
or UO_1102 (O_1102,N_29611,N_29143);
and UO_1103 (O_1103,N_29145,N_29121);
or UO_1104 (O_1104,N_29207,N_29802);
xnor UO_1105 (O_1105,N_29477,N_29062);
and UO_1106 (O_1106,N_29689,N_29905);
nand UO_1107 (O_1107,N_29756,N_29041);
or UO_1108 (O_1108,N_29926,N_29846);
xnor UO_1109 (O_1109,N_29579,N_29995);
xnor UO_1110 (O_1110,N_29995,N_29244);
nor UO_1111 (O_1111,N_29092,N_29674);
nand UO_1112 (O_1112,N_29887,N_29438);
nand UO_1113 (O_1113,N_29203,N_29284);
nor UO_1114 (O_1114,N_29811,N_29108);
nor UO_1115 (O_1115,N_29207,N_29796);
and UO_1116 (O_1116,N_29530,N_29308);
and UO_1117 (O_1117,N_29697,N_29378);
or UO_1118 (O_1118,N_29122,N_29993);
nor UO_1119 (O_1119,N_29592,N_29187);
or UO_1120 (O_1120,N_29227,N_29027);
nand UO_1121 (O_1121,N_29230,N_29575);
and UO_1122 (O_1122,N_29392,N_29459);
xor UO_1123 (O_1123,N_29752,N_29194);
nand UO_1124 (O_1124,N_29323,N_29061);
xor UO_1125 (O_1125,N_29555,N_29297);
and UO_1126 (O_1126,N_29149,N_29414);
xnor UO_1127 (O_1127,N_29895,N_29589);
nand UO_1128 (O_1128,N_29121,N_29551);
and UO_1129 (O_1129,N_29651,N_29516);
nor UO_1130 (O_1130,N_29406,N_29002);
or UO_1131 (O_1131,N_29685,N_29280);
and UO_1132 (O_1132,N_29832,N_29640);
or UO_1133 (O_1133,N_29692,N_29141);
or UO_1134 (O_1134,N_29943,N_29426);
and UO_1135 (O_1135,N_29827,N_29527);
nand UO_1136 (O_1136,N_29478,N_29577);
or UO_1137 (O_1137,N_29581,N_29678);
nor UO_1138 (O_1138,N_29176,N_29555);
and UO_1139 (O_1139,N_29301,N_29377);
or UO_1140 (O_1140,N_29693,N_29739);
xor UO_1141 (O_1141,N_29317,N_29536);
xor UO_1142 (O_1142,N_29578,N_29165);
or UO_1143 (O_1143,N_29629,N_29068);
xnor UO_1144 (O_1144,N_29658,N_29079);
nand UO_1145 (O_1145,N_29675,N_29290);
nand UO_1146 (O_1146,N_29039,N_29138);
or UO_1147 (O_1147,N_29471,N_29516);
or UO_1148 (O_1148,N_29476,N_29801);
nand UO_1149 (O_1149,N_29510,N_29799);
nand UO_1150 (O_1150,N_29852,N_29992);
xnor UO_1151 (O_1151,N_29368,N_29230);
nand UO_1152 (O_1152,N_29589,N_29606);
xor UO_1153 (O_1153,N_29557,N_29718);
xor UO_1154 (O_1154,N_29215,N_29549);
nor UO_1155 (O_1155,N_29520,N_29549);
nand UO_1156 (O_1156,N_29481,N_29249);
or UO_1157 (O_1157,N_29725,N_29136);
and UO_1158 (O_1158,N_29396,N_29679);
or UO_1159 (O_1159,N_29273,N_29645);
and UO_1160 (O_1160,N_29805,N_29108);
nor UO_1161 (O_1161,N_29980,N_29504);
xor UO_1162 (O_1162,N_29675,N_29543);
xnor UO_1163 (O_1163,N_29703,N_29423);
or UO_1164 (O_1164,N_29400,N_29704);
or UO_1165 (O_1165,N_29131,N_29154);
or UO_1166 (O_1166,N_29070,N_29648);
or UO_1167 (O_1167,N_29376,N_29178);
nor UO_1168 (O_1168,N_29203,N_29408);
nor UO_1169 (O_1169,N_29502,N_29912);
and UO_1170 (O_1170,N_29743,N_29838);
and UO_1171 (O_1171,N_29832,N_29465);
or UO_1172 (O_1172,N_29575,N_29434);
or UO_1173 (O_1173,N_29818,N_29928);
or UO_1174 (O_1174,N_29608,N_29111);
xnor UO_1175 (O_1175,N_29698,N_29431);
or UO_1176 (O_1176,N_29049,N_29446);
or UO_1177 (O_1177,N_29017,N_29409);
nand UO_1178 (O_1178,N_29588,N_29093);
nand UO_1179 (O_1179,N_29795,N_29395);
or UO_1180 (O_1180,N_29279,N_29676);
xnor UO_1181 (O_1181,N_29780,N_29056);
and UO_1182 (O_1182,N_29725,N_29475);
or UO_1183 (O_1183,N_29709,N_29718);
xnor UO_1184 (O_1184,N_29609,N_29860);
nor UO_1185 (O_1185,N_29600,N_29547);
xor UO_1186 (O_1186,N_29606,N_29242);
and UO_1187 (O_1187,N_29946,N_29507);
and UO_1188 (O_1188,N_29237,N_29043);
xor UO_1189 (O_1189,N_29982,N_29912);
nand UO_1190 (O_1190,N_29254,N_29313);
or UO_1191 (O_1191,N_29057,N_29538);
nand UO_1192 (O_1192,N_29588,N_29877);
or UO_1193 (O_1193,N_29988,N_29694);
nand UO_1194 (O_1194,N_29003,N_29656);
or UO_1195 (O_1195,N_29535,N_29414);
and UO_1196 (O_1196,N_29270,N_29165);
xnor UO_1197 (O_1197,N_29506,N_29058);
or UO_1198 (O_1198,N_29761,N_29140);
nand UO_1199 (O_1199,N_29463,N_29634);
or UO_1200 (O_1200,N_29619,N_29558);
nor UO_1201 (O_1201,N_29587,N_29816);
xor UO_1202 (O_1202,N_29364,N_29174);
xor UO_1203 (O_1203,N_29766,N_29957);
xor UO_1204 (O_1204,N_29658,N_29832);
xnor UO_1205 (O_1205,N_29413,N_29891);
nor UO_1206 (O_1206,N_29696,N_29491);
xor UO_1207 (O_1207,N_29644,N_29130);
and UO_1208 (O_1208,N_29542,N_29340);
or UO_1209 (O_1209,N_29697,N_29344);
xnor UO_1210 (O_1210,N_29499,N_29798);
and UO_1211 (O_1211,N_29804,N_29219);
xnor UO_1212 (O_1212,N_29999,N_29900);
or UO_1213 (O_1213,N_29351,N_29026);
xor UO_1214 (O_1214,N_29002,N_29156);
xor UO_1215 (O_1215,N_29534,N_29628);
nor UO_1216 (O_1216,N_29729,N_29284);
or UO_1217 (O_1217,N_29253,N_29279);
nand UO_1218 (O_1218,N_29617,N_29436);
nand UO_1219 (O_1219,N_29129,N_29203);
and UO_1220 (O_1220,N_29906,N_29352);
nor UO_1221 (O_1221,N_29778,N_29974);
or UO_1222 (O_1222,N_29292,N_29334);
nand UO_1223 (O_1223,N_29115,N_29910);
nand UO_1224 (O_1224,N_29097,N_29965);
nor UO_1225 (O_1225,N_29383,N_29519);
nand UO_1226 (O_1226,N_29348,N_29509);
or UO_1227 (O_1227,N_29283,N_29404);
nand UO_1228 (O_1228,N_29074,N_29817);
nand UO_1229 (O_1229,N_29397,N_29443);
and UO_1230 (O_1230,N_29131,N_29751);
nor UO_1231 (O_1231,N_29080,N_29045);
and UO_1232 (O_1232,N_29626,N_29541);
xnor UO_1233 (O_1233,N_29434,N_29198);
nor UO_1234 (O_1234,N_29761,N_29859);
nand UO_1235 (O_1235,N_29873,N_29136);
or UO_1236 (O_1236,N_29608,N_29616);
or UO_1237 (O_1237,N_29938,N_29788);
and UO_1238 (O_1238,N_29976,N_29530);
and UO_1239 (O_1239,N_29280,N_29013);
nor UO_1240 (O_1240,N_29553,N_29892);
xnor UO_1241 (O_1241,N_29796,N_29541);
or UO_1242 (O_1242,N_29429,N_29417);
nor UO_1243 (O_1243,N_29448,N_29352);
or UO_1244 (O_1244,N_29098,N_29089);
xor UO_1245 (O_1245,N_29753,N_29979);
xnor UO_1246 (O_1246,N_29155,N_29200);
and UO_1247 (O_1247,N_29309,N_29802);
and UO_1248 (O_1248,N_29266,N_29841);
xor UO_1249 (O_1249,N_29273,N_29387);
and UO_1250 (O_1250,N_29219,N_29490);
nor UO_1251 (O_1251,N_29161,N_29675);
and UO_1252 (O_1252,N_29592,N_29316);
xnor UO_1253 (O_1253,N_29502,N_29754);
xnor UO_1254 (O_1254,N_29589,N_29668);
and UO_1255 (O_1255,N_29026,N_29221);
nor UO_1256 (O_1256,N_29050,N_29413);
nand UO_1257 (O_1257,N_29375,N_29954);
nand UO_1258 (O_1258,N_29246,N_29834);
nor UO_1259 (O_1259,N_29202,N_29468);
or UO_1260 (O_1260,N_29675,N_29619);
and UO_1261 (O_1261,N_29880,N_29355);
nor UO_1262 (O_1262,N_29100,N_29276);
and UO_1263 (O_1263,N_29800,N_29529);
and UO_1264 (O_1264,N_29040,N_29510);
xnor UO_1265 (O_1265,N_29691,N_29288);
xnor UO_1266 (O_1266,N_29643,N_29362);
nand UO_1267 (O_1267,N_29123,N_29523);
xnor UO_1268 (O_1268,N_29708,N_29924);
nand UO_1269 (O_1269,N_29771,N_29560);
xor UO_1270 (O_1270,N_29793,N_29908);
or UO_1271 (O_1271,N_29103,N_29552);
nand UO_1272 (O_1272,N_29321,N_29198);
nand UO_1273 (O_1273,N_29354,N_29938);
nor UO_1274 (O_1274,N_29022,N_29685);
xor UO_1275 (O_1275,N_29656,N_29222);
nor UO_1276 (O_1276,N_29641,N_29292);
or UO_1277 (O_1277,N_29340,N_29990);
nand UO_1278 (O_1278,N_29137,N_29455);
xor UO_1279 (O_1279,N_29328,N_29661);
and UO_1280 (O_1280,N_29542,N_29501);
or UO_1281 (O_1281,N_29084,N_29029);
xor UO_1282 (O_1282,N_29407,N_29950);
nand UO_1283 (O_1283,N_29932,N_29803);
and UO_1284 (O_1284,N_29247,N_29211);
xor UO_1285 (O_1285,N_29886,N_29511);
nand UO_1286 (O_1286,N_29720,N_29068);
nor UO_1287 (O_1287,N_29615,N_29966);
and UO_1288 (O_1288,N_29533,N_29149);
xnor UO_1289 (O_1289,N_29346,N_29008);
nor UO_1290 (O_1290,N_29292,N_29518);
and UO_1291 (O_1291,N_29339,N_29293);
nor UO_1292 (O_1292,N_29436,N_29359);
and UO_1293 (O_1293,N_29601,N_29554);
nor UO_1294 (O_1294,N_29397,N_29379);
nand UO_1295 (O_1295,N_29602,N_29700);
nand UO_1296 (O_1296,N_29885,N_29622);
or UO_1297 (O_1297,N_29278,N_29553);
or UO_1298 (O_1298,N_29057,N_29243);
nand UO_1299 (O_1299,N_29637,N_29693);
and UO_1300 (O_1300,N_29700,N_29188);
and UO_1301 (O_1301,N_29736,N_29080);
and UO_1302 (O_1302,N_29034,N_29925);
nor UO_1303 (O_1303,N_29756,N_29765);
and UO_1304 (O_1304,N_29209,N_29027);
xor UO_1305 (O_1305,N_29112,N_29768);
nor UO_1306 (O_1306,N_29036,N_29178);
and UO_1307 (O_1307,N_29747,N_29177);
nor UO_1308 (O_1308,N_29883,N_29215);
or UO_1309 (O_1309,N_29481,N_29791);
or UO_1310 (O_1310,N_29619,N_29347);
nand UO_1311 (O_1311,N_29117,N_29493);
nor UO_1312 (O_1312,N_29185,N_29000);
xnor UO_1313 (O_1313,N_29026,N_29673);
or UO_1314 (O_1314,N_29572,N_29581);
or UO_1315 (O_1315,N_29791,N_29108);
nor UO_1316 (O_1316,N_29411,N_29485);
nand UO_1317 (O_1317,N_29405,N_29051);
and UO_1318 (O_1318,N_29442,N_29908);
and UO_1319 (O_1319,N_29704,N_29005);
nand UO_1320 (O_1320,N_29764,N_29220);
or UO_1321 (O_1321,N_29169,N_29523);
xnor UO_1322 (O_1322,N_29937,N_29203);
or UO_1323 (O_1323,N_29672,N_29386);
nor UO_1324 (O_1324,N_29706,N_29182);
nand UO_1325 (O_1325,N_29045,N_29513);
and UO_1326 (O_1326,N_29112,N_29336);
xor UO_1327 (O_1327,N_29764,N_29058);
nand UO_1328 (O_1328,N_29298,N_29314);
nand UO_1329 (O_1329,N_29788,N_29129);
or UO_1330 (O_1330,N_29082,N_29224);
or UO_1331 (O_1331,N_29649,N_29234);
or UO_1332 (O_1332,N_29468,N_29318);
and UO_1333 (O_1333,N_29072,N_29826);
nand UO_1334 (O_1334,N_29539,N_29289);
xor UO_1335 (O_1335,N_29926,N_29119);
and UO_1336 (O_1336,N_29613,N_29215);
or UO_1337 (O_1337,N_29689,N_29101);
xnor UO_1338 (O_1338,N_29776,N_29360);
nor UO_1339 (O_1339,N_29726,N_29906);
and UO_1340 (O_1340,N_29679,N_29568);
and UO_1341 (O_1341,N_29927,N_29460);
or UO_1342 (O_1342,N_29844,N_29132);
nor UO_1343 (O_1343,N_29068,N_29205);
nor UO_1344 (O_1344,N_29339,N_29108);
nand UO_1345 (O_1345,N_29177,N_29158);
nand UO_1346 (O_1346,N_29723,N_29782);
and UO_1347 (O_1347,N_29963,N_29394);
or UO_1348 (O_1348,N_29047,N_29023);
xor UO_1349 (O_1349,N_29163,N_29195);
or UO_1350 (O_1350,N_29684,N_29377);
and UO_1351 (O_1351,N_29949,N_29648);
xor UO_1352 (O_1352,N_29992,N_29337);
or UO_1353 (O_1353,N_29607,N_29215);
or UO_1354 (O_1354,N_29679,N_29297);
nand UO_1355 (O_1355,N_29097,N_29708);
nand UO_1356 (O_1356,N_29533,N_29102);
xor UO_1357 (O_1357,N_29353,N_29064);
or UO_1358 (O_1358,N_29849,N_29137);
nand UO_1359 (O_1359,N_29202,N_29999);
nand UO_1360 (O_1360,N_29632,N_29895);
xor UO_1361 (O_1361,N_29743,N_29160);
nor UO_1362 (O_1362,N_29456,N_29064);
or UO_1363 (O_1363,N_29327,N_29810);
nor UO_1364 (O_1364,N_29218,N_29424);
xnor UO_1365 (O_1365,N_29265,N_29341);
and UO_1366 (O_1366,N_29908,N_29960);
or UO_1367 (O_1367,N_29628,N_29693);
and UO_1368 (O_1368,N_29533,N_29359);
nand UO_1369 (O_1369,N_29116,N_29443);
and UO_1370 (O_1370,N_29668,N_29743);
nand UO_1371 (O_1371,N_29943,N_29626);
or UO_1372 (O_1372,N_29097,N_29903);
nor UO_1373 (O_1373,N_29305,N_29287);
or UO_1374 (O_1374,N_29992,N_29554);
or UO_1375 (O_1375,N_29817,N_29750);
or UO_1376 (O_1376,N_29757,N_29717);
xor UO_1377 (O_1377,N_29340,N_29905);
nand UO_1378 (O_1378,N_29919,N_29700);
xnor UO_1379 (O_1379,N_29018,N_29671);
nand UO_1380 (O_1380,N_29955,N_29705);
and UO_1381 (O_1381,N_29285,N_29150);
and UO_1382 (O_1382,N_29662,N_29159);
or UO_1383 (O_1383,N_29302,N_29457);
and UO_1384 (O_1384,N_29143,N_29139);
xnor UO_1385 (O_1385,N_29972,N_29380);
xnor UO_1386 (O_1386,N_29890,N_29758);
nand UO_1387 (O_1387,N_29923,N_29064);
nor UO_1388 (O_1388,N_29673,N_29596);
or UO_1389 (O_1389,N_29147,N_29676);
xor UO_1390 (O_1390,N_29977,N_29704);
nor UO_1391 (O_1391,N_29180,N_29957);
or UO_1392 (O_1392,N_29810,N_29267);
nor UO_1393 (O_1393,N_29230,N_29588);
or UO_1394 (O_1394,N_29865,N_29506);
or UO_1395 (O_1395,N_29667,N_29035);
nand UO_1396 (O_1396,N_29896,N_29486);
and UO_1397 (O_1397,N_29212,N_29720);
nor UO_1398 (O_1398,N_29537,N_29387);
or UO_1399 (O_1399,N_29735,N_29321);
xor UO_1400 (O_1400,N_29442,N_29926);
and UO_1401 (O_1401,N_29272,N_29170);
nor UO_1402 (O_1402,N_29872,N_29611);
and UO_1403 (O_1403,N_29422,N_29856);
xor UO_1404 (O_1404,N_29105,N_29667);
and UO_1405 (O_1405,N_29835,N_29150);
xnor UO_1406 (O_1406,N_29314,N_29418);
or UO_1407 (O_1407,N_29032,N_29633);
xor UO_1408 (O_1408,N_29587,N_29910);
nor UO_1409 (O_1409,N_29423,N_29481);
nor UO_1410 (O_1410,N_29825,N_29903);
or UO_1411 (O_1411,N_29014,N_29044);
xor UO_1412 (O_1412,N_29025,N_29887);
nand UO_1413 (O_1413,N_29681,N_29464);
or UO_1414 (O_1414,N_29024,N_29668);
nor UO_1415 (O_1415,N_29764,N_29386);
or UO_1416 (O_1416,N_29400,N_29538);
and UO_1417 (O_1417,N_29224,N_29627);
nand UO_1418 (O_1418,N_29405,N_29846);
nand UO_1419 (O_1419,N_29893,N_29119);
xor UO_1420 (O_1420,N_29069,N_29237);
nor UO_1421 (O_1421,N_29937,N_29341);
nor UO_1422 (O_1422,N_29069,N_29454);
nor UO_1423 (O_1423,N_29442,N_29727);
nor UO_1424 (O_1424,N_29855,N_29912);
and UO_1425 (O_1425,N_29587,N_29514);
xnor UO_1426 (O_1426,N_29228,N_29360);
xor UO_1427 (O_1427,N_29019,N_29639);
and UO_1428 (O_1428,N_29449,N_29863);
nor UO_1429 (O_1429,N_29454,N_29443);
nor UO_1430 (O_1430,N_29149,N_29085);
nand UO_1431 (O_1431,N_29166,N_29508);
nor UO_1432 (O_1432,N_29881,N_29744);
nor UO_1433 (O_1433,N_29553,N_29608);
and UO_1434 (O_1434,N_29638,N_29681);
nand UO_1435 (O_1435,N_29410,N_29325);
nand UO_1436 (O_1436,N_29928,N_29141);
nor UO_1437 (O_1437,N_29829,N_29727);
and UO_1438 (O_1438,N_29681,N_29879);
xnor UO_1439 (O_1439,N_29321,N_29924);
or UO_1440 (O_1440,N_29497,N_29631);
xnor UO_1441 (O_1441,N_29674,N_29225);
and UO_1442 (O_1442,N_29117,N_29958);
nand UO_1443 (O_1443,N_29781,N_29934);
nor UO_1444 (O_1444,N_29895,N_29416);
and UO_1445 (O_1445,N_29262,N_29883);
nor UO_1446 (O_1446,N_29993,N_29596);
nor UO_1447 (O_1447,N_29275,N_29371);
or UO_1448 (O_1448,N_29572,N_29979);
xor UO_1449 (O_1449,N_29196,N_29202);
xor UO_1450 (O_1450,N_29326,N_29439);
and UO_1451 (O_1451,N_29260,N_29105);
and UO_1452 (O_1452,N_29850,N_29891);
nand UO_1453 (O_1453,N_29489,N_29481);
nand UO_1454 (O_1454,N_29571,N_29317);
nor UO_1455 (O_1455,N_29569,N_29870);
and UO_1456 (O_1456,N_29564,N_29337);
xnor UO_1457 (O_1457,N_29861,N_29052);
xnor UO_1458 (O_1458,N_29121,N_29842);
nand UO_1459 (O_1459,N_29574,N_29358);
and UO_1460 (O_1460,N_29047,N_29719);
nor UO_1461 (O_1461,N_29331,N_29985);
and UO_1462 (O_1462,N_29471,N_29487);
nand UO_1463 (O_1463,N_29530,N_29884);
nand UO_1464 (O_1464,N_29187,N_29192);
nand UO_1465 (O_1465,N_29119,N_29554);
xor UO_1466 (O_1466,N_29942,N_29642);
and UO_1467 (O_1467,N_29555,N_29604);
nor UO_1468 (O_1468,N_29601,N_29062);
nand UO_1469 (O_1469,N_29463,N_29167);
nand UO_1470 (O_1470,N_29078,N_29566);
and UO_1471 (O_1471,N_29482,N_29689);
or UO_1472 (O_1472,N_29637,N_29621);
xnor UO_1473 (O_1473,N_29217,N_29562);
and UO_1474 (O_1474,N_29513,N_29429);
nor UO_1475 (O_1475,N_29520,N_29504);
xnor UO_1476 (O_1476,N_29360,N_29516);
nor UO_1477 (O_1477,N_29869,N_29157);
and UO_1478 (O_1478,N_29229,N_29662);
and UO_1479 (O_1479,N_29009,N_29585);
or UO_1480 (O_1480,N_29192,N_29009);
nor UO_1481 (O_1481,N_29495,N_29718);
or UO_1482 (O_1482,N_29193,N_29053);
nor UO_1483 (O_1483,N_29029,N_29798);
or UO_1484 (O_1484,N_29126,N_29362);
nand UO_1485 (O_1485,N_29477,N_29849);
nand UO_1486 (O_1486,N_29588,N_29250);
or UO_1487 (O_1487,N_29198,N_29140);
nor UO_1488 (O_1488,N_29541,N_29580);
or UO_1489 (O_1489,N_29034,N_29951);
xor UO_1490 (O_1490,N_29206,N_29802);
nor UO_1491 (O_1491,N_29400,N_29215);
or UO_1492 (O_1492,N_29017,N_29592);
nor UO_1493 (O_1493,N_29769,N_29859);
xnor UO_1494 (O_1494,N_29281,N_29492);
or UO_1495 (O_1495,N_29538,N_29864);
or UO_1496 (O_1496,N_29320,N_29025);
nand UO_1497 (O_1497,N_29578,N_29721);
xor UO_1498 (O_1498,N_29794,N_29293);
nor UO_1499 (O_1499,N_29664,N_29123);
or UO_1500 (O_1500,N_29232,N_29338);
nand UO_1501 (O_1501,N_29727,N_29510);
nand UO_1502 (O_1502,N_29938,N_29814);
and UO_1503 (O_1503,N_29479,N_29352);
nor UO_1504 (O_1504,N_29084,N_29614);
nand UO_1505 (O_1505,N_29696,N_29761);
nand UO_1506 (O_1506,N_29218,N_29423);
nand UO_1507 (O_1507,N_29373,N_29432);
and UO_1508 (O_1508,N_29878,N_29532);
nand UO_1509 (O_1509,N_29280,N_29955);
nand UO_1510 (O_1510,N_29761,N_29447);
nor UO_1511 (O_1511,N_29674,N_29849);
nor UO_1512 (O_1512,N_29634,N_29137);
xnor UO_1513 (O_1513,N_29926,N_29323);
or UO_1514 (O_1514,N_29074,N_29398);
nand UO_1515 (O_1515,N_29234,N_29587);
nor UO_1516 (O_1516,N_29137,N_29071);
xor UO_1517 (O_1517,N_29876,N_29591);
or UO_1518 (O_1518,N_29873,N_29172);
xnor UO_1519 (O_1519,N_29864,N_29866);
nand UO_1520 (O_1520,N_29013,N_29177);
and UO_1521 (O_1521,N_29274,N_29857);
or UO_1522 (O_1522,N_29305,N_29450);
nor UO_1523 (O_1523,N_29037,N_29077);
and UO_1524 (O_1524,N_29701,N_29836);
xor UO_1525 (O_1525,N_29663,N_29519);
and UO_1526 (O_1526,N_29675,N_29366);
and UO_1527 (O_1527,N_29275,N_29738);
nand UO_1528 (O_1528,N_29290,N_29967);
and UO_1529 (O_1529,N_29925,N_29911);
nor UO_1530 (O_1530,N_29315,N_29252);
and UO_1531 (O_1531,N_29968,N_29799);
and UO_1532 (O_1532,N_29153,N_29590);
and UO_1533 (O_1533,N_29757,N_29989);
and UO_1534 (O_1534,N_29133,N_29393);
xnor UO_1535 (O_1535,N_29018,N_29131);
xor UO_1536 (O_1536,N_29728,N_29528);
nor UO_1537 (O_1537,N_29067,N_29268);
nor UO_1538 (O_1538,N_29870,N_29952);
nor UO_1539 (O_1539,N_29649,N_29386);
nor UO_1540 (O_1540,N_29085,N_29419);
or UO_1541 (O_1541,N_29726,N_29719);
and UO_1542 (O_1542,N_29162,N_29403);
and UO_1543 (O_1543,N_29658,N_29737);
nand UO_1544 (O_1544,N_29548,N_29355);
or UO_1545 (O_1545,N_29274,N_29273);
nor UO_1546 (O_1546,N_29265,N_29895);
xor UO_1547 (O_1547,N_29850,N_29941);
nand UO_1548 (O_1548,N_29677,N_29609);
nand UO_1549 (O_1549,N_29571,N_29814);
nor UO_1550 (O_1550,N_29357,N_29908);
or UO_1551 (O_1551,N_29644,N_29896);
and UO_1552 (O_1552,N_29546,N_29114);
nand UO_1553 (O_1553,N_29832,N_29654);
or UO_1554 (O_1554,N_29243,N_29854);
or UO_1555 (O_1555,N_29522,N_29479);
nand UO_1556 (O_1556,N_29563,N_29700);
nor UO_1557 (O_1557,N_29704,N_29175);
nor UO_1558 (O_1558,N_29029,N_29987);
and UO_1559 (O_1559,N_29018,N_29773);
nor UO_1560 (O_1560,N_29031,N_29931);
nand UO_1561 (O_1561,N_29645,N_29419);
or UO_1562 (O_1562,N_29408,N_29711);
nand UO_1563 (O_1563,N_29055,N_29759);
or UO_1564 (O_1564,N_29294,N_29829);
xor UO_1565 (O_1565,N_29659,N_29926);
and UO_1566 (O_1566,N_29867,N_29059);
xnor UO_1567 (O_1567,N_29009,N_29270);
nand UO_1568 (O_1568,N_29085,N_29139);
xnor UO_1569 (O_1569,N_29975,N_29925);
nand UO_1570 (O_1570,N_29889,N_29300);
and UO_1571 (O_1571,N_29448,N_29646);
xnor UO_1572 (O_1572,N_29439,N_29952);
and UO_1573 (O_1573,N_29068,N_29365);
and UO_1574 (O_1574,N_29409,N_29157);
or UO_1575 (O_1575,N_29664,N_29285);
nor UO_1576 (O_1576,N_29116,N_29940);
or UO_1577 (O_1577,N_29526,N_29917);
xnor UO_1578 (O_1578,N_29922,N_29486);
and UO_1579 (O_1579,N_29461,N_29626);
or UO_1580 (O_1580,N_29779,N_29187);
nand UO_1581 (O_1581,N_29596,N_29028);
nor UO_1582 (O_1582,N_29446,N_29284);
or UO_1583 (O_1583,N_29930,N_29521);
or UO_1584 (O_1584,N_29443,N_29811);
or UO_1585 (O_1585,N_29161,N_29983);
or UO_1586 (O_1586,N_29861,N_29104);
nand UO_1587 (O_1587,N_29386,N_29348);
xor UO_1588 (O_1588,N_29529,N_29297);
or UO_1589 (O_1589,N_29479,N_29359);
or UO_1590 (O_1590,N_29950,N_29440);
xor UO_1591 (O_1591,N_29755,N_29439);
nor UO_1592 (O_1592,N_29067,N_29296);
xnor UO_1593 (O_1593,N_29990,N_29413);
nor UO_1594 (O_1594,N_29228,N_29491);
and UO_1595 (O_1595,N_29188,N_29195);
xor UO_1596 (O_1596,N_29058,N_29442);
xor UO_1597 (O_1597,N_29896,N_29546);
or UO_1598 (O_1598,N_29588,N_29715);
and UO_1599 (O_1599,N_29244,N_29403);
nand UO_1600 (O_1600,N_29692,N_29978);
nor UO_1601 (O_1601,N_29946,N_29231);
nor UO_1602 (O_1602,N_29419,N_29317);
or UO_1603 (O_1603,N_29464,N_29663);
nor UO_1604 (O_1604,N_29280,N_29863);
nand UO_1605 (O_1605,N_29002,N_29689);
nand UO_1606 (O_1606,N_29285,N_29508);
xor UO_1607 (O_1607,N_29342,N_29230);
or UO_1608 (O_1608,N_29314,N_29482);
nand UO_1609 (O_1609,N_29947,N_29586);
and UO_1610 (O_1610,N_29664,N_29113);
and UO_1611 (O_1611,N_29490,N_29075);
nor UO_1612 (O_1612,N_29320,N_29028);
or UO_1613 (O_1613,N_29785,N_29338);
or UO_1614 (O_1614,N_29769,N_29911);
nor UO_1615 (O_1615,N_29749,N_29187);
xnor UO_1616 (O_1616,N_29006,N_29866);
nand UO_1617 (O_1617,N_29464,N_29021);
nand UO_1618 (O_1618,N_29566,N_29230);
nor UO_1619 (O_1619,N_29675,N_29454);
nor UO_1620 (O_1620,N_29626,N_29408);
nand UO_1621 (O_1621,N_29090,N_29284);
xor UO_1622 (O_1622,N_29302,N_29369);
and UO_1623 (O_1623,N_29174,N_29794);
xnor UO_1624 (O_1624,N_29022,N_29354);
and UO_1625 (O_1625,N_29122,N_29088);
and UO_1626 (O_1626,N_29941,N_29745);
and UO_1627 (O_1627,N_29783,N_29600);
xor UO_1628 (O_1628,N_29556,N_29440);
and UO_1629 (O_1629,N_29283,N_29397);
xnor UO_1630 (O_1630,N_29678,N_29322);
or UO_1631 (O_1631,N_29272,N_29020);
or UO_1632 (O_1632,N_29040,N_29639);
xor UO_1633 (O_1633,N_29867,N_29318);
or UO_1634 (O_1634,N_29613,N_29691);
nor UO_1635 (O_1635,N_29087,N_29383);
xnor UO_1636 (O_1636,N_29800,N_29266);
and UO_1637 (O_1637,N_29230,N_29456);
or UO_1638 (O_1638,N_29690,N_29208);
and UO_1639 (O_1639,N_29422,N_29749);
and UO_1640 (O_1640,N_29917,N_29554);
nor UO_1641 (O_1641,N_29344,N_29924);
nor UO_1642 (O_1642,N_29111,N_29865);
nor UO_1643 (O_1643,N_29266,N_29194);
or UO_1644 (O_1644,N_29318,N_29371);
xnor UO_1645 (O_1645,N_29731,N_29651);
nand UO_1646 (O_1646,N_29860,N_29571);
nor UO_1647 (O_1647,N_29776,N_29431);
nor UO_1648 (O_1648,N_29802,N_29413);
xor UO_1649 (O_1649,N_29216,N_29368);
nand UO_1650 (O_1650,N_29686,N_29672);
or UO_1651 (O_1651,N_29494,N_29578);
and UO_1652 (O_1652,N_29790,N_29175);
xnor UO_1653 (O_1653,N_29232,N_29018);
xnor UO_1654 (O_1654,N_29510,N_29630);
nor UO_1655 (O_1655,N_29017,N_29485);
nor UO_1656 (O_1656,N_29976,N_29790);
nand UO_1657 (O_1657,N_29892,N_29787);
nor UO_1658 (O_1658,N_29910,N_29017);
xor UO_1659 (O_1659,N_29101,N_29450);
or UO_1660 (O_1660,N_29299,N_29562);
nor UO_1661 (O_1661,N_29482,N_29795);
nor UO_1662 (O_1662,N_29620,N_29369);
nor UO_1663 (O_1663,N_29170,N_29221);
xor UO_1664 (O_1664,N_29935,N_29825);
or UO_1665 (O_1665,N_29609,N_29561);
xor UO_1666 (O_1666,N_29664,N_29879);
xor UO_1667 (O_1667,N_29974,N_29964);
nand UO_1668 (O_1668,N_29012,N_29422);
or UO_1669 (O_1669,N_29130,N_29269);
or UO_1670 (O_1670,N_29062,N_29078);
nand UO_1671 (O_1671,N_29101,N_29074);
or UO_1672 (O_1672,N_29713,N_29295);
or UO_1673 (O_1673,N_29928,N_29273);
and UO_1674 (O_1674,N_29892,N_29599);
or UO_1675 (O_1675,N_29037,N_29723);
nor UO_1676 (O_1676,N_29081,N_29924);
nor UO_1677 (O_1677,N_29708,N_29425);
nand UO_1678 (O_1678,N_29233,N_29178);
nor UO_1679 (O_1679,N_29234,N_29366);
nor UO_1680 (O_1680,N_29620,N_29904);
or UO_1681 (O_1681,N_29946,N_29860);
or UO_1682 (O_1682,N_29700,N_29332);
xor UO_1683 (O_1683,N_29618,N_29115);
nor UO_1684 (O_1684,N_29333,N_29467);
and UO_1685 (O_1685,N_29481,N_29609);
nor UO_1686 (O_1686,N_29379,N_29011);
or UO_1687 (O_1687,N_29854,N_29464);
nand UO_1688 (O_1688,N_29659,N_29535);
xnor UO_1689 (O_1689,N_29326,N_29237);
nand UO_1690 (O_1690,N_29914,N_29785);
and UO_1691 (O_1691,N_29600,N_29865);
or UO_1692 (O_1692,N_29393,N_29210);
or UO_1693 (O_1693,N_29640,N_29178);
or UO_1694 (O_1694,N_29424,N_29661);
nand UO_1695 (O_1695,N_29938,N_29912);
nand UO_1696 (O_1696,N_29120,N_29844);
nor UO_1697 (O_1697,N_29489,N_29971);
nand UO_1698 (O_1698,N_29406,N_29522);
nand UO_1699 (O_1699,N_29262,N_29512);
nor UO_1700 (O_1700,N_29903,N_29004);
or UO_1701 (O_1701,N_29416,N_29575);
nand UO_1702 (O_1702,N_29403,N_29646);
nand UO_1703 (O_1703,N_29670,N_29325);
and UO_1704 (O_1704,N_29201,N_29415);
and UO_1705 (O_1705,N_29019,N_29800);
nor UO_1706 (O_1706,N_29967,N_29407);
nand UO_1707 (O_1707,N_29759,N_29074);
or UO_1708 (O_1708,N_29770,N_29784);
or UO_1709 (O_1709,N_29642,N_29237);
nand UO_1710 (O_1710,N_29354,N_29905);
nor UO_1711 (O_1711,N_29763,N_29855);
and UO_1712 (O_1712,N_29948,N_29661);
nand UO_1713 (O_1713,N_29478,N_29552);
and UO_1714 (O_1714,N_29348,N_29411);
xor UO_1715 (O_1715,N_29454,N_29768);
nand UO_1716 (O_1716,N_29115,N_29720);
nor UO_1717 (O_1717,N_29760,N_29147);
and UO_1718 (O_1718,N_29573,N_29011);
nand UO_1719 (O_1719,N_29851,N_29045);
xnor UO_1720 (O_1720,N_29934,N_29605);
or UO_1721 (O_1721,N_29953,N_29252);
nor UO_1722 (O_1722,N_29160,N_29385);
xnor UO_1723 (O_1723,N_29960,N_29159);
and UO_1724 (O_1724,N_29038,N_29692);
and UO_1725 (O_1725,N_29296,N_29665);
or UO_1726 (O_1726,N_29860,N_29274);
nand UO_1727 (O_1727,N_29024,N_29311);
or UO_1728 (O_1728,N_29813,N_29780);
xnor UO_1729 (O_1729,N_29541,N_29549);
or UO_1730 (O_1730,N_29111,N_29883);
xor UO_1731 (O_1731,N_29540,N_29947);
nand UO_1732 (O_1732,N_29579,N_29521);
nor UO_1733 (O_1733,N_29269,N_29180);
nand UO_1734 (O_1734,N_29219,N_29068);
and UO_1735 (O_1735,N_29325,N_29005);
xor UO_1736 (O_1736,N_29404,N_29590);
nand UO_1737 (O_1737,N_29446,N_29022);
or UO_1738 (O_1738,N_29914,N_29705);
nor UO_1739 (O_1739,N_29501,N_29965);
nor UO_1740 (O_1740,N_29044,N_29453);
and UO_1741 (O_1741,N_29116,N_29455);
nand UO_1742 (O_1742,N_29562,N_29390);
xnor UO_1743 (O_1743,N_29381,N_29977);
and UO_1744 (O_1744,N_29723,N_29902);
nand UO_1745 (O_1745,N_29293,N_29334);
and UO_1746 (O_1746,N_29754,N_29940);
xor UO_1747 (O_1747,N_29139,N_29613);
nor UO_1748 (O_1748,N_29739,N_29820);
nor UO_1749 (O_1749,N_29722,N_29725);
and UO_1750 (O_1750,N_29711,N_29353);
or UO_1751 (O_1751,N_29434,N_29111);
or UO_1752 (O_1752,N_29572,N_29605);
nand UO_1753 (O_1753,N_29970,N_29264);
nand UO_1754 (O_1754,N_29861,N_29887);
xor UO_1755 (O_1755,N_29124,N_29623);
or UO_1756 (O_1756,N_29886,N_29108);
or UO_1757 (O_1757,N_29098,N_29152);
and UO_1758 (O_1758,N_29305,N_29490);
nand UO_1759 (O_1759,N_29951,N_29124);
or UO_1760 (O_1760,N_29537,N_29449);
nand UO_1761 (O_1761,N_29796,N_29226);
nand UO_1762 (O_1762,N_29650,N_29499);
nand UO_1763 (O_1763,N_29913,N_29599);
and UO_1764 (O_1764,N_29854,N_29899);
or UO_1765 (O_1765,N_29573,N_29544);
and UO_1766 (O_1766,N_29834,N_29901);
nand UO_1767 (O_1767,N_29011,N_29457);
xor UO_1768 (O_1768,N_29087,N_29155);
or UO_1769 (O_1769,N_29091,N_29367);
nand UO_1770 (O_1770,N_29417,N_29136);
xnor UO_1771 (O_1771,N_29839,N_29980);
and UO_1772 (O_1772,N_29330,N_29747);
and UO_1773 (O_1773,N_29679,N_29080);
nor UO_1774 (O_1774,N_29047,N_29751);
nand UO_1775 (O_1775,N_29975,N_29787);
or UO_1776 (O_1776,N_29534,N_29897);
or UO_1777 (O_1777,N_29714,N_29353);
xor UO_1778 (O_1778,N_29335,N_29641);
or UO_1779 (O_1779,N_29883,N_29362);
xor UO_1780 (O_1780,N_29692,N_29135);
or UO_1781 (O_1781,N_29857,N_29623);
nor UO_1782 (O_1782,N_29241,N_29364);
and UO_1783 (O_1783,N_29232,N_29317);
and UO_1784 (O_1784,N_29230,N_29376);
or UO_1785 (O_1785,N_29678,N_29460);
xnor UO_1786 (O_1786,N_29034,N_29516);
nand UO_1787 (O_1787,N_29994,N_29323);
nand UO_1788 (O_1788,N_29606,N_29103);
nand UO_1789 (O_1789,N_29738,N_29509);
xor UO_1790 (O_1790,N_29969,N_29959);
and UO_1791 (O_1791,N_29057,N_29386);
nor UO_1792 (O_1792,N_29780,N_29298);
or UO_1793 (O_1793,N_29637,N_29610);
nand UO_1794 (O_1794,N_29778,N_29832);
and UO_1795 (O_1795,N_29195,N_29411);
xor UO_1796 (O_1796,N_29411,N_29010);
nor UO_1797 (O_1797,N_29758,N_29941);
xnor UO_1798 (O_1798,N_29218,N_29152);
nor UO_1799 (O_1799,N_29164,N_29705);
nand UO_1800 (O_1800,N_29531,N_29216);
or UO_1801 (O_1801,N_29914,N_29726);
and UO_1802 (O_1802,N_29402,N_29796);
xnor UO_1803 (O_1803,N_29384,N_29682);
nand UO_1804 (O_1804,N_29241,N_29439);
xnor UO_1805 (O_1805,N_29840,N_29561);
or UO_1806 (O_1806,N_29330,N_29439);
nand UO_1807 (O_1807,N_29775,N_29415);
or UO_1808 (O_1808,N_29959,N_29887);
nand UO_1809 (O_1809,N_29090,N_29064);
and UO_1810 (O_1810,N_29234,N_29553);
or UO_1811 (O_1811,N_29494,N_29513);
nor UO_1812 (O_1812,N_29797,N_29171);
or UO_1813 (O_1813,N_29621,N_29002);
nand UO_1814 (O_1814,N_29463,N_29743);
xnor UO_1815 (O_1815,N_29669,N_29416);
nor UO_1816 (O_1816,N_29707,N_29642);
xnor UO_1817 (O_1817,N_29814,N_29897);
nor UO_1818 (O_1818,N_29050,N_29427);
nand UO_1819 (O_1819,N_29114,N_29142);
nand UO_1820 (O_1820,N_29253,N_29881);
nand UO_1821 (O_1821,N_29355,N_29581);
and UO_1822 (O_1822,N_29190,N_29805);
and UO_1823 (O_1823,N_29526,N_29996);
nand UO_1824 (O_1824,N_29853,N_29725);
xor UO_1825 (O_1825,N_29702,N_29283);
xor UO_1826 (O_1826,N_29868,N_29588);
xnor UO_1827 (O_1827,N_29989,N_29746);
xor UO_1828 (O_1828,N_29741,N_29332);
xor UO_1829 (O_1829,N_29027,N_29490);
xor UO_1830 (O_1830,N_29455,N_29495);
xnor UO_1831 (O_1831,N_29736,N_29907);
and UO_1832 (O_1832,N_29694,N_29023);
and UO_1833 (O_1833,N_29182,N_29737);
nand UO_1834 (O_1834,N_29532,N_29102);
nor UO_1835 (O_1835,N_29400,N_29283);
nand UO_1836 (O_1836,N_29838,N_29053);
or UO_1837 (O_1837,N_29119,N_29273);
nand UO_1838 (O_1838,N_29237,N_29535);
nand UO_1839 (O_1839,N_29043,N_29452);
nor UO_1840 (O_1840,N_29328,N_29292);
or UO_1841 (O_1841,N_29778,N_29620);
nor UO_1842 (O_1842,N_29539,N_29439);
nand UO_1843 (O_1843,N_29606,N_29985);
or UO_1844 (O_1844,N_29119,N_29395);
and UO_1845 (O_1845,N_29171,N_29376);
xnor UO_1846 (O_1846,N_29668,N_29058);
xnor UO_1847 (O_1847,N_29539,N_29221);
nor UO_1848 (O_1848,N_29154,N_29251);
or UO_1849 (O_1849,N_29147,N_29751);
xnor UO_1850 (O_1850,N_29090,N_29524);
nor UO_1851 (O_1851,N_29125,N_29229);
xnor UO_1852 (O_1852,N_29271,N_29875);
or UO_1853 (O_1853,N_29732,N_29943);
and UO_1854 (O_1854,N_29304,N_29713);
or UO_1855 (O_1855,N_29499,N_29665);
nand UO_1856 (O_1856,N_29835,N_29659);
or UO_1857 (O_1857,N_29792,N_29202);
xor UO_1858 (O_1858,N_29818,N_29498);
and UO_1859 (O_1859,N_29876,N_29448);
or UO_1860 (O_1860,N_29545,N_29178);
nor UO_1861 (O_1861,N_29967,N_29528);
nor UO_1862 (O_1862,N_29171,N_29853);
xnor UO_1863 (O_1863,N_29621,N_29664);
nor UO_1864 (O_1864,N_29319,N_29291);
or UO_1865 (O_1865,N_29661,N_29611);
and UO_1866 (O_1866,N_29522,N_29683);
nor UO_1867 (O_1867,N_29772,N_29729);
nor UO_1868 (O_1868,N_29612,N_29405);
nor UO_1869 (O_1869,N_29040,N_29231);
xor UO_1870 (O_1870,N_29567,N_29651);
nor UO_1871 (O_1871,N_29131,N_29819);
or UO_1872 (O_1872,N_29772,N_29553);
or UO_1873 (O_1873,N_29739,N_29550);
xnor UO_1874 (O_1874,N_29074,N_29321);
nand UO_1875 (O_1875,N_29565,N_29479);
or UO_1876 (O_1876,N_29825,N_29679);
and UO_1877 (O_1877,N_29456,N_29796);
nor UO_1878 (O_1878,N_29280,N_29559);
nand UO_1879 (O_1879,N_29352,N_29399);
xnor UO_1880 (O_1880,N_29567,N_29450);
nand UO_1881 (O_1881,N_29725,N_29894);
nand UO_1882 (O_1882,N_29420,N_29857);
xor UO_1883 (O_1883,N_29115,N_29404);
and UO_1884 (O_1884,N_29099,N_29511);
nor UO_1885 (O_1885,N_29675,N_29223);
or UO_1886 (O_1886,N_29222,N_29438);
and UO_1887 (O_1887,N_29216,N_29572);
nand UO_1888 (O_1888,N_29904,N_29417);
or UO_1889 (O_1889,N_29630,N_29053);
or UO_1890 (O_1890,N_29608,N_29885);
or UO_1891 (O_1891,N_29233,N_29287);
xor UO_1892 (O_1892,N_29089,N_29804);
and UO_1893 (O_1893,N_29425,N_29546);
xor UO_1894 (O_1894,N_29874,N_29986);
nor UO_1895 (O_1895,N_29931,N_29567);
nor UO_1896 (O_1896,N_29881,N_29585);
or UO_1897 (O_1897,N_29704,N_29247);
and UO_1898 (O_1898,N_29915,N_29189);
nor UO_1899 (O_1899,N_29898,N_29815);
or UO_1900 (O_1900,N_29651,N_29576);
xnor UO_1901 (O_1901,N_29361,N_29267);
or UO_1902 (O_1902,N_29057,N_29148);
and UO_1903 (O_1903,N_29255,N_29306);
or UO_1904 (O_1904,N_29529,N_29444);
nor UO_1905 (O_1905,N_29251,N_29027);
xor UO_1906 (O_1906,N_29585,N_29174);
nor UO_1907 (O_1907,N_29770,N_29334);
and UO_1908 (O_1908,N_29776,N_29012);
or UO_1909 (O_1909,N_29005,N_29951);
nand UO_1910 (O_1910,N_29960,N_29525);
nand UO_1911 (O_1911,N_29881,N_29902);
and UO_1912 (O_1912,N_29912,N_29146);
and UO_1913 (O_1913,N_29050,N_29829);
nor UO_1914 (O_1914,N_29079,N_29380);
and UO_1915 (O_1915,N_29482,N_29547);
and UO_1916 (O_1916,N_29676,N_29574);
nor UO_1917 (O_1917,N_29194,N_29972);
or UO_1918 (O_1918,N_29563,N_29163);
nand UO_1919 (O_1919,N_29373,N_29639);
nand UO_1920 (O_1920,N_29053,N_29766);
nand UO_1921 (O_1921,N_29375,N_29545);
nor UO_1922 (O_1922,N_29608,N_29033);
and UO_1923 (O_1923,N_29453,N_29238);
nor UO_1924 (O_1924,N_29461,N_29892);
nand UO_1925 (O_1925,N_29262,N_29746);
xnor UO_1926 (O_1926,N_29814,N_29464);
nor UO_1927 (O_1927,N_29795,N_29667);
xnor UO_1928 (O_1928,N_29712,N_29746);
nand UO_1929 (O_1929,N_29464,N_29268);
nor UO_1930 (O_1930,N_29162,N_29569);
nor UO_1931 (O_1931,N_29992,N_29139);
nor UO_1932 (O_1932,N_29184,N_29334);
nor UO_1933 (O_1933,N_29498,N_29812);
and UO_1934 (O_1934,N_29205,N_29142);
nor UO_1935 (O_1935,N_29372,N_29173);
and UO_1936 (O_1936,N_29848,N_29380);
or UO_1937 (O_1937,N_29285,N_29609);
nor UO_1938 (O_1938,N_29806,N_29670);
xnor UO_1939 (O_1939,N_29077,N_29218);
nor UO_1940 (O_1940,N_29833,N_29462);
or UO_1941 (O_1941,N_29094,N_29732);
nor UO_1942 (O_1942,N_29968,N_29109);
and UO_1943 (O_1943,N_29193,N_29683);
xor UO_1944 (O_1944,N_29615,N_29652);
and UO_1945 (O_1945,N_29030,N_29810);
or UO_1946 (O_1946,N_29261,N_29403);
and UO_1947 (O_1947,N_29026,N_29634);
and UO_1948 (O_1948,N_29005,N_29077);
nand UO_1949 (O_1949,N_29682,N_29147);
or UO_1950 (O_1950,N_29026,N_29929);
nor UO_1951 (O_1951,N_29939,N_29782);
or UO_1952 (O_1952,N_29825,N_29939);
and UO_1953 (O_1953,N_29601,N_29565);
nand UO_1954 (O_1954,N_29360,N_29940);
nand UO_1955 (O_1955,N_29608,N_29122);
nand UO_1956 (O_1956,N_29969,N_29784);
xnor UO_1957 (O_1957,N_29000,N_29449);
and UO_1958 (O_1958,N_29369,N_29547);
and UO_1959 (O_1959,N_29308,N_29630);
or UO_1960 (O_1960,N_29607,N_29104);
nand UO_1961 (O_1961,N_29378,N_29132);
or UO_1962 (O_1962,N_29606,N_29081);
and UO_1963 (O_1963,N_29350,N_29102);
nor UO_1964 (O_1964,N_29046,N_29777);
xor UO_1965 (O_1965,N_29875,N_29369);
or UO_1966 (O_1966,N_29813,N_29606);
nand UO_1967 (O_1967,N_29123,N_29872);
nor UO_1968 (O_1968,N_29059,N_29103);
xor UO_1969 (O_1969,N_29534,N_29673);
and UO_1970 (O_1970,N_29337,N_29166);
and UO_1971 (O_1971,N_29055,N_29086);
nor UO_1972 (O_1972,N_29424,N_29677);
nand UO_1973 (O_1973,N_29789,N_29295);
and UO_1974 (O_1974,N_29686,N_29157);
nor UO_1975 (O_1975,N_29744,N_29867);
xnor UO_1976 (O_1976,N_29241,N_29863);
nand UO_1977 (O_1977,N_29364,N_29797);
or UO_1978 (O_1978,N_29549,N_29029);
nor UO_1979 (O_1979,N_29579,N_29544);
and UO_1980 (O_1980,N_29610,N_29407);
and UO_1981 (O_1981,N_29247,N_29655);
nand UO_1982 (O_1982,N_29090,N_29175);
and UO_1983 (O_1983,N_29824,N_29989);
and UO_1984 (O_1984,N_29197,N_29384);
nand UO_1985 (O_1985,N_29468,N_29136);
xnor UO_1986 (O_1986,N_29219,N_29670);
nand UO_1987 (O_1987,N_29910,N_29136);
and UO_1988 (O_1988,N_29245,N_29081);
and UO_1989 (O_1989,N_29778,N_29845);
or UO_1990 (O_1990,N_29803,N_29568);
nand UO_1991 (O_1991,N_29003,N_29802);
nor UO_1992 (O_1992,N_29963,N_29420);
nor UO_1993 (O_1993,N_29539,N_29581);
nand UO_1994 (O_1994,N_29579,N_29949);
or UO_1995 (O_1995,N_29192,N_29970);
and UO_1996 (O_1996,N_29376,N_29725);
or UO_1997 (O_1997,N_29585,N_29268);
nand UO_1998 (O_1998,N_29454,N_29967);
nand UO_1999 (O_1999,N_29254,N_29910);
xnor UO_2000 (O_2000,N_29966,N_29433);
or UO_2001 (O_2001,N_29109,N_29684);
and UO_2002 (O_2002,N_29846,N_29720);
nand UO_2003 (O_2003,N_29848,N_29251);
nor UO_2004 (O_2004,N_29363,N_29188);
and UO_2005 (O_2005,N_29676,N_29049);
and UO_2006 (O_2006,N_29667,N_29948);
or UO_2007 (O_2007,N_29146,N_29692);
xnor UO_2008 (O_2008,N_29327,N_29446);
and UO_2009 (O_2009,N_29851,N_29316);
nor UO_2010 (O_2010,N_29107,N_29855);
and UO_2011 (O_2011,N_29791,N_29973);
xnor UO_2012 (O_2012,N_29259,N_29896);
or UO_2013 (O_2013,N_29238,N_29120);
xor UO_2014 (O_2014,N_29417,N_29075);
nor UO_2015 (O_2015,N_29135,N_29417);
nand UO_2016 (O_2016,N_29974,N_29463);
xnor UO_2017 (O_2017,N_29949,N_29090);
nand UO_2018 (O_2018,N_29475,N_29541);
nor UO_2019 (O_2019,N_29151,N_29684);
and UO_2020 (O_2020,N_29560,N_29311);
xnor UO_2021 (O_2021,N_29822,N_29736);
nand UO_2022 (O_2022,N_29423,N_29583);
xnor UO_2023 (O_2023,N_29463,N_29796);
and UO_2024 (O_2024,N_29181,N_29608);
nand UO_2025 (O_2025,N_29595,N_29007);
nor UO_2026 (O_2026,N_29162,N_29206);
or UO_2027 (O_2027,N_29869,N_29606);
xor UO_2028 (O_2028,N_29864,N_29558);
and UO_2029 (O_2029,N_29745,N_29162);
nand UO_2030 (O_2030,N_29899,N_29588);
xor UO_2031 (O_2031,N_29724,N_29185);
nand UO_2032 (O_2032,N_29019,N_29099);
and UO_2033 (O_2033,N_29998,N_29370);
and UO_2034 (O_2034,N_29498,N_29069);
nand UO_2035 (O_2035,N_29484,N_29151);
xnor UO_2036 (O_2036,N_29779,N_29396);
nor UO_2037 (O_2037,N_29581,N_29432);
or UO_2038 (O_2038,N_29385,N_29525);
nor UO_2039 (O_2039,N_29905,N_29355);
nand UO_2040 (O_2040,N_29296,N_29045);
nand UO_2041 (O_2041,N_29360,N_29412);
or UO_2042 (O_2042,N_29239,N_29720);
and UO_2043 (O_2043,N_29579,N_29608);
nor UO_2044 (O_2044,N_29116,N_29247);
or UO_2045 (O_2045,N_29861,N_29206);
nor UO_2046 (O_2046,N_29879,N_29232);
nor UO_2047 (O_2047,N_29294,N_29249);
and UO_2048 (O_2048,N_29334,N_29795);
xnor UO_2049 (O_2049,N_29880,N_29644);
or UO_2050 (O_2050,N_29423,N_29558);
nand UO_2051 (O_2051,N_29228,N_29310);
nor UO_2052 (O_2052,N_29698,N_29432);
or UO_2053 (O_2053,N_29351,N_29067);
xor UO_2054 (O_2054,N_29769,N_29134);
and UO_2055 (O_2055,N_29020,N_29400);
nand UO_2056 (O_2056,N_29899,N_29036);
nor UO_2057 (O_2057,N_29411,N_29681);
and UO_2058 (O_2058,N_29519,N_29134);
nor UO_2059 (O_2059,N_29589,N_29532);
and UO_2060 (O_2060,N_29615,N_29372);
nand UO_2061 (O_2061,N_29326,N_29288);
or UO_2062 (O_2062,N_29710,N_29377);
nor UO_2063 (O_2063,N_29226,N_29695);
and UO_2064 (O_2064,N_29775,N_29472);
xor UO_2065 (O_2065,N_29108,N_29266);
or UO_2066 (O_2066,N_29972,N_29636);
and UO_2067 (O_2067,N_29695,N_29241);
nor UO_2068 (O_2068,N_29381,N_29442);
nand UO_2069 (O_2069,N_29480,N_29854);
xnor UO_2070 (O_2070,N_29035,N_29993);
xor UO_2071 (O_2071,N_29840,N_29603);
nor UO_2072 (O_2072,N_29551,N_29420);
nand UO_2073 (O_2073,N_29784,N_29968);
and UO_2074 (O_2074,N_29610,N_29224);
nand UO_2075 (O_2075,N_29408,N_29540);
nor UO_2076 (O_2076,N_29792,N_29051);
nand UO_2077 (O_2077,N_29616,N_29029);
nor UO_2078 (O_2078,N_29910,N_29499);
and UO_2079 (O_2079,N_29814,N_29259);
and UO_2080 (O_2080,N_29146,N_29515);
or UO_2081 (O_2081,N_29887,N_29910);
nand UO_2082 (O_2082,N_29939,N_29745);
xor UO_2083 (O_2083,N_29289,N_29562);
xnor UO_2084 (O_2084,N_29824,N_29961);
nand UO_2085 (O_2085,N_29876,N_29243);
xnor UO_2086 (O_2086,N_29391,N_29956);
or UO_2087 (O_2087,N_29977,N_29827);
nor UO_2088 (O_2088,N_29279,N_29263);
nand UO_2089 (O_2089,N_29595,N_29606);
nor UO_2090 (O_2090,N_29792,N_29611);
and UO_2091 (O_2091,N_29951,N_29663);
or UO_2092 (O_2092,N_29855,N_29553);
nor UO_2093 (O_2093,N_29536,N_29346);
nor UO_2094 (O_2094,N_29743,N_29629);
nand UO_2095 (O_2095,N_29846,N_29946);
nor UO_2096 (O_2096,N_29181,N_29950);
nor UO_2097 (O_2097,N_29382,N_29439);
or UO_2098 (O_2098,N_29354,N_29275);
nor UO_2099 (O_2099,N_29239,N_29715);
and UO_2100 (O_2100,N_29066,N_29167);
nor UO_2101 (O_2101,N_29088,N_29688);
nand UO_2102 (O_2102,N_29575,N_29342);
nor UO_2103 (O_2103,N_29970,N_29181);
xor UO_2104 (O_2104,N_29598,N_29251);
nand UO_2105 (O_2105,N_29944,N_29046);
or UO_2106 (O_2106,N_29470,N_29474);
xor UO_2107 (O_2107,N_29539,N_29010);
or UO_2108 (O_2108,N_29215,N_29980);
nand UO_2109 (O_2109,N_29923,N_29893);
or UO_2110 (O_2110,N_29932,N_29151);
nand UO_2111 (O_2111,N_29188,N_29889);
xor UO_2112 (O_2112,N_29546,N_29348);
xor UO_2113 (O_2113,N_29742,N_29296);
and UO_2114 (O_2114,N_29095,N_29379);
nor UO_2115 (O_2115,N_29971,N_29973);
nand UO_2116 (O_2116,N_29021,N_29416);
nand UO_2117 (O_2117,N_29884,N_29609);
or UO_2118 (O_2118,N_29609,N_29866);
or UO_2119 (O_2119,N_29290,N_29736);
or UO_2120 (O_2120,N_29020,N_29177);
nand UO_2121 (O_2121,N_29668,N_29106);
xor UO_2122 (O_2122,N_29962,N_29805);
nor UO_2123 (O_2123,N_29540,N_29475);
nor UO_2124 (O_2124,N_29553,N_29376);
nor UO_2125 (O_2125,N_29119,N_29156);
nand UO_2126 (O_2126,N_29451,N_29495);
nand UO_2127 (O_2127,N_29989,N_29568);
nor UO_2128 (O_2128,N_29410,N_29036);
and UO_2129 (O_2129,N_29993,N_29833);
xnor UO_2130 (O_2130,N_29187,N_29560);
or UO_2131 (O_2131,N_29104,N_29395);
and UO_2132 (O_2132,N_29715,N_29689);
nor UO_2133 (O_2133,N_29081,N_29022);
xnor UO_2134 (O_2134,N_29694,N_29905);
nand UO_2135 (O_2135,N_29955,N_29856);
nor UO_2136 (O_2136,N_29022,N_29758);
nor UO_2137 (O_2137,N_29021,N_29580);
xnor UO_2138 (O_2138,N_29695,N_29605);
or UO_2139 (O_2139,N_29685,N_29996);
xor UO_2140 (O_2140,N_29157,N_29895);
nor UO_2141 (O_2141,N_29781,N_29908);
and UO_2142 (O_2142,N_29228,N_29005);
xnor UO_2143 (O_2143,N_29958,N_29980);
nand UO_2144 (O_2144,N_29593,N_29383);
nor UO_2145 (O_2145,N_29031,N_29807);
and UO_2146 (O_2146,N_29391,N_29698);
nand UO_2147 (O_2147,N_29608,N_29074);
or UO_2148 (O_2148,N_29771,N_29170);
nand UO_2149 (O_2149,N_29463,N_29277);
or UO_2150 (O_2150,N_29407,N_29894);
nor UO_2151 (O_2151,N_29711,N_29046);
xnor UO_2152 (O_2152,N_29332,N_29545);
and UO_2153 (O_2153,N_29535,N_29723);
xor UO_2154 (O_2154,N_29418,N_29728);
xnor UO_2155 (O_2155,N_29369,N_29674);
or UO_2156 (O_2156,N_29651,N_29983);
or UO_2157 (O_2157,N_29754,N_29012);
nand UO_2158 (O_2158,N_29455,N_29013);
xor UO_2159 (O_2159,N_29907,N_29710);
xor UO_2160 (O_2160,N_29525,N_29576);
xor UO_2161 (O_2161,N_29185,N_29759);
or UO_2162 (O_2162,N_29249,N_29373);
nor UO_2163 (O_2163,N_29555,N_29710);
xnor UO_2164 (O_2164,N_29548,N_29308);
xor UO_2165 (O_2165,N_29994,N_29148);
xnor UO_2166 (O_2166,N_29092,N_29883);
nor UO_2167 (O_2167,N_29808,N_29943);
xor UO_2168 (O_2168,N_29986,N_29377);
xnor UO_2169 (O_2169,N_29214,N_29209);
or UO_2170 (O_2170,N_29353,N_29806);
or UO_2171 (O_2171,N_29893,N_29672);
nand UO_2172 (O_2172,N_29617,N_29719);
and UO_2173 (O_2173,N_29992,N_29445);
and UO_2174 (O_2174,N_29365,N_29073);
or UO_2175 (O_2175,N_29600,N_29951);
xor UO_2176 (O_2176,N_29875,N_29108);
nor UO_2177 (O_2177,N_29887,N_29182);
xor UO_2178 (O_2178,N_29744,N_29129);
or UO_2179 (O_2179,N_29436,N_29742);
or UO_2180 (O_2180,N_29246,N_29766);
nand UO_2181 (O_2181,N_29030,N_29651);
xnor UO_2182 (O_2182,N_29082,N_29712);
nand UO_2183 (O_2183,N_29783,N_29136);
nand UO_2184 (O_2184,N_29005,N_29449);
nor UO_2185 (O_2185,N_29560,N_29944);
or UO_2186 (O_2186,N_29586,N_29416);
nand UO_2187 (O_2187,N_29221,N_29040);
nand UO_2188 (O_2188,N_29829,N_29652);
xor UO_2189 (O_2189,N_29750,N_29425);
and UO_2190 (O_2190,N_29269,N_29683);
nor UO_2191 (O_2191,N_29211,N_29815);
xnor UO_2192 (O_2192,N_29764,N_29311);
or UO_2193 (O_2193,N_29654,N_29862);
nor UO_2194 (O_2194,N_29358,N_29172);
xnor UO_2195 (O_2195,N_29300,N_29051);
nand UO_2196 (O_2196,N_29711,N_29279);
nor UO_2197 (O_2197,N_29122,N_29923);
nor UO_2198 (O_2198,N_29450,N_29737);
xor UO_2199 (O_2199,N_29656,N_29465);
or UO_2200 (O_2200,N_29606,N_29046);
nand UO_2201 (O_2201,N_29373,N_29944);
xnor UO_2202 (O_2202,N_29497,N_29139);
and UO_2203 (O_2203,N_29235,N_29467);
nand UO_2204 (O_2204,N_29302,N_29052);
and UO_2205 (O_2205,N_29250,N_29087);
xnor UO_2206 (O_2206,N_29234,N_29104);
xnor UO_2207 (O_2207,N_29640,N_29324);
or UO_2208 (O_2208,N_29943,N_29950);
or UO_2209 (O_2209,N_29114,N_29291);
xor UO_2210 (O_2210,N_29697,N_29601);
nand UO_2211 (O_2211,N_29328,N_29271);
nor UO_2212 (O_2212,N_29232,N_29376);
or UO_2213 (O_2213,N_29111,N_29047);
nor UO_2214 (O_2214,N_29369,N_29357);
nand UO_2215 (O_2215,N_29908,N_29162);
or UO_2216 (O_2216,N_29919,N_29714);
xor UO_2217 (O_2217,N_29231,N_29488);
or UO_2218 (O_2218,N_29472,N_29799);
xor UO_2219 (O_2219,N_29660,N_29937);
nand UO_2220 (O_2220,N_29333,N_29953);
nor UO_2221 (O_2221,N_29250,N_29711);
xor UO_2222 (O_2222,N_29593,N_29497);
and UO_2223 (O_2223,N_29225,N_29841);
or UO_2224 (O_2224,N_29696,N_29443);
xor UO_2225 (O_2225,N_29884,N_29978);
or UO_2226 (O_2226,N_29466,N_29167);
and UO_2227 (O_2227,N_29918,N_29916);
nor UO_2228 (O_2228,N_29909,N_29139);
nor UO_2229 (O_2229,N_29998,N_29038);
nand UO_2230 (O_2230,N_29010,N_29061);
nor UO_2231 (O_2231,N_29466,N_29463);
nand UO_2232 (O_2232,N_29376,N_29395);
nand UO_2233 (O_2233,N_29430,N_29681);
or UO_2234 (O_2234,N_29177,N_29490);
or UO_2235 (O_2235,N_29205,N_29241);
or UO_2236 (O_2236,N_29728,N_29475);
and UO_2237 (O_2237,N_29050,N_29854);
and UO_2238 (O_2238,N_29562,N_29732);
and UO_2239 (O_2239,N_29648,N_29103);
nand UO_2240 (O_2240,N_29352,N_29827);
nand UO_2241 (O_2241,N_29475,N_29079);
xor UO_2242 (O_2242,N_29772,N_29838);
nor UO_2243 (O_2243,N_29794,N_29691);
xor UO_2244 (O_2244,N_29973,N_29599);
and UO_2245 (O_2245,N_29424,N_29317);
and UO_2246 (O_2246,N_29054,N_29080);
xnor UO_2247 (O_2247,N_29475,N_29675);
xor UO_2248 (O_2248,N_29021,N_29492);
nor UO_2249 (O_2249,N_29304,N_29318);
nand UO_2250 (O_2250,N_29578,N_29853);
nor UO_2251 (O_2251,N_29313,N_29992);
xnor UO_2252 (O_2252,N_29324,N_29442);
or UO_2253 (O_2253,N_29995,N_29836);
nand UO_2254 (O_2254,N_29158,N_29659);
and UO_2255 (O_2255,N_29902,N_29005);
or UO_2256 (O_2256,N_29990,N_29739);
and UO_2257 (O_2257,N_29315,N_29764);
and UO_2258 (O_2258,N_29453,N_29325);
nand UO_2259 (O_2259,N_29592,N_29042);
xor UO_2260 (O_2260,N_29578,N_29872);
xor UO_2261 (O_2261,N_29321,N_29033);
xnor UO_2262 (O_2262,N_29719,N_29192);
or UO_2263 (O_2263,N_29077,N_29951);
nand UO_2264 (O_2264,N_29044,N_29167);
or UO_2265 (O_2265,N_29603,N_29256);
xor UO_2266 (O_2266,N_29940,N_29211);
or UO_2267 (O_2267,N_29315,N_29686);
and UO_2268 (O_2268,N_29376,N_29539);
xnor UO_2269 (O_2269,N_29005,N_29267);
nor UO_2270 (O_2270,N_29133,N_29652);
and UO_2271 (O_2271,N_29146,N_29796);
xor UO_2272 (O_2272,N_29131,N_29279);
and UO_2273 (O_2273,N_29468,N_29292);
nand UO_2274 (O_2274,N_29287,N_29481);
nand UO_2275 (O_2275,N_29478,N_29696);
nor UO_2276 (O_2276,N_29644,N_29114);
xnor UO_2277 (O_2277,N_29813,N_29343);
nand UO_2278 (O_2278,N_29236,N_29508);
nand UO_2279 (O_2279,N_29604,N_29587);
and UO_2280 (O_2280,N_29824,N_29808);
or UO_2281 (O_2281,N_29796,N_29268);
nor UO_2282 (O_2282,N_29358,N_29221);
and UO_2283 (O_2283,N_29887,N_29519);
xnor UO_2284 (O_2284,N_29072,N_29515);
nor UO_2285 (O_2285,N_29638,N_29517);
nand UO_2286 (O_2286,N_29345,N_29411);
or UO_2287 (O_2287,N_29365,N_29926);
nand UO_2288 (O_2288,N_29276,N_29184);
or UO_2289 (O_2289,N_29134,N_29386);
xnor UO_2290 (O_2290,N_29601,N_29520);
or UO_2291 (O_2291,N_29345,N_29413);
nand UO_2292 (O_2292,N_29393,N_29149);
and UO_2293 (O_2293,N_29261,N_29273);
xnor UO_2294 (O_2294,N_29333,N_29710);
nand UO_2295 (O_2295,N_29396,N_29341);
or UO_2296 (O_2296,N_29611,N_29983);
xnor UO_2297 (O_2297,N_29303,N_29215);
nor UO_2298 (O_2298,N_29412,N_29117);
or UO_2299 (O_2299,N_29434,N_29252);
xor UO_2300 (O_2300,N_29397,N_29028);
nand UO_2301 (O_2301,N_29458,N_29772);
xnor UO_2302 (O_2302,N_29493,N_29888);
nand UO_2303 (O_2303,N_29638,N_29417);
xor UO_2304 (O_2304,N_29342,N_29353);
nor UO_2305 (O_2305,N_29224,N_29597);
nand UO_2306 (O_2306,N_29984,N_29718);
nor UO_2307 (O_2307,N_29619,N_29923);
and UO_2308 (O_2308,N_29493,N_29809);
and UO_2309 (O_2309,N_29398,N_29097);
xnor UO_2310 (O_2310,N_29003,N_29282);
or UO_2311 (O_2311,N_29725,N_29257);
and UO_2312 (O_2312,N_29200,N_29964);
xor UO_2313 (O_2313,N_29958,N_29023);
nor UO_2314 (O_2314,N_29175,N_29707);
or UO_2315 (O_2315,N_29652,N_29708);
xnor UO_2316 (O_2316,N_29065,N_29617);
nor UO_2317 (O_2317,N_29744,N_29877);
nand UO_2318 (O_2318,N_29210,N_29375);
and UO_2319 (O_2319,N_29920,N_29070);
and UO_2320 (O_2320,N_29070,N_29965);
xnor UO_2321 (O_2321,N_29615,N_29811);
nand UO_2322 (O_2322,N_29522,N_29455);
xnor UO_2323 (O_2323,N_29088,N_29164);
xor UO_2324 (O_2324,N_29552,N_29505);
or UO_2325 (O_2325,N_29635,N_29052);
xnor UO_2326 (O_2326,N_29614,N_29658);
and UO_2327 (O_2327,N_29161,N_29411);
and UO_2328 (O_2328,N_29816,N_29318);
and UO_2329 (O_2329,N_29759,N_29115);
and UO_2330 (O_2330,N_29917,N_29755);
or UO_2331 (O_2331,N_29238,N_29583);
and UO_2332 (O_2332,N_29116,N_29034);
nor UO_2333 (O_2333,N_29499,N_29506);
nand UO_2334 (O_2334,N_29735,N_29112);
nand UO_2335 (O_2335,N_29916,N_29998);
nand UO_2336 (O_2336,N_29164,N_29198);
or UO_2337 (O_2337,N_29783,N_29168);
xnor UO_2338 (O_2338,N_29040,N_29663);
nand UO_2339 (O_2339,N_29929,N_29299);
nor UO_2340 (O_2340,N_29547,N_29015);
nor UO_2341 (O_2341,N_29596,N_29639);
and UO_2342 (O_2342,N_29376,N_29019);
nand UO_2343 (O_2343,N_29305,N_29386);
nor UO_2344 (O_2344,N_29883,N_29774);
or UO_2345 (O_2345,N_29865,N_29018);
xor UO_2346 (O_2346,N_29863,N_29861);
nand UO_2347 (O_2347,N_29373,N_29787);
nand UO_2348 (O_2348,N_29759,N_29526);
or UO_2349 (O_2349,N_29924,N_29907);
nor UO_2350 (O_2350,N_29345,N_29294);
and UO_2351 (O_2351,N_29802,N_29444);
nor UO_2352 (O_2352,N_29138,N_29752);
and UO_2353 (O_2353,N_29673,N_29544);
nand UO_2354 (O_2354,N_29402,N_29455);
xnor UO_2355 (O_2355,N_29677,N_29234);
xnor UO_2356 (O_2356,N_29119,N_29391);
xor UO_2357 (O_2357,N_29224,N_29070);
nor UO_2358 (O_2358,N_29704,N_29190);
xnor UO_2359 (O_2359,N_29700,N_29443);
xnor UO_2360 (O_2360,N_29752,N_29169);
xnor UO_2361 (O_2361,N_29294,N_29793);
nand UO_2362 (O_2362,N_29189,N_29810);
nand UO_2363 (O_2363,N_29246,N_29049);
xor UO_2364 (O_2364,N_29583,N_29083);
and UO_2365 (O_2365,N_29798,N_29084);
nor UO_2366 (O_2366,N_29962,N_29241);
and UO_2367 (O_2367,N_29925,N_29356);
and UO_2368 (O_2368,N_29536,N_29610);
or UO_2369 (O_2369,N_29055,N_29805);
or UO_2370 (O_2370,N_29724,N_29045);
and UO_2371 (O_2371,N_29828,N_29075);
or UO_2372 (O_2372,N_29288,N_29145);
or UO_2373 (O_2373,N_29789,N_29315);
xor UO_2374 (O_2374,N_29797,N_29271);
xor UO_2375 (O_2375,N_29407,N_29748);
nor UO_2376 (O_2376,N_29265,N_29379);
and UO_2377 (O_2377,N_29281,N_29305);
nand UO_2378 (O_2378,N_29248,N_29809);
and UO_2379 (O_2379,N_29803,N_29589);
and UO_2380 (O_2380,N_29717,N_29637);
or UO_2381 (O_2381,N_29683,N_29208);
and UO_2382 (O_2382,N_29249,N_29402);
nor UO_2383 (O_2383,N_29158,N_29776);
or UO_2384 (O_2384,N_29180,N_29646);
nor UO_2385 (O_2385,N_29767,N_29929);
and UO_2386 (O_2386,N_29666,N_29407);
xor UO_2387 (O_2387,N_29074,N_29501);
nand UO_2388 (O_2388,N_29351,N_29080);
nor UO_2389 (O_2389,N_29944,N_29405);
xor UO_2390 (O_2390,N_29088,N_29636);
xor UO_2391 (O_2391,N_29964,N_29055);
nand UO_2392 (O_2392,N_29348,N_29138);
nand UO_2393 (O_2393,N_29390,N_29655);
or UO_2394 (O_2394,N_29384,N_29345);
and UO_2395 (O_2395,N_29584,N_29973);
or UO_2396 (O_2396,N_29044,N_29467);
and UO_2397 (O_2397,N_29340,N_29572);
nand UO_2398 (O_2398,N_29222,N_29081);
and UO_2399 (O_2399,N_29311,N_29726);
nor UO_2400 (O_2400,N_29773,N_29386);
xor UO_2401 (O_2401,N_29063,N_29284);
and UO_2402 (O_2402,N_29700,N_29072);
or UO_2403 (O_2403,N_29491,N_29070);
nand UO_2404 (O_2404,N_29626,N_29236);
nand UO_2405 (O_2405,N_29437,N_29802);
nor UO_2406 (O_2406,N_29239,N_29434);
and UO_2407 (O_2407,N_29767,N_29789);
nand UO_2408 (O_2408,N_29769,N_29858);
nor UO_2409 (O_2409,N_29869,N_29528);
or UO_2410 (O_2410,N_29109,N_29550);
and UO_2411 (O_2411,N_29614,N_29670);
nand UO_2412 (O_2412,N_29543,N_29258);
nand UO_2413 (O_2413,N_29741,N_29098);
nor UO_2414 (O_2414,N_29210,N_29388);
and UO_2415 (O_2415,N_29338,N_29479);
nand UO_2416 (O_2416,N_29199,N_29672);
nand UO_2417 (O_2417,N_29468,N_29722);
nand UO_2418 (O_2418,N_29104,N_29306);
nand UO_2419 (O_2419,N_29191,N_29765);
nand UO_2420 (O_2420,N_29107,N_29472);
nor UO_2421 (O_2421,N_29630,N_29750);
or UO_2422 (O_2422,N_29383,N_29008);
xnor UO_2423 (O_2423,N_29408,N_29080);
nand UO_2424 (O_2424,N_29655,N_29145);
nand UO_2425 (O_2425,N_29080,N_29722);
nand UO_2426 (O_2426,N_29878,N_29213);
xor UO_2427 (O_2427,N_29422,N_29947);
nand UO_2428 (O_2428,N_29768,N_29681);
nand UO_2429 (O_2429,N_29446,N_29915);
nor UO_2430 (O_2430,N_29588,N_29122);
and UO_2431 (O_2431,N_29019,N_29462);
or UO_2432 (O_2432,N_29410,N_29442);
and UO_2433 (O_2433,N_29272,N_29411);
xor UO_2434 (O_2434,N_29529,N_29133);
or UO_2435 (O_2435,N_29187,N_29628);
or UO_2436 (O_2436,N_29750,N_29824);
xor UO_2437 (O_2437,N_29682,N_29829);
and UO_2438 (O_2438,N_29453,N_29514);
nor UO_2439 (O_2439,N_29995,N_29097);
nand UO_2440 (O_2440,N_29375,N_29145);
or UO_2441 (O_2441,N_29797,N_29214);
nand UO_2442 (O_2442,N_29788,N_29747);
nand UO_2443 (O_2443,N_29452,N_29842);
nand UO_2444 (O_2444,N_29049,N_29550);
xnor UO_2445 (O_2445,N_29232,N_29730);
xor UO_2446 (O_2446,N_29771,N_29683);
xor UO_2447 (O_2447,N_29073,N_29470);
or UO_2448 (O_2448,N_29631,N_29297);
nand UO_2449 (O_2449,N_29886,N_29087);
or UO_2450 (O_2450,N_29531,N_29777);
or UO_2451 (O_2451,N_29267,N_29548);
nor UO_2452 (O_2452,N_29913,N_29732);
nand UO_2453 (O_2453,N_29892,N_29487);
and UO_2454 (O_2454,N_29885,N_29796);
nor UO_2455 (O_2455,N_29236,N_29171);
or UO_2456 (O_2456,N_29678,N_29500);
nand UO_2457 (O_2457,N_29437,N_29541);
nand UO_2458 (O_2458,N_29456,N_29952);
nand UO_2459 (O_2459,N_29107,N_29493);
nand UO_2460 (O_2460,N_29127,N_29057);
and UO_2461 (O_2461,N_29352,N_29410);
or UO_2462 (O_2462,N_29144,N_29118);
xnor UO_2463 (O_2463,N_29361,N_29302);
nor UO_2464 (O_2464,N_29299,N_29758);
nor UO_2465 (O_2465,N_29460,N_29875);
nor UO_2466 (O_2466,N_29088,N_29472);
nor UO_2467 (O_2467,N_29537,N_29254);
nor UO_2468 (O_2468,N_29817,N_29895);
nor UO_2469 (O_2469,N_29230,N_29721);
and UO_2470 (O_2470,N_29048,N_29922);
and UO_2471 (O_2471,N_29908,N_29716);
xor UO_2472 (O_2472,N_29563,N_29165);
or UO_2473 (O_2473,N_29800,N_29717);
xnor UO_2474 (O_2474,N_29416,N_29914);
xnor UO_2475 (O_2475,N_29936,N_29463);
and UO_2476 (O_2476,N_29293,N_29845);
nor UO_2477 (O_2477,N_29593,N_29909);
xor UO_2478 (O_2478,N_29590,N_29676);
or UO_2479 (O_2479,N_29764,N_29721);
nand UO_2480 (O_2480,N_29132,N_29667);
xor UO_2481 (O_2481,N_29702,N_29526);
nor UO_2482 (O_2482,N_29366,N_29259);
nand UO_2483 (O_2483,N_29492,N_29932);
or UO_2484 (O_2484,N_29616,N_29580);
and UO_2485 (O_2485,N_29804,N_29379);
nor UO_2486 (O_2486,N_29021,N_29132);
or UO_2487 (O_2487,N_29766,N_29870);
and UO_2488 (O_2488,N_29610,N_29216);
xor UO_2489 (O_2489,N_29135,N_29445);
and UO_2490 (O_2490,N_29626,N_29164);
or UO_2491 (O_2491,N_29042,N_29487);
nor UO_2492 (O_2492,N_29064,N_29248);
xor UO_2493 (O_2493,N_29361,N_29418);
nand UO_2494 (O_2494,N_29469,N_29240);
or UO_2495 (O_2495,N_29905,N_29533);
nand UO_2496 (O_2496,N_29083,N_29019);
nand UO_2497 (O_2497,N_29122,N_29786);
nor UO_2498 (O_2498,N_29902,N_29818);
xnor UO_2499 (O_2499,N_29462,N_29908);
nand UO_2500 (O_2500,N_29734,N_29448);
or UO_2501 (O_2501,N_29338,N_29589);
or UO_2502 (O_2502,N_29250,N_29025);
or UO_2503 (O_2503,N_29232,N_29596);
nor UO_2504 (O_2504,N_29942,N_29106);
and UO_2505 (O_2505,N_29488,N_29579);
xor UO_2506 (O_2506,N_29484,N_29620);
xnor UO_2507 (O_2507,N_29067,N_29613);
nor UO_2508 (O_2508,N_29177,N_29846);
or UO_2509 (O_2509,N_29391,N_29690);
nand UO_2510 (O_2510,N_29654,N_29433);
and UO_2511 (O_2511,N_29100,N_29955);
or UO_2512 (O_2512,N_29855,N_29911);
and UO_2513 (O_2513,N_29236,N_29786);
and UO_2514 (O_2514,N_29033,N_29284);
or UO_2515 (O_2515,N_29372,N_29008);
and UO_2516 (O_2516,N_29766,N_29646);
xor UO_2517 (O_2517,N_29750,N_29235);
or UO_2518 (O_2518,N_29936,N_29045);
or UO_2519 (O_2519,N_29045,N_29665);
and UO_2520 (O_2520,N_29329,N_29501);
and UO_2521 (O_2521,N_29053,N_29957);
and UO_2522 (O_2522,N_29076,N_29287);
nor UO_2523 (O_2523,N_29944,N_29803);
xnor UO_2524 (O_2524,N_29315,N_29392);
or UO_2525 (O_2525,N_29054,N_29395);
nor UO_2526 (O_2526,N_29944,N_29274);
xnor UO_2527 (O_2527,N_29754,N_29018);
nand UO_2528 (O_2528,N_29444,N_29863);
nor UO_2529 (O_2529,N_29458,N_29925);
and UO_2530 (O_2530,N_29847,N_29584);
or UO_2531 (O_2531,N_29678,N_29248);
nor UO_2532 (O_2532,N_29399,N_29115);
nor UO_2533 (O_2533,N_29952,N_29491);
and UO_2534 (O_2534,N_29417,N_29029);
or UO_2535 (O_2535,N_29443,N_29829);
xnor UO_2536 (O_2536,N_29129,N_29544);
xor UO_2537 (O_2537,N_29361,N_29512);
xor UO_2538 (O_2538,N_29846,N_29624);
or UO_2539 (O_2539,N_29248,N_29583);
nor UO_2540 (O_2540,N_29538,N_29817);
or UO_2541 (O_2541,N_29905,N_29348);
xor UO_2542 (O_2542,N_29167,N_29287);
or UO_2543 (O_2543,N_29849,N_29582);
and UO_2544 (O_2544,N_29020,N_29549);
and UO_2545 (O_2545,N_29425,N_29410);
or UO_2546 (O_2546,N_29092,N_29579);
and UO_2547 (O_2547,N_29404,N_29607);
xor UO_2548 (O_2548,N_29709,N_29987);
and UO_2549 (O_2549,N_29953,N_29537);
and UO_2550 (O_2550,N_29905,N_29843);
nand UO_2551 (O_2551,N_29168,N_29449);
xor UO_2552 (O_2552,N_29897,N_29812);
xor UO_2553 (O_2553,N_29313,N_29719);
nor UO_2554 (O_2554,N_29867,N_29369);
and UO_2555 (O_2555,N_29855,N_29508);
xnor UO_2556 (O_2556,N_29200,N_29957);
and UO_2557 (O_2557,N_29081,N_29901);
xnor UO_2558 (O_2558,N_29986,N_29823);
and UO_2559 (O_2559,N_29409,N_29902);
xnor UO_2560 (O_2560,N_29420,N_29803);
and UO_2561 (O_2561,N_29545,N_29035);
nor UO_2562 (O_2562,N_29374,N_29111);
xor UO_2563 (O_2563,N_29006,N_29324);
or UO_2564 (O_2564,N_29441,N_29827);
nor UO_2565 (O_2565,N_29976,N_29308);
nor UO_2566 (O_2566,N_29036,N_29539);
and UO_2567 (O_2567,N_29881,N_29018);
nor UO_2568 (O_2568,N_29317,N_29712);
nand UO_2569 (O_2569,N_29095,N_29621);
or UO_2570 (O_2570,N_29217,N_29196);
nor UO_2571 (O_2571,N_29952,N_29246);
nand UO_2572 (O_2572,N_29697,N_29107);
xor UO_2573 (O_2573,N_29429,N_29328);
and UO_2574 (O_2574,N_29244,N_29204);
and UO_2575 (O_2575,N_29794,N_29265);
or UO_2576 (O_2576,N_29681,N_29538);
or UO_2577 (O_2577,N_29504,N_29192);
nor UO_2578 (O_2578,N_29143,N_29877);
nand UO_2579 (O_2579,N_29919,N_29928);
nand UO_2580 (O_2580,N_29877,N_29079);
xor UO_2581 (O_2581,N_29095,N_29784);
and UO_2582 (O_2582,N_29888,N_29107);
and UO_2583 (O_2583,N_29341,N_29610);
nand UO_2584 (O_2584,N_29949,N_29453);
nor UO_2585 (O_2585,N_29378,N_29931);
nand UO_2586 (O_2586,N_29395,N_29443);
xor UO_2587 (O_2587,N_29129,N_29584);
nor UO_2588 (O_2588,N_29525,N_29639);
nor UO_2589 (O_2589,N_29412,N_29921);
and UO_2590 (O_2590,N_29713,N_29041);
and UO_2591 (O_2591,N_29781,N_29573);
xnor UO_2592 (O_2592,N_29644,N_29166);
xnor UO_2593 (O_2593,N_29290,N_29951);
nor UO_2594 (O_2594,N_29953,N_29783);
and UO_2595 (O_2595,N_29396,N_29889);
xor UO_2596 (O_2596,N_29676,N_29966);
nand UO_2597 (O_2597,N_29764,N_29477);
or UO_2598 (O_2598,N_29273,N_29367);
nand UO_2599 (O_2599,N_29281,N_29324);
nor UO_2600 (O_2600,N_29498,N_29064);
and UO_2601 (O_2601,N_29326,N_29695);
or UO_2602 (O_2602,N_29762,N_29879);
nand UO_2603 (O_2603,N_29218,N_29514);
nor UO_2604 (O_2604,N_29222,N_29456);
nor UO_2605 (O_2605,N_29148,N_29815);
nand UO_2606 (O_2606,N_29866,N_29278);
and UO_2607 (O_2607,N_29771,N_29378);
or UO_2608 (O_2608,N_29351,N_29034);
and UO_2609 (O_2609,N_29395,N_29090);
xor UO_2610 (O_2610,N_29729,N_29490);
xor UO_2611 (O_2611,N_29595,N_29794);
nand UO_2612 (O_2612,N_29250,N_29685);
nand UO_2613 (O_2613,N_29959,N_29006);
nor UO_2614 (O_2614,N_29429,N_29355);
nor UO_2615 (O_2615,N_29807,N_29664);
or UO_2616 (O_2616,N_29617,N_29703);
and UO_2617 (O_2617,N_29100,N_29204);
nor UO_2618 (O_2618,N_29511,N_29006);
or UO_2619 (O_2619,N_29452,N_29655);
or UO_2620 (O_2620,N_29321,N_29286);
nor UO_2621 (O_2621,N_29089,N_29144);
and UO_2622 (O_2622,N_29967,N_29102);
and UO_2623 (O_2623,N_29119,N_29327);
or UO_2624 (O_2624,N_29454,N_29734);
and UO_2625 (O_2625,N_29578,N_29675);
and UO_2626 (O_2626,N_29801,N_29669);
xor UO_2627 (O_2627,N_29811,N_29610);
nor UO_2628 (O_2628,N_29519,N_29510);
nand UO_2629 (O_2629,N_29245,N_29265);
and UO_2630 (O_2630,N_29385,N_29071);
or UO_2631 (O_2631,N_29797,N_29297);
xor UO_2632 (O_2632,N_29220,N_29971);
nor UO_2633 (O_2633,N_29060,N_29100);
xor UO_2634 (O_2634,N_29756,N_29389);
nand UO_2635 (O_2635,N_29010,N_29265);
or UO_2636 (O_2636,N_29698,N_29378);
nand UO_2637 (O_2637,N_29213,N_29727);
xnor UO_2638 (O_2638,N_29088,N_29215);
or UO_2639 (O_2639,N_29277,N_29664);
or UO_2640 (O_2640,N_29870,N_29455);
nand UO_2641 (O_2641,N_29962,N_29551);
xor UO_2642 (O_2642,N_29436,N_29344);
or UO_2643 (O_2643,N_29120,N_29785);
xnor UO_2644 (O_2644,N_29445,N_29348);
xnor UO_2645 (O_2645,N_29114,N_29487);
nand UO_2646 (O_2646,N_29972,N_29944);
or UO_2647 (O_2647,N_29890,N_29038);
or UO_2648 (O_2648,N_29670,N_29768);
or UO_2649 (O_2649,N_29458,N_29394);
and UO_2650 (O_2650,N_29200,N_29034);
or UO_2651 (O_2651,N_29284,N_29254);
nand UO_2652 (O_2652,N_29221,N_29457);
and UO_2653 (O_2653,N_29806,N_29587);
nand UO_2654 (O_2654,N_29570,N_29826);
nand UO_2655 (O_2655,N_29392,N_29557);
or UO_2656 (O_2656,N_29655,N_29073);
nand UO_2657 (O_2657,N_29371,N_29083);
or UO_2658 (O_2658,N_29533,N_29427);
and UO_2659 (O_2659,N_29052,N_29165);
nor UO_2660 (O_2660,N_29691,N_29733);
and UO_2661 (O_2661,N_29661,N_29905);
nand UO_2662 (O_2662,N_29363,N_29051);
nand UO_2663 (O_2663,N_29320,N_29170);
xor UO_2664 (O_2664,N_29537,N_29962);
and UO_2665 (O_2665,N_29681,N_29862);
or UO_2666 (O_2666,N_29381,N_29031);
nand UO_2667 (O_2667,N_29817,N_29027);
or UO_2668 (O_2668,N_29892,N_29854);
nand UO_2669 (O_2669,N_29888,N_29203);
or UO_2670 (O_2670,N_29492,N_29273);
xor UO_2671 (O_2671,N_29558,N_29733);
or UO_2672 (O_2672,N_29435,N_29879);
xnor UO_2673 (O_2673,N_29604,N_29038);
nand UO_2674 (O_2674,N_29864,N_29369);
nand UO_2675 (O_2675,N_29265,N_29543);
and UO_2676 (O_2676,N_29700,N_29805);
nand UO_2677 (O_2677,N_29086,N_29879);
nand UO_2678 (O_2678,N_29956,N_29408);
nor UO_2679 (O_2679,N_29703,N_29119);
or UO_2680 (O_2680,N_29872,N_29107);
nand UO_2681 (O_2681,N_29843,N_29706);
and UO_2682 (O_2682,N_29589,N_29853);
nor UO_2683 (O_2683,N_29982,N_29773);
xor UO_2684 (O_2684,N_29522,N_29267);
nand UO_2685 (O_2685,N_29842,N_29155);
nor UO_2686 (O_2686,N_29682,N_29054);
or UO_2687 (O_2687,N_29526,N_29481);
xor UO_2688 (O_2688,N_29373,N_29873);
nor UO_2689 (O_2689,N_29284,N_29453);
nand UO_2690 (O_2690,N_29898,N_29426);
nand UO_2691 (O_2691,N_29980,N_29416);
nand UO_2692 (O_2692,N_29760,N_29700);
or UO_2693 (O_2693,N_29958,N_29912);
nor UO_2694 (O_2694,N_29241,N_29320);
or UO_2695 (O_2695,N_29357,N_29873);
and UO_2696 (O_2696,N_29023,N_29151);
nor UO_2697 (O_2697,N_29528,N_29072);
nand UO_2698 (O_2698,N_29323,N_29246);
xnor UO_2699 (O_2699,N_29949,N_29778);
or UO_2700 (O_2700,N_29500,N_29397);
xor UO_2701 (O_2701,N_29508,N_29947);
xnor UO_2702 (O_2702,N_29566,N_29700);
xor UO_2703 (O_2703,N_29811,N_29716);
and UO_2704 (O_2704,N_29577,N_29364);
or UO_2705 (O_2705,N_29141,N_29170);
nand UO_2706 (O_2706,N_29057,N_29059);
nand UO_2707 (O_2707,N_29725,N_29652);
and UO_2708 (O_2708,N_29197,N_29131);
xor UO_2709 (O_2709,N_29934,N_29804);
xnor UO_2710 (O_2710,N_29318,N_29648);
xor UO_2711 (O_2711,N_29221,N_29556);
and UO_2712 (O_2712,N_29804,N_29729);
nand UO_2713 (O_2713,N_29718,N_29694);
and UO_2714 (O_2714,N_29832,N_29555);
nor UO_2715 (O_2715,N_29995,N_29861);
and UO_2716 (O_2716,N_29331,N_29241);
nor UO_2717 (O_2717,N_29439,N_29843);
nor UO_2718 (O_2718,N_29543,N_29089);
or UO_2719 (O_2719,N_29347,N_29480);
xnor UO_2720 (O_2720,N_29349,N_29385);
xnor UO_2721 (O_2721,N_29196,N_29615);
or UO_2722 (O_2722,N_29034,N_29291);
or UO_2723 (O_2723,N_29439,N_29887);
or UO_2724 (O_2724,N_29900,N_29815);
nor UO_2725 (O_2725,N_29143,N_29544);
xor UO_2726 (O_2726,N_29961,N_29954);
and UO_2727 (O_2727,N_29512,N_29132);
nor UO_2728 (O_2728,N_29417,N_29886);
and UO_2729 (O_2729,N_29815,N_29564);
xnor UO_2730 (O_2730,N_29133,N_29272);
nor UO_2731 (O_2731,N_29025,N_29750);
and UO_2732 (O_2732,N_29808,N_29096);
xnor UO_2733 (O_2733,N_29366,N_29689);
and UO_2734 (O_2734,N_29546,N_29324);
nand UO_2735 (O_2735,N_29565,N_29486);
or UO_2736 (O_2736,N_29247,N_29069);
and UO_2737 (O_2737,N_29971,N_29550);
nor UO_2738 (O_2738,N_29515,N_29918);
and UO_2739 (O_2739,N_29081,N_29618);
nor UO_2740 (O_2740,N_29068,N_29834);
nor UO_2741 (O_2741,N_29145,N_29367);
xnor UO_2742 (O_2742,N_29090,N_29227);
nor UO_2743 (O_2743,N_29610,N_29746);
xor UO_2744 (O_2744,N_29220,N_29039);
xnor UO_2745 (O_2745,N_29921,N_29950);
xor UO_2746 (O_2746,N_29076,N_29542);
nand UO_2747 (O_2747,N_29120,N_29649);
nand UO_2748 (O_2748,N_29235,N_29048);
or UO_2749 (O_2749,N_29773,N_29328);
xnor UO_2750 (O_2750,N_29208,N_29012);
and UO_2751 (O_2751,N_29621,N_29645);
or UO_2752 (O_2752,N_29833,N_29586);
and UO_2753 (O_2753,N_29512,N_29826);
or UO_2754 (O_2754,N_29589,N_29850);
nand UO_2755 (O_2755,N_29813,N_29428);
nor UO_2756 (O_2756,N_29474,N_29382);
and UO_2757 (O_2757,N_29620,N_29682);
xnor UO_2758 (O_2758,N_29404,N_29760);
and UO_2759 (O_2759,N_29459,N_29258);
xnor UO_2760 (O_2760,N_29756,N_29648);
xnor UO_2761 (O_2761,N_29147,N_29375);
nand UO_2762 (O_2762,N_29223,N_29474);
nand UO_2763 (O_2763,N_29518,N_29509);
or UO_2764 (O_2764,N_29586,N_29215);
nor UO_2765 (O_2765,N_29585,N_29209);
xnor UO_2766 (O_2766,N_29459,N_29509);
nand UO_2767 (O_2767,N_29637,N_29832);
or UO_2768 (O_2768,N_29296,N_29168);
or UO_2769 (O_2769,N_29626,N_29358);
or UO_2770 (O_2770,N_29703,N_29772);
nor UO_2771 (O_2771,N_29648,N_29203);
nor UO_2772 (O_2772,N_29358,N_29482);
nand UO_2773 (O_2773,N_29225,N_29932);
or UO_2774 (O_2774,N_29694,N_29983);
nor UO_2775 (O_2775,N_29269,N_29987);
and UO_2776 (O_2776,N_29872,N_29899);
nand UO_2777 (O_2777,N_29870,N_29312);
nand UO_2778 (O_2778,N_29579,N_29905);
or UO_2779 (O_2779,N_29005,N_29763);
nor UO_2780 (O_2780,N_29235,N_29889);
or UO_2781 (O_2781,N_29119,N_29164);
xor UO_2782 (O_2782,N_29347,N_29097);
xnor UO_2783 (O_2783,N_29771,N_29734);
nor UO_2784 (O_2784,N_29042,N_29541);
and UO_2785 (O_2785,N_29358,N_29068);
and UO_2786 (O_2786,N_29800,N_29297);
nor UO_2787 (O_2787,N_29971,N_29832);
nand UO_2788 (O_2788,N_29012,N_29175);
nor UO_2789 (O_2789,N_29615,N_29478);
or UO_2790 (O_2790,N_29424,N_29225);
or UO_2791 (O_2791,N_29204,N_29721);
or UO_2792 (O_2792,N_29008,N_29150);
nor UO_2793 (O_2793,N_29625,N_29838);
nor UO_2794 (O_2794,N_29554,N_29327);
nor UO_2795 (O_2795,N_29290,N_29839);
or UO_2796 (O_2796,N_29981,N_29304);
xnor UO_2797 (O_2797,N_29582,N_29098);
and UO_2798 (O_2798,N_29219,N_29472);
nand UO_2799 (O_2799,N_29860,N_29340);
nor UO_2800 (O_2800,N_29388,N_29473);
nand UO_2801 (O_2801,N_29180,N_29615);
or UO_2802 (O_2802,N_29249,N_29092);
nand UO_2803 (O_2803,N_29597,N_29903);
and UO_2804 (O_2804,N_29591,N_29592);
xnor UO_2805 (O_2805,N_29716,N_29476);
nor UO_2806 (O_2806,N_29010,N_29929);
nor UO_2807 (O_2807,N_29005,N_29625);
xnor UO_2808 (O_2808,N_29313,N_29158);
or UO_2809 (O_2809,N_29607,N_29733);
xor UO_2810 (O_2810,N_29824,N_29379);
or UO_2811 (O_2811,N_29497,N_29733);
xnor UO_2812 (O_2812,N_29475,N_29484);
xor UO_2813 (O_2813,N_29161,N_29587);
nor UO_2814 (O_2814,N_29365,N_29156);
nand UO_2815 (O_2815,N_29764,N_29194);
and UO_2816 (O_2816,N_29915,N_29113);
nor UO_2817 (O_2817,N_29587,N_29969);
nand UO_2818 (O_2818,N_29352,N_29712);
nor UO_2819 (O_2819,N_29662,N_29550);
or UO_2820 (O_2820,N_29618,N_29262);
xnor UO_2821 (O_2821,N_29521,N_29890);
and UO_2822 (O_2822,N_29953,N_29458);
or UO_2823 (O_2823,N_29569,N_29939);
xor UO_2824 (O_2824,N_29666,N_29560);
nor UO_2825 (O_2825,N_29637,N_29184);
nand UO_2826 (O_2826,N_29662,N_29316);
nand UO_2827 (O_2827,N_29627,N_29031);
xor UO_2828 (O_2828,N_29398,N_29671);
and UO_2829 (O_2829,N_29152,N_29361);
nor UO_2830 (O_2830,N_29552,N_29514);
and UO_2831 (O_2831,N_29091,N_29070);
nand UO_2832 (O_2832,N_29459,N_29762);
xnor UO_2833 (O_2833,N_29157,N_29390);
xor UO_2834 (O_2834,N_29652,N_29687);
and UO_2835 (O_2835,N_29926,N_29387);
or UO_2836 (O_2836,N_29688,N_29458);
or UO_2837 (O_2837,N_29476,N_29350);
and UO_2838 (O_2838,N_29161,N_29326);
nor UO_2839 (O_2839,N_29426,N_29895);
or UO_2840 (O_2840,N_29222,N_29523);
and UO_2841 (O_2841,N_29166,N_29295);
nor UO_2842 (O_2842,N_29727,N_29552);
or UO_2843 (O_2843,N_29170,N_29031);
nand UO_2844 (O_2844,N_29865,N_29897);
xnor UO_2845 (O_2845,N_29431,N_29544);
xnor UO_2846 (O_2846,N_29615,N_29164);
or UO_2847 (O_2847,N_29662,N_29578);
nand UO_2848 (O_2848,N_29356,N_29226);
nand UO_2849 (O_2849,N_29279,N_29510);
or UO_2850 (O_2850,N_29425,N_29421);
and UO_2851 (O_2851,N_29692,N_29807);
and UO_2852 (O_2852,N_29734,N_29256);
nor UO_2853 (O_2853,N_29359,N_29652);
and UO_2854 (O_2854,N_29081,N_29920);
and UO_2855 (O_2855,N_29413,N_29639);
xor UO_2856 (O_2856,N_29045,N_29340);
xor UO_2857 (O_2857,N_29563,N_29658);
and UO_2858 (O_2858,N_29592,N_29404);
nor UO_2859 (O_2859,N_29702,N_29954);
nand UO_2860 (O_2860,N_29027,N_29885);
and UO_2861 (O_2861,N_29217,N_29520);
nand UO_2862 (O_2862,N_29701,N_29752);
or UO_2863 (O_2863,N_29635,N_29900);
nor UO_2864 (O_2864,N_29371,N_29850);
nand UO_2865 (O_2865,N_29505,N_29190);
and UO_2866 (O_2866,N_29828,N_29845);
nor UO_2867 (O_2867,N_29394,N_29401);
nand UO_2868 (O_2868,N_29388,N_29094);
nand UO_2869 (O_2869,N_29742,N_29402);
xnor UO_2870 (O_2870,N_29446,N_29846);
nor UO_2871 (O_2871,N_29179,N_29311);
xor UO_2872 (O_2872,N_29331,N_29108);
xor UO_2873 (O_2873,N_29704,N_29632);
or UO_2874 (O_2874,N_29889,N_29641);
or UO_2875 (O_2875,N_29640,N_29413);
xor UO_2876 (O_2876,N_29316,N_29226);
and UO_2877 (O_2877,N_29203,N_29724);
xnor UO_2878 (O_2878,N_29610,N_29537);
nor UO_2879 (O_2879,N_29103,N_29750);
or UO_2880 (O_2880,N_29620,N_29426);
nor UO_2881 (O_2881,N_29370,N_29664);
xor UO_2882 (O_2882,N_29193,N_29090);
or UO_2883 (O_2883,N_29278,N_29485);
nor UO_2884 (O_2884,N_29695,N_29779);
and UO_2885 (O_2885,N_29179,N_29583);
nor UO_2886 (O_2886,N_29009,N_29617);
nor UO_2887 (O_2887,N_29132,N_29618);
xor UO_2888 (O_2888,N_29180,N_29949);
or UO_2889 (O_2889,N_29774,N_29890);
xnor UO_2890 (O_2890,N_29310,N_29888);
nand UO_2891 (O_2891,N_29344,N_29047);
nand UO_2892 (O_2892,N_29007,N_29463);
nand UO_2893 (O_2893,N_29903,N_29861);
and UO_2894 (O_2894,N_29806,N_29181);
or UO_2895 (O_2895,N_29240,N_29124);
nor UO_2896 (O_2896,N_29597,N_29163);
nor UO_2897 (O_2897,N_29456,N_29517);
or UO_2898 (O_2898,N_29389,N_29567);
xnor UO_2899 (O_2899,N_29357,N_29743);
nand UO_2900 (O_2900,N_29337,N_29693);
and UO_2901 (O_2901,N_29614,N_29976);
xor UO_2902 (O_2902,N_29137,N_29101);
nand UO_2903 (O_2903,N_29435,N_29587);
xor UO_2904 (O_2904,N_29822,N_29939);
or UO_2905 (O_2905,N_29456,N_29662);
or UO_2906 (O_2906,N_29450,N_29198);
and UO_2907 (O_2907,N_29827,N_29207);
nor UO_2908 (O_2908,N_29405,N_29777);
nand UO_2909 (O_2909,N_29560,N_29021);
nor UO_2910 (O_2910,N_29980,N_29837);
xor UO_2911 (O_2911,N_29964,N_29001);
nand UO_2912 (O_2912,N_29504,N_29953);
and UO_2913 (O_2913,N_29139,N_29304);
xnor UO_2914 (O_2914,N_29385,N_29045);
or UO_2915 (O_2915,N_29618,N_29658);
nand UO_2916 (O_2916,N_29520,N_29540);
xor UO_2917 (O_2917,N_29944,N_29936);
nor UO_2918 (O_2918,N_29426,N_29715);
nand UO_2919 (O_2919,N_29891,N_29344);
or UO_2920 (O_2920,N_29204,N_29503);
and UO_2921 (O_2921,N_29016,N_29401);
nor UO_2922 (O_2922,N_29771,N_29952);
xor UO_2923 (O_2923,N_29909,N_29377);
and UO_2924 (O_2924,N_29607,N_29084);
and UO_2925 (O_2925,N_29754,N_29538);
nor UO_2926 (O_2926,N_29196,N_29707);
and UO_2927 (O_2927,N_29949,N_29669);
or UO_2928 (O_2928,N_29251,N_29333);
nand UO_2929 (O_2929,N_29449,N_29240);
xor UO_2930 (O_2930,N_29576,N_29175);
or UO_2931 (O_2931,N_29194,N_29706);
nand UO_2932 (O_2932,N_29855,N_29856);
or UO_2933 (O_2933,N_29884,N_29219);
nor UO_2934 (O_2934,N_29165,N_29959);
nor UO_2935 (O_2935,N_29636,N_29075);
nor UO_2936 (O_2936,N_29633,N_29099);
or UO_2937 (O_2937,N_29866,N_29979);
nand UO_2938 (O_2938,N_29175,N_29070);
or UO_2939 (O_2939,N_29053,N_29594);
and UO_2940 (O_2940,N_29920,N_29907);
nand UO_2941 (O_2941,N_29682,N_29845);
or UO_2942 (O_2942,N_29087,N_29826);
or UO_2943 (O_2943,N_29251,N_29038);
xnor UO_2944 (O_2944,N_29436,N_29787);
and UO_2945 (O_2945,N_29586,N_29892);
nor UO_2946 (O_2946,N_29005,N_29889);
or UO_2947 (O_2947,N_29151,N_29573);
and UO_2948 (O_2948,N_29443,N_29381);
or UO_2949 (O_2949,N_29286,N_29012);
nand UO_2950 (O_2950,N_29800,N_29678);
nor UO_2951 (O_2951,N_29508,N_29378);
nor UO_2952 (O_2952,N_29630,N_29131);
xnor UO_2953 (O_2953,N_29859,N_29848);
or UO_2954 (O_2954,N_29079,N_29094);
nand UO_2955 (O_2955,N_29642,N_29988);
and UO_2956 (O_2956,N_29675,N_29754);
nand UO_2957 (O_2957,N_29123,N_29993);
xnor UO_2958 (O_2958,N_29838,N_29093);
nand UO_2959 (O_2959,N_29042,N_29360);
or UO_2960 (O_2960,N_29594,N_29587);
nand UO_2961 (O_2961,N_29600,N_29531);
xnor UO_2962 (O_2962,N_29297,N_29423);
xor UO_2963 (O_2963,N_29418,N_29517);
or UO_2964 (O_2964,N_29341,N_29291);
nor UO_2965 (O_2965,N_29217,N_29426);
and UO_2966 (O_2966,N_29811,N_29962);
xnor UO_2967 (O_2967,N_29179,N_29021);
nor UO_2968 (O_2968,N_29121,N_29907);
or UO_2969 (O_2969,N_29407,N_29602);
nor UO_2970 (O_2970,N_29954,N_29763);
and UO_2971 (O_2971,N_29407,N_29060);
xor UO_2972 (O_2972,N_29639,N_29839);
nor UO_2973 (O_2973,N_29384,N_29847);
or UO_2974 (O_2974,N_29997,N_29955);
xor UO_2975 (O_2975,N_29704,N_29883);
and UO_2976 (O_2976,N_29761,N_29671);
and UO_2977 (O_2977,N_29997,N_29225);
or UO_2978 (O_2978,N_29024,N_29622);
nand UO_2979 (O_2979,N_29450,N_29157);
and UO_2980 (O_2980,N_29482,N_29435);
xnor UO_2981 (O_2981,N_29090,N_29736);
and UO_2982 (O_2982,N_29145,N_29909);
or UO_2983 (O_2983,N_29903,N_29875);
nand UO_2984 (O_2984,N_29708,N_29478);
and UO_2985 (O_2985,N_29594,N_29432);
xnor UO_2986 (O_2986,N_29084,N_29177);
or UO_2987 (O_2987,N_29390,N_29025);
nor UO_2988 (O_2988,N_29864,N_29099);
and UO_2989 (O_2989,N_29798,N_29490);
xnor UO_2990 (O_2990,N_29285,N_29422);
or UO_2991 (O_2991,N_29406,N_29120);
nor UO_2992 (O_2992,N_29283,N_29756);
nand UO_2993 (O_2993,N_29055,N_29448);
xor UO_2994 (O_2994,N_29920,N_29468);
nand UO_2995 (O_2995,N_29261,N_29140);
and UO_2996 (O_2996,N_29991,N_29145);
and UO_2997 (O_2997,N_29067,N_29680);
nand UO_2998 (O_2998,N_29059,N_29163);
nand UO_2999 (O_2999,N_29351,N_29909);
or UO_3000 (O_3000,N_29174,N_29475);
nand UO_3001 (O_3001,N_29624,N_29457);
and UO_3002 (O_3002,N_29290,N_29869);
and UO_3003 (O_3003,N_29310,N_29435);
nand UO_3004 (O_3004,N_29295,N_29256);
nor UO_3005 (O_3005,N_29263,N_29629);
nor UO_3006 (O_3006,N_29935,N_29747);
and UO_3007 (O_3007,N_29380,N_29910);
or UO_3008 (O_3008,N_29012,N_29751);
nor UO_3009 (O_3009,N_29443,N_29175);
and UO_3010 (O_3010,N_29370,N_29942);
xnor UO_3011 (O_3011,N_29747,N_29631);
and UO_3012 (O_3012,N_29849,N_29917);
xnor UO_3013 (O_3013,N_29345,N_29610);
or UO_3014 (O_3014,N_29697,N_29511);
nor UO_3015 (O_3015,N_29537,N_29388);
xnor UO_3016 (O_3016,N_29088,N_29981);
nor UO_3017 (O_3017,N_29308,N_29836);
and UO_3018 (O_3018,N_29740,N_29910);
nand UO_3019 (O_3019,N_29201,N_29439);
xnor UO_3020 (O_3020,N_29481,N_29743);
nor UO_3021 (O_3021,N_29864,N_29938);
and UO_3022 (O_3022,N_29475,N_29822);
nand UO_3023 (O_3023,N_29167,N_29755);
nor UO_3024 (O_3024,N_29798,N_29848);
and UO_3025 (O_3025,N_29030,N_29374);
and UO_3026 (O_3026,N_29131,N_29615);
and UO_3027 (O_3027,N_29973,N_29712);
xnor UO_3028 (O_3028,N_29832,N_29784);
nor UO_3029 (O_3029,N_29328,N_29316);
xor UO_3030 (O_3030,N_29210,N_29667);
xnor UO_3031 (O_3031,N_29411,N_29763);
xor UO_3032 (O_3032,N_29942,N_29205);
nand UO_3033 (O_3033,N_29969,N_29644);
xor UO_3034 (O_3034,N_29296,N_29569);
nand UO_3035 (O_3035,N_29426,N_29530);
and UO_3036 (O_3036,N_29620,N_29146);
and UO_3037 (O_3037,N_29938,N_29307);
nand UO_3038 (O_3038,N_29569,N_29779);
or UO_3039 (O_3039,N_29327,N_29125);
xor UO_3040 (O_3040,N_29258,N_29846);
and UO_3041 (O_3041,N_29821,N_29581);
xnor UO_3042 (O_3042,N_29893,N_29086);
and UO_3043 (O_3043,N_29244,N_29419);
or UO_3044 (O_3044,N_29995,N_29518);
nor UO_3045 (O_3045,N_29431,N_29981);
and UO_3046 (O_3046,N_29512,N_29866);
or UO_3047 (O_3047,N_29703,N_29236);
xor UO_3048 (O_3048,N_29709,N_29693);
and UO_3049 (O_3049,N_29105,N_29759);
and UO_3050 (O_3050,N_29275,N_29035);
and UO_3051 (O_3051,N_29982,N_29289);
xor UO_3052 (O_3052,N_29791,N_29072);
xor UO_3053 (O_3053,N_29369,N_29895);
or UO_3054 (O_3054,N_29748,N_29212);
xnor UO_3055 (O_3055,N_29948,N_29812);
nand UO_3056 (O_3056,N_29859,N_29367);
nor UO_3057 (O_3057,N_29354,N_29157);
or UO_3058 (O_3058,N_29527,N_29136);
nand UO_3059 (O_3059,N_29017,N_29883);
or UO_3060 (O_3060,N_29760,N_29705);
and UO_3061 (O_3061,N_29656,N_29719);
xnor UO_3062 (O_3062,N_29384,N_29323);
or UO_3063 (O_3063,N_29875,N_29898);
nand UO_3064 (O_3064,N_29096,N_29190);
nand UO_3065 (O_3065,N_29595,N_29224);
xnor UO_3066 (O_3066,N_29765,N_29341);
and UO_3067 (O_3067,N_29479,N_29499);
nand UO_3068 (O_3068,N_29181,N_29512);
and UO_3069 (O_3069,N_29002,N_29465);
nor UO_3070 (O_3070,N_29918,N_29247);
and UO_3071 (O_3071,N_29945,N_29150);
and UO_3072 (O_3072,N_29791,N_29819);
nor UO_3073 (O_3073,N_29850,N_29016);
nor UO_3074 (O_3074,N_29740,N_29240);
nand UO_3075 (O_3075,N_29992,N_29778);
nor UO_3076 (O_3076,N_29893,N_29772);
and UO_3077 (O_3077,N_29369,N_29484);
nand UO_3078 (O_3078,N_29537,N_29121);
nor UO_3079 (O_3079,N_29555,N_29450);
and UO_3080 (O_3080,N_29193,N_29504);
nand UO_3081 (O_3081,N_29222,N_29748);
and UO_3082 (O_3082,N_29399,N_29820);
nand UO_3083 (O_3083,N_29135,N_29936);
xor UO_3084 (O_3084,N_29372,N_29890);
and UO_3085 (O_3085,N_29538,N_29654);
nand UO_3086 (O_3086,N_29196,N_29321);
xor UO_3087 (O_3087,N_29947,N_29924);
nor UO_3088 (O_3088,N_29011,N_29174);
xnor UO_3089 (O_3089,N_29982,N_29166);
nand UO_3090 (O_3090,N_29471,N_29354);
nor UO_3091 (O_3091,N_29827,N_29222);
nand UO_3092 (O_3092,N_29330,N_29774);
xor UO_3093 (O_3093,N_29329,N_29074);
and UO_3094 (O_3094,N_29441,N_29171);
xor UO_3095 (O_3095,N_29480,N_29115);
xor UO_3096 (O_3096,N_29079,N_29631);
nand UO_3097 (O_3097,N_29711,N_29869);
and UO_3098 (O_3098,N_29556,N_29948);
nor UO_3099 (O_3099,N_29824,N_29940);
xnor UO_3100 (O_3100,N_29699,N_29378);
or UO_3101 (O_3101,N_29170,N_29811);
and UO_3102 (O_3102,N_29090,N_29813);
or UO_3103 (O_3103,N_29438,N_29764);
xor UO_3104 (O_3104,N_29580,N_29327);
and UO_3105 (O_3105,N_29131,N_29255);
xnor UO_3106 (O_3106,N_29384,N_29069);
xnor UO_3107 (O_3107,N_29503,N_29271);
nor UO_3108 (O_3108,N_29981,N_29413);
or UO_3109 (O_3109,N_29934,N_29708);
and UO_3110 (O_3110,N_29117,N_29083);
or UO_3111 (O_3111,N_29009,N_29936);
and UO_3112 (O_3112,N_29214,N_29659);
nand UO_3113 (O_3113,N_29941,N_29057);
or UO_3114 (O_3114,N_29702,N_29212);
xnor UO_3115 (O_3115,N_29952,N_29530);
and UO_3116 (O_3116,N_29268,N_29671);
nand UO_3117 (O_3117,N_29075,N_29094);
xor UO_3118 (O_3118,N_29918,N_29601);
or UO_3119 (O_3119,N_29496,N_29434);
nand UO_3120 (O_3120,N_29792,N_29511);
nand UO_3121 (O_3121,N_29788,N_29275);
or UO_3122 (O_3122,N_29797,N_29990);
and UO_3123 (O_3123,N_29247,N_29436);
and UO_3124 (O_3124,N_29711,N_29000);
or UO_3125 (O_3125,N_29179,N_29383);
or UO_3126 (O_3126,N_29642,N_29168);
or UO_3127 (O_3127,N_29161,N_29501);
xnor UO_3128 (O_3128,N_29228,N_29094);
nor UO_3129 (O_3129,N_29905,N_29604);
xor UO_3130 (O_3130,N_29334,N_29977);
nand UO_3131 (O_3131,N_29027,N_29468);
or UO_3132 (O_3132,N_29118,N_29776);
nor UO_3133 (O_3133,N_29908,N_29431);
and UO_3134 (O_3134,N_29211,N_29706);
xor UO_3135 (O_3135,N_29840,N_29589);
nor UO_3136 (O_3136,N_29553,N_29939);
nor UO_3137 (O_3137,N_29882,N_29822);
nor UO_3138 (O_3138,N_29127,N_29285);
nor UO_3139 (O_3139,N_29637,N_29430);
nand UO_3140 (O_3140,N_29181,N_29159);
nor UO_3141 (O_3141,N_29425,N_29495);
or UO_3142 (O_3142,N_29117,N_29831);
and UO_3143 (O_3143,N_29318,N_29402);
and UO_3144 (O_3144,N_29838,N_29424);
nor UO_3145 (O_3145,N_29568,N_29251);
nor UO_3146 (O_3146,N_29990,N_29689);
and UO_3147 (O_3147,N_29536,N_29567);
or UO_3148 (O_3148,N_29193,N_29180);
xnor UO_3149 (O_3149,N_29274,N_29410);
nand UO_3150 (O_3150,N_29382,N_29222);
nand UO_3151 (O_3151,N_29094,N_29577);
and UO_3152 (O_3152,N_29632,N_29206);
xnor UO_3153 (O_3153,N_29391,N_29334);
xor UO_3154 (O_3154,N_29442,N_29500);
and UO_3155 (O_3155,N_29030,N_29403);
xnor UO_3156 (O_3156,N_29638,N_29164);
xor UO_3157 (O_3157,N_29758,N_29854);
xnor UO_3158 (O_3158,N_29040,N_29352);
and UO_3159 (O_3159,N_29968,N_29525);
xnor UO_3160 (O_3160,N_29900,N_29786);
nand UO_3161 (O_3161,N_29046,N_29212);
and UO_3162 (O_3162,N_29676,N_29020);
nand UO_3163 (O_3163,N_29098,N_29884);
nor UO_3164 (O_3164,N_29374,N_29292);
xor UO_3165 (O_3165,N_29783,N_29468);
nand UO_3166 (O_3166,N_29456,N_29933);
xnor UO_3167 (O_3167,N_29920,N_29113);
nand UO_3168 (O_3168,N_29585,N_29851);
nor UO_3169 (O_3169,N_29656,N_29591);
or UO_3170 (O_3170,N_29027,N_29325);
or UO_3171 (O_3171,N_29236,N_29367);
nor UO_3172 (O_3172,N_29882,N_29464);
and UO_3173 (O_3173,N_29219,N_29987);
or UO_3174 (O_3174,N_29873,N_29564);
xnor UO_3175 (O_3175,N_29000,N_29293);
xor UO_3176 (O_3176,N_29800,N_29102);
xnor UO_3177 (O_3177,N_29912,N_29279);
xor UO_3178 (O_3178,N_29996,N_29370);
xnor UO_3179 (O_3179,N_29403,N_29889);
nand UO_3180 (O_3180,N_29772,N_29135);
and UO_3181 (O_3181,N_29140,N_29547);
nor UO_3182 (O_3182,N_29307,N_29106);
nand UO_3183 (O_3183,N_29911,N_29062);
xnor UO_3184 (O_3184,N_29742,N_29896);
nor UO_3185 (O_3185,N_29753,N_29443);
or UO_3186 (O_3186,N_29850,N_29086);
nor UO_3187 (O_3187,N_29563,N_29928);
nand UO_3188 (O_3188,N_29177,N_29565);
and UO_3189 (O_3189,N_29126,N_29109);
nor UO_3190 (O_3190,N_29806,N_29118);
nand UO_3191 (O_3191,N_29526,N_29173);
xor UO_3192 (O_3192,N_29516,N_29968);
and UO_3193 (O_3193,N_29374,N_29979);
or UO_3194 (O_3194,N_29331,N_29607);
nor UO_3195 (O_3195,N_29454,N_29389);
nor UO_3196 (O_3196,N_29544,N_29255);
and UO_3197 (O_3197,N_29594,N_29665);
xnor UO_3198 (O_3198,N_29911,N_29444);
nand UO_3199 (O_3199,N_29689,N_29343);
or UO_3200 (O_3200,N_29985,N_29178);
or UO_3201 (O_3201,N_29036,N_29447);
and UO_3202 (O_3202,N_29342,N_29621);
and UO_3203 (O_3203,N_29213,N_29001);
or UO_3204 (O_3204,N_29683,N_29870);
or UO_3205 (O_3205,N_29250,N_29583);
nand UO_3206 (O_3206,N_29035,N_29052);
nand UO_3207 (O_3207,N_29222,N_29953);
nor UO_3208 (O_3208,N_29580,N_29047);
nand UO_3209 (O_3209,N_29625,N_29313);
nand UO_3210 (O_3210,N_29223,N_29854);
or UO_3211 (O_3211,N_29695,N_29761);
nor UO_3212 (O_3212,N_29927,N_29993);
xnor UO_3213 (O_3213,N_29955,N_29409);
xor UO_3214 (O_3214,N_29574,N_29683);
nor UO_3215 (O_3215,N_29505,N_29104);
xnor UO_3216 (O_3216,N_29588,N_29268);
nand UO_3217 (O_3217,N_29091,N_29015);
or UO_3218 (O_3218,N_29581,N_29443);
and UO_3219 (O_3219,N_29275,N_29467);
nor UO_3220 (O_3220,N_29917,N_29670);
nor UO_3221 (O_3221,N_29683,N_29994);
or UO_3222 (O_3222,N_29319,N_29561);
or UO_3223 (O_3223,N_29629,N_29438);
nand UO_3224 (O_3224,N_29274,N_29522);
nor UO_3225 (O_3225,N_29017,N_29788);
and UO_3226 (O_3226,N_29380,N_29047);
and UO_3227 (O_3227,N_29965,N_29285);
nand UO_3228 (O_3228,N_29400,N_29787);
nor UO_3229 (O_3229,N_29037,N_29036);
or UO_3230 (O_3230,N_29257,N_29100);
nand UO_3231 (O_3231,N_29418,N_29965);
nor UO_3232 (O_3232,N_29121,N_29594);
nor UO_3233 (O_3233,N_29201,N_29946);
and UO_3234 (O_3234,N_29477,N_29603);
nor UO_3235 (O_3235,N_29047,N_29476);
nor UO_3236 (O_3236,N_29783,N_29407);
nand UO_3237 (O_3237,N_29232,N_29630);
or UO_3238 (O_3238,N_29890,N_29639);
nand UO_3239 (O_3239,N_29615,N_29186);
nor UO_3240 (O_3240,N_29519,N_29736);
nand UO_3241 (O_3241,N_29222,N_29226);
xnor UO_3242 (O_3242,N_29656,N_29482);
nor UO_3243 (O_3243,N_29340,N_29312);
nor UO_3244 (O_3244,N_29234,N_29252);
nor UO_3245 (O_3245,N_29915,N_29857);
nand UO_3246 (O_3246,N_29374,N_29691);
nor UO_3247 (O_3247,N_29249,N_29581);
xnor UO_3248 (O_3248,N_29839,N_29121);
or UO_3249 (O_3249,N_29076,N_29722);
xnor UO_3250 (O_3250,N_29360,N_29650);
xnor UO_3251 (O_3251,N_29175,N_29085);
xnor UO_3252 (O_3252,N_29469,N_29264);
nand UO_3253 (O_3253,N_29377,N_29080);
and UO_3254 (O_3254,N_29045,N_29671);
and UO_3255 (O_3255,N_29257,N_29091);
xor UO_3256 (O_3256,N_29118,N_29163);
nand UO_3257 (O_3257,N_29642,N_29779);
and UO_3258 (O_3258,N_29576,N_29783);
and UO_3259 (O_3259,N_29651,N_29620);
or UO_3260 (O_3260,N_29873,N_29838);
xnor UO_3261 (O_3261,N_29523,N_29235);
and UO_3262 (O_3262,N_29133,N_29155);
nand UO_3263 (O_3263,N_29305,N_29629);
nor UO_3264 (O_3264,N_29398,N_29808);
xor UO_3265 (O_3265,N_29448,N_29834);
or UO_3266 (O_3266,N_29513,N_29710);
xnor UO_3267 (O_3267,N_29263,N_29846);
xor UO_3268 (O_3268,N_29227,N_29629);
nor UO_3269 (O_3269,N_29281,N_29138);
nor UO_3270 (O_3270,N_29218,N_29566);
and UO_3271 (O_3271,N_29219,N_29815);
xnor UO_3272 (O_3272,N_29045,N_29982);
xor UO_3273 (O_3273,N_29877,N_29847);
xor UO_3274 (O_3274,N_29601,N_29236);
and UO_3275 (O_3275,N_29718,N_29292);
and UO_3276 (O_3276,N_29481,N_29528);
or UO_3277 (O_3277,N_29077,N_29374);
and UO_3278 (O_3278,N_29574,N_29237);
nand UO_3279 (O_3279,N_29966,N_29530);
nand UO_3280 (O_3280,N_29850,N_29239);
and UO_3281 (O_3281,N_29598,N_29293);
nor UO_3282 (O_3282,N_29700,N_29362);
nor UO_3283 (O_3283,N_29528,N_29970);
nand UO_3284 (O_3284,N_29095,N_29617);
or UO_3285 (O_3285,N_29644,N_29955);
nor UO_3286 (O_3286,N_29835,N_29020);
and UO_3287 (O_3287,N_29502,N_29629);
and UO_3288 (O_3288,N_29842,N_29293);
nand UO_3289 (O_3289,N_29442,N_29973);
xor UO_3290 (O_3290,N_29287,N_29607);
xnor UO_3291 (O_3291,N_29279,N_29515);
xnor UO_3292 (O_3292,N_29900,N_29501);
or UO_3293 (O_3293,N_29189,N_29515);
nor UO_3294 (O_3294,N_29849,N_29952);
nor UO_3295 (O_3295,N_29581,N_29850);
nor UO_3296 (O_3296,N_29186,N_29534);
nand UO_3297 (O_3297,N_29677,N_29162);
xor UO_3298 (O_3298,N_29978,N_29012);
xor UO_3299 (O_3299,N_29686,N_29567);
nand UO_3300 (O_3300,N_29092,N_29182);
or UO_3301 (O_3301,N_29309,N_29140);
xnor UO_3302 (O_3302,N_29754,N_29972);
nand UO_3303 (O_3303,N_29536,N_29766);
nand UO_3304 (O_3304,N_29943,N_29799);
or UO_3305 (O_3305,N_29937,N_29714);
xor UO_3306 (O_3306,N_29163,N_29571);
nor UO_3307 (O_3307,N_29387,N_29719);
and UO_3308 (O_3308,N_29084,N_29634);
nand UO_3309 (O_3309,N_29515,N_29137);
nand UO_3310 (O_3310,N_29456,N_29520);
and UO_3311 (O_3311,N_29149,N_29363);
nand UO_3312 (O_3312,N_29082,N_29097);
xor UO_3313 (O_3313,N_29253,N_29653);
or UO_3314 (O_3314,N_29872,N_29128);
xor UO_3315 (O_3315,N_29260,N_29762);
nand UO_3316 (O_3316,N_29389,N_29855);
xnor UO_3317 (O_3317,N_29822,N_29624);
xor UO_3318 (O_3318,N_29210,N_29976);
nor UO_3319 (O_3319,N_29512,N_29579);
and UO_3320 (O_3320,N_29431,N_29823);
and UO_3321 (O_3321,N_29845,N_29120);
nand UO_3322 (O_3322,N_29196,N_29482);
or UO_3323 (O_3323,N_29439,N_29205);
nor UO_3324 (O_3324,N_29334,N_29228);
xor UO_3325 (O_3325,N_29724,N_29663);
nand UO_3326 (O_3326,N_29510,N_29990);
and UO_3327 (O_3327,N_29819,N_29601);
nor UO_3328 (O_3328,N_29207,N_29804);
nand UO_3329 (O_3329,N_29041,N_29921);
and UO_3330 (O_3330,N_29257,N_29765);
and UO_3331 (O_3331,N_29010,N_29853);
nor UO_3332 (O_3332,N_29728,N_29617);
nor UO_3333 (O_3333,N_29032,N_29758);
nor UO_3334 (O_3334,N_29838,N_29998);
or UO_3335 (O_3335,N_29068,N_29601);
xnor UO_3336 (O_3336,N_29150,N_29232);
or UO_3337 (O_3337,N_29074,N_29088);
xnor UO_3338 (O_3338,N_29452,N_29875);
or UO_3339 (O_3339,N_29918,N_29885);
or UO_3340 (O_3340,N_29624,N_29558);
nor UO_3341 (O_3341,N_29305,N_29953);
and UO_3342 (O_3342,N_29575,N_29807);
and UO_3343 (O_3343,N_29897,N_29456);
nand UO_3344 (O_3344,N_29130,N_29839);
nand UO_3345 (O_3345,N_29484,N_29472);
and UO_3346 (O_3346,N_29023,N_29738);
or UO_3347 (O_3347,N_29029,N_29422);
and UO_3348 (O_3348,N_29299,N_29309);
nor UO_3349 (O_3349,N_29357,N_29424);
nor UO_3350 (O_3350,N_29212,N_29136);
or UO_3351 (O_3351,N_29399,N_29080);
and UO_3352 (O_3352,N_29596,N_29573);
or UO_3353 (O_3353,N_29351,N_29774);
xnor UO_3354 (O_3354,N_29717,N_29748);
and UO_3355 (O_3355,N_29448,N_29446);
xnor UO_3356 (O_3356,N_29804,N_29733);
or UO_3357 (O_3357,N_29329,N_29566);
nor UO_3358 (O_3358,N_29485,N_29657);
or UO_3359 (O_3359,N_29770,N_29567);
and UO_3360 (O_3360,N_29877,N_29775);
and UO_3361 (O_3361,N_29601,N_29022);
nor UO_3362 (O_3362,N_29189,N_29479);
and UO_3363 (O_3363,N_29473,N_29185);
and UO_3364 (O_3364,N_29450,N_29647);
or UO_3365 (O_3365,N_29611,N_29109);
and UO_3366 (O_3366,N_29261,N_29244);
and UO_3367 (O_3367,N_29539,N_29910);
nand UO_3368 (O_3368,N_29828,N_29865);
and UO_3369 (O_3369,N_29480,N_29011);
xnor UO_3370 (O_3370,N_29622,N_29553);
nor UO_3371 (O_3371,N_29434,N_29149);
xor UO_3372 (O_3372,N_29835,N_29091);
nor UO_3373 (O_3373,N_29342,N_29301);
nand UO_3374 (O_3374,N_29197,N_29786);
and UO_3375 (O_3375,N_29986,N_29201);
and UO_3376 (O_3376,N_29742,N_29989);
xnor UO_3377 (O_3377,N_29187,N_29781);
and UO_3378 (O_3378,N_29098,N_29745);
or UO_3379 (O_3379,N_29360,N_29849);
xnor UO_3380 (O_3380,N_29476,N_29050);
or UO_3381 (O_3381,N_29980,N_29471);
and UO_3382 (O_3382,N_29742,N_29047);
and UO_3383 (O_3383,N_29735,N_29777);
nand UO_3384 (O_3384,N_29859,N_29318);
and UO_3385 (O_3385,N_29686,N_29302);
nand UO_3386 (O_3386,N_29643,N_29639);
xor UO_3387 (O_3387,N_29769,N_29585);
or UO_3388 (O_3388,N_29048,N_29694);
and UO_3389 (O_3389,N_29719,N_29769);
and UO_3390 (O_3390,N_29172,N_29087);
xnor UO_3391 (O_3391,N_29459,N_29088);
xor UO_3392 (O_3392,N_29252,N_29824);
nand UO_3393 (O_3393,N_29496,N_29533);
nand UO_3394 (O_3394,N_29056,N_29658);
and UO_3395 (O_3395,N_29226,N_29775);
nor UO_3396 (O_3396,N_29015,N_29457);
xor UO_3397 (O_3397,N_29019,N_29570);
nand UO_3398 (O_3398,N_29379,N_29828);
and UO_3399 (O_3399,N_29234,N_29985);
and UO_3400 (O_3400,N_29199,N_29924);
and UO_3401 (O_3401,N_29501,N_29292);
nand UO_3402 (O_3402,N_29606,N_29403);
and UO_3403 (O_3403,N_29944,N_29857);
or UO_3404 (O_3404,N_29396,N_29069);
and UO_3405 (O_3405,N_29404,N_29274);
xor UO_3406 (O_3406,N_29802,N_29251);
xor UO_3407 (O_3407,N_29473,N_29595);
nand UO_3408 (O_3408,N_29005,N_29414);
or UO_3409 (O_3409,N_29613,N_29484);
or UO_3410 (O_3410,N_29053,N_29722);
and UO_3411 (O_3411,N_29916,N_29633);
xor UO_3412 (O_3412,N_29481,N_29618);
nand UO_3413 (O_3413,N_29125,N_29382);
xor UO_3414 (O_3414,N_29692,N_29936);
and UO_3415 (O_3415,N_29884,N_29276);
nand UO_3416 (O_3416,N_29608,N_29602);
and UO_3417 (O_3417,N_29156,N_29901);
and UO_3418 (O_3418,N_29002,N_29158);
and UO_3419 (O_3419,N_29566,N_29890);
xnor UO_3420 (O_3420,N_29204,N_29386);
or UO_3421 (O_3421,N_29464,N_29564);
and UO_3422 (O_3422,N_29337,N_29355);
nor UO_3423 (O_3423,N_29142,N_29198);
and UO_3424 (O_3424,N_29817,N_29567);
nor UO_3425 (O_3425,N_29515,N_29181);
nand UO_3426 (O_3426,N_29618,N_29074);
xor UO_3427 (O_3427,N_29693,N_29254);
and UO_3428 (O_3428,N_29381,N_29683);
nand UO_3429 (O_3429,N_29428,N_29953);
xor UO_3430 (O_3430,N_29694,N_29663);
or UO_3431 (O_3431,N_29038,N_29767);
nand UO_3432 (O_3432,N_29093,N_29879);
xor UO_3433 (O_3433,N_29995,N_29368);
nor UO_3434 (O_3434,N_29235,N_29721);
xor UO_3435 (O_3435,N_29269,N_29426);
nor UO_3436 (O_3436,N_29974,N_29022);
nand UO_3437 (O_3437,N_29542,N_29197);
or UO_3438 (O_3438,N_29464,N_29934);
and UO_3439 (O_3439,N_29264,N_29980);
nor UO_3440 (O_3440,N_29082,N_29239);
or UO_3441 (O_3441,N_29840,N_29321);
and UO_3442 (O_3442,N_29390,N_29372);
nor UO_3443 (O_3443,N_29385,N_29249);
nand UO_3444 (O_3444,N_29149,N_29715);
nand UO_3445 (O_3445,N_29773,N_29354);
nor UO_3446 (O_3446,N_29456,N_29706);
nor UO_3447 (O_3447,N_29269,N_29748);
nor UO_3448 (O_3448,N_29932,N_29081);
nor UO_3449 (O_3449,N_29520,N_29049);
and UO_3450 (O_3450,N_29484,N_29578);
nand UO_3451 (O_3451,N_29459,N_29242);
nand UO_3452 (O_3452,N_29524,N_29878);
xnor UO_3453 (O_3453,N_29649,N_29048);
nand UO_3454 (O_3454,N_29556,N_29466);
and UO_3455 (O_3455,N_29089,N_29400);
or UO_3456 (O_3456,N_29033,N_29751);
nor UO_3457 (O_3457,N_29763,N_29701);
or UO_3458 (O_3458,N_29323,N_29502);
nor UO_3459 (O_3459,N_29859,N_29874);
xnor UO_3460 (O_3460,N_29437,N_29030);
or UO_3461 (O_3461,N_29694,N_29661);
or UO_3462 (O_3462,N_29890,N_29046);
nor UO_3463 (O_3463,N_29722,N_29440);
nor UO_3464 (O_3464,N_29798,N_29800);
nor UO_3465 (O_3465,N_29800,N_29144);
and UO_3466 (O_3466,N_29151,N_29402);
nor UO_3467 (O_3467,N_29940,N_29591);
and UO_3468 (O_3468,N_29327,N_29603);
nand UO_3469 (O_3469,N_29097,N_29454);
nor UO_3470 (O_3470,N_29906,N_29843);
nand UO_3471 (O_3471,N_29077,N_29899);
nand UO_3472 (O_3472,N_29612,N_29368);
or UO_3473 (O_3473,N_29830,N_29293);
xnor UO_3474 (O_3474,N_29882,N_29800);
nor UO_3475 (O_3475,N_29426,N_29881);
nor UO_3476 (O_3476,N_29751,N_29872);
nor UO_3477 (O_3477,N_29107,N_29280);
nor UO_3478 (O_3478,N_29001,N_29949);
nor UO_3479 (O_3479,N_29430,N_29222);
xnor UO_3480 (O_3480,N_29110,N_29341);
xor UO_3481 (O_3481,N_29739,N_29750);
nor UO_3482 (O_3482,N_29075,N_29767);
and UO_3483 (O_3483,N_29330,N_29178);
nor UO_3484 (O_3484,N_29141,N_29103);
and UO_3485 (O_3485,N_29965,N_29705);
and UO_3486 (O_3486,N_29627,N_29941);
xnor UO_3487 (O_3487,N_29340,N_29665);
nand UO_3488 (O_3488,N_29852,N_29910);
and UO_3489 (O_3489,N_29223,N_29669);
xnor UO_3490 (O_3490,N_29076,N_29810);
xor UO_3491 (O_3491,N_29516,N_29437);
or UO_3492 (O_3492,N_29141,N_29479);
nand UO_3493 (O_3493,N_29830,N_29021);
nand UO_3494 (O_3494,N_29145,N_29732);
or UO_3495 (O_3495,N_29167,N_29675);
xnor UO_3496 (O_3496,N_29303,N_29244);
and UO_3497 (O_3497,N_29628,N_29158);
nor UO_3498 (O_3498,N_29529,N_29222);
xor UO_3499 (O_3499,N_29190,N_29800);
endmodule