module basic_500_3000_500_6_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_37,In_187);
and U1 (N_1,In_462,In_138);
or U2 (N_2,In_381,In_130);
nor U3 (N_3,In_109,In_283);
nor U4 (N_4,In_95,In_90);
nand U5 (N_5,In_239,In_326);
nand U6 (N_6,In_473,In_20);
and U7 (N_7,In_420,In_416);
or U8 (N_8,In_364,In_98);
and U9 (N_9,In_447,In_267);
nor U10 (N_10,In_202,In_218);
or U11 (N_11,In_278,In_212);
and U12 (N_12,In_241,In_96);
xor U13 (N_13,In_0,In_105);
and U14 (N_14,In_397,In_426);
nor U15 (N_15,In_336,In_143);
xor U16 (N_16,In_262,In_357);
and U17 (N_17,In_128,In_348);
or U18 (N_18,In_135,In_404);
nor U19 (N_19,In_53,In_162);
or U20 (N_20,In_340,In_117);
and U21 (N_21,In_395,In_131);
and U22 (N_22,In_303,In_298);
nand U23 (N_23,In_295,In_172);
nor U24 (N_24,In_484,In_42);
or U25 (N_25,In_479,In_240);
nand U26 (N_26,In_290,In_341);
and U27 (N_27,In_101,In_358);
or U28 (N_28,In_166,In_398);
and U29 (N_29,In_246,In_31);
or U30 (N_30,In_439,In_39);
nand U31 (N_31,In_294,In_17);
nor U32 (N_32,In_275,In_235);
or U33 (N_33,In_476,In_459);
nand U34 (N_34,In_421,In_427);
nor U35 (N_35,In_45,In_26);
xor U36 (N_36,In_180,In_111);
and U37 (N_37,In_141,In_145);
or U38 (N_38,In_6,In_50);
and U39 (N_39,In_441,In_196);
nand U40 (N_40,In_237,In_8);
or U41 (N_41,In_337,In_440);
or U42 (N_42,In_7,In_207);
and U43 (N_43,In_216,In_300);
and U44 (N_44,In_149,In_322);
nor U45 (N_45,In_64,In_346);
and U46 (N_46,In_169,In_311);
nor U47 (N_47,In_82,In_81);
and U48 (N_48,In_119,In_460);
or U49 (N_49,In_274,In_467);
and U50 (N_50,In_469,In_38);
and U51 (N_51,In_52,In_120);
nand U52 (N_52,In_386,In_270);
or U53 (N_53,In_59,In_384);
nand U54 (N_54,In_150,In_254);
or U55 (N_55,In_279,In_214);
and U56 (N_56,In_123,In_151);
nand U57 (N_57,In_265,In_10);
xnor U58 (N_58,In_253,In_181);
or U59 (N_59,In_297,In_104);
and U60 (N_60,In_134,In_291);
or U61 (N_61,In_174,In_312);
nor U62 (N_62,In_137,In_284);
nor U63 (N_63,In_32,In_425);
and U64 (N_64,In_259,In_107);
and U65 (N_65,In_478,In_227);
nand U66 (N_66,In_142,In_195);
and U67 (N_67,In_88,In_489);
or U68 (N_68,In_179,In_176);
nand U69 (N_69,In_448,In_412);
nor U70 (N_70,In_83,In_2);
and U71 (N_71,In_354,In_175);
and U72 (N_72,In_375,In_446);
and U73 (N_73,In_18,In_156);
nor U74 (N_74,In_62,In_490);
nor U75 (N_75,In_238,In_126);
nand U76 (N_76,In_436,In_451);
and U77 (N_77,In_79,In_396);
and U78 (N_78,In_315,In_407);
nor U79 (N_79,In_417,In_268);
nand U80 (N_80,In_68,In_296);
or U81 (N_81,In_173,In_338);
nand U82 (N_82,In_261,In_276);
or U83 (N_83,In_465,In_273);
nor U84 (N_84,In_380,In_220);
nand U85 (N_85,In_61,In_51);
nand U86 (N_86,In_71,In_406);
nand U87 (N_87,In_122,In_411);
nor U88 (N_88,In_112,In_229);
or U89 (N_89,In_167,In_301);
or U90 (N_90,In_495,In_3);
or U91 (N_91,In_219,In_30);
nand U92 (N_92,In_60,In_497);
or U93 (N_93,In_438,In_80);
nor U94 (N_94,In_182,In_194);
and U95 (N_95,In_49,In_46);
nand U96 (N_96,In_387,In_103);
nor U97 (N_97,In_333,In_247);
and U98 (N_98,In_217,In_74);
nand U99 (N_99,In_23,In_437);
or U100 (N_100,In_472,In_189);
nor U101 (N_101,In_255,In_76);
nand U102 (N_102,In_245,In_370);
nor U103 (N_103,In_385,In_309);
nor U104 (N_104,In_21,In_486);
nor U105 (N_105,In_153,In_363);
and U106 (N_106,In_266,In_400);
nor U107 (N_107,In_299,In_402);
nand U108 (N_108,In_445,In_328);
nor U109 (N_109,In_342,In_54);
nand U110 (N_110,In_356,In_263);
xnor U111 (N_111,In_443,In_100);
nand U112 (N_112,In_133,In_75);
nand U113 (N_113,In_1,In_429);
nor U114 (N_114,In_92,In_331);
nand U115 (N_115,In_292,In_77);
xor U116 (N_116,In_376,In_147);
and U117 (N_117,In_391,In_413);
or U118 (N_118,In_35,In_401);
or U119 (N_119,In_230,In_491);
nor U120 (N_120,In_178,In_482);
and U121 (N_121,In_91,In_316);
nor U122 (N_122,In_22,In_428);
or U123 (N_123,In_118,In_457);
nor U124 (N_124,In_410,In_474);
and U125 (N_125,In_223,In_488);
nor U126 (N_126,In_125,In_372);
nand U127 (N_127,In_409,In_414);
nor U128 (N_128,In_127,In_197);
nor U129 (N_129,In_305,In_66);
nor U130 (N_130,In_158,In_392);
xor U131 (N_131,In_163,In_164);
or U132 (N_132,In_63,In_4);
nor U133 (N_133,In_444,In_466);
and U134 (N_134,In_29,In_69);
nor U135 (N_135,In_224,In_67);
or U136 (N_136,In_25,In_302);
and U137 (N_137,In_190,In_165);
and U138 (N_138,In_377,In_359);
nor U139 (N_139,In_14,In_424);
nand U140 (N_140,In_121,In_132);
or U141 (N_141,In_144,In_277);
or U142 (N_142,In_499,In_85);
and U143 (N_143,In_360,In_399);
nor U144 (N_144,In_204,In_403);
nor U145 (N_145,In_361,In_226);
or U146 (N_146,In_373,In_192);
or U147 (N_147,In_41,In_99);
nor U148 (N_148,In_168,In_324);
or U149 (N_149,In_36,In_345);
nor U150 (N_150,In_113,In_293);
and U151 (N_151,In_55,In_350);
nor U152 (N_152,In_244,In_5);
nand U153 (N_153,In_199,In_250);
and U154 (N_154,In_355,In_222);
and U155 (N_155,In_487,In_269);
nand U156 (N_156,In_256,In_191);
nor U157 (N_157,In_308,In_264);
nor U158 (N_158,In_282,In_366);
or U159 (N_159,In_12,In_468);
or U160 (N_160,In_110,In_87);
or U161 (N_161,In_48,In_464);
or U162 (N_162,In_236,In_200);
and U163 (N_163,In_86,In_215);
and U164 (N_164,In_475,In_435);
nand U165 (N_165,In_494,In_24);
nor U166 (N_166,In_430,In_347);
and U167 (N_167,In_492,In_188);
and U168 (N_168,In_160,In_232);
and U169 (N_169,In_442,In_323);
nand U170 (N_170,In_458,In_433);
or U171 (N_171,In_184,In_390);
or U172 (N_172,In_234,In_471);
or U173 (N_173,In_139,In_432);
nor U174 (N_174,In_313,In_304);
nor U175 (N_175,In_203,In_28);
and U176 (N_176,In_243,In_454);
nand U177 (N_177,In_453,In_257);
or U178 (N_178,In_288,In_483);
nand U179 (N_179,In_231,In_102);
and U180 (N_180,In_485,In_285);
nand U181 (N_181,In_58,In_78);
nand U182 (N_182,In_70,In_94);
or U183 (N_183,In_44,In_9);
and U184 (N_184,In_198,In_335);
nor U185 (N_185,In_280,In_325);
or U186 (N_186,In_252,In_177);
and U187 (N_187,In_73,In_43);
nor U188 (N_188,In_106,In_154);
and U189 (N_189,In_415,In_205);
or U190 (N_190,In_251,In_260);
or U191 (N_191,In_493,In_463);
or U192 (N_192,In_456,In_431);
or U193 (N_193,In_140,In_171);
nand U194 (N_194,In_378,In_210);
and U195 (N_195,In_33,In_65);
or U196 (N_196,In_16,In_157);
nand U197 (N_197,In_449,In_108);
or U198 (N_198,In_367,In_56);
and U199 (N_199,In_152,In_408);
nand U200 (N_200,In_480,In_344);
and U201 (N_201,In_334,In_159);
nand U202 (N_202,In_146,In_136);
nor U203 (N_203,In_362,In_89);
nand U204 (N_204,In_161,In_374);
nor U205 (N_205,In_40,In_185);
nand U206 (N_206,In_394,In_155);
nor U207 (N_207,In_388,In_317);
or U208 (N_208,In_209,In_19);
nand U209 (N_209,In_319,In_286);
nand U210 (N_210,In_383,In_148);
or U211 (N_211,In_271,In_34);
or U212 (N_212,In_249,In_221);
nor U213 (N_213,In_306,In_393);
nor U214 (N_214,In_477,In_72);
nor U215 (N_215,In_330,In_84);
or U216 (N_216,In_365,In_418);
nand U217 (N_217,In_450,In_201);
nor U218 (N_218,In_186,In_389);
nand U219 (N_219,In_289,In_461);
and U220 (N_220,In_327,In_498);
nand U221 (N_221,In_368,In_272);
or U222 (N_222,In_233,In_452);
or U223 (N_223,In_183,In_206);
nand U224 (N_224,In_332,In_352);
nor U225 (N_225,In_321,In_287);
nand U226 (N_226,In_11,In_15);
nand U227 (N_227,In_343,In_307);
or U228 (N_228,In_314,In_379);
or U229 (N_229,In_349,In_481);
and U230 (N_230,In_351,In_318);
and U231 (N_231,In_129,In_193);
or U232 (N_232,In_434,In_57);
and U233 (N_233,In_422,In_225);
and U234 (N_234,In_496,In_115);
and U235 (N_235,In_423,In_353);
and U236 (N_236,In_242,In_455);
and U237 (N_237,In_419,In_228);
and U238 (N_238,In_258,In_97);
nand U239 (N_239,In_27,In_371);
or U240 (N_240,In_116,In_213);
and U241 (N_241,In_310,In_248);
nor U242 (N_242,In_47,In_211);
and U243 (N_243,In_320,In_329);
or U244 (N_244,In_339,In_124);
and U245 (N_245,In_93,In_13);
nand U246 (N_246,In_170,In_114);
nand U247 (N_247,In_470,In_405);
nand U248 (N_248,In_382,In_281);
nand U249 (N_249,In_208,In_369);
or U250 (N_250,In_102,In_126);
nand U251 (N_251,In_26,In_472);
or U252 (N_252,In_356,In_419);
nand U253 (N_253,In_71,In_60);
nand U254 (N_254,In_183,In_133);
nor U255 (N_255,In_280,In_42);
or U256 (N_256,In_128,In_275);
nand U257 (N_257,In_459,In_408);
nand U258 (N_258,In_51,In_105);
nand U259 (N_259,In_115,In_129);
nor U260 (N_260,In_300,In_103);
and U261 (N_261,In_245,In_206);
or U262 (N_262,In_19,In_4);
nor U263 (N_263,In_99,In_150);
or U264 (N_264,In_51,In_166);
nand U265 (N_265,In_110,In_483);
nor U266 (N_266,In_378,In_182);
or U267 (N_267,In_351,In_230);
or U268 (N_268,In_290,In_89);
nor U269 (N_269,In_189,In_107);
nor U270 (N_270,In_237,In_70);
nand U271 (N_271,In_277,In_384);
or U272 (N_272,In_442,In_266);
or U273 (N_273,In_378,In_322);
and U274 (N_274,In_310,In_466);
or U275 (N_275,In_284,In_51);
nor U276 (N_276,In_159,In_21);
nand U277 (N_277,In_440,In_314);
or U278 (N_278,In_3,In_112);
nor U279 (N_279,In_292,In_436);
nor U280 (N_280,In_260,In_281);
or U281 (N_281,In_415,In_137);
and U282 (N_282,In_49,In_318);
nand U283 (N_283,In_214,In_200);
nor U284 (N_284,In_128,In_319);
or U285 (N_285,In_442,In_33);
nand U286 (N_286,In_287,In_34);
or U287 (N_287,In_88,In_190);
nand U288 (N_288,In_100,In_320);
xor U289 (N_289,In_274,In_260);
nand U290 (N_290,In_14,In_361);
xnor U291 (N_291,In_197,In_496);
nand U292 (N_292,In_366,In_484);
nor U293 (N_293,In_65,In_478);
and U294 (N_294,In_71,In_248);
or U295 (N_295,In_66,In_278);
or U296 (N_296,In_79,In_102);
nor U297 (N_297,In_457,In_119);
or U298 (N_298,In_287,In_8);
nand U299 (N_299,In_324,In_140);
nor U300 (N_300,In_493,In_461);
nand U301 (N_301,In_232,In_148);
or U302 (N_302,In_336,In_53);
nor U303 (N_303,In_24,In_422);
nor U304 (N_304,In_484,In_256);
or U305 (N_305,In_255,In_485);
nor U306 (N_306,In_114,In_37);
nand U307 (N_307,In_305,In_418);
nand U308 (N_308,In_208,In_465);
or U309 (N_309,In_369,In_44);
or U310 (N_310,In_220,In_423);
and U311 (N_311,In_83,In_104);
nor U312 (N_312,In_104,In_400);
or U313 (N_313,In_346,In_369);
nor U314 (N_314,In_306,In_181);
nor U315 (N_315,In_456,In_370);
and U316 (N_316,In_288,In_433);
or U317 (N_317,In_383,In_260);
xnor U318 (N_318,In_340,In_360);
or U319 (N_319,In_378,In_472);
and U320 (N_320,In_340,In_173);
nor U321 (N_321,In_131,In_475);
nand U322 (N_322,In_213,In_353);
nor U323 (N_323,In_194,In_403);
or U324 (N_324,In_18,In_228);
nor U325 (N_325,In_263,In_308);
nand U326 (N_326,In_221,In_325);
and U327 (N_327,In_335,In_138);
nand U328 (N_328,In_249,In_494);
nand U329 (N_329,In_255,In_67);
nand U330 (N_330,In_476,In_142);
nor U331 (N_331,In_491,In_69);
nand U332 (N_332,In_373,In_235);
nand U333 (N_333,In_320,In_459);
or U334 (N_334,In_419,In_454);
nor U335 (N_335,In_96,In_297);
or U336 (N_336,In_260,In_486);
and U337 (N_337,In_79,In_6);
nor U338 (N_338,In_60,In_436);
and U339 (N_339,In_245,In_328);
nand U340 (N_340,In_153,In_63);
nand U341 (N_341,In_249,In_171);
nand U342 (N_342,In_110,In_153);
nand U343 (N_343,In_367,In_374);
nor U344 (N_344,In_250,In_291);
nand U345 (N_345,In_318,In_93);
or U346 (N_346,In_225,In_18);
nor U347 (N_347,In_316,In_269);
or U348 (N_348,In_290,In_356);
and U349 (N_349,In_143,In_30);
xnor U350 (N_350,In_203,In_101);
nand U351 (N_351,In_195,In_242);
nand U352 (N_352,In_300,In_423);
nand U353 (N_353,In_75,In_95);
nor U354 (N_354,In_434,In_367);
or U355 (N_355,In_482,In_140);
nand U356 (N_356,In_413,In_378);
or U357 (N_357,In_38,In_146);
nand U358 (N_358,In_105,In_346);
nand U359 (N_359,In_61,In_9);
nor U360 (N_360,In_381,In_193);
or U361 (N_361,In_150,In_1);
or U362 (N_362,In_89,In_33);
or U363 (N_363,In_195,In_345);
nor U364 (N_364,In_307,In_397);
or U365 (N_365,In_229,In_80);
nor U366 (N_366,In_364,In_69);
nand U367 (N_367,In_209,In_149);
nand U368 (N_368,In_312,In_367);
nand U369 (N_369,In_240,In_443);
nor U370 (N_370,In_320,In_120);
nand U371 (N_371,In_125,In_185);
or U372 (N_372,In_479,In_111);
or U373 (N_373,In_442,In_316);
nand U374 (N_374,In_474,In_360);
or U375 (N_375,In_219,In_295);
and U376 (N_376,In_6,In_461);
nor U377 (N_377,In_5,In_353);
or U378 (N_378,In_67,In_385);
and U379 (N_379,In_110,In_280);
nor U380 (N_380,In_283,In_226);
nand U381 (N_381,In_302,In_75);
nor U382 (N_382,In_369,In_81);
and U383 (N_383,In_109,In_121);
nand U384 (N_384,In_353,In_6);
and U385 (N_385,In_328,In_87);
nor U386 (N_386,In_371,In_243);
and U387 (N_387,In_96,In_294);
or U388 (N_388,In_78,In_95);
nor U389 (N_389,In_58,In_39);
and U390 (N_390,In_5,In_381);
and U391 (N_391,In_434,In_216);
xnor U392 (N_392,In_25,In_345);
or U393 (N_393,In_301,In_273);
nand U394 (N_394,In_270,In_60);
nor U395 (N_395,In_241,In_175);
nand U396 (N_396,In_298,In_376);
nor U397 (N_397,In_355,In_147);
nor U398 (N_398,In_427,In_48);
nand U399 (N_399,In_284,In_300);
nor U400 (N_400,In_236,In_86);
and U401 (N_401,In_177,In_462);
nand U402 (N_402,In_482,In_197);
xnor U403 (N_403,In_135,In_266);
and U404 (N_404,In_237,In_125);
nand U405 (N_405,In_347,In_441);
or U406 (N_406,In_60,In_344);
and U407 (N_407,In_278,In_218);
nor U408 (N_408,In_307,In_252);
nand U409 (N_409,In_354,In_222);
xor U410 (N_410,In_471,In_185);
nand U411 (N_411,In_380,In_280);
or U412 (N_412,In_195,In_316);
nand U413 (N_413,In_85,In_122);
and U414 (N_414,In_311,In_352);
and U415 (N_415,In_57,In_42);
nand U416 (N_416,In_79,In_224);
nor U417 (N_417,In_110,In_459);
and U418 (N_418,In_220,In_169);
nand U419 (N_419,In_133,In_121);
or U420 (N_420,In_378,In_441);
nand U421 (N_421,In_445,In_19);
or U422 (N_422,In_238,In_17);
or U423 (N_423,In_363,In_27);
nand U424 (N_424,In_172,In_487);
xor U425 (N_425,In_217,In_331);
or U426 (N_426,In_235,In_394);
and U427 (N_427,In_44,In_262);
xor U428 (N_428,In_134,In_216);
or U429 (N_429,In_191,In_116);
and U430 (N_430,In_393,In_36);
and U431 (N_431,In_335,In_471);
and U432 (N_432,In_111,In_423);
nor U433 (N_433,In_52,In_34);
nand U434 (N_434,In_407,In_392);
or U435 (N_435,In_338,In_179);
and U436 (N_436,In_439,In_226);
xnor U437 (N_437,In_256,In_401);
nand U438 (N_438,In_302,In_419);
nand U439 (N_439,In_73,In_364);
nand U440 (N_440,In_144,In_261);
xor U441 (N_441,In_327,In_89);
nand U442 (N_442,In_340,In_311);
nand U443 (N_443,In_123,In_0);
or U444 (N_444,In_291,In_12);
and U445 (N_445,In_382,In_22);
or U446 (N_446,In_255,In_269);
nand U447 (N_447,In_45,In_18);
nand U448 (N_448,In_378,In_81);
nor U449 (N_449,In_392,In_33);
nor U450 (N_450,In_208,In_187);
nand U451 (N_451,In_43,In_357);
and U452 (N_452,In_159,In_341);
and U453 (N_453,In_299,In_389);
and U454 (N_454,In_424,In_259);
and U455 (N_455,In_305,In_198);
nand U456 (N_456,In_212,In_385);
or U457 (N_457,In_32,In_28);
nor U458 (N_458,In_97,In_64);
or U459 (N_459,In_327,In_491);
nor U460 (N_460,In_369,In_116);
nand U461 (N_461,In_345,In_10);
and U462 (N_462,In_312,In_206);
or U463 (N_463,In_195,In_441);
or U464 (N_464,In_115,In_371);
or U465 (N_465,In_353,In_419);
nand U466 (N_466,In_427,In_236);
and U467 (N_467,In_350,In_248);
nand U468 (N_468,In_342,In_429);
or U469 (N_469,In_349,In_106);
nor U470 (N_470,In_467,In_153);
or U471 (N_471,In_298,In_194);
or U472 (N_472,In_217,In_390);
or U473 (N_473,In_299,In_353);
or U474 (N_474,In_404,In_24);
nor U475 (N_475,In_432,In_71);
nand U476 (N_476,In_213,In_99);
nand U477 (N_477,In_232,In_498);
nor U478 (N_478,In_140,In_158);
and U479 (N_479,In_35,In_122);
or U480 (N_480,In_436,In_299);
nand U481 (N_481,In_426,In_384);
nand U482 (N_482,In_469,In_447);
nor U483 (N_483,In_188,In_311);
nand U484 (N_484,In_366,In_451);
or U485 (N_485,In_318,In_347);
nand U486 (N_486,In_214,In_54);
or U487 (N_487,In_11,In_258);
or U488 (N_488,In_196,In_382);
and U489 (N_489,In_389,In_319);
nand U490 (N_490,In_242,In_114);
and U491 (N_491,In_263,In_344);
nor U492 (N_492,In_185,In_5);
or U493 (N_493,In_13,In_267);
nor U494 (N_494,In_281,In_177);
and U495 (N_495,In_436,In_70);
and U496 (N_496,In_475,In_484);
or U497 (N_497,In_427,In_142);
nand U498 (N_498,In_116,In_89);
or U499 (N_499,In_406,In_282);
nand U500 (N_500,N_107,N_257);
nor U501 (N_501,N_279,N_209);
or U502 (N_502,N_317,N_97);
and U503 (N_503,N_134,N_73);
nor U504 (N_504,N_408,N_241);
and U505 (N_505,N_150,N_264);
nand U506 (N_506,N_68,N_113);
nand U507 (N_507,N_219,N_263);
nor U508 (N_508,N_410,N_136);
and U509 (N_509,N_67,N_230);
or U510 (N_510,N_470,N_424);
nand U511 (N_511,N_80,N_307);
or U512 (N_512,N_192,N_425);
xnor U513 (N_513,N_320,N_308);
nor U514 (N_514,N_315,N_297);
and U515 (N_515,N_208,N_288);
nand U516 (N_516,N_329,N_350);
or U517 (N_517,N_0,N_343);
and U518 (N_518,N_498,N_409);
xnor U519 (N_519,N_205,N_149);
or U520 (N_520,N_194,N_490);
nand U521 (N_521,N_277,N_471);
nor U522 (N_522,N_49,N_405);
and U523 (N_523,N_316,N_265);
nand U524 (N_524,N_167,N_383);
nand U525 (N_525,N_162,N_413);
nor U526 (N_526,N_355,N_132);
and U527 (N_527,N_457,N_300);
nor U528 (N_528,N_353,N_301);
nand U529 (N_529,N_431,N_43);
nor U530 (N_530,N_414,N_261);
nand U531 (N_531,N_191,N_356);
or U532 (N_532,N_156,N_10);
nand U533 (N_533,N_227,N_47);
nor U534 (N_534,N_337,N_294);
nor U535 (N_535,N_17,N_369);
nand U536 (N_536,N_181,N_296);
xor U537 (N_537,N_114,N_63);
nand U538 (N_538,N_90,N_333);
nor U539 (N_539,N_22,N_217);
and U540 (N_540,N_18,N_218);
nand U541 (N_541,N_228,N_171);
nand U542 (N_542,N_488,N_469);
nand U543 (N_543,N_378,N_165);
or U544 (N_544,N_478,N_458);
or U545 (N_545,N_441,N_210);
nor U546 (N_546,N_324,N_185);
nor U547 (N_547,N_422,N_313);
nand U548 (N_548,N_411,N_276);
nor U549 (N_549,N_286,N_254);
nand U550 (N_550,N_95,N_161);
or U551 (N_551,N_399,N_499);
or U552 (N_552,N_1,N_388);
nand U553 (N_553,N_391,N_119);
and U554 (N_554,N_60,N_474);
nand U555 (N_555,N_14,N_323);
nor U556 (N_556,N_236,N_403);
nand U557 (N_557,N_66,N_332);
xnor U558 (N_558,N_328,N_271);
or U559 (N_559,N_137,N_222);
and U560 (N_560,N_312,N_131);
and U561 (N_561,N_4,N_238);
nand U562 (N_562,N_443,N_120);
and U563 (N_563,N_168,N_292);
or U564 (N_564,N_34,N_445);
nor U565 (N_565,N_75,N_448);
nor U566 (N_566,N_489,N_198);
nor U567 (N_567,N_148,N_269);
or U568 (N_568,N_495,N_394);
or U569 (N_569,N_78,N_253);
or U570 (N_570,N_237,N_273);
or U571 (N_571,N_460,N_121);
xnor U572 (N_572,N_486,N_89);
and U573 (N_573,N_59,N_325);
or U574 (N_574,N_64,N_427);
or U575 (N_575,N_406,N_81);
or U576 (N_576,N_494,N_289);
nand U577 (N_577,N_311,N_177);
or U578 (N_578,N_466,N_157);
nor U579 (N_579,N_326,N_340);
and U580 (N_580,N_147,N_415);
nor U581 (N_581,N_418,N_44);
nor U582 (N_582,N_246,N_429);
nand U583 (N_583,N_461,N_46);
nand U584 (N_584,N_366,N_215);
and U585 (N_585,N_373,N_39);
nor U586 (N_586,N_176,N_154);
nand U587 (N_587,N_491,N_25);
nand U588 (N_588,N_472,N_235);
nor U589 (N_589,N_272,N_480);
and U590 (N_590,N_145,N_188);
nor U591 (N_591,N_248,N_184);
nor U592 (N_592,N_281,N_464);
nor U593 (N_593,N_314,N_493);
nand U594 (N_594,N_193,N_396);
nor U595 (N_595,N_23,N_242);
and U596 (N_596,N_36,N_249);
or U597 (N_597,N_335,N_50);
and U598 (N_598,N_224,N_117);
nor U599 (N_599,N_30,N_166);
and U600 (N_600,N_104,N_20);
and U601 (N_601,N_140,N_99);
or U602 (N_602,N_196,N_432);
xnor U603 (N_603,N_342,N_155);
and U604 (N_604,N_267,N_13);
xnor U605 (N_605,N_250,N_372);
nor U606 (N_606,N_344,N_33);
and U607 (N_607,N_86,N_213);
nor U608 (N_608,N_361,N_293);
nor U609 (N_609,N_65,N_479);
or U610 (N_610,N_153,N_82);
and U611 (N_611,N_142,N_375);
and U612 (N_612,N_357,N_7);
or U613 (N_613,N_363,N_280);
nor U614 (N_614,N_42,N_275);
nand U615 (N_615,N_346,N_69);
or U616 (N_616,N_310,N_27);
and U617 (N_617,N_182,N_359);
and U618 (N_618,N_212,N_12);
and U619 (N_619,N_256,N_306);
nor U620 (N_620,N_92,N_303);
and U621 (N_621,N_94,N_169);
and U622 (N_622,N_106,N_260);
nand U623 (N_623,N_282,N_226);
nand U624 (N_624,N_477,N_206);
nor U625 (N_625,N_473,N_115);
or U626 (N_626,N_216,N_362);
nor U627 (N_627,N_144,N_365);
or U628 (N_628,N_62,N_348);
nor U629 (N_629,N_183,N_243);
or U630 (N_630,N_164,N_118);
or U631 (N_631,N_354,N_291);
or U632 (N_632,N_225,N_455);
nand U633 (N_633,N_393,N_245);
and U634 (N_634,N_103,N_454);
or U635 (N_635,N_453,N_298);
and U636 (N_636,N_108,N_255);
or U637 (N_637,N_72,N_52);
nand U638 (N_638,N_270,N_266);
or U639 (N_639,N_6,N_28);
and U640 (N_640,N_347,N_70);
or U641 (N_641,N_51,N_24);
and U642 (N_642,N_331,N_349);
or U643 (N_643,N_160,N_274);
nand U644 (N_644,N_201,N_122);
nand U645 (N_645,N_133,N_109);
or U646 (N_646,N_377,N_38);
or U647 (N_647,N_233,N_26);
and U648 (N_648,N_85,N_345);
and U649 (N_649,N_3,N_364);
xor U650 (N_650,N_139,N_98);
or U651 (N_651,N_420,N_387);
and U652 (N_652,N_336,N_295);
nor U653 (N_653,N_305,N_199);
nor U654 (N_654,N_214,N_444);
nand U655 (N_655,N_400,N_35);
and U656 (N_656,N_41,N_417);
nor U657 (N_657,N_385,N_426);
nor U658 (N_658,N_452,N_438);
nor U659 (N_659,N_476,N_423);
and U660 (N_660,N_190,N_111);
and U661 (N_661,N_404,N_371);
nor U662 (N_662,N_382,N_84);
xor U663 (N_663,N_268,N_392);
nand U664 (N_664,N_397,N_492);
or U665 (N_665,N_170,N_462);
nand U666 (N_666,N_220,N_11);
or U667 (N_667,N_302,N_61);
and U668 (N_668,N_287,N_437);
nor U669 (N_669,N_229,N_71);
and U670 (N_670,N_211,N_231);
or U671 (N_671,N_283,N_436);
and U672 (N_672,N_151,N_368);
or U673 (N_673,N_128,N_299);
nand U674 (N_674,N_398,N_76);
nor U675 (N_675,N_126,N_8);
or U676 (N_676,N_401,N_402);
nor U677 (N_677,N_379,N_55);
or U678 (N_678,N_130,N_9);
nor U679 (N_679,N_2,N_58);
and U680 (N_680,N_123,N_407);
nor U681 (N_681,N_322,N_465);
and U682 (N_682,N_386,N_428);
xor U683 (N_683,N_15,N_29);
xnor U684 (N_684,N_32,N_53);
nor U685 (N_685,N_330,N_374);
or U686 (N_686,N_221,N_152);
and U687 (N_687,N_79,N_370);
or U688 (N_688,N_497,N_304);
or U689 (N_689,N_419,N_102);
and U690 (N_690,N_484,N_352);
xnor U691 (N_691,N_251,N_16);
nor U692 (N_692,N_442,N_179);
and U693 (N_693,N_258,N_463);
and U694 (N_694,N_390,N_487);
or U695 (N_695,N_240,N_338);
nand U696 (N_696,N_48,N_434);
xor U697 (N_697,N_31,N_327);
or U698 (N_698,N_376,N_93);
nor U699 (N_699,N_87,N_37);
nand U700 (N_700,N_135,N_321);
or U701 (N_701,N_5,N_449);
nor U702 (N_702,N_389,N_309);
nor U703 (N_703,N_341,N_367);
nor U704 (N_704,N_339,N_189);
and U705 (N_705,N_252,N_483);
or U706 (N_706,N_175,N_232);
nand U707 (N_707,N_440,N_45);
and U708 (N_708,N_239,N_381);
and U709 (N_709,N_360,N_262);
nor U710 (N_710,N_101,N_143);
nor U711 (N_711,N_450,N_163);
nor U712 (N_712,N_96,N_173);
and U713 (N_713,N_412,N_197);
and U714 (N_714,N_112,N_125);
and U715 (N_715,N_204,N_416);
nor U716 (N_716,N_468,N_451);
nor U717 (N_717,N_195,N_172);
nor U718 (N_718,N_247,N_482);
nand U719 (N_719,N_290,N_380);
nor U720 (N_720,N_358,N_447);
nand U721 (N_721,N_57,N_138);
and U722 (N_722,N_202,N_467);
and U723 (N_723,N_278,N_207);
nand U724 (N_724,N_430,N_223);
nand U725 (N_725,N_77,N_384);
nor U726 (N_726,N_116,N_40);
or U727 (N_727,N_475,N_496);
nand U728 (N_728,N_234,N_141);
and U729 (N_729,N_318,N_83);
nor U730 (N_730,N_284,N_439);
nor U731 (N_731,N_456,N_174);
nand U732 (N_732,N_56,N_319);
nand U733 (N_733,N_187,N_180);
nor U734 (N_734,N_459,N_259);
and U735 (N_735,N_351,N_186);
nand U736 (N_736,N_19,N_124);
or U737 (N_737,N_433,N_203);
nor U738 (N_738,N_127,N_395);
and U739 (N_739,N_110,N_74);
nor U740 (N_740,N_105,N_421);
or U741 (N_741,N_91,N_146);
or U742 (N_742,N_129,N_178);
nor U743 (N_743,N_285,N_334);
nor U744 (N_744,N_100,N_244);
nor U745 (N_745,N_481,N_435);
nor U746 (N_746,N_54,N_446);
or U747 (N_747,N_158,N_88);
or U748 (N_748,N_200,N_21);
nand U749 (N_749,N_485,N_159);
and U750 (N_750,N_19,N_391);
or U751 (N_751,N_438,N_105);
nand U752 (N_752,N_229,N_468);
and U753 (N_753,N_59,N_0);
and U754 (N_754,N_45,N_316);
and U755 (N_755,N_344,N_182);
nor U756 (N_756,N_229,N_467);
or U757 (N_757,N_204,N_294);
and U758 (N_758,N_18,N_305);
xor U759 (N_759,N_392,N_166);
xor U760 (N_760,N_163,N_415);
nand U761 (N_761,N_424,N_304);
nand U762 (N_762,N_445,N_204);
nor U763 (N_763,N_95,N_424);
and U764 (N_764,N_25,N_425);
nand U765 (N_765,N_465,N_181);
nor U766 (N_766,N_30,N_214);
or U767 (N_767,N_447,N_110);
nand U768 (N_768,N_441,N_425);
nor U769 (N_769,N_284,N_41);
nand U770 (N_770,N_251,N_235);
nand U771 (N_771,N_363,N_277);
nand U772 (N_772,N_419,N_21);
nand U773 (N_773,N_403,N_45);
and U774 (N_774,N_342,N_159);
and U775 (N_775,N_295,N_243);
or U776 (N_776,N_246,N_152);
nand U777 (N_777,N_292,N_318);
nand U778 (N_778,N_46,N_380);
nor U779 (N_779,N_360,N_6);
nand U780 (N_780,N_223,N_260);
or U781 (N_781,N_366,N_73);
and U782 (N_782,N_343,N_322);
nand U783 (N_783,N_238,N_324);
xnor U784 (N_784,N_146,N_225);
nand U785 (N_785,N_207,N_121);
nor U786 (N_786,N_478,N_287);
nor U787 (N_787,N_437,N_389);
nor U788 (N_788,N_135,N_398);
nor U789 (N_789,N_294,N_423);
nor U790 (N_790,N_105,N_394);
nor U791 (N_791,N_313,N_377);
nand U792 (N_792,N_110,N_238);
and U793 (N_793,N_224,N_11);
or U794 (N_794,N_373,N_268);
nand U795 (N_795,N_59,N_209);
or U796 (N_796,N_205,N_215);
and U797 (N_797,N_155,N_367);
or U798 (N_798,N_167,N_212);
or U799 (N_799,N_10,N_353);
or U800 (N_800,N_490,N_151);
or U801 (N_801,N_161,N_48);
and U802 (N_802,N_204,N_3);
nor U803 (N_803,N_392,N_97);
and U804 (N_804,N_257,N_275);
or U805 (N_805,N_444,N_16);
nor U806 (N_806,N_54,N_496);
nand U807 (N_807,N_16,N_141);
nor U808 (N_808,N_33,N_154);
and U809 (N_809,N_241,N_298);
nand U810 (N_810,N_492,N_454);
nor U811 (N_811,N_188,N_23);
or U812 (N_812,N_236,N_95);
and U813 (N_813,N_148,N_467);
or U814 (N_814,N_61,N_341);
or U815 (N_815,N_411,N_105);
nand U816 (N_816,N_449,N_458);
or U817 (N_817,N_131,N_19);
and U818 (N_818,N_18,N_279);
nor U819 (N_819,N_336,N_76);
nand U820 (N_820,N_431,N_482);
nand U821 (N_821,N_480,N_308);
nand U822 (N_822,N_492,N_85);
and U823 (N_823,N_10,N_450);
or U824 (N_824,N_443,N_387);
nor U825 (N_825,N_472,N_240);
and U826 (N_826,N_205,N_488);
or U827 (N_827,N_59,N_144);
or U828 (N_828,N_367,N_96);
nor U829 (N_829,N_205,N_366);
nand U830 (N_830,N_284,N_440);
or U831 (N_831,N_20,N_118);
or U832 (N_832,N_156,N_41);
and U833 (N_833,N_65,N_158);
xnor U834 (N_834,N_485,N_110);
nand U835 (N_835,N_387,N_200);
or U836 (N_836,N_131,N_30);
nor U837 (N_837,N_272,N_0);
or U838 (N_838,N_388,N_62);
xnor U839 (N_839,N_187,N_436);
xnor U840 (N_840,N_456,N_78);
and U841 (N_841,N_371,N_425);
and U842 (N_842,N_343,N_244);
nor U843 (N_843,N_322,N_493);
and U844 (N_844,N_331,N_435);
nand U845 (N_845,N_300,N_104);
nand U846 (N_846,N_469,N_309);
and U847 (N_847,N_71,N_186);
nor U848 (N_848,N_204,N_44);
nand U849 (N_849,N_191,N_3);
nor U850 (N_850,N_16,N_250);
nor U851 (N_851,N_388,N_2);
nor U852 (N_852,N_198,N_56);
nor U853 (N_853,N_390,N_28);
nand U854 (N_854,N_9,N_428);
or U855 (N_855,N_270,N_141);
nor U856 (N_856,N_85,N_393);
or U857 (N_857,N_171,N_333);
and U858 (N_858,N_474,N_484);
nor U859 (N_859,N_67,N_186);
and U860 (N_860,N_186,N_77);
nor U861 (N_861,N_173,N_467);
nor U862 (N_862,N_347,N_332);
and U863 (N_863,N_15,N_406);
nand U864 (N_864,N_177,N_386);
nor U865 (N_865,N_176,N_280);
nor U866 (N_866,N_65,N_329);
or U867 (N_867,N_485,N_220);
and U868 (N_868,N_16,N_468);
nand U869 (N_869,N_78,N_303);
or U870 (N_870,N_385,N_235);
or U871 (N_871,N_313,N_375);
nor U872 (N_872,N_416,N_159);
xnor U873 (N_873,N_453,N_151);
and U874 (N_874,N_367,N_423);
xor U875 (N_875,N_477,N_161);
xor U876 (N_876,N_448,N_471);
or U877 (N_877,N_415,N_203);
and U878 (N_878,N_256,N_1);
nor U879 (N_879,N_203,N_26);
nor U880 (N_880,N_295,N_479);
nand U881 (N_881,N_342,N_337);
or U882 (N_882,N_194,N_55);
nand U883 (N_883,N_212,N_145);
nand U884 (N_884,N_127,N_295);
or U885 (N_885,N_296,N_333);
or U886 (N_886,N_96,N_487);
and U887 (N_887,N_382,N_243);
or U888 (N_888,N_495,N_308);
and U889 (N_889,N_365,N_496);
nand U890 (N_890,N_37,N_29);
nand U891 (N_891,N_218,N_32);
or U892 (N_892,N_85,N_115);
nand U893 (N_893,N_488,N_310);
and U894 (N_894,N_356,N_180);
and U895 (N_895,N_246,N_331);
nand U896 (N_896,N_496,N_265);
or U897 (N_897,N_48,N_24);
and U898 (N_898,N_485,N_202);
and U899 (N_899,N_489,N_82);
or U900 (N_900,N_453,N_10);
nor U901 (N_901,N_37,N_260);
and U902 (N_902,N_296,N_167);
nor U903 (N_903,N_345,N_191);
nor U904 (N_904,N_252,N_235);
xor U905 (N_905,N_437,N_311);
and U906 (N_906,N_240,N_487);
nand U907 (N_907,N_476,N_216);
nand U908 (N_908,N_339,N_147);
nor U909 (N_909,N_273,N_360);
and U910 (N_910,N_28,N_361);
nor U911 (N_911,N_104,N_18);
or U912 (N_912,N_385,N_369);
or U913 (N_913,N_461,N_275);
nand U914 (N_914,N_340,N_433);
or U915 (N_915,N_484,N_390);
nor U916 (N_916,N_297,N_102);
nand U917 (N_917,N_410,N_113);
and U918 (N_918,N_389,N_294);
and U919 (N_919,N_445,N_366);
or U920 (N_920,N_48,N_236);
and U921 (N_921,N_422,N_10);
nor U922 (N_922,N_46,N_7);
or U923 (N_923,N_66,N_37);
xnor U924 (N_924,N_47,N_48);
and U925 (N_925,N_174,N_131);
nand U926 (N_926,N_190,N_182);
or U927 (N_927,N_324,N_103);
nor U928 (N_928,N_73,N_448);
and U929 (N_929,N_200,N_36);
nor U930 (N_930,N_88,N_13);
nand U931 (N_931,N_207,N_7);
nand U932 (N_932,N_30,N_189);
and U933 (N_933,N_354,N_178);
or U934 (N_934,N_277,N_164);
nand U935 (N_935,N_379,N_73);
or U936 (N_936,N_208,N_30);
nor U937 (N_937,N_215,N_447);
nor U938 (N_938,N_352,N_374);
nor U939 (N_939,N_265,N_115);
nand U940 (N_940,N_19,N_70);
and U941 (N_941,N_390,N_333);
nor U942 (N_942,N_70,N_304);
nor U943 (N_943,N_134,N_298);
nand U944 (N_944,N_218,N_462);
or U945 (N_945,N_30,N_390);
nor U946 (N_946,N_309,N_87);
nor U947 (N_947,N_470,N_449);
or U948 (N_948,N_88,N_101);
nand U949 (N_949,N_273,N_187);
and U950 (N_950,N_484,N_12);
or U951 (N_951,N_484,N_154);
or U952 (N_952,N_466,N_459);
nor U953 (N_953,N_159,N_196);
nor U954 (N_954,N_73,N_477);
or U955 (N_955,N_211,N_281);
xor U956 (N_956,N_483,N_354);
and U957 (N_957,N_456,N_477);
nor U958 (N_958,N_453,N_100);
and U959 (N_959,N_38,N_157);
and U960 (N_960,N_191,N_184);
xnor U961 (N_961,N_418,N_238);
nor U962 (N_962,N_276,N_153);
or U963 (N_963,N_294,N_86);
and U964 (N_964,N_143,N_234);
and U965 (N_965,N_362,N_95);
and U966 (N_966,N_458,N_271);
nand U967 (N_967,N_259,N_238);
nor U968 (N_968,N_71,N_426);
nand U969 (N_969,N_85,N_16);
nor U970 (N_970,N_470,N_62);
nand U971 (N_971,N_146,N_325);
or U972 (N_972,N_281,N_233);
or U973 (N_973,N_137,N_240);
or U974 (N_974,N_474,N_477);
nor U975 (N_975,N_124,N_360);
and U976 (N_976,N_331,N_351);
nor U977 (N_977,N_328,N_129);
nand U978 (N_978,N_145,N_290);
and U979 (N_979,N_491,N_94);
nand U980 (N_980,N_134,N_369);
or U981 (N_981,N_238,N_305);
and U982 (N_982,N_447,N_100);
or U983 (N_983,N_174,N_368);
and U984 (N_984,N_16,N_155);
or U985 (N_985,N_198,N_157);
or U986 (N_986,N_344,N_256);
and U987 (N_987,N_397,N_495);
and U988 (N_988,N_133,N_176);
or U989 (N_989,N_218,N_415);
nor U990 (N_990,N_212,N_357);
nor U991 (N_991,N_335,N_265);
nor U992 (N_992,N_182,N_74);
and U993 (N_993,N_484,N_33);
and U994 (N_994,N_162,N_303);
nor U995 (N_995,N_194,N_25);
and U996 (N_996,N_454,N_89);
nand U997 (N_997,N_245,N_63);
and U998 (N_998,N_344,N_440);
or U999 (N_999,N_135,N_356);
nor U1000 (N_1000,N_636,N_651);
xnor U1001 (N_1001,N_828,N_569);
and U1002 (N_1002,N_504,N_936);
or U1003 (N_1003,N_550,N_744);
or U1004 (N_1004,N_517,N_613);
and U1005 (N_1005,N_638,N_626);
xor U1006 (N_1006,N_601,N_890);
or U1007 (N_1007,N_742,N_657);
nor U1008 (N_1008,N_928,N_854);
or U1009 (N_1009,N_946,N_720);
nand U1010 (N_1010,N_740,N_948);
or U1011 (N_1011,N_749,N_732);
or U1012 (N_1012,N_896,N_977);
nor U1013 (N_1013,N_899,N_993);
nor U1014 (N_1014,N_566,N_759);
xor U1015 (N_1015,N_688,N_888);
or U1016 (N_1016,N_575,N_739);
or U1017 (N_1017,N_653,N_757);
or U1018 (N_1018,N_856,N_881);
nor U1019 (N_1019,N_996,N_608);
or U1020 (N_1020,N_589,N_889);
nand U1021 (N_1021,N_719,N_611);
nor U1022 (N_1022,N_958,N_672);
nor U1023 (N_1023,N_760,N_943);
or U1024 (N_1024,N_844,N_635);
or U1025 (N_1025,N_523,N_603);
nand U1026 (N_1026,N_803,N_598);
or U1027 (N_1027,N_827,N_982);
nor U1028 (N_1028,N_779,N_606);
and U1029 (N_1029,N_585,N_787);
or U1030 (N_1030,N_694,N_634);
nor U1031 (N_1031,N_614,N_780);
and U1032 (N_1032,N_628,N_869);
or U1033 (N_1033,N_750,N_661);
nor U1034 (N_1034,N_766,N_887);
nor U1035 (N_1035,N_870,N_850);
and U1036 (N_1036,N_617,N_811);
nor U1037 (N_1037,N_515,N_913);
nor U1038 (N_1038,N_677,N_519);
nor U1039 (N_1039,N_537,N_902);
or U1040 (N_1040,N_724,N_616);
nor U1041 (N_1041,N_786,N_640);
nand U1042 (N_1042,N_914,N_510);
nor U1043 (N_1043,N_755,N_654);
nand U1044 (N_1044,N_745,N_738);
nand U1045 (N_1045,N_736,N_952);
nor U1046 (N_1046,N_639,N_524);
nand U1047 (N_1047,N_590,N_622);
and U1048 (N_1048,N_637,N_901);
nand U1049 (N_1049,N_935,N_907);
or U1050 (N_1050,N_641,N_705);
nor U1051 (N_1051,N_775,N_772);
nand U1052 (N_1052,N_737,N_885);
nand U1053 (N_1053,N_546,N_602);
and U1054 (N_1054,N_686,N_992);
nand U1055 (N_1055,N_625,N_691);
or U1056 (N_1056,N_893,N_747);
and U1057 (N_1057,N_858,N_554);
nand U1058 (N_1058,N_868,N_607);
nand U1059 (N_1059,N_697,N_551);
nor U1060 (N_1060,N_599,N_666);
xor U1061 (N_1061,N_839,N_833);
and U1062 (N_1062,N_624,N_781);
and U1063 (N_1063,N_712,N_802);
or U1064 (N_1064,N_764,N_931);
and U1065 (N_1065,N_904,N_961);
or U1066 (N_1066,N_695,N_723);
nand U1067 (N_1067,N_967,N_704);
nand U1068 (N_1068,N_728,N_880);
xor U1069 (N_1069,N_610,N_648);
and U1070 (N_1070,N_891,N_646);
and U1071 (N_1071,N_942,N_937);
and U1072 (N_1072,N_658,N_584);
or U1073 (N_1073,N_746,N_808);
and U1074 (N_1074,N_792,N_925);
nand U1075 (N_1075,N_684,N_619);
nand U1076 (N_1076,N_698,N_511);
or U1077 (N_1077,N_903,N_615);
nor U1078 (N_1078,N_886,N_900);
and U1079 (N_1079,N_915,N_748);
nand U1080 (N_1080,N_514,N_919);
nand U1081 (N_1081,N_970,N_796);
and U1082 (N_1082,N_908,N_852);
and U1083 (N_1083,N_593,N_592);
nand U1084 (N_1084,N_795,N_556);
nand U1085 (N_1085,N_703,N_951);
and U1086 (N_1086,N_862,N_756);
nand U1087 (N_1087,N_843,N_999);
or U1088 (N_1088,N_820,N_539);
and U1089 (N_1089,N_733,N_784);
nand U1090 (N_1090,N_949,N_957);
nor U1091 (N_1091,N_754,N_543);
or U1092 (N_1092,N_679,N_620);
nor U1093 (N_1093,N_867,N_954);
nand U1094 (N_1094,N_910,N_699);
nand U1095 (N_1095,N_591,N_557);
xnor U1096 (N_1096,N_562,N_962);
or U1097 (N_1097,N_894,N_707);
and U1098 (N_1098,N_960,N_767);
nand U1099 (N_1099,N_831,N_830);
xnor U1100 (N_1100,N_979,N_560);
and U1101 (N_1101,N_669,N_841);
nand U1102 (N_1102,N_674,N_995);
or U1103 (N_1103,N_508,N_525);
or U1104 (N_1104,N_561,N_503);
nor U1105 (N_1105,N_700,N_687);
and U1106 (N_1106,N_909,N_770);
or U1107 (N_1107,N_807,N_998);
nor U1108 (N_1108,N_813,N_944);
or U1109 (N_1109,N_673,N_667);
nand U1110 (N_1110,N_863,N_729);
nand U1111 (N_1111,N_597,N_758);
or U1112 (N_1112,N_581,N_652);
nor U1113 (N_1113,N_980,N_917);
or U1114 (N_1114,N_941,N_570);
xnor U1115 (N_1115,N_576,N_778);
and U1116 (N_1116,N_547,N_647);
nand U1117 (N_1117,N_822,N_845);
nor U1118 (N_1118,N_826,N_665);
nand U1119 (N_1119,N_834,N_974);
nand U1120 (N_1120,N_512,N_768);
nand U1121 (N_1121,N_549,N_801);
nand U1122 (N_1122,N_545,N_753);
nand U1123 (N_1123,N_788,N_824);
nand U1124 (N_1124,N_955,N_629);
and U1125 (N_1125,N_959,N_924);
or U1126 (N_1126,N_920,N_631);
or U1127 (N_1127,N_987,N_540);
and U1128 (N_1128,N_701,N_765);
nand U1129 (N_1129,N_644,N_725);
nor U1130 (N_1130,N_685,N_580);
and U1131 (N_1131,N_777,N_535);
nand U1132 (N_1132,N_662,N_763);
nor U1133 (N_1133,N_897,N_817);
or U1134 (N_1134,N_507,N_573);
nor U1135 (N_1135,N_553,N_873);
nand U1136 (N_1136,N_655,N_994);
and U1137 (N_1137,N_534,N_815);
nand U1138 (N_1138,N_950,N_632);
nand U1139 (N_1139,N_769,N_572);
nor U1140 (N_1140,N_835,N_877);
nand U1141 (N_1141,N_846,N_975);
nand U1142 (N_1142,N_709,N_513);
and U1143 (N_1143,N_876,N_898);
nor U1144 (N_1144,N_574,N_805);
and U1145 (N_1145,N_548,N_583);
or U1146 (N_1146,N_741,N_642);
or U1147 (N_1147,N_509,N_789);
xor U1148 (N_1148,N_563,N_762);
nor U1149 (N_1149,N_743,N_664);
nor U1150 (N_1150,N_857,N_633);
and U1151 (N_1151,N_866,N_823);
or U1152 (N_1152,N_717,N_895);
and U1153 (N_1153,N_971,N_934);
and U1154 (N_1154,N_538,N_600);
and U1155 (N_1155,N_558,N_623);
and U1156 (N_1156,N_670,N_663);
or U1157 (N_1157,N_671,N_659);
nand U1158 (N_1158,N_505,N_922);
or U1159 (N_1159,N_676,N_579);
nor U1160 (N_1160,N_710,N_520);
and U1161 (N_1161,N_568,N_500);
nand U1162 (N_1162,N_594,N_798);
or U1163 (N_1163,N_927,N_675);
or U1164 (N_1164,N_849,N_978);
nor U1165 (N_1165,N_878,N_800);
and U1166 (N_1166,N_596,N_726);
or U1167 (N_1167,N_618,N_721);
or U1168 (N_1168,N_986,N_533);
or U1169 (N_1169,N_882,N_861);
nand U1170 (N_1170,N_783,N_809);
and U1171 (N_1171,N_711,N_506);
and U1172 (N_1172,N_860,N_577);
nor U1173 (N_1173,N_650,N_649);
and U1174 (N_1174,N_825,N_926);
xnor U1175 (N_1175,N_832,N_794);
and U1176 (N_1176,N_851,N_945);
nor U1177 (N_1177,N_988,N_968);
and U1178 (N_1178,N_761,N_656);
nor U1179 (N_1179,N_879,N_645);
and U1180 (N_1180,N_713,N_604);
or U1181 (N_1181,N_791,N_836);
and U1182 (N_1182,N_612,N_953);
nand U1183 (N_1183,N_848,N_722);
nand U1184 (N_1184,N_643,N_715);
or U1185 (N_1185,N_541,N_559);
and U1186 (N_1186,N_588,N_923);
nor U1187 (N_1187,N_526,N_730);
nand U1188 (N_1188,N_716,N_938);
nor U1189 (N_1189,N_678,N_947);
or U1190 (N_1190,N_985,N_930);
and U1191 (N_1191,N_530,N_621);
or U1192 (N_1192,N_921,N_829);
and U1193 (N_1193,N_518,N_586);
nand U1194 (N_1194,N_812,N_929);
nand U1195 (N_1195,N_689,N_785);
or U1196 (N_1196,N_799,N_911);
nand U1197 (N_1197,N_865,N_842);
or U1198 (N_1198,N_932,N_578);
nand U1199 (N_1199,N_544,N_991);
nor U1200 (N_1200,N_972,N_816);
nand U1201 (N_1201,N_956,N_536);
nor U1202 (N_1202,N_682,N_696);
and U1203 (N_1203,N_690,N_681);
nand U1204 (N_1204,N_912,N_531);
xnor U1205 (N_1205,N_660,N_751);
or U1206 (N_1206,N_693,N_874);
nand U1207 (N_1207,N_771,N_804);
or U1208 (N_1208,N_702,N_964);
or U1209 (N_1209,N_564,N_939);
nand U1210 (N_1210,N_965,N_818);
nor U1211 (N_1211,N_528,N_532);
or U1212 (N_1212,N_521,N_872);
and U1213 (N_1213,N_814,N_727);
and U1214 (N_1214,N_567,N_522);
nand U1215 (N_1215,N_680,N_853);
nand U1216 (N_1216,N_776,N_552);
xnor U1217 (N_1217,N_892,N_582);
or U1218 (N_1218,N_906,N_529);
xnor U1219 (N_1219,N_933,N_731);
nand U1220 (N_1220,N_734,N_918);
or U1221 (N_1221,N_773,N_864);
xor U1222 (N_1222,N_692,N_516);
or U1223 (N_1223,N_668,N_840);
and U1224 (N_1224,N_838,N_683);
or U1225 (N_1225,N_806,N_555);
nand U1226 (N_1226,N_595,N_708);
and U1227 (N_1227,N_963,N_627);
and U1228 (N_1228,N_797,N_847);
nand U1229 (N_1229,N_605,N_973);
nand U1230 (N_1230,N_855,N_630);
nor U1231 (N_1231,N_859,N_837);
or U1232 (N_1232,N_981,N_782);
nand U1233 (N_1233,N_984,N_983);
or U1234 (N_1234,N_718,N_905);
nand U1235 (N_1235,N_871,N_916);
or U1236 (N_1236,N_565,N_501);
nand U1237 (N_1237,N_735,N_706);
nand U1238 (N_1238,N_875,N_969);
nor U1239 (N_1239,N_884,N_819);
or U1240 (N_1240,N_571,N_714);
nand U1241 (N_1241,N_752,N_989);
or U1242 (N_1242,N_883,N_587);
nor U1243 (N_1243,N_810,N_609);
nand U1244 (N_1244,N_990,N_790);
nand U1245 (N_1245,N_774,N_542);
or U1246 (N_1246,N_976,N_793);
and U1247 (N_1247,N_940,N_527);
nand U1248 (N_1248,N_997,N_502);
or U1249 (N_1249,N_821,N_966);
and U1250 (N_1250,N_869,N_996);
and U1251 (N_1251,N_825,N_781);
or U1252 (N_1252,N_541,N_999);
nand U1253 (N_1253,N_653,N_820);
or U1254 (N_1254,N_701,N_913);
or U1255 (N_1255,N_857,N_801);
nand U1256 (N_1256,N_648,N_541);
nor U1257 (N_1257,N_518,N_712);
nand U1258 (N_1258,N_993,N_580);
or U1259 (N_1259,N_650,N_771);
or U1260 (N_1260,N_644,N_712);
nand U1261 (N_1261,N_544,N_879);
nand U1262 (N_1262,N_635,N_734);
nor U1263 (N_1263,N_758,N_737);
nor U1264 (N_1264,N_616,N_952);
nor U1265 (N_1265,N_786,N_592);
nand U1266 (N_1266,N_708,N_589);
nor U1267 (N_1267,N_774,N_877);
nor U1268 (N_1268,N_619,N_527);
nor U1269 (N_1269,N_517,N_866);
and U1270 (N_1270,N_738,N_975);
or U1271 (N_1271,N_996,N_560);
nand U1272 (N_1272,N_737,N_966);
nand U1273 (N_1273,N_848,N_514);
or U1274 (N_1274,N_878,N_983);
nor U1275 (N_1275,N_862,N_705);
xnor U1276 (N_1276,N_667,N_883);
nor U1277 (N_1277,N_953,N_877);
or U1278 (N_1278,N_509,N_817);
nor U1279 (N_1279,N_586,N_855);
or U1280 (N_1280,N_781,N_853);
and U1281 (N_1281,N_622,N_553);
or U1282 (N_1282,N_785,N_709);
and U1283 (N_1283,N_662,N_508);
and U1284 (N_1284,N_714,N_578);
nand U1285 (N_1285,N_889,N_902);
or U1286 (N_1286,N_934,N_561);
or U1287 (N_1287,N_698,N_729);
or U1288 (N_1288,N_786,N_796);
nor U1289 (N_1289,N_746,N_947);
nand U1290 (N_1290,N_608,N_551);
and U1291 (N_1291,N_730,N_959);
or U1292 (N_1292,N_713,N_804);
nand U1293 (N_1293,N_757,N_617);
nand U1294 (N_1294,N_942,N_589);
nor U1295 (N_1295,N_921,N_957);
and U1296 (N_1296,N_564,N_510);
xnor U1297 (N_1297,N_918,N_503);
nor U1298 (N_1298,N_775,N_649);
or U1299 (N_1299,N_652,N_644);
and U1300 (N_1300,N_588,N_632);
nand U1301 (N_1301,N_630,N_862);
and U1302 (N_1302,N_807,N_761);
nand U1303 (N_1303,N_920,N_745);
and U1304 (N_1304,N_859,N_586);
and U1305 (N_1305,N_784,N_746);
nand U1306 (N_1306,N_991,N_865);
and U1307 (N_1307,N_996,N_620);
and U1308 (N_1308,N_883,N_804);
or U1309 (N_1309,N_828,N_898);
nor U1310 (N_1310,N_869,N_969);
nand U1311 (N_1311,N_646,N_581);
nand U1312 (N_1312,N_981,N_887);
nor U1313 (N_1313,N_600,N_850);
and U1314 (N_1314,N_607,N_991);
and U1315 (N_1315,N_975,N_905);
and U1316 (N_1316,N_759,N_920);
and U1317 (N_1317,N_649,N_923);
nand U1318 (N_1318,N_906,N_558);
nor U1319 (N_1319,N_601,N_939);
or U1320 (N_1320,N_630,N_561);
nand U1321 (N_1321,N_622,N_679);
or U1322 (N_1322,N_748,N_643);
nor U1323 (N_1323,N_634,N_791);
and U1324 (N_1324,N_535,N_660);
or U1325 (N_1325,N_627,N_834);
xnor U1326 (N_1326,N_580,N_546);
nand U1327 (N_1327,N_521,N_540);
or U1328 (N_1328,N_644,N_749);
nand U1329 (N_1329,N_836,N_531);
and U1330 (N_1330,N_581,N_708);
and U1331 (N_1331,N_822,N_922);
or U1332 (N_1332,N_881,N_586);
nor U1333 (N_1333,N_686,N_919);
and U1334 (N_1334,N_791,N_627);
nor U1335 (N_1335,N_587,N_801);
or U1336 (N_1336,N_845,N_693);
or U1337 (N_1337,N_619,N_905);
or U1338 (N_1338,N_656,N_777);
nor U1339 (N_1339,N_693,N_866);
or U1340 (N_1340,N_971,N_947);
or U1341 (N_1341,N_660,N_845);
and U1342 (N_1342,N_759,N_823);
and U1343 (N_1343,N_873,N_563);
or U1344 (N_1344,N_887,N_987);
or U1345 (N_1345,N_787,N_806);
and U1346 (N_1346,N_630,N_736);
or U1347 (N_1347,N_892,N_743);
and U1348 (N_1348,N_751,N_783);
nor U1349 (N_1349,N_641,N_954);
nor U1350 (N_1350,N_790,N_666);
or U1351 (N_1351,N_934,N_987);
and U1352 (N_1352,N_835,N_528);
or U1353 (N_1353,N_726,N_602);
and U1354 (N_1354,N_696,N_941);
nand U1355 (N_1355,N_923,N_904);
nor U1356 (N_1356,N_704,N_674);
nand U1357 (N_1357,N_713,N_775);
nand U1358 (N_1358,N_683,N_600);
nand U1359 (N_1359,N_829,N_549);
and U1360 (N_1360,N_935,N_627);
or U1361 (N_1361,N_974,N_792);
and U1362 (N_1362,N_953,N_723);
or U1363 (N_1363,N_848,N_564);
and U1364 (N_1364,N_634,N_560);
or U1365 (N_1365,N_842,N_525);
xnor U1366 (N_1366,N_853,N_524);
nand U1367 (N_1367,N_536,N_903);
or U1368 (N_1368,N_601,N_524);
or U1369 (N_1369,N_639,N_803);
nand U1370 (N_1370,N_619,N_867);
or U1371 (N_1371,N_760,N_905);
and U1372 (N_1372,N_948,N_709);
and U1373 (N_1373,N_684,N_696);
and U1374 (N_1374,N_908,N_923);
nor U1375 (N_1375,N_875,N_949);
nand U1376 (N_1376,N_606,N_961);
nand U1377 (N_1377,N_745,N_578);
nor U1378 (N_1378,N_577,N_715);
nor U1379 (N_1379,N_754,N_969);
nand U1380 (N_1380,N_948,N_611);
xnor U1381 (N_1381,N_559,N_663);
or U1382 (N_1382,N_546,N_767);
or U1383 (N_1383,N_517,N_921);
and U1384 (N_1384,N_769,N_555);
or U1385 (N_1385,N_778,N_613);
nor U1386 (N_1386,N_795,N_987);
xnor U1387 (N_1387,N_550,N_817);
nand U1388 (N_1388,N_563,N_619);
and U1389 (N_1389,N_570,N_992);
and U1390 (N_1390,N_807,N_819);
nor U1391 (N_1391,N_797,N_845);
nand U1392 (N_1392,N_752,N_901);
nand U1393 (N_1393,N_785,N_975);
nand U1394 (N_1394,N_876,N_669);
or U1395 (N_1395,N_544,N_870);
xor U1396 (N_1396,N_993,N_506);
xor U1397 (N_1397,N_915,N_946);
nor U1398 (N_1398,N_756,N_743);
and U1399 (N_1399,N_906,N_626);
nand U1400 (N_1400,N_941,N_971);
nor U1401 (N_1401,N_633,N_813);
or U1402 (N_1402,N_825,N_729);
nor U1403 (N_1403,N_518,N_550);
nand U1404 (N_1404,N_895,N_536);
or U1405 (N_1405,N_632,N_909);
nor U1406 (N_1406,N_961,N_622);
nor U1407 (N_1407,N_681,N_710);
nor U1408 (N_1408,N_690,N_827);
and U1409 (N_1409,N_517,N_770);
or U1410 (N_1410,N_712,N_759);
or U1411 (N_1411,N_694,N_725);
nand U1412 (N_1412,N_685,N_824);
nand U1413 (N_1413,N_960,N_576);
nand U1414 (N_1414,N_844,N_898);
or U1415 (N_1415,N_605,N_869);
and U1416 (N_1416,N_615,N_576);
nand U1417 (N_1417,N_770,N_563);
nand U1418 (N_1418,N_794,N_528);
or U1419 (N_1419,N_655,N_592);
nor U1420 (N_1420,N_764,N_614);
and U1421 (N_1421,N_678,N_696);
nor U1422 (N_1422,N_539,N_669);
nor U1423 (N_1423,N_984,N_866);
nor U1424 (N_1424,N_936,N_749);
nor U1425 (N_1425,N_733,N_855);
nor U1426 (N_1426,N_610,N_966);
nand U1427 (N_1427,N_589,N_508);
nand U1428 (N_1428,N_650,N_580);
and U1429 (N_1429,N_571,N_635);
or U1430 (N_1430,N_822,N_912);
and U1431 (N_1431,N_949,N_888);
nor U1432 (N_1432,N_775,N_949);
nor U1433 (N_1433,N_883,N_931);
and U1434 (N_1434,N_572,N_901);
and U1435 (N_1435,N_758,N_700);
nor U1436 (N_1436,N_780,N_639);
nand U1437 (N_1437,N_656,N_693);
nor U1438 (N_1438,N_504,N_533);
nor U1439 (N_1439,N_879,N_563);
or U1440 (N_1440,N_917,N_631);
and U1441 (N_1441,N_918,N_707);
nand U1442 (N_1442,N_718,N_541);
or U1443 (N_1443,N_989,N_873);
or U1444 (N_1444,N_737,N_704);
nor U1445 (N_1445,N_824,N_543);
nor U1446 (N_1446,N_969,N_586);
or U1447 (N_1447,N_777,N_905);
nand U1448 (N_1448,N_733,N_826);
and U1449 (N_1449,N_512,N_647);
nor U1450 (N_1450,N_689,N_912);
nor U1451 (N_1451,N_659,N_579);
nor U1452 (N_1452,N_760,N_894);
or U1453 (N_1453,N_977,N_917);
and U1454 (N_1454,N_858,N_737);
nand U1455 (N_1455,N_989,N_696);
nand U1456 (N_1456,N_870,N_743);
and U1457 (N_1457,N_502,N_521);
xnor U1458 (N_1458,N_631,N_720);
nor U1459 (N_1459,N_897,N_762);
nor U1460 (N_1460,N_630,N_771);
nor U1461 (N_1461,N_676,N_872);
or U1462 (N_1462,N_915,N_849);
nor U1463 (N_1463,N_946,N_512);
nor U1464 (N_1464,N_797,N_624);
and U1465 (N_1465,N_545,N_841);
nor U1466 (N_1466,N_582,N_904);
nand U1467 (N_1467,N_688,N_979);
and U1468 (N_1468,N_985,N_724);
nand U1469 (N_1469,N_655,N_656);
and U1470 (N_1470,N_987,N_960);
and U1471 (N_1471,N_648,N_582);
nor U1472 (N_1472,N_657,N_975);
and U1473 (N_1473,N_746,N_526);
nand U1474 (N_1474,N_633,N_852);
or U1475 (N_1475,N_736,N_716);
nand U1476 (N_1476,N_544,N_817);
or U1477 (N_1477,N_700,N_668);
or U1478 (N_1478,N_717,N_666);
or U1479 (N_1479,N_956,N_621);
and U1480 (N_1480,N_908,N_513);
or U1481 (N_1481,N_692,N_731);
xor U1482 (N_1482,N_526,N_680);
nand U1483 (N_1483,N_987,N_900);
or U1484 (N_1484,N_504,N_729);
or U1485 (N_1485,N_622,N_687);
and U1486 (N_1486,N_609,N_597);
nand U1487 (N_1487,N_548,N_785);
xor U1488 (N_1488,N_737,N_689);
or U1489 (N_1489,N_590,N_858);
and U1490 (N_1490,N_994,N_701);
nor U1491 (N_1491,N_978,N_880);
and U1492 (N_1492,N_946,N_959);
or U1493 (N_1493,N_823,N_640);
and U1494 (N_1494,N_577,N_619);
and U1495 (N_1495,N_999,N_638);
and U1496 (N_1496,N_860,N_825);
nand U1497 (N_1497,N_930,N_544);
nand U1498 (N_1498,N_924,N_911);
nand U1499 (N_1499,N_724,N_988);
and U1500 (N_1500,N_1150,N_1308);
xor U1501 (N_1501,N_1028,N_1186);
nand U1502 (N_1502,N_1174,N_1219);
nor U1503 (N_1503,N_1426,N_1417);
and U1504 (N_1504,N_1194,N_1310);
nand U1505 (N_1505,N_1156,N_1299);
or U1506 (N_1506,N_1175,N_1303);
and U1507 (N_1507,N_1343,N_1055);
nand U1508 (N_1508,N_1189,N_1233);
and U1509 (N_1509,N_1119,N_1063);
and U1510 (N_1510,N_1406,N_1444);
or U1511 (N_1511,N_1439,N_1448);
nor U1512 (N_1512,N_1145,N_1167);
and U1513 (N_1513,N_1155,N_1226);
and U1514 (N_1514,N_1181,N_1024);
or U1515 (N_1515,N_1239,N_1487);
nand U1516 (N_1516,N_1093,N_1405);
nand U1517 (N_1517,N_1411,N_1441);
or U1518 (N_1518,N_1260,N_1038);
and U1519 (N_1519,N_1330,N_1252);
nand U1520 (N_1520,N_1435,N_1270);
and U1521 (N_1521,N_1068,N_1296);
nor U1522 (N_1522,N_1169,N_1446);
nand U1523 (N_1523,N_1277,N_1424);
and U1524 (N_1524,N_1412,N_1257);
nand U1525 (N_1525,N_1345,N_1229);
or U1526 (N_1526,N_1264,N_1042);
or U1527 (N_1527,N_1211,N_1004);
nand U1528 (N_1528,N_1022,N_1153);
nor U1529 (N_1529,N_1466,N_1123);
and U1530 (N_1530,N_1176,N_1165);
or U1531 (N_1531,N_1253,N_1146);
nand U1532 (N_1532,N_1114,N_1320);
or U1533 (N_1533,N_1416,N_1212);
nand U1534 (N_1534,N_1242,N_1287);
or U1535 (N_1535,N_1368,N_1421);
or U1536 (N_1536,N_1402,N_1099);
nand U1537 (N_1537,N_1104,N_1065);
or U1538 (N_1538,N_1061,N_1127);
nor U1539 (N_1539,N_1386,N_1143);
xnor U1540 (N_1540,N_1428,N_1216);
and U1541 (N_1541,N_1003,N_1274);
or U1542 (N_1542,N_1295,N_1147);
or U1543 (N_1543,N_1465,N_1327);
nand U1544 (N_1544,N_1305,N_1263);
nor U1545 (N_1545,N_1018,N_1034);
or U1546 (N_1546,N_1497,N_1125);
nand U1547 (N_1547,N_1318,N_1098);
nor U1548 (N_1548,N_1076,N_1188);
nor U1549 (N_1549,N_1362,N_1047);
nand U1550 (N_1550,N_1383,N_1302);
nand U1551 (N_1551,N_1333,N_1053);
or U1552 (N_1552,N_1050,N_1381);
and U1553 (N_1553,N_1095,N_1471);
nor U1554 (N_1554,N_1431,N_1283);
and U1555 (N_1555,N_1344,N_1020);
nor U1556 (N_1556,N_1185,N_1377);
or U1557 (N_1557,N_1373,N_1397);
or U1558 (N_1558,N_1342,N_1290);
and U1559 (N_1559,N_1225,N_1467);
nor U1560 (N_1560,N_1419,N_1403);
and U1561 (N_1561,N_1463,N_1245);
nand U1562 (N_1562,N_1473,N_1140);
or U1563 (N_1563,N_1315,N_1170);
or U1564 (N_1564,N_1039,N_1035);
and U1565 (N_1565,N_1021,N_1031);
and U1566 (N_1566,N_1009,N_1255);
and U1567 (N_1567,N_1361,N_1187);
and U1568 (N_1568,N_1273,N_1027);
nor U1569 (N_1569,N_1112,N_1321);
nand U1570 (N_1570,N_1470,N_1158);
nor U1571 (N_1571,N_1414,N_1026);
or U1572 (N_1572,N_1477,N_1399);
nor U1573 (N_1573,N_1340,N_1266);
nor U1574 (N_1574,N_1429,N_1457);
nand U1575 (N_1575,N_1173,N_1032);
or U1576 (N_1576,N_1415,N_1083);
nor U1577 (N_1577,N_1152,N_1409);
and U1578 (N_1578,N_1102,N_1052);
and U1579 (N_1579,N_1336,N_1496);
nor U1580 (N_1580,N_1218,N_1197);
or U1581 (N_1581,N_1058,N_1071);
or U1582 (N_1582,N_1331,N_1030);
nor U1583 (N_1583,N_1060,N_1408);
and U1584 (N_1584,N_1351,N_1199);
nand U1585 (N_1585,N_1434,N_1319);
and U1586 (N_1586,N_1012,N_1278);
and U1587 (N_1587,N_1388,N_1232);
or U1588 (N_1588,N_1371,N_1097);
nand U1589 (N_1589,N_1171,N_1349);
or U1590 (N_1590,N_1258,N_1442);
and U1591 (N_1591,N_1350,N_1096);
and U1592 (N_1592,N_1235,N_1285);
and U1593 (N_1593,N_1248,N_1089);
and U1594 (N_1594,N_1142,N_1490);
nand U1595 (N_1595,N_1224,N_1328);
or U1596 (N_1596,N_1043,N_1198);
and U1597 (N_1597,N_1276,N_1046);
and U1598 (N_1598,N_1067,N_1495);
nor U1599 (N_1599,N_1370,N_1352);
or U1600 (N_1600,N_1369,N_1192);
or U1601 (N_1601,N_1432,N_1313);
nor U1602 (N_1602,N_1385,N_1182);
and U1603 (N_1603,N_1390,N_1491);
nor U1604 (N_1604,N_1124,N_1401);
nor U1605 (N_1605,N_1019,N_1375);
nor U1606 (N_1606,N_1374,N_1324);
and U1607 (N_1607,N_1100,N_1433);
nand U1608 (N_1608,N_1016,N_1472);
nor U1609 (N_1609,N_1163,N_1438);
and U1610 (N_1610,N_1382,N_1037);
nor U1611 (N_1611,N_1480,N_1279);
nand U1612 (N_1612,N_1304,N_1400);
and U1613 (N_1613,N_1291,N_1025);
and U1614 (N_1614,N_1110,N_1256);
or U1615 (N_1615,N_1307,N_1081);
and U1616 (N_1616,N_1230,N_1062);
xnor U1617 (N_1617,N_1306,N_1418);
or U1618 (N_1618,N_1059,N_1006);
nor U1619 (N_1619,N_1001,N_1474);
nor U1620 (N_1620,N_1014,N_1184);
nand U1621 (N_1621,N_1479,N_1178);
and U1622 (N_1622,N_1348,N_1384);
nand U1623 (N_1623,N_1222,N_1109);
nand U1624 (N_1624,N_1316,N_1422);
or U1625 (N_1625,N_1073,N_1389);
nor U1626 (N_1626,N_1183,N_1223);
and U1627 (N_1627,N_1492,N_1300);
nor U1628 (N_1628,N_1293,N_1393);
nand U1629 (N_1629,N_1332,N_1440);
nand U1630 (N_1630,N_1215,N_1107);
and U1631 (N_1631,N_1135,N_1423);
or U1632 (N_1632,N_1129,N_1164);
or U1633 (N_1633,N_1051,N_1262);
and U1634 (N_1634,N_1378,N_1002);
or U1635 (N_1635,N_1337,N_1115);
nand U1636 (N_1636,N_1220,N_1354);
and U1637 (N_1637,N_1066,N_1040);
nor U1638 (N_1638,N_1103,N_1111);
nand U1639 (N_1639,N_1407,N_1070);
or U1640 (N_1640,N_1149,N_1338);
nand U1641 (N_1641,N_1138,N_1203);
nor U1642 (N_1642,N_1394,N_1092);
nor U1643 (N_1643,N_1484,N_1395);
nand U1644 (N_1644,N_1254,N_1353);
and U1645 (N_1645,N_1054,N_1010);
and U1646 (N_1646,N_1478,N_1207);
or U1647 (N_1647,N_1271,N_1284);
or U1648 (N_1648,N_1269,N_1227);
xnor U1649 (N_1649,N_1005,N_1447);
nor U1650 (N_1650,N_1317,N_1468);
and U1651 (N_1651,N_1455,N_1168);
xnor U1652 (N_1652,N_1234,N_1380);
or U1653 (N_1653,N_1159,N_1392);
and U1654 (N_1654,N_1202,N_1161);
nand U1655 (N_1655,N_1275,N_1136);
nand U1656 (N_1656,N_1160,N_1072);
and U1657 (N_1657,N_1281,N_1356);
or U1658 (N_1658,N_1221,N_1476);
nand U1659 (N_1659,N_1339,N_1325);
nand U1660 (N_1660,N_1048,N_1108);
or U1661 (N_1661,N_1311,N_1133);
nor U1662 (N_1662,N_1355,N_1341);
and U1663 (N_1663,N_1314,N_1210);
nor U1664 (N_1664,N_1461,N_1036);
nor U1665 (N_1665,N_1334,N_1425);
or U1666 (N_1666,N_1074,N_1292);
or U1667 (N_1667,N_1286,N_1236);
nand U1668 (N_1668,N_1458,N_1017);
nand U1669 (N_1669,N_1195,N_1204);
nor U1670 (N_1670,N_1301,N_1106);
nor U1671 (N_1671,N_1118,N_1084);
nor U1672 (N_1672,N_1462,N_1090);
nand U1673 (N_1673,N_1113,N_1193);
nor U1674 (N_1674,N_1452,N_1259);
or U1675 (N_1675,N_1445,N_1086);
or U1676 (N_1676,N_1120,N_1213);
nor U1677 (N_1677,N_1075,N_1488);
and U1678 (N_1678,N_1045,N_1064);
nor U1679 (N_1679,N_1029,N_1240);
nand U1680 (N_1680,N_1359,N_1312);
or U1681 (N_1681,N_1126,N_1196);
nand U1682 (N_1682,N_1117,N_1346);
and U1683 (N_1683,N_1366,N_1007);
nor U1684 (N_1684,N_1464,N_1105);
and U1685 (N_1685,N_1116,N_1033);
nand U1686 (N_1686,N_1011,N_1294);
nor U1687 (N_1687,N_1357,N_1451);
nor U1688 (N_1688,N_1238,N_1217);
nor U1689 (N_1689,N_1231,N_1122);
and U1690 (N_1690,N_1326,N_1200);
and U1691 (N_1691,N_1398,N_1130);
nor U1692 (N_1692,N_1134,N_1413);
or U1693 (N_1693,N_1453,N_1372);
nor U1694 (N_1694,N_1044,N_1209);
nand U1695 (N_1695,N_1013,N_1282);
nand U1696 (N_1696,N_1128,N_1085);
nor U1697 (N_1697,N_1154,N_1148);
nor U1698 (N_1698,N_1469,N_1094);
or U1699 (N_1699,N_1190,N_1481);
and U1700 (N_1700,N_1244,N_1243);
or U1701 (N_1701,N_1079,N_1191);
nor U1702 (N_1702,N_1347,N_1077);
or U1703 (N_1703,N_1486,N_1499);
and U1704 (N_1704,N_1268,N_1437);
xor U1705 (N_1705,N_1162,N_1443);
and U1706 (N_1706,N_1379,N_1267);
or U1707 (N_1707,N_1228,N_1214);
nor U1708 (N_1708,N_1206,N_1475);
nand U1709 (N_1709,N_1420,N_1121);
nand U1710 (N_1710,N_1289,N_1251);
nor U1711 (N_1711,N_1323,N_1141);
or U1712 (N_1712,N_1404,N_1363);
nand U1713 (N_1713,N_1456,N_1131);
and U1714 (N_1714,N_1396,N_1460);
nor U1715 (N_1715,N_1023,N_1201);
and U1716 (N_1716,N_1087,N_1246);
and U1717 (N_1717,N_1483,N_1205);
or U1718 (N_1718,N_1008,N_1049);
and U1719 (N_1719,N_1391,N_1247);
nand U1720 (N_1720,N_1335,N_1288);
nand U1721 (N_1721,N_1265,N_1069);
and U1722 (N_1722,N_1137,N_1241);
and U1723 (N_1723,N_1272,N_1322);
and U1724 (N_1724,N_1482,N_1151);
or U1725 (N_1725,N_1298,N_1056);
nor U1726 (N_1726,N_1365,N_1015);
and U1727 (N_1727,N_1427,N_1489);
or U1728 (N_1728,N_1367,N_1080);
xnor U1729 (N_1729,N_1494,N_1376);
or U1730 (N_1730,N_1430,N_1387);
nand U1731 (N_1731,N_1208,N_1261);
nand U1732 (N_1732,N_1180,N_1091);
nor U1733 (N_1733,N_1249,N_1329);
nand U1734 (N_1734,N_1360,N_1493);
nand U1735 (N_1735,N_1041,N_1078);
nor U1736 (N_1736,N_1177,N_1450);
nand U1737 (N_1737,N_1157,N_1358);
nand U1738 (N_1738,N_1139,N_1449);
and U1739 (N_1739,N_1309,N_1082);
and U1740 (N_1740,N_1459,N_1237);
and U1741 (N_1741,N_1088,N_1297);
and U1742 (N_1742,N_1364,N_1498);
and U1743 (N_1743,N_1144,N_1280);
xor U1744 (N_1744,N_1179,N_1057);
nand U1745 (N_1745,N_1101,N_1132);
nand U1746 (N_1746,N_1436,N_1454);
or U1747 (N_1747,N_1410,N_1000);
nor U1748 (N_1748,N_1250,N_1172);
and U1749 (N_1749,N_1485,N_1166);
nand U1750 (N_1750,N_1384,N_1060);
or U1751 (N_1751,N_1397,N_1151);
or U1752 (N_1752,N_1422,N_1040);
nor U1753 (N_1753,N_1184,N_1331);
nor U1754 (N_1754,N_1185,N_1109);
or U1755 (N_1755,N_1494,N_1030);
nand U1756 (N_1756,N_1406,N_1123);
nand U1757 (N_1757,N_1250,N_1010);
nand U1758 (N_1758,N_1468,N_1390);
nand U1759 (N_1759,N_1204,N_1093);
and U1760 (N_1760,N_1055,N_1382);
nand U1761 (N_1761,N_1108,N_1295);
nor U1762 (N_1762,N_1069,N_1206);
xor U1763 (N_1763,N_1053,N_1171);
and U1764 (N_1764,N_1335,N_1092);
or U1765 (N_1765,N_1182,N_1264);
nor U1766 (N_1766,N_1488,N_1479);
and U1767 (N_1767,N_1260,N_1051);
nand U1768 (N_1768,N_1148,N_1303);
nor U1769 (N_1769,N_1324,N_1499);
nand U1770 (N_1770,N_1030,N_1001);
or U1771 (N_1771,N_1082,N_1182);
nor U1772 (N_1772,N_1222,N_1326);
and U1773 (N_1773,N_1288,N_1458);
nor U1774 (N_1774,N_1115,N_1093);
nor U1775 (N_1775,N_1230,N_1135);
and U1776 (N_1776,N_1400,N_1461);
nor U1777 (N_1777,N_1378,N_1474);
nor U1778 (N_1778,N_1368,N_1073);
nand U1779 (N_1779,N_1294,N_1049);
or U1780 (N_1780,N_1108,N_1063);
and U1781 (N_1781,N_1129,N_1093);
nor U1782 (N_1782,N_1158,N_1446);
nand U1783 (N_1783,N_1117,N_1227);
or U1784 (N_1784,N_1136,N_1072);
xor U1785 (N_1785,N_1323,N_1271);
and U1786 (N_1786,N_1217,N_1288);
and U1787 (N_1787,N_1408,N_1440);
or U1788 (N_1788,N_1234,N_1019);
and U1789 (N_1789,N_1481,N_1110);
nor U1790 (N_1790,N_1438,N_1420);
xnor U1791 (N_1791,N_1424,N_1042);
and U1792 (N_1792,N_1221,N_1375);
or U1793 (N_1793,N_1087,N_1138);
nand U1794 (N_1794,N_1480,N_1036);
nor U1795 (N_1795,N_1294,N_1042);
nand U1796 (N_1796,N_1477,N_1320);
and U1797 (N_1797,N_1064,N_1370);
or U1798 (N_1798,N_1407,N_1152);
and U1799 (N_1799,N_1378,N_1365);
nand U1800 (N_1800,N_1409,N_1053);
nand U1801 (N_1801,N_1124,N_1254);
nor U1802 (N_1802,N_1474,N_1471);
or U1803 (N_1803,N_1205,N_1123);
nor U1804 (N_1804,N_1294,N_1210);
or U1805 (N_1805,N_1473,N_1498);
and U1806 (N_1806,N_1467,N_1173);
nor U1807 (N_1807,N_1275,N_1185);
nor U1808 (N_1808,N_1164,N_1390);
and U1809 (N_1809,N_1070,N_1041);
xor U1810 (N_1810,N_1038,N_1171);
and U1811 (N_1811,N_1377,N_1166);
or U1812 (N_1812,N_1272,N_1253);
nor U1813 (N_1813,N_1289,N_1472);
nand U1814 (N_1814,N_1021,N_1076);
and U1815 (N_1815,N_1476,N_1088);
nand U1816 (N_1816,N_1224,N_1473);
nand U1817 (N_1817,N_1296,N_1036);
nand U1818 (N_1818,N_1419,N_1395);
nor U1819 (N_1819,N_1467,N_1187);
or U1820 (N_1820,N_1096,N_1316);
nand U1821 (N_1821,N_1465,N_1467);
nand U1822 (N_1822,N_1396,N_1044);
or U1823 (N_1823,N_1258,N_1111);
nand U1824 (N_1824,N_1141,N_1153);
and U1825 (N_1825,N_1486,N_1497);
nor U1826 (N_1826,N_1049,N_1396);
nor U1827 (N_1827,N_1017,N_1181);
nand U1828 (N_1828,N_1040,N_1419);
or U1829 (N_1829,N_1159,N_1190);
or U1830 (N_1830,N_1361,N_1329);
or U1831 (N_1831,N_1210,N_1143);
or U1832 (N_1832,N_1284,N_1010);
and U1833 (N_1833,N_1294,N_1262);
and U1834 (N_1834,N_1324,N_1104);
or U1835 (N_1835,N_1229,N_1254);
and U1836 (N_1836,N_1247,N_1356);
and U1837 (N_1837,N_1109,N_1333);
or U1838 (N_1838,N_1126,N_1163);
nand U1839 (N_1839,N_1158,N_1285);
or U1840 (N_1840,N_1237,N_1204);
and U1841 (N_1841,N_1316,N_1054);
xnor U1842 (N_1842,N_1242,N_1113);
nand U1843 (N_1843,N_1475,N_1461);
nand U1844 (N_1844,N_1059,N_1003);
or U1845 (N_1845,N_1494,N_1331);
nand U1846 (N_1846,N_1392,N_1200);
nor U1847 (N_1847,N_1160,N_1046);
nand U1848 (N_1848,N_1490,N_1394);
nand U1849 (N_1849,N_1080,N_1002);
or U1850 (N_1850,N_1429,N_1080);
or U1851 (N_1851,N_1425,N_1459);
xnor U1852 (N_1852,N_1320,N_1333);
and U1853 (N_1853,N_1425,N_1055);
or U1854 (N_1854,N_1265,N_1381);
or U1855 (N_1855,N_1016,N_1020);
or U1856 (N_1856,N_1325,N_1170);
and U1857 (N_1857,N_1046,N_1303);
or U1858 (N_1858,N_1291,N_1311);
and U1859 (N_1859,N_1415,N_1443);
nand U1860 (N_1860,N_1278,N_1180);
xnor U1861 (N_1861,N_1496,N_1081);
and U1862 (N_1862,N_1395,N_1150);
nor U1863 (N_1863,N_1157,N_1214);
and U1864 (N_1864,N_1188,N_1176);
nor U1865 (N_1865,N_1447,N_1253);
nor U1866 (N_1866,N_1470,N_1336);
or U1867 (N_1867,N_1242,N_1411);
nand U1868 (N_1868,N_1312,N_1097);
or U1869 (N_1869,N_1104,N_1066);
nor U1870 (N_1870,N_1125,N_1495);
nor U1871 (N_1871,N_1454,N_1439);
xor U1872 (N_1872,N_1443,N_1463);
nor U1873 (N_1873,N_1484,N_1384);
or U1874 (N_1874,N_1035,N_1163);
and U1875 (N_1875,N_1471,N_1345);
or U1876 (N_1876,N_1148,N_1027);
nor U1877 (N_1877,N_1245,N_1103);
and U1878 (N_1878,N_1029,N_1050);
nor U1879 (N_1879,N_1468,N_1320);
or U1880 (N_1880,N_1208,N_1136);
and U1881 (N_1881,N_1173,N_1351);
and U1882 (N_1882,N_1412,N_1304);
xor U1883 (N_1883,N_1398,N_1353);
or U1884 (N_1884,N_1270,N_1399);
xor U1885 (N_1885,N_1425,N_1085);
nor U1886 (N_1886,N_1467,N_1228);
and U1887 (N_1887,N_1066,N_1402);
nor U1888 (N_1888,N_1056,N_1121);
or U1889 (N_1889,N_1057,N_1008);
and U1890 (N_1890,N_1428,N_1143);
nand U1891 (N_1891,N_1283,N_1007);
nand U1892 (N_1892,N_1277,N_1156);
or U1893 (N_1893,N_1137,N_1022);
nand U1894 (N_1894,N_1230,N_1148);
nor U1895 (N_1895,N_1051,N_1386);
or U1896 (N_1896,N_1307,N_1213);
or U1897 (N_1897,N_1062,N_1322);
or U1898 (N_1898,N_1048,N_1055);
or U1899 (N_1899,N_1054,N_1423);
or U1900 (N_1900,N_1447,N_1055);
nor U1901 (N_1901,N_1009,N_1010);
nand U1902 (N_1902,N_1010,N_1296);
and U1903 (N_1903,N_1462,N_1042);
nor U1904 (N_1904,N_1165,N_1412);
and U1905 (N_1905,N_1299,N_1066);
or U1906 (N_1906,N_1282,N_1425);
and U1907 (N_1907,N_1164,N_1297);
nor U1908 (N_1908,N_1087,N_1079);
and U1909 (N_1909,N_1283,N_1337);
nand U1910 (N_1910,N_1223,N_1149);
xor U1911 (N_1911,N_1073,N_1429);
or U1912 (N_1912,N_1402,N_1465);
and U1913 (N_1913,N_1065,N_1187);
nor U1914 (N_1914,N_1074,N_1460);
xnor U1915 (N_1915,N_1130,N_1127);
or U1916 (N_1916,N_1125,N_1295);
nand U1917 (N_1917,N_1221,N_1004);
and U1918 (N_1918,N_1354,N_1219);
or U1919 (N_1919,N_1278,N_1283);
nor U1920 (N_1920,N_1156,N_1313);
or U1921 (N_1921,N_1375,N_1435);
nand U1922 (N_1922,N_1018,N_1250);
nand U1923 (N_1923,N_1386,N_1351);
or U1924 (N_1924,N_1171,N_1088);
nor U1925 (N_1925,N_1362,N_1116);
nor U1926 (N_1926,N_1471,N_1234);
or U1927 (N_1927,N_1190,N_1253);
or U1928 (N_1928,N_1040,N_1090);
or U1929 (N_1929,N_1088,N_1129);
and U1930 (N_1930,N_1456,N_1476);
or U1931 (N_1931,N_1330,N_1496);
xor U1932 (N_1932,N_1218,N_1384);
nor U1933 (N_1933,N_1122,N_1352);
nor U1934 (N_1934,N_1043,N_1112);
nor U1935 (N_1935,N_1059,N_1104);
or U1936 (N_1936,N_1002,N_1205);
nor U1937 (N_1937,N_1361,N_1432);
nand U1938 (N_1938,N_1200,N_1017);
nor U1939 (N_1939,N_1158,N_1387);
and U1940 (N_1940,N_1062,N_1201);
xnor U1941 (N_1941,N_1120,N_1188);
nand U1942 (N_1942,N_1279,N_1495);
xnor U1943 (N_1943,N_1236,N_1467);
nand U1944 (N_1944,N_1424,N_1097);
and U1945 (N_1945,N_1045,N_1385);
and U1946 (N_1946,N_1270,N_1442);
nand U1947 (N_1947,N_1196,N_1084);
and U1948 (N_1948,N_1006,N_1009);
and U1949 (N_1949,N_1437,N_1160);
and U1950 (N_1950,N_1255,N_1141);
nor U1951 (N_1951,N_1022,N_1207);
and U1952 (N_1952,N_1348,N_1401);
nor U1953 (N_1953,N_1402,N_1248);
xor U1954 (N_1954,N_1124,N_1025);
nor U1955 (N_1955,N_1044,N_1114);
and U1956 (N_1956,N_1269,N_1137);
or U1957 (N_1957,N_1049,N_1302);
or U1958 (N_1958,N_1443,N_1366);
nor U1959 (N_1959,N_1324,N_1313);
and U1960 (N_1960,N_1073,N_1021);
nor U1961 (N_1961,N_1471,N_1179);
or U1962 (N_1962,N_1489,N_1385);
and U1963 (N_1963,N_1046,N_1104);
or U1964 (N_1964,N_1324,N_1441);
or U1965 (N_1965,N_1364,N_1086);
or U1966 (N_1966,N_1251,N_1163);
or U1967 (N_1967,N_1047,N_1048);
or U1968 (N_1968,N_1013,N_1388);
or U1969 (N_1969,N_1415,N_1356);
or U1970 (N_1970,N_1043,N_1268);
and U1971 (N_1971,N_1324,N_1248);
nand U1972 (N_1972,N_1447,N_1024);
or U1973 (N_1973,N_1434,N_1404);
nand U1974 (N_1974,N_1291,N_1163);
nand U1975 (N_1975,N_1142,N_1198);
nand U1976 (N_1976,N_1146,N_1429);
nor U1977 (N_1977,N_1082,N_1221);
nor U1978 (N_1978,N_1415,N_1243);
nor U1979 (N_1979,N_1333,N_1281);
or U1980 (N_1980,N_1113,N_1233);
or U1981 (N_1981,N_1095,N_1042);
and U1982 (N_1982,N_1033,N_1417);
or U1983 (N_1983,N_1226,N_1305);
nand U1984 (N_1984,N_1196,N_1261);
nor U1985 (N_1985,N_1469,N_1352);
and U1986 (N_1986,N_1090,N_1049);
or U1987 (N_1987,N_1451,N_1057);
nand U1988 (N_1988,N_1308,N_1432);
nor U1989 (N_1989,N_1466,N_1394);
or U1990 (N_1990,N_1312,N_1059);
nand U1991 (N_1991,N_1113,N_1403);
and U1992 (N_1992,N_1093,N_1239);
nand U1993 (N_1993,N_1360,N_1125);
nor U1994 (N_1994,N_1058,N_1285);
or U1995 (N_1995,N_1112,N_1144);
nand U1996 (N_1996,N_1131,N_1110);
nand U1997 (N_1997,N_1177,N_1127);
nor U1998 (N_1998,N_1439,N_1007);
or U1999 (N_1999,N_1317,N_1268);
nor U2000 (N_2000,N_1847,N_1723);
or U2001 (N_2001,N_1815,N_1729);
or U2002 (N_2002,N_1687,N_1613);
nand U2003 (N_2003,N_1580,N_1572);
or U2004 (N_2004,N_1955,N_1849);
nor U2005 (N_2005,N_1953,N_1792);
nand U2006 (N_2006,N_1652,N_1625);
or U2007 (N_2007,N_1900,N_1670);
nand U2008 (N_2008,N_1904,N_1990);
and U2009 (N_2009,N_1969,N_1543);
or U2010 (N_2010,N_1784,N_1974);
or U2011 (N_2011,N_1957,N_1938);
nor U2012 (N_2012,N_1759,N_1602);
or U2013 (N_2013,N_1802,N_1735);
nor U2014 (N_2014,N_1901,N_1721);
and U2015 (N_2015,N_1516,N_1888);
nor U2016 (N_2016,N_1728,N_1762);
and U2017 (N_2017,N_1632,N_1547);
nand U2018 (N_2018,N_1563,N_1982);
and U2019 (N_2019,N_1908,N_1927);
or U2020 (N_2020,N_1737,N_1750);
and U2021 (N_2021,N_1756,N_1923);
nand U2022 (N_2022,N_1656,N_1817);
nor U2023 (N_2023,N_1752,N_1520);
or U2024 (N_2024,N_1624,N_1658);
nor U2025 (N_2025,N_1761,N_1626);
or U2026 (N_2026,N_1716,N_1555);
nand U2027 (N_2027,N_1584,N_1781);
or U2028 (N_2028,N_1882,N_1896);
nor U2029 (N_2029,N_1623,N_1913);
or U2030 (N_2030,N_1910,N_1780);
and U2031 (N_2031,N_1607,N_1892);
or U2032 (N_2032,N_1612,N_1726);
nand U2033 (N_2033,N_1573,N_1834);
nand U2034 (N_2034,N_1525,N_1961);
and U2035 (N_2035,N_1918,N_1783);
nor U2036 (N_2036,N_1664,N_1706);
xnor U2037 (N_2037,N_1978,N_1599);
nor U2038 (N_2038,N_1770,N_1765);
and U2039 (N_2039,N_1799,N_1659);
nor U2040 (N_2040,N_1522,N_1775);
or U2041 (N_2041,N_1585,N_1715);
nor U2042 (N_2042,N_1876,N_1504);
nand U2043 (N_2043,N_1546,N_1711);
nor U2044 (N_2044,N_1618,N_1707);
nand U2045 (N_2045,N_1686,N_1965);
xor U2046 (N_2046,N_1785,N_1942);
nor U2047 (N_2047,N_1844,N_1870);
xor U2048 (N_2048,N_1746,N_1542);
nor U2049 (N_2049,N_1669,N_1840);
or U2050 (N_2050,N_1578,N_1651);
nor U2051 (N_2051,N_1524,N_1851);
nand U2052 (N_2052,N_1672,N_1883);
or U2053 (N_2053,N_1601,N_1742);
or U2054 (N_2054,N_1583,N_1515);
nand U2055 (N_2055,N_1631,N_1809);
nor U2056 (N_2056,N_1738,N_1979);
and U2057 (N_2057,N_1821,N_1699);
or U2058 (N_2058,N_1692,N_1899);
or U2059 (N_2059,N_1710,N_1768);
xnor U2060 (N_2060,N_1694,N_1992);
nor U2061 (N_2061,N_1581,N_1588);
and U2062 (N_2062,N_1528,N_1997);
and U2063 (N_2063,N_1649,N_1675);
and U2064 (N_2064,N_1713,N_1943);
or U2065 (N_2065,N_1506,N_1634);
nand U2066 (N_2066,N_1907,N_1502);
nor U2067 (N_2067,N_1920,N_1884);
and U2068 (N_2068,N_1645,N_1782);
nor U2069 (N_2069,N_1696,N_1887);
and U2070 (N_2070,N_1564,N_1608);
nand U2071 (N_2071,N_1944,N_1552);
nand U2072 (N_2072,N_1655,N_1676);
xor U2073 (N_2073,N_1947,N_1657);
or U2074 (N_2074,N_1791,N_1591);
nor U2075 (N_2075,N_1966,N_1637);
or U2076 (N_2076,N_1987,N_1709);
or U2077 (N_2077,N_1951,N_1984);
nand U2078 (N_2078,N_1697,N_1806);
and U2079 (N_2079,N_1550,N_1642);
and U2080 (N_2080,N_1681,N_1939);
nor U2081 (N_2081,N_1587,N_1703);
nor U2082 (N_2082,N_1948,N_1946);
or U2083 (N_2083,N_1507,N_1671);
nand U2084 (N_2084,N_1663,N_1776);
nor U2085 (N_2085,N_1789,N_1508);
nand U2086 (N_2086,N_1644,N_1596);
or U2087 (N_2087,N_1902,N_1926);
and U2088 (N_2088,N_1921,N_1647);
xor U2089 (N_2089,N_1639,N_1680);
nor U2090 (N_2090,N_1717,N_1832);
nand U2091 (N_2091,N_1861,N_1995);
nand U2092 (N_2092,N_1766,N_1929);
and U2093 (N_2093,N_1545,N_1816);
or U2094 (N_2094,N_1886,N_1996);
nor U2095 (N_2095,N_1731,N_1863);
and U2096 (N_2096,N_1648,N_1855);
nor U2097 (N_2097,N_1733,N_1682);
and U2098 (N_2098,N_1895,N_1823);
or U2099 (N_2099,N_1769,N_1852);
and U2100 (N_2100,N_1745,N_1646);
and U2101 (N_2101,N_1879,N_1814);
nand U2102 (N_2102,N_1890,N_1749);
nor U2103 (N_2103,N_1569,N_1967);
xnor U2104 (N_2104,N_1985,N_1568);
nand U2105 (N_2105,N_1539,N_1662);
nor U2106 (N_2106,N_1641,N_1793);
nand U2107 (N_2107,N_1604,N_1541);
and U2108 (N_2108,N_1922,N_1805);
nand U2109 (N_2109,N_1600,N_1937);
and U2110 (N_2110,N_1872,N_1619);
nor U2111 (N_2111,N_1977,N_1548);
or U2112 (N_2112,N_1773,N_1511);
or U2113 (N_2113,N_1877,N_1889);
nand U2114 (N_2114,N_1695,N_1875);
or U2115 (N_2115,N_1754,N_1813);
nor U2116 (N_2116,N_1576,N_1565);
nor U2117 (N_2117,N_1536,N_1748);
nor U2118 (N_2118,N_1952,N_1537);
nand U2119 (N_2119,N_1559,N_1758);
nand U2120 (N_2120,N_1930,N_1730);
or U2121 (N_2121,N_1945,N_1931);
and U2122 (N_2122,N_1854,N_1743);
or U2123 (N_2123,N_1871,N_1828);
nor U2124 (N_2124,N_1771,N_1598);
nand U2125 (N_2125,N_1795,N_1983);
or U2126 (N_2126,N_1843,N_1856);
and U2127 (N_2127,N_1829,N_1794);
nor U2128 (N_2128,N_1653,N_1700);
nor U2129 (N_2129,N_1800,N_1531);
or U2130 (N_2130,N_1660,N_1734);
or U2131 (N_2131,N_1501,N_1963);
or U2132 (N_2132,N_1841,N_1741);
and U2133 (N_2133,N_1796,N_1858);
or U2134 (N_2134,N_1705,N_1810);
nor U2135 (N_2135,N_1954,N_1898);
or U2136 (N_2136,N_1740,N_1736);
or U2137 (N_2137,N_1956,N_1636);
nand U2138 (N_2138,N_1708,N_1933);
and U2139 (N_2139,N_1683,N_1595);
nor U2140 (N_2140,N_1757,N_1797);
and U2141 (N_2141,N_1812,N_1869);
and U2142 (N_2142,N_1751,N_1894);
nor U2143 (N_2143,N_1912,N_1991);
nor U2144 (N_2144,N_1914,N_1558);
and U2145 (N_2145,N_1744,N_1819);
nor U2146 (N_2146,N_1936,N_1688);
nand U2147 (N_2147,N_1989,N_1579);
nor U2148 (N_2148,N_1928,N_1772);
nand U2149 (N_2149,N_1747,N_1808);
nor U2150 (N_2150,N_1620,N_1562);
nand U2151 (N_2151,N_1897,N_1827);
or U2152 (N_2152,N_1891,N_1874);
nand U2153 (N_2153,N_1732,N_1862);
nor U2154 (N_2154,N_1950,N_1845);
or U2155 (N_2155,N_1627,N_1693);
and U2156 (N_2156,N_1880,N_1582);
and U2157 (N_2157,N_1790,N_1919);
nor U2158 (N_2158,N_1534,N_1704);
xor U2159 (N_2159,N_1574,N_1577);
or U2160 (N_2160,N_1935,N_1557);
or U2161 (N_2161,N_1690,N_1622);
and U2162 (N_2162,N_1725,N_1535);
nand U2163 (N_2163,N_1820,N_1885);
nor U2164 (N_2164,N_1962,N_1925);
nand U2165 (N_2165,N_1893,N_1529);
nor U2166 (N_2166,N_1714,N_1980);
nor U2167 (N_2167,N_1566,N_1553);
nor U2168 (N_2168,N_1594,N_1586);
nor U2169 (N_2169,N_1701,N_1777);
and U2170 (N_2170,N_1760,N_1727);
nor U2171 (N_2171,N_1590,N_1881);
nor U2172 (N_2172,N_1857,N_1527);
nand U2173 (N_2173,N_1850,N_1679);
or U2174 (N_2174,N_1818,N_1973);
and U2175 (N_2175,N_1673,N_1788);
and U2176 (N_2176,N_1575,N_1767);
and U2177 (N_2177,N_1968,N_1661);
nand U2178 (N_2178,N_1807,N_1822);
nand U2179 (N_2179,N_1867,N_1691);
and U2180 (N_2180,N_1722,N_1975);
nor U2181 (N_2181,N_1860,N_1833);
or U2182 (N_2182,N_1971,N_1512);
and U2183 (N_2183,N_1824,N_1610);
and U2184 (N_2184,N_1830,N_1972);
nor U2185 (N_2185,N_1864,N_1570);
or U2186 (N_2186,N_1753,N_1835);
nand U2187 (N_2187,N_1500,N_1629);
nand U2188 (N_2188,N_1940,N_1831);
nand U2189 (N_2189,N_1606,N_1518);
and U2190 (N_2190,N_1970,N_1801);
and U2191 (N_2191,N_1532,N_1517);
and U2192 (N_2192,N_1698,N_1853);
or U2193 (N_2193,N_1778,N_1611);
nand U2194 (N_2194,N_1556,N_1934);
nor U2195 (N_2195,N_1526,N_1593);
nor U2196 (N_2196,N_1533,N_1804);
or U2197 (N_2197,N_1712,N_1826);
nor U2198 (N_2198,N_1633,N_1685);
nand U2199 (N_2199,N_1787,N_1906);
and U2200 (N_2200,N_1905,N_1615);
or U2201 (N_2201,N_1865,N_1635);
nor U2202 (N_2202,N_1779,N_1916);
or U2203 (N_2203,N_1640,N_1628);
or U2204 (N_2204,N_1837,N_1560);
nand U2205 (N_2205,N_1998,N_1786);
or U2206 (N_2206,N_1668,N_1994);
or U2207 (N_2207,N_1614,N_1915);
and U2208 (N_2208,N_1763,N_1702);
and U2209 (N_2209,N_1609,N_1678);
and U2210 (N_2210,N_1616,N_1621);
or U2211 (N_2211,N_1924,N_1510);
nand U2212 (N_2212,N_1665,N_1868);
and U2213 (N_2213,N_1719,N_1811);
nand U2214 (N_2214,N_1911,N_1571);
and U2215 (N_2215,N_1774,N_1993);
or U2216 (N_2216,N_1513,N_1597);
or U2217 (N_2217,N_1917,N_1677);
xor U2218 (N_2218,N_1848,N_1949);
nand U2219 (N_2219,N_1999,N_1519);
nand U2220 (N_2220,N_1739,N_1838);
nor U2221 (N_2221,N_1958,N_1798);
nand U2222 (N_2222,N_1503,N_1684);
or U2223 (N_2223,N_1718,N_1981);
and U2224 (N_2224,N_1514,N_1667);
nor U2225 (N_2225,N_1603,N_1643);
and U2226 (N_2226,N_1960,N_1988);
and U2227 (N_2227,N_1986,N_1567);
and U2228 (N_2228,N_1589,N_1964);
nand U2229 (N_2229,N_1549,N_1551);
and U2230 (N_2230,N_1842,N_1866);
nor U2231 (N_2231,N_1941,N_1846);
and U2232 (N_2232,N_1859,N_1724);
or U2233 (N_2233,N_1605,N_1505);
or U2234 (N_2234,N_1764,N_1755);
and U2235 (N_2235,N_1530,N_1654);
nand U2236 (N_2236,N_1630,N_1521);
nor U2237 (N_2237,N_1873,N_1561);
xor U2238 (N_2238,N_1903,N_1540);
nor U2239 (N_2239,N_1544,N_1554);
or U2240 (N_2240,N_1825,N_1803);
nor U2241 (N_2241,N_1617,N_1509);
or U2242 (N_2242,N_1638,N_1650);
or U2243 (N_2243,N_1959,N_1666);
nor U2244 (N_2244,N_1836,N_1523);
nor U2245 (N_2245,N_1689,N_1976);
or U2246 (N_2246,N_1909,N_1674);
nor U2247 (N_2247,N_1592,N_1878);
or U2248 (N_2248,N_1538,N_1839);
or U2249 (N_2249,N_1932,N_1720);
or U2250 (N_2250,N_1671,N_1806);
nor U2251 (N_2251,N_1751,N_1968);
xor U2252 (N_2252,N_1544,N_1615);
nand U2253 (N_2253,N_1701,N_1943);
nor U2254 (N_2254,N_1938,N_1667);
xor U2255 (N_2255,N_1644,N_1783);
nand U2256 (N_2256,N_1915,N_1808);
and U2257 (N_2257,N_1916,N_1754);
nand U2258 (N_2258,N_1703,N_1889);
nand U2259 (N_2259,N_1940,N_1776);
nor U2260 (N_2260,N_1894,N_1867);
or U2261 (N_2261,N_1902,N_1546);
nor U2262 (N_2262,N_1721,N_1503);
xnor U2263 (N_2263,N_1597,N_1890);
and U2264 (N_2264,N_1796,N_1946);
nor U2265 (N_2265,N_1793,N_1961);
nor U2266 (N_2266,N_1556,N_1662);
and U2267 (N_2267,N_1649,N_1954);
or U2268 (N_2268,N_1647,N_1810);
nand U2269 (N_2269,N_1648,N_1519);
or U2270 (N_2270,N_1866,N_1992);
and U2271 (N_2271,N_1693,N_1968);
or U2272 (N_2272,N_1992,N_1775);
nand U2273 (N_2273,N_1957,N_1890);
and U2274 (N_2274,N_1904,N_1583);
nand U2275 (N_2275,N_1540,N_1625);
and U2276 (N_2276,N_1741,N_1755);
or U2277 (N_2277,N_1505,N_1518);
nand U2278 (N_2278,N_1764,N_1754);
nand U2279 (N_2279,N_1701,N_1651);
or U2280 (N_2280,N_1682,N_1535);
and U2281 (N_2281,N_1753,N_1938);
or U2282 (N_2282,N_1676,N_1992);
nor U2283 (N_2283,N_1638,N_1532);
nand U2284 (N_2284,N_1974,N_1723);
nor U2285 (N_2285,N_1858,N_1736);
or U2286 (N_2286,N_1816,N_1740);
nand U2287 (N_2287,N_1515,N_1834);
nor U2288 (N_2288,N_1548,N_1916);
nand U2289 (N_2289,N_1569,N_1932);
or U2290 (N_2290,N_1625,N_1707);
or U2291 (N_2291,N_1836,N_1539);
xnor U2292 (N_2292,N_1684,N_1679);
nand U2293 (N_2293,N_1897,N_1511);
nand U2294 (N_2294,N_1596,N_1875);
nand U2295 (N_2295,N_1821,N_1601);
xor U2296 (N_2296,N_1622,N_1599);
and U2297 (N_2297,N_1525,N_1557);
and U2298 (N_2298,N_1932,N_1925);
nand U2299 (N_2299,N_1602,N_1913);
nor U2300 (N_2300,N_1851,N_1761);
nand U2301 (N_2301,N_1760,N_1840);
and U2302 (N_2302,N_1704,N_1977);
nor U2303 (N_2303,N_1873,N_1741);
nand U2304 (N_2304,N_1753,N_1529);
nand U2305 (N_2305,N_1967,N_1955);
and U2306 (N_2306,N_1925,N_1750);
nand U2307 (N_2307,N_1686,N_1640);
nor U2308 (N_2308,N_1626,N_1698);
nor U2309 (N_2309,N_1910,N_1673);
nand U2310 (N_2310,N_1933,N_1822);
nor U2311 (N_2311,N_1833,N_1531);
nand U2312 (N_2312,N_1691,N_1510);
and U2313 (N_2313,N_1512,N_1747);
nor U2314 (N_2314,N_1805,N_1762);
or U2315 (N_2315,N_1913,N_1711);
and U2316 (N_2316,N_1991,N_1700);
or U2317 (N_2317,N_1737,N_1787);
nand U2318 (N_2318,N_1644,N_1815);
nand U2319 (N_2319,N_1725,N_1590);
nand U2320 (N_2320,N_1999,N_1643);
nor U2321 (N_2321,N_1788,N_1615);
nor U2322 (N_2322,N_1831,N_1713);
nand U2323 (N_2323,N_1523,N_1994);
and U2324 (N_2324,N_1702,N_1876);
nor U2325 (N_2325,N_1688,N_1729);
or U2326 (N_2326,N_1616,N_1581);
or U2327 (N_2327,N_1859,N_1955);
or U2328 (N_2328,N_1559,N_1647);
xor U2329 (N_2329,N_1814,N_1564);
and U2330 (N_2330,N_1518,N_1972);
or U2331 (N_2331,N_1597,N_1964);
nand U2332 (N_2332,N_1991,N_1825);
xor U2333 (N_2333,N_1642,N_1639);
nand U2334 (N_2334,N_1600,N_1547);
nand U2335 (N_2335,N_1540,N_1910);
nand U2336 (N_2336,N_1684,N_1694);
or U2337 (N_2337,N_1920,N_1552);
or U2338 (N_2338,N_1640,N_1631);
or U2339 (N_2339,N_1907,N_1522);
or U2340 (N_2340,N_1886,N_1564);
or U2341 (N_2341,N_1983,N_1917);
xnor U2342 (N_2342,N_1508,N_1612);
and U2343 (N_2343,N_1852,N_1579);
nand U2344 (N_2344,N_1823,N_1598);
or U2345 (N_2345,N_1869,N_1690);
and U2346 (N_2346,N_1703,N_1831);
nand U2347 (N_2347,N_1503,N_1834);
nor U2348 (N_2348,N_1994,N_1705);
nor U2349 (N_2349,N_1999,N_1685);
and U2350 (N_2350,N_1593,N_1718);
nor U2351 (N_2351,N_1914,N_1864);
nand U2352 (N_2352,N_1889,N_1774);
xor U2353 (N_2353,N_1948,N_1622);
and U2354 (N_2354,N_1740,N_1598);
nand U2355 (N_2355,N_1841,N_1778);
and U2356 (N_2356,N_1918,N_1703);
and U2357 (N_2357,N_1516,N_1858);
and U2358 (N_2358,N_1720,N_1939);
nand U2359 (N_2359,N_1502,N_1969);
and U2360 (N_2360,N_1619,N_1618);
nor U2361 (N_2361,N_1934,N_1557);
nand U2362 (N_2362,N_1594,N_1632);
nand U2363 (N_2363,N_1824,N_1636);
nand U2364 (N_2364,N_1619,N_1696);
and U2365 (N_2365,N_1590,N_1866);
nor U2366 (N_2366,N_1572,N_1946);
nand U2367 (N_2367,N_1818,N_1613);
or U2368 (N_2368,N_1543,N_1578);
nand U2369 (N_2369,N_1586,N_1678);
and U2370 (N_2370,N_1960,N_1621);
nand U2371 (N_2371,N_1949,N_1906);
xor U2372 (N_2372,N_1779,N_1935);
or U2373 (N_2373,N_1749,N_1898);
nor U2374 (N_2374,N_1976,N_1903);
or U2375 (N_2375,N_1722,N_1673);
or U2376 (N_2376,N_1686,N_1529);
and U2377 (N_2377,N_1887,N_1991);
nand U2378 (N_2378,N_1942,N_1701);
nand U2379 (N_2379,N_1557,N_1836);
or U2380 (N_2380,N_1874,N_1695);
and U2381 (N_2381,N_1848,N_1549);
and U2382 (N_2382,N_1669,N_1757);
or U2383 (N_2383,N_1894,N_1860);
nor U2384 (N_2384,N_1947,N_1615);
or U2385 (N_2385,N_1779,N_1690);
or U2386 (N_2386,N_1975,N_1524);
nor U2387 (N_2387,N_1523,N_1652);
nor U2388 (N_2388,N_1652,N_1751);
xnor U2389 (N_2389,N_1933,N_1724);
and U2390 (N_2390,N_1530,N_1569);
and U2391 (N_2391,N_1868,N_1713);
nand U2392 (N_2392,N_1912,N_1679);
nand U2393 (N_2393,N_1633,N_1544);
or U2394 (N_2394,N_1836,N_1689);
or U2395 (N_2395,N_1742,N_1990);
or U2396 (N_2396,N_1722,N_1610);
nand U2397 (N_2397,N_1741,N_1977);
nand U2398 (N_2398,N_1537,N_1535);
and U2399 (N_2399,N_1644,N_1587);
nand U2400 (N_2400,N_1880,N_1735);
nand U2401 (N_2401,N_1777,N_1757);
or U2402 (N_2402,N_1717,N_1966);
nand U2403 (N_2403,N_1719,N_1845);
or U2404 (N_2404,N_1847,N_1918);
nand U2405 (N_2405,N_1693,N_1971);
and U2406 (N_2406,N_1741,N_1653);
nand U2407 (N_2407,N_1972,N_1913);
and U2408 (N_2408,N_1813,N_1636);
nand U2409 (N_2409,N_1982,N_1579);
nor U2410 (N_2410,N_1905,N_1983);
and U2411 (N_2411,N_1642,N_1536);
nor U2412 (N_2412,N_1707,N_1939);
or U2413 (N_2413,N_1604,N_1686);
nand U2414 (N_2414,N_1930,N_1938);
or U2415 (N_2415,N_1948,N_1760);
and U2416 (N_2416,N_1886,N_1933);
nand U2417 (N_2417,N_1551,N_1657);
and U2418 (N_2418,N_1659,N_1664);
xnor U2419 (N_2419,N_1561,N_1669);
or U2420 (N_2420,N_1707,N_1979);
nand U2421 (N_2421,N_1981,N_1729);
or U2422 (N_2422,N_1903,N_1595);
nand U2423 (N_2423,N_1705,N_1884);
or U2424 (N_2424,N_1811,N_1622);
or U2425 (N_2425,N_1705,N_1632);
and U2426 (N_2426,N_1523,N_1634);
nand U2427 (N_2427,N_1568,N_1816);
nor U2428 (N_2428,N_1947,N_1835);
or U2429 (N_2429,N_1949,N_1965);
nor U2430 (N_2430,N_1792,N_1990);
nor U2431 (N_2431,N_1815,N_1563);
and U2432 (N_2432,N_1942,N_1714);
nand U2433 (N_2433,N_1705,N_1965);
or U2434 (N_2434,N_1593,N_1994);
or U2435 (N_2435,N_1891,N_1832);
and U2436 (N_2436,N_1709,N_1785);
or U2437 (N_2437,N_1964,N_1622);
nand U2438 (N_2438,N_1805,N_1780);
and U2439 (N_2439,N_1677,N_1630);
and U2440 (N_2440,N_1768,N_1922);
nor U2441 (N_2441,N_1712,N_1857);
or U2442 (N_2442,N_1610,N_1772);
nor U2443 (N_2443,N_1763,N_1879);
and U2444 (N_2444,N_1653,N_1715);
and U2445 (N_2445,N_1926,N_1647);
nand U2446 (N_2446,N_1591,N_1518);
nand U2447 (N_2447,N_1630,N_1764);
or U2448 (N_2448,N_1586,N_1756);
nand U2449 (N_2449,N_1578,N_1778);
nor U2450 (N_2450,N_1679,N_1943);
nand U2451 (N_2451,N_1875,N_1893);
or U2452 (N_2452,N_1659,N_1898);
or U2453 (N_2453,N_1918,N_1518);
nand U2454 (N_2454,N_1965,N_1590);
nand U2455 (N_2455,N_1742,N_1818);
and U2456 (N_2456,N_1666,N_1844);
and U2457 (N_2457,N_1602,N_1932);
or U2458 (N_2458,N_1848,N_1901);
and U2459 (N_2459,N_1511,N_1776);
or U2460 (N_2460,N_1744,N_1986);
xor U2461 (N_2461,N_1764,N_1769);
and U2462 (N_2462,N_1749,N_1742);
or U2463 (N_2463,N_1838,N_1554);
nor U2464 (N_2464,N_1911,N_1860);
and U2465 (N_2465,N_1662,N_1599);
nor U2466 (N_2466,N_1617,N_1651);
nor U2467 (N_2467,N_1516,N_1844);
nor U2468 (N_2468,N_1515,N_1652);
nor U2469 (N_2469,N_1847,N_1595);
nand U2470 (N_2470,N_1549,N_1999);
nor U2471 (N_2471,N_1989,N_1848);
and U2472 (N_2472,N_1763,N_1789);
nor U2473 (N_2473,N_1775,N_1875);
or U2474 (N_2474,N_1748,N_1611);
or U2475 (N_2475,N_1734,N_1860);
and U2476 (N_2476,N_1771,N_1889);
nor U2477 (N_2477,N_1935,N_1737);
nor U2478 (N_2478,N_1732,N_1846);
nand U2479 (N_2479,N_1960,N_1806);
or U2480 (N_2480,N_1706,N_1974);
and U2481 (N_2481,N_1993,N_1933);
nand U2482 (N_2482,N_1920,N_1614);
and U2483 (N_2483,N_1673,N_1882);
nand U2484 (N_2484,N_1771,N_1593);
nand U2485 (N_2485,N_1901,N_1853);
or U2486 (N_2486,N_1847,N_1657);
and U2487 (N_2487,N_1849,N_1816);
and U2488 (N_2488,N_1808,N_1694);
nand U2489 (N_2489,N_1668,N_1847);
or U2490 (N_2490,N_1560,N_1887);
nor U2491 (N_2491,N_1555,N_1941);
nand U2492 (N_2492,N_1713,N_1974);
nor U2493 (N_2493,N_1556,N_1910);
or U2494 (N_2494,N_1610,N_1541);
and U2495 (N_2495,N_1810,N_1645);
nor U2496 (N_2496,N_1880,N_1729);
nor U2497 (N_2497,N_1564,N_1803);
and U2498 (N_2498,N_1944,N_1960);
nor U2499 (N_2499,N_1558,N_1659);
or U2500 (N_2500,N_2499,N_2455);
xor U2501 (N_2501,N_2182,N_2129);
nor U2502 (N_2502,N_2336,N_2193);
nor U2503 (N_2503,N_2364,N_2253);
or U2504 (N_2504,N_2376,N_2196);
or U2505 (N_2505,N_2289,N_2201);
or U2506 (N_2506,N_2489,N_2218);
and U2507 (N_2507,N_2103,N_2297);
nand U2508 (N_2508,N_2255,N_2216);
or U2509 (N_2509,N_2144,N_2473);
xnor U2510 (N_2510,N_2314,N_2279);
or U2511 (N_2511,N_2340,N_2256);
or U2512 (N_2512,N_2323,N_2269);
and U2513 (N_2513,N_2322,N_2342);
or U2514 (N_2514,N_2185,N_2292);
xnor U2515 (N_2515,N_2210,N_2331);
nor U2516 (N_2516,N_2385,N_2449);
nor U2517 (N_2517,N_2397,N_2059);
nand U2518 (N_2518,N_2258,N_2001);
nor U2519 (N_2519,N_2360,N_2410);
nor U2520 (N_2520,N_2174,N_2171);
nand U2521 (N_2521,N_2147,N_2306);
or U2522 (N_2522,N_2157,N_2008);
and U2523 (N_2523,N_2183,N_2444);
and U2524 (N_2524,N_2353,N_2142);
or U2525 (N_2525,N_2075,N_2354);
and U2526 (N_2526,N_2112,N_2398);
nand U2527 (N_2527,N_2486,N_2382);
nand U2528 (N_2528,N_2022,N_2287);
nand U2529 (N_2529,N_2180,N_2457);
xor U2530 (N_2530,N_2346,N_2370);
nand U2531 (N_2531,N_2214,N_2295);
and U2532 (N_2532,N_2320,N_2321);
and U2533 (N_2533,N_2053,N_2260);
nand U2534 (N_2534,N_2245,N_2036);
or U2535 (N_2535,N_2371,N_2395);
or U2536 (N_2536,N_2073,N_2149);
nor U2537 (N_2537,N_2386,N_2278);
nand U2538 (N_2538,N_2220,N_2367);
or U2539 (N_2539,N_2337,N_2143);
nand U2540 (N_2540,N_2072,N_2126);
and U2541 (N_2541,N_2019,N_2023);
nand U2542 (N_2542,N_2136,N_2389);
and U2543 (N_2543,N_2078,N_2105);
nand U2544 (N_2544,N_2421,N_2135);
and U2545 (N_2545,N_2328,N_2197);
or U2546 (N_2546,N_2474,N_2497);
and U2547 (N_2547,N_2282,N_2228);
nand U2548 (N_2548,N_2217,N_2261);
nand U2549 (N_2549,N_2424,N_2044);
and U2550 (N_2550,N_2130,N_2158);
nor U2551 (N_2551,N_2037,N_2338);
and U2552 (N_2552,N_2264,N_2071);
or U2553 (N_2553,N_2451,N_2358);
nor U2554 (N_2554,N_2178,N_2476);
nor U2555 (N_2555,N_2368,N_2191);
and U2556 (N_2556,N_2408,N_2088);
or U2557 (N_2557,N_2361,N_2453);
nand U2558 (N_2558,N_2239,N_2039);
xnor U2559 (N_2559,N_2265,N_2280);
and U2560 (N_2560,N_2042,N_2000);
nand U2561 (N_2561,N_2168,N_2091);
and U2562 (N_2562,N_2082,N_2485);
and U2563 (N_2563,N_2004,N_2288);
nand U2564 (N_2564,N_2428,N_2468);
xor U2565 (N_2565,N_2035,N_2469);
nand U2566 (N_2566,N_2263,N_2415);
and U2567 (N_2567,N_2167,N_2335);
nor U2568 (N_2568,N_2325,N_2043);
xor U2569 (N_2569,N_2475,N_2404);
and U2570 (N_2570,N_2401,N_2419);
nor U2571 (N_2571,N_2271,N_2111);
nor U2572 (N_2572,N_2118,N_2387);
xnor U2573 (N_2573,N_2057,N_2454);
or U2574 (N_2574,N_2466,N_2285);
or U2575 (N_2575,N_2231,N_2006);
or U2576 (N_2576,N_2206,N_2181);
or U2577 (N_2577,N_2267,N_2133);
nor U2578 (N_2578,N_2281,N_2391);
nor U2579 (N_2579,N_2259,N_2430);
or U2580 (N_2580,N_2127,N_2249);
nand U2581 (N_2581,N_2375,N_2162);
or U2582 (N_2582,N_2076,N_2140);
or U2583 (N_2583,N_2450,N_2313);
nor U2584 (N_2584,N_2377,N_2029);
nor U2585 (N_2585,N_2123,N_2380);
and U2586 (N_2586,N_2479,N_2352);
or U2587 (N_2587,N_2283,N_2032);
nor U2588 (N_2588,N_2002,N_2341);
or U2589 (N_2589,N_2339,N_2012);
nand U2590 (N_2590,N_2190,N_2117);
or U2591 (N_2591,N_2212,N_2242);
and U2592 (N_2592,N_2384,N_2429);
nor U2593 (N_2593,N_2199,N_2120);
and U2594 (N_2594,N_2366,N_2363);
nor U2595 (N_2595,N_2495,N_2477);
nand U2596 (N_2596,N_2134,N_2308);
and U2597 (N_2597,N_2095,N_2422);
nand U2598 (N_2598,N_2262,N_2173);
nor U2599 (N_2599,N_2176,N_2194);
nor U2600 (N_2600,N_2471,N_2431);
nor U2601 (N_2601,N_2009,N_2392);
or U2602 (N_2602,N_2491,N_2296);
or U2603 (N_2603,N_2251,N_2356);
or U2604 (N_2604,N_2152,N_2060);
or U2605 (N_2605,N_2324,N_2309);
or U2606 (N_2606,N_2452,N_2319);
or U2607 (N_2607,N_2165,N_2205);
and U2608 (N_2608,N_2304,N_2318);
or U2609 (N_2609,N_2438,N_2098);
nand U2610 (N_2610,N_2050,N_2014);
nor U2611 (N_2611,N_2099,N_2235);
and U2612 (N_2612,N_2104,N_2225);
or U2613 (N_2613,N_2403,N_2224);
or U2614 (N_2614,N_2092,N_2423);
nand U2615 (N_2615,N_2040,N_2482);
and U2616 (N_2616,N_2139,N_2492);
or U2617 (N_2617,N_2277,N_2274);
or U2618 (N_2618,N_2232,N_2124);
xor U2619 (N_2619,N_2478,N_2378);
nor U2620 (N_2620,N_2446,N_2122);
or U2621 (N_2621,N_2222,N_2275);
and U2622 (N_2622,N_2412,N_2350);
nor U2623 (N_2623,N_2458,N_2192);
nand U2624 (N_2624,N_2464,N_2100);
nand U2625 (N_2625,N_2425,N_2238);
nand U2626 (N_2626,N_2327,N_2445);
nor U2627 (N_2627,N_2187,N_2399);
nor U2628 (N_2628,N_2204,N_2393);
or U2629 (N_2629,N_2208,N_2219);
and U2630 (N_2630,N_2163,N_2400);
nor U2631 (N_2631,N_2286,N_2065);
and U2632 (N_2632,N_2020,N_2443);
nor U2633 (N_2633,N_2317,N_2198);
nand U2634 (N_2634,N_2487,N_2433);
and U2635 (N_2635,N_2115,N_2200);
nor U2636 (N_2636,N_2013,N_2357);
nand U2637 (N_2637,N_2347,N_2155);
and U2638 (N_2638,N_2034,N_2442);
or U2639 (N_2639,N_2237,N_2330);
nor U2640 (N_2640,N_2097,N_2113);
and U2641 (N_2641,N_2298,N_2148);
or U2642 (N_2642,N_2017,N_2435);
or U2643 (N_2643,N_2186,N_2329);
nor U2644 (N_2644,N_2077,N_2164);
and U2645 (N_2645,N_2064,N_2085);
nand U2646 (N_2646,N_2247,N_2426);
nor U2647 (N_2647,N_2069,N_2343);
or U2648 (N_2648,N_2021,N_2015);
nand U2649 (N_2649,N_2351,N_2096);
nand U2650 (N_2650,N_2244,N_2373);
and U2651 (N_2651,N_2405,N_2272);
or U2652 (N_2652,N_2153,N_2056);
or U2653 (N_2653,N_2101,N_2303);
nor U2654 (N_2654,N_2418,N_2106);
nand U2655 (N_2655,N_2307,N_2240);
nand U2656 (N_2656,N_2390,N_2062);
nor U2657 (N_2657,N_2349,N_2290);
nor U2658 (N_2658,N_2055,N_2388);
or U2659 (N_2659,N_2081,N_2243);
and U2660 (N_2660,N_2299,N_2334);
nand U2661 (N_2661,N_2131,N_2047);
or U2662 (N_2662,N_2052,N_2114);
nand U2663 (N_2663,N_2102,N_2417);
and U2664 (N_2664,N_2496,N_2276);
or U2665 (N_2665,N_2160,N_2437);
nand U2666 (N_2666,N_2010,N_2344);
xor U2667 (N_2667,N_2456,N_2179);
and U2668 (N_2668,N_2137,N_2250);
and U2669 (N_2669,N_2223,N_2470);
and U2670 (N_2670,N_2362,N_2432);
and U2671 (N_2671,N_2301,N_2484);
nor U2672 (N_2672,N_2480,N_2046);
and U2673 (N_2673,N_2156,N_2440);
nor U2674 (N_2674,N_2159,N_2058);
nand U2675 (N_2675,N_2184,N_2436);
or U2676 (N_2676,N_2266,N_2049);
nor U2677 (N_2677,N_2402,N_2414);
nor U2678 (N_2678,N_2302,N_2170);
nor U2679 (N_2679,N_2086,N_2005);
or U2680 (N_2680,N_2316,N_2119);
nand U2681 (N_2681,N_2026,N_2121);
and U2682 (N_2682,N_2448,N_2093);
nand U2683 (N_2683,N_2300,N_2166);
or U2684 (N_2684,N_2061,N_2369);
or U2685 (N_2685,N_2333,N_2236);
nand U2686 (N_2686,N_2063,N_2483);
and U2687 (N_2687,N_2409,N_2125);
and U2688 (N_2688,N_2359,N_2145);
or U2689 (N_2689,N_2411,N_2230);
nand U2690 (N_2690,N_2463,N_2177);
nor U2691 (N_2691,N_2268,N_2203);
and U2692 (N_2692,N_2248,N_2284);
nor U2693 (N_2693,N_2355,N_2080);
nor U2694 (N_2694,N_2209,N_2107);
and U2695 (N_2695,N_2427,N_2447);
nor U2696 (N_2696,N_2233,N_2045);
xnor U2697 (N_2697,N_2054,N_2068);
nor U2698 (N_2698,N_2493,N_2048);
nor U2699 (N_2699,N_2490,N_2345);
nand U2700 (N_2700,N_2024,N_2221);
nor U2701 (N_2701,N_2089,N_2332);
and U2702 (N_2702,N_2270,N_2465);
or U2703 (N_2703,N_2215,N_2472);
nand U2704 (N_2704,N_2348,N_2372);
nor U2705 (N_2705,N_2406,N_2202);
nor U2706 (N_2706,N_2027,N_2146);
nand U2707 (N_2707,N_2041,N_2003);
and U2708 (N_2708,N_2273,N_2108);
and U2709 (N_2709,N_2383,N_2257);
or U2710 (N_2710,N_2213,N_2151);
xnor U2711 (N_2711,N_2407,N_2462);
nand U2712 (N_2712,N_2488,N_2420);
nor U2713 (N_2713,N_2326,N_2116);
or U2714 (N_2714,N_2441,N_2413);
and U2715 (N_2715,N_2211,N_2312);
nand U2716 (N_2716,N_2459,N_2311);
nand U2717 (N_2717,N_2460,N_2067);
nand U2718 (N_2718,N_2132,N_2439);
or U2719 (N_2719,N_2234,N_2090);
and U2720 (N_2720,N_2074,N_2154);
nor U2721 (N_2721,N_2207,N_2246);
or U2722 (N_2722,N_2038,N_2379);
or U2723 (N_2723,N_2481,N_2087);
nand U2724 (N_2724,N_2018,N_2229);
or U2725 (N_2725,N_2051,N_2305);
and U2726 (N_2726,N_2195,N_2365);
or U2727 (N_2727,N_2161,N_2252);
xnor U2728 (N_2728,N_2011,N_2241);
or U2729 (N_2729,N_2189,N_2381);
nand U2730 (N_2730,N_2374,N_2310);
nor U2731 (N_2731,N_2188,N_2110);
and U2732 (N_2732,N_2070,N_2227);
and U2733 (N_2733,N_2394,N_2138);
nor U2734 (N_2734,N_2294,N_2254);
nand U2735 (N_2735,N_2094,N_2128);
and U2736 (N_2736,N_2175,N_2109);
nor U2737 (N_2737,N_2169,N_2172);
and U2738 (N_2738,N_2007,N_2025);
nand U2739 (N_2739,N_2461,N_2396);
nor U2740 (N_2740,N_2028,N_2033);
nor U2741 (N_2741,N_2150,N_2494);
or U2742 (N_2742,N_2141,N_2066);
xor U2743 (N_2743,N_2030,N_2291);
nand U2744 (N_2744,N_2434,N_2498);
or U2745 (N_2745,N_2416,N_2226);
or U2746 (N_2746,N_2031,N_2315);
xnor U2747 (N_2747,N_2016,N_2083);
nand U2748 (N_2748,N_2467,N_2084);
or U2749 (N_2749,N_2079,N_2293);
nor U2750 (N_2750,N_2483,N_2035);
nor U2751 (N_2751,N_2025,N_2454);
or U2752 (N_2752,N_2426,N_2411);
nor U2753 (N_2753,N_2338,N_2444);
nor U2754 (N_2754,N_2076,N_2467);
or U2755 (N_2755,N_2022,N_2111);
or U2756 (N_2756,N_2228,N_2268);
nor U2757 (N_2757,N_2209,N_2015);
xor U2758 (N_2758,N_2026,N_2029);
nand U2759 (N_2759,N_2076,N_2488);
nor U2760 (N_2760,N_2042,N_2184);
nor U2761 (N_2761,N_2326,N_2449);
nor U2762 (N_2762,N_2364,N_2130);
and U2763 (N_2763,N_2474,N_2388);
or U2764 (N_2764,N_2069,N_2113);
and U2765 (N_2765,N_2300,N_2020);
or U2766 (N_2766,N_2411,N_2169);
xor U2767 (N_2767,N_2348,N_2274);
and U2768 (N_2768,N_2470,N_2374);
xor U2769 (N_2769,N_2122,N_2466);
or U2770 (N_2770,N_2390,N_2034);
nand U2771 (N_2771,N_2118,N_2249);
nand U2772 (N_2772,N_2079,N_2217);
and U2773 (N_2773,N_2438,N_2039);
nor U2774 (N_2774,N_2154,N_2387);
nor U2775 (N_2775,N_2167,N_2313);
and U2776 (N_2776,N_2057,N_2470);
nor U2777 (N_2777,N_2036,N_2113);
nand U2778 (N_2778,N_2155,N_2011);
and U2779 (N_2779,N_2205,N_2443);
nand U2780 (N_2780,N_2294,N_2278);
nand U2781 (N_2781,N_2336,N_2188);
or U2782 (N_2782,N_2381,N_2035);
and U2783 (N_2783,N_2490,N_2237);
nor U2784 (N_2784,N_2474,N_2465);
nor U2785 (N_2785,N_2274,N_2244);
nor U2786 (N_2786,N_2286,N_2430);
and U2787 (N_2787,N_2082,N_2387);
nor U2788 (N_2788,N_2094,N_2206);
xor U2789 (N_2789,N_2446,N_2321);
and U2790 (N_2790,N_2206,N_2463);
or U2791 (N_2791,N_2065,N_2236);
and U2792 (N_2792,N_2370,N_2057);
xnor U2793 (N_2793,N_2062,N_2491);
and U2794 (N_2794,N_2488,N_2434);
and U2795 (N_2795,N_2214,N_2320);
nand U2796 (N_2796,N_2196,N_2379);
and U2797 (N_2797,N_2440,N_2414);
or U2798 (N_2798,N_2037,N_2079);
nor U2799 (N_2799,N_2292,N_2295);
nand U2800 (N_2800,N_2493,N_2106);
nand U2801 (N_2801,N_2292,N_2283);
nor U2802 (N_2802,N_2261,N_2054);
and U2803 (N_2803,N_2366,N_2038);
or U2804 (N_2804,N_2368,N_2371);
or U2805 (N_2805,N_2349,N_2300);
nor U2806 (N_2806,N_2000,N_2393);
and U2807 (N_2807,N_2101,N_2097);
nand U2808 (N_2808,N_2014,N_2108);
nor U2809 (N_2809,N_2383,N_2476);
nor U2810 (N_2810,N_2498,N_2411);
or U2811 (N_2811,N_2115,N_2297);
nor U2812 (N_2812,N_2365,N_2445);
and U2813 (N_2813,N_2085,N_2024);
or U2814 (N_2814,N_2477,N_2438);
or U2815 (N_2815,N_2387,N_2259);
nand U2816 (N_2816,N_2318,N_2019);
and U2817 (N_2817,N_2054,N_2327);
or U2818 (N_2818,N_2242,N_2240);
or U2819 (N_2819,N_2384,N_2303);
or U2820 (N_2820,N_2291,N_2153);
nand U2821 (N_2821,N_2203,N_2325);
and U2822 (N_2822,N_2275,N_2303);
or U2823 (N_2823,N_2083,N_2113);
nor U2824 (N_2824,N_2443,N_2481);
xnor U2825 (N_2825,N_2449,N_2090);
and U2826 (N_2826,N_2370,N_2153);
and U2827 (N_2827,N_2019,N_2411);
nand U2828 (N_2828,N_2188,N_2455);
or U2829 (N_2829,N_2041,N_2257);
or U2830 (N_2830,N_2299,N_2482);
and U2831 (N_2831,N_2069,N_2061);
nor U2832 (N_2832,N_2066,N_2421);
or U2833 (N_2833,N_2071,N_2379);
nand U2834 (N_2834,N_2219,N_2416);
or U2835 (N_2835,N_2291,N_2330);
and U2836 (N_2836,N_2472,N_2143);
nand U2837 (N_2837,N_2356,N_2009);
nand U2838 (N_2838,N_2422,N_2466);
nand U2839 (N_2839,N_2253,N_2002);
nor U2840 (N_2840,N_2395,N_2461);
nor U2841 (N_2841,N_2476,N_2067);
xnor U2842 (N_2842,N_2406,N_2180);
nand U2843 (N_2843,N_2499,N_2039);
nor U2844 (N_2844,N_2227,N_2397);
nand U2845 (N_2845,N_2089,N_2017);
and U2846 (N_2846,N_2093,N_2426);
and U2847 (N_2847,N_2474,N_2054);
or U2848 (N_2848,N_2393,N_2301);
and U2849 (N_2849,N_2152,N_2161);
nor U2850 (N_2850,N_2403,N_2391);
or U2851 (N_2851,N_2070,N_2278);
nand U2852 (N_2852,N_2418,N_2207);
and U2853 (N_2853,N_2249,N_2130);
nor U2854 (N_2854,N_2226,N_2020);
nor U2855 (N_2855,N_2013,N_2233);
nor U2856 (N_2856,N_2150,N_2255);
or U2857 (N_2857,N_2177,N_2349);
nand U2858 (N_2858,N_2358,N_2242);
nand U2859 (N_2859,N_2191,N_2097);
xnor U2860 (N_2860,N_2312,N_2459);
and U2861 (N_2861,N_2412,N_2422);
nor U2862 (N_2862,N_2256,N_2111);
nor U2863 (N_2863,N_2156,N_2289);
nand U2864 (N_2864,N_2417,N_2114);
and U2865 (N_2865,N_2061,N_2094);
or U2866 (N_2866,N_2220,N_2075);
nand U2867 (N_2867,N_2410,N_2180);
xor U2868 (N_2868,N_2183,N_2202);
or U2869 (N_2869,N_2245,N_2321);
nor U2870 (N_2870,N_2381,N_2026);
or U2871 (N_2871,N_2152,N_2413);
or U2872 (N_2872,N_2295,N_2098);
xnor U2873 (N_2873,N_2276,N_2148);
and U2874 (N_2874,N_2022,N_2367);
or U2875 (N_2875,N_2417,N_2088);
nand U2876 (N_2876,N_2463,N_2244);
or U2877 (N_2877,N_2450,N_2162);
and U2878 (N_2878,N_2040,N_2276);
or U2879 (N_2879,N_2125,N_2350);
xnor U2880 (N_2880,N_2137,N_2117);
nand U2881 (N_2881,N_2179,N_2430);
or U2882 (N_2882,N_2384,N_2431);
nand U2883 (N_2883,N_2065,N_2201);
or U2884 (N_2884,N_2185,N_2024);
and U2885 (N_2885,N_2411,N_2078);
nor U2886 (N_2886,N_2045,N_2188);
or U2887 (N_2887,N_2445,N_2393);
nand U2888 (N_2888,N_2235,N_2278);
or U2889 (N_2889,N_2387,N_2226);
or U2890 (N_2890,N_2145,N_2055);
or U2891 (N_2891,N_2373,N_2174);
nor U2892 (N_2892,N_2188,N_2124);
or U2893 (N_2893,N_2038,N_2136);
nand U2894 (N_2894,N_2025,N_2090);
nand U2895 (N_2895,N_2481,N_2206);
nand U2896 (N_2896,N_2338,N_2038);
or U2897 (N_2897,N_2056,N_2163);
or U2898 (N_2898,N_2405,N_2330);
and U2899 (N_2899,N_2307,N_2089);
nand U2900 (N_2900,N_2213,N_2338);
and U2901 (N_2901,N_2482,N_2063);
nor U2902 (N_2902,N_2493,N_2126);
nand U2903 (N_2903,N_2353,N_2024);
nand U2904 (N_2904,N_2389,N_2409);
nand U2905 (N_2905,N_2079,N_2077);
nand U2906 (N_2906,N_2364,N_2019);
nand U2907 (N_2907,N_2145,N_2159);
or U2908 (N_2908,N_2075,N_2290);
nor U2909 (N_2909,N_2416,N_2047);
nand U2910 (N_2910,N_2241,N_2463);
nor U2911 (N_2911,N_2069,N_2374);
or U2912 (N_2912,N_2390,N_2064);
nand U2913 (N_2913,N_2132,N_2427);
nand U2914 (N_2914,N_2382,N_2187);
or U2915 (N_2915,N_2414,N_2282);
and U2916 (N_2916,N_2317,N_2034);
nor U2917 (N_2917,N_2466,N_2114);
nand U2918 (N_2918,N_2318,N_2475);
and U2919 (N_2919,N_2038,N_2290);
nor U2920 (N_2920,N_2390,N_2375);
or U2921 (N_2921,N_2008,N_2009);
nor U2922 (N_2922,N_2139,N_2443);
nand U2923 (N_2923,N_2104,N_2349);
and U2924 (N_2924,N_2156,N_2406);
nor U2925 (N_2925,N_2160,N_2058);
and U2926 (N_2926,N_2181,N_2255);
or U2927 (N_2927,N_2084,N_2332);
nor U2928 (N_2928,N_2340,N_2275);
or U2929 (N_2929,N_2440,N_2024);
or U2930 (N_2930,N_2481,N_2112);
and U2931 (N_2931,N_2354,N_2198);
nor U2932 (N_2932,N_2036,N_2491);
nor U2933 (N_2933,N_2275,N_2288);
and U2934 (N_2934,N_2417,N_2098);
nand U2935 (N_2935,N_2352,N_2011);
and U2936 (N_2936,N_2319,N_2316);
and U2937 (N_2937,N_2345,N_2407);
nand U2938 (N_2938,N_2255,N_2424);
nor U2939 (N_2939,N_2439,N_2483);
and U2940 (N_2940,N_2117,N_2254);
and U2941 (N_2941,N_2474,N_2125);
nor U2942 (N_2942,N_2488,N_2448);
nand U2943 (N_2943,N_2473,N_2226);
nor U2944 (N_2944,N_2352,N_2159);
nor U2945 (N_2945,N_2303,N_2402);
nor U2946 (N_2946,N_2132,N_2370);
or U2947 (N_2947,N_2084,N_2219);
and U2948 (N_2948,N_2007,N_2450);
nor U2949 (N_2949,N_2001,N_2325);
nand U2950 (N_2950,N_2065,N_2396);
nor U2951 (N_2951,N_2242,N_2257);
or U2952 (N_2952,N_2014,N_2022);
nand U2953 (N_2953,N_2234,N_2190);
nand U2954 (N_2954,N_2005,N_2105);
nand U2955 (N_2955,N_2456,N_2098);
or U2956 (N_2956,N_2357,N_2152);
nand U2957 (N_2957,N_2354,N_2009);
and U2958 (N_2958,N_2378,N_2222);
nand U2959 (N_2959,N_2118,N_2417);
and U2960 (N_2960,N_2437,N_2050);
or U2961 (N_2961,N_2126,N_2343);
or U2962 (N_2962,N_2002,N_2456);
nand U2963 (N_2963,N_2014,N_2337);
or U2964 (N_2964,N_2105,N_2053);
nor U2965 (N_2965,N_2375,N_2408);
xor U2966 (N_2966,N_2135,N_2252);
nand U2967 (N_2967,N_2148,N_2092);
nand U2968 (N_2968,N_2331,N_2168);
nor U2969 (N_2969,N_2016,N_2444);
nand U2970 (N_2970,N_2416,N_2003);
nor U2971 (N_2971,N_2488,N_2056);
xor U2972 (N_2972,N_2177,N_2008);
and U2973 (N_2973,N_2264,N_2079);
nor U2974 (N_2974,N_2260,N_2102);
or U2975 (N_2975,N_2086,N_2360);
or U2976 (N_2976,N_2445,N_2234);
and U2977 (N_2977,N_2087,N_2237);
nor U2978 (N_2978,N_2488,N_2157);
nor U2979 (N_2979,N_2412,N_2170);
or U2980 (N_2980,N_2158,N_2461);
nor U2981 (N_2981,N_2040,N_2449);
nand U2982 (N_2982,N_2355,N_2449);
nand U2983 (N_2983,N_2404,N_2369);
and U2984 (N_2984,N_2334,N_2068);
or U2985 (N_2985,N_2344,N_2166);
or U2986 (N_2986,N_2496,N_2139);
or U2987 (N_2987,N_2367,N_2047);
or U2988 (N_2988,N_2375,N_2195);
nand U2989 (N_2989,N_2452,N_2056);
nand U2990 (N_2990,N_2096,N_2302);
xor U2991 (N_2991,N_2019,N_2016);
nor U2992 (N_2992,N_2069,N_2118);
nand U2993 (N_2993,N_2428,N_2003);
xor U2994 (N_2994,N_2224,N_2073);
and U2995 (N_2995,N_2316,N_2052);
or U2996 (N_2996,N_2003,N_2252);
nand U2997 (N_2997,N_2278,N_2445);
and U2998 (N_2998,N_2016,N_2132);
nor U2999 (N_2999,N_2458,N_2405);
nor UO_0 (O_0,N_2900,N_2714);
and UO_1 (O_1,N_2561,N_2565);
and UO_2 (O_2,N_2623,N_2612);
and UO_3 (O_3,N_2556,N_2605);
xor UO_4 (O_4,N_2684,N_2628);
xnor UO_5 (O_5,N_2555,N_2888);
or UO_6 (O_6,N_2810,N_2506);
or UO_7 (O_7,N_2809,N_2698);
and UO_8 (O_8,N_2727,N_2598);
nor UO_9 (O_9,N_2877,N_2513);
nand UO_10 (O_10,N_2510,N_2652);
nand UO_11 (O_11,N_2795,N_2544);
and UO_12 (O_12,N_2878,N_2545);
nand UO_13 (O_13,N_2537,N_2525);
or UO_14 (O_14,N_2854,N_2531);
nand UO_15 (O_15,N_2630,N_2646);
and UO_16 (O_16,N_2892,N_2847);
nand UO_17 (O_17,N_2955,N_2585);
and UO_18 (O_18,N_2702,N_2905);
nand UO_19 (O_19,N_2532,N_2800);
nor UO_20 (O_20,N_2777,N_2781);
and UO_21 (O_21,N_2797,N_2944);
or UO_22 (O_22,N_2830,N_2601);
nand UO_23 (O_23,N_2660,N_2917);
nand UO_24 (O_24,N_2954,N_2577);
nor UO_25 (O_25,N_2583,N_2901);
or UO_26 (O_26,N_2975,N_2844);
or UO_27 (O_27,N_2642,N_2602);
and UO_28 (O_28,N_2857,N_2938);
nor UO_29 (O_29,N_2618,N_2841);
nor UO_30 (O_30,N_2693,N_2734);
nor UO_31 (O_31,N_2580,N_2672);
nand UO_32 (O_32,N_2657,N_2837);
or UO_33 (O_33,N_2502,N_2568);
nand UO_34 (O_34,N_2690,N_2984);
nor UO_35 (O_35,N_2989,N_2681);
nand UO_36 (O_36,N_2564,N_2974);
and UO_37 (O_37,N_2579,N_2875);
and UO_38 (O_38,N_2910,N_2551);
and UO_39 (O_39,N_2633,N_2922);
nand UO_40 (O_40,N_2807,N_2895);
nand UO_41 (O_41,N_2696,N_2839);
or UO_42 (O_42,N_2593,N_2645);
or UO_43 (O_43,N_2870,N_2739);
and UO_44 (O_44,N_2833,N_2767);
nor UO_45 (O_45,N_2629,N_2803);
and UO_46 (O_46,N_2559,N_2615);
or UO_47 (O_47,N_2759,N_2838);
and UO_48 (O_48,N_2906,N_2625);
or UO_49 (O_49,N_2653,N_2829);
and UO_50 (O_50,N_2526,N_2997);
or UO_51 (O_51,N_2884,N_2707);
or UO_52 (O_52,N_2921,N_2783);
and UO_53 (O_53,N_2762,N_2654);
nor UO_54 (O_54,N_2998,N_2950);
or UO_55 (O_55,N_2740,N_2587);
nand UO_56 (O_56,N_2514,N_2907);
or UO_57 (O_57,N_2924,N_2624);
nand UO_58 (O_58,N_2933,N_2791);
nand UO_59 (O_59,N_2988,N_2869);
nand UO_60 (O_60,N_2687,N_2616);
or UO_61 (O_61,N_2661,N_2966);
nor UO_62 (O_62,N_2603,N_2852);
nor UO_63 (O_63,N_2765,N_2971);
and UO_64 (O_64,N_2972,N_2996);
and UO_65 (O_65,N_2617,N_2717);
or UO_66 (O_66,N_2929,N_2804);
or UO_67 (O_67,N_2599,N_2927);
and UO_68 (O_68,N_2918,N_2539);
nand UO_69 (O_69,N_2963,N_2814);
nor UO_70 (O_70,N_2578,N_2648);
xnor UO_71 (O_71,N_2744,N_2610);
xor UO_72 (O_72,N_2597,N_2865);
nand UO_73 (O_73,N_2862,N_2903);
nor UO_74 (O_74,N_2755,N_2764);
and UO_75 (O_75,N_2771,N_2571);
or UO_76 (O_76,N_2641,N_2656);
and UO_77 (O_77,N_2926,N_2674);
nand UO_78 (O_78,N_2512,N_2941);
and UO_79 (O_79,N_2812,N_2775);
and UO_80 (O_80,N_2978,N_2980);
nand UO_81 (O_81,N_2589,N_2779);
nand UO_82 (O_82,N_2991,N_2529);
nand UO_83 (O_83,N_2705,N_2915);
or UO_84 (O_84,N_2826,N_2746);
and UO_85 (O_85,N_2890,N_2643);
and UO_86 (O_86,N_2688,N_2521);
and UO_87 (O_87,N_2703,N_2673);
nand UO_88 (O_88,N_2823,N_2967);
or UO_89 (O_89,N_2650,N_2945);
or UO_90 (O_90,N_2520,N_2621);
or UO_91 (O_91,N_2749,N_2784);
or UO_92 (O_92,N_2956,N_2840);
nor UO_93 (O_93,N_2543,N_2936);
and UO_94 (O_94,N_2715,N_2663);
nor UO_95 (O_95,N_2942,N_2581);
nor UO_96 (O_96,N_2756,N_2776);
nor UO_97 (O_97,N_2914,N_2994);
and UO_98 (O_98,N_2596,N_2773);
or UO_99 (O_99,N_2524,N_2738);
nand UO_100 (O_100,N_2821,N_2939);
nor UO_101 (O_101,N_2752,N_2832);
nor UO_102 (O_102,N_2874,N_2557);
and UO_103 (O_103,N_2894,N_2518);
or UO_104 (O_104,N_2952,N_2848);
nand UO_105 (O_105,N_2897,N_2572);
or UO_106 (O_106,N_2889,N_2552);
nor UO_107 (O_107,N_2965,N_2588);
nand UO_108 (O_108,N_2763,N_2730);
nor UO_109 (O_109,N_2569,N_2753);
and UO_110 (O_110,N_2778,N_2716);
and UO_111 (O_111,N_2573,N_2508);
xor UO_112 (O_112,N_2668,N_2882);
nand UO_113 (O_113,N_2570,N_2636);
or UO_114 (O_114,N_2947,N_2757);
and UO_115 (O_115,N_2644,N_2970);
nor UO_116 (O_116,N_2879,N_2611);
or UO_117 (O_117,N_2788,N_2806);
and UO_118 (O_118,N_2600,N_2866);
or UO_119 (O_119,N_2567,N_2834);
nor UO_120 (O_120,N_2920,N_2949);
or UO_121 (O_121,N_2535,N_2962);
and UO_122 (O_122,N_2522,N_2799);
nand UO_123 (O_123,N_2808,N_2576);
nor UO_124 (O_124,N_2842,N_2566);
nand UO_125 (O_125,N_2675,N_2986);
nand UO_126 (O_126,N_2981,N_2768);
nand UO_127 (O_127,N_2733,N_2639);
nor UO_128 (O_128,N_2726,N_2904);
or UO_129 (O_129,N_2563,N_2881);
and UO_130 (O_130,N_2880,N_2898);
nand UO_131 (O_131,N_2912,N_2849);
or UO_132 (O_132,N_2590,N_2632);
nor UO_133 (O_133,N_2902,N_2586);
or UO_134 (O_134,N_2943,N_2729);
nand UO_135 (O_135,N_2640,N_2990);
or UO_136 (O_136,N_2747,N_2613);
nor UO_137 (O_137,N_2536,N_2719);
nor UO_138 (O_138,N_2604,N_2527);
and UO_139 (O_139,N_2699,N_2546);
nand UO_140 (O_140,N_2709,N_2973);
nor UO_141 (O_141,N_2509,N_2504);
nor UO_142 (O_142,N_2824,N_2876);
or UO_143 (O_143,N_2780,N_2669);
nor UO_144 (O_144,N_2995,N_2958);
nor UO_145 (O_145,N_2712,N_2846);
nor UO_146 (O_146,N_2953,N_2792);
nor UO_147 (O_147,N_2761,N_2893);
nor UO_148 (O_148,N_2793,N_2999);
nand UO_149 (O_149,N_2886,N_2503);
or UO_150 (O_150,N_2622,N_2883);
nand UO_151 (O_151,N_2718,N_2885);
nand UO_152 (O_152,N_2620,N_2549);
or UO_153 (O_153,N_2523,N_2679);
nor UO_154 (O_154,N_2860,N_2969);
nand UO_155 (O_155,N_2676,N_2934);
and UO_156 (O_156,N_2811,N_2711);
nor UO_157 (O_157,N_2731,N_2871);
or UO_158 (O_158,N_2548,N_2750);
or UO_159 (O_159,N_2519,N_2850);
and UO_160 (O_160,N_2946,N_2592);
or UO_161 (O_161,N_2798,N_2964);
nor UO_162 (O_162,N_2951,N_2932);
or UO_163 (O_163,N_2528,N_2720);
or UO_164 (O_164,N_2968,N_2634);
nor UO_165 (O_165,N_2626,N_2627);
and UO_166 (O_166,N_2856,N_2710);
nand UO_167 (O_167,N_2851,N_2819);
nor UO_168 (O_168,N_2701,N_2913);
nand UO_169 (O_169,N_2706,N_2655);
or UO_170 (O_170,N_2813,N_2948);
nor UO_171 (O_171,N_2659,N_2722);
xor UO_172 (O_172,N_2993,N_2591);
nand UO_173 (O_173,N_2560,N_2649);
and UO_174 (O_174,N_2836,N_2916);
and UO_175 (O_175,N_2959,N_2501);
nor UO_176 (O_176,N_2670,N_2515);
nand UO_177 (O_177,N_2831,N_2985);
nor UO_178 (O_178,N_2500,N_2682);
nor UO_179 (O_179,N_2743,N_2737);
and UO_180 (O_180,N_2664,N_2540);
and UO_181 (O_181,N_2665,N_2516);
nor UO_182 (O_182,N_2911,N_2606);
and UO_183 (O_183,N_2671,N_2787);
nand UO_184 (O_184,N_2541,N_2935);
nor UO_185 (O_185,N_2631,N_2694);
or UO_186 (O_186,N_2957,N_2827);
nand UO_187 (O_187,N_2662,N_2635);
nand UO_188 (O_188,N_2925,N_2802);
or UO_189 (O_189,N_2721,N_2796);
and UO_190 (O_190,N_2562,N_2908);
and UO_191 (O_191,N_2864,N_2651);
and UO_192 (O_192,N_2695,N_2517);
and UO_193 (O_193,N_2760,N_2547);
nand UO_194 (O_194,N_2822,N_2863);
nor UO_195 (O_195,N_2751,N_2774);
and UO_196 (O_196,N_2724,N_2584);
and UO_197 (O_197,N_2977,N_2937);
nor UO_198 (O_198,N_2553,N_2741);
nand UO_199 (O_199,N_2960,N_2982);
and UO_200 (O_200,N_2683,N_2692);
and UO_201 (O_201,N_2538,N_2614);
nor UO_202 (O_202,N_2554,N_2872);
and UO_203 (O_203,N_2825,N_2896);
or UO_204 (O_204,N_2708,N_2845);
or UO_205 (O_205,N_2891,N_2859);
nor UO_206 (O_206,N_2766,N_2818);
nand UO_207 (O_207,N_2505,N_2919);
nor UO_208 (O_208,N_2930,N_2992);
nand UO_209 (O_209,N_2507,N_2732);
xor UO_210 (O_210,N_2782,N_2940);
or UO_211 (O_211,N_2976,N_2533);
nor UO_212 (O_212,N_2909,N_2686);
nor UO_213 (O_213,N_2697,N_2638);
and UO_214 (O_214,N_2758,N_2542);
nor UO_215 (O_215,N_2658,N_2887);
nor UO_216 (O_216,N_2828,N_2595);
or UO_217 (O_217,N_2608,N_2790);
and UO_218 (O_218,N_2855,N_2785);
nor UO_219 (O_219,N_2723,N_2979);
or UO_220 (O_220,N_2728,N_2769);
or UO_221 (O_221,N_2691,N_2574);
nor UO_222 (O_222,N_2637,N_2923);
nand UO_223 (O_223,N_2736,N_2689);
or UO_224 (O_224,N_2786,N_2867);
and UO_225 (O_225,N_2899,N_2680);
nand UO_226 (O_226,N_2594,N_2609);
nor UO_227 (O_227,N_2511,N_2861);
or UO_228 (O_228,N_2745,N_2835);
and UO_229 (O_229,N_2754,N_2748);
and UO_230 (O_230,N_2704,N_2607);
xnor UO_231 (O_231,N_2713,N_2805);
and UO_232 (O_232,N_2873,N_2853);
nand UO_233 (O_233,N_2817,N_2685);
nor UO_234 (O_234,N_2735,N_2868);
or UO_235 (O_235,N_2987,N_2858);
and UO_236 (O_236,N_2666,N_2647);
nor UO_237 (O_237,N_2550,N_2725);
or UO_238 (O_238,N_2772,N_2677);
nand UO_239 (O_239,N_2534,N_2678);
nand UO_240 (O_240,N_2530,N_2843);
nand UO_241 (O_241,N_2770,N_2815);
nand UO_242 (O_242,N_2801,N_2667);
or UO_243 (O_243,N_2558,N_2582);
and UO_244 (O_244,N_2742,N_2794);
nand UO_245 (O_245,N_2931,N_2789);
xor UO_246 (O_246,N_2961,N_2816);
and UO_247 (O_247,N_2619,N_2575);
nand UO_248 (O_248,N_2820,N_2983);
or UO_249 (O_249,N_2700,N_2928);
and UO_250 (O_250,N_2701,N_2917);
nor UO_251 (O_251,N_2877,N_2669);
nand UO_252 (O_252,N_2869,N_2634);
or UO_253 (O_253,N_2696,N_2644);
nor UO_254 (O_254,N_2650,N_2958);
nor UO_255 (O_255,N_2851,N_2739);
nand UO_256 (O_256,N_2641,N_2850);
nand UO_257 (O_257,N_2514,N_2960);
nor UO_258 (O_258,N_2683,N_2992);
nor UO_259 (O_259,N_2821,N_2500);
or UO_260 (O_260,N_2548,N_2720);
and UO_261 (O_261,N_2693,N_2982);
and UO_262 (O_262,N_2558,N_2914);
or UO_263 (O_263,N_2644,N_2791);
nand UO_264 (O_264,N_2902,N_2692);
xor UO_265 (O_265,N_2617,N_2692);
and UO_266 (O_266,N_2720,N_2553);
nor UO_267 (O_267,N_2626,N_2529);
and UO_268 (O_268,N_2667,N_2671);
nor UO_269 (O_269,N_2526,N_2844);
and UO_270 (O_270,N_2841,N_2770);
or UO_271 (O_271,N_2956,N_2837);
and UO_272 (O_272,N_2526,N_2655);
and UO_273 (O_273,N_2708,N_2863);
and UO_274 (O_274,N_2577,N_2574);
or UO_275 (O_275,N_2565,N_2548);
and UO_276 (O_276,N_2738,N_2601);
nor UO_277 (O_277,N_2511,N_2546);
and UO_278 (O_278,N_2747,N_2921);
nand UO_279 (O_279,N_2830,N_2751);
or UO_280 (O_280,N_2871,N_2826);
nand UO_281 (O_281,N_2694,N_2848);
and UO_282 (O_282,N_2846,N_2715);
nor UO_283 (O_283,N_2628,N_2589);
or UO_284 (O_284,N_2782,N_2907);
and UO_285 (O_285,N_2540,N_2945);
nand UO_286 (O_286,N_2868,N_2980);
and UO_287 (O_287,N_2941,N_2858);
nor UO_288 (O_288,N_2624,N_2704);
xnor UO_289 (O_289,N_2565,N_2633);
nand UO_290 (O_290,N_2993,N_2979);
or UO_291 (O_291,N_2503,N_2858);
and UO_292 (O_292,N_2609,N_2943);
or UO_293 (O_293,N_2506,N_2531);
and UO_294 (O_294,N_2743,N_2886);
nand UO_295 (O_295,N_2847,N_2758);
or UO_296 (O_296,N_2713,N_2902);
nor UO_297 (O_297,N_2512,N_2623);
nor UO_298 (O_298,N_2689,N_2651);
or UO_299 (O_299,N_2667,N_2630);
nor UO_300 (O_300,N_2904,N_2933);
or UO_301 (O_301,N_2907,N_2503);
or UO_302 (O_302,N_2833,N_2976);
and UO_303 (O_303,N_2922,N_2965);
nor UO_304 (O_304,N_2698,N_2730);
and UO_305 (O_305,N_2701,N_2763);
and UO_306 (O_306,N_2727,N_2589);
nand UO_307 (O_307,N_2572,N_2981);
nor UO_308 (O_308,N_2606,N_2505);
xnor UO_309 (O_309,N_2786,N_2502);
nand UO_310 (O_310,N_2712,N_2974);
nand UO_311 (O_311,N_2588,N_2540);
or UO_312 (O_312,N_2644,N_2624);
nor UO_313 (O_313,N_2961,N_2951);
nand UO_314 (O_314,N_2552,N_2512);
nor UO_315 (O_315,N_2503,N_2586);
nand UO_316 (O_316,N_2976,N_2879);
or UO_317 (O_317,N_2832,N_2726);
nand UO_318 (O_318,N_2987,N_2702);
or UO_319 (O_319,N_2868,N_2988);
nand UO_320 (O_320,N_2771,N_2933);
and UO_321 (O_321,N_2618,N_2808);
nand UO_322 (O_322,N_2739,N_2727);
nand UO_323 (O_323,N_2512,N_2895);
and UO_324 (O_324,N_2605,N_2917);
and UO_325 (O_325,N_2667,N_2780);
xnor UO_326 (O_326,N_2657,N_2711);
or UO_327 (O_327,N_2890,N_2988);
and UO_328 (O_328,N_2906,N_2762);
or UO_329 (O_329,N_2711,N_2610);
and UO_330 (O_330,N_2524,N_2583);
nor UO_331 (O_331,N_2670,N_2917);
nor UO_332 (O_332,N_2743,N_2891);
nor UO_333 (O_333,N_2952,N_2781);
and UO_334 (O_334,N_2649,N_2593);
nand UO_335 (O_335,N_2593,N_2944);
nand UO_336 (O_336,N_2620,N_2650);
nor UO_337 (O_337,N_2761,N_2592);
and UO_338 (O_338,N_2652,N_2591);
nand UO_339 (O_339,N_2698,N_2891);
or UO_340 (O_340,N_2624,N_2712);
nand UO_341 (O_341,N_2871,N_2869);
nor UO_342 (O_342,N_2619,N_2525);
xor UO_343 (O_343,N_2940,N_2502);
and UO_344 (O_344,N_2730,N_2555);
and UO_345 (O_345,N_2537,N_2755);
or UO_346 (O_346,N_2966,N_2858);
or UO_347 (O_347,N_2686,N_2868);
or UO_348 (O_348,N_2686,N_2689);
or UO_349 (O_349,N_2976,N_2501);
or UO_350 (O_350,N_2872,N_2637);
and UO_351 (O_351,N_2638,N_2968);
or UO_352 (O_352,N_2564,N_2815);
and UO_353 (O_353,N_2951,N_2999);
nor UO_354 (O_354,N_2859,N_2524);
nor UO_355 (O_355,N_2679,N_2650);
nor UO_356 (O_356,N_2665,N_2889);
nand UO_357 (O_357,N_2791,N_2885);
nand UO_358 (O_358,N_2594,N_2902);
xor UO_359 (O_359,N_2811,N_2830);
or UO_360 (O_360,N_2540,N_2981);
nor UO_361 (O_361,N_2986,N_2814);
and UO_362 (O_362,N_2831,N_2703);
xor UO_363 (O_363,N_2511,N_2971);
and UO_364 (O_364,N_2672,N_2794);
and UO_365 (O_365,N_2633,N_2748);
nor UO_366 (O_366,N_2716,N_2511);
and UO_367 (O_367,N_2707,N_2796);
or UO_368 (O_368,N_2564,N_2812);
nand UO_369 (O_369,N_2627,N_2706);
or UO_370 (O_370,N_2966,N_2845);
nor UO_371 (O_371,N_2783,N_2835);
nand UO_372 (O_372,N_2907,N_2681);
or UO_373 (O_373,N_2879,N_2653);
nor UO_374 (O_374,N_2877,N_2578);
and UO_375 (O_375,N_2780,N_2860);
nand UO_376 (O_376,N_2924,N_2599);
nand UO_377 (O_377,N_2746,N_2795);
nand UO_378 (O_378,N_2958,N_2814);
or UO_379 (O_379,N_2691,N_2865);
and UO_380 (O_380,N_2712,N_2937);
nor UO_381 (O_381,N_2635,N_2655);
nor UO_382 (O_382,N_2866,N_2554);
or UO_383 (O_383,N_2733,N_2561);
nand UO_384 (O_384,N_2979,N_2827);
or UO_385 (O_385,N_2676,N_2848);
nand UO_386 (O_386,N_2698,N_2830);
or UO_387 (O_387,N_2669,N_2864);
or UO_388 (O_388,N_2891,N_2932);
nor UO_389 (O_389,N_2702,N_2811);
and UO_390 (O_390,N_2765,N_2681);
nor UO_391 (O_391,N_2735,N_2794);
or UO_392 (O_392,N_2795,N_2988);
or UO_393 (O_393,N_2920,N_2567);
or UO_394 (O_394,N_2632,N_2763);
and UO_395 (O_395,N_2812,N_2856);
nor UO_396 (O_396,N_2705,N_2988);
nand UO_397 (O_397,N_2623,N_2617);
nand UO_398 (O_398,N_2541,N_2661);
and UO_399 (O_399,N_2872,N_2535);
nor UO_400 (O_400,N_2668,N_2899);
nor UO_401 (O_401,N_2579,N_2720);
nand UO_402 (O_402,N_2709,N_2688);
nand UO_403 (O_403,N_2996,N_2740);
or UO_404 (O_404,N_2984,N_2726);
nand UO_405 (O_405,N_2853,N_2675);
nand UO_406 (O_406,N_2989,N_2866);
or UO_407 (O_407,N_2642,N_2715);
nor UO_408 (O_408,N_2717,N_2978);
nand UO_409 (O_409,N_2604,N_2885);
nand UO_410 (O_410,N_2760,N_2708);
nor UO_411 (O_411,N_2684,N_2565);
or UO_412 (O_412,N_2972,N_2533);
and UO_413 (O_413,N_2775,N_2997);
nor UO_414 (O_414,N_2854,N_2656);
or UO_415 (O_415,N_2673,N_2847);
nand UO_416 (O_416,N_2698,N_2653);
nor UO_417 (O_417,N_2541,N_2543);
and UO_418 (O_418,N_2943,N_2739);
and UO_419 (O_419,N_2615,N_2545);
nor UO_420 (O_420,N_2971,N_2622);
or UO_421 (O_421,N_2955,N_2749);
nor UO_422 (O_422,N_2688,N_2869);
or UO_423 (O_423,N_2875,N_2848);
and UO_424 (O_424,N_2682,N_2659);
nor UO_425 (O_425,N_2797,N_2872);
and UO_426 (O_426,N_2987,N_2697);
nand UO_427 (O_427,N_2765,N_2957);
or UO_428 (O_428,N_2602,N_2758);
nor UO_429 (O_429,N_2613,N_2516);
and UO_430 (O_430,N_2666,N_2546);
nor UO_431 (O_431,N_2539,N_2839);
or UO_432 (O_432,N_2740,N_2783);
or UO_433 (O_433,N_2719,N_2926);
nor UO_434 (O_434,N_2956,N_2724);
nor UO_435 (O_435,N_2550,N_2731);
nand UO_436 (O_436,N_2620,N_2622);
xnor UO_437 (O_437,N_2537,N_2594);
or UO_438 (O_438,N_2532,N_2827);
nor UO_439 (O_439,N_2551,N_2594);
nand UO_440 (O_440,N_2513,N_2563);
or UO_441 (O_441,N_2667,N_2879);
or UO_442 (O_442,N_2502,N_2839);
nor UO_443 (O_443,N_2652,N_2628);
and UO_444 (O_444,N_2851,N_2594);
or UO_445 (O_445,N_2639,N_2974);
and UO_446 (O_446,N_2580,N_2934);
nor UO_447 (O_447,N_2609,N_2763);
and UO_448 (O_448,N_2753,N_2588);
and UO_449 (O_449,N_2966,N_2877);
and UO_450 (O_450,N_2820,N_2515);
xnor UO_451 (O_451,N_2560,N_2672);
nand UO_452 (O_452,N_2796,N_2677);
nand UO_453 (O_453,N_2551,N_2607);
and UO_454 (O_454,N_2981,N_2961);
nand UO_455 (O_455,N_2589,N_2817);
nand UO_456 (O_456,N_2795,N_2817);
nor UO_457 (O_457,N_2673,N_2979);
xor UO_458 (O_458,N_2521,N_2665);
and UO_459 (O_459,N_2755,N_2767);
xnor UO_460 (O_460,N_2743,N_2828);
and UO_461 (O_461,N_2820,N_2864);
or UO_462 (O_462,N_2645,N_2580);
and UO_463 (O_463,N_2858,N_2995);
or UO_464 (O_464,N_2674,N_2795);
nand UO_465 (O_465,N_2840,N_2920);
or UO_466 (O_466,N_2753,N_2700);
or UO_467 (O_467,N_2961,N_2892);
and UO_468 (O_468,N_2729,N_2715);
or UO_469 (O_469,N_2912,N_2525);
and UO_470 (O_470,N_2702,N_2998);
and UO_471 (O_471,N_2907,N_2904);
or UO_472 (O_472,N_2783,N_2544);
and UO_473 (O_473,N_2992,N_2853);
nand UO_474 (O_474,N_2832,N_2600);
and UO_475 (O_475,N_2855,N_2694);
nand UO_476 (O_476,N_2810,N_2707);
nor UO_477 (O_477,N_2708,N_2513);
nor UO_478 (O_478,N_2597,N_2728);
or UO_479 (O_479,N_2820,N_2613);
or UO_480 (O_480,N_2738,N_2672);
or UO_481 (O_481,N_2677,N_2709);
or UO_482 (O_482,N_2916,N_2544);
nand UO_483 (O_483,N_2507,N_2825);
or UO_484 (O_484,N_2978,N_2798);
and UO_485 (O_485,N_2721,N_2781);
or UO_486 (O_486,N_2970,N_2856);
nor UO_487 (O_487,N_2617,N_2968);
or UO_488 (O_488,N_2850,N_2966);
or UO_489 (O_489,N_2967,N_2791);
and UO_490 (O_490,N_2837,N_2966);
nor UO_491 (O_491,N_2971,N_2628);
and UO_492 (O_492,N_2537,N_2893);
nand UO_493 (O_493,N_2748,N_2556);
or UO_494 (O_494,N_2793,N_2786);
nor UO_495 (O_495,N_2660,N_2839);
nand UO_496 (O_496,N_2969,N_2831);
nor UO_497 (O_497,N_2921,N_2681);
and UO_498 (O_498,N_2506,N_2990);
nor UO_499 (O_499,N_2962,N_2675);
endmodule