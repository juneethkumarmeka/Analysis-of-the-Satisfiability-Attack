module basic_500_3000_500_6_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_262,In_241);
nand U1 (N_1,In_282,In_470);
and U2 (N_2,In_63,In_450);
or U3 (N_3,In_461,In_74);
or U4 (N_4,In_269,In_96);
and U5 (N_5,In_34,In_300);
nand U6 (N_6,In_477,In_42);
or U7 (N_7,In_29,In_65);
nand U8 (N_8,In_260,In_204);
nand U9 (N_9,In_255,In_71);
nor U10 (N_10,In_18,In_379);
nor U11 (N_11,In_38,In_484);
nor U12 (N_12,In_105,In_87);
or U13 (N_13,In_208,In_181);
or U14 (N_14,In_438,In_133);
and U15 (N_15,In_197,In_32);
nor U16 (N_16,In_7,In_367);
xor U17 (N_17,In_271,In_344);
nor U18 (N_18,In_298,In_354);
nand U19 (N_19,In_26,In_369);
xor U20 (N_20,In_377,In_424);
nand U21 (N_21,In_160,In_136);
xnor U22 (N_22,In_313,In_53);
nand U23 (N_23,In_246,In_419);
and U24 (N_24,In_153,In_61);
nor U25 (N_25,In_414,In_340);
or U26 (N_26,In_99,In_259);
or U27 (N_27,In_326,In_10);
or U28 (N_28,In_283,In_47);
nand U29 (N_29,In_104,In_244);
or U30 (N_30,In_270,In_49);
and U31 (N_31,In_485,In_207);
xor U32 (N_32,In_209,In_199);
and U33 (N_33,In_368,In_51);
nand U34 (N_34,In_84,In_107);
nor U35 (N_35,In_472,In_458);
and U36 (N_36,In_124,In_41);
nand U37 (N_37,In_120,In_219);
or U38 (N_38,In_94,In_141);
and U39 (N_39,In_119,In_329);
or U40 (N_40,In_79,In_406);
or U41 (N_41,In_169,In_400);
and U42 (N_42,In_361,In_195);
nand U43 (N_43,In_426,In_146);
xor U44 (N_44,In_425,In_218);
and U45 (N_45,In_495,In_234);
nor U46 (N_46,In_48,In_278);
nor U47 (N_47,In_455,In_43);
nand U48 (N_48,In_410,In_158);
nand U49 (N_49,In_135,In_205);
and U50 (N_50,In_242,In_436);
nand U51 (N_51,In_92,In_266);
or U52 (N_52,In_265,In_371);
or U53 (N_53,In_452,In_147);
or U54 (N_54,In_186,In_295);
or U55 (N_55,In_106,In_356);
nor U56 (N_56,In_75,In_491);
nand U57 (N_57,In_392,In_6);
and U58 (N_58,In_114,In_433);
nor U59 (N_59,In_319,In_474);
nand U60 (N_60,In_466,In_468);
or U61 (N_61,In_301,In_479);
nor U62 (N_62,In_162,In_129);
and U63 (N_63,In_232,In_274);
xnor U64 (N_64,In_441,In_78);
nand U65 (N_65,In_353,In_446);
or U66 (N_66,In_76,In_396);
xor U67 (N_67,In_183,In_413);
nor U68 (N_68,In_365,In_200);
nor U69 (N_69,In_364,In_148);
or U70 (N_70,In_467,In_276);
xor U71 (N_71,In_193,In_291);
and U72 (N_72,In_486,In_56);
and U73 (N_73,In_203,In_151);
nand U74 (N_74,In_268,In_417);
or U75 (N_75,In_206,In_130);
or U76 (N_76,In_173,In_494);
or U77 (N_77,In_152,In_316);
xor U78 (N_78,In_496,In_334);
and U79 (N_79,In_166,In_388);
or U80 (N_80,In_385,In_220);
and U81 (N_81,In_349,In_13);
nor U82 (N_82,In_412,In_40);
or U83 (N_83,In_460,In_297);
xnor U84 (N_84,In_277,In_342);
nor U85 (N_85,In_302,In_256);
and U86 (N_86,In_73,In_284);
or U87 (N_87,In_225,In_435);
xnor U88 (N_88,In_437,In_311);
and U89 (N_89,In_192,In_488);
and U90 (N_90,In_101,In_222);
nand U91 (N_91,In_428,In_381);
xor U92 (N_92,In_176,In_336);
xor U93 (N_93,In_123,In_386);
xor U94 (N_94,In_1,In_25);
or U95 (N_95,In_387,In_66);
nand U96 (N_96,In_185,In_170);
nor U97 (N_97,In_231,In_355);
and U98 (N_98,In_235,In_167);
or U99 (N_99,In_240,In_211);
and U100 (N_100,In_161,In_493);
and U101 (N_101,In_214,In_462);
and U102 (N_102,In_407,In_352);
nor U103 (N_103,In_475,In_389);
or U104 (N_104,In_445,In_402);
and U105 (N_105,In_469,In_331);
nor U106 (N_106,In_212,In_20);
and U107 (N_107,In_159,In_325);
nor U108 (N_108,In_37,In_126);
nand U109 (N_109,In_382,In_131);
nand U110 (N_110,In_247,In_90);
nor U111 (N_111,In_337,In_22);
nor U112 (N_112,In_254,In_431);
nor U113 (N_113,In_62,In_314);
xnor U114 (N_114,In_332,In_14);
and U115 (N_115,In_363,In_45);
and U116 (N_116,In_459,In_21);
and U117 (N_117,In_60,In_83);
nand U118 (N_118,In_238,In_2);
and U119 (N_119,In_86,In_157);
nor U120 (N_120,In_272,In_116);
and U121 (N_121,In_453,In_328);
and U122 (N_122,In_113,In_24);
nand U123 (N_123,In_150,In_97);
and U124 (N_124,In_343,In_154);
nor U125 (N_125,In_429,In_285);
or U126 (N_126,In_70,In_286);
nand U127 (N_127,In_121,In_196);
or U128 (N_128,In_401,In_165);
or U129 (N_129,In_499,In_399);
nor U130 (N_130,In_308,In_346);
and U131 (N_131,In_391,In_492);
nor U132 (N_132,In_11,In_201);
and U133 (N_133,In_28,In_471);
or U134 (N_134,In_187,In_180);
and U135 (N_135,In_109,In_481);
xor U136 (N_136,In_476,In_44);
or U137 (N_137,In_293,In_434);
nor U138 (N_138,In_454,In_68);
and U139 (N_139,In_306,In_226);
nand U140 (N_140,In_320,In_67);
and U141 (N_141,In_134,In_447);
nand U142 (N_142,In_373,In_350);
or U143 (N_143,In_296,In_395);
nor U144 (N_144,In_415,In_178);
or U145 (N_145,In_432,In_357);
nor U146 (N_146,In_210,In_305);
nand U147 (N_147,In_184,In_375);
and U148 (N_148,In_215,In_341);
nand U149 (N_149,In_138,In_118);
or U150 (N_150,In_245,In_478);
xnor U151 (N_151,In_439,In_289);
or U152 (N_152,In_190,In_102);
nand U153 (N_153,In_122,In_405);
xor U154 (N_154,In_80,In_292);
xor U155 (N_155,In_403,In_318);
and U156 (N_156,In_27,In_82);
and U157 (N_157,In_50,In_339);
nand U158 (N_158,In_487,In_132);
nor U159 (N_159,In_422,In_125);
and U160 (N_160,In_451,In_448);
nand U161 (N_161,In_465,In_128);
or U162 (N_162,In_348,In_224);
or U163 (N_163,In_54,In_281);
nor U164 (N_164,In_294,In_213);
or U165 (N_165,In_366,In_117);
nand U166 (N_166,In_228,In_91);
nand U167 (N_167,In_110,In_248);
and U168 (N_168,In_252,In_52);
and U169 (N_169,In_16,In_243);
or U170 (N_170,In_93,In_15);
xor U171 (N_171,In_310,In_394);
or U172 (N_172,In_444,In_279);
and U173 (N_173,In_250,In_17);
and U174 (N_174,In_333,In_347);
nand U175 (N_175,In_194,In_89);
nor U176 (N_176,In_239,In_483);
xnor U177 (N_177,In_380,In_236);
nand U178 (N_178,In_497,In_108);
nor U179 (N_179,In_189,In_449);
and U180 (N_180,In_33,In_23);
nand U181 (N_181,In_140,In_249);
nor U182 (N_182,In_490,In_57);
nand U183 (N_183,In_217,In_95);
nand U184 (N_184,In_409,In_175);
and U185 (N_185,In_299,In_430);
or U186 (N_186,In_88,In_230);
nor U187 (N_187,In_288,In_427);
nand U188 (N_188,In_489,In_30);
or U189 (N_189,In_19,In_482);
xor U190 (N_190,In_223,In_345);
or U191 (N_191,In_251,In_317);
nor U192 (N_192,In_418,In_72);
and U193 (N_193,In_0,In_473);
xor U194 (N_194,In_8,In_290);
and U195 (N_195,In_35,In_36);
nor U196 (N_196,In_145,In_216);
and U197 (N_197,In_237,In_221);
and U198 (N_198,In_174,In_359);
xnor U199 (N_199,In_351,In_307);
or U200 (N_200,In_440,In_198);
or U201 (N_201,In_335,In_398);
nand U202 (N_202,In_4,In_182);
and U203 (N_203,In_423,In_55);
and U204 (N_204,In_64,In_315);
nand U205 (N_205,In_5,In_227);
or U206 (N_206,In_139,In_163);
or U207 (N_207,In_287,In_112);
or U208 (N_208,In_143,In_498);
or U209 (N_209,In_233,In_393);
and U210 (N_210,In_383,In_3);
nor U211 (N_211,In_358,In_172);
and U212 (N_212,In_321,In_312);
and U213 (N_213,In_384,In_327);
or U214 (N_214,In_155,In_144);
or U215 (N_215,In_263,In_179);
xnor U216 (N_216,In_273,In_324);
nor U217 (N_217,In_416,In_456);
or U218 (N_218,In_258,In_59);
nand U219 (N_219,In_442,In_275);
nand U220 (N_220,In_330,In_111);
nor U221 (N_221,In_370,In_463);
nand U222 (N_222,In_77,In_164);
nor U223 (N_223,In_421,In_127);
or U224 (N_224,In_257,In_304);
nor U225 (N_225,In_378,In_374);
and U226 (N_226,In_156,In_31);
or U227 (N_227,In_168,In_397);
nand U228 (N_228,In_360,In_85);
nand U229 (N_229,In_480,In_81);
nor U230 (N_230,In_253,In_69);
and U231 (N_231,In_390,In_303);
nor U232 (N_232,In_408,In_362);
xor U233 (N_233,In_100,In_12);
nor U234 (N_234,In_376,In_137);
and U235 (N_235,In_457,In_264);
nand U236 (N_236,In_229,In_372);
nand U237 (N_237,In_267,In_177);
nor U238 (N_238,In_149,In_188);
or U239 (N_239,In_323,In_420);
and U240 (N_240,In_58,In_46);
xnor U241 (N_241,In_171,In_338);
or U242 (N_242,In_98,In_39);
or U243 (N_243,In_115,In_309);
and U244 (N_244,In_404,In_411);
nor U245 (N_245,In_191,In_322);
nand U246 (N_246,In_9,In_464);
and U247 (N_247,In_202,In_280);
xor U248 (N_248,In_261,In_103);
nor U249 (N_249,In_142,In_443);
xnor U250 (N_250,In_429,In_492);
or U251 (N_251,In_461,In_18);
nor U252 (N_252,In_301,In_77);
or U253 (N_253,In_293,In_205);
or U254 (N_254,In_35,In_106);
and U255 (N_255,In_447,In_43);
and U256 (N_256,In_373,In_411);
nor U257 (N_257,In_47,In_415);
or U258 (N_258,In_494,In_279);
and U259 (N_259,In_218,In_234);
xnor U260 (N_260,In_474,In_202);
or U261 (N_261,In_489,In_308);
nand U262 (N_262,In_123,In_138);
and U263 (N_263,In_467,In_278);
or U264 (N_264,In_389,In_1);
and U265 (N_265,In_76,In_74);
nand U266 (N_266,In_448,In_440);
or U267 (N_267,In_425,In_198);
xor U268 (N_268,In_187,In_311);
nor U269 (N_269,In_247,In_26);
nor U270 (N_270,In_429,In_401);
xnor U271 (N_271,In_376,In_396);
nor U272 (N_272,In_149,In_139);
nor U273 (N_273,In_432,In_437);
xor U274 (N_274,In_280,In_248);
xor U275 (N_275,In_238,In_120);
nand U276 (N_276,In_56,In_215);
nand U277 (N_277,In_378,In_201);
nor U278 (N_278,In_449,In_131);
nand U279 (N_279,In_421,In_163);
and U280 (N_280,In_161,In_333);
or U281 (N_281,In_293,In_202);
nor U282 (N_282,In_333,In_75);
nand U283 (N_283,In_53,In_461);
or U284 (N_284,In_436,In_303);
nand U285 (N_285,In_65,In_237);
and U286 (N_286,In_275,In_39);
and U287 (N_287,In_244,In_9);
nor U288 (N_288,In_451,In_44);
nor U289 (N_289,In_131,In_463);
nand U290 (N_290,In_376,In_112);
or U291 (N_291,In_135,In_235);
or U292 (N_292,In_7,In_47);
nor U293 (N_293,In_458,In_166);
xor U294 (N_294,In_95,In_170);
or U295 (N_295,In_57,In_41);
or U296 (N_296,In_85,In_463);
nand U297 (N_297,In_435,In_197);
nor U298 (N_298,In_390,In_339);
or U299 (N_299,In_254,In_334);
xnor U300 (N_300,In_440,In_269);
and U301 (N_301,In_395,In_312);
and U302 (N_302,In_196,In_252);
nor U303 (N_303,In_238,In_84);
nand U304 (N_304,In_437,In_134);
nor U305 (N_305,In_262,In_428);
nand U306 (N_306,In_341,In_224);
nor U307 (N_307,In_95,In_45);
or U308 (N_308,In_181,In_354);
xor U309 (N_309,In_152,In_353);
and U310 (N_310,In_28,In_293);
or U311 (N_311,In_454,In_304);
nand U312 (N_312,In_272,In_456);
nand U313 (N_313,In_85,In_444);
nor U314 (N_314,In_475,In_488);
and U315 (N_315,In_106,In_46);
and U316 (N_316,In_443,In_45);
nor U317 (N_317,In_67,In_233);
nand U318 (N_318,In_104,In_364);
and U319 (N_319,In_482,In_33);
nand U320 (N_320,In_276,In_325);
nor U321 (N_321,In_26,In_43);
or U322 (N_322,In_187,In_156);
nand U323 (N_323,In_412,In_331);
nand U324 (N_324,In_414,In_107);
nor U325 (N_325,In_229,In_125);
nor U326 (N_326,In_391,In_488);
or U327 (N_327,In_30,In_179);
nand U328 (N_328,In_421,In_432);
or U329 (N_329,In_484,In_195);
or U330 (N_330,In_260,In_417);
nor U331 (N_331,In_195,In_67);
nand U332 (N_332,In_117,In_401);
and U333 (N_333,In_177,In_154);
nor U334 (N_334,In_391,In_54);
or U335 (N_335,In_153,In_384);
and U336 (N_336,In_437,In_281);
nor U337 (N_337,In_104,In_82);
nor U338 (N_338,In_293,In_3);
nand U339 (N_339,In_172,In_92);
or U340 (N_340,In_15,In_190);
xnor U341 (N_341,In_470,In_91);
nand U342 (N_342,In_100,In_474);
nand U343 (N_343,In_267,In_391);
and U344 (N_344,In_385,In_187);
or U345 (N_345,In_346,In_240);
nor U346 (N_346,In_495,In_57);
nor U347 (N_347,In_266,In_439);
nand U348 (N_348,In_260,In_439);
nand U349 (N_349,In_404,In_333);
and U350 (N_350,In_449,In_308);
and U351 (N_351,In_69,In_286);
and U352 (N_352,In_367,In_383);
or U353 (N_353,In_64,In_240);
xor U354 (N_354,In_184,In_151);
xnor U355 (N_355,In_209,In_109);
xnor U356 (N_356,In_165,In_152);
nor U357 (N_357,In_287,In_201);
or U358 (N_358,In_466,In_56);
and U359 (N_359,In_175,In_461);
nand U360 (N_360,In_260,In_326);
nand U361 (N_361,In_4,In_200);
nor U362 (N_362,In_317,In_241);
xnor U363 (N_363,In_87,In_396);
or U364 (N_364,In_65,In_57);
xor U365 (N_365,In_471,In_166);
nor U366 (N_366,In_39,In_78);
nand U367 (N_367,In_414,In_468);
or U368 (N_368,In_154,In_17);
and U369 (N_369,In_465,In_491);
and U370 (N_370,In_489,In_249);
or U371 (N_371,In_441,In_237);
xnor U372 (N_372,In_200,In_136);
and U373 (N_373,In_397,In_91);
or U374 (N_374,In_405,In_268);
nor U375 (N_375,In_411,In_16);
or U376 (N_376,In_499,In_79);
xnor U377 (N_377,In_359,In_406);
nand U378 (N_378,In_25,In_394);
nand U379 (N_379,In_242,In_464);
and U380 (N_380,In_93,In_493);
xor U381 (N_381,In_57,In_475);
nor U382 (N_382,In_150,In_192);
and U383 (N_383,In_189,In_245);
or U384 (N_384,In_353,In_240);
nand U385 (N_385,In_329,In_331);
nand U386 (N_386,In_413,In_198);
and U387 (N_387,In_310,In_171);
nor U388 (N_388,In_436,In_441);
nor U389 (N_389,In_197,In_479);
nand U390 (N_390,In_71,In_365);
xnor U391 (N_391,In_206,In_265);
nand U392 (N_392,In_438,In_366);
nand U393 (N_393,In_61,In_90);
nor U394 (N_394,In_479,In_407);
and U395 (N_395,In_295,In_279);
or U396 (N_396,In_103,In_148);
nand U397 (N_397,In_56,In_192);
nand U398 (N_398,In_20,In_358);
nand U399 (N_399,In_108,In_444);
nand U400 (N_400,In_381,In_267);
nor U401 (N_401,In_151,In_362);
and U402 (N_402,In_324,In_270);
nand U403 (N_403,In_459,In_498);
nand U404 (N_404,In_109,In_164);
and U405 (N_405,In_209,In_91);
nor U406 (N_406,In_301,In_133);
or U407 (N_407,In_315,In_387);
or U408 (N_408,In_264,In_399);
xor U409 (N_409,In_499,In_117);
nor U410 (N_410,In_373,In_286);
and U411 (N_411,In_394,In_126);
and U412 (N_412,In_331,In_428);
and U413 (N_413,In_157,In_321);
xnor U414 (N_414,In_374,In_22);
nand U415 (N_415,In_114,In_214);
nor U416 (N_416,In_344,In_57);
nand U417 (N_417,In_490,In_360);
or U418 (N_418,In_107,In_132);
nor U419 (N_419,In_483,In_472);
or U420 (N_420,In_391,In_245);
and U421 (N_421,In_164,In_372);
and U422 (N_422,In_425,In_135);
nor U423 (N_423,In_369,In_319);
and U424 (N_424,In_50,In_126);
and U425 (N_425,In_274,In_96);
nand U426 (N_426,In_39,In_436);
and U427 (N_427,In_484,In_452);
and U428 (N_428,In_332,In_128);
or U429 (N_429,In_463,In_270);
xnor U430 (N_430,In_153,In_333);
nand U431 (N_431,In_126,In_259);
nor U432 (N_432,In_293,In_31);
nand U433 (N_433,In_173,In_127);
or U434 (N_434,In_21,In_84);
nor U435 (N_435,In_336,In_175);
or U436 (N_436,In_120,In_197);
nand U437 (N_437,In_81,In_429);
and U438 (N_438,In_335,In_408);
nor U439 (N_439,In_373,In_492);
and U440 (N_440,In_195,In_285);
nor U441 (N_441,In_400,In_433);
or U442 (N_442,In_494,In_153);
nand U443 (N_443,In_419,In_7);
and U444 (N_444,In_423,In_199);
nand U445 (N_445,In_125,In_45);
nor U446 (N_446,In_137,In_114);
nand U447 (N_447,In_186,In_114);
nor U448 (N_448,In_270,In_24);
nor U449 (N_449,In_381,In_250);
nor U450 (N_450,In_260,In_252);
nor U451 (N_451,In_499,In_255);
nor U452 (N_452,In_190,In_483);
nor U453 (N_453,In_138,In_139);
or U454 (N_454,In_145,In_382);
nand U455 (N_455,In_386,In_252);
or U456 (N_456,In_421,In_454);
nand U457 (N_457,In_469,In_172);
nor U458 (N_458,In_406,In_222);
nand U459 (N_459,In_117,In_289);
and U460 (N_460,In_132,In_29);
or U461 (N_461,In_3,In_437);
and U462 (N_462,In_322,In_41);
and U463 (N_463,In_342,In_444);
xor U464 (N_464,In_264,In_58);
nor U465 (N_465,In_238,In_80);
nand U466 (N_466,In_434,In_397);
and U467 (N_467,In_392,In_65);
and U468 (N_468,In_465,In_158);
xnor U469 (N_469,In_332,In_155);
and U470 (N_470,In_425,In_40);
and U471 (N_471,In_401,In_494);
and U472 (N_472,In_114,In_295);
or U473 (N_473,In_131,In_363);
xor U474 (N_474,In_496,In_255);
or U475 (N_475,In_315,In_159);
nor U476 (N_476,In_13,In_369);
or U477 (N_477,In_78,In_272);
nor U478 (N_478,In_110,In_400);
and U479 (N_479,In_140,In_238);
nor U480 (N_480,In_82,In_100);
or U481 (N_481,In_340,In_449);
nor U482 (N_482,In_111,In_163);
nand U483 (N_483,In_477,In_149);
or U484 (N_484,In_148,In_150);
nor U485 (N_485,In_473,In_164);
xnor U486 (N_486,In_287,In_198);
nand U487 (N_487,In_150,In_390);
nand U488 (N_488,In_391,In_363);
and U489 (N_489,In_1,In_450);
or U490 (N_490,In_86,In_80);
nand U491 (N_491,In_355,In_178);
nor U492 (N_492,In_261,In_78);
nand U493 (N_493,In_368,In_233);
or U494 (N_494,In_379,In_239);
or U495 (N_495,In_289,In_93);
nor U496 (N_496,In_467,In_265);
xor U497 (N_497,In_201,In_173);
nand U498 (N_498,In_101,In_428);
or U499 (N_499,In_385,In_273);
or U500 (N_500,N_263,N_464);
nand U501 (N_501,N_53,N_272);
nand U502 (N_502,N_148,N_219);
and U503 (N_503,N_349,N_155);
nand U504 (N_504,N_322,N_83);
and U505 (N_505,N_20,N_249);
or U506 (N_506,N_316,N_56);
nor U507 (N_507,N_454,N_361);
nand U508 (N_508,N_437,N_269);
nor U509 (N_509,N_352,N_23);
nor U510 (N_510,N_26,N_142);
nand U511 (N_511,N_439,N_154);
nor U512 (N_512,N_446,N_462);
or U513 (N_513,N_65,N_177);
or U514 (N_514,N_78,N_150);
nand U515 (N_515,N_164,N_206);
nand U516 (N_516,N_425,N_135);
and U517 (N_517,N_100,N_258);
xnor U518 (N_518,N_318,N_18);
and U519 (N_519,N_212,N_240);
or U520 (N_520,N_242,N_82);
or U521 (N_521,N_160,N_239);
and U522 (N_522,N_119,N_41);
nor U523 (N_523,N_88,N_380);
or U524 (N_524,N_338,N_185);
and U525 (N_525,N_441,N_399);
nor U526 (N_526,N_490,N_93);
nand U527 (N_527,N_336,N_398);
or U528 (N_528,N_77,N_59);
and U529 (N_529,N_278,N_498);
nor U530 (N_530,N_294,N_482);
nand U531 (N_531,N_205,N_444);
xnor U532 (N_532,N_51,N_25);
or U533 (N_533,N_306,N_410);
nor U534 (N_534,N_492,N_428);
nor U535 (N_535,N_459,N_286);
nand U536 (N_536,N_46,N_408);
or U537 (N_537,N_394,N_447);
nor U538 (N_538,N_98,N_369);
or U539 (N_539,N_213,N_268);
nor U540 (N_540,N_413,N_94);
nor U541 (N_541,N_404,N_167);
nand U542 (N_542,N_16,N_378);
nor U543 (N_543,N_309,N_126);
or U544 (N_544,N_234,N_442);
nand U545 (N_545,N_97,N_312);
nand U546 (N_546,N_305,N_431);
xor U547 (N_547,N_334,N_128);
nand U548 (N_548,N_270,N_450);
or U549 (N_549,N_362,N_189);
or U550 (N_550,N_191,N_427);
xnor U551 (N_551,N_342,N_6);
nand U552 (N_552,N_114,N_455);
and U553 (N_553,N_124,N_477);
or U554 (N_554,N_147,N_152);
nand U555 (N_555,N_19,N_196);
nand U556 (N_556,N_420,N_344);
and U557 (N_557,N_287,N_480);
or U558 (N_558,N_58,N_143);
nand U559 (N_559,N_329,N_434);
and U560 (N_560,N_472,N_71);
nor U561 (N_561,N_445,N_357);
or U562 (N_562,N_188,N_491);
xnor U563 (N_563,N_17,N_111);
nand U564 (N_564,N_350,N_300);
and U565 (N_565,N_359,N_421);
or U566 (N_566,N_488,N_192);
xor U567 (N_567,N_168,N_245);
and U568 (N_568,N_202,N_130);
or U569 (N_569,N_400,N_220);
or U570 (N_570,N_366,N_264);
or U571 (N_571,N_418,N_273);
or U572 (N_572,N_481,N_495);
and U573 (N_573,N_304,N_162);
or U574 (N_574,N_463,N_232);
or U575 (N_575,N_9,N_303);
nor U576 (N_576,N_393,N_457);
or U577 (N_577,N_64,N_422);
nand U578 (N_578,N_458,N_34);
nor U579 (N_579,N_499,N_214);
nor U580 (N_580,N_317,N_370);
nor U581 (N_581,N_365,N_190);
xor U582 (N_582,N_251,N_341);
xnor U583 (N_583,N_123,N_243);
nor U584 (N_584,N_324,N_246);
nor U585 (N_585,N_260,N_487);
nand U586 (N_586,N_103,N_347);
and U587 (N_587,N_426,N_440);
nand U588 (N_588,N_435,N_112);
nand U589 (N_589,N_416,N_63);
nor U590 (N_590,N_368,N_384);
or U591 (N_591,N_346,N_382);
and U592 (N_592,N_397,N_2);
nand U593 (N_593,N_43,N_301);
nand U594 (N_594,N_265,N_238);
nand U595 (N_595,N_283,N_390);
nor U596 (N_596,N_121,N_171);
or U597 (N_597,N_35,N_372);
nor U598 (N_598,N_424,N_153);
nor U599 (N_599,N_96,N_113);
or U600 (N_600,N_308,N_37);
nor U601 (N_601,N_320,N_101);
or U602 (N_602,N_335,N_351);
or U603 (N_603,N_348,N_62);
or U604 (N_604,N_118,N_178);
nand U605 (N_605,N_373,N_307);
nand U606 (N_606,N_173,N_227);
nor U607 (N_607,N_356,N_201);
nor U608 (N_608,N_337,N_129);
nand U609 (N_609,N_292,N_222);
nand U610 (N_610,N_131,N_267);
nor U611 (N_611,N_248,N_250);
nand U612 (N_612,N_208,N_451);
nor U613 (N_613,N_45,N_470);
nor U614 (N_614,N_453,N_132);
and U615 (N_615,N_471,N_375);
or U616 (N_616,N_266,N_279);
or U617 (N_617,N_169,N_289);
or U618 (N_618,N_314,N_414);
nor U619 (N_619,N_186,N_49);
nor U620 (N_620,N_354,N_387);
and U621 (N_621,N_383,N_407);
nor U622 (N_622,N_438,N_215);
nand U623 (N_623,N_31,N_313);
nand U624 (N_624,N_449,N_494);
or U625 (N_625,N_330,N_8);
and U626 (N_626,N_187,N_325);
xnor U627 (N_627,N_194,N_221);
nor U628 (N_628,N_10,N_180);
or U629 (N_629,N_137,N_237);
xor U630 (N_630,N_381,N_75);
and U631 (N_631,N_203,N_298);
and U632 (N_632,N_281,N_328);
or U633 (N_633,N_211,N_469);
and U634 (N_634,N_315,N_133);
or U635 (N_635,N_66,N_15);
and U636 (N_636,N_376,N_30);
xnor U637 (N_637,N_299,N_106);
or U638 (N_638,N_417,N_271);
or U639 (N_639,N_385,N_109);
nand U640 (N_640,N_38,N_290);
or U641 (N_641,N_388,N_403);
or U642 (N_642,N_448,N_149);
or U643 (N_643,N_339,N_332);
and U644 (N_644,N_467,N_419);
and U645 (N_645,N_92,N_36);
nor U646 (N_646,N_40,N_433);
nand U647 (N_647,N_236,N_183);
nand U648 (N_648,N_172,N_497);
and U649 (N_649,N_331,N_345);
nand U650 (N_650,N_193,N_430);
xnor U651 (N_651,N_468,N_379);
nor U652 (N_652,N_99,N_116);
or U653 (N_653,N_0,N_218);
nor U654 (N_654,N_184,N_395);
nand U655 (N_655,N_241,N_415);
or U656 (N_656,N_117,N_364);
and U657 (N_657,N_4,N_355);
xnor U658 (N_658,N_224,N_412);
nor U659 (N_659,N_76,N_443);
nor U660 (N_660,N_29,N_138);
or U661 (N_661,N_12,N_174);
and U662 (N_662,N_200,N_209);
and U663 (N_663,N_274,N_89);
nand U664 (N_664,N_198,N_52);
or U665 (N_665,N_353,N_108);
nand U666 (N_666,N_24,N_87);
nand U667 (N_667,N_295,N_493);
nand U668 (N_668,N_343,N_73);
nand U669 (N_669,N_229,N_466);
and U670 (N_670,N_14,N_217);
and U671 (N_671,N_296,N_120);
and U672 (N_672,N_33,N_166);
and U673 (N_673,N_310,N_207);
and U674 (N_674,N_105,N_401);
nand U675 (N_675,N_68,N_473);
or U676 (N_676,N_91,N_452);
nor U677 (N_677,N_39,N_107);
nor U678 (N_678,N_489,N_474);
nor U679 (N_679,N_85,N_80);
nand U680 (N_680,N_284,N_157);
or U681 (N_681,N_475,N_282);
and U682 (N_682,N_277,N_140);
and U683 (N_683,N_371,N_275);
or U684 (N_684,N_363,N_392);
or U685 (N_685,N_461,N_326);
or U686 (N_686,N_297,N_476);
and U687 (N_687,N_262,N_389);
and U688 (N_688,N_141,N_84);
xnor U689 (N_689,N_293,N_159);
nor U690 (N_690,N_195,N_67);
nor U691 (N_691,N_161,N_235);
nor U692 (N_692,N_176,N_86);
or U693 (N_693,N_69,N_57);
nor U694 (N_694,N_7,N_146);
nand U695 (N_695,N_429,N_47);
xnor U696 (N_696,N_170,N_483);
and U697 (N_697,N_115,N_230);
nor U698 (N_698,N_197,N_479);
or U699 (N_699,N_102,N_406);
nor U700 (N_700,N_386,N_233);
or U701 (N_701,N_456,N_90);
and U702 (N_702,N_391,N_151);
and U703 (N_703,N_55,N_311);
or U704 (N_704,N_175,N_210);
nor U705 (N_705,N_374,N_5);
and U706 (N_706,N_134,N_228);
and U707 (N_707,N_436,N_110);
and U708 (N_708,N_32,N_156);
nor U709 (N_709,N_42,N_259);
nand U710 (N_710,N_253,N_223);
nor U711 (N_711,N_405,N_13);
nand U712 (N_712,N_225,N_199);
nor U713 (N_713,N_122,N_104);
and U714 (N_714,N_396,N_165);
or U715 (N_715,N_261,N_81);
nand U716 (N_716,N_61,N_484);
nand U717 (N_717,N_44,N_163);
or U718 (N_718,N_145,N_333);
or U719 (N_719,N_244,N_285);
and U720 (N_720,N_280,N_321);
or U721 (N_721,N_423,N_252);
nor U722 (N_722,N_247,N_340);
nor U723 (N_723,N_1,N_79);
nand U724 (N_724,N_496,N_72);
and U725 (N_725,N_276,N_367);
or U726 (N_726,N_358,N_60);
and U727 (N_727,N_179,N_27);
and U728 (N_728,N_257,N_139);
nor U729 (N_729,N_256,N_54);
or U730 (N_730,N_432,N_70);
nor U731 (N_731,N_182,N_323);
nand U732 (N_732,N_409,N_21);
or U733 (N_733,N_158,N_3);
or U734 (N_734,N_22,N_327);
nor U735 (N_735,N_28,N_136);
nand U736 (N_736,N_204,N_255);
or U737 (N_737,N_50,N_302);
or U738 (N_738,N_377,N_216);
xnor U739 (N_739,N_11,N_95);
nor U740 (N_740,N_48,N_402);
nor U741 (N_741,N_254,N_319);
nor U742 (N_742,N_181,N_127);
or U743 (N_743,N_486,N_485);
or U744 (N_744,N_74,N_288);
nor U745 (N_745,N_226,N_478);
nor U746 (N_746,N_465,N_460);
xor U747 (N_747,N_125,N_411);
or U748 (N_748,N_360,N_291);
or U749 (N_749,N_144,N_231);
or U750 (N_750,N_70,N_484);
nor U751 (N_751,N_172,N_53);
xor U752 (N_752,N_161,N_392);
and U753 (N_753,N_494,N_240);
or U754 (N_754,N_160,N_209);
nor U755 (N_755,N_2,N_17);
nand U756 (N_756,N_64,N_126);
and U757 (N_757,N_214,N_102);
xor U758 (N_758,N_141,N_368);
nand U759 (N_759,N_115,N_177);
nand U760 (N_760,N_46,N_24);
or U761 (N_761,N_392,N_499);
nor U762 (N_762,N_148,N_104);
or U763 (N_763,N_417,N_378);
and U764 (N_764,N_46,N_417);
or U765 (N_765,N_392,N_397);
xor U766 (N_766,N_422,N_338);
xnor U767 (N_767,N_386,N_131);
or U768 (N_768,N_418,N_243);
or U769 (N_769,N_203,N_242);
nand U770 (N_770,N_86,N_136);
nor U771 (N_771,N_291,N_224);
or U772 (N_772,N_457,N_438);
nor U773 (N_773,N_50,N_301);
and U774 (N_774,N_70,N_402);
and U775 (N_775,N_38,N_45);
and U776 (N_776,N_261,N_7);
and U777 (N_777,N_382,N_404);
or U778 (N_778,N_98,N_120);
and U779 (N_779,N_245,N_219);
and U780 (N_780,N_103,N_349);
or U781 (N_781,N_282,N_462);
and U782 (N_782,N_146,N_303);
and U783 (N_783,N_180,N_189);
and U784 (N_784,N_262,N_122);
and U785 (N_785,N_76,N_270);
or U786 (N_786,N_491,N_258);
xnor U787 (N_787,N_100,N_218);
nor U788 (N_788,N_213,N_27);
or U789 (N_789,N_252,N_310);
nor U790 (N_790,N_374,N_49);
nand U791 (N_791,N_167,N_367);
nor U792 (N_792,N_49,N_63);
nand U793 (N_793,N_268,N_9);
nor U794 (N_794,N_293,N_151);
nand U795 (N_795,N_186,N_260);
xor U796 (N_796,N_78,N_361);
xor U797 (N_797,N_465,N_84);
nor U798 (N_798,N_471,N_486);
or U799 (N_799,N_349,N_11);
nor U800 (N_800,N_388,N_464);
nor U801 (N_801,N_368,N_341);
nand U802 (N_802,N_269,N_238);
or U803 (N_803,N_201,N_274);
or U804 (N_804,N_369,N_119);
or U805 (N_805,N_167,N_405);
or U806 (N_806,N_84,N_96);
nand U807 (N_807,N_131,N_201);
and U808 (N_808,N_256,N_464);
or U809 (N_809,N_209,N_272);
and U810 (N_810,N_80,N_499);
xor U811 (N_811,N_382,N_344);
nand U812 (N_812,N_96,N_67);
nor U813 (N_813,N_122,N_376);
nand U814 (N_814,N_270,N_96);
and U815 (N_815,N_91,N_283);
nand U816 (N_816,N_164,N_430);
nor U817 (N_817,N_287,N_188);
and U818 (N_818,N_338,N_290);
nor U819 (N_819,N_30,N_240);
and U820 (N_820,N_242,N_63);
or U821 (N_821,N_131,N_341);
nand U822 (N_822,N_263,N_41);
and U823 (N_823,N_315,N_294);
or U824 (N_824,N_69,N_250);
xor U825 (N_825,N_146,N_473);
nand U826 (N_826,N_332,N_223);
nor U827 (N_827,N_313,N_296);
nand U828 (N_828,N_440,N_189);
or U829 (N_829,N_192,N_102);
or U830 (N_830,N_271,N_266);
nor U831 (N_831,N_44,N_5);
or U832 (N_832,N_340,N_114);
or U833 (N_833,N_493,N_446);
nand U834 (N_834,N_494,N_239);
nor U835 (N_835,N_194,N_337);
or U836 (N_836,N_179,N_228);
nor U837 (N_837,N_44,N_90);
nor U838 (N_838,N_294,N_53);
or U839 (N_839,N_59,N_427);
nor U840 (N_840,N_462,N_423);
and U841 (N_841,N_64,N_17);
or U842 (N_842,N_30,N_303);
xor U843 (N_843,N_295,N_291);
or U844 (N_844,N_409,N_375);
nor U845 (N_845,N_471,N_272);
nand U846 (N_846,N_437,N_76);
and U847 (N_847,N_463,N_347);
nand U848 (N_848,N_179,N_243);
nand U849 (N_849,N_407,N_379);
nand U850 (N_850,N_366,N_136);
nor U851 (N_851,N_450,N_343);
and U852 (N_852,N_491,N_486);
and U853 (N_853,N_488,N_180);
xor U854 (N_854,N_342,N_447);
or U855 (N_855,N_67,N_212);
or U856 (N_856,N_189,N_377);
or U857 (N_857,N_191,N_320);
nor U858 (N_858,N_360,N_23);
and U859 (N_859,N_344,N_95);
nand U860 (N_860,N_381,N_129);
nor U861 (N_861,N_357,N_429);
and U862 (N_862,N_213,N_120);
nor U863 (N_863,N_47,N_112);
or U864 (N_864,N_211,N_490);
and U865 (N_865,N_104,N_159);
nand U866 (N_866,N_101,N_392);
nand U867 (N_867,N_458,N_436);
nor U868 (N_868,N_312,N_65);
nand U869 (N_869,N_410,N_101);
nand U870 (N_870,N_382,N_302);
xor U871 (N_871,N_14,N_260);
nand U872 (N_872,N_155,N_401);
nand U873 (N_873,N_331,N_14);
xnor U874 (N_874,N_410,N_328);
nor U875 (N_875,N_50,N_480);
and U876 (N_876,N_304,N_310);
nand U877 (N_877,N_444,N_307);
and U878 (N_878,N_256,N_159);
or U879 (N_879,N_477,N_71);
nand U880 (N_880,N_108,N_461);
nor U881 (N_881,N_163,N_433);
and U882 (N_882,N_286,N_154);
and U883 (N_883,N_208,N_318);
and U884 (N_884,N_162,N_351);
nor U885 (N_885,N_169,N_444);
and U886 (N_886,N_459,N_163);
and U887 (N_887,N_483,N_44);
and U888 (N_888,N_279,N_109);
xor U889 (N_889,N_431,N_395);
or U890 (N_890,N_230,N_231);
and U891 (N_891,N_245,N_170);
nand U892 (N_892,N_139,N_400);
nand U893 (N_893,N_213,N_57);
nand U894 (N_894,N_256,N_1);
nor U895 (N_895,N_477,N_399);
and U896 (N_896,N_451,N_437);
and U897 (N_897,N_430,N_497);
or U898 (N_898,N_151,N_458);
nor U899 (N_899,N_184,N_103);
or U900 (N_900,N_423,N_83);
nor U901 (N_901,N_331,N_24);
nor U902 (N_902,N_205,N_319);
and U903 (N_903,N_230,N_381);
and U904 (N_904,N_197,N_225);
nor U905 (N_905,N_109,N_24);
nor U906 (N_906,N_319,N_342);
and U907 (N_907,N_487,N_12);
nor U908 (N_908,N_131,N_491);
nor U909 (N_909,N_210,N_387);
nor U910 (N_910,N_357,N_145);
and U911 (N_911,N_103,N_376);
and U912 (N_912,N_375,N_68);
nor U913 (N_913,N_262,N_251);
xor U914 (N_914,N_54,N_210);
nand U915 (N_915,N_377,N_35);
or U916 (N_916,N_406,N_411);
nand U917 (N_917,N_214,N_168);
and U918 (N_918,N_107,N_467);
nor U919 (N_919,N_169,N_373);
and U920 (N_920,N_435,N_89);
or U921 (N_921,N_307,N_55);
nor U922 (N_922,N_339,N_271);
or U923 (N_923,N_324,N_390);
or U924 (N_924,N_70,N_450);
or U925 (N_925,N_120,N_38);
nor U926 (N_926,N_424,N_190);
nor U927 (N_927,N_397,N_296);
xnor U928 (N_928,N_48,N_135);
nor U929 (N_929,N_212,N_296);
and U930 (N_930,N_225,N_260);
nor U931 (N_931,N_262,N_384);
nor U932 (N_932,N_361,N_270);
nand U933 (N_933,N_441,N_298);
nand U934 (N_934,N_431,N_481);
or U935 (N_935,N_82,N_152);
and U936 (N_936,N_174,N_30);
nor U937 (N_937,N_400,N_80);
and U938 (N_938,N_343,N_362);
or U939 (N_939,N_373,N_485);
nor U940 (N_940,N_354,N_312);
or U941 (N_941,N_458,N_470);
nand U942 (N_942,N_107,N_103);
nor U943 (N_943,N_97,N_335);
and U944 (N_944,N_281,N_309);
nand U945 (N_945,N_449,N_214);
xnor U946 (N_946,N_462,N_322);
or U947 (N_947,N_30,N_304);
nand U948 (N_948,N_170,N_488);
or U949 (N_949,N_249,N_285);
nand U950 (N_950,N_310,N_65);
xor U951 (N_951,N_454,N_89);
and U952 (N_952,N_286,N_280);
and U953 (N_953,N_276,N_158);
or U954 (N_954,N_283,N_34);
nand U955 (N_955,N_91,N_332);
or U956 (N_956,N_335,N_157);
and U957 (N_957,N_435,N_309);
and U958 (N_958,N_37,N_433);
and U959 (N_959,N_311,N_397);
nor U960 (N_960,N_388,N_261);
nand U961 (N_961,N_229,N_338);
or U962 (N_962,N_353,N_157);
or U963 (N_963,N_344,N_339);
and U964 (N_964,N_233,N_35);
and U965 (N_965,N_103,N_327);
and U966 (N_966,N_391,N_456);
nand U967 (N_967,N_379,N_93);
nor U968 (N_968,N_121,N_241);
nand U969 (N_969,N_268,N_47);
xnor U970 (N_970,N_112,N_292);
nand U971 (N_971,N_409,N_157);
nor U972 (N_972,N_382,N_170);
nand U973 (N_973,N_459,N_465);
nand U974 (N_974,N_54,N_391);
nand U975 (N_975,N_345,N_318);
and U976 (N_976,N_449,N_101);
and U977 (N_977,N_411,N_481);
or U978 (N_978,N_154,N_471);
xnor U979 (N_979,N_260,N_228);
nor U980 (N_980,N_19,N_276);
nor U981 (N_981,N_70,N_311);
and U982 (N_982,N_140,N_204);
and U983 (N_983,N_481,N_499);
or U984 (N_984,N_320,N_116);
nor U985 (N_985,N_398,N_428);
nor U986 (N_986,N_120,N_308);
or U987 (N_987,N_454,N_317);
nand U988 (N_988,N_107,N_105);
and U989 (N_989,N_442,N_333);
and U990 (N_990,N_456,N_179);
nand U991 (N_991,N_364,N_295);
and U992 (N_992,N_180,N_85);
and U993 (N_993,N_242,N_447);
nor U994 (N_994,N_445,N_421);
nand U995 (N_995,N_52,N_480);
nand U996 (N_996,N_136,N_26);
or U997 (N_997,N_13,N_35);
nand U998 (N_998,N_161,N_19);
nor U999 (N_999,N_35,N_19);
and U1000 (N_1000,N_762,N_816);
nand U1001 (N_1001,N_931,N_884);
or U1002 (N_1002,N_834,N_589);
nor U1003 (N_1003,N_768,N_627);
xor U1004 (N_1004,N_876,N_728);
nand U1005 (N_1005,N_909,N_915);
or U1006 (N_1006,N_978,N_901);
and U1007 (N_1007,N_656,N_775);
nand U1008 (N_1008,N_683,N_546);
nand U1009 (N_1009,N_729,N_996);
nand U1010 (N_1010,N_992,N_612);
nor U1011 (N_1011,N_899,N_894);
nor U1012 (N_1012,N_934,N_848);
nor U1013 (N_1013,N_817,N_935);
nand U1014 (N_1014,N_942,N_639);
and U1015 (N_1015,N_515,N_549);
or U1016 (N_1016,N_688,N_970);
or U1017 (N_1017,N_785,N_720);
nand U1018 (N_1018,N_766,N_773);
and U1019 (N_1019,N_708,N_622);
or U1020 (N_1020,N_841,N_780);
and U1021 (N_1021,N_822,N_913);
and U1022 (N_1022,N_677,N_956);
or U1023 (N_1023,N_795,N_937);
or U1024 (N_1024,N_593,N_799);
and U1025 (N_1025,N_678,N_797);
xnor U1026 (N_1026,N_916,N_505);
nor U1027 (N_1027,N_924,N_998);
xnor U1028 (N_1028,N_990,N_824);
and U1029 (N_1029,N_890,N_953);
xnor U1030 (N_1030,N_947,N_682);
or U1031 (N_1031,N_963,N_642);
nand U1032 (N_1032,N_705,N_929);
nand U1033 (N_1033,N_769,N_553);
nor U1034 (N_1034,N_845,N_840);
xor U1035 (N_1035,N_760,N_551);
nand U1036 (N_1036,N_662,N_626);
and U1037 (N_1037,N_812,N_644);
nand U1038 (N_1038,N_865,N_857);
and U1039 (N_1039,N_689,N_623);
and U1040 (N_1040,N_727,N_987);
nand U1041 (N_1041,N_735,N_741);
nand U1042 (N_1042,N_684,N_950);
xnor U1043 (N_1043,N_617,N_979);
nor U1044 (N_1044,N_949,N_738);
and U1045 (N_1045,N_534,N_779);
nor U1046 (N_1046,N_517,N_648);
or U1047 (N_1047,N_791,N_667);
nor U1048 (N_1048,N_844,N_948);
xor U1049 (N_1049,N_601,N_615);
nor U1050 (N_1050,N_701,N_962);
or U1051 (N_1051,N_744,N_896);
nand U1052 (N_1052,N_582,N_930);
nor U1053 (N_1053,N_945,N_537);
or U1054 (N_1054,N_620,N_995);
or U1055 (N_1055,N_540,N_629);
nand U1056 (N_1056,N_800,N_763);
or U1057 (N_1057,N_568,N_693);
xor U1058 (N_1058,N_983,N_597);
nand U1059 (N_1059,N_842,N_887);
or U1060 (N_1060,N_831,N_634);
and U1061 (N_1061,N_714,N_628);
or U1062 (N_1062,N_837,N_721);
xor U1063 (N_1063,N_751,N_508);
or U1064 (N_1064,N_843,N_655);
or U1065 (N_1065,N_801,N_715);
nor U1066 (N_1066,N_621,N_969);
or U1067 (N_1067,N_748,N_658);
nand U1068 (N_1068,N_700,N_527);
or U1069 (N_1069,N_521,N_793);
or U1070 (N_1070,N_681,N_624);
or U1071 (N_1071,N_679,N_997);
nand U1072 (N_1072,N_504,N_587);
nor U1073 (N_1073,N_570,N_828);
and U1074 (N_1074,N_509,N_805);
and U1075 (N_1075,N_820,N_988);
or U1076 (N_1076,N_923,N_783);
nor U1077 (N_1077,N_854,N_583);
nand U1078 (N_1078,N_758,N_588);
xor U1079 (N_1079,N_788,N_542);
and U1080 (N_1080,N_900,N_567);
and U1081 (N_1081,N_502,N_918);
nor U1082 (N_1082,N_859,N_984);
and U1083 (N_1083,N_586,N_936);
and U1084 (N_1084,N_807,N_737);
nand U1085 (N_1085,N_536,N_754);
or U1086 (N_1086,N_882,N_591);
or U1087 (N_1087,N_577,N_647);
nand U1088 (N_1088,N_966,N_977);
or U1089 (N_1089,N_552,N_993);
nor U1090 (N_1090,N_631,N_740);
and U1091 (N_1091,N_922,N_767);
nand U1092 (N_1092,N_618,N_921);
and U1093 (N_1093,N_892,N_897);
xnor U1094 (N_1094,N_704,N_598);
xor U1095 (N_1095,N_860,N_514);
nor U1096 (N_1096,N_917,N_566);
or U1097 (N_1097,N_630,N_616);
or U1098 (N_1098,N_671,N_723);
and U1099 (N_1099,N_874,N_964);
nor U1100 (N_1100,N_852,N_666);
or U1101 (N_1101,N_559,N_725);
xor U1102 (N_1102,N_694,N_895);
nor U1103 (N_1103,N_604,N_712);
or U1104 (N_1104,N_510,N_823);
or U1105 (N_1105,N_782,N_975);
nand U1106 (N_1106,N_753,N_646);
xor U1107 (N_1107,N_849,N_872);
and U1108 (N_1108,N_886,N_933);
xnor U1109 (N_1109,N_562,N_599);
or U1110 (N_1110,N_529,N_839);
nor U1111 (N_1111,N_576,N_742);
xor U1112 (N_1112,N_802,N_806);
and U1113 (N_1113,N_611,N_919);
nor U1114 (N_1114,N_691,N_573);
or U1115 (N_1115,N_600,N_696);
nand U1116 (N_1116,N_520,N_524);
and U1117 (N_1117,N_981,N_713);
nand U1118 (N_1118,N_770,N_608);
or U1119 (N_1119,N_905,N_675);
and U1120 (N_1120,N_784,N_994);
and U1121 (N_1121,N_833,N_657);
or U1122 (N_1122,N_660,N_986);
xor U1123 (N_1123,N_500,N_703);
nor U1124 (N_1124,N_563,N_716);
nand U1125 (N_1125,N_697,N_665);
nand U1126 (N_1126,N_757,N_939);
nand U1127 (N_1127,N_745,N_506);
nand U1128 (N_1128,N_847,N_541);
or U1129 (N_1129,N_771,N_804);
xnor U1130 (N_1130,N_717,N_813);
and U1131 (N_1131,N_571,N_535);
or U1132 (N_1132,N_772,N_965);
nand U1133 (N_1133,N_761,N_580);
or U1134 (N_1134,N_796,N_528);
nor U1135 (N_1135,N_825,N_991);
and U1136 (N_1136,N_569,N_554);
and U1137 (N_1137,N_853,N_814);
xor U1138 (N_1138,N_878,N_522);
xnor U1139 (N_1139,N_989,N_869);
and U1140 (N_1140,N_827,N_596);
and U1141 (N_1141,N_908,N_579);
nor U1142 (N_1142,N_513,N_850);
nand U1143 (N_1143,N_883,N_651);
and U1144 (N_1144,N_669,N_609);
nand U1145 (N_1145,N_533,N_578);
nand U1146 (N_1146,N_531,N_759);
xor U1147 (N_1147,N_711,N_706);
nand U1148 (N_1148,N_614,N_652);
or U1149 (N_1149,N_695,N_523);
nand U1150 (N_1150,N_507,N_879);
and U1151 (N_1151,N_707,N_889);
nand U1152 (N_1152,N_613,N_556);
and U1153 (N_1153,N_815,N_592);
nor U1154 (N_1154,N_764,N_643);
or U1155 (N_1155,N_584,N_606);
and U1156 (N_1156,N_856,N_687);
and U1157 (N_1157,N_794,N_654);
and U1158 (N_1158,N_602,N_944);
and U1159 (N_1159,N_550,N_982);
or U1160 (N_1160,N_544,N_603);
and U1161 (N_1161,N_855,N_972);
nand U1162 (N_1162,N_664,N_739);
or U1163 (N_1163,N_548,N_561);
xnor U1164 (N_1164,N_532,N_786);
and U1165 (N_1165,N_730,N_955);
and U1166 (N_1166,N_946,N_719);
nor U1167 (N_1167,N_893,N_838);
nand U1168 (N_1168,N_875,N_585);
and U1169 (N_1169,N_776,N_595);
and U1170 (N_1170,N_518,N_866);
nor U1171 (N_1171,N_932,N_685);
nor U1172 (N_1172,N_765,N_830);
xor U1173 (N_1173,N_575,N_752);
or U1174 (N_1174,N_891,N_526);
xnor U1175 (N_1175,N_558,N_726);
nor U1176 (N_1176,N_686,N_943);
nor U1177 (N_1177,N_709,N_871);
or U1178 (N_1178,N_952,N_951);
xnor U1179 (N_1179,N_906,N_590);
or U1180 (N_1180,N_904,N_787);
or U1181 (N_1181,N_680,N_818);
nand U1182 (N_1182,N_668,N_640);
nand U1183 (N_1183,N_503,N_867);
and U1184 (N_1184,N_861,N_722);
and U1185 (N_1185,N_826,N_958);
or U1186 (N_1186,N_985,N_663);
nor U1187 (N_1187,N_625,N_974);
and U1188 (N_1188,N_880,N_954);
nor U1189 (N_1189,N_755,N_911);
nand U1190 (N_1190,N_961,N_574);
nand U1191 (N_1191,N_732,N_545);
nand U1192 (N_1192,N_710,N_750);
xor U1193 (N_1193,N_543,N_690);
nor U1194 (N_1194,N_976,N_938);
nand U1195 (N_1195,N_835,N_692);
nor U1196 (N_1196,N_743,N_888);
and U1197 (N_1197,N_925,N_798);
and U1198 (N_1198,N_594,N_810);
nand U1199 (N_1199,N_698,N_980);
xnor U1200 (N_1200,N_610,N_530);
and U1201 (N_1201,N_957,N_724);
or U1202 (N_1202,N_516,N_659);
nand U1203 (N_1203,N_650,N_676);
or U1204 (N_1204,N_898,N_968);
and U1205 (N_1205,N_885,N_653);
or U1206 (N_1206,N_778,N_673);
nor U1207 (N_1207,N_519,N_846);
and U1208 (N_1208,N_699,N_512);
nor U1209 (N_1209,N_999,N_547);
nand U1210 (N_1210,N_809,N_907);
nor U1211 (N_1211,N_836,N_511);
nand U1212 (N_1212,N_862,N_649);
xor U1213 (N_1213,N_973,N_674);
or U1214 (N_1214,N_557,N_636);
nand U1215 (N_1215,N_774,N_736);
xor U1216 (N_1216,N_959,N_638);
nand U1217 (N_1217,N_821,N_863);
and U1218 (N_1218,N_877,N_781);
or U1219 (N_1219,N_501,N_927);
nand U1220 (N_1220,N_555,N_910);
and U1221 (N_1221,N_718,N_637);
nor U1222 (N_1222,N_733,N_565);
nand U1223 (N_1223,N_912,N_581);
or U1224 (N_1224,N_731,N_971);
and U1225 (N_1225,N_756,N_564);
nor U1226 (N_1226,N_633,N_645);
nand U1227 (N_1227,N_790,N_632);
nand U1228 (N_1228,N_819,N_572);
nor U1229 (N_1229,N_525,N_539);
and U1230 (N_1230,N_881,N_928);
nor U1231 (N_1231,N_873,N_941);
and U1232 (N_1232,N_864,N_870);
or U1233 (N_1233,N_670,N_641);
nor U1234 (N_1234,N_808,N_747);
nand U1235 (N_1235,N_789,N_607);
or U1236 (N_1236,N_926,N_777);
nor U1237 (N_1237,N_903,N_914);
nor U1238 (N_1238,N_749,N_868);
or U1239 (N_1239,N_605,N_538);
nor U1240 (N_1240,N_635,N_858);
nand U1241 (N_1241,N_734,N_702);
or U1242 (N_1242,N_792,N_920);
nor U1243 (N_1243,N_560,N_902);
nor U1244 (N_1244,N_661,N_746);
or U1245 (N_1245,N_803,N_967);
nor U1246 (N_1246,N_851,N_940);
nand U1247 (N_1247,N_811,N_960);
or U1248 (N_1248,N_832,N_619);
nor U1249 (N_1249,N_672,N_829);
nand U1250 (N_1250,N_885,N_884);
or U1251 (N_1251,N_760,N_556);
or U1252 (N_1252,N_653,N_553);
or U1253 (N_1253,N_809,N_975);
nor U1254 (N_1254,N_577,N_854);
and U1255 (N_1255,N_984,N_666);
and U1256 (N_1256,N_949,N_735);
and U1257 (N_1257,N_632,N_830);
or U1258 (N_1258,N_729,N_630);
or U1259 (N_1259,N_658,N_549);
and U1260 (N_1260,N_567,N_605);
or U1261 (N_1261,N_795,N_837);
nor U1262 (N_1262,N_763,N_508);
nor U1263 (N_1263,N_564,N_597);
nor U1264 (N_1264,N_617,N_856);
nor U1265 (N_1265,N_524,N_779);
and U1266 (N_1266,N_591,N_640);
and U1267 (N_1267,N_902,N_519);
or U1268 (N_1268,N_806,N_582);
and U1269 (N_1269,N_709,N_637);
nand U1270 (N_1270,N_638,N_860);
or U1271 (N_1271,N_849,N_822);
and U1272 (N_1272,N_615,N_949);
or U1273 (N_1273,N_639,N_598);
nand U1274 (N_1274,N_531,N_586);
or U1275 (N_1275,N_715,N_552);
or U1276 (N_1276,N_818,N_649);
nand U1277 (N_1277,N_927,N_603);
or U1278 (N_1278,N_662,N_570);
and U1279 (N_1279,N_890,N_815);
nor U1280 (N_1280,N_626,N_759);
xnor U1281 (N_1281,N_760,N_614);
nand U1282 (N_1282,N_770,N_506);
nand U1283 (N_1283,N_577,N_670);
or U1284 (N_1284,N_881,N_707);
and U1285 (N_1285,N_879,N_963);
nor U1286 (N_1286,N_911,N_650);
or U1287 (N_1287,N_763,N_980);
and U1288 (N_1288,N_877,N_745);
or U1289 (N_1289,N_617,N_752);
nand U1290 (N_1290,N_759,N_793);
and U1291 (N_1291,N_700,N_519);
nand U1292 (N_1292,N_792,N_678);
nand U1293 (N_1293,N_657,N_599);
nand U1294 (N_1294,N_558,N_950);
or U1295 (N_1295,N_893,N_662);
and U1296 (N_1296,N_533,N_677);
xor U1297 (N_1297,N_695,N_702);
nand U1298 (N_1298,N_621,N_791);
and U1299 (N_1299,N_820,N_778);
xor U1300 (N_1300,N_878,N_871);
nand U1301 (N_1301,N_601,N_844);
and U1302 (N_1302,N_509,N_861);
and U1303 (N_1303,N_704,N_769);
nand U1304 (N_1304,N_547,N_610);
and U1305 (N_1305,N_663,N_822);
or U1306 (N_1306,N_584,N_508);
or U1307 (N_1307,N_802,N_919);
xnor U1308 (N_1308,N_861,N_923);
nand U1309 (N_1309,N_960,N_872);
nand U1310 (N_1310,N_925,N_957);
and U1311 (N_1311,N_797,N_973);
nor U1312 (N_1312,N_809,N_673);
or U1313 (N_1313,N_825,N_915);
nor U1314 (N_1314,N_527,N_873);
and U1315 (N_1315,N_602,N_567);
nor U1316 (N_1316,N_926,N_693);
nand U1317 (N_1317,N_806,N_786);
and U1318 (N_1318,N_835,N_621);
xnor U1319 (N_1319,N_913,N_622);
and U1320 (N_1320,N_574,N_827);
or U1321 (N_1321,N_709,N_769);
xnor U1322 (N_1322,N_793,N_943);
and U1323 (N_1323,N_873,N_623);
and U1324 (N_1324,N_956,N_632);
nand U1325 (N_1325,N_937,N_718);
nand U1326 (N_1326,N_910,N_991);
and U1327 (N_1327,N_673,N_709);
and U1328 (N_1328,N_664,N_722);
nor U1329 (N_1329,N_547,N_648);
and U1330 (N_1330,N_656,N_833);
nand U1331 (N_1331,N_971,N_509);
and U1332 (N_1332,N_897,N_736);
and U1333 (N_1333,N_712,N_747);
nand U1334 (N_1334,N_920,N_596);
nand U1335 (N_1335,N_568,N_893);
or U1336 (N_1336,N_923,N_876);
or U1337 (N_1337,N_944,N_608);
nor U1338 (N_1338,N_600,N_846);
xnor U1339 (N_1339,N_871,N_510);
nor U1340 (N_1340,N_589,N_977);
xnor U1341 (N_1341,N_870,N_807);
nand U1342 (N_1342,N_804,N_993);
nor U1343 (N_1343,N_901,N_645);
nand U1344 (N_1344,N_903,N_533);
nor U1345 (N_1345,N_732,N_638);
nor U1346 (N_1346,N_703,N_902);
and U1347 (N_1347,N_927,N_525);
or U1348 (N_1348,N_945,N_669);
nand U1349 (N_1349,N_682,N_915);
and U1350 (N_1350,N_654,N_979);
xnor U1351 (N_1351,N_589,N_710);
or U1352 (N_1352,N_619,N_992);
nor U1353 (N_1353,N_919,N_632);
nand U1354 (N_1354,N_705,N_662);
nor U1355 (N_1355,N_646,N_583);
or U1356 (N_1356,N_986,N_744);
nand U1357 (N_1357,N_955,N_737);
or U1358 (N_1358,N_830,N_545);
and U1359 (N_1359,N_530,N_942);
or U1360 (N_1360,N_708,N_939);
or U1361 (N_1361,N_877,N_827);
nor U1362 (N_1362,N_846,N_939);
or U1363 (N_1363,N_820,N_973);
or U1364 (N_1364,N_811,N_681);
and U1365 (N_1365,N_583,N_894);
nor U1366 (N_1366,N_676,N_658);
or U1367 (N_1367,N_625,N_514);
nor U1368 (N_1368,N_805,N_766);
and U1369 (N_1369,N_972,N_996);
and U1370 (N_1370,N_663,N_858);
nor U1371 (N_1371,N_946,N_981);
and U1372 (N_1372,N_525,N_900);
nand U1373 (N_1373,N_731,N_654);
xor U1374 (N_1374,N_537,N_613);
or U1375 (N_1375,N_841,N_852);
and U1376 (N_1376,N_605,N_924);
nor U1377 (N_1377,N_603,N_941);
or U1378 (N_1378,N_556,N_903);
nor U1379 (N_1379,N_881,N_991);
nor U1380 (N_1380,N_708,N_834);
and U1381 (N_1381,N_998,N_703);
or U1382 (N_1382,N_958,N_969);
nand U1383 (N_1383,N_508,N_687);
nand U1384 (N_1384,N_568,N_986);
nor U1385 (N_1385,N_740,N_674);
or U1386 (N_1386,N_535,N_811);
or U1387 (N_1387,N_589,N_633);
nand U1388 (N_1388,N_584,N_729);
nand U1389 (N_1389,N_629,N_537);
or U1390 (N_1390,N_566,N_914);
and U1391 (N_1391,N_852,N_574);
nand U1392 (N_1392,N_614,N_769);
or U1393 (N_1393,N_955,N_924);
or U1394 (N_1394,N_983,N_767);
nand U1395 (N_1395,N_942,N_712);
or U1396 (N_1396,N_576,N_517);
and U1397 (N_1397,N_700,N_893);
and U1398 (N_1398,N_676,N_549);
xor U1399 (N_1399,N_558,N_673);
and U1400 (N_1400,N_815,N_792);
nor U1401 (N_1401,N_826,N_585);
or U1402 (N_1402,N_783,N_581);
nor U1403 (N_1403,N_640,N_745);
nor U1404 (N_1404,N_985,N_846);
nor U1405 (N_1405,N_687,N_569);
or U1406 (N_1406,N_587,N_919);
or U1407 (N_1407,N_743,N_648);
nor U1408 (N_1408,N_651,N_688);
nor U1409 (N_1409,N_759,N_782);
or U1410 (N_1410,N_744,N_674);
nor U1411 (N_1411,N_852,N_928);
nor U1412 (N_1412,N_978,N_613);
nor U1413 (N_1413,N_954,N_534);
xor U1414 (N_1414,N_659,N_948);
or U1415 (N_1415,N_820,N_808);
and U1416 (N_1416,N_865,N_752);
and U1417 (N_1417,N_627,N_909);
and U1418 (N_1418,N_937,N_502);
nor U1419 (N_1419,N_609,N_784);
and U1420 (N_1420,N_669,N_519);
nand U1421 (N_1421,N_971,N_981);
and U1422 (N_1422,N_864,N_575);
or U1423 (N_1423,N_672,N_610);
nand U1424 (N_1424,N_523,N_551);
xor U1425 (N_1425,N_737,N_730);
nand U1426 (N_1426,N_554,N_966);
and U1427 (N_1427,N_524,N_832);
or U1428 (N_1428,N_740,N_761);
xor U1429 (N_1429,N_590,N_520);
and U1430 (N_1430,N_901,N_874);
nand U1431 (N_1431,N_759,N_677);
nand U1432 (N_1432,N_760,N_588);
xor U1433 (N_1433,N_679,N_809);
or U1434 (N_1434,N_579,N_957);
or U1435 (N_1435,N_721,N_826);
nand U1436 (N_1436,N_936,N_575);
nand U1437 (N_1437,N_950,N_848);
nand U1438 (N_1438,N_848,N_886);
xnor U1439 (N_1439,N_868,N_662);
nand U1440 (N_1440,N_850,N_507);
nand U1441 (N_1441,N_806,N_579);
nor U1442 (N_1442,N_556,N_502);
and U1443 (N_1443,N_779,N_973);
or U1444 (N_1444,N_776,N_750);
nand U1445 (N_1445,N_732,N_930);
or U1446 (N_1446,N_824,N_641);
or U1447 (N_1447,N_855,N_552);
nand U1448 (N_1448,N_626,N_849);
and U1449 (N_1449,N_672,N_995);
and U1450 (N_1450,N_549,N_525);
nand U1451 (N_1451,N_514,N_567);
nand U1452 (N_1452,N_503,N_868);
nand U1453 (N_1453,N_556,N_608);
xor U1454 (N_1454,N_619,N_788);
nand U1455 (N_1455,N_513,N_884);
nor U1456 (N_1456,N_583,N_746);
and U1457 (N_1457,N_835,N_924);
and U1458 (N_1458,N_575,N_686);
and U1459 (N_1459,N_846,N_602);
nand U1460 (N_1460,N_857,N_848);
and U1461 (N_1461,N_661,N_707);
or U1462 (N_1462,N_945,N_659);
nor U1463 (N_1463,N_950,N_656);
nor U1464 (N_1464,N_555,N_795);
or U1465 (N_1465,N_988,N_868);
nand U1466 (N_1466,N_712,N_597);
nand U1467 (N_1467,N_879,N_851);
or U1468 (N_1468,N_713,N_602);
and U1469 (N_1469,N_761,N_966);
xor U1470 (N_1470,N_515,N_712);
nor U1471 (N_1471,N_752,N_926);
and U1472 (N_1472,N_969,N_832);
nor U1473 (N_1473,N_980,N_744);
nand U1474 (N_1474,N_753,N_580);
nand U1475 (N_1475,N_875,N_583);
nor U1476 (N_1476,N_561,N_936);
nor U1477 (N_1477,N_986,N_842);
nor U1478 (N_1478,N_651,N_606);
nor U1479 (N_1479,N_587,N_514);
or U1480 (N_1480,N_627,N_817);
nand U1481 (N_1481,N_584,N_671);
nor U1482 (N_1482,N_612,N_874);
nor U1483 (N_1483,N_865,N_891);
nand U1484 (N_1484,N_888,N_930);
nand U1485 (N_1485,N_932,N_573);
xnor U1486 (N_1486,N_899,N_501);
and U1487 (N_1487,N_859,N_772);
nor U1488 (N_1488,N_739,N_514);
or U1489 (N_1489,N_769,N_541);
and U1490 (N_1490,N_686,N_939);
or U1491 (N_1491,N_961,N_701);
or U1492 (N_1492,N_667,N_548);
xnor U1493 (N_1493,N_573,N_930);
xnor U1494 (N_1494,N_755,N_614);
nand U1495 (N_1495,N_888,N_738);
nand U1496 (N_1496,N_605,N_552);
nor U1497 (N_1497,N_668,N_601);
or U1498 (N_1498,N_587,N_843);
nor U1499 (N_1499,N_623,N_755);
nor U1500 (N_1500,N_1056,N_1220);
nor U1501 (N_1501,N_1118,N_1017);
or U1502 (N_1502,N_1000,N_1120);
or U1503 (N_1503,N_1013,N_1351);
and U1504 (N_1504,N_1398,N_1063);
and U1505 (N_1505,N_1238,N_1306);
nand U1506 (N_1506,N_1083,N_1280);
and U1507 (N_1507,N_1248,N_1035);
and U1508 (N_1508,N_1284,N_1037);
nor U1509 (N_1509,N_1080,N_1146);
nor U1510 (N_1510,N_1036,N_1413);
nand U1511 (N_1511,N_1336,N_1138);
nand U1512 (N_1512,N_1365,N_1086);
nor U1513 (N_1513,N_1370,N_1444);
or U1514 (N_1514,N_1497,N_1340);
and U1515 (N_1515,N_1230,N_1414);
xor U1516 (N_1516,N_1430,N_1258);
nor U1517 (N_1517,N_1437,N_1202);
nor U1518 (N_1518,N_1117,N_1127);
nand U1519 (N_1519,N_1221,N_1331);
nand U1520 (N_1520,N_1304,N_1227);
nor U1521 (N_1521,N_1462,N_1344);
nor U1522 (N_1522,N_1463,N_1052);
nand U1523 (N_1523,N_1373,N_1456);
and U1524 (N_1524,N_1106,N_1379);
and U1525 (N_1525,N_1156,N_1267);
nand U1526 (N_1526,N_1183,N_1113);
xnor U1527 (N_1527,N_1493,N_1041);
nand U1528 (N_1528,N_1405,N_1049);
nor U1529 (N_1529,N_1428,N_1167);
nand U1530 (N_1530,N_1445,N_1194);
nor U1531 (N_1531,N_1421,N_1150);
or U1532 (N_1532,N_1476,N_1051);
and U1533 (N_1533,N_1261,N_1390);
nor U1534 (N_1534,N_1125,N_1378);
nor U1535 (N_1535,N_1326,N_1459);
or U1536 (N_1536,N_1122,N_1406);
nor U1537 (N_1537,N_1403,N_1498);
and U1538 (N_1538,N_1188,N_1055);
or U1539 (N_1539,N_1019,N_1020);
and U1540 (N_1540,N_1341,N_1302);
and U1541 (N_1541,N_1237,N_1287);
nor U1542 (N_1542,N_1468,N_1333);
and U1543 (N_1543,N_1047,N_1295);
nor U1544 (N_1544,N_1093,N_1256);
nor U1545 (N_1545,N_1193,N_1027);
and U1546 (N_1546,N_1034,N_1288);
nor U1547 (N_1547,N_1165,N_1148);
nor U1548 (N_1548,N_1025,N_1099);
nor U1549 (N_1549,N_1350,N_1422);
and U1550 (N_1550,N_1451,N_1094);
or U1551 (N_1551,N_1477,N_1263);
nand U1552 (N_1552,N_1048,N_1186);
or U1553 (N_1553,N_1152,N_1383);
and U1554 (N_1554,N_1315,N_1210);
or U1555 (N_1555,N_1065,N_1352);
xor U1556 (N_1556,N_1259,N_1207);
or U1557 (N_1557,N_1439,N_1469);
xor U1558 (N_1558,N_1411,N_1323);
and U1559 (N_1559,N_1197,N_1143);
nor U1560 (N_1560,N_1192,N_1322);
nor U1561 (N_1561,N_1184,N_1294);
nor U1562 (N_1562,N_1408,N_1296);
nor U1563 (N_1563,N_1397,N_1454);
or U1564 (N_1564,N_1461,N_1180);
nor U1565 (N_1565,N_1391,N_1426);
nor U1566 (N_1566,N_1088,N_1129);
nor U1567 (N_1567,N_1402,N_1485);
or U1568 (N_1568,N_1236,N_1182);
and U1569 (N_1569,N_1077,N_1301);
nor U1570 (N_1570,N_1009,N_1457);
or U1571 (N_1571,N_1166,N_1039);
xnor U1572 (N_1572,N_1139,N_1442);
nand U1573 (N_1573,N_1268,N_1211);
and U1574 (N_1574,N_1472,N_1367);
or U1575 (N_1575,N_1031,N_1092);
nand U1576 (N_1576,N_1475,N_1418);
nand U1577 (N_1577,N_1345,N_1307);
xor U1578 (N_1578,N_1064,N_1262);
nand U1579 (N_1579,N_1254,N_1229);
or U1580 (N_1580,N_1400,N_1347);
nor U1581 (N_1581,N_1251,N_1091);
and U1582 (N_1582,N_1054,N_1104);
nor U1583 (N_1583,N_1161,N_1410);
and U1584 (N_1584,N_1382,N_1429);
or U1585 (N_1585,N_1226,N_1154);
nor U1586 (N_1586,N_1327,N_1053);
nor U1587 (N_1587,N_1277,N_1200);
or U1588 (N_1588,N_1177,N_1082);
nand U1589 (N_1589,N_1495,N_1396);
or U1590 (N_1590,N_1431,N_1225);
or U1591 (N_1591,N_1486,N_1003);
nand U1592 (N_1592,N_1241,N_1325);
nand U1593 (N_1593,N_1160,N_1298);
nor U1594 (N_1594,N_1195,N_1044);
and U1595 (N_1595,N_1356,N_1278);
nand U1596 (N_1596,N_1436,N_1089);
and U1597 (N_1597,N_1204,N_1059);
nand U1598 (N_1598,N_1242,N_1107);
nor U1599 (N_1599,N_1409,N_1386);
nor U1600 (N_1600,N_1257,N_1416);
and U1601 (N_1601,N_1108,N_1417);
nand U1602 (N_1602,N_1272,N_1291);
nor U1603 (N_1603,N_1464,N_1448);
xnor U1604 (N_1604,N_1234,N_1337);
nand U1605 (N_1605,N_1453,N_1343);
and U1606 (N_1606,N_1374,N_1050);
and U1607 (N_1607,N_1141,N_1008);
and U1608 (N_1608,N_1187,N_1021);
and U1609 (N_1609,N_1024,N_1358);
nand U1610 (N_1610,N_1140,N_1199);
and U1611 (N_1611,N_1076,N_1179);
and U1612 (N_1612,N_1032,N_1474);
nor U1613 (N_1613,N_1338,N_1109);
and U1614 (N_1614,N_1218,N_1126);
xnor U1615 (N_1615,N_1171,N_1433);
or U1616 (N_1616,N_1040,N_1329);
xnor U1617 (N_1617,N_1102,N_1283);
or U1618 (N_1618,N_1355,N_1281);
or U1619 (N_1619,N_1299,N_1213);
or U1620 (N_1620,N_1062,N_1393);
nor U1621 (N_1621,N_1070,N_1145);
and U1622 (N_1622,N_1133,N_1312);
nand U1623 (N_1623,N_1098,N_1208);
nor U1624 (N_1624,N_1018,N_1381);
and U1625 (N_1625,N_1311,N_1144);
xor U1626 (N_1626,N_1101,N_1201);
nand U1627 (N_1627,N_1371,N_1363);
nor U1628 (N_1628,N_1191,N_1404);
xnor U1629 (N_1629,N_1282,N_1185);
nor U1630 (N_1630,N_1420,N_1249);
nand U1631 (N_1631,N_1205,N_1216);
nand U1632 (N_1632,N_1030,N_1119);
or U1633 (N_1633,N_1232,N_1206);
or U1634 (N_1634,N_1087,N_1438);
or U1635 (N_1635,N_1084,N_1389);
nor U1636 (N_1636,N_1470,N_1484);
nand U1637 (N_1637,N_1198,N_1314);
nand U1638 (N_1638,N_1388,N_1116);
nand U1639 (N_1639,N_1481,N_1375);
and U1640 (N_1640,N_1330,N_1111);
or U1641 (N_1641,N_1103,N_1467);
xnor U1642 (N_1642,N_1427,N_1190);
and U1643 (N_1643,N_1362,N_1487);
and U1644 (N_1644,N_1380,N_1112);
nor U1645 (N_1645,N_1328,N_1435);
and U1646 (N_1646,N_1392,N_1460);
or U1647 (N_1647,N_1449,N_1247);
nand U1648 (N_1648,N_1105,N_1006);
and U1649 (N_1649,N_1270,N_1316);
xnor U1650 (N_1650,N_1387,N_1369);
xor U1651 (N_1651,N_1022,N_1292);
xor U1652 (N_1652,N_1494,N_1060);
or U1653 (N_1653,N_1372,N_1224);
nand U1654 (N_1654,N_1203,N_1465);
nor U1655 (N_1655,N_1239,N_1214);
nor U1656 (N_1656,N_1033,N_1029);
and U1657 (N_1657,N_1181,N_1466);
nor U1658 (N_1658,N_1320,N_1339);
nand U1659 (N_1659,N_1342,N_1308);
or U1660 (N_1660,N_1360,N_1136);
xor U1661 (N_1661,N_1240,N_1243);
and U1662 (N_1662,N_1483,N_1384);
nor U1663 (N_1663,N_1271,N_1023);
and U1664 (N_1664,N_1447,N_1407);
xor U1665 (N_1665,N_1172,N_1149);
nand U1666 (N_1666,N_1354,N_1273);
xor U1667 (N_1667,N_1130,N_1349);
nor U1668 (N_1668,N_1385,N_1434);
nand U1669 (N_1669,N_1212,N_1255);
nand U1670 (N_1670,N_1376,N_1073);
and U1671 (N_1671,N_1010,N_1115);
xnor U1672 (N_1672,N_1132,N_1489);
nand U1673 (N_1673,N_1346,N_1097);
nor U1674 (N_1674,N_1415,N_1310);
nand U1675 (N_1675,N_1067,N_1252);
nor U1676 (N_1676,N_1289,N_1155);
and U1677 (N_1677,N_1364,N_1219);
and U1678 (N_1678,N_1028,N_1491);
and U1679 (N_1679,N_1012,N_1260);
and U1680 (N_1680,N_1335,N_1110);
and U1681 (N_1681,N_1178,N_1164);
nand U1682 (N_1682,N_1228,N_1279);
nand U1683 (N_1683,N_1222,N_1235);
nand U1684 (N_1684,N_1123,N_1223);
or U1685 (N_1685,N_1274,N_1450);
nor U1686 (N_1686,N_1319,N_1121);
nand U1687 (N_1687,N_1042,N_1090);
xor U1688 (N_1688,N_1419,N_1057);
or U1689 (N_1689,N_1074,N_1153);
xor U1690 (N_1690,N_1423,N_1245);
or U1691 (N_1691,N_1163,N_1432);
xor U1692 (N_1692,N_1081,N_1368);
xnor U1693 (N_1693,N_1366,N_1004);
or U1694 (N_1694,N_1276,N_1078);
and U1695 (N_1695,N_1348,N_1401);
or U1696 (N_1696,N_1394,N_1359);
or U1697 (N_1697,N_1159,N_1478);
or U1698 (N_1698,N_1071,N_1305);
or U1699 (N_1699,N_1290,N_1266);
nor U1700 (N_1700,N_1309,N_1002);
and U1701 (N_1701,N_1443,N_1174);
nand U1702 (N_1702,N_1317,N_1162);
and U1703 (N_1703,N_1011,N_1334);
and U1704 (N_1704,N_1170,N_1209);
or U1705 (N_1705,N_1096,N_1499);
nor U1706 (N_1706,N_1357,N_1488);
and U1707 (N_1707,N_1458,N_1095);
and U1708 (N_1708,N_1068,N_1131);
nand U1709 (N_1709,N_1321,N_1332);
nor U1710 (N_1710,N_1045,N_1001);
and U1711 (N_1711,N_1069,N_1168);
nor U1712 (N_1712,N_1038,N_1250);
nand U1713 (N_1713,N_1079,N_1007);
or U1714 (N_1714,N_1157,N_1473);
nand U1715 (N_1715,N_1471,N_1173);
or U1716 (N_1716,N_1425,N_1135);
and U1717 (N_1717,N_1015,N_1482);
or U1718 (N_1718,N_1399,N_1061);
xnor U1719 (N_1719,N_1446,N_1043);
nand U1720 (N_1720,N_1134,N_1269);
nand U1721 (N_1721,N_1137,N_1395);
or U1722 (N_1722,N_1014,N_1016);
nand U1723 (N_1723,N_1176,N_1318);
nor U1724 (N_1724,N_1128,N_1151);
nor U1725 (N_1725,N_1265,N_1303);
nor U1726 (N_1726,N_1286,N_1005);
and U1727 (N_1727,N_1085,N_1353);
nand U1728 (N_1728,N_1377,N_1253);
nor U1729 (N_1729,N_1293,N_1075);
nor U1730 (N_1730,N_1215,N_1196);
nor U1731 (N_1731,N_1026,N_1158);
or U1732 (N_1732,N_1233,N_1313);
nor U1733 (N_1733,N_1479,N_1217);
nand U1734 (N_1734,N_1297,N_1440);
and U1735 (N_1735,N_1455,N_1058);
xor U1736 (N_1736,N_1300,N_1124);
or U1737 (N_1737,N_1285,N_1169);
nor U1738 (N_1738,N_1147,N_1231);
or U1739 (N_1739,N_1175,N_1361);
nor U1740 (N_1740,N_1424,N_1496);
nor U1741 (N_1741,N_1189,N_1480);
or U1742 (N_1742,N_1066,N_1275);
nand U1743 (N_1743,N_1246,N_1441);
and U1744 (N_1744,N_1492,N_1100);
nand U1745 (N_1745,N_1452,N_1412);
and U1746 (N_1746,N_1264,N_1142);
and U1747 (N_1747,N_1046,N_1490);
nand U1748 (N_1748,N_1072,N_1324);
xnor U1749 (N_1749,N_1244,N_1114);
nand U1750 (N_1750,N_1426,N_1325);
or U1751 (N_1751,N_1436,N_1034);
nand U1752 (N_1752,N_1353,N_1076);
or U1753 (N_1753,N_1030,N_1102);
or U1754 (N_1754,N_1436,N_1238);
and U1755 (N_1755,N_1431,N_1220);
or U1756 (N_1756,N_1139,N_1176);
and U1757 (N_1757,N_1136,N_1316);
nor U1758 (N_1758,N_1051,N_1223);
nand U1759 (N_1759,N_1211,N_1235);
xor U1760 (N_1760,N_1366,N_1050);
nor U1761 (N_1761,N_1447,N_1300);
nor U1762 (N_1762,N_1296,N_1291);
nand U1763 (N_1763,N_1000,N_1274);
or U1764 (N_1764,N_1373,N_1332);
and U1765 (N_1765,N_1010,N_1042);
and U1766 (N_1766,N_1382,N_1329);
xor U1767 (N_1767,N_1214,N_1412);
nand U1768 (N_1768,N_1310,N_1154);
xnor U1769 (N_1769,N_1230,N_1150);
nand U1770 (N_1770,N_1320,N_1326);
or U1771 (N_1771,N_1021,N_1357);
or U1772 (N_1772,N_1483,N_1230);
and U1773 (N_1773,N_1480,N_1361);
nand U1774 (N_1774,N_1451,N_1283);
nand U1775 (N_1775,N_1392,N_1271);
nand U1776 (N_1776,N_1060,N_1241);
nand U1777 (N_1777,N_1453,N_1299);
xor U1778 (N_1778,N_1337,N_1348);
nand U1779 (N_1779,N_1303,N_1393);
and U1780 (N_1780,N_1330,N_1312);
and U1781 (N_1781,N_1413,N_1082);
nor U1782 (N_1782,N_1077,N_1368);
nand U1783 (N_1783,N_1046,N_1280);
or U1784 (N_1784,N_1423,N_1151);
and U1785 (N_1785,N_1174,N_1259);
nand U1786 (N_1786,N_1056,N_1370);
or U1787 (N_1787,N_1450,N_1428);
nor U1788 (N_1788,N_1233,N_1351);
or U1789 (N_1789,N_1456,N_1029);
and U1790 (N_1790,N_1305,N_1486);
nor U1791 (N_1791,N_1002,N_1267);
and U1792 (N_1792,N_1299,N_1232);
and U1793 (N_1793,N_1476,N_1029);
or U1794 (N_1794,N_1021,N_1274);
nand U1795 (N_1795,N_1178,N_1226);
nor U1796 (N_1796,N_1005,N_1059);
nor U1797 (N_1797,N_1110,N_1395);
nor U1798 (N_1798,N_1313,N_1152);
and U1799 (N_1799,N_1086,N_1232);
or U1800 (N_1800,N_1115,N_1402);
or U1801 (N_1801,N_1008,N_1374);
nand U1802 (N_1802,N_1178,N_1253);
or U1803 (N_1803,N_1245,N_1429);
and U1804 (N_1804,N_1092,N_1055);
nand U1805 (N_1805,N_1448,N_1364);
nand U1806 (N_1806,N_1099,N_1475);
and U1807 (N_1807,N_1371,N_1277);
nor U1808 (N_1808,N_1052,N_1159);
nor U1809 (N_1809,N_1334,N_1305);
nand U1810 (N_1810,N_1184,N_1369);
nand U1811 (N_1811,N_1101,N_1073);
xor U1812 (N_1812,N_1348,N_1072);
xor U1813 (N_1813,N_1113,N_1335);
and U1814 (N_1814,N_1132,N_1078);
or U1815 (N_1815,N_1392,N_1134);
or U1816 (N_1816,N_1124,N_1032);
nor U1817 (N_1817,N_1246,N_1409);
xor U1818 (N_1818,N_1133,N_1107);
and U1819 (N_1819,N_1189,N_1370);
or U1820 (N_1820,N_1073,N_1343);
xor U1821 (N_1821,N_1314,N_1182);
nor U1822 (N_1822,N_1495,N_1187);
and U1823 (N_1823,N_1258,N_1438);
and U1824 (N_1824,N_1355,N_1250);
or U1825 (N_1825,N_1243,N_1211);
or U1826 (N_1826,N_1278,N_1170);
and U1827 (N_1827,N_1020,N_1030);
nand U1828 (N_1828,N_1119,N_1253);
and U1829 (N_1829,N_1098,N_1162);
or U1830 (N_1830,N_1036,N_1059);
and U1831 (N_1831,N_1271,N_1202);
and U1832 (N_1832,N_1425,N_1200);
or U1833 (N_1833,N_1282,N_1409);
nor U1834 (N_1834,N_1452,N_1486);
and U1835 (N_1835,N_1015,N_1021);
and U1836 (N_1836,N_1031,N_1483);
nor U1837 (N_1837,N_1122,N_1013);
nand U1838 (N_1838,N_1393,N_1014);
nand U1839 (N_1839,N_1069,N_1082);
nand U1840 (N_1840,N_1172,N_1483);
xor U1841 (N_1841,N_1225,N_1337);
nand U1842 (N_1842,N_1248,N_1152);
and U1843 (N_1843,N_1404,N_1067);
nand U1844 (N_1844,N_1492,N_1238);
nor U1845 (N_1845,N_1348,N_1015);
nand U1846 (N_1846,N_1293,N_1001);
and U1847 (N_1847,N_1068,N_1241);
xnor U1848 (N_1848,N_1167,N_1497);
nand U1849 (N_1849,N_1268,N_1071);
or U1850 (N_1850,N_1204,N_1276);
xnor U1851 (N_1851,N_1488,N_1208);
nor U1852 (N_1852,N_1376,N_1259);
nand U1853 (N_1853,N_1424,N_1380);
xor U1854 (N_1854,N_1413,N_1330);
or U1855 (N_1855,N_1380,N_1353);
nor U1856 (N_1856,N_1433,N_1439);
nand U1857 (N_1857,N_1083,N_1100);
nand U1858 (N_1858,N_1486,N_1436);
nand U1859 (N_1859,N_1455,N_1074);
xor U1860 (N_1860,N_1460,N_1091);
xnor U1861 (N_1861,N_1039,N_1016);
nor U1862 (N_1862,N_1253,N_1248);
and U1863 (N_1863,N_1281,N_1172);
nor U1864 (N_1864,N_1269,N_1045);
or U1865 (N_1865,N_1272,N_1496);
xor U1866 (N_1866,N_1410,N_1154);
xnor U1867 (N_1867,N_1257,N_1490);
or U1868 (N_1868,N_1030,N_1417);
and U1869 (N_1869,N_1014,N_1254);
nor U1870 (N_1870,N_1342,N_1388);
and U1871 (N_1871,N_1081,N_1006);
or U1872 (N_1872,N_1177,N_1194);
or U1873 (N_1873,N_1213,N_1016);
or U1874 (N_1874,N_1275,N_1426);
and U1875 (N_1875,N_1113,N_1247);
nor U1876 (N_1876,N_1244,N_1352);
and U1877 (N_1877,N_1468,N_1282);
nand U1878 (N_1878,N_1122,N_1329);
and U1879 (N_1879,N_1254,N_1032);
nand U1880 (N_1880,N_1297,N_1420);
xnor U1881 (N_1881,N_1110,N_1006);
and U1882 (N_1882,N_1173,N_1193);
nand U1883 (N_1883,N_1469,N_1130);
nor U1884 (N_1884,N_1141,N_1074);
and U1885 (N_1885,N_1240,N_1485);
or U1886 (N_1886,N_1294,N_1169);
or U1887 (N_1887,N_1440,N_1104);
nand U1888 (N_1888,N_1139,N_1357);
or U1889 (N_1889,N_1057,N_1317);
nor U1890 (N_1890,N_1380,N_1469);
nor U1891 (N_1891,N_1294,N_1010);
or U1892 (N_1892,N_1164,N_1485);
xnor U1893 (N_1893,N_1324,N_1289);
nand U1894 (N_1894,N_1171,N_1029);
nor U1895 (N_1895,N_1423,N_1059);
nor U1896 (N_1896,N_1091,N_1173);
and U1897 (N_1897,N_1201,N_1273);
and U1898 (N_1898,N_1315,N_1291);
xor U1899 (N_1899,N_1393,N_1234);
or U1900 (N_1900,N_1440,N_1352);
xor U1901 (N_1901,N_1151,N_1485);
nand U1902 (N_1902,N_1294,N_1098);
and U1903 (N_1903,N_1215,N_1293);
or U1904 (N_1904,N_1121,N_1084);
nand U1905 (N_1905,N_1308,N_1477);
or U1906 (N_1906,N_1402,N_1112);
nor U1907 (N_1907,N_1096,N_1135);
or U1908 (N_1908,N_1429,N_1185);
and U1909 (N_1909,N_1116,N_1180);
nand U1910 (N_1910,N_1360,N_1447);
xnor U1911 (N_1911,N_1064,N_1285);
nand U1912 (N_1912,N_1131,N_1002);
nand U1913 (N_1913,N_1048,N_1197);
or U1914 (N_1914,N_1325,N_1359);
or U1915 (N_1915,N_1102,N_1013);
or U1916 (N_1916,N_1165,N_1173);
and U1917 (N_1917,N_1177,N_1340);
xor U1918 (N_1918,N_1453,N_1177);
nor U1919 (N_1919,N_1197,N_1324);
xor U1920 (N_1920,N_1254,N_1242);
or U1921 (N_1921,N_1104,N_1191);
nand U1922 (N_1922,N_1151,N_1161);
xnor U1923 (N_1923,N_1120,N_1022);
nor U1924 (N_1924,N_1210,N_1132);
nor U1925 (N_1925,N_1319,N_1173);
and U1926 (N_1926,N_1091,N_1379);
nor U1927 (N_1927,N_1477,N_1239);
xor U1928 (N_1928,N_1009,N_1053);
nor U1929 (N_1929,N_1058,N_1167);
nor U1930 (N_1930,N_1155,N_1041);
or U1931 (N_1931,N_1163,N_1433);
nor U1932 (N_1932,N_1438,N_1193);
or U1933 (N_1933,N_1462,N_1457);
and U1934 (N_1934,N_1174,N_1031);
nand U1935 (N_1935,N_1045,N_1334);
nand U1936 (N_1936,N_1019,N_1467);
and U1937 (N_1937,N_1476,N_1117);
nor U1938 (N_1938,N_1140,N_1301);
and U1939 (N_1939,N_1063,N_1313);
xor U1940 (N_1940,N_1243,N_1414);
nor U1941 (N_1941,N_1227,N_1442);
nor U1942 (N_1942,N_1293,N_1000);
nor U1943 (N_1943,N_1350,N_1272);
nor U1944 (N_1944,N_1323,N_1097);
nor U1945 (N_1945,N_1096,N_1000);
or U1946 (N_1946,N_1109,N_1427);
nor U1947 (N_1947,N_1294,N_1250);
and U1948 (N_1948,N_1309,N_1191);
nand U1949 (N_1949,N_1381,N_1021);
nor U1950 (N_1950,N_1268,N_1257);
or U1951 (N_1951,N_1283,N_1335);
xnor U1952 (N_1952,N_1457,N_1325);
nand U1953 (N_1953,N_1092,N_1386);
xnor U1954 (N_1954,N_1155,N_1388);
and U1955 (N_1955,N_1259,N_1477);
nor U1956 (N_1956,N_1233,N_1201);
nor U1957 (N_1957,N_1202,N_1171);
nand U1958 (N_1958,N_1344,N_1342);
or U1959 (N_1959,N_1486,N_1156);
nand U1960 (N_1960,N_1153,N_1310);
nor U1961 (N_1961,N_1233,N_1038);
and U1962 (N_1962,N_1447,N_1384);
nand U1963 (N_1963,N_1448,N_1288);
or U1964 (N_1964,N_1292,N_1442);
and U1965 (N_1965,N_1177,N_1307);
nand U1966 (N_1966,N_1235,N_1282);
and U1967 (N_1967,N_1088,N_1038);
nand U1968 (N_1968,N_1160,N_1422);
nor U1969 (N_1969,N_1085,N_1297);
and U1970 (N_1970,N_1180,N_1217);
nand U1971 (N_1971,N_1237,N_1402);
or U1972 (N_1972,N_1031,N_1207);
xor U1973 (N_1973,N_1402,N_1139);
nor U1974 (N_1974,N_1498,N_1322);
xor U1975 (N_1975,N_1248,N_1057);
nand U1976 (N_1976,N_1333,N_1021);
nor U1977 (N_1977,N_1203,N_1223);
and U1978 (N_1978,N_1279,N_1039);
xor U1979 (N_1979,N_1121,N_1001);
or U1980 (N_1980,N_1434,N_1160);
xor U1981 (N_1981,N_1214,N_1358);
xor U1982 (N_1982,N_1469,N_1078);
nor U1983 (N_1983,N_1405,N_1119);
nor U1984 (N_1984,N_1126,N_1241);
nor U1985 (N_1985,N_1011,N_1315);
xor U1986 (N_1986,N_1370,N_1197);
nor U1987 (N_1987,N_1492,N_1065);
or U1988 (N_1988,N_1141,N_1090);
or U1989 (N_1989,N_1260,N_1288);
nand U1990 (N_1990,N_1007,N_1278);
nand U1991 (N_1991,N_1084,N_1263);
nand U1992 (N_1992,N_1054,N_1035);
xnor U1993 (N_1993,N_1172,N_1433);
xnor U1994 (N_1994,N_1258,N_1177);
and U1995 (N_1995,N_1464,N_1499);
nor U1996 (N_1996,N_1151,N_1056);
nand U1997 (N_1997,N_1311,N_1027);
and U1998 (N_1998,N_1219,N_1321);
nor U1999 (N_1999,N_1195,N_1213);
and U2000 (N_2000,N_1580,N_1661);
nand U2001 (N_2001,N_1507,N_1584);
or U2002 (N_2002,N_1505,N_1648);
and U2003 (N_2003,N_1998,N_1705);
nor U2004 (N_2004,N_1793,N_1950);
nand U2005 (N_2005,N_1889,N_1916);
or U2006 (N_2006,N_1698,N_1955);
nor U2007 (N_2007,N_1603,N_1904);
and U2008 (N_2008,N_1837,N_1772);
nand U2009 (N_2009,N_1780,N_1754);
or U2010 (N_2010,N_1631,N_1579);
nand U2011 (N_2011,N_1724,N_1795);
nor U2012 (N_2012,N_1746,N_1536);
or U2013 (N_2013,N_1851,N_1583);
or U2014 (N_2014,N_1991,N_1739);
and U2015 (N_2015,N_1903,N_1737);
and U2016 (N_2016,N_1758,N_1978);
nand U2017 (N_2017,N_1573,N_1764);
and U2018 (N_2018,N_1800,N_1864);
or U2019 (N_2019,N_1568,N_1627);
nand U2020 (N_2020,N_1894,N_1517);
nand U2021 (N_2021,N_1594,N_1918);
and U2022 (N_2022,N_1662,N_1528);
and U2023 (N_2023,N_1628,N_1763);
and U2024 (N_2024,N_1714,N_1860);
xnor U2025 (N_2025,N_1741,N_1686);
nand U2026 (N_2026,N_1944,N_1613);
and U2027 (N_2027,N_1824,N_1880);
and U2028 (N_2028,N_1823,N_1570);
nor U2029 (N_2029,N_1975,N_1666);
or U2030 (N_2030,N_1711,N_1592);
nand U2031 (N_2031,N_1940,N_1876);
nor U2032 (N_2032,N_1817,N_1827);
and U2033 (N_2033,N_1512,N_1738);
nand U2034 (N_2034,N_1921,N_1912);
nand U2035 (N_2035,N_1706,N_1989);
or U2036 (N_2036,N_1777,N_1830);
nor U2037 (N_2037,N_1722,N_1601);
nand U2038 (N_2038,N_1976,N_1548);
nand U2039 (N_2039,N_1890,N_1668);
and U2040 (N_2040,N_1923,N_1832);
and U2041 (N_2041,N_1759,N_1813);
nor U2042 (N_2042,N_1665,N_1966);
nor U2043 (N_2043,N_1563,N_1770);
or U2044 (N_2044,N_1617,N_1854);
and U2045 (N_2045,N_1957,N_1997);
and U2046 (N_2046,N_1969,N_1858);
and U2047 (N_2047,N_1914,N_1620);
nor U2048 (N_2048,N_1659,N_1637);
and U2049 (N_2049,N_1942,N_1586);
nor U2050 (N_2050,N_1525,N_1762);
nand U2051 (N_2051,N_1929,N_1947);
nand U2052 (N_2052,N_1681,N_1547);
and U2053 (N_2053,N_1938,N_1778);
or U2054 (N_2054,N_1862,N_1751);
nor U2055 (N_2055,N_1590,N_1588);
and U2056 (N_2056,N_1514,N_1671);
nor U2057 (N_2057,N_1885,N_1905);
or U2058 (N_2058,N_1895,N_1605);
nand U2059 (N_2059,N_1878,N_1844);
nand U2060 (N_2060,N_1527,N_1526);
xnor U2061 (N_2061,N_1719,N_1756);
or U2062 (N_2062,N_1682,N_1883);
or U2063 (N_2063,N_1587,N_1589);
nor U2064 (N_2064,N_1853,N_1888);
or U2065 (N_2065,N_1638,N_1755);
and U2066 (N_2066,N_1608,N_1930);
nand U2067 (N_2067,N_1546,N_1537);
and U2068 (N_2068,N_1875,N_1656);
nor U2069 (N_2069,N_1731,N_1810);
nand U2070 (N_2070,N_1531,N_1806);
nand U2071 (N_2071,N_1664,N_1700);
xnor U2072 (N_2072,N_1977,N_1776);
or U2073 (N_2073,N_1708,N_1909);
nand U2074 (N_2074,N_1652,N_1769);
xor U2075 (N_2075,N_1692,N_1654);
or U2076 (N_2076,N_1999,N_1882);
xor U2077 (N_2077,N_1796,N_1683);
and U2078 (N_2078,N_1863,N_1971);
nand U2079 (N_2079,N_1768,N_1560);
and U2080 (N_2080,N_1632,N_1848);
or U2081 (N_2081,N_1612,N_1629);
or U2082 (N_2082,N_1650,N_1967);
nor U2083 (N_2083,N_1825,N_1742);
nor U2084 (N_2084,N_1616,N_1834);
and U2085 (N_2085,N_1840,N_1680);
xor U2086 (N_2086,N_1753,N_1729);
nand U2087 (N_2087,N_1639,N_1716);
or U2088 (N_2088,N_1979,N_1922);
and U2089 (N_2089,N_1633,N_1676);
or U2090 (N_2090,N_1933,N_1907);
nand U2091 (N_2091,N_1713,N_1785);
or U2092 (N_2092,N_1812,N_1747);
and U2093 (N_2093,N_1710,N_1784);
nand U2094 (N_2094,N_1841,N_1609);
or U2095 (N_2095,N_1718,N_1958);
and U2096 (N_2096,N_1582,N_1630);
xnor U2097 (N_2097,N_1732,N_1712);
and U2098 (N_2098,N_1773,N_1543);
or U2099 (N_2099,N_1757,N_1550);
nand U2100 (N_2100,N_1625,N_1677);
nor U2101 (N_2101,N_1591,N_1624);
nor U2102 (N_2102,N_1985,N_1786);
or U2103 (N_2103,N_1911,N_1760);
or U2104 (N_2104,N_1618,N_1994);
xor U2105 (N_2105,N_1565,N_1927);
and U2106 (N_2106,N_1635,N_1670);
and U2107 (N_2107,N_1807,N_1926);
nor U2108 (N_2108,N_1881,N_1693);
or U2109 (N_2109,N_1646,N_1736);
nand U2110 (N_2110,N_1564,N_1816);
nor U2111 (N_2111,N_1685,N_1687);
and U2112 (N_2112,N_1541,N_1782);
or U2113 (N_2113,N_1576,N_1986);
nor U2114 (N_2114,N_1524,N_1554);
or U2115 (N_2115,N_1581,N_1574);
nor U2116 (N_2116,N_1811,N_1996);
and U2117 (N_2117,N_1622,N_1644);
nand U2118 (N_2118,N_1963,N_1794);
and U2119 (N_2119,N_1752,N_1897);
and U2120 (N_2120,N_1669,N_1917);
or U2121 (N_2121,N_1879,N_1538);
and U2122 (N_2122,N_1822,N_1783);
and U2123 (N_2123,N_1750,N_1697);
and U2124 (N_2124,N_1691,N_1870);
and U2125 (N_2125,N_1804,N_1509);
xnor U2126 (N_2126,N_1765,N_1694);
xor U2127 (N_2127,N_1688,N_1936);
or U2128 (N_2128,N_1913,N_1906);
nand U2129 (N_2129,N_1571,N_1634);
xor U2130 (N_2130,N_1707,N_1699);
nor U2131 (N_2131,N_1809,N_1835);
or U2132 (N_2132,N_1521,N_1552);
or U2133 (N_2133,N_1826,N_1900);
or U2134 (N_2134,N_1566,N_1740);
or U2135 (N_2135,N_1856,N_1798);
and U2136 (N_2136,N_1529,N_1720);
and U2137 (N_2137,N_1744,N_1596);
nand U2138 (N_2138,N_1690,N_1910);
and U2139 (N_2139,N_1645,N_1867);
or U2140 (N_2140,N_1855,N_1619);
and U2141 (N_2141,N_1802,N_1803);
and U2142 (N_2142,N_1558,N_1761);
and U2143 (N_2143,N_1674,N_1501);
nand U2144 (N_2144,N_1775,N_1701);
xor U2145 (N_2145,N_1519,N_1653);
or U2146 (N_2146,N_1684,N_1974);
and U2147 (N_2147,N_1962,N_1606);
nand U2148 (N_2148,N_1919,N_1831);
nor U2149 (N_2149,N_1988,N_1726);
and U2150 (N_2150,N_1607,N_1611);
or U2151 (N_2151,N_1873,N_1987);
or U2152 (N_2152,N_1925,N_1839);
nor U2153 (N_2153,N_1504,N_1932);
xor U2154 (N_2154,N_1503,N_1931);
nand U2155 (N_2155,N_1555,N_1748);
and U2156 (N_2156,N_1673,N_1551);
or U2157 (N_2157,N_1728,N_1949);
nor U2158 (N_2158,N_1604,N_1893);
nand U2159 (N_2159,N_1792,N_1920);
or U2160 (N_2160,N_1600,N_1544);
or U2161 (N_2161,N_1790,N_1959);
nand U2162 (N_2162,N_1679,N_1928);
xnor U2163 (N_2163,N_1805,N_1866);
nor U2164 (N_2164,N_1557,N_1845);
or U2165 (N_2165,N_1973,N_1672);
xor U2166 (N_2166,N_1717,N_1857);
and U2167 (N_2167,N_1621,N_1941);
or U2168 (N_2168,N_1956,N_1833);
nand U2169 (N_2169,N_1945,N_1970);
nor U2170 (N_2170,N_1992,N_1801);
and U2171 (N_2171,N_1774,N_1508);
nand U2172 (N_2172,N_1651,N_1561);
and U2173 (N_2173,N_1636,N_1715);
or U2174 (N_2174,N_1852,N_1982);
and U2175 (N_2175,N_1943,N_1952);
nand U2176 (N_2176,N_1791,N_1868);
and U2177 (N_2177,N_1532,N_1559);
or U2178 (N_2178,N_1721,N_1808);
nand U2179 (N_2179,N_1815,N_1735);
and U2180 (N_2180,N_1766,N_1539);
nor U2181 (N_2181,N_1908,N_1533);
nor U2182 (N_2182,N_1954,N_1953);
nand U2183 (N_2183,N_1585,N_1595);
xor U2184 (N_2184,N_1695,N_1540);
nand U2185 (N_2185,N_1983,N_1877);
and U2186 (N_2186,N_1829,N_1658);
and U2187 (N_2187,N_1647,N_1614);
xor U2188 (N_2188,N_1667,N_1597);
nor U2189 (N_2189,N_1599,N_1643);
and U2190 (N_2190,N_1884,N_1678);
or U2191 (N_2191,N_1787,N_1641);
nand U2192 (N_2192,N_1838,N_1655);
nand U2193 (N_2193,N_1623,N_1513);
nand U2194 (N_2194,N_1924,N_1502);
nand U2195 (N_2195,N_1556,N_1578);
nand U2196 (N_2196,N_1534,N_1523);
and U2197 (N_2197,N_1510,N_1569);
nor U2198 (N_2198,N_1704,N_1610);
xnor U2199 (N_2199,N_1788,N_1993);
xnor U2200 (N_2200,N_1887,N_1902);
nor U2201 (N_2201,N_1771,N_1553);
xor U2202 (N_2202,N_1730,N_1500);
nand U2203 (N_2203,N_1935,N_1663);
nand U2204 (N_2204,N_1951,N_1934);
nor U2205 (N_2205,N_1821,N_1828);
or U2206 (N_2206,N_1859,N_1734);
nor U2207 (N_2207,N_1847,N_1886);
or U2208 (N_2208,N_1915,N_1995);
nor U2209 (N_2209,N_1948,N_1520);
or U2210 (N_2210,N_1745,N_1572);
or U2211 (N_2211,N_1549,N_1577);
xor U2212 (N_2212,N_1602,N_1615);
nor U2213 (N_2213,N_1980,N_1965);
nand U2214 (N_2214,N_1836,N_1842);
nand U2215 (N_2215,N_1640,N_1749);
nand U2216 (N_2216,N_1872,N_1522);
or U2217 (N_2217,N_1545,N_1797);
and U2218 (N_2218,N_1767,N_1598);
nand U2219 (N_2219,N_1515,N_1937);
and U2220 (N_2220,N_1725,N_1575);
and U2221 (N_2221,N_1593,N_1898);
nor U2222 (N_2222,N_1506,N_1530);
xor U2223 (N_2223,N_1901,N_1518);
xnor U2224 (N_2224,N_1946,N_1703);
nor U2225 (N_2225,N_1723,N_1727);
and U2226 (N_2226,N_1843,N_1891);
nor U2227 (N_2227,N_1849,N_1516);
or U2228 (N_2228,N_1789,N_1850);
nor U2229 (N_2229,N_1871,N_1675);
and U2230 (N_2230,N_1865,N_1899);
nand U2231 (N_2231,N_1567,N_1626);
xor U2232 (N_2232,N_1660,N_1961);
or U2233 (N_2233,N_1799,N_1984);
nand U2234 (N_2234,N_1535,N_1657);
and U2235 (N_2235,N_1892,N_1896);
nand U2236 (N_2236,N_1733,N_1696);
or U2237 (N_2237,N_1562,N_1781);
or U2238 (N_2238,N_1820,N_1702);
nor U2239 (N_2239,N_1874,N_1846);
nand U2240 (N_2240,N_1968,N_1649);
and U2241 (N_2241,N_1960,N_1981);
xor U2242 (N_2242,N_1542,N_1861);
and U2243 (N_2243,N_1779,N_1689);
nor U2244 (N_2244,N_1972,N_1814);
xor U2245 (N_2245,N_1964,N_1642);
xnor U2246 (N_2246,N_1869,N_1743);
or U2247 (N_2247,N_1511,N_1709);
nor U2248 (N_2248,N_1819,N_1818);
nand U2249 (N_2249,N_1939,N_1990);
nand U2250 (N_2250,N_1536,N_1997);
or U2251 (N_2251,N_1554,N_1704);
nor U2252 (N_2252,N_1573,N_1944);
or U2253 (N_2253,N_1881,N_1650);
nand U2254 (N_2254,N_1810,N_1866);
and U2255 (N_2255,N_1946,N_1867);
nand U2256 (N_2256,N_1999,N_1895);
or U2257 (N_2257,N_1817,N_1692);
or U2258 (N_2258,N_1974,N_1614);
and U2259 (N_2259,N_1709,N_1628);
and U2260 (N_2260,N_1726,N_1820);
or U2261 (N_2261,N_1964,N_1916);
nand U2262 (N_2262,N_1510,N_1988);
nand U2263 (N_2263,N_1550,N_1766);
or U2264 (N_2264,N_1957,N_1612);
and U2265 (N_2265,N_1981,N_1514);
or U2266 (N_2266,N_1917,N_1716);
xnor U2267 (N_2267,N_1562,N_1980);
or U2268 (N_2268,N_1918,N_1844);
or U2269 (N_2269,N_1531,N_1601);
or U2270 (N_2270,N_1776,N_1832);
nor U2271 (N_2271,N_1573,N_1794);
and U2272 (N_2272,N_1705,N_1679);
or U2273 (N_2273,N_1504,N_1920);
nand U2274 (N_2274,N_1599,N_1764);
or U2275 (N_2275,N_1895,N_1545);
nand U2276 (N_2276,N_1777,N_1980);
nand U2277 (N_2277,N_1762,N_1519);
nor U2278 (N_2278,N_1835,N_1938);
or U2279 (N_2279,N_1838,N_1531);
xor U2280 (N_2280,N_1618,N_1731);
or U2281 (N_2281,N_1776,N_1981);
or U2282 (N_2282,N_1673,N_1883);
nand U2283 (N_2283,N_1605,N_1939);
nand U2284 (N_2284,N_1755,N_1529);
or U2285 (N_2285,N_1533,N_1749);
or U2286 (N_2286,N_1944,N_1777);
nor U2287 (N_2287,N_1573,N_1669);
and U2288 (N_2288,N_1794,N_1846);
xnor U2289 (N_2289,N_1799,N_1857);
nor U2290 (N_2290,N_1560,N_1590);
nor U2291 (N_2291,N_1819,N_1589);
nor U2292 (N_2292,N_1713,N_1929);
xor U2293 (N_2293,N_1660,N_1851);
nand U2294 (N_2294,N_1887,N_1578);
or U2295 (N_2295,N_1549,N_1656);
and U2296 (N_2296,N_1811,N_1642);
or U2297 (N_2297,N_1740,N_1771);
nand U2298 (N_2298,N_1770,N_1829);
nor U2299 (N_2299,N_1500,N_1687);
and U2300 (N_2300,N_1619,N_1898);
and U2301 (N_2301,N_1747,N_1697);
and U2302 (N_2302,N_1710,N_1720);
nor U2303 (N_2303,N_1778,N_1779);
nor U2304 (N_2304,N_1778,N_1576);
xnor U2305 (N_2305,N_1677,N_1809);
nor U2306 (N_2306,N_1694,N_1522);
nor U2307 (N_2307,N_1526,N_1659);
nor U2308 (N_2308,N_1744,N_1707);
and U2309 (N_2309,N_1831,N_1583);
or U2310 (N_2310,N_1552,N_1602);
xnor U2311 (N_2311,N_1922,N_1897);
nand U2312 (N_2312,N_1704,N_1782);
and U2313 (N_2313,N_1951,N_1851);
and U2314 (N_2314,N_1608,N_1886);
and U2315 (N_2315,N_1753,N_1631);
and U2316 (N_2316,N_1663,N_1996);
and U2317 (N_2317,N_1690,N_1913);
nand U2318 (N_2318,N_1646,N_1971);
or U2319 (N_2319,N_1844,N_1600);
or U2320 (N_2320,N_1734,N_1714);
or U2321 (N_2321,N_1662,N_1530);
nand U2322 (N_2322,N_1751,N_1554);
nor U2323 (N_2323,N_1591,N_1808);
nand U2324 (N_2324,N_1703,N_1994);
nor U2325 (N_2325,N_1653,N_1727);
or U2326 (N_2326,N_1715,N_1956);
nand U2327 (N_2327,N_1706,N_1897);
and U2328 (N_2328,N_1604,N_1563);
or U2329 (N_2329,N_1914,N_1777);
or U2330 (N_2330,N_1694,N_1552);
or U2331 (N_2331,N_1873,N_1523);
nor U2332 (N_2332,N_1967,N_1973);
and U2333 (N_2333,N_1726,N_1662);
nand U2334 (N_2334,N_1986,N_1518);
nand U2335 (N_2335,N_1976,N_1641);
and U2336 (N_2336,N_1817,N_1717);
xnor U2337 (N_2337,N_1576,N_1506);
nand U2338 (N_2338,N_1890,N_1726);
nand U2339 (N_2339,N_1909,N_1896);
or U2340 (N_2340,N_1843,N_1540);
or U2341 (N_2341,N_1917,N_1553);
or U2342 (N_2342,N_1653,N_1601);
nor U2343 (N_2343,N_1971,N_1785);
xor U2344 (N_2344,N_1721,N_1907);
nand U2345 (N_2345,N_1628,N_1764);
or U2346 (N_2346,N_1572,N_1907);
nand U2347 (N_2347,N_1905,N_1632);
and U2348 (N_2348,N_1591,N_1887);
nor U2349 (N_2349,N_1710,N_1554);
or U2350 (N_2350,N_1987,N_1632);
nand U2351 (N_2351,N_1906,N_1504);
and U2352 (N_2352,N_1549,N_1757);
and U2353 (N_2353,N_1649,N_1643);
or U2354 (N_2354,N_1797,N_1809);
nor U2355 (N_2355,N_1989,N_1590);
nand U2356 (N_2356,N_1958,N_1962);
and U2357 (N_2357,N_1909,N_1971);
xnor U2358 (N_2358,N_1533,N_1876);
xnor U2359 (N_2359,N_1558,N_1896);
nor U2360 (N_2360,N_1553,N_1624);
nor U2361 (N_2361,N_1729,N_1927);
or U2362 (N_2362,N_1784,N_1863);
and U2363 (N_2363,N_1907,N_1765);
and U2364 (N_2364,N_1586,N_1763);
nor U2365 (N_2365,N_1918,N_1756);
and U2366 (N_2366,N_1964,N_1996);
or U2367 (N_2367,N_1538,N_1665);
or U2368 (N_2368,N_1526,N_1825);
nand U2369 (N_2369,N_1912,N_1753);
nand U2370 (N_2370,N_1668,N_1907);
nor U2371 (N_2371,N_1913,N_1702);
and U2372 (N_2372,N_1830,N_1553);
nand U2373 (N_2373,N_1540,N_1567);
nand U2374 (N_2374,N_1518,N_1948);
xnor U2375 (N_2375,N_1947,N_1525);
xnor U2376 (N_2376,N_1676,N_1923);
nor U2377 (N_2377,N_1779,N_1734);
nor U2378 (N_2378,N_1516,N_1760);
nor U2379 (N_2379,N_1849,N_1644);
nor U2380 (N_2380,N_1798,N_1672);
nand U2381 (N_2381,N_1557,N_1986);
and U2382 (N_2382,N_1596,N_1754);
nand U2383 (N_2383,N_1969,N_1632);
nor U2384 (N_2384,N_1524,N_1857);
nor U2385 (N_2385,N_1554,N_1581);
and U2386 (N_2386,N_1552,N_1943);
nor U2387 (N_2387,N_1981,N_1868);
or U2388 (N_2388,N_1818,N_1640);
nand U2389 (N_2389,N_1674,N_1520);
or U2390 (N_2390,N_1999,N_1564);
or U2391 (N_2391,N_1683,N_1658);
and U2392 (N_2392,N_1959,N_1672);
and U2393 (N_2393,N_1521,N_1717);
nand U2394 (N_2394,N_1539,N_1631);
xor U2395 (N_2395,N_1528,N_1977);
xnor U2396 (N_2396,N_1543,N_1554);
or U2397 (N_2397,N_1558,N_1677);
nor U2398 (N_2398,N_1981,N_1978);
nand U2399 (N_2399,N_1640,N_1888);
xor U2400 (N_2400,N_1865,N_1867);
or U2401 (N_2401,N_1613,N_1775);
nand U2402 (N_2402,N_1845,N_1953);
nor U2403 (N_2403,N_1942,N_1871);
and U2404 (N_2404,N_1702,N_1677);
or U2405 (N_2405,N_1563,N_1902);
xnor U2406 (N_2406,N_1643,N_1589);
nand U2407 (N_2407,N_1768,N_1767);
and U2408 (N_2408,N_1724,N_1978);
and U2409 (N_2409,N_1757,N_1614);
or U2410 (N_2410,N_1588,N_1664);
nor U2411 (N_2411,N_1615,N_1593);
or U2412 (N_2412,N_1928,N_1501);
xor U2413 (N_2413,N_1585,N_1946);
xor U2414 (N_2414,N_1834,N_1635);
nand U2415 (N_2415,N_1776,N_1796);
or U2416 (N_2416,N_1904,N_1889);
and U2417 (N_2417,N_1938,N_1826);
or U2418 (N_2418,N_1665,N_1883);
or U2419 (N_2419,N_1597,N_1655);
nor U2420 (N_2420,N_1750,N_1560);
or U2421 (N_2421,N_1864,N_1953);
nand U2422 (N_2422,N_1957,N_1675);
nand U2423 (N_2423,N_1691,N_1887);
nor U2424 (N_2424,N_1675,N_1714);
nor U2425 (N_2425,N_1545,N_1510);
nand U2426 (N_2426,N_1856,N_1824);
nor U2427 (N_2427,N_1796,N_1711);
nand U2428 (N_2428,N_1732,N_1811);
and U2429 (N_2429,N_1507,N_1847);
nor U2430 (N_2430,N_1732,N_1503);
or U2431 (N_2431,N_1899,N_1575);
nor U2432 (N_2432,N_1641,N_1511);
or U2433 (N_2433,N_1673,N_1854);
nor U2434 (N_2434,N_1673,N_1578);
nor U2435 (N_2435,N_1606,N_1698);
or U2436 (N_2436,N_1756,N_1529);
nand U2437 (N_2437,N_1778,N_1692);
or U2438 (N_2438,N_1512,N_1749);
nand U2439 (N_2439,N_1770,N_1962);
or U2440 (N_2440,N_1730,N_1917);
nand U2441 (N_2441,N_1835,N_1710);
nand U2442 (N_2442,N_1558,N_1577);
and U2443 (N_2443,N_1820,N_1848);
nor U2444 (N_2444,N_1595,N_1940);
or U2445 (N_2445,N_1518,N_1800);
or U2446 (N_2446,N_1846,N_1851);
nand U2447 (N_2447,N_1624,N_1697);
or U2448 (N_2448,N_1989,N_1512);
nand U2449 (N_2449,N_1979,N_1857);
xnor U2450 (N_2450,N_1882,N_1608);
nand U2451 (N_2451,N_1856,N_1609);
nand U2452 (N_2452,N_1973,N_1656);
and U2453 (N_2453,N_1619,N_1837);
xnor U2454 (N_2454,N_1786,N_1704);
nor U2455 (N_2455,N_1901,N_1752);
or U2456 (N_2456,N_1938,N_1534);
or U2457 (N_2457,N_1569,N_1960);
or U2458 (N_2458,N_1589,N_1522);
or U2459 (N_2459,N_1849,N_1783);
or U2460 (N_2460,N_1635,N_1763);
xnor U2461 (N_2461,N_1836,N_1975);
xor U2462 (N_2462,N_1509,N_1578);
xor U2463 (N_2463,N_1515,N_1881);
or U2464 (N_2464,N_1763,N_1940);
nor U2465 (N_2465,N_1993,N_1701);
nand U2466 (N_2466,N_1889,N_1696);
or U2467 (N_2467,N_1767,N_1884);
nor U2468 (N_2468,N_1984,N_1819);
xor U2469 (N_2469,N_1628,N_1608);
nand U2470 (N_2470,N_1732,N_1726);
nand U2471 (N_2471,N_1558,N_1792);
nand U2472 (N_2472,N_1713,N_1830);
nor U2473 (N_2473,N_1893,N_1961);
and U2474 (N_2474,N_1813,N_1752);
nand U2475 (N_2475,N_1816,N_1906);
nor U2476 (N_2476,N_1571,N_1848);
nand U2477 (N_2477,N_1981,N_1895);
and U2478 (N_2478,N_1743,N_1823);
xor U2479 (N_2479,N_1720,N_1501);
and U2480 (N_2480,N_1795,N_1866);
nand U2481 (N_2481,N_1756,N_1938);
and U2482 (N_2482,N_1969,N_1785);
or U2483 (N_2483,N_1833,N_1628);
and U2484 (N_2484,N_1629,N_1792);
nand U2485 (N_2485,N_1896,N_1676);
nand U2486 (N_2486,N_1955,N_1959);
and U2487 (N_2487,N_1772,N_1525);
and U2488 (N_2488,N_1981,N_1940);
and U2489 (N_2489,N_1502,N_1709);
and U2490 (N_2490,N_1712,N_1749);
and U2491 (N_2491,N_1828,N_1639);
nand U2492 (N_2492,N_1633,N_1513);
or U2493 (N_2493,N_1948,N_1647);
or U2494 (N_2494,N_1717,N_1535);
and U2495 (N_2495,N_1698,N_1792);
or U2496 (N_2496,N_1941,N_1861);
and U2497 (N_2497,N_1979,N_1976);
nor U2498 (N_2498,N_1829,N_1824);
and U2499 (N_2499,N_1702,N_1907);
or U2500 (N_2500,N_2160,N_2470);
or U2501 (N_2501,N_2419,N_2050);
or U2502 (N_2502,N_2319,N_2130);
nand U2503 (N_2503,N_2210,N_2161);
or U2504 (N_2504,N_2110,N_2424);
nor U2505 (N_2505,N_2144,N_2201);
and U2506 (N_2506,N_2458,N_2312);
and U2507 (N_2507,N_2003,N_2199);
or U2508 (N_2508,N_2062,N_2125);
and U2509 (N_2509,N_2432,N_2163);
nor U2510 (N_2510,N_2485,N_2385);
or U2511 (N_2511,N_2445,N_2299);
nand U2512 (N_2512,N_2353,N_2084);
nand U2513 (N_2513,N_2051,N_2472);
nor U2514 (N_2514,N_2049,N_2309);
or U2515 (N_2515,N_2376,N_2268);
and U2516 (N_2516,N_2406,N_2282);
nor U2517 (N_2517,N_2134,N_2303);
nor U2518 (N_2518,N_2129,N_2178);
or U2519 (N_2519,N_2039,N_2416);
xnor U2520 (N_2520,N_2434,N_2459);
and U2521 (N_2521,N_2214,N_2088);
or U2522 (N_2522,N_2090,N_2253);
or U2523 (N_2523,N_2438,N_2141);
or U2524 (N_2524,N_2055,N_2227);
and U2525 (N_2525,N_2043,N_2495);
and U2526 (N_2526,N_2415,N_2232);
nor U2527 (N_2527,N_2302,N_2234);
nor U2528 (N_2528,N_2475,N_2258);
nand U2529 (N_2529,N_2273,N_2159);
nand U2530 (N_2530,N_2468,N_2208);
and U2531 (N_2531,N_2063,N_2143);
or U2532 (N_2532,N_2339,N_2118);
nand U2533 (N_2533,N_2379,N_2193);
nor U2534 (N_2534,N_2436,N_2198);
or U2535 (N_2535,N_2386,N_2172);
xor U2536 (N_2536,N_2173,N_2204);
and U2537 (N_2537,N_2481,N_2333);
nor U2538 (N_2538,N_2146,N_2133);
xnor U2539 (N_2539,N_2292,N_2285);
and U2540 (N_2540,N_2311,N_2287);
nor U2541 (N_2541,N_2404,N_2132);
and U2542 (N_2542,N_2382,N_2097);
or U2543 (N_2543,N_2412,N_2023);
nor U2544 (N_2544,N_2346,N_2449);
xnor U2545 (N_2545,N_2479,N_2196);
nand U2546 (N_2546,N_2408,N_2200);
xnor U2547 (N_2547,N_2126,N_2493);
or U2548 (N_2548,N_2153,N_2070);
nor U2549 (N_2549,N_2447,N_2036);
and U2550 (N_2550,N_2068,N_2295);
nor U2551 (N_2551,N_2325,N_2454);
and U2552 (N_2552,N_2139,N_2212);
nor U2553 (N_2553,N_2409,N_2174);
or U2554 (N_2554,N_2347,N_2122);
nor U2555 (N_2555,N_2188,N_2136);
nand U2556 (N_2556,N_2367,N_2168);
nor U2557 (N_2557,N_2250,N_2306);
xor U2558 (N_2558,N_2262,N_2082);
or U2559 (N_2559,N_2357,N_2237);
or U2560 (N_2560,N_2446,N_2444);
and U2561 (N_2561,N_2344,N_2140);
or U2562 (N_2562,N_2042,N_2358);
nand U2563 (N_2563,N_2076,N_2480);
nand U2564 (N_2564,N_2016,N_2102);
nor U2565 (N_2565,N_2395,N_2158);
and U2566 (N_2566,N_2451,N_2297);
and U2567 (N_2567,N_2332,N_2079);
nor U2568 (N_2568,N_2226,N_2289);
nand U2569 (N_2569,N_2047,N_2330);
xor U2570 (N_2570,N_2264,N_2027);
nor U2571 (N_2571,N_2114,N_2372);
nor U2572 (N_2572,N_2064,N_2067);
xnor U2573 (N_2573,N_2467,N_2370);
and U2574 (N_2574,N_2059,N_2457);
nand U2575 (N_2575,N_2257,N_2298);
xnor U2576 (N_2576,N_2041,N_2286);
or U2577 (N_2577,N_2336,N_2222);
or U2578 (N_2578,N_2120,N_2383);
xor U2579 (N_2579,N_2279,N_2020);
nor U2580 (N_2580,N_2243,N_2101);
or U2581 (N_2581,N_2033,N_2487);
and U2582 (N_2582,N_2037,N_2006);
nand U2583 (N_2583,N_2350,N_2320);
nand U2584 (N_2584,N_2075,N_2281);
nand U2585 (N_2585,N_2308,N_2327);
nand U2586 (N_2586,N_2443,N_2260);
and U2587 (N_2587,N_2414,N_2440);
and U2588 (N_2588,N_2078,N_2484);
nor U2589 (N_2589,N_2307,N_2486);
nand U2590 (N_2590,N_2028,N_2058);
nor U2591 (N_2591,N_2491,N_2393);
or U2592 (N_2592,N_2013,N_2164);
or U2593 (N_2593,N_2032,N_2496);
xnor U2594 (N_2594,N_2004,N_2124);
nand U2595 (N_2595,N_2329,N_2239);
or U2596 (N_2596,N_2489,N_2442);
and U2597 (N_2597,N_2430,N_2038);
nor U2598 (N_2598,N_2046,N_2280);
and U2599 (N_2599,N_2396,N_2324);
and U2600 (N_2600,N_2207,N_2151);
or U2601 (N_2601,N_2190,N_2394);
xor U2602 (N_2602,N_2462,N_2147);
or U2603 (N_2603,N_2411,N_2015);
and U2604 (N_2604,N_2398,N_2321);
or U2605 (N_2605,N_2202,N_2094);
nand U2606 (N_2606,N_2313,N_2030);
nor U2607 (N_2607,N_2403,N_2065);
xor U2608 (N_2608,N_2235,N_2351);
nand U2609 (N_2609,N_2345,N_2213);
nor U2610 (N_2610,N_2230,N_2040);
and U2611 (N_2611,N_2490,N_2275);
and U2612 (N_2612,N_2310,N_2294);
or U2613 (N_2613,N_2269,N_2053);
nor U2614 (N_2614,N_2123,N_2099);
nor U2615 (N_2615,N_2209,N_2181);
xnor U2616 (N_2616,N_2361,N_2035);
or U2617 (N_2617,N_2420,N_2087);
or U2618 (N_2618,N_2267,N_2244);
nand U2619 (N_2619,N_2219,N_2096);
xor U2620 (N_2620,N_2340,N_2450);
nor U2621 (N_2621,N_2005,N_2331);
or U2622 (N_2622,N_2113,N_2375);
nand U2623 (N_2623,N_2391,N_2228);
or U2624 (N_2624,N_2138,N_2407);
and U2625 (N_2625,N_2381,N_2453);
nor U2626 (N_2626,N_2107,N_2322);
or U2627 (N_2627,N_2056,N_2211);
or U2628 (N_2628,N_2012,N_2413);
nand U2629 (N_2629,N_2195,N_2492);
or U2630 (N_2630,N_2483,N_2494);
nand U2631 (N_2631,N_2441,N_2261);
nand U2632 (N_2632,N_2352,N_2182);
or U2633 (N_2633,N_2187,N_2334);
and U2634 (N_2634,N_2137,N_2074);
nand U2635 (N_2635,N_2240,N_2488);
or U2636 (N_2636,N_2417,N_2498);
and U2637 (N_2637,N_2354,N_2265);
nor U2638 (N_2638,N_2000,N_2176);
nor U2639 (N_2639,N_2103,N_2247);
and U2640 (N_2640,N_2460,N_2183);
nand U2641 (N_2641,N_2014,N_2474);
nand U2642 (N_2642,N_2105,N_2071);
nor U2643 (N_2643,N_2439,N_2116);
nand U2644 (N_2644,N_2184,N_2337);
or U2645 (N_2645,N_2215,N_2373);
xor U2646 (N_2646,N_2166,N_2288);
nor U2647 (N_2647,N_2425,N_2377);
and U2648 (N_2648,N_2085,N_2127);
or U2649 (N_2649,N_2363,N_2115);
or U2650 (N_2650,N_2206,N_2044);
or U2651 (N_2651,N_2179,N_2384);
or U2652 (N_2652,N_2314,N_2323);
nand U2653 (N_2653,N_2301,N_2304);
xnor U2654 (N_2654,N_2152,N_2343);
or U2655 (N_2655,N_2186,N_2316);
and U2656 (N_2656,N_2368,N_2400);
or U2657 (N_2657,N_2429,N_2223);
or U2658 (N_2658,N_2111,N_2131);
and U2659 (N_2659,N_2191,N_2401);
or U2660 (N_2660,N_2052,N_2119);
or U2661 (N_2661,N_2469,N_2095);
and U2662 (N_2662,N_2410,N_2142);
nand U2663 (N_2663,N_2177,N_2477);
or U2664 (N_2664,N_2271,N_2335);
nand U2665 (N_2665,N_2045,N_2274);
nor U2666 (N_2666,N_2418,N_2388);
or U2667 (N_2667,N_2093,N_2326);
and U2668 (N_2668,N_2380,N_2389);
nor U2669 (N_2669,N_2248,N_2175);
xnor U2670 (N_2670,N_2154,N_2010);
and U2671 (N_2671,N_2318,N_2399);
nor U2672 (N_2672,N_2100,N_2378);
nand U2673 (N_2673,N_2149,N_2435);
nand U2674 (N_2674,N_2021,N_2083);
and U2675 (N_2675,N_2364,N_2162);
and U2676 (N_2676,N_2251,N_2155);
nor U2677 (N_2677,N_2465,N_2148);
nand U2678 (N_2678,N_2192,N_2048);
or U2679 (N_2679,N_2092,N_2291);
nand U2680 (N_2680,N_2236,N_2098);
nor U2681 (N_2681,N_2106,N_2001);
or U2682 (N_2682,N_2205,N_2077);
and U2683 (N_2683,N_2073,N_2194);
or U2684 (N_2684,N_2255,N_2342);
and U2685 (N_2685,N_2348,N_2349);
and U2686 (N_2686,N_2017,N_2089);
or U2687 (N_2687,N_2448,N_2167);
and U2688 (N_2688,N_2437,N_2170);
and U2689 (N_2689,N_2455,N_2217);
nor U2690 (N_2690,N_2452,N_2290);
nor U2691 (N_2691,N_2428,N_2026);
nand U2692 (N_2692,N_2225,N_2054);
nor U2693 (N_2693,N_2360,N_2189);
and U2694 (N_2694,N_2220,N_2296);
and U2695 (N_2695,N_2397,N_2293);
nor U2696 (N_2696,N_2266,N_2072);
nand U2697 (N_2697,N_2390,N_2471);
nor U2698 (N_2698,N_2008,N_2387);
and U2699 (N_2699,N_2157,N_2366);
and U2700 (N_2700,N_2229,N_2371);
nand U2701 (N_2701,N_2018,N_2423);
xor U2702 (N_2702,N_2185,N_2081);
or U2703 (N_2703,N_2150,N_2007);
nand U2704 (N_2704,N_2080,N_2060);
and U2705 (N_2705,N_2197,N_2109);
and U2706 (N_2706,N_2238,N_2405);
and U2707 (N_2707,N_2218,N_2019);
or U2708 (N_2708,N_2277,N_2476);
and U2709 (N_2709,N_2482,N_2104);
nand U2710 (N_2710,N_2369,N_2433);
nor U2711 (N_2711,N_2402,N_2135);
or U2712 (N_2712,N_2112,N_2431);
and U2713 (N_2713,N_2057,N_2025);
nand U2714 (N_2714,N_2252,N_2233);
nand U2715 (N_2715,N_2221,N_2022);
or U2716 (N_2716,N_2422,N_2355);
and U2717 (N_2717,N_2463,N_2338);
nand U2718 (N_2718,N_2362,N_2421);
xnor U2719 (N_2719,N_2203,N_2456);
nor U2720 (N_2720,N_2263,N_2478);
and U2721 (N_2721,N_2091,N_2254);
or U2722 (N_2722,N_2359,N_2128);
nor U2723 (N_2723,N_2024,N_2117);
and U2724 (N_2724,N_2121,N_2328);
nand U2725 (N_2725,N_2108,N_2246);
and U2726 (N_2726,N_2034,N_2061);
or U2727 (N_2727,N_2029,N_2245);
and U2728 (N_2728,N_2171,N_2317);
nand U2729 (N_2729,N_2165,N_2392);
nand U2730 (N_2730,N_2278,N_2341);
and U2731 (N_2731,N_2241,N_2300);
nand U2732 (N_2732,N_2315,N_2169);
nor U2733 (N_2733,N_2069,N_2066);
nand U2734 (N_2734,N_2283,N_2466);
nor U2735 (N_2735,N_2002,N_2374);
or U2736 (N_2736,N_2497,N_2009);
and U2737 (N_2737,N_2231,N_2270);
nand U2738 (N_2738,N_2461,N_2305);
xnor U2739 (N_2739,N_2276,N_2180);
or U2740 (N_2740,N_2272,N_2499);
or U2741 (N_2741,N_2256,N_2464);
and U2742 (N_2742,N_2216,N_2242);
nand U2743 (N_2743,N_2284,N_2145);
nand U2744 (N_2744,N_2249,N_2259);
nor U2745 (N_2745,N_2427,N_2365);
nand U2746 (N_2746,N_2426,N_2473);
or U2747 (N_2747,N_2356,N_2156);
nor U2748 (N_2748,N_2011,N_2224);
or U2749 (N_2749,N_2086,N_2031);
or U2750 (N_2750,N_2271,N_2387);
and U2751 (N_2751,N_2173,N_2045);
or U2752 (N_2752,N_2376,N_2467);
and U2753 (N_2753,N_2380,N_2075);
nand U2754 (N_2754,N_2128,N_2459);
and U2755 (N_2755,N_2186,N_2276);
xnor U2756 (N_2756,N_2305,N_2224);
xor U2757 (N_2757,N_2059,N_2233);
nand U2758 (N_2758,N_2306,N_2149);
nor U2759 (N_2759,N_2146,N_2399);
xor U2760 (N_2760,N_2360,N_2391);
nand U2761 (N_2761,N_2288,N_2259);
nor U2762 (N_2762,N_2447,N_2058);
and U2763 (N_2763,N_2255,N_2340);
nand U2764 (N_2764,N_2232,N_2310);
nand U2765 (N_2765,N_2003,N_2190);
xnor U2766 (N_2766,N_2444,N_2127);
or U2767 (N_2767,N_2233,N_2015);
or U2768 (N_2768,N_2232,N_2465);
nand U2769 (N_2769,N_2474,N_2402);
nor U2770 (N_2770,N_2314,N_2405);
nor U2771 (N_2771,N_2337,N_2089);
or U2772 (N_2772,N_2148,N_2269);
xnor U2773 (N_2773,N_2227,N_2413);
xnor U2774 (N_2774,N_2309,N_2492);
and U2775 (N_2775,N_2479,N_2269);
or U2776 (N_2776,N_2499,N_2443);
nand U2777 (N_2777,N_2162,N_2065);
or U2778 (N_2778,N_2181,N_2244);
and U2779 (N_2779,N_2011,N_2316);
nand U2780 (N_2780,N_2453,N_2290);
xnor U2781 (N_2781,N_2216,N_2063);
nor U2782 (N_2782,N_2018,N_2122);
and U2783 (N_2783,N_2337,N_2125);
nor U2784 (N_2784,N_2130,N_2089);
nand U2785 (N_2785,N_2002,N_2214);
and U2786 (N_2786,N_2374,N_2040);
and U2787 (N_2787,N_2199,N_2014);
and U2788 (N_2788,N_2417,N_2042);
and U2789 (N_2789,N_2453,N_2437);
nor U2790 (N_2790,N_2385,N_2251);
and U2791 (N_2791,N_2092,N_2116);
nand U2792 (N_2792,N_2053,N_2083);
or U2793 (N_2793,N_2486,N_2179);
and U2794 (N_2794,N_2233,N_2022);
nor U2795 (N_2795,N_2493,N_2102);
and U2796 (N_2796,N_2478,N_2296);
and U2797 (N_2797,N_2273,N_2118);
or U2798 (N_2798,N_2077,N_2377);
and U2799 (N_2799,N_2069,N_2243);
and U2800 (N_2800,N_2078,N_2279);
nor U2801 (N_2801,N_2177,N_2156);
nand U2802 (N_2802,N_2476,N_2058);
and U2803 (N_2803,N_2057,N_2080);
or U2804 (N_2804,N_2479,N_2092);
or U2805 (N_2805,N_2290,N_2221);
nand U2806 (N_2806,N_2192,N_2056);
and U2807 (N_2807,N_2461,N_2044);
or U2808 (N_2808,N_2396,N_2472);
xor U2809 (N_2809,N_2123,N_2263);
and U2810 (N_2810,N_2080,N_2261);
nand U2811 (N_2811,N_2421,N_2414);
and U2812 (N_2812,N_2183,N_2360);
xnor U2813 (N_2813,N_2117,N_2356);
nand U2814 (N_2814,N_2041,N_2302);
or U2815 (N_2815,N_2216,N_2145);
nand U2816 (N_2816,N_2127,N_2317);
nor U2817 (N_2817,N_2299,N_2123);
or U2818 (N_2818,N_2265,N_2102);
and U2819 (N_2819,N_2475,N_2260);
or U2820 (N_2820,N_2253,N_2122);
nand U2821 (N_2821,N_2143,N_2171);
and U2822 (N_2822,N_2294,N_2484);
or U2823 (N_2823,N_2287,N_2231);
xnor U2824 (N_2824,N_2197,N_2322);
and U2825 (N_2825,N_2134,N_2389);
nor U2826 (N_2826,N_2460,N_2177);
nand U2827 (N_2827,N_2341,N_2440);
nand U2828 (N_2828,N_2044,N_2221);
nor U2829 (N_2829,N_2476,N_2089);
and U2830 (N_2830,N_2004,N_2154);
and U2831 (N_2831,N_2436,N_2183);
or U2832 (N_2832,N_2450,N_2240);
and U2833 (N_2833,N_2036,N_2428);
nand U2834 (N_2834,N_2053,N_2107);
nand U2835 (N_2835,N_2135,N_2328);
nand U2836 (N_2836,N_2138,N_2218);
and U2837 (N_2837,N_2377,N_2476);
nor U2838 (N_2838,N_2069,N_2005);
nand U2839 (N_2839,N_2019,N_2327);
or U2840 (N_2840,N_2109,N_2291);
nand U2841 (N_2841,N_2154,N_2037);
nand U2842 (N_2842,N_2073,N_2101);
and U2843 (N_2843,N_2135,N_2373);
or U2844 (N_2844,N_2064,N_2217);
nand U2845 (N_2845,N_2415,N_2330);
nand U2846 (N_2846,N_2488,N_2232);
nor U2847 (N_2847,N_2492,N_2168);
nor U2848 (N_2848,N_2470,N_2053);
or U2849 (N_2849,N_2453,N_2386);
or U2850 (N_2850,N_2491,N_2490);
and U2851 (N_2851,N_2474,N_2060);
nor U2852 (N_2852,N_2374,N_2321);
and U2853 (N_2853,N_2364,N_2470);
or U2854 (N_2854,N_2200,N_2220);
or U2855 (N_2855,N_2109,N_2248);
and U2856 (N_2856,N_2429,N_2492);
and U2857 (N_2857,N_2372,N_2191);
or U2858 (N_2858,N_2447,N_2418);
nand U2859 (N_2859,N_2064,N_2159);
xnor U2860 (N_2860,N_2156,N_2060);
nor U2861 (N_2861,N_2487,N_2272);
or U2862 (N_2862,N_2120,N_2166);
or U2863 (N_2863,N_2167,N_2228);
nand U2864 (N_2864,N_2140,N_2313);
or U2865 (N_2865,N_2453,N_2317);
or U2866 (N_2866,N_2268,N_2083);
and U2867 (N_2867,N_2091,N_2281);
and U2868 (N_2868,N_2481,N_2241);
nand U2869 (N_2869,N_2484,N_2456);
and U2870 (N_2870,N_2163,N_2442);
or U2871 (N_2871,N_2412,N_2464);
xnor U2872 (N_2872,N_2278,N_2297);
nor U2873 (N_2873,N_2467,N_2225);
and U2874 (N_2874,N_2234,N_2478);
nor U2875 (N_2875,N_2190,N_2336);
or U2876 (N_2876,N_2217,N_2202);
and U2877 (N_2877,N_2046,N_2076);
nand U2878 (N_2878,N_2032,N_2029);
xor U2879 (N_2879,N_2408,N_2106);
nor U2880 (N_2880,N_2152,N_2055);
or U2881 (N_2881,N_2010,N_2406);
nor U2882 (N_2882,N_2038,N_2259);
or U2883 (N_2883,N_2233,N_2281);
or U2884 (N_2884,N_2222,N_2340);
or U2885 (N_2885,N_2407,N_2012);
nand U2886 (N_2886,N_2463,N_2485);
xor U2887 (N_2887,N_2473,N_2369);
and U2888 (N_2888,N_2467,N_2154);
or U2889 (N_2889,N_2088,N_2393);
nor U2890 (N_2890,N_2387,N_2405);
nand U2891 (N_2891,N_2049,N_2202);
or U2892 (N_2892,N_2346,N_2470);
nor U2893 (N_2893,N_2399,N_2008);
nand U2894 (N_2894,N_2355,N_2475);
and U2895 (N_2895,N_2459,N_2082);
and U2896 (N_2896,N_2442,N_2329);
nand U2897 (N_2897,N_2464,N_2175);
nand U2898 (N_2898,N_2079,N_2336);
and U2899 (N_2899,N_2105,N_2198);
and U2900 (N_2900,N_2192,N_2449);
nor U2901 (N_2901,N_2153,N_2268);
and U2902 (N_2902,N_2158,N_2108);
and U2903 (N_2903,N_2491,N_2249);
or U2904 (N_2904,N_2024,N_2278);
or U2905 (N_2905,N_2148,N_2357);
and U2906 (N_2906,N_2066,N_2202);
or U2907 (N_2907,N_2454,N_2194);
nand U2908 (N_2908,N_2179,N_2365);
nand U2909 (N_2909,N_2262,N_2063);
xor U2910 (N_2910,N_2097,N_2297);
nand U2911 (N_2911,N_2131,N_2459);
or U2912 (N_2912,N_2304,N_2276);
xor U2913 (N_2913,N_2436,N_2026);
nand U2914 (N_2914,N_2427,N_2020);
xnor U2915 (N_2915,N_2216,N_2059);
xnor U2916 (N_2916,N_2072,N_2042);
and U2917 (N_2917,N_2402,N_2371);
nor U2918 (N_2918,N_2342,N_2260);
nand U2919 (N_2919,N_2167,N_2332);
or U2920 (N_2920,N_2306,N_2449);
xnor U2921 (N_2921,N_2290,N_2340);
and U2922 (N_2922,N_2336,N_2424);
and U2923 (N_2923,N_2272,N_2396);
or U2924 (N_2924,N_2278,N_2008);
or U2925 (N_2925,N_2091,N_2111);
and U2926 (N_2926,N_2003,N_2191);
nor U2927 (N_2927,N_2440,N_2284);
nand U2928 (N_2928,N_2278,N_2326);
nor U2929 (N_2929,N_2089,N_2438);
and U2930 (N_2930,N_2328,N_2006);
nand U2931 (N_2931,N_2079,N_2115);
nand U2932 (N_2932,N_2431,N_2297);
and U2933 (N_2933,N_2432,N_2067);
nor U2934 (N_2934,N_2254,N_2140);
and U2935 (N_2935,N_2450,N_2380);
nor U2936 (N_2936,N_2347,N_2224);
and U2937 (N_2937,N_2386,N_2416);
or U2938 (N_2938,N_2025,N_2089);
and U2939 (N_2939,N_2113,N_2351);
nand U2940 (N_2940,N_2335,N_2081);
and U2941 (N_2941,N_2323,N_2335);
nand U2942 (N_2942,N_2466,N_2039);
and U2943 (N_2943,N_2068,N_2327);
nor U2944 (N_2944,N_2018,N_2184);
or U2945 (N_2945,N_2291,N_2360);
nor U2946 (N_2946,N_2263,N_2063);
or U2947 (N_2947,N_2429,N_2338);
xnor U2948 (N_2948,N_2212,N_2405);
nor U2949 (N_2949,N_2337,N_2378);
and U2950 (N_2950,N_2319,N_2350);
or U2951 (N_2951,N_2322,N_2075);
xnor U2952 (N_2952,N_2455,N_2261);
xnor U2953 (N_2953,N_2164,N_2337);
and U2954 (N_2954,N_2220,N_2034);
or U2955 (N_2955,N_2328,N_2046);
nor U2956 (N_2956,N_2023,N_2409);
or U2957 (N_2957,N_2251,N_2073);
nor U2958 (N_2958,N_2009,N_2364);
or U2959 (N_2959,N_2488,N_2188);
xor U2960 (N_2960,N_2401,N_2017);
or U2961 (N_2961,N_2285,N_2488);
nor U2962 (N_2962,N_2366,N_2392);
or U2963 (N_2963,N_2082,N_2449);
xor U2964 (N_2964,N_2473,N_2305);
xnor U2965 (N_2965,N_2490,N_2225);
or U2966 (N_2966,N_2487,N_2040);
and U2967 (N_2967,N_2088,N_2007);
xor U2968 (N_2968,N_2395,N_2088);
or U2969 (N_2969,N_2294,N_2252);
nor U2970 (N_2970,N_2240,N_2296);
nand U2971 (N_2971,N_2454,N_2341);
nand U2972 (N_2972,N_2387,N_2350);
or U2973 (N_2973,N_2371,N_2208);
or U2974 (N_2974,N_2208,N_2017);
xor U2975 (N_2975,N_2282,N_2148);
nor U2976 (N_2976,N_2022,N_2167);
nand U2977 (N_2977,N_2305,N_2338);
or U2978 (N_2978,N_2466,N_2158);
or U2979 (N_2979,N_2134,N_2214);
and U2980 (N_2980,N_2227,N_2193);
or U2981 (N_2981,N_2401,N_2371);
nand U2982 (N_2982,N_2285,N_2229);
and U2983 (N_2983,N_2290,N_2450);
or U2984 (N_2984,N_2247,N_2156);
nand U2985 (N_2985,N_2012,N_2326);
and U2986 (N_2986,N_2178,N_2031);
nor U2987 (N_2987,N_2208,N_2305);
xor U2988 (N_2988,N_2311,N_2007);
nor U2989 (N_2989,N_2139,N_2374);
and U2990 (N_2990,N_2314,N_2340);
nor U2991 (N_2991,N_2278,N_2128);
xor U2992 (N_2992,N_2090,N_2220);
and U2993 (N_2993,N_2018,N_2491);
nand U2994 (N_2994,N_2259,N_2155);
or U2995 (N_2995,N_2304,N_2385);
nor U2996 (N_2996,N_2406,N_2078);
and U2997 (N_2997,N_2402,N_2113);
nor U2998 (N_2998,N_2384,N_2256);
nor U2999 (N_2999,N_2482,N_2312);
nand UO_0 (O_0,N_2586,N_2560);
or UO_1 (O_1,N_2922,N_2698);
or UO_2 (O_2,N_2642,N_2915);
nand UO_3 (O_3,N_2873,N_2722);
or UO_4 (O_4,N_2601,N_2739);
xnor UO_5 (O_5,N_2983,N_2847);
nand UO_6 (O_6,N_2743,N_2605);
nand UO_7 (O_7,N_2748,N_2853);
and UO_8 (O_8,N_2704,N_2762);
and UO_9 (O_9,N_2726,N_2639);
or UO_10 (O_10,N_2819,N_2582);
and UO_11 (O_11,N_2737,N_2815);
and UO_12 (O_12,N_2969,N_2868);
xnor UO_13 (O_13,N_2970,N_2745);
nand UO_14 (O_14,N_2565,N_2747);
or UO_15 (O_15,N_2643,N_2651);
xor UO_16 (O_16,N_2557,N_2519);
xor UO_17 (O_17,N_2856,N_2555);
or UO_18 (O_18,N_2545,N_2501);
and UO_19 (O_19,N_2968,N_2829);
nor UO_20 (O_20,N_2988,N_2625);
and UO_21 (O_21,N_2547,N_2857);
and UO_22 (O_22,N_2621,N_2526);
nand UO_23 (O_23,N_2686,N_2575);
nor UO_24 (O_24,N_2966,N_2649);
nor UO_25 (O_25,N_2977,N_2691);
and UO_26 (O_26,N_2742,N_2578);
nand UO_27 (O_27,N_2515,N_2825);
nand UO_28 (O_28,N_2684,N_2832);
nand UO_29 (O_29,N_2725,N_2685);
and UO_30 (O_30,N_2812,N_2618);
xnor UO_31 (O_31,N_2690,N_2697);
or UO_32 (O_32,N_2602,N_2583);
and UO_33 (O_33,N_2597,N_2883);
nand UO_34 (O_34,N_2824,N_2965);
and UO_35 (O_35,N_2630,N_2727);
nor UO_36 (O_36,N_2718,N_2633);
nand UO_37 (O_37,N_2620,N_2660);
and UO_38 (O_38,N_2914,N_2559);
and UO_39 (O_39,N_2773,N_2652);
and UO_40 (O_40,N_2769,N_2913);
and UO_41 (O_41,N_2524,N_2801);
nor UO_42 (O_42,N_2837,N_2783);
nand UO_43 (O_43,N_2663,N_2779);
and UO_44 (O_44,N_2518,N_2667);
nor UO_45 (O_45,N_2821,N_2527);
and UO_46 (O_46,N_2796,N_2918);
and UO_47 (O_47,N_2880,N_2656);
xnor UO_48 (O_48,N_2994,N_2535);
and UO_49 (O_49,N_2788,N_2860);
and UO_50 (O_50,N_2755,N_2967);
and UO_51 (O_51,N_2613,N_2808);
nand UO_52 (O_52,N_2612,N_2644);
or UO_53 (O_53,N_2717,N_2973);
xnor UO_54 (O_54,N_2681,N_2648);
and UO_55 (O_55,N_2786,N_2710);
nor UO_56 (O_56,N_2525,N_2843);
xnor UO_57 (O_57,N_2879,N_2931);
nor UO_58 (O_58,N_2658,N_2987);
and UO_59 (O_59,N_2713,N_2768);
or UO_60 (O_60,N_2870,N_2905);
xor UO_61 (O_61,N_2841,N_2534);
xor UO_62 (O_62,N_2544,N_2834);
nor UO_63 (O_63,N_2816,N_2619);
or UO_64 (O_64,N_2731,N_2842);
and UO_65 (O_65,N_2509,N_2767);
nand UO_66 (O_66,N_2823,N_2705);
or UO_67 (O_67,N_2510,N_2886);
and UO_68 (O_68,N_2876,N_2603);
nand UO_69 (O_69,N_2916,N_2553);
or UO_70 (O_70,N_2673,N_2539);
and UO_71 (O_71,N_2887,N_2921);
nor UO_72 (O_72,N_2811,N_2571);
nand UO_73 (O_73,N_2687,N_2566);
or UO_74 (O_74,N_2599,N_2724);
nor UO_75 (O_75,N_2736,N_2871);
and UO_76 (O_76,N_2759,N_2982);
nand UO_77 (O_77,N_2807,N_2946);
and UO_78 (O_78,N_2814,N_2863);
nand UO_79 (O_79,N_2513,N_2588);
or UO_80 (O_80,N_2923,N_2953);
nand UO_81 (O_81,N_2984,N_2756);
nor UO_82 (O_82,N_2791,N_2949);
nor UO_83 (O_83,N_2552,N_2978);
nand UO_84 (O_84,N_2980,N_2934);
nor UO_85 (O_85,N_2865,N_2774);
and UO_86 (O_86,N_2634,N_2763);
nand UO_87 (O_87,N_2793,N_2610);
nor UO_88 (O_88,N_2794,N_2795);
and UO_89 (O_89,N_2878,N_2638);
nor UO_90 (O_90,N_2540,N_2720);
xnor UO_91 (O_91,N_2657,N_2666);
nand UO_92 (O_92,N_2912,N_2723);
nor UO_93 (O_93,N_2751,N_2520);
xnor UO_94 (O_94,N_2789,N_2888);
or UO_95 (O_95,N_2558,N_2668);
nor UO_96 (O_96,N_2563,N_2707);
and UO_97 (O_97,N_2805,N_2650);
nand UO_98 (O_98,N_2990,N_2584);
or UO_99 (O_99,N_2728,N_2986);
and UO_100 (O_100,N_2611,N_2874);
or UO_101 (O_101,N_2770,N_2564);
and UO_102 (O_102,N_2750,N_2875);
or UO_103 (O_103,N_2771,N_2904);
nand UO_104 (O_104,N_2647,N_2716);
and UO_105 (O_105,N_2766,N_2590);
and UO_106 (O_106,N_2901,N_2645);
xnor UO_107 (O_107,N_2662,N_2749);
and UO_108 (O_108,N_2635,N_2729);
nand UO_109 (O_109,N_2692,N_2682);
nand UO_110 (O_110,N_2730,N_2592);
nor UO_111 (O_111,N_2924,N_2993);
nand UO_112 (O_112,N_2721,N_2538);
xnor UO_113 (O_113,N_2975,N_2714);
nand UO_114 (O_114,N_2775,N_2679);
xor UO_115 (O_115,N_2587,N_2869);
or UO_116 (O_116,N_2971,N_2840);
and UO_117 (O_117,N_2581,N_2703);
or UO_118 (O_118,N_2764,N_2933);
or UO_119 (O_119,N_2694,N_2803);
and UO_120 (O_120,N_2542,N_2757);
or UO_121 (O_121,N_2778,N_2568);
nand UO_122 (O_122,N_2570,N_2661);
nand UO_123 (O_123,N_2595,N_2802);
or UO_124 (O_124,N_2699,N_2573);
xnor UO_125 (O_125,N_2740,N_2537);
nor UO_126 (O_126,N_2838,N_2689);
xnor UO_127 (O_127,N_2550,N_2974);
nand UO_128 (O_128,N_2512,N_2800);
nand UO_129 (O_129,N_2752,N_2855);
nand UO_130 (O_130,N_2503,N_2877);
and UO_131 (O_131,N_2623,N_2640);
xnor UO_132 (O_132,N_2511,N_2646);
nand UO_133 (O_133,N_2963,N_2893);
nand UO_134 (O_134,N_2835,N_2549);
and UO_135 (O_135,N_2958,N_2799);
nor UO_136 (O_136,N_2899,N_2536);
xnor UO_137 (O_137,N_2523,N_2678);
nand UO_138 (O_138,N_2909,N_2927);
and UO_139 (O_139,N_2693,N_2507);
and UO_140 (O_140,N_2517,N_2939);
or UO_141 (O_141,N_2632,N_2641);
nor UO_142 (O_142,N_2792,N_2891);
and UO_143 (O_143,N_2719,N_2996);
or UO_144 (O_144,N_2818,N_2735);
or UO_145 (O_145,N_2911,N_2906);
or UO_146 (O_146,N_2945,N_2700);
or UO_147 (O_147,N_2956,N_2827);
or UO_148 (O_148,N_2787,N_2951);
or UO_149 (O_149,N_2806,N_2695);
or UO_150 (O_150,N_2561,N_2947);
nand UO_151 (O_151,N_2920,N_2989);
and UO_152 (O_152,N_2585,N_2908);
or UO_153 (O_153,N_2896,N_2514);
nand UO_154 (O_154,N_2734,N_2627);
and UO_155 (O_155,N_2895,N_2972);
nand UO_156 (O_156,N_2543,N_2940);
and UO_157 (O_157,N_2897,N_2785);
and UO_158 (O_158,N_2894,N_2955);
xor UO_159 (O_159,N_2615,N_2741);
and UO_160 (O_160,N_2944,N_2579);
xnor UO_161 (O_161,N_2985,N_2997);
nor UO_162 (O_162,N_2839,N_2761);
xnor UO_163 (O_163,N_2950,N_2701);
nor UO_164 (O_164,N_2680,N_2859);
or UO_165 (O_165,N_2593,N_2861);
or UO_166 (O_166,N_2781,N_2554);
nand UO_167 (O_167,N_2851,N_2889);
and UO_168 (O_168,N_2532,N_2952);
and UO_169 (O_169,N_2797,N_2505);
or UO_170 (O_170,N_2903,N_2948);
nand UO_171 (O_171,N_2677,N_2674);
and UO_172 (O_172,N_2862,N_2754);
nor UO_173 (O_173,N_2589,N_2609);
nand UO_174 (O_174,N_2782,N_2919);
and UO_175 (O_175,N_2892,N_2683);
and UO_176 (O_176,N_2746,N_2500);
and UO_177 (O_177,N_2551,N_2910);
nand UO_178 (O_178,N_2932,N_2777);
nand UO_179 (O_179,N_2614,N_2577);
nand UO_180 (O_180,N_2607,N_2753);
nor UO_181 (O_181,N_2508,N_2772);
nor UO_182 (O_182,N_2846,N_2572);
nand UO_183 (O_183,N_2960,N_2935);
and UO_184 (O_184,N_2902,N_2964);
nand UO_185 (O_185,N_2715,N_2798);
and UO_186 (O_186,N_2784,N_2898);
nand UO_187 (O_187,N_2670,N_2959);
xor UO_188 (O_188,N_2676,N_2576);
or UO_189 (O_189,N_2654,N_2556);
nand UO_190 (O_190,N_2858,N_2521);
and UO_191 (O_191,N_2954,N_2885);
or UO_192 (O_192,N_2636,N_2849);
nand UO_193 (O_193,N_2999,N_2529);
nand UO_194 (O_194,N_2672,N_2907);
and UO_195 (O_195,N_2979,N_2991);
xnor UO_196 (O_196,N_2606,N_2900);
and UO_197 (O_197,N_2962,N_2598);
nor UO_198 (O_198,N_2830,N_2957);
nor UO_199 (O_199,N_2655,N_2569);
nor UO_200 (O_200,N_2995,N_2712);
nor UO_201 (O_201,N_2653,N_2810);
or UO_202 (O_202,N_2929,N_2664);
and UO_203 (O_203,N_2938,N_2502);
or UO_204 (O_204,N_2596,N_2702);
or UO_205 (O_205,N_2854,N_2516);
and UO_206 (O_206,N_2844,N_2930);
nor UO_207 (O_207,N_2659,N_2696);
and UO_208 (O_208,N_2976,N_2890);
and UO_209 (O_209,N_2675,N_2732);
or UO_210 (O_210,N_2617,N_2506);
nand UO_211 (O_211,N_2822,N_2594);
and UO_212 (O_212,N_2604,N_2917);
and UO_213 (O_213,N_2884,N_2671);
or UO_214 (O_214,N_2998,N_2942);
nand UO_215 (O_215,N_2608,N_2817);
and UO_216 (O_216,N_2925,N_2809);
nand UO_217 (O_217,N_2836,N_2541);
and UO_218 (O_218,N_2864,N_2733);
or UO_219 (O_219,N_2591,N_2928);
or UO_220 (O_220,N_2831,N_2531);
and UO_221 (O_221,N_2826,N_2937);
or UO_222 (O_222,N_2706,N_2626);
and UO_223 (O_223,N_2845,N_2562);
xnor UO_224 (O_224,N_2926,N_2738);
nand UO_225 (O_225,N_2629,N_2881);
nand UO_226 (O_226,N_2711,N_2504);
or UO_227 (O_227,N_2961,N_2804);
xnor UO_228 (O_228,N_2867,N_2981);
and UO_229 (O_229,N_2600,N_2850);
xnor UO_230 (O_230,N_2628,N_2624);
xor UO_231 (O_231,N_2872,N_2580);
nand UO_232 (O_232,N_2574,N_2522);
or UO_233 (O_233,N_2780,N_2665);
nor UO_234 (O_234,N_2709,N_2744);
or UO_235 (O_235,N_2828,N_2992);
nand UO_236 (O_236,N_2760,N_2882);
nand UO_237 (O_237,N_2776,N_2688);
or UO_238 (O_238,N_2813,N_2669);
or UO_239 (O_239,N_2790,N_2941);
and UO_240 (O_240,N_2533,N_2548);
nor UO_241 (O_241,N_2936,N_2852);
nand UO_242 (O_242,N_2765,N_2848);
nor UO_243 (O_243,N_2616,N_2567);
or UO_244 (O_244,N_2833,N_2631);
xnor UO_245 (O_245,N_2528,N_2820);
or UO_246 (O_246,N_2943,N_2530);
and UO_247 (O_247,N_2637,N_2866);
and UO_248 (O_248,N_2758,N_2708);
or UO_249 (O_249,N_2546,N_2622);
and UO_250 (O_250,N_2522,N_2774);
or UO_251 (O_251,N_2661,N_2546);
nand UO_252 (O_252,N_2712,N_2893);
or UO_253 (O_253,N_2588,N_2901);
and UO_254 (O_254,N_2756,N_2690);
and UO_255 (O_255,N_2544,N_2946);
and UO_256 (O_256,N_2582,N_2516);
nand UO_257 (O_257,N_2920,N_2977);
and UO_258 (O_258,N_2530,N_2622);
nor UO_259 (O_259,N_2637,N_2516);
nor UO_260 (O_260,N_2686,N_2568);
and UO_261 (O_261,N_2591,N_2651);
and UO_262 (O_262,N_2733,N_2567);
xor UO_263 (O_263,N_2673,N_2724);
or UO_264 (O_264,N_2787,N_2652);
nand UO_265 (O_265,N_2582,N_2909);
or UO_266 (O_266,N_2840,N_2681);
xnor UO_267 (O_267,N_2862,N_2611);
nor UO_268 (O_268,N_2703,N_2827);
and UO_269 (O_269,N_2896,N_2500);
xor UO_270 (O_270,N_2869,N_2638);
nor UO_271 (O_271,N_2858,N_2565);
nor UO_272 (O_272,N_2947,N_2558);
and UO_273 (O_273,N_2928,N_2833);
or UO_274 (O_274,N_2823,N_2698);
or UO_275 (O_275,N_2749,N_2631);
nand UO_276 (O_276,N_2931,N_2565);
and UO_277 (O_277,N_2595,N_2790);
nand UO_278 (O_278,N_2753,N_2573);
nor UO_279 (O_279,N_2815,N_2839);
or UO_280 (O_280,N_2830,N_2839);
and UO_281 (O_281,N_2559,N_2600);
or UO_282 (O_282,N_2982,N_2862);
or UO_283 (O_283,N_2920,N_2594);
xnor UO_284 (O_284,N_2959,N_2871);
nand UO_285 (O_285,N_2945,N_2820);
nand UO_286 (O_286,N_2783,N_2855);
nor UO_287 (O_287,N_2618,N_2769);
nand UO_288 (O_288,N_2577,N_2793);
xnor UO_289 (O_289,N_2962,N_2765);
nand UO_290 (O_290,N_2875,N_2517);
and UO_291 (O_291,N_2837,N_2705);
nor UO_292 (O_292,N_2751,N_2853);
or UO_293 (O_293,N_2791,N_2657);
xnor UO_294 (O_294,N_2590,N_2774);
nand UO_295 (O_295,N_2783,N_2925);
nand UO_296 (O_296,N_2597,N_2893);
nand UO_297 (O_297,N_2946,N_2799);
or UO_298 (O_298,N_2823,N_2806);
and UO_299 (O_299,N_2779,N_2710);
nor UO_300 (O_300,N_2950,N_2550);
nand UO_301 (O_301,N_2641,N_2939);
or UO_302 (O_302,N_2759,N_2904);
nor UO_303 (O_303,N_2686,N_2981);
or UO_304 (O_304,N_2966,N_2847);
or UO_305 (O_305,N_2980,N_2697);
nor UO_306 (O_306,N_2693,N_2801);
or UO_307 (O_307,N_2826,N_2676);
and UO_308 (O_308,N_2729,N_2963);
or UO_309 (O_309,N_2721,N_2946);
nand UO_310 (O_310,N_2509,N_2503);
nor UO_311 (O_311,N_2714,N_2583);
nand UO_312 (O_312,N_2989,N_2721);
nor UO_313 (O_313,N_2836,N_2543);
or UO_314 (O_314,N_2554,N_2610);
nor UO_315 (O_315,N_2504,N_2874);
or UO_316 (O_316,N_2967,N_2864);
or UO_317 (O_317,N_2766,N_2575);
nand UO_318 (O_318,N_2911,N_2613);
and UO_319 (O_319,N_2993,N_2913);
and UO_320 (O_320,N_2609,N_2939);
nand UO_321 (O_321,N_2951,N_2685);
and UO_322 (O_322,N_2955,N_2630);
nand UO_323 (O_323,N_2575,N_2813);
or UO_324 (O_324,N_2978,N_2886);
and UO_325 (O_325,N_2874,N_2549);
nor UO_326 (O_326,N_2599,N_2742);
and UO_327 (O_327,N_2714,N_2829);
nand UO_328 (O_328,N_2764,N_2854);
or UO_329 (O_329,N_2711,N_2789);
or UO_330 (O_330,N_2597,N_2948);
nand UO_331 (O_331,N_2811,N_2590);
and UO_332 (O_332,N_2731,N_2574);
nor UO_333 (O_333,N_2891,N_2573);
or UO_334 (O_334,N_2712,N_2555);
nor UO_335 (O_335,N_2870,N_2757);
xor UO_336 (O_336,N_2679,N_2823);
and UO_337 (O_337,N_2736,N_2514);
and UO_338 (O_338,N_2990,N_2891);
or UO_339 (O_339,N_2931,N_2537);
and UO_340 (O_340,N_2999,N_2780);
xnor UO_341 (O_341,N_2949,N_2642);
nand UO_342 (O_342,N_2926,N_2965);
and UO_343 (O_343,N_2732,N_2536);
nor UO_344 (O_344,N_2709,N_2600);
nand UO_345 (O_345,N_2534,N_2930);
xnor UO_346 (O_346,N_2657,N_2845);
or UO_347 (O_347,N_2819,N_2667);
nand UO_348 (O_348,N_2891,N_2529);
and UO_349 (O_349,N_2815,N_2538);
nand UO_350 (O_350,N_2978,N_2760);
nor UO_351 (O_351,N_2501,N_2616);
nand UO_352 (O_352,N_2716,N_2589);
nand UO_353 (O_353,N_2605,N_2928);
and UO_354 (O_354,N_2758,N_2743);
and UO_355 (O_355,N_2729,N_2849);
or UO_356 (O_356,N_2653,N_2564);
nor UO_357 (O_357,N_2777,N_2708);
nand UO_358 (O_358,N_2882,N_2969);
nand UO_359 (O_359,N_2944,N_2928);
nand UO_360 (O_360,N_2957,N_2561);
nor UO_361 (O_361,N_2592,N_2815);
nand UO_362 (O_362,N_2765,N_2724);
xor UO_363 (O_363,N_2977,N_2863);
or UO_364 (O_364,N_2738,N_2650);
nor UO_365 (O_365,N_2984,N_2874);
and UO_366 (O_366,N_2751,N_2878);
nor UO_367 (O_367,N_2898,N_2762);
nor UO_368 (O_368,N_2923,N_2838);
nand UO_369 (O_369,N_2514,N_2970);
nor UO_370 (O_370,N_2761,N_2939);
nand UO_371 (O_371,N_2890,N_2811);
or UO_372 (O_372,N_2537,N_2689);
nor UO_373 (O_373,N_2758,N_2647);
nand UO_374 (O_374,N_2967,N_2573);
xnor UO_375 (O_375,N_2732,N_2669);
or UO_376 (O_376,N_2572,N_2809);
nor UO_377 (O_377,N_2861,N_2618);
and UO_378 (O_378,N_2971,N_2987);
nor UO_379 (O_379,N_2651,N_2677);
or UO_380 (O_380,N_2814,N_2859);
or UO_381 (O_381,N_2657,N_2565);
or UO_382 (O_382,N_2915,N_2806);
or UO_383 (O_383,N_2684,N_2600);
nand UO_384 (O_384,N_2928,N_2702);
or UO_385 (O_385,N_2544,N_2634);
and UO_386 (O_386,N_2859,N_2511);
and UO_387 (O_387,N_2774,N_2868);
xnor UO_388 (O_388,N_2550,N_2609);
xor UO_389 (O_389,N_2694,N_2560);
xnor UO_390 (O_390,N_2918,N_2525);
nor UO_391 (O_391,N_2523,N_2593);
nor UO_392 (O_392,N_2802,N_2826);
nand UO_393 (O_393,N_2721,N_2662);
and UO_394 (O_394,N_2684,N_2646);
nand UO_395 (O_395,N_2997,N_2938);
or UO_396 (O_396,N_2742,N_2817);
xor UO_397 (O_397,N_2915,N_2810);
and UO_398 (O_398,N_2625,N_2676);
nor UO_399 (O_399,N_2683,N_2703);
or UO_400 (O_400,N_2518,N_2543);
and UO_401 (O_401,N_2623,N_2801);
and UO_402 (O_402,N_2700,N_2650);
nand UO_403 (O_403,N_2887,N_2843);
and UO_404 (O_404,N_2967,N_2983);
or UO_405 (O_405,N_2679,N_2898);
and UO_406 (O_406,N_2600,N_2941);
or UO_407 (O_407,N_2862,N_2980);
and UO_408 (O_408,N_2584,N_2681);
or UO_409 (O_409,N_2926,N_2960);
xnor UO_410 (O_410,N_2801,N_2898);
and UO_411 (O_411,N_2668,N_2876);
nor UO_412 (O_412,N_2859,N_2632);
or UO_413 (O_413,N_2637,N_2638);
xnor UO_414 (O_414,N_2547,N_2675);
or UO_415 (O_415,N_2638,N_2861);
nand UO_416 (O_416,N_2812,N_2819);
and UO_417 (O_417,N_2575,N_2828);
and UO_418 (O_418,N_2550,N_2694);
nor UO_419 (O_419,N_2607,N_2617);
nor UO_420 (O_420,N_2843,N_2953);
or UO_421 (O_421,N_2793,N_2777);
and UO_422 (O_422,N_2513,N_2775);
nand UO_423 (O_423,N_2734,N_2581);
or UO_424 (O_424,N_2924,N_2591);
or UO_425 (O_425,N_2939,N_2814);
or UO_426 (O_426,N_2709,N_2623);
nor UO_427 (O_427,N_2578,N_2616);
or UO_428 (O_428,N_2646,N_2790);
nor UO_429 (O_429,N_2974,N_2896);
or UO_430 (O_430,N_2575,N_2869);
or UO_431 (O_431,N_2975,N_2990);
or UO_432 (O_432,N_2711,N_2718);
or UO_433 (O_433,N_2513,N_2516);
and UO_434 (O_434,N_2952,N_2525);
and UO_435 (O_435,N_2984,N_2951);
nand UO_436 (O_436,N_2600,N_2802);
xor UO_437 (O_437,N_2753,N_2925);
nand UO_438 (O_438,N_2768,N_2668);
nor UO_439 (O_439,N_2502,N_2861);
nand UO_440 (O_440,N_2757,N_2911);
or UO_441 (O_441,N_2874,N_2827);
and UO_442 (O_442,N_2862,N_2523);
and UO_443 (O_443,N_2651,N_2834);
and UO_444 (O_444,N_2539,N_2779);
and UO_445 (O_445,N_2641,N_2938);
nor UO_446 (O_446,N_2702,N_2938);
nand UO_447 (O_447,N_2532,N_2894);
or UO_448 (O_448,N_2590,N_2578);
xor UO_449 (O_449,N_2911,N_2553);
nor UO_450 (O_450,N_2699,N_2714);
or UO_451 (O_451,N_2702,N_2792);
nor UO_452 (O_452,N_2549,N_2815);
nor UO_453 (O_453,N_2530,N_2708);
or UO_454 (O_454,N_2597,N_2695);
xnor UO_455 (O_455,N_2796,N_2693);
nor UO_456 (O_456,N_2670,N_2751);
nor UO_457 (O_457,N_2954,N_2825);
and UO_458 (O_458,N_2634,N_2823);
nand UO_459 (O_459,N_2885,N_2951);
or UO_460 (O_460,N_2601,N_2717);
and UO_461 (O_461,N_2861,N_2816);
xor UO_462 (O_462,N_2606,N_2767);
nand UO_463 (O_463,N_2617,N_2733);
and UO_464 (O_464,N_2590,N_2603);
and UO_465 (O_465,N_2687,N_2558);
nand UO_466 (O_466,N_2843,N_2906);
nand UO_467 (O_467,N_2564,N_2976);
or UO_468 (O_468,N_2826,N_2870);
or UO_469 (O_469,N_2910,N_2919);
nor UO_470 (O_470,N_2562,N_2675);
nand UO_471 (O_471,N_2545,N_2698);
nand UO_472 (O_472,N_2620,N_2510);
and UO_473 (O_473,N_2615,N_2913);
xor UO_474 (O_474,N_2518,N_2728);
nand UO_475 (O_475,N_2876,N_2651);
nor UO_476 (O_476,N_2643,N_2803);
nand UO_477 (O_477,N_2614,N_2972);
nand UO_478 (O_478,N_2857,N_2878);
and UO_479 (O_479,N_2926,N_2829);
nand UO_480 (O_480,N_2742,N_2664);
nand UO_481 (O_481,N_2764,N_2776);
nand UO_482 (O_482,N_2500,N_2881);
nand UO_483 (O_483,N_2876,N_2680);
nand UO_484 (O_484,N_2628,N_2733);
and UO_485 (O_485,N_2935,N_2967);
nor UO_486 (O_486,N_2693,N_2733);
nor UO_487 (O_487,N_2539,N_2811);
or UO_488 (O_488,N_2984,N_2576);
and UO_489 (O_489,N_2819,N_2862);
nand UO_490 (O_490,N_2670,N_2942);
nor UO_491 (O_491,N_2789,N_2600);
and UO_492 (O_492,N_2759,N_2528);
nand UO_493 (O_493,N_2833,N_2960);
xor UO_494 (O_494,N_2939,N_2960);
nand UO_495 (O_495,N_2881,N_2800);
xnor UO_496 (O_496,N_2568,N_2965);
or UO_497 (O_497,N_2536,N_2728);
nand UO_498 (O_498,N_2592,N_2610);
xnor UO_499 (O_499,N_2693,N_2795);
endmodule