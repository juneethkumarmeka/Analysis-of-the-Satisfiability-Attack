module basic_500_3000_500_6_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_303,In_473);
nand U1 (N_1,In_19,In_465);
or U2 (N_2,In_190,In_459);
nand U3 (N_3,In_67,In_396);
or U4 (N_4,In_362,In_429);
nand U5 (N_5,In_295,In_225);
or U6 (N_6,In_351,In_317);
and U7 (N_7,In_358,In_420);
and U8 (N_8,In_71,In_316);
nor U9 (N_9,In_361,In_187);
or U10 (N_10,In_308,In_155);
and U11 (N_11,In_436,In_109);
nor U12 (N_12,In_215,In_365);
or U13 (N_13,In_88,In_64);
and U14 (N_14,In_46,In_151);
or U15 (N_15,In_398,In_201);
nor U16 (N_16,In_68,In_194);
xnor U17 (N_17,In_57,In_17);
and U18 (N_18,In_205,In_291);
or U19 (N_19,In_179,In_206);
or U20 (N_20,In_412,In_258);
nor U21 (N_21,In_492,In_160);
xor U22 (N_22,In_448,In_402);
or U23 (N_23,In_350,In_241);
and U24 (N_24,In_52,In_18);
nor U25 (N_25,In_233,In_445);
nand U26 (N_26,In_208,In_313);
nand U27 (N_27,In_277,In_388);
and U28 (N_28,In_372,In_463);
and U29 (N_29,In_343,In_280);
and U30 (N_30,In_219,In_379);
or U31 (N_31,In_259,In_301);
nor U32 (N_32,In_103,In_374);
or U33 (N_33,In_2,In_76);
nor U34 (N_34,In_323,In_193);
and U35 (N_35,In_345,In_227);
nand U36 (N_36,In_127,In_83);
nand U37 (N_37,In_245,In_173);
nor U38 (N_38,In_477,In_276);
or U39 (N_39,In_421,In_114);
nor U40 (N_40,In_156,In_33);
or U41 (N_41,In_328,In_357);
nand U42 (N_42,In_407,In_55);
nand U43 (N_43,In_13,In_391);
nand U44 (N_44,In_457,In_380);
or U45 (N_45,In_441,In_311);
nand U46 (N_46,In_342,In_154);
and U47 (N_47,In_212,In_462);
nor U48 (N_48,In_229,In_352);
or U49 (N_49,In_108,In_366);
nand U50 (N_50,In_107,In_112);
or U51 (N_51,In_279,In_368);
and U52 (N_52,In_20,In_117);
nand U53 (N_53,In_326,In_369);
and U54 (N_54,In_164,In_24);
xnor U55 (N_55,In_135,In_221);
nand U56 (N_56,In_120,In_381);
or U57 (N_57,In_106,In_77);
and U58 (N_58,In_331,In_116);
or U59 (N_59,In_403,In_341);
xor U60 (N_60,In_228,In_296);
nor U61 (N_61,In_248,In_319);
and U62 (N_62,In_370,In_272);
nor U63 (N_63,In_257,In_184);
nand U64 (N_64,In_204,In_39);
nor U65 (N_65,In_455,In_192);
and U66 (N_66,In_183,In_200);
or U67 (N_67,In_474,In_26);
and U68 (N_68,In_485,In_386);
nand U69 (N_69,In_422,In_479);
nand U70 (N_70,In_136,In_314);
or U71 (N_71,In_25,In_143);
nand U72 (N_72,In_121,In_392);
or U73 (N_73,In_15,In_480);
nand U74 (N_74,In_446,In_415);
or U75 (N_75,In_167,In_254);
and U76 (N_76,In_253,In_373);
and U77 (N_77,In_125,In_191);
and U78 (N_78,In_393,In_409);
xor U79 (N_79,In_339,In_8);
xor U80 (N_80,In_82,In_250);
nor U81 (N_81,In_300,In_428);
or U82 (N_82,In_163,In_242);
and U83 (N_83,In_188,In_185);
nand U84 (N_84,In_130,In_483);
or U85 (N_85,In_476,In_261);
xor U86 (N_86,In_247,In_211);
and U87 (N_87,In_148,In_14);
or U88 (N_88,In_249,In_287);
or U89 (N_89,In_29,In_70);
and U90 (N_90,In_438,In_105);
nand U91 (N_91,In_404,In_62);
nand U92 (N_92,In_298,In_400);
nor U93 (N_93,In_307,In_213);
or U94 (N_94,In_84,In_499);
nor U95 (N_95,In_43,In_38);
and U96 (N_96,In_152,In_174);
nand U97 (N_97,In_81,In_222);
nor U98 (N_98,In_449,In_399);
nor U99 (N_99,In_431,In_115);
nand U100 (N_100,In_454,In_378);
or U101 (N_101,In_99,In_417);
nor U102 (N_102,In_195,In_432);
and U103 (N_103,In_51,In_90);
and U104 (N_104,In_496,In_58);
or U105 (N_105,In_230,In_356);
or U106 (N_106,In_210,In_390);
and U107 (N_107,In_299,In_59);
nor U108 (N_108,In_375,In_86);
nand U109 (N_109,In_158,In_85);
or U110 (N_110,In_377,In_203);
nand U111 (N_111,In_397,In_235);
or U112 (N_112,In_282,In_246);
nand U113 (N_113,In_10,In_270);
xor U114 (N_114,In_354,In_353);
nor U115 (N_115,In_267,In_252);
nand U116 (N_116,In_284,In_274);
or U117 (N_117,In_144,In_364);
nand U118 (N_118,In_433,In_336);
or U119 (N_119,In_478,In_294);
nand U120 (N_120,In_469,In_1);
or U121 (N_121,In_256,In_440);
nor U122 (N_122,In_31,In_132);
or U123 (N_123,In_334,In_425);
and U124 (N_124,In_110,In_202);
and U125 (N_125,In_292,In_170);
and U126 (N_126,In_122,In_315);
nor U127 (N_127,In_488,In_147);
or U128 (N_128,In_36,In_325);
nor U129 (N_129,In_118,In_444);
nand U130 (N_130,In_333,In_278);
and U131 (N_131,In_337,In_293);
or U132 (N_132,In_285,In_34);
or U133 (N_133,In_490,In_471);
and U134 (N_134,In_238,In_346);
nor U135 (N_135,In_489,In_74);
or U136 (N_136,In_56,In_162);
nor U137 (N_137,In_395,In_427);
and U138 (N_138,In_41,In_50);
or U139 (N_139,In_149,In_240);
nand U140 (N_140,In_451,In_54);
nand U141 (N_141,In_189,In_263);
or U142 (N_142,In_423,In_159);
nor U143 (N_143,In_80,In_217);
nor U144 (N_144,In_97,In_322);
nand U145 (N_145,In_165,In_452);
nand U146 (N_146,In_94,In_199);
xnor U147 (N_147,In_224,In_371);
and U148 (N_148,In_171,In_119);
nor U149 (N_149,In_239,In_231);
xor U150 (N_150,In_491,In_416);
or U151 (N_151,In_177,In_306);
and U152 (N_152,In_146,In_426);
or U153 (N_153,In_150,In_244);
nor U154 (N_154,In_61,In_321);
or U155 (N_155,In_102,In_157);
nor U156 (N_156,In_359,In_269);
nand U157 (N_157,In_45,In_35);
and U158 (N_158,In_63,In_218);
nor U159 (N_159,In_197,In_475);
and U160 (N_160,In_401,In_142);
nand U161 (N_161,In_139,In_271);
nand U162 (N_162,In_405,In_226);
nor U163 (N_163,In_23,In_140);
nor U164 (N_164,In_283,In_93);
or U165 (N_165,In_419,In_16);
or U166 (N_166,In_335,In_27);
nand U167 (N_167,In_141,In_349);
and U168 (N_168,In_22,In_338);
or U169 (N_169,In_355,In_12);
and U170 (N_170,In_464,In_42);
nor U171 (N_171,In_360,In_216);
or U172 (N_172,In_435,In_72);
or U173 (N_173,In_466,In_181);
or U174 (N_174,In_497,In_243);
nor U175 (N_175,In_30,In_264);
xnor U176 (N_176,In_53,In_6);
nand U177 (N_177,In_330,In_347);
and U178 (N_178,In_98,In_384);
and U179 (N_179,In_439,In_126);
and U180 (N_180,In_456,In_4);
and U181 (N_181,In_363,In_176);
or U182 (N_182,In_468,In_286);
nor U183 (N_183,In_430,In_289);
and U184 (N_184,In_234,In_111);
nor U185 (N_185,In_89,In_166);
xnor U186 (N_186,In_367,In_413);
or U187 (N_187,In_101,In_443);
xnor U188 (N_188,In_5,In_169);
or U189 (N_189,In_467,In_408);
or U190 (N_190,In_266,In_310);
or U191 (N_191,In_304,In_288);
or U192 (N_192,In_498,In_411);
nor U193 (N_193,In_66,In_268);
nand U194 (N_194,In_418,In_340);
xor U195 (N_195,In_251,In_410);
and U196 (N_196,In_133,In_145);
or U197 (N_197,In_137,In_214);
nor U198 (N_198,In_344,In_329);
xor U199 (N_199,In_182,In_387);
nor U200 (N_200,In_96,In_21);
and U201 (N_201,In_78,In_297);
nor U202 (N_202,In_186,In_79);
nand U203 (N_203,In_487,In_376);
nand U204 (N_204,In_450,In_494);
and U205 (N_205,In_232,In_32);
nand U206 (N_206,In_324,In_91);
or U207 (N_207,In_37,In_44);
and U208 (N_208,In_168,In_47);
or U209 (N_209,In_180,In_447);
nor U210 (N_210,In_442,In_394);
nor U211 (N_211,In_484,In_495);
nand U212 (N_212,In_262,In_95);
and U213 (N_213,In_255,In_138);
nor U214 (N_214,In_198,In_131);
nor U215 (N_215,In_220,In_123);
and U216 (N_216,In_223,In_458);
nand U217 (N_217,In_290,In_104);
or U218 (N_218,In_332,In_385);
nor U219 (N_219,In_237,In_172);
nand U220 (N_220,In_481,In_196);
nand U221 (N_221,In_461,In_178);
or U222 (N_222,In_320,In_327);
nand U223 (N_223,In_40,In_129);
and U224 (N_224,In_124,In_0);
nor U225 (N_225,In_73,In_100);
and U226 (N_226,In_48,In_348);
and U227 (N_227,In_28,In_414);
nand U228 (N_228,In_265,In_305);
nand U229 (N_229,In_434,In_209);
or U230 (N_230,In_134,In_312);
nor U231 (N_231,In_486,In_460);
or U232 (N_232,In_482,In_60);
nand U233 (N_233,In_383,In_406);
nand U234 (N_234,In_302,In_493);
and U235 (N_235,In_49,In_9);
and U236 (N_236,In_318,In_75);
or U237 (N_237,In_453,In_472);
or U238 (N_238,In_175,In_69);
nand U239 (N_239,In_161,In_113);
and U240 (N_240,In_207,In_309);
nand U241 (N_241,In_87,In_389);
or U242 (N_242,In_153,In_128);
nand U243 (N_243,In_470,In_65);
nor U244 (N_244,In_273,In_11);
or U245 (N_245,In_275,In_236);
and U246 (N_246,In_382,In_281);
or U247 (N_247,In_7,In_3);
nand U248 (N_248,In_92,In_437);
nor U249 (N_249,In_260,In_424);
and U250 (N_250,In_364,In_46);
or U251 (N_251,In_300,In_421);
or U252 (N_252,In_95,In_168);
or U253 (N_253,In_224,In_159);
nor U254 (N_254,In_21,In_112);
and U255 (N_255,In_274,In_489);
or U256 (N_256,In_462,In_348);
nand U257 (N_257,In_165,In_356);
nor U258 (N_258,In_105,In_335);
nor U259 (N_259,In_269,In_440);
or U260 (N_260,In_186,In_85);
and U261 (N_261,In_317,In_393);
nor U262 (N_262,In_80,In_396);
or U263 (N_263,In_335,In_237);
nor U264 (N_264,In_498,In_150);
and U265 (N_265,In_418,In_237);
nor U266 (N_266,In_371,In_50);
and U267 (N_267,In_188,In_13);
nand U268 (N_268,In_467,In_263);
and U269 (N_269,In_51,In_447);
nor U270 (N_270,In_342,In_110);
nand U271 (N_271,In_390,In_441);
nand U272 (N_272,In_490,In_179);
nand U273 (N_273,In_453,In_262);
and U274 (N_274,In_54,In_201);
xnor U275 (N_275,In_95,In_412);
or U276 (N_276,In_437,In_238);
and U277 (N_277,In_344,In_144);
nor U278 (N_278,In_152,In_76);
nand U279 (N_279,In_353,In_495);
or U280 (N_280,In_220,In_154);
and U281 (N_281,In_361,In_217);
nor U282 (N_282,In_282,In_446);
nand U283 (N_283,In_7,In_469);
nand U284 (N_284,In_407,In_169);
nand U285 (N_285,In_381,In_293);
or U286 (N_286,In_52,In_378);
nor U287 (N_287,In_121,In_260);
nand U288 (N_288,In_437,In_37);
and U289 (N_289,In_5,In_27);
nand U290 (N_290,In_186,In_377);
nor U291 (N_291,In_128,In_63);
nor U292 (N_292,In_83,In_203);
nand U293 (N_293,In_496,In_305);
and U294 (N_294,In_288,In_487);
and U295 (N_295,In_489,In_496);
nand U296 (N_296,In_307,In_178);
or U297 (N_297,In_109,In_271);
nor U298 (N_298,In_428,In_376);
nor U299 (N_299,In_94,In_53);
or U300 (N_300,In_75,In_57);
nor U301 (N_301,In_323,In_352);
or U302 (N_302,In_205,In_210);
or U303 (N_303,In_88,In_190);
nor U304 (N_304,In_481,In_220);
nor U305 (N_305,In_174,In_20);
and U306 (N_306,In_470,In_176);
or U307 (N_307,In_29,In_453);
and U308 (N_308,In_169,In_196);
and U309 (N_309,In_427,In_183);
and U310 (N_310,In_467,In_310);
nand U311 (N_311,In_132,In_251);
nor U312 (N_312,In_186,In_301);
and U313 (N_313,In_105,In_24);
or U314 (N_314,In_33,In_425);
and U315 (N_315,In_49,In_138);
and U316 (N_316,In_129,In_208);
or U317 (N_317,In_38,In_80);
and U318 (N_318,In_223,In_314);
and U319 (N_319,In_230,In_69);
or U320 (N_320,In_27,In_466);
nor U321 (N_321,In_410,In_133);
nand U322 (N_322,In_118,In_91);
and U323 (N_323,In_295,In_145);
xnor U324 (N_324,In_270,In_402);
and U325 (N_325,In_361,In_455);
or U326 (N_326,In_424,In_263);
or U327 (N_327,In_306,In_391);
and U328 (N_328,In_167,In_88);
and U329 (N_329,In_437,In_352);
or U330 (N_330,In_436,In_96);
nand U331 (N_331,In_223,In_57);
or U332 (N_332,In_427,In_420);
nand U333 (N_333,In_323,In_415);
nor U334 (N_334,In_492,In_361);
nand U335 (N_335,In_266,In_431);
or U336 (N_336,In_116,In_470);
nand U337 (N_337,In_137,In_361);
nor U338 (N_338,In_191,In_304);
and U339 (N_339,In_153,In_331);
nor U340 (N_340,In_147,In_156);
and U341 (N_341,In_309,In_32);
and U342 (N_342,In_196,In_417);
nand U343 (N_343,In_494,In_300);
or U344 (N_344,In_428,In_499);
and U345 (N_345,In_204,In_11);
or U346 (N_346,In_422,In_156);
nand U347 (N_347,In_237,In_191);
xnor U348 (N_348,In_384,In_465);
or U349 (N_349,In_97,In_329);
xor U350 (N_350,In_164,In_54);
and U351 (N_351,In_324,In_497);
and U352 (N_352,In_315,In_331);
or U353 (N_353,In_231,In_94);
and U354 (N_354,In_109,In_152);
or U355 (N_355,In_238,In_421);
or U356 (N_356,In_372,In_442);
or U357 (N_357,In_388,In_18);
and U358 (N_358,In_206,In_2);
nor U359 (N_359,In_80,In_92);
and U360 (N_360,In_354,In_109);
nand U361 (N_361,In_70,In_291);
and U362 (N_362,In_496,In_332);
or U363 (N_363,In_44,In_123);
and U364 (N_364,In_31,In_495);
nor U365 (N_365,In_174,In_345);
nor U366 (N_366,In_210,In_40);
and U367 (N_367,In_144,In_399);
nor U368 (N_368,In_293,In_499);
and U369 (N_369,In_424,In_98);
or U370 (N_370,In_239,In_94);
or U371 (N_371,In_401,In_317);
or U372 (N_372,In_105,In_88);
or U373 (N_373,In_272,In_141);
and U374 (N_374,In_476,In_9);
or U375 (N_375,In_406,In_213);
nor U376 (N_376,In_392,In_405);
and U377 (N_377,In_124,In_495);
and U378 (N_378,In_259,In_214);
or U379 (N_379,In_389,In_133);
and U380 (N_380,In_122,In_37);
nand U381 (N_381,In_320,In_193);
nor U382 (N_382,In_367,In_443);
nor U383 (N_383,In_228,In_176);
and U384 (N_384,In_454,In_87);
and U385 (N_385,In_310,In_427);
or U386 (N_386,In_494,In_383);
or U387 (N_387,In_139,In_39);
and U388 (N_388,In_301,In_253);
or U389 (N_389,In_6,In_191);
nand U390 (N_390,In_185,In_458);
and U391 (N_391,In_25,In_10);
nand U392 (N_392,In_160,In_190);
nor U393 (N_393,In_17,In_79);
nor U394 (N_394,In_218,In_246);
or U395 (N_395,In_311,In_444);
or U396 (N_396,In_161,In_246);
and U397 (N_397,In_64,In_415);
and U398 (N_398,In_460,In_70);
nand U399 (N_399,In_377,In_48);
nand U400 (N_400,In_222,In_145);
or U401 (N_401,In_221,In_433);
nor U402 (N_402,In_316,In_490);
nor U403 (N_403,In_370,In_177);
nor U404 (N_404,In_20,In_379);
nor U405 (N_405,In_212,In_68);
xor U406 (N_406,In_206,In_367);
nand U407 (N_407,In_408,In_343);
and U408 (N_408,In_208,In_334);
and U409 (N_409,In_143,In_294);
and U410 (N_410,In_280,In_77);
and U411 (N_411,In_278,In_389);
nand U412 (N_412,In_339,In_142);
and U413 (N_413,In_24,In_249);
nand U414 (N_414,In_421,In_412);
or U415 (N_415,In_301,In_267);
nand U416 (N_416,In_269,In_141);
nand U417 (N_417,In_386,In_263);
or U418 (N_418,In_313,In_97);
xor U419 (N_419,In_163,In_257);
nand U420 (N_420,In_496,In_471);
nand U421 (N_421,In_355,In_440);
nor U422 (N_422,In_280,In_250);
or U423 (N_423,In_122,In_422);
nor U424 (N_424,In_336,In_209);
and U425 (N_425,In_223,In_254);
or U426 (N_426,In_45,In_107);
xor U427 (N_427,In_113,In_288);
and U428 (N_428,In_369,In_395);
and U429 (N_429,In_452,In_225);
xnor U430 (N_430,In_382,In_266);
nor U431 (N_431,In_42,In_78);
and U432 (N_432,In_198,In_85);
and U433 (N_433,In_194,In_132);
xor U434 (N_434,In_365,In_324);
nand U435 (N_435,In_312,In_493);
nor U436 (N_436,In_231,In_222);
nand U437 (N_437,In_461,In_189);
nor U438 (N_438,In_407,In_368);
nand U439 (N_439,In_280,In_204);
or U440 (N_440,In_125,In_494);
or U441 (N_441,In_422,In_183);
and U442 (N_442,In_258,In_126);
and U443 (N_443,In_134,In_142);
nand U444 (N_444,In_92,In_7);
xnor U445 (N_445,In_487,In_341);
nor U446 (N_446,In_179,In_427);
nand U447 (N_447,In_342,In_407);
or U448 (N_448,In_320,In_287);
or U449 (N_449,In_203,In_412);
nand U450 (N_450,In_29,In_499);
or U451 (N_451,In_282,In_323);
and U452 (N_452,In_280,In_463);
nor U453 (N_453,In_247,In_256);
nor U454 (N_454,In_485,In_203);
or U455 (N_455,In_409,In_231);
or U456 (N_456,In_254,In_377);
or U457 (N_457,In_50,In_4);
nor U458 (N_458,In_183,In_79);
or U459 (N_459,In_8,In_93);
nor U460 (N_460,In_2,In_155);
nor U461 (N_461,In_409,In_462);
nand U462 (N_462,In_27,In_400);
and U463 (N_463,In_329,In_245);
xor U464 (N_464,In_65,In_122);
nor U465 (N_465,In_134,In_410);
nand U466 (N_466,In_306,In_349);
nor U467 (N_467,In_47,In_392);
nor U468 (N_468,In_254,In_486);
nand U469 (N_469,In_181,In_195);
nor U470 (N_470,In_386,In_423);
and U471 (N_471,In_15,In_87);
or U472 (N_472,In_427,In_86);
and U473 (N_473,In_376,In_273);
nand U474 (N_474,In_29,In_459);
or U475 (N_475,In_326,In_151);
and U476 (N_476,In_48,In_472);
nor U477 (N_477,In_256,In_372);
and U478 (N_478,In_405,In_255);
xor U479 (N_479,In_264,In_134);
and U480 (N_480,In_277,In_473);
or U481 (N_481,In_188,In_446);
and U482 (N_482,In_180,In_128);
nand U483 (N_483,In_50,In_110);
and U484 (N_484,In_94,In_291);
or U485 (N_485,In_137,In_396);
nand U486 (N_486,In_387,In_445);
nand U487 (N_487,In_107,In_455);
or U488 (N_488,In_22,In_176);
and U489 (N_489,In_329,In_58);
nor U490 (N_490,In_202,In_74);
nand U491 (N_491,In_95,In_14);
nand U492 (N_492,In_253,In_350);
nand U493 (N_493,In_257,In_122);
nand U494 (N_494,In_323,In_468);
and U495 (N_495,In_380,In_110);
nand U496 (N_496,In_476,In_429);
nand U497 (N_497,In_234,In_94);
nand U498 (N_498,In_121,In_302);
and U499 (N_499,In_324,In_158);
nand U500 (N_500,N_331,N_340);
or U501 (N_501,N_334,N_82);
nand U502 (N_502,N_227,N_115);
nor U503 (N_503,N_215,N_0);
xor U504 (N_504,N_420,N_299);
or U505 (N_505,N_399,N_353);
nor U506 (N_506,N_377,N_103);
nor U507 (N_507,N_152,N_188);
nand U508 (N_508,N_428,N_43);
nor U509 (N_509,N_276,N_211);
or U510 (N_510,N_277,N_443);
nand U511 (N_511,N_8,N_56);
nand U512 (N_512,N_427,N_327);
nand U513 (N_513,N_436,N_96);
and U514 (N_514,N_167,N_355);
or U515 (N_515,N_16,N_415);
xnor U516 (N_516,N_454,N_243);
nor U517 (N_517,N_136,N_287);
nor U518 (N_518,N_366,N_107);
and U519 (N_519,N_361,N_269);
and U520 (N_520,N_265,N_49);
and U521 (N_521,N_142,N_359);
or U522 (N_522,N_122,N_477);
nand U523 (N_523,N_316,N_230);
nor U524 (N_524,N_134,N_15);
and U525 (N_525,N_404,N_109);
xor U526 (N_526,N_387,N_275);
nand U527 (N_527,N_406,N_348);
and U528 (N_528,N_6,N_455);
nand U529 (N_529,N_68,N_46);
nor U530 (N_530,N_249,N_321);
nor U531 (N_531,N_172,N_129);
nor U532 (N_532,N_384,N_171);
nor U533 (N_533,N_54,N_432);
or U534 (N_534,N_157,N_468);
nor U535 (N_535,N_89,N_294);
and U536 (N_536,N_290,N_281);
nor U537 (N_537,N_449,N_291);
nand U538 (N_538,N_197,N_280);
or U539 (N_539,N_23,N_10);
and U540 (N_540,N_419,N_319);
nand U541 (N_541,N_322,N_424);
and U542 (N_542,N_250,N_228);
nor U543 (N_543,N_124,N_60);
or U544 (N_544,N_199,N_177);
and U545 (N_545,N_206,N_271);
and U546 (N_546,N_37,N_426);
and U547 (N_547,N_195,N_255);
nor U548 (N_548,N_339,N_58);
or U549 (N_549,N_482,N_397);
or U550 (N_550,N_72,N_52);
nor U551 (N_551,N_24,N_492);
xnor U552 (N_552,N_110,N_472);
or U553 (N_553,N_99,N_145);
and U554 (N_554,N_80,N_100);
and U555 (N_555,N_7,N_317);
or U556 (N_556,N_112,N_416);
and U557 (N_557,N_64,N_252);
or U558 (N_558,N_141,N_200);
nand U559 (N_559,N_45,N_13);
nor U560 (N_560,N_184,N_232);
nor U561 (N_561,N_288,N_474);
or U562 (N_562,N_373,N_226);
or U563 (N_563,N_266,N_479);
nor U564 (N_564,N_106,N_370);
or U565 (N_565,N_182,N_5);
nor U566 (N_566,N_241,N_310);
xor U567 (N_567,N_117,N_178);
or U568 (N_568,N_111,N_11);
nand U569 (N_569,N_409,N_450);
or U570 (N_570,N_475,N_459);
nand U571 (N_571,N_304,N_4);
or U572 (N_572,N_238,N_364);
nor U573 (N_573,N_311,N_125);
and U574 (N_574,N_263,N_421);
nor U575 (N_575,N_201,N_388);
and U576 (N_576,N_382,N_254);
or U577 (N_577,N_91,N_491);
nand U578 (N_578,N_191,N_34);
nor U579 (N_579,N_9,N_435);
and U580 (N_580,N_408,N_389);
or U581 (N_581,N_307,N_76);
or U582 (N_582,N_116,N_289);
nor U583 (N_583,N_347,N_351);
nand U584 (N_584,N_374,N_36);
nor U585 (N_585,N_457,N_278);
and U586 (N_586,N_149,N_465);
nand U587 (N_587,N_494,N_485);
and U588 (N_588,N_417,N_140);
or U589 (N_589,N_218,N_22);
and U590 (N_590,N_335,N_297);
xor U591 (N_591,N_356,N_77);
or U592 (N_592,N_371,N_376);
xor U593 (N_593,N_405,N_246);
nand U594 (N_594,N_32,N_248);
nor U595 (N_595,N_27,N_44);
and U596 (N_596,N_495,N_401);
or U597 (N_597,N_101,N_402);
and U598 (N_598,N_239,N_84);
nor U599 (N_599,N_471,N_40);
xnor U600 (N_600,N_413,N_253);
nand U601 (N_601,N_127,N_394);
nand U602 (N_602,N_367,N_194);
nor U603 (N_603,N_189,N_193);
and U604 (N_604,N_393,N_187);
and U605 (N_605,N_490,N_108);
or U606 (N_606,N_126,N_164);
and U607 (N_607,N_221,N_113);
or U608 (N_608,N_293,N_180);
or U609 (N_609,N_323,N_487);
and U610 (N_610,N_222,N_497);
nand U611 (N_611,N_314,N_229);
or U612 (N_612,N_53,N_308);
and U613 (N_613,N_301,N_456);
or U614 (N_614,N_458,N_75);
nand U615 (N_615,N_131,N_363);
or U616 (N_616,N_224,N_20);
nor U617 (N_617,N_441,N_210);
nand U618 (N_618,N_483,N_330);
nand U619 (N_619,N_29,N_85);
nand U620 (N_620,N_79,N_395);
nand U621 (N_621,N_162,N_38);
and U622 (N_622,N_168,N_119);
nand U623 (N_623,N_235,N_65);
nand U624 (N_624,N_242,N_219);
nor U625 (N_625,N_257,N_181);
or U626 (N_626,N_305,N_165);
nor U627 (N_627,N_344,N_360);
or U628 (N_628,N_422,N_453);
or U629 (N_629,N_163,N_260);
and U630 (N_630,N_245,N_480);
and U631 (N_631,N_273,N_154);
or U632 (N_632,N_352,N_220);
and U633 (N_633,N_452,N_247);
nor U634 (N_634,N_442,N_333);
or U635 (N_635,N_212,N_346);
and U636 (N_636,N_489,N_486);
and U637 (N_637,N_258,N_237);
and U638 (N_638,N_496,N_158);
or U639 (N_639,N_190,N_196);
nor U640 (N_640,N_262,N_137);
nand U641 (N_641,N_192,N_41);
or U642 (N_642,N_386,N_223);
nand U643 (N_643,N_161,N_28);
nor U644 (N_644,N_12,N_270);
nor U645 (N_645,N_179,N_92);
nand U646 (N_646,N_14,N_469);
nand U647 (N_647,N_473,N_205);
nand U648 (N_648,N_59,N_274);
nand U649 (N_649,N_286,N_315);
and U650 (N_650,N_71,N_204);
nor U651 (N_651,N_214,N_233);
or U652 (N_652,N_70,N_17);
or U653 (N_653,N_244,N_412);
or U654 (N_654,N_216,N_292);
nand U655 (N_655,N_138,N_375);
nor U656 (N_656,N_95,N_498);
nand U657 (N_657,N_398,N_411);
nor U658 (N_658,N_217,N_396);
nand U659 (N_659,N_381,N_198);
nor U660 (N_660,N_306,N_336);
and U661 (N_661,N_488,N_51);
nor U662 (N_662,N_87,N_121);
nor U663 (N_663,N_337,N_354);
and U664 (N_664,N_251,N_231);
nor U665 (N_665,N_341,N_21);
or U666 (N_666,N_423,N_392);
nand U667 (N_667,N_313,N_185);
nand U668 (N_668,N_57,N_328);
or U669 (N_669,N_114,N_447);
nand U670 (N_670,N_169,N_128);
and U671 (N_671,N_151,N_1);
or U672 (N_672,N_368,N_342);
nor U673 (N_673,N_94,N_362);
nand U674 (N_674,N_439,N_26);
or U675 (N_675,N_176,N_300);
or U676 (N_676,N_343,N_466);
nor U677 (N_677,N_476,N_464);
nand U678 (N_678,N_31,N_2);
nand U679 (N_679,N_470,N_104);
or U680 (N_680,N_30,N_400);
and U681 (N_681,N_50,N_484);
xor U682 (N_682,N_47,N_63);
and U683 (N_683,N_202,N_148);
nor U684 (N_684,N_98,N_448);
nand U685 (N_685,N_160,N_478);
nor U686 (N_686,N_268,N_159);
nand U687 (N_687,N_285,N_207);
or U688 (N_688,N_296,N_378);
nand U689 (N_689,N_430,N_135);
or U690 (N_690,N_120,N_139);
nor U691 (N_691,N_463,N_55);
nor U692 (N_692,N_320,N_295);
and U693 (N_693,N_18,N_358);
nand U694 (N_694,N_379,N_48);
and U695 (N_695,N_166,N_261);
nand U696 (N_696,N_88,N_130);
and U697 (N_697,N_105,N_329);
or U698 (N_698,N_284,N_170);
nand U699 (N_699,N_25,N_19);
or U700 (N_700,N_272,N_410);
nand U701 (N_701,N_345,N_390);
nand U702 (N_702,N_446,N_86);
xnor U703 (N_703,N_81,N_203);
nand U704 (N_704,N_35,N_225);
nor U705 (N_705,N_462,N_467);
nor U706 (N_706,N_282,N_155);
nor U707 (N_707,N_186,N_481);
nand U708 (N_708,N_431,N_460);
or U709 (N_709,N_83,N_62);
nand U710 (N_710,N_302,N_144);
or U711 (N_711,N_434,N_391);
nor U712 (N_712,N_499,N_150);
nand U713 (N_713,N_324,N_326);
xor U714 (N_714,N_259,N_61);
nor U715 (N_715,N_264,N_66);
and U716 (N_716,N_173,N_213);
or U717 (N_717,N_118,N_146);
nand U718 (N_718,N_380,N_153);
and U719 (N_719,N_338,N_383);
nor U720 (N_720,N_208,N_451);
nand U721 (N_721,N_175,N_493);
or U722 (N_722,N_312,N_102);
nor U723 (N_723,N_74,N_461);
and U724 (N_724,N_143,N_433);
and U725 (N_725,N_240,N_349);
and U726 (N_726,N_325,N_318);
xnor U727 (N_727,N_33,N_156);
and U728 (N_728,N_309,N_147);
nand U729 (N_729,N_69,N_418);
xnor U730 (N_730,N_236,N_183);
and U731 (N_731,N_267,N_256);
or U732 (N_732,N_425,N_78);
nand U733 (N_733,N_97,N_67);
nor U734 (N_734,N_283,N_298);
xnor U735 (N_735,N_445,N_73);
nor U736 (N_736,N_279,N_429);
nand U737 (N_737,N_42,N_385);
nand U738 (N_738,N_90,N_209);
nand U739 (N_739,N_234,N_39);
or U740 (N_740,N_414,N_403);
and U741 (N_741,N_133,N_357);
and U742 (N_742,N_369,N_174);
or U743 (N_743,N_3,N_123);
nor U744 (N_744,N_438,N_437);
nand U745 (N_745,N_303,N_365);
nor U746 (N_746,N_350,N_407);
nand U747 (N_747,N_332,N_444);
xor U748 (N_748,N_372,N_440);
nor U749 (N_749,N_132,N_93);
nor U750 (N_750,N_227,N_132);
nand U751 (N_751,N_242,N_13);
nor U752 (N_752,N_113,N_89);
nor U753 (N_753,N_73,N_60);
and U754 (N_754,N_359,N_458);
or U755 (N_755,N_188,N_34);
nand U756 (N_756,N_372,N_215);
and U757 (N_757,N_138,N_226);
nor U758 (N_758,N_237,N_272);
and U759 (N_759,N_354,N_375);
or U760 (N_760,N_169,N_53);
nor U761 (N_761,N_457,N_39);
nand U762 (N_762,N_266,N_493);
or U763 (N_763,N_219,N_473);
nand U764 (N_764,N_450,N_127);
and U765 (N_765,N_434,N_31);
and U766 (N_766,N_329,N_145);
or U767 (N_767,N_435,N_484);
nand U768 (N_768,N_184,N_317);
and U769 (N_769,N_53,N_426);
nand U770 (N_770,N_293,N_54);
nand U771 (N_771,N_307,N_450);
or U772 (N_772,N_478,N_466);
xnor U773 (N_773,N_270,N_195);
or U774 (N_774,N_368,N_495);
and U775 (N_775,N_183,N_454);
or U776 (N_776,N_47,N_445);
nand U777 (N_777,N_215,N_60);
nand U778 (N_778,N_127,N_280);
nor U779 (N_779,N_397,N_105);
nand U780 (N_780,N_434,N_84);
xnor U781 (N_781,N_451,N_108);
nor U782 (N_782,N_386,N_241);
or U783 (N_783,N_321,N_381);
nand U784 (N_784,N_473,N_28);
or U785 (N_785,N_411,N_281);
and U786 (N_786,N_498,N_50);
or U787 (N_787,N_388,N_492);
and U788 (N_788,N_387,N_78);
or U789 (N_789,N_424,N_469);
or U790 (N_790,N_25,N_370);
and U791 (N_791,N_21,N_493);
or U792 (N_792,N_377,N_141);
and U793 (N_793,N_42,N_376);
nor U794 (N_794,N_464,N_167);
and U795 (N_795,N_108,N_420);
and U796 (N_796,N_390,N_244);
or U797 (N_797,N_290,N_85);
nand U798 (N_798,N_389,N_129);
or U799 (N_799,N_137,N_36);
and U800 (N_800,N_3,N_394);
nor U801 (N_801,N_498,N_211);
and U802 (N_802,N_222,N_253);
and U803 (N_803,N_17,N_374);
nand U804 (N_804,N_100,N_257);
or U805 (N_805,N_253,N_232);
nand U806 (N_806,N_446,N_288);
or U807 (N_807,N_178,N_367);
nand U808 (N_808,N_264,N_245);
nor U809 (N_809,N_376,N_106);
or U810 (N_810,N_318,N_303);
nand U811 (N_811,N_99,N_324);
nand U812 (N_812,N_53,N_401);
and U813 (N_813,N_91,N_315);
nor U814 (N_814,N_343,N_235);
or U815 (N_815,N_50,N_305);
and U816 (N_816,N_133,N_88);
nor U817 (N_817,N_434,N_294);
or U818 (N_818,N_27,N_369);
and U819 (N_819,N_476,N_70);
nor U820 (N_820,N_66,N_331);
nor U821 (N_821,N_363,N_7);
nand U822 (N_822,N_432,N_469);
and U823 (N_823,N_161,N_269);
or U824 (N_824,N_218,N_429);
and U825 (N_825,N_292,N_171);
or U826 (N_826,N_249,N_436);
nor U827 (N_827,N_130,N_459);
or U828 (N_828,N_195,N_117);
nor U829 (N_829,N_261,N_490);
nor U830 (N_830,N_471,N_149);
nand U831 (N_831,N_29,N_269);
and U832 (N_832,N_391,N_472);
and U833 (N_833,N_446,N_57);
xor U834 (N_834,N_365,N_44);
xor U835 (N_835,N_304,N_331);
nand U836 (N_836,N_489,N_140);
or U837 (N_837,N_83,N_2);
nand U838 (N_838,N_63,N_187);
and U839 (N_839,N_458,N_101);
nand U840 (N_840,N_69,N_295);
or U841 (N_841,N_55,N_205);
or U842 (N_842,N_172,N_127);
or U843 (N_843,N_383,N_290);
nand U844 (N_844,N_404,N_463);
and U845 (N_845,N_498,N_3);
nor U846 (N_846,N_228,N_7);
nor U847 (N_847,N_59,N_265);
or U848 (N_848,N_314,N_65);
nor U849 (N_849,N_22,N_74);
nor U850 (N_850,N_107,N_329);
and U851 (N_851,N_222,N_232);
nor U852 (N_852,N_112,N_223);
nand U853 (N_853,N_412,N_488);
and U854 (N_854,N_211,N_274);
nor U855 (N_855,N_201,N_104);
nor U856 (N_856,N_19,N_57);
and U857 (N_857,N_246,N_166);
or U858 (N_858,N_453,N_238);
nand U859 (N_859,N_431,N_467);
and U860 (N_860,N_148,N_397);
or U861 (N_861,N_416,N_304);
and U862 (N_862,N_296,N_481);
nand U863 (N_863,N_289,N_383);
nor U864 (N_864,N_4,N_147);
nor U865 (N_865,N_438,N_495);
and U866 (N_866,N_30,N_190);
nand U867 (N_867,N_375,N_262);
nor U868 (N_868,N_21,N_451);
nor U869 (N_869,N_469,N_322);
or U870 (N_870,N_349,N_205);
and U871 (N_871,N_324,N_244);
and U872 (N_872,N_334,N_204);
and U873 (N_873,N_163,N_333);
and U874 (N_874,N_426,N_288);
nor U875 (N_875,N_179,N_427);
nand U876 (N_876,N_240,N_406);
nor U877 (N_877,N_398,N_480);
nor U878 (N_878,N_296,N_204);
or U879 (N_879,N_77,N_160);
or U880 (N_880,N_480,N_445);
or U881 (N_881,N_331,N_116);
nand U882 (N_882,N_134,N_167);
nand U883 (N_883,N_112,N_476);
and U884 (N_884,N_21,N_0);
nand U885 (N_885,N_443,N_418);
xor U886 (N_886,N_289,N_361);
or U887 (N_887,N_82,N_196);
and U888 (N_888,N_387,N_40);
nand U889 (N_889,N_313,N_20);
nand U890 (N_890,N_132,N_144);
nand U891 (N_891,N_459,N_208);
or U892 (N_892,N_108,N_304);
nand U893 (N_893,N_427,N_351);
or U894 (N_894,N_243,N_127);
and U895 (N_895,N_488,N_292);
nor U896 (N_896,N_169,N_208);
nor U897 (N_897,N_317,N_371);
or U898 (N_898,N_407,N_127);
nand U899 (N_899,N_199,N_179);
nand U900 (N_900,N_107,N_307);
nor U901 (N_901,N_31,N_349);
nand U902 (N_902,N_422,N_436);
nor U903 (N_903,N_316,N_253);
and U904 (N_904,N_214,N_364);
nor U905 (N_905,N_87,N_321);
nand U906 (N_906,N_210,N_1);
and U907 (N_907,N_301,N_144);
and U908 (N_908,N_360,N_129);
and U909 (N_909,N_208,N_476);
nand U910 (N_910,N_355,N_221);
nor U911 (N_911,N_104,N_273);
or U912 (N_912,N_180,N_78);
nor U913 (N_913,N_70,N_168);
or U914 (N_914,N_107,N_343);
and U915 (N_915,N_249,N_274);
or U916 (N_916,N_207,N_27);
or U917 (N_917,N_142,N_322);
nor U918 (N_918,N_302,N_325);
and U919 (N_919,N_44,N_130);
or U920 (N_920,N_23,N_205);
and U921 (N_921,N_327,N_205);
nand U922 (N_922,N_414,N_373);
or U923 (N_923,N_332,N_113);
nor U924 (N_924,N_51,N_20);
nor U925 (N_925,N_431,N_64);
xor U926 (N_926,N_45,N_149);
nand U927 (N_927,N_447,N_391);
and U928 (N_928,N_383,N_12);
nand U929 (N_929,N_450,N_257);
or U930 (N_930,N_168,N_126);
and U931 (N_931,N_439,N_2);
or U932 (N_932,N_118,N_86);
nor U933 (N_933,N_91,N_274);
or U934 (N_934,N_96,N_483);
nand U935 (N_935,N_498,N_99);
nand U936 (N_936,N_217,N_283);
nor U937 (N_937,N_151,N_164);
nand U938 (N_938,N_104,N_27);
nand U939 (N_939,N_357,N_104);
and U940 (N_940,N_99,N_184);
and U941 (N_941,N_253,N_385);
and U942 (N_942,N_144,N_163);
or U943 (N_943,N_490,N_237);
and U944 (N_944,N_137,N_376);
nor U945 (N_945,N_122,N_49);
nand U946 (N_946,N_243,N_392);
nor U947 (N_947,N_2,N_430);
nor U948 (N_948,N_218,N_132);
nand U949 (N_949,N_216,N_486);
nor U950 (N_950,N_124,N_450);
nor U951 (N_951,N_292,N_389);
nor U952 (N_952,N_261,N_139);
and U953 (N_953,N_9,N_471);
or U954 (N_954,N_231,N_349);
and U955 (N_955,N_313,N_116);
and U956 (N_956,N_387,N_233);
and U957 (N_957,N_185,N_178);
nor U958 (N_958,N_137,N_322);
nor U959 (N_959,N_2,N_29);
nor U960 (N_960,N_284,N_305);
nand U961 (N_961,N_67,N_493);
nor U962 (N_962,N_398,N_498);
nand U963 (N_963,N_492,N_90);
or U964 (N_964,N_260,N_291);
or U965 (N_965,N_214,N_166);
and U966 (N_966,N_177,N_264);
and U967 (N_967,N_23,N_284);
nand U968 (N_968,N_59,N_473);
or U969 (N_969,N_99,N_354);
nor U970 (N_970,N_76,N_57);
or U971 (N_971,N_271,N_351);
and U972 (N_972,N_359,N_443);
and U973 (N_973,N_242,N_344);
and U974 (N_974,N_472,N_29);
and U975 (N_975,N_431,N_311);
and U976 (N_976,N_204,N_491);
nor U977 (N_977,N_479,N_22);
nand U978 (N_978,N_93,N_222);
or U979 (N_979,N_311,N_14);
nor U980 (N_980,N_370,N_125);
or U981 (N_981,N_227,N_162);
and U982 (N_982,N_251,N_212);
nor U983 (N_983,N_104,N_432);
nand U984 (N_984,N_6,N_8);
and U985 (N_985,N_21,N_178);
and U986 (N_986,N_215,N_2);
and U987 (N_987,N_403,N_142);
nand U988 (N_988,N_428,N_45);
nand U989 (N_989,N_217,N_22);
nor U990 (N_990,N_410,N_439);
or U991 (N_991,N_7,N_343);
and U992 (N_992,N_491,N_245);
and U993 (N_993,N_370,N_203);
nand U994 (N_994,N_393,N_105);
nor U995 (N_995,N_156,N_469);
nor U996 (N_996,N_19,N_199);
and U997 (N_997,N_240,N_455);
nor U998 (N_998,N_64,N_194);
and U999 (N_999,N_17,N_298);
nor U1000 (N_1000,N_781,N_599);
nor U1001 (N_1001,N_880,N_907);
and U1002 (N_1002,N_940,N_856);
and U1003 (N_1003,N_683,N_593);
and U1004 (N_1004,N_580,N_903);
or U1005 (N_1005,N_701,N_978);
nor U1006 (N_1006,N_990,N_804);
nor U1007 (N_1007,N_642,N_959);
nand U1008 (N_1008,N_560,N_971);
or U1009 (N_1009,N_760,N_906);
nor U1010 (N_1010,N_779,N_689);
nand U1011 (N_1011,N_551,N_645);
or U1012 (N_1012,N_525,N_882);
nand U1013 (N_1013,N_658,N_944);
nand U1014 (N_1014,N_711,N_843);
or U1015 (N_1015,N_970,N_867);
nand U1016 (N_1016,N_647,N_974);
or U1017 (N_1017,N_900,N_696);
and U1018 (N_1018,N_932,N_590);
nand U1019 (N_1019,N_628,N_799);
nor U1020 (N_1020,N_646,N_584);
and U1021 (N_1021,N_574,N_730);
nand U1022 (N_1022,N_747,N_668);
and U1023 (N_1023,N_953,N_518);
nor U1024 (N_1024,N_715,N_663);
nor U1025 (N_1025,N_719,N_841);
nor U1026 (N_1026,N_744,N_566);
or U1027 (N_1027,N_594,N_875);
nand U1028 (N_1028,N_596,N_809);
nand U1029 (N_1029,N_772,N_515);
nor U1030 (N_1030,N_775,N_678);
and U1031 (N_1031,N_888,N_697);
nor U1032 (N_1032,N_999,N_676);
nand U1033 (N_1033,N_948,N_890);
and U1034 (N_1034,N_557,N_922);
or U1035 (N_1035,N_579,N_854);
and U1036 (N_1036,N_502,N_756);
or U1037 (N_1037,N_936,N_534);
nor U1038 (N_1038,N_649,N_904);
and U1039 (N_1039,N_549,N_898);
and U1040 (N_1040,N_975,N_636);
and U1041 (N_1041,N_881,N_994);
and U1042 (N_1042,N_825,N_895);
or U1043 (N_1043,N_894,N_535);
xor U1044 (N_1044,N_896,N_694);
or U1045 (N_1045,N_846,N_726);
and U1046 (N_1046,N_553,N_533);
nor U1047 (N_1047,N_988,N_968);
nand U1048 (N_1048,N_769,N_877);
nor U1049 (N_1049,N_759,N_823);
and U1050 (N_1050,N_538,N_790);
or U1051 (N_1051,N_752,N_679);
and U1052 (N_1052,N_749,N_996);
or U1053 (N_1053,N_523,N_659);
xnor U1054 (N_1054,N_556,N_632);
or U1055 (N_1055,N_876,N_864);
nand U1056 (N_1056,N_774,N_615);
and U1057 (N_1057,N_812,N_851);
nand U1058 (N_1058,N_808,N_589);
and U1059 (N_1059,N_861,N_942);
nor U1060 (N_1060,N_688,N_572);
or U1061 (N_1061,N_949,N_662);
nor U1062 (N_1062,N_828,N_567);
nand U1063 (N_1063,N_600,N_609);
and U1064 (N_1064,N_737,N_705);
or U1065 (N_1065,N_935,N_588);
nor U1066 (N_1066,N_723,N_575);
nor U1067 (N_1067,N_690,N_813);
and U1068 (N_1068,N_559,N_914);
nand U1069 (N_1069,N_530,N_651);
and U1070 (N_1070,N_674,N_902);
or U1071 (N_1071,N_699,N_921);
nor U1072 (N_1072,N_728,N_563);
nand U1073 (N_1073,N_717,N_669);
nand U1074 (N_1074,N_827,N_513);
nand U1075 (N_1075,N_789,N_865);
or U1076 (N_1076,N_507,N_576);
nor U1077 (N_1077,N_629,N_810);
and U1078 (N_1078,N_866,N_592);
nand U1079 (N_1079,N_545,N_765);
and U1080 (N_1080,N_795,N_884);
and U1081 (N_1081,N_739,N_562);
nor U1082 (N_1082,N_704,N_550);
and U1083 (N_1083,N_635,N_976);
or U1084 (N_1084,N_686,N_729);
and U1085 (N_1085,N_630,N_623);
nand U1086 (N_1086,N_616,N_956);
and U1087 (N_1087,N_571,N_989);
and U1088 (N_1088,N_660,N_770);
nor U1089 (N_1089,N_505,N_801);
or U1090 (N_1090,N_783,N_621);
and U1091 (N_1091,N_582,N_692);
nand U1092 (N_1092,N_708,N_529);
nand U1093 (N_1093,N_815,N_622);
and U1094 (N_1094,N_703,N_735);
and U1095 (N_1095,N_901,N_691);
nand U1096 (N_1096,N_840,N_657);
nand U1097 (N_1097,N_984,N_987);
nor U1098 (N_1098,N_947,N_754);
or U1099 (N_1099,N_603,N_964);
and U1100 (N_1100,N_541,N_652);
or U1101 (N_1101,N_780,N_638);
or U1102 (N_1102,N_830,N_870);
nand U1103 (N_1103,N_937,N_977);
nand U1104 (N_1104,N_934,N_991);
xor U1105 (N_1105,N_792,N_595);
nor U1106 (N_1106,N_506,N_643);
nor U1107 (N_1107,N_508,N_733);
or U1108 (N_1108,N_913,N_995);
nor U1109 (N_1109,N_569,N_526);
and U1110 (N_1110,N_724,N_552);
nand U1111 (N_1111,N_542,N_540);
or U1112 (N_1112,N_785,N_879);
and U1113 (N_1113,N_546,N_819);
and U1114 (N_1114,N_682,N_793);
xor U1115 (N_1115,N_943,N_834);
nand U1116 (N_1116,N_554,N_547);
or U1117 (N_1117,N_727,N_712);
or U1118 (N_1118,N_811,N_665);
or U1119 (N_1119,N_748,N_555);
xnor U1120 (N_1120,N_655,N_997);
nand U1121 (N_1121,N_814,N_763);
nor U1122 (N_1122,N_982,N_514);
or U1123 (N_1123,N_771,N_802);
and U1124 (N_1124,N_952,N_874);
or U1125 (N_1125,N_998,N_661);
or U1126 (N_1126,N_909,N_720);
nand U1127 (N_1127,N_966,N_577);
nor U1128 (N_1128,N_565,N_503);
nor U1129 (N_1129,N_738,N_761);
nand U1130 (N_1130,N_641,N_803);
or U1131 (N_1131,N_543,N_915);
nand U1132 (N_1132,N_656,N_608);
nor U1133 (N_1133,N_916,N_776);
or U1134 (N_1134,N_905,N_611);
and U1135 (N_1135,N_972,N_923);
or U1136 (N_1136,N_681,N_753);
and U1137 (N_1137,N_672,N_664);
and U1138 (N_1138,N_500,N_601);
and U1139 (N_1139,N_667,N_707);
or U1140 (N_1140,N_796,N_743);
nand U1141 (N_1141,N_787,N_993);
nor U1142 (N_1142,N_741,N_524);
or U1143 (N_1143,N_528,N_564);
nor U1144 (N_1144,N_633,N_631);
nor U1145 (N_1145,N_722,N_951);
or U1146 (N_1146,N_927,N_666);
nand U1147 (N_1147,N_605,N_986);
nand U1148 (N_1148,N_736,N_849);
or U1149 (N_1149,N_887,N_673);
nand U1150 (N_1150,N_831,N_568);
nand U1151 (N_1151,N_857,N_858);
or U1152 (N_1152,N_821,N_710);
nand U1153 (N_1153,N_511,N_919);
nor U1154 (N_1154,N_725,N_677);
and U1155 (N_1155,N_822,N_899);
nand U1156 (N_1156,N_816,N_695);
nand U1157 (N_1157,N_740,N_745);
xnor U1158 (N_1158,N_832,N_624);
nor U1159 (N_1159,N_967,N_750);
nor U1160 (N_1160,N_850,N_732);
or U1161 (N_1161,N_818,N_521);
or U1162 (N_1162,N_981,N_862);
nor U1163 (N_1163,N_602,N_536);
xor U1164 (N_1164,N_805,N_941);
or U1165 (N_1165,N_532,N_924);
nor U1166 (N_1166,N_886,N_908);
nor U1167 (N_1167,N_578,N_680);
or U1168 (N_1168,N_871,N_979);
nor U1169 (N_1169,N_950,N_527);
nand U1170 (N_1170,N_878,N_852);
nand U1171 (N_1171,N_845,N_910);
and U1172 (N_1172,N_892,N_509);
or U1173 (N_1173,N_838,N_925);
or U1174 (N_1174,N_911,N_782);
and U1175 (N_1175,N_519,N_965);
or U1176 (N_1176,N_734,N_639);
and U1177 (N_1177,N_853,N_614);
nand U1178 (N_1178,N_610,N_648);
nor U1179 (N_1179,N_620,N_654);
or U1180 (N_1180,N_847,N_591);
nand U1181 (N_1181,N_872,N_955);
and U1182 (N_1182,N_606,N_824);
and U1183 (N_1183,N_835,N_837);
and U1184 (N_1184,N_912,N_983);
or U1185 (N_1185,N_826,N_859);
nand U1186 (N_1186,N_558,N_992);
and U1187 (N_1187,N_985,N_512);
or U1188 (N_1188,N_746,N_798);
and U1189 (N_1189,N_714,N_762);
or U1190 (N_1190,N_939,N_917);
nor U1191 (N_1191,N_522,N_848);
nor U1192 (N_1192,N_931,N_791);
or U1193 (N_1193,N_946,N_548);
nand U1194 (N_1194,N_625,N_767);
and U1195 (N_1195,N_570,N_731);
nand U1196 (N_1196,N_926,N_501);
nor U1197 (N_1197,N_561,N_531);
nor U1198 (N_1198,N_918,N_597);
xor U1199 (N_1199,N_758,N_929);
or U1200 (N_1200,N_675,N_960);
nor U1201 (N_1201,N_980,N_897);
nor U1202 (N_1202,N_958,N_961);
or U1203 (N_1203,N_751,N_684);
nand U1204 (N_1204,N_963,N_716);
nand U1205 (N_1205,N_670,N_671);
nor U1206 (N_1206,N_516,N_930);
nand U1207 (N_1207,N_957,N_693);
and U1208 (N_1208,N_634,N_585);
xnor U1209 (N_1209,N_653,N_766);
or U1210 (N_1210,N_768,N_784);
nor U1211 (N_1211,N_698,N_598);
and U1212 (N_1212,N_573,N_778);
or U1213 (N_1213,N_860,N_928);
nor U1214 (N_1214,N_721,N_954);
and U1215 (N_1215,N_607,N_626);
nor U1216 (N_1216,N_650,N_842);
nor U1217 (N_1217,N_794,N_869);
nand U1218 (N_1218,N_800,N_604);
and U1219 (N_1219,N_889,N_933);
or U1220 (N_1220,N_713,N_587);
or U1221 (N_1221,N_788,N_855);
nor U1222 (N_1222,N_581,N_510);
and U1223 (N_1223,N_613,N_777);
nand U1224 (N_1224,N_786,N_817);
or U1225 (N_1225,N_644,N_700);
nor U1226 (N_1226,N_973,N_702);
or U1227 (N_1227,N_807,N_504);
nor U1228 (N_1228,N_891,N_839);
or U1229 (N_1229,N_873,N_829);
or U1230 (N_1230,N_583,N_517);
nor U1231 (N_1231,N_640,N_627);
and U1232 (N_1232,N_685,N_544);
or U1233 (N_1233,N_764,N_962);
and U1234 (N_1234,N_969,N_773);
nand U1235 (N_1235,N_806,N_945);
and U1236 (N_1236,N_844,N_687);
and U1237 (N_1237,N_885,N_618);
nand U1238 (N_1238,N_742,N_709);
xnor U1239 (N_1239,N_520,N_863);
nand U1240 (N_1240,N_617,N_797);
or U1241 (N_1241,N_537,N_706);
and U1242 (N_1242,N_539,N_755);
and U1243 (N_1243,N_938,N_820);
and U1244 (N_1244,N_757,N_868);
nand U1245 (N_1245,N_586,N_893);
or U1246 (N_1246,N_920,N_612);
or U1247 (N_1247,N_619,N_836);
and U1248 (N_1248,N_883,N_833);
nand U1249 (N_1249,N_718,N_637);
or U1250 (N_1250,N_594,N_776);
or U1251 (N_1251,N_758,N_578);
xor U1252 (N_1252,N_712,N_917);
nor U1253 (N_1253,N_803,N_907);
nor U1254 (N_1254,N_583,N_655);
nand U1255 (N_1255,N_994,N_766);
nor U1256 (N_1256,N_884,N_867);
or U1257 (N_1257,N_654,N_954);
and U1258 (N_1258,N_805,N_795);
and U1259 (N_1259,N_909,N_661);
nor U1260 (N_1260,N_609,N_591);
nand U1261 (N_1261,N_574,N_719);
or U1262 (N_1262,N_706,N_966);
nand U1263 (N_1263,N_597,N_619);
and U1264 (N_1264,N_971,N_898);
nor U1265 (N_1265,N_729,N_697);
nand U1266 (N_1266,N_885,N_741);
nor U1267 (N_1267,N_659,N_790);
or U1268 (N_1268,N_694,N_712);
and U1269 (N_1269,N_567,N_893);
and U1270 (N_1270,N_916,N_871);
or U1271 (N_1271,N_735,N_588);
nand U1272 (N_1272,N_980,N_753);
nor U1273 (N_1273,N_863,N_918);
nand U1274 (N_1274,N_514,N_925);
nand U1275 (N_1275,N_585,N_954);
nand U1276 (N_1276,N_990,N_933);
or U1277 (N_1277,N_534,N_853);
or U1278 (N_1278,N_788,N_920);
nand U1279 (N_1279,N_554,N_784);
nand U1280 (N_1280,N_971,N_577);
and U1281 (N_1281,N_769,N_674);
nand U1282 (N_1282,N_899,N_645);
or U1283 (N_1283,N_536,N_753);
nor U1284 (N_1284,N_617,N_753);
and U1285 (N_1285,N_994,N_754);
and U1286 (N_1286,N_920,N_663);
and U1287 (N_1287,N_921,N_572);
and U1288 (N_1288,N_700,N_699);
and U1289 (N_1289,N_650,N_776);
nand U1290 (N_1290,N_516,N_555);
and U1291 (N_1291,N_705,N_723);
nand U1292 (N_1292,N_885,N_909);
and U1293 (N_1293,N_923,N_818);
and U1294 (N_1294,N_652,N_703);
xor U1295 (N_1295,N_703,N_824);
nand U1296 (N_1296,N_959,N_569);
and U1297 (N_1297,N_560,N_948);
nor U1298 (N_1298,N_724,N_678);
nor U1299 (N_1299,N_524,N_717);
or U1300 (N_1300,N_559,N_524);
or U1301 (N_1301,N_968,N_830);
and U1302 (N_1302,N_732,N_695);
nand U1303 (N_1303,N_676,N_771);
nor U1304 (N_1304,N_642,N_648);
or U1305 (N_1305,N_941,N_848);
or U1306 (N_1306,N_910,N_867);
nor U1307 (N_1307,N_932,N_956);
nand U1308 (N_1308,N_607,N_563);
or U1309 (N_1309,N_583,N_534);
nor U1310 (N_1310,N_996,N_637);
and U1311 (N_1311,N_626,N_879);
nor U1312 (N_1312,N_813,N_796);
nor U1313 (N_1313,N_678,N_572);
and U1314 (N_1314,N_642,N_575);
and U1315 (N_1315,N_625,N_782);
or U1316 (N_1316,N_861,N_614);
nand U1317 (N_1317,N_805,N_807);
or U1318 (N_1318,N_613,N_650);
or U1319 (N_1319,N_739,N_842);
nand U1320 (N_1320,N_754,N_565);
and U1321 (N_1321,N_869,N_532);
nand U1322 (N_1322,N_505,N_602);
nor U1323 (N_1323,N_693,N_980);
or U1324 (N_1324,N_589,N_937);
or U1325 (N_1325,N_609,N_955);
and U1326 (N_1326,N_616,N_884);
nand U1327 (N_1327,N_797,N_930);
nand U1328 (N_1328,N_808,N_539);
or U1329 (N_1329,N_587,N_922);
or U1330 (N_1330,N_789,N_774);
nor U1331 (N_1331,N_865,N_776);
xnor U1332 (N_1332,N_572,N_743);
nand U1333 (N_1333,N_619,N_821);
and U1334 (N_1334,N_501,N_764);
or U1335 (N_1335,N_786,N_858);
and U1336 (N_1336,N_649,N_884);
or U1337 (N_1337,N_758,N_862);
nand U1338 (N_1338,N_677,N_858);
or U1339 (N_1339,N_881,N_713);
nor U1340 (N_1340,N_574,N_994);
nor U1341 (N_1341,N_801,N_554);
and U1342 (N_1342,N_985,N_940);
or U1343 (N_1343,N_583,N_812);
nand U1344 (N_1344,N_828,N_531);
and U1345 (N_1345,N_578,N_806);
nand U1346 (N_1346,N_620,N_544);
nor U1347 (N_1347,N_516,N_539);
nor U1348 (N_1348,N_561,N_729);
nor U1349 (N_1349,N_945,N_683);
nor U1350 (N_1350,N_989,N_772);
or U1351 (N_1351,N_638,N_994);
and U1352 (N_1352,N_603,N_577);
nand U1353 (N_1353,N_549,N_661);
nand U1354 (N_1354,N_960,N_882);
or U1355 (N_1355,N_942,N_953);
and U1356 (N_1356,N_531,N_932);
nor U1357 (N_1357,N_538,N_641);
and U1358 (N_1358,N_585,N_615);
or U1359 (N_1359,N_796,N_817);
and U1360 (N_1360,N_612,N_895);
nand U1361 (N_1361,N_846,N_965);
nand U1362 (N_1362,N_569,N_631);
nand U1363 (N_1363,N_655,N_560);
and U1364 (N_1364,N_819,N_521);
nor U1365 (N_1365,N_659,N_938);
nor U1366 (N_1366,N_891,N_852);
or U1367 (N_1367,N_762,N_944);
nor U1368 (N_1368,N_821,N_862);
nor U1369 (N_1369,N_755,N_716);
nand U1370 (N_1370,N_963,N_834);
nand U1371 (N_1371,N_524,N_843);
nor U1372 (N_1372,N_909,N_873);
nand U1373 (N_1373,N_538,N_630);
or U1374 (N_1374,N_597,N_797);
and U1375 (N_1375,N_913,N_757);
nor U1376 (N_1376,N_864,N_809);
nand U1377 (N_1377,N_921,N_815);
or U1378 (N_1378,N_766,N_613);
and U1379 (N_1379,N_593,N_971);
nor U1380 (N_1380,N_520,N_842);
and U1381 (N_1381,N_738,N_945);
nor U1382 (N_1382,N_992,N_631);
or U1383 (N_1383,N_826,N_893);
nor U1384 (N_1384,N_985,N_621);
nor U1385 (N_1385,N_802,N_917);
and U1386 (N_1386,N_525,N_715);
or U1387 (N_1387,N_830,N_728);
xor U1388 (N_1388,N_627,N_716);
and U1389 (N_1389,N_924,N_636);
and U1390 (N_1390,N_540,N_965);
nor U1391 (N_1391,N_529,N_660);
nor U1392 (N_1392,N_664,N_711);
and U1393 (N_1393,N_883,N_792);
and U1394 (N_1394,N_996,N_818);
or U1395 (N_1395,N_586,N_799);
nand U1396 (N_1396,N_942,N_827);
xor U1397 (N_1397,N_919,N_529);
and U1398 (N_1398,N_931,N_964);
and U1399 (N_1399,N_931,N_761);
or U1400 (N_1400,N_767,N_623);
nor U1401 (N_1401,N_545,N_950);
nand U1402 (N_1402,N_959,N_660);
or U1403 (N_1403,N_562,N_831);
nor U1404 (N_1404,N_815,N_690);
nand U1405 (N_1405,N_612,N_698);
nor U1406 (N_1406,N_879,N_596);
and U1407 (N_1407,N_738,N_901);
nand U1408 (N_1408,N_992,N_587);
nand U1409 (N_1409,N_690,N_994);
xnor U1410 (N_1410,N_856,N_931);
nand U1411 (N_1411,N_667,N_932);
nor U1412 (N_1412,N_639,N_746);
or U1413 (N_1413,N_585,N_654);
nand U1414 (N_1414,N_603,N_512);
nor U1415 (N_1415,N_808,N_626);
nand U1416 (N_1416,N_896,N_514);
or U1417 (N_1417,N_547,N_765);
nand U1418 (N_1418,N_811,N_509);
and U1419 (N_1419,N_840,N_707);
or U1420 (N_1420,N_503,N_590);
nor U1421 (N_1421,N_812,N_759);
or U1422 (N_1422,N_904,N_838);
and U1423 (N_1423,N_619,N_598);
nor U1424 (N_1424,N_704,N_829);
xnor U1425 (N_1425,N_732,N_968);
and U1426 (N_1426,N_734,N_769);
nand U1427 (N_1427,N_586,N_909);
nor U1428 (N_1428,N_999,N_796);
or U1429 (N_1429,N_908,N_766);
nor U1430 (N_1430,N_840,N_720);
and U1431 (N_1431,N_558,N_589);
nor U1432 (N_1432,N_539,N_920);
nand U1433 (N_1433,N_721,N_661);
and U1434 (N_1434,N_704,N_913);
or U1435 (N_1435,N_729,N_549);
nand U1436 (N_1436,N_508,N_665);
nor U1437 (N_1437,N_755,N_632);
and U1438 (N_1438,N_950,N_564);
or U1439 (N_1439,N_539,N_767);
or U1440 (N_1440,N_805,N_931);
nand U1441 (N_1441,N_644,N_966);
or U1442 (N_1442,N_609,N_930);
and U1443 (N_1443,N_933,N_729);
nand U1444 (N_1444,N_936,N_766);
and U1445 (N_1445,N_764,N_721);
or U1446 (N_1446,N_731,N_999);
and U1447 (N_1447,N_981,N_665);
and U1448 (N_1448,N_669,N_627);
and U1449 (N_1449,N_568,N_727);
nand U1450 (N_1450,N_621,N_778);
nor U1451 (N_1451,N_614,N_785);
nand U1452 (N_1452,N_571,N_815);
nand U1453 (N_1453,N_985,N_967);
and U1454 (N_1454,N_595,N_720);
or U1455 (N_1455,N_514,N_641);
xor U1456 (N_1456,N_503,N_554);
nor U1457 (N_1457,N_950,N_977);
and U1458 (N_1458,N_761,N_746);
nor U1459 (N_1459,N_775,N_614);
and U1460 (N_1460,N_685,N_994);
or U1461 (N_1461,N_519,N_573);
nand U1462 (N_1462,N_627,N_641);
nor U1463 (N_1463,N_910,N_961);
or U1464 (N_1464,N_747,N_623);
nor U1465 (N_1465,N_790,N_713);
or U1466 (N_1466,N_975,N_542);
or U1467 (N_1467,N_869,N_563);
or U1468 (N_1468,N_784,N_723);
nand U1469 (N_1469,N_699,N_572);
and U1470 (N_1470,N_781,N_663);
or U1471 (N_1471,N_721,N_600);
and U1472 (N_1472,N_802,N_873);
nor U1473 (N_1473,N_761,N_708);
nand U1474 (N_1474,N_738,N_633);
or U1475 (N_1475,N_888,N_564);
nand U1476 (N_1476,N_705,N_984);
nand U1477 (N_1477,N_820,N_880);
and U1478 (N_1478,N_595,N_526);
nand U1479 (N_1479,N_846,N_668);
nand U1480 (N_1480,N_608,N_971);
nor U1481 (N_1481,N_651,N_832);
or U1482 (N_1482,N_754,N_681);
nand U1483 (N_1483,N_795,N_543);
nor U1484 (N_1484,N_864,N_916);
or U1485 (N_1485,N_778,N_996);
xnor U1486 (N_1486,N_510,N_634);
nand U1487 (N_1487,N_568,N_613);
nand U1488 (N_1488,N_844,N_619);
nor U1489 (N_1489,N_654,N_625);
and U1490 (N_1490,N_617,N_507);
nand U1491 (N_1491,N_760,N_962);
or U1492 (N_1492,N_686,N_996);
or U1493 (N_1493,N_758,N_884);
and U1494 (N_1494,N_948,N_529);
xor U1495 (N_1495,N_722,N_973);
and U1496 (N_1496,N_517,N_870);
and U1497 (N_1497,N_957,N_937);
and U1498 (N_1498,N_824,N_582);
and U1499 (N_1499,N_528,N_698);
or U1500 (N_1500,N_1295,N_1072);
or U1501 (N_1501,N_1177,N_1008);
and U1502 (N_1502,N_1034,N_1422);
nor U1503 (N_1503,N_1122,N_1420);
and U1504 (N_1504,N_1194,N_1103);
nand U1505 (N_1505,N_1233,N_1038);
nand U1506 (N_1506,N_1151,N_1173);
or U1507 (N_1507,N_1412,N_1240);
and U1508 (N_1508,N_1459,N_1465);
or U1509 (N_1509,N_1478,N_1395);
and U1510 (N_1510,N_1277,N_1332);
nor U1511 (N_1511,N_1148,N_1017);
nand U1512 (N_1512,N_1481,N_1182);
and U1513 (N_1513,N_1153,N_1399);
nand U1514 (N_1514,N_1101,N_1146);
or U1515 (N_1515,N_1162,N_1089);
and U1516 (N_1516,N_1268,N_1102);
and U1517 (N_1517,N_1386,N_1090);
or U1518 (N_1518,N_1473,N_1061);
nor U1519 (N_1519,N_1362,N_1178);
nand U1520 (N_1520,N_1002,N_1293);
or U1521 (N_1521,N_1346,N_1476);
and U1522 (N_1522,N_1470,N_1227);
nor U1523 (N_1523,N_1498,N_1324);
nor U1524 (N_1524,N_1396,N_1036);
xor U1525 (N_1525,N_1201,N_1385);
nand U1526 (N_1526,N_1248,N_1445);
xor U1527 (N_1527,N_1147,N_1000);
nand U1528 (N_1528,N_1064,N_1118);
nand U1529 (N_1529,N_1025,N_1311);
and U1530 (N_1530,N_1126,N_1220);
nor U1531 (N_1531,N_1406,N_1214);
nor U1532 (N_1532,N_1207,N_1373);
nand U1533 (N_1533,N_1022,N_1097);
nand U1534 (N_1534,N_1106,N_1184);
or U1535 (N_1535,N_1360,N_1047);
nand U1536 (N_1536,N_1109,N_1345);
and U1537 (N_1537,N_1342,N_1289);
xor U1538 (N_1538,N_1046,N_1026);
or U1539 (N_1539,N_1461,N_1474);
nor U1540 (N_1540,N_1050,N_1483);
and U1541 (N_1541,N_1125,N_1265);
nor U1542 (N_1542,N_1379,N_1041);
or U1543 (N_1543,N_1204,N_1247);
nand U1544 (N_1544,N_1413,N_1108);
or U1545 (N_1545,N_1161,N_1490);
nor U1546 (N_1546,N_1222,N_1279);
or U1547 (N_1547,N_1016,N_1131);
nor U1548 (N_1548,N_1305,N_1359);
nor U1549 (N_1549,N_1056,N_1155);
or U1550 (N_1550,N_1171,N_1384);
xor U1551 (N_1551,N_1226,N_1331);
nor U1552 (N_1552,N_1377,N_1111);
and U1553 (N_1553,N_1009,N_1033);
nor U1554 (N_1554,N_1258,N_1310);
nor U1555 (N_1555,N_1129,N_1340);
nor U1556 (N_1556,N_1285,N_1313);
nand U1557 (N_1557,N_1048,N_1320);
and U1558 (N_1558,N_1416,N_1011);
nand U1559 (N_1559,N_1397,N_1492);
nand U1560 (N_1560,N_1244,N_1253);
nand U1561 (N_1561,N_1349,N_1426);
nor U1562 (N_1562,N_1128,N_1449);
nor U1563 (N_1563,N_1057,N_1354);
nand U1564 (N_1564,N_1484,N_1007);
and U1565 (N_1565,N_1319,N_1428);
nand U1566 (N_1566,N_1304,N_1032);
and U1567 (N_1567,N_1499,N_1193);
nor U1568 (N_1568,N_1452,N_1356);
nor U1569 (N_1569,N_1215,N_1035);
nor U1570 (N_1570,N_1460,N_1100);
nor U1571 (N_1571,N_1315,N_1479);
nand U1572 (N_1572,N_1180,N_1437);
and U1573 (N_1573,N_1328,N_1183);
nand U1574 (N_1574,N_1443,N_1429);
and U1575 (N_1575,N_1043,N_1040);
or U1576 (N_1576,N_1191,N_1239);
or U1577 (N_1577,N_1343,N_1059);
nand U1578 (N_1578,N_1286,N_1369);
nand U1579 (N_1579,N_1221,N_1276);
or U1580 (N_1580,N_1158,N_1486);
nor U1581 (N_1581,N_1453,N_1387);
and U1582 (N_1582,N_1283,N_1140);
and U1583 (N_1583,N_1317,N_1485);
nand U1584 (N_1584,N_1440,N_1175);
nand U1585 (N_1585,N_1497,N_1080);
nand U1586 (N_1586,N_1230,N_1083);
xnor U1587 (N_1587,N_1023,N_1092);
nand U1588 (N_1588,N_1077,N_1053);
and U1589 (N_1589,N_1348,N_1495);
xnor U1590 (N_1590,N_1307,N_1325);
nand U1591 (N_1591,N_1364,N_1394);
nor U1592 (N_1592,N_1403,N_1401);
or U1593 (N_1593,N_1363,N_1375);
nor U1594 (N_1594,N_1071,N_1219);
or U1595 (N_1595,N_1278,N_1493);
and U1596 (N_1596,N_1120,N_1154);
or U1597 (N_1597,N_1436,N_1149);
or U1598 (N_1598,N_1255,N_1110);
nand U1599 (N_1599,N_1294,N_1361);
or U1600 (N_1600,N_1303,N_1318);
nand U1601 (N_1601,N_1296,N_1257);
nand U1602 (N_1602,N_1438,N_1241);
nor U1603 (N_1603,N_1063,N_1482);
nand U1604 (N_1604,N_1112,N_1351);
or U1605 (N_1605,N_1344,N_1167);
nand U1606 (N_1606,N_1078,N_1085);
and U1607 (N_1607,N_1446,N_1243);
or U1608 (N_1608,N_1271,N_1469);
or U1609 (N_1609,N_1073,N_1068);
or U1610 (N_1610,N_1411,N_1049);
nor U1611 (N_1611,N_1389,N_1280);
or U1612 (N_1612,N_1138,N_1339);
and U1613 (N_1613,N_1462,N_1251);
or U1614 (N_1614,N_1334,N_1388);
nand U1615 (N_1615,N_1245,N_1018);
or U1616 (N_1616,N_1150,N_1358);
nand U1617 (N_1617,N_1455,N_1383);
nor U1618 (N_1618,N_1086,N_1402);
nor U1619 (N_1619,N_1199,N_1019);
nor U1620 (N_1620,N_1076,N_1234);
nand U1621 (N_1621,N_1404,N_1435);
nor U1622 (N_1622,N_1329,N_1269);
and U1623 (N_1623,N_1135,N_1054);
and U1624 (N_1624,N_1454,N_1312);
or U1625 (N_1625,N_1421,N_1231);
and U1626 (N_1626,N_1192,N_1165);
nor U1627 (N_1627,N_1235,N_1205);
nor U1628 (N_1628,N_1288,N_1316);
nand U1629 (N_1629,N_1466,N_1210);
nand U1630 (N_1630,N_1039,N_1355);
nand U1631 (N_1631,N_1274,N_1442);
nor U1632 (N_1632,N_1260,N_1062);
and U1633 (N_1633,N_1143,N_1130);
nor U1634 (N_1634,N_1003,N_1471);
or U1635 (N_1635,N_1489,N_1004);
and U1636 (N_1636,N_1121,N_1353);
and U1637 (N_1637,N_1202,N_1099);
nor U1638 (N_1638,N_1475,N_1393);
nor U1639 (N_1639,N_1432,N_1472);
and U1640 (N_1640,N_1093,N_1189);
or U1641 (N_1641,N_1433,N_1414);
and U1642 (N_1642,N_1374,N_1390);
or U1643 (N_1643,N_1213,N_1211);
or U1644 (N_1644,N_1250,N_1232);
nand U1645 (N_1645,N_1263,N_1037);
nor U1646 (N_1646,N_1190,N_1238);
nor U1647 (N_1647,N_1308,N_1378);
and U1648 (N_1648,N_1156,N_1176);
nand U1649 (N_1649,N_1246,N_1081);
nand U1650 (N_1650,N_1115,N_1463);
nand U1651 (N_1651,N_1309,N_1292);
nor U1652 (N_1652,N_1336,N_1398);
and U1653 (N_1653,N_1427,N_1267);
nor U1654 (N_1654,N_1335,N_1030);
nand U1655 (N_1655,N_1074,N_1141);
and U1656 (N_1656,N_1287,N_1005);
nor U1657 (N_1657,N_1487,N_1382);
and U1658 (N_1658,N_1347,N_1249);
nor U1659 (N_1659,N_1082,N_1418);
or U1660 (N_1660,N_1366,N_1488);
and U1661 (N_1661,N_1188,N_1075);
or U1662 (N_1662,N_1290,N_1006);
and U1663 (N_1663,N_1291,N_1114);
nor U1664 (N_1664,N_1259,N_1262);
or U1665 (N_1665,N_1273,N_1477);
nor U1666 (N_1666,N_1372,N_1001);
or U1667 (N_1667,N_1237,N_1113);
nand U1668 (N_1668,N_1323,N_1203);
and U1669 (N_1669,N_1337,N_1104);
nand U1670 (N_1670,N_1069,N_1163);
nand U1671 (N_1671,N_1098,N_1272);
and U1672 (N_1672,N_1058,N_1242);
and U1673 (N_1673,N_1208,N_1236);
and U1674 (N_1674,N_1144,N_1254);
nand U1675 (N_1675,N_1468,N_1430);
nand U1676 (N_1676,N_1451,N_1370);
or U1677 (N_1677,N_1051,N_1195);
nand U1678 (N_1678,N_1169,N_1480);
or U1679 (N_1679,N_1060,N_1217);
nand U1680 (N_1680,N_1168,N_1256);
nor U1681 (N_1681,N_1124,N_1132);
or U1682 (N_1682,N_1070,N_1179);
or U1683 (N_1683,N_1300,N_1264);
or U1684 (N_1684,N_1170,N_1014);
nor U1685 (N_1685,N_1371,N_1134);
nor U1686 (N_1686,N_1333,N_1496);
nand U1687 (N_1687,N_1145,N_1447);
xor U1688 (N_1688,N_1434,N_1270);
and U1689 (N_1689,N_1096,N_1065);
or U1690 (N_1690,N_1365,N_1261);
and U1691 (N_1691,N_1327,N_1407);
and U1692 (N_1692,N_1298,N_1450);
nor U1693 (N_1693,N_1028,N_1095);
or U1694 (N_1694,N_1456,N_1314);
or U1695 (N_1695,N_1172,N_1027);
or U1696 (N_1696,N_1087,N_1448);
and U1697 (N_1697,N_1229,N_1417);
nor U1698 (N_1698,N_1088,N_1031);
nor U1699 (N_1699,N_1218,N_1423);
nor U1700 (N_1700,N_1458,N_1431);
xnor U1701 (N_1701,N_1223,N_1367);
nor U1702 (N_1702,N_1187,N_1302);
nor U1703 (N_1703,N_1392,N_1159);
nor U1704 (N_1704,N_1196,N_1094);
and U1705 (N_1705,N_1198,N_1044);
or U1706 (N_1706,N_1326,N_1301);
nor U1707 (N_1707,N_1136,N_1225);
nor U1708 (N_1708,N_1186,N_1441);
and U1709 (N_1709,N_1029,N_1457);
nand U1710 (N_1710,N_1067,N_1400);
or U1711 (N_1711,N_1127,N_1408);
nand U1712 (N_1712,N_1012,N_1055);
or U1713 (N_1713,N_1381,N_1152);
and U1714 (N_1714,N_1042,N_1425);
or U1715 (N_1715,N_1424,N_1020);
and U1716 (N_1716,N_1282,N_1297);
nor U1717 (N_1717,N_1010,N_1133);
nor U1718 (N_1718,N_1185,N_1091);
or U1719 (N_1719,N_1107,N_1224);
nor U1720 (N_1720,N_1321,N_1015);
and U1721 (N_1721,N_1174,N_1380);
or U1722 (N_1722,N_1341,N_1252);
nor U1723 (N_1723,N_1299,N_1052);
or U1724 (N_1724,N_1024,N_1228);
nand U1725 (N_1725,N_1200,N_1119);
nor U1726 (N_1726,N_1350,N_1181);
and U1727 (N_1727,N_1197,N_1021);
nand U1728 (N_1728,N_1439,N_1157);
nand U1729 (N_1729,N_1444,N_1117);
xor U1730 (N_1730,N_1066,N_1352);
or U1731 (N_1731,N_1045,N_1281);
and U1732 (N_1732,N_1275,N_1216);
nor U1733 (N_1733,N_1409,N_1306);
nor U1734 (N_1734,N_1419,N_1137);
or U1735 (N_1735,N_1105,N_1116);
or U1736 (N_1736,N_1467,N_1266);
and U1737 (N_1737,N_1322,N_1166);
nand U1738 (N_1738,N_1376,N_1284);
nand U1739 (N_1739,N_1464,N_1209);
or U1740 (N_1740,N_1123,N_1494);
or U1741 (N_1741,N_1212,N_1084);
and U1742 (N_1742,N_1330,N_1357);
nand U1743 (N_1743,N_1160,N_1338);
and U1744 (N_1744,N_1491,N_1206);
and U1745 (N_1745,N_1142,N_1410);
or U1746 (N_1746,N_1415,N_1164);
nand U1747 (N_1747,N_1079,N_1013);
or U1748 (N_1748,N_1405,N_1139);
nor U1749 (N_1749,N_1368,N_1391);
nor U1750 (N_1750,N_1248,N_1300);
nor U1751 (N_1751,N_1010,N_1407);
xnor U1752 (N_1752,N_1142,N_1317);
or U1753 (N_1753,N_1441,N_1294);
and U1754 (N_1754,N_1368,N_1327);
nand U1755 (N_1755,N_1376,N_1161);
or U1756 (N_1756,N_1307,N_1243);
and U1757 (N_1757,N_1097,N_1327);
or U1758 (N_1758,N_1171,N_1066);
nor U1759 (N_1759,N_1123,N_1409);
and U1760 (N_1760,N_1114,N_1223);
nand U1761 (N_1761,N_1127,N_1486);
and U1762 (N_1762,N_1003,N_1393);
and U1763 (N_1763,N_1081,N_1015);
nand U1764 (N_1764,N_1278,N_1091);
or U1765 (N_1765,N_1402,N_1459);
and U1766 (N_1766,N_1232,N_1242);
nor U1767 (N_1767,N_1112,N_1404);
nand U1768 (N_1768,N_1154,N_1015);
nand U1769 (N_1769,N_1227,N_1193);
nor U1770 (N_1770,N_1464,N_1120);
nor U1771 (N_1771,N_1083,N_1336);
nand U1772 (N_1772,N_1372,N_1380);
nand U1773 (N_1773,N_1479,N_1179);
nand U1774 (N_1774,N_1435,N_1392);
nor U1775 (N_1775,N_1063,N_1070);
nor U1776 (N_1776,N_1041,N_1236);
nor U1777 (N_1777,N_1138,N_1378);
nor U1778 (N_1778,N_1280,N_1039);
nor U1779 (N_1779,N_1267,N_1121);
or U1780 (N_1780,N_1061,N_1188);
nor U1781 (N_1781,N_1148,N_1456);
or U1782 (N_1782,N_1355,N_1152);
and U1783 (N_1783,N_1412,N_1107);
and U1784 (N_1784,N_1106,N_1111);
nand U1785 (N_1785,N_1211,N_1391);
nor U1786 (N_1786,N_1398,N_1420);
nor U1787 (N_1787,N_1484,N_1457);
and U1788 (N_1788,N_1133,N_1258);
or U1789 (N_1789,N_1073,N_1129);
nand U1790 (N_1790,N_1180,N_1345);
nand U1791 (N_1791,N_1081,N_1053);
and U1792 (N_1792,N_1187,N_1455);
nand U1793 (N_1793,N_1114,N_1441);
and U1794 (N_1794,N_1074,N_1010);
or U1795 (N_1795,N_1071,N_1307);
or U1796 (N_1796,N_1163,N_1150);
nor U1797 (N_1797,N_1274,N_1392);
nor U1798 (N_1798,N_1224,N_1346);
or U1799 (N_1799,N_1029,N_1313);
nor U1800 (N_1800,N_1066,N_1114);
nand U1801 (N_1801,N_1095,N_1020);
nand U1802 (N_1802,N_1209,N_1093);
or U1803 (N_1803,N_1089,N_1178);
and U1804 (N_1804,N_1007,N_1319);
and U1805 (N_1805,N_1353,N_1096);
or U1806 (N_1806,N_1021,N_1422);
or U1807 (N_1807,N_1081,N_1236);
or U1808 (N_1808,N_1456,N_1484);
and U1809 (N_1809,N_1058,N_1248);
nor U1810 (N_1810,N_1047,N_1019);
nor U1811 (N_1811,N_1257,N_1073);
nor U1812 (N_1812,N_1314,N_1278);
nand U1813 (N_1813,N_1210,N_1198);
and U1814 (N_1814,N_1085,N_1426);
nand U1815 (N_1815,N_1327,N_1487);
or U1816 (N_1816,N_1133,N_1354);
or U1817 (N_1817,N_1232,N_1170);
nor U1818 (N_1818,N_1236,N_1426);
nand U1819 (N_1819,N_1291,N_1264);
nor U1820 (N_1820,N_1383,N_1227);
nand U1821 (N_1821,N_1488,N_1017);
and U1822 (N_1822,N_1295,N_1110);
or U1823 (N_1823,N_1037,N_1067);
or U1824 (N_1824,N_1151,N_1385);
nand U1825 (N_1825,N_1034,N_1379);
or U1826 (N_1826,N_1475,N_1470);
nor U1827 (N_1827,N_1307,N_1214);
and U1828 (N_1828,N_1376,N_1438);
and U1829 (N_1829,N_1482,N_1311);
or U1830 (N_1830,N_1285,N_1494);
or U1831 (N_1831,N_1401,N_1272);
and U1832 (N_1832,N_1203,N_1141);
or U1833 (N_1833,N_1496,N_1403);
or U1834 (N_1834,N_1187,N_1183);
or U1835 (N_1835,N_1291,N_1394);
nor U1836 (N_1836,N_1012,N_1140);
and U1837 (N_1837,N_1176,N_1059);
nor U1838 (N_1838,N_1379,N_1209);
and U1839 (N_1839,N_1017,N_1437);
nor U1840 (N_1840,N_1380,N_1359);
nand U1841 (N_1841,N_1477,N_1224);
nor U1842 (N_1842,N_1146,N_1302);
nand U1843 (N_1843,N_1150,N_1290);
and U1844 (N_1844,N_1181,N_1150);
or U1845 (N_1845,N_1297,N_1195);
or U1846 (N_1846,N_1466,N_1228);
and U1847 (N_1847,N_1289,N_1058);
nor U1848 (N_1848,N_1302,N_1216);
nand U1849 (N_1849,N_1446,N_1463);
or U1850 (N_1850,N_1303,N_1179);
and U1851 (N_1851,N_1166,N_1048);
or U1852 (N_1852,N_1185,N_1249);
nor U1853 (N_1853,N_1129,N_1462);
xnor U1854 (N_1854,N_1236,N_1401);
or U1855 (N_1855,N_1300,N_1058);
or U1856 (N_1856,N_1296,N_1474);
nor U1857 (N_1857,N_1092,N_1114);
nand U1858 (N_1858,N_1158,N_1220);
nand U1859 (N_1859,N_1448,N_1195);
xor U1860 (N_1860,N_1290,N_1037);
nor U1861 (N_1861,N_1358,N_1221);
or U1862 (N_1862,N_1442,N_1348);
nor U1863 (N_1863,N_1397,N_1214);
or U1864 (N_1864,N_1316,N_1319);
and U1865 (N_1865,N_1018,N_1037);
and U1866 (N_1866,N_1404,N_1092);
and U1867 (N_1867,N_1376,N_1107);
or U1868 (N_1868,N_1195,N_1214);
nor U1869 (N_1869,N_1338,N_1389);
nand U1870 (N_1870,N_1407,N_1321);
nand U1871 (N_1871,N_1242,N_1342);
or U1872 (N_1872,N_1325,N_1036);
and U1873 (N_1873,N_1458,N_1317);
nand U1874 (N_1874,N_1270,N_1308);
nor U1875 (N_1875,N_1463,N_1195);
or U1876 (N_1876,N_1224,N_1184);
nand U1877 (N_1877,N_1062,N_1071);
and U1878 (N_1878,N_1275,N_1494);
nor U1879 (N_1879,N_1240,N_1062);
and U1880 (N_1880,N_1112,N_1345);
or U1881 (N_1881,N_1316,N_1248);
or U1882 (N_1882,N_1348,N_1049);
xor U1883 (N_1883,N_1028,N_1090);
nor U1884 (N_1884,N_1171,N_1183);
nor U1885 (N_1885,N_1132,N_1196);
or U1886 (N_1886,N_1121,N_1406);
or U1887 (N_1887,N_1377,N_1044);
and U1888 (N_1888,N_1368,N_1264);
nor U1889 (N_1889,N_1324,N_1089);
or U1890 (N_1890,N_1377,N_1048);
and U1891 (N_1891,N_1291,N_1414);
and U1892 (N_1892,N_1449,N_1237);
and U1893 (N_1893,N_1316,N_1171);
nor U1894 (N_1894,N_1040,N_1014);
or U1895 (N_1895,N_1280,N_1453);
and U1896 (N_1896,N_1260,N_1076);
and U1897 (N_1897,N_1303,N_1171);
nor U1898 (N_1898,N_1043,N_1251);
nor U1899 (N_1899,N_1322,N_1494);
and U1900 (N_1900,N_1294,N_1050);
and U1901 (N_1901,N_1274,N_1086);
nor U1902 (N_1902,N_1381,N_1204);
or U1903 (N_1903,N_1163,N_1215);
xnor U1904 (N_1904,N_1415,N_1170);
nor U1905 (N_1905,N_1053,N_1496);
and U1906 (N_1906,N_1337,N_1451);
nand U1907 (N_1907,N_1426,N_1481);
or U1908 (N_1908,N_1032,N_1355);
nor U1909 (N_1909,N_1314,N_1174);
nor U1910 (N_1910,N_1406,N_1023);
nor U1911 (N_1911,N_1088,N_1363);
and U1912 (N_1912,N_1449,N_1058);
or U1913 (N_1913,N_1022,N_1440);
nor U1914 (N_1914,N_1357,N_1153);
nor U1915 (N_1915,N_1190,N_1021);
nand U1916 (N_1916,N_1485,N_1073);
xor U1917 (N_1917,N_1249,N_1245);
nor U1918 (N_1918,N_1236,N_1398);
or U1919 (N_1919,N_1127,N_1041);
and U1920 (N_1920,N_1100,N_1459);
xnor U1921 (N_1921,N_1458,N_1291);
and U1922 (N_1922,N_1155,N_1423);
nor U1923 (N_1923,N_1383,N_1054);
nand U1924 (N_1924,N_1233,N_1163);
xnor U1925 (N_1925,N_1415,N_1392);
nand U1926 (N_1926,N_1151,N_1061);
or U1927 (N_1927,N_1351,N_1449);
nand U1928 (N_1928,N_1135,N_1225);
nor U1929 (N_1929,N_1082,N_1307);
and U1930 (N_1930,N_1165,N_1353);
nor U1931 (N_1931,N_1163,N_1266);
or U1932 (N_1932,N_1321,N_1167);
nand U1933 (N_1933,N_1260,N_1353);
or U1934 (N_1934,N_1157,N_1469);
nor U1935 (N_1935,N_1401,N_1182);
nor U1936 (N_1936,N_1234,N_1364);
nand U1937 (N_1937,N_1079,N_1413);
and U1938 (N_1938,N_1324,N_1242);
and U1939 (N_1939,N_1113,N_1172);
nand U1940 (N_1940,N_1213,N_1311);
or U1941 (N_1941,N_1425,N_1165);
nand U1942 (N_1942,N_1385,N_1081);
nand U1943 (N_1943,N_1287,N_1039);
nand U1944 (N_1944,N_1306,N_1131);
and U1945 (N_1945,N_1000,N_1376);
nand U1946 (N_1946,N_1266,N_1476);
or U1947 (N_1947,N_1323,N_1224);
nor U1948 (N_1948,N_1452,N_1257);
or U1949 (N_1949,N_1301,N_1121);
nand U1950 (N_1950,N_1293,N_1306);
and U1951 (N_1951,N_1132,N_1053);
or U1952 (N_1952,N_1238,N_1342);
and U1953 (N_1953,N_1205,N_1029);
and U1954 (N_1954,N_1484,N_1378);
and U1955 (N_1955,N_1003,N_1497);
and U1956 (N_1956,N_1163,N_1433);
nor U1957 (N_1957,N_1281,N_1193);
nor U1958 (N_1958,N_1256,N_1290);
nor U1959 (N_1959,N_1467,N_1443);
nand U1960 (N_1960,N_1001,N_1065);
nand U1961 (N_1961,N_1455,N_1416);
nand U1962 (N_1962,N_1359,N_1107);
or U1963 (N_1963,N_1030,N_1264);
and U1964 (N_1964,N_1171,N_1425);
nand U1965 (N_1965,N_1326,N_1207);
nor U1966 (N_1966,N_1057,N_1399);
and U1967 (N_1967,N_1005,N_1075);
nor U1968 (N_1968,N_1342,N_1356);
nor U1969 (N_1969,N_1104,N_1256);
and U1970 (N_1970,N_1203,N_1068);
nor U1971 (N_1971,N_1011,N_1241);
or U1972 (N_1972,N_1268,N_1206);
or U1973 (N_1973,N_1025,N_1068);
and U1974 (N_1974,N_1034,N_1145);
nand U1975 (N_1975,N_1473,N_1269);
and U1976 (N_1976,N_1410,N_1388);
or U1977 (N_1977,N_1382,N_1381);
or U1978 (N_1978,N_1095,N_1449);
or U1979 (N_1979,N_1108,N_1383);
nand U1980 (N_1980,N_1006,N_1166);
nand U1981 (N_1981,N_1415,N_1372);
or U1982 (N_1982,N_1082,N_1028);
nand U1983 (N_1983,N_1490,N_1198);
and U1984 (N_1984,N_1030,N_1180);
nand U1985 (N_1985,N_1084,N_1444);
and U1986 (N_1986,N_1263,N_1246);
nand U1987 (N_1987,N_1127,N_1411);
or U1988 (N_1988,N_1112,N_1360);
nand U1989 (N_1989,N_1047,N_1379);
nand U1990 (N_1990,N_1385,N_1491);
and U1991 (N_1991,N_1428,N_1004);
or U1992 (N_1992,N_1439,N_1396);
and U1993 (N_1993,N_1064,N_1407);
and U1994 (N_1994,N_1259,N_1417);
or U1995 (N_1995,N_1032,N_1305);
or U1996 (N_1996,N_1332,N_1134);
nor U1997 (N_1997,N_1215,N_1451);
nand U1998 (N_1998,N_1078,N_1327);
or U1999 (N_1999,N_1017,N_1416);
nand U2000 (N_2000,N_1951,N_1925);
or U2001 (N_2001,N_1840,N_1740);
xor U2002 (N_2002,N_1723,N_1659);
nand U2003 (N_2003,N_1743,N_1835);
xnor U2004 (N_2004,N_1790,N_1749);
and U2005 (N_2005,N_1858,N_1941);
or U2006 (N_2006,N_1530,N_1898);
or U2007 (N_2007,N_1515,N_1847);
or U2008 (N_2008,N_1757,N_1953);
or U2009 (N_2009,N_1714,N_1682);
and U2010 (N_2010,N_1828,N_1514);
xnor U2011 (N_2011,N_1764,N_1708);
xor U2012 (N_2012,N_1785,N_1725);
and U2013 (N_2013,N_1859,N_1888);
nor U2014 (N_2014,N_1756,N_1526);
nand U2015 (N_2015,N_1961,N_1942);
and U2016 (N_2016,N_1831,N_1967);
and U2017 (N_2017,N_1510,N_1674);
or U2018 (N_2018,N_1626,N_1860);
or U2019 (N_2019,N_1927,N_1545);
and U2020 (N_2020,N_1878,N_1923);
and U2021 (N_2021,N_1706,N_1633);
xnor U2022 (N_2022,N_1766,N_1973);
nand U2023 (N_2023,N_1807,N_1728);
and U2024 (N_2024,N_1541,N_1734);
nor U2025 (N_2025,N_1738,N_1853);
nand U2026 (N_2026,N_1901,N_1652);
nand U2027 (N_2027,N_1508,N_1623);
nor U2028 (N_2028,N_1534,N_1803);
and U2029 (N_2029,N_1993,N_1575);
or U2030 (N_2030,N_1727,N_1819);
nand U2031 (N_2031,N_1531,N_1643);
nor U2032 (N_2032,N_1730,N_1569);
and U2033 (N_2033,N_1665,N_1809);
nand U2034 (N_2034,N_1795,N_1874);
nand U2035 (N_2035,N_1722,N_1978);
nand U2036 (N_2036,N_1981,N_1532);
nand U2037 (N_2037,N_1673,N_1671);
and U2038 (N_2038,N_1509,N_1876);
and U2039 (N_2039,N_1637,N_1754);
nand U2040 (N_2040,N_1767,N_1871);
nand U2041 (N_2041,N_1994,N_1924);
nor U2042 (N_2042,N_1592,N_1873);
or U2043 (N_2043,N_1815,N_1947);
nor U2044 (N_2044,N_1695,N_1669);
or U2045 (N_2045,N_1755,N_1829);
nand U2046 (N_2046,N_1857,N_1559);
nor U2047 (N_2047,N_1564,N_1917);
xor U2048 (N_2048,N_1940,N_1655);
or U2049 (N_2049,N_1833,N_1500);
nor U2050 (N_2050,N_1550,N_1970);
and U2051 (N_2051,N_1957,N_1883);
or U2052 (N_2052,N_1679,N_1590);
or U2053 (N_2053,N_1784,N_1931);
nor U2054 (N_2054,N_1991,N_1612);
nand U2055 (N_2055,N_1576,N_1890);
and U2056 (N_2056,N_1960,N_1557);
nor U2057 (N_2057,N_1697,N_1919);
nand U2058 (N_2058,N_1748,N_1701);
or U2059 (N_2059,N_1689,N_1782);
or U2060 (N_2060,N_1816,N_1971);
nor U2061 (N_2061,N_1818,N_1913);
nand U2062 (N_2062,N_1989,N_1851);
or U2063 (N_2063,N_1928,N_1711);
and U2064 (N_2064,N_1737,N_1963);
and U2065 (N_2065,N_1794,N_1584);
nand U2066 (N_2066,N_1600,N_1547);
or U2067 (N_2067,N_1583,N_1826);
nand U2068 (N_2068,N_1911,N_1769);
and U2069 (N_2069,N_1724,N_1691);
nor U2070 (N_2070,N_1909,N_1745);
nand U2071 (N_2071,N_1624,N_1812);
nor U2072 (N_2072,N_1715,N_1506);
and U2073 (N_2073,N_1915,N_1990);
nor U2074 (N_2074,N_1558,N_1548);
and U2075 (N_2075,N_1863,N_1955);
and U2076 (N_2076,N_1642,N_1774);
or U2077 (N_2077,N_1739,N_1634);
nand U2078 (N_2078,N_1950,N_1735);
and U2079 (N_2079,N_1975,N_1553);
nor U2080 (N_2080,N_1908,N_1627);
nor U2081 (N_2081,N_1638,N_1586);
nor U2082 (N_2082,N_1597,N_1690);
nor U2083 (N_2083,N_1983,N_1882);
nand U2084 (N_2084,N_1503,N_1716);
nor U2085 (N_2085,N_1629,N_1646);
and U2086 (N_2086,N_1688,N_1854);
nor U2087 (N_2087,N_1992,N_1881);
nand U2088 (N_2088,N_1662,N_1587);
nand U2089 (N_2089,N_1588,N_1800);
or U2090 (N_2090,N_1952,N_1733);
or U2091 (N_2091,N_1704,N_1647);
and U2092 (N_2092,N_1964,N_1920);
nor U2093 (N_2093,N_1772,N_1799);
or U2094 (N_2094,N_1912,N_1841);
nand U2095 (N_2095,N_1804,N_1793);
nand U2096 (N_2096,N_1930,N_1958);
or U2097 (N_2097,N_1683,N_1519);
and U2098 (N_2098,N_1520,N_1618);
xor U2099 (N_2099,N_1698,N_1666);
or U2100 (N_2100,N_1864,N_1788);
and U2101 (N_2101,N_1904,N_1792);
or U2102 (N_2102,N_1705,N_1591);
nor U2103 (N_2103,N_1773,N_1949);
nand U2104 (N_2104,N_1645,N_1877);
nand U2105 (N_2105,N_1677,N_1731);
nand U2106 (N_2106,N_1806,N_1846);
or U2107 (N_2107,N_1893,N_1903);
and U2108 (N_2108,N_1744,N_1501);
nand U2109 (N_2109,N_1729,N_1937);
nor U2110 (N_2110,N_1533,N_1850);
or U2111 (N_2111,N_1896,N_1721);
nand U2112 (N_2112,N_1502,N_1566);
nor U2113 (N_2113,N_1517,N_1599);
nand U2114 (N_2114,N_1929,N_1867);
nor U2115 (N_2115,N_1985,N_1632);
nor U2116 (N_2116,N_1573,N_1692);
or U2117 (N_2117,N_1540,N_1649);
and U2118 (N_2118,N_1598,N_1855);
and U2119 (N_2119,N_1604,N_1563);
nor U2120 (N_2120,N_1605,N_1570);
or U2121 (N_2121,N_1603,N_1822);
and U2122 (N_2122,N_1763,N_1658);
or U2123 (N_2123,N_1551,N_1768);
nand U2124 (N_2124,N_1751,N_1617);
and U2125 (N_2125,N_1752,N_1988);
or U2126 (N_2126,N_1577,N_1965);
nor U2127 (N_2127,N_1518,N_1758);
nor U2128 (N_2128,N_1918,N_1676);
xnor U2129 (N_2129,N_1562,N_1717);
or U2130 (N_2130,N_1808,N_1943);
nand U2131 (N_2131,N_1589,N_1552);
nor U2132 (N_2132,N_1567,N_1650);
nor U2133 (N_2133,N_1885,N_1895);
xnor U2134 (N_2134,N_1686,N_1865);
nor U2135 (N_2135,N_1891,N_1775);
or U2136 (N_2136,N_1777,N_1596);
nor U2137 (N_2137,N_1856,N_1844);
or U2138 (N_2138,N_1644,N_1842);
xnor U2139 (N_2139,N_1922,N_1839);
nor U2140 (N_2140,N_1933,N_1787);
or U2141 (N_2141,N_1999,N_1830);
nor U2142 (N_2142,N_1838,N_1977);
and U2143 (N_2143,N_1998,N_1672);
xor U2144 (N_2144,N_1611,N_1972);
nand U2145 (N_2145,N_1578,N_1700);
nand U2146 (N_2146,N_1636,N_1779);
nor U2147 (N_2147,N_1640,N_1580);
and U2148 (N_2148,N_1535,N_1762);
nor U2149 (N_2149,N_1761,N_1974);
nand U2150 (N_2150,N_1810,N_1709);
and U2151 (N_2151,N_1944,N_1561);
nor U2152 (N_2152,N_1668,N_1742);
nand U2153 (N_2153,N_1870,N_1910);
nand U2154 (N_2154,N_1710,N_1529);
nand U2155 (N_2155,N_1796,N_1980);
and U2156 (N_2156,N_1581,N_1505);
and U2157 (N_2157,N_1760,N_1987);
or U2158 (N_2158,N_1837,N_1568);
and U2159 (N_2159,N_1525,N_1619);
xnor U2160 (N_2160,N_1820,N_1954);
nor U2161 (N_2161,N_1979,N_1556);
and U2162 (N_2162,N_1694,N_1622);
xor U2163 (N_2163,N_1783,N_1513);
nor U2164 (N_2164,N_1906,N_1916);
and U2165 (N_2165,N_1511,N_1696);
or U2166 (N_2166,N_1607,N_1608);
or U2167 (N_2167,N_1834,N_1832);
or U2168 (N_2168,N_1641,N_1613);
nand U2169 (N_2169,N_1574,N_1778);
nand U2170 (N_2170,N_1719,N_1902);
or U2171 (N_2171,N_1681,N_1825);
nor U2172 (N_2172,N_1921,N_1610);
and U2173 (N_2173,N_1811,N_1889);
nand U2174 (N_2174,N_1544,N_1621);
nor U2175 (N_2175,N_1938,N_1663);
and U2176 (N_2176,N_1635,N_1892);
or U2177 (N_2177,N_1936,N_1897);
xnor U2178 (N_2178,N_1523,N_1542);
or U2179 (N_2179,N_1886,N_1956);
nor U2180 (N_2180,N_1746,N_1817);
or U2181 (N_2181,N_1713,N_1685);
nor U2182 (N_2182,N_1875,N_1654);
nor U2183 (N_2183,N_1880,N_1702);
nand U2184 (N_2184,N_1770,N_1821);
nor U2185 (N_2185,N_1934,N_1879);
and U2186 (N_2186,N_1914,N_1848);
or U2187 (N_2187,N_1948,N_1747);
nand U2188 (N_2188,N_1926,N_1554);
nor U2189 (N_2189,N_1862,N_1741);
and U2190 (N_2190,N_1797,N_1823);
nand U2191 (N_2191,N_1594,N_1661);
nor U2192 (N_2192,N_1750,N_1565);
and U2193 (N_2193,N_1616,N_1620);
and U2194 (N_2194,N_1720,N_1585);
or U2195 (N_2195,N_1968,N_1726);
nor U2196 (N_2196,N_1602,N_1572);
nor U2197 (N_2197,N_1639,N_1884);
and U2198 (N_2198,N_1900,N_1656);
or U2199 (N_2199,N_1836,N_1615);
and U2200 (N_2200,N_1693,N_1571);
nand U2201 (N_2201,N_1664,N_1776);
nand U2202 (N_2202,N_1606,N_1814);
or U2203 (N_2203,N_1982,N_1527);
and U2204 (N_2204,N_1524,N_1849);
and U2205 (N_2205,N_1805,N_1504);
nor U2206 (N_2206,N_1543,N_1824);
or U2207 (N_2207,N_1962,N_1595);
and U2208 (N_2208,N_1887,N_1614);
and U2209 (N_2209,N_1997,N_1648);
nor U2210 (N_2210,N_1507,N_1765);
nor U2211 (N_2211,N_1707,N_1732);
nor U2212 (N_2212,N_1630,N_1687);
or U2213 (N_2213,N_1905,N_1539);
nor U2214 (N_2214,N_1582,N_1699);
nor U2215 (N_2215,N_1932,N_1736);
nor U2216 (N_2216,N_1966,N_1660);
nor U2217 (N_2217,N_1852,N_1555);
nand U2218 (N_2218,N_1869,N_1675);
nor U2219 (N_2219,N_1653,N_1680);
nand U2220 (N_2220,N_1609,N_1868);
and U2221 (N_2221,N_1786,N_1780);
or U2222 (N_2222,N_1791,N_1560);
nand U2223 (N_2223,N_1986,N_1866);
xor U2224 (N_2224,N_1845,N_1802);
nand U2225 (N_2225,N_1512,N_1536);
or U2226 (N_2226,N_1945,N_1537);
nor U2227 (N_2227,N_1522,N_1894);
nor U2228 (N_2228,N_1861,N_1946);
or U2229 (N_2229,N_1969,N_1789);
or U2230 (N_2230,N_1813,N_1798);
or U2231 (N_2231,N_1899,N_1976);
or U2232 (N_2232,N_1546,N_1549);
and U2233 (N_2233,N_1684,N_1538);
nand U2234 (N_2234,N_1781,N_1601);
or U2235 (N_2235,N_1712,N_1843);
and U2236 (N_2236,N_1801,N_1753);
or U2237 (N_2237,N_1593,N_1678);
and U2238 (N_2238,N_1625,N_1631);
and U2239 (N_2239,N_1657,N_1651);
or U2240 (N_2240,N_1759,N_1628);
and U2241 (N_2241,N_1718,N_1516);
or U2242 (N_2242,N_1872,N_1521);
nor U2243 (N_2243,N_1528,N_1771);
and U2244 (N_2244,N_1703,N_1935);
or U2245 (N_2245,N_1996,N_1579);
or U2246 (N_2246,N_1827,N_1959);
nand U2247 (N_2247,N_1939,N_1670);
and U2248 (N_2248,N_1984,N_1995);
or U2249 (N_2249,N_1667,N_1907);
or U2250 (N_2250,N_1914,N_1751);
and U2251 (N_2251,N_1524,N_1880);
nand U2252 (N_2252,N_1596,N_1852);
nand U2253 (N_2253,N_1793,N_1663);
and U2254 (N_2254,N_1695,N_1846);
and U2255 (N_2255,N_1924,N_1533);
nor U2256 (N_2256,N_1939,N_1706);
or U2257 (N_2257,N_1749,N_1904);
nor U2258 (N_2258,N_1917,N_1890);
and U2259 (N_2259,N_1553,N_1529);
nor U2260 (N_2260,N_1586,N_1501);
nor U2261 (N_2261,N_1976,N_1678);
nand U2262 (N_2262,N_1595,N_1946);
nand U2263 (N_2263,N_1868,N_1644);
or U2264 (N_2264,N_1852,N_1883);
xor U2265 (N_2265,N_1611,N_1930);
nor U2266 (N_2266,N_1793,N_1886);
and U2267 (N_2267,N_1581,N_1925);
or U2268 (N_2268,N_1938,N_1924);
nor U2269 (N_2269,N_1932,N_1900);
nand U2270 (N_2270,N_1975,N_1661);
nor U2271 (N_2271,N_1880,N_1947);
and U2272 (N_2272,N_1540,N_1641);
nor U2273 (N_2273,N_1717,N_1892);
or U2274 (N_2274,N_1702,N_1859);
or U2275 (N_2275,N_1939,N_1821);
or U2276 (N_2276,N_1743,N_1508);
and U2277 (N_2277,N_1947,N_1592);
nand U2278 (N_2278,N_1552,N_1895);
or U2279 (N_2279,N_1953,N_1699);
and U2280 (N_2280,N_1953,N_1989);
and U2281 (N_2281,N_1983,N_1859);
xnor U2282 (N_2282,N_1752,N_1571);
nand U2283 (N_2283,N_1994,N_1908);
and U2284 (N_2284,N_1613,N_1985);
xor U2285 (N_2285,N_1527,N_1538);
nand U2286 (N_2286,N_1706,N_1784);
and U2287 (N_2287,N_1983,N_1913);
nand U2288 (N_2288,N_1998,N_1806);
and U2289 (N_2289,N_1651,N_1818);
xnor U2290 (N_2290,N_1875,N_1818);
nand U2291 (N_2291,N_1962,N_1632);
nor U2292 (N_2292,N_1525,N_1797);
or U2293 (N_2293,N_1792,N_1617);
nor U2294 (N_2294,N_1735,N_1906);
and U2295 (N_2295,N_1533,N_1650);
nand U2296 (N_2296,N_1996,N_1938);
or U2297 (N_2297,N_1758,N_1874);
or U2298 (N_2298,N_1960,N_1535);
nand U2299 (N_2299,N_1617,N_1652);
nand U2300 (N_2300,N_1661,N_1658);
or U2301 (N_2301,N_1760,N_1685);
nor U2302 (N_2302,N_1708,N_1595);
nor U2303 (N_2303,N_1612,N_1983);
nand U2304 (N_2304,N_1946,N_1821);
nand U2305 (N_2305,N_1892,N_1876);
nand U2306 (N_2306,N_1645,N_1833);
nor U2307 (N_2307,N_1989,N_1602);
nand U2308 (N_2308,N_1646,N_1764);
nand U2309 (N_2309,N_1775,N_1519);
nor U2310 (N_2310,N_1616,N_1996);
nand U2311 (N_2311,N_1927,N_1850);
and U2312 (N_2312,N_1577,N_1699);
and U2313 (N_2313,N_1993,N_1960);
nor U2314 (N_2314,N_1791,N_1589);
and U2315 (N_2315,N_1873,N_1710);
nand U2316 (N_2316,N_1605,N_1842);
nand U2317 (N_2317,N_1811,N_1992);
or U2318 (N_2318,N_1617,N_1507);
nand U2319 (N_2319,N_1685,N_1997);
or U2320 (N_2320,N_1663,N_1651);
and U2321 (N_2321,N_1690,N_1624);
nor U2322 (N_2322,N_1865,N_1670);
or U2323 (N_2323,N_1760,N_1704);
and U2324 (N_2324,N_1771,N_1879);
and U2325 (N_2325,N_1502,N_1685);
nand U2326 (N_2326,N_1739,N_1762);
nand U2327 (N_2327,N_1730,N_1941);
and U2328 (N_2328,N_1795,N_1565);
nand U2329 (N_2329,N_1643,N_1941);
nor U2330 (N_2330,N_1612,N_1740);
or U2331 (N_2331,N_1888,N_1974);
nor U2332 (N_2332,N_1735,N_1917);
nor U2333 (N_2333,N_1718,N_1824);
nor U2334 (N_2334,N_1840,N_1626);
and U2335 (N_2335,N_1829,N_1814);
nand U2336 (N_2336,N_1865,N_1721);
nor U2337 (N_2337,N_1783,N_1593);
or U2338 (N_2338,N_1875,N_1963);
nand U2339 (N_2339,N_1568,N_1728);
nor U2340 (N_2340,N_1563,N_1981);
or U2341 (N_2341,N_1837,N_1865);
nand U2342 (N_2342,N_1988,N_1773);
and U2343 (N_2343,N_1728,N_1925);
nor U2344 (N_2344,N_1873,N_1605);
and U2345 (N_2345,N_1937,N_1588);
or U2346 (N_2346,N_1599,N_1671);
or U2347 (N_2347,N_1544,N_1584);
and U2348 (N_2348,N_1594,N_1838);
or U2349 (N_2349,N_1921,N_1973);
and U2350 (N_2350,N_1574,N_1811);
or U2351 (N_2351,N_1609,N_1719);
or U2352 (N_2352,N_1996,N_1869);
xnor U2353 (N_2353,N_1514,N_1842);
nand U2354 (N_2354,N_1693,N_1718);
or U2355 (N_2355,N_1687,N_1545);
nor U2356 (N_2356,N_1896,N_1624);
or U2357 (N_2357,N_1576,N_1884);
or U2358 (N_2358,N_1690,N_1621);
and U2359 (N_2359,N_1943,N_1834);
or U2360 (N_2360,N_1684,N_1870);
nand U2361 (N_2361,N_1774,N_1789);
nand U2362 (N_2362,N_1868,N_1883);
nand U2363 (N_2363,N_1902,N_1767);
and U2364 (N_2364,N_1860,N_1952);
and U2365 (N_2365,N_1980,N_1731);
nor U2366 (N_2366,N_1520,N_1661);
and U2367 (N_2367,N_1839,N_1988);
and U2368 (N_2368,N_1615,N_1662);
nand U2369 (N_2369,N_1744,N_1503);
nand U2370 (N_2370,N_1774,N_1870);
nand U2371 (N_2371,N_1603,N_1519);
or U2372 (N_2372,N_1784,N_1770);
and U2373 (N_2373,N_1941,N_1673);
or U2374 (N_2374,N_1599,N_1959);
nand U2375 (N_2375,N_1849,N_1694);
and U2376 (N_2376,N_1648,N_1774);
or U2377 (N_2377,N_1527,N_1615);
and U2378 (N_2378,N_1957,N_1751);
nor U2379 (N_2379,N_1730,N_1763);
and U2380 (N_2380,N_1562,N_1914);
and U2381 (N_2381,N_1568,N_1607);
nor U2382 (N_2382,N_1902,N_1557);
or U2383 (N_2383,N_1618,N_1807);
nor U2384 (N_2384,N_1756,N_1874);
or U2385 (N_2385,N_1893,N_1705);
or U2386 (N_2386,N_1559,N_1830);
or U2387 (N_2387,N_1992,N_1999);
xnor U2388 (N_2388,N_1914,N_1829);
xnor U2389 (N_2389,N_1801,N_1891);
nand U2390 (N_2390,N_1850,N_1814);
or U2391 (N_2391,N_1593,N_1893);
and U2392 (N_2392,N_1922,N_1717);
nor U2393 (N_2393,N_1870,N_1934);
nand U2394 (N_2394,N_1526,N_1505);
nand U2395 (N_2395,N_1704,N_1795);
or U2396 (N_2396,N_1735,N_1649);
or U2397 (N_2397,N_1517,N_1710);
nor U2398 (N_2398,N_1972,N_1671);
xnor U2399 (N_2399,N_1547,N_1695);
and U2400 (N_2400,N_1535,N_1809);
or U2401 (N_2401,N_1538,N_1648);
or U2402 (N_2402,N_1563,N_1573);
or U2403 (N_2403,N_1885,N_1766);
and U2404 (N_2404,N_1739,N_1733);
nand U2405 (N_2405,N_1564,N_1807);
nand U2406 (N_2406,N_1636,N_1684);
and U2407 (N_2407,N_1769,N_1865);
and U2408 (N_2408,N_1627,N_1961);
and U2409 (N_2409,N_1962,N_1932);
or U2410 (N_2410,N_1977,N_1879);
nand U2411 (N_2411,N_1689,N_1712);
nor U2412 (N_2412,N_1537,N_1599);
nor U2413 (N_2413,N_1731,N_1769);
nand U2414 (N_2414,N_1811,N_1581);
and U2415 (N_2415,N_1924,N_1904);
nand U2416 (N_2416,N_1547,N_1951);
or U2417 (N_2417,N_1568,N_1788);
or U2418 (N_2418,N_1750,N_1628);
nand U2419 (N_2419,N_1533,N_1539);
or U2420 (N_2420,N_1835,N_1723);
nor U2421 (N_2421,N_1967,N_1939);
nor U2422 (N_2422,N_1573,N_1831);
or U2423 (N_2423,N_1602,N_1885);
nor U2424 (N_2424,N_1744,N_1649);
or U2425 (N_2425,N_1663,N_1706);
and U2426 (N_2426,N_1740,N_1771);
and U2427 (N_2427,N_1898,N_1772);
nand U2428 (N_2428,N_1683,N_1984);
or U2429 (N_2429,N_1610,N_1854);
nor U2430 (N_2430,N_1958,N_1802);
and U2431 (N_2431,N_1978,N_1588);
and U2432 (N_2432,N_1615,N_1502);
or U2433 (N_2433,N_1782,N_1805);
or U2434 (N_2434,N_1823,N_1565);
or U2435 (N_2435,N_1972,N_1737);
or U2436 (N_2436,N_1828,N_1696);
or U2437 (N_2437,N_1658,N_1521);
nor U2438 (N_2438,N_1999,N_1952);
or U2439 (N_2439,N_1633,N_1978);
and U2440 (N_2440,N_1563,N_1917);
or U2441 (N_2441,N_1923,N_1851);
or U2442 (N_2442,N_1985,N_1899);
nand U2443 (N_2443,N_1944,N_1590);
and U2444 (N_2444,N_1792,N_1948);
nand U2445 (N_2445,N_1782,N_1983);
nand U2446 (N_2446,N_1509,N_1937);
nor U2447 (N_2447,N_1665,N_1810);
xnor U2448 (N_2448,N_1727,N_1617);
or U2449 (N_2449,N_1944,N_1584);
nand U2450 (N_2450,N_1727,N_1958);
or U2451 (N_2451,N_1724,N_1798);
nor U2452 (N_2452,N_1701,N_1843);
nor U2453 (N_2453,N_1983,N_1528);
nand U2454 (N_2454,N_1812,N_1942);
and U2455 (N_2455,N_1653,N_1804);
and U2456 (N_2456,N_1750,N_1904);
and U2457 (N_2457,N_1794,N_1763);
nor U2458 (N_2458,N_1525,N_1722);
or U2459 (N_2459,N_1562,N_1803);
nand U2460 (N_2460,N_1804,N_1910);
or U2461 (N_2461,N_1553,N_1913);
and U2462 (N_2462,N_1619,N_1956);
nand U2463 (N_2463,N_1798,N_1716);
nand U2464 (N_2464,N_1536,N_1809);
or U2465 (N_2465,N_1952,N_1937);
nor U2466 (N_2466,N_1909,N_1577);
or U2467 (N_2467,N_1503,N_1796);
and U2468 (N_2468,N_1655,N_1589);
or U2469 (N_2469,N_1739,N_1995);
nand U2470 (N_2470,N_1971,N_1968);
nand U2471 (N_2471,N_1701,N_1945);
and U2472 (N_2472,N_1736,N_1833);
and U2473 (N_2473,N_1609,N_1568);
nand U2474 (N_2474,N_1631,N_1918);
or U2475 (N_2475,N_1594,N_1739);
nand U2476 (N_2476,N_1635,N_1611);
nand U2477 (N_2477,N_1837,N_1839);
and U2478 (N_2478,N_1556,N_1587);
nand U2479 (N_2479,N_1833,N_1765);
and U2480 (N_2480,N_1843,N_1870);
and U2481 (N_2481,N_1807,N_1650);
and U2482 (N_2482,N_1548,N_1896);
and U2483 (N_2483,N_1972,N_1830);
nor U2484 (N_2484,N_1932,N_1537);
and U2485 (N_2485,N_1565,N_1690);
nand U2486 (N_2486,N_1992,N_1894);
or U2487 (N_2487,N_1555,N_1831);
and U2488 (N_2488,N_1818,N_1903);
or U2489 (N_2489,N_1734,N_1925);
and U2490 (N_2490,N_1544,N_1812);
nand U2491 (N_2491,N_1631,N_1564);
or U2492 (N_2492,N_1896,N_1581);
or U2493 (N_2493,N_1623,N_1523);
or U2494 (N_2494,N_1901,N_1615);
nor U2495 (N_2495,N_1670,N_1963);
or U2496 (N_2496,N_1751,N_1741);
or U2497 (N_2497,N_1556,N_1908);
nor U2498 (N_2498,N_1765,N_1788);
nand U2499 (N_2499,N_1841,N_1955);
or U2500 (N_2500,N_2100,N_2337);
nor U2501 (N_2501,N_2260,N_2247);
or U2502 (N_2502,N_2188,N_2072);
nor U2503 (N_2503,N_2369,N_2138);
nand U2504 (N_2504,N_2114,N_2011);
nand U2505 (N_2505,N_2439,N_2020);
and U2506 (N_2506,N_2403,N_2264);
or U2507 (N_2507,N_2293,N_2469);
or U2508 (N_2508,N_2098,N_2161);
nand U2509 (N_2509,N_2480,N_2354);
and U2510 (N_2510,N_2099,N_2318);
or U2511 (N_2511,N_2300,N_2307);
nand U2512 (N_2512,N_2401,N_2249);
nor U2513 (N_2513,N_2071,N_2172);
nand U2514 (N_2514,N_2149,N_2066);
nor U2515 (N_2515,N_2039,N_2431);
or U2516 (N_2516,N_2177,N_2385);
and U2517 (N_2517,N_2267,N_2498);
xor U2518 (N_2518,N_2268,N_2007);
and U2519 (N_2519,N_2437,N_2196);
and U2520 (N_2520,N_2438,N_2010);
nor U2521 (N_2521,N_2362,N_2009);
nor U2522 (N_2522,N_2287,N_2468);
nor U2523 (N_2523,N_2269,N_2113);
and U2524 (N_2524,N_2005,N_2124);
and U2525 (N_2525,N_2187,N_2453);
and U2526 (N_2526,N_2340,N_2008);
nor U2527 (N_2527,N_2356,N_2237);
or U2528 (N_2528,N_2434,N_2065);
nor U2529 (N_2529,N_2279,N_2118);
nand U2530 (N_2530,N_2145,N_2359);
nand U2531 (N_2531,N_2165,N_2398);
or U2532 (N_2532,N_2430,N_2331);
nor U2533 (N_2533,N_2167,N_2125);
or U2534 (N_2534,N_2364,N_2189);
and U2535 (N_2535,N_2341,N_2421);
xor U2536 (N_2536,N_2240,N_2329);
nor U2537 (N_2537,N_2313,N_2069);
nor U2538 (N_2538,N_2164,N_2484);
xor U2539 (N_2539,N_2327,N_2326);
nand U2540 (N_2540,N_2408,N_2075);
nor U2541 (N_2541,N_2257,N_2224);
or U2542 (N_2542,N_2083,N_2481);
or U2543 (N_2543,N_2241,N_2054);
nor U2544 (N_2544,N_2328,N_2272);
nand U2545 (N_2545,N_2001,N_2197);
and U2546 (N_2546,N_2201,N_2088);
and U2547 (N_2547,N_2076,N_2162);
nor U2548 (N_2548,N_2312,N_2345);
and U2549 (N_2549,N_2030,N_2393);
nor U2550 (N_2550,N_2184,N_2414);
or U2551 (N_2551,N_2296,N_2425);
and U2552 (N_2552,N_2426,N_2049);
and U2553 (N_2553,N_2116,N_2226);
nor U2554 (N_2554,N_2253,N_2238);
nand U2555 (N_2555,N_2127,N_2455);
or U2556 (N_2556,N_2220,N_2308);
or U2557 (N_2557,N_2281,N_2420);
nand U2558 (N_2558,N_2277,N_2415);
and U2559 (N_2559,N_2466,N_2360);
and U2560 (N_2560,N_2064,N_2273);
nand U2561 (N_2561,N_2274,N_2015);
nand U2562 (N_2562,N_2407,N_2367);
or U2563 (N_2563,N_2129,N_2440);
and U2564 (N_2564,N_2456,N_2255);
nor U2565 (N_2565,N_2106,N_2024);
nand U2566 (N_2566,N_2060,N_2085);
nand U2567 (N_2567,N_2244,N_2034);
or U2568 (N_2568,N_2306,N_2488);
and U2569 (N_2569,N_2483,N_2057);
and U2570 (N_2570,N_2284,N_2094);
or U2571 (N_2571,N_2235,N_2265);
nand U2572 (N_2572,N_2061,N_2482);
and U2573 (N_2573,N_2233,N_2042);
nand U2574 (N_2574,N_2381,N_2006);
nand U2575 (N_2575,N_2448,N_2317);
nor U2576 (N_2576,N_2454,N_2387);
or U2577 (N_2577,N_2150,N_2459);
nand U2578 (N_2578,N_2029,N_2128);
or U2579 (N_2579,N_2082,N_2391);
and U2580 (N_2580,N_2019,N_2036);
nand U2581 (N_2581,N_2266,N_2144);
or U2582 (N_2582,N_2147,N_2378);
and U2583 (N_2583,N_2014,N_2348);
nand U2584 (N_2584,N_2027,N_2262);
and U2585 (N_2585,N_2117,N_2315);
or U2586 (N_2586,N_2092,N_2351);
nor U2587 (N_2587,N_2416,N_2256);
and U2588 (N_2588,N_2396,N_2368);
xor U2589 (N_2589,N_2097,N_2462);
xor U2590 (N_2590,N_2428,N_2413);
nand U2591 (N_2591,N_2436,N_2151);
and U2592 (N_2592,N_2176,N_2204);
nor U2593 (N_2593,N_2397,N_2089);
and U2594 (N_2594,N_2031,N_2294);
or U2595 (N_2595,N_2347,N_2219);
or U2596 (N_2596,N_2342,N_2336);
nand U2597 (N_2597,N_2242,N_2423);
nand U2598 (N_2598,N_2160,N_2230);
nand U2599 (N_2599,N_2195,N_2377);
and U2600 (N_2600,N_2252,N_2355);
nor U2601 (N_2601,N_2166,N_2101);
or U2602 (N_2602,N_2035,N_2451);
nor U2603 (N_2603,N_2096,N_2363);
and U2604 (N_2604,N_2000,N_2492);
or U2605 (N_2605,N_2334,N_2146);
and U2606 (N_2606,N_2429,N_2032);
or U2607 (N_2607,N_2221,N_2476);
nand U2608 (N_2608,N_2003,N_2074);
or U2609 (N_2609,N_2048,N_2209);
or U2610 (N_2610,N_2471,N_2215);
xor U2611 (N_2611,N_2495,N_2297);
or U2612 (N_2612,N_2087,N_2133);
nor U2613 (N_2613,N_2119,N_2388);
nand U2614 (N_2614,N_2109,N_2173);
or U2615 (N_2615,N_2491,N_2270);
nor U2616 (N_2616,N_2142,N_2384);
xor U2617 (N_2617,N_2446,N_2325);
nor U2618 (N_2618,N_2283,N_2261);
or U2619 (N_2619,N_2419,N_2225);
or U2620 (N_2620,N_2395,N_2250);
and U2621 (N_2621,N_2460,N_2207);
nand U2622 (N_2622,N_2223,N_2135);
and U2623 (N_2623,N_2494,N_2344);
and U2624 (N_2624,N_2259,N_2289);
nor U2625 (N_2625,N_2450,N_2159);
and U2626 (N_2626,N_2322,N_2357);
nor U2627 (N_2627,N_2153,N_2409);
nor U2628 (N_2628,N_2121,N_2496);
and U2629 (N_2629,N_2246,N_2120);
nand U2630 (N_2630,N_2465,N_2012);
nor U2631 (N_2631,N_2406,N_2132);
nor U2632 (N_2632,N_2021,N_2490);
or U2633 (N_2633,N_2339,N_2070);
nor U2634 (N_2634,N_2411,N_2206);
and U2635 (N_2635,N_2033,N_2234);
or U2636 (N_2636,N_2126,N_2123);
or U2637 (N_2637,N_2473,N_2055);
nand U2638 (N_2638,N_2093,N_2169);
or U2639 (N_2639,N_2485,N_2077);
and U2640 (N_2640,N_2371,N_2479);
nand U2641 (N_2641,N_2102,N_2467);
and U2642 (N_2642,N_2280,N_2143);
nor U2643 (N_2643,N_2067,N_2245);
and U2644 (N_2644,N_2276,N_2310);
or U2645 (N_2645,N_2137,N_2464);
or U2646 (N_2646,N_2412,N_2386);
and U2647 (N_2647,N_2227,N_2474);
or U2648 (N_2648,N_2078,N_2158);
nand U2649 (N_2649,N_2285,N_2047);
nand U2650 (N_2650,N_2002,N_2194);
nand U2651 (N_2651,N_2497,N_2410);
nand U2652 (N_2652,N_2258,N_2489);
or U2653 (N_2653,N_2185,N_2402);
nor U2654 (N_2654,N_2372,N_2288);
and U2655 (N_2655,N_2040,N_2292);
nor U2656 (N_2656,N_2190,N_2346);
nor U2657 (N_2657,N_2263,N_2290);
xor U2658 (N_2658,N_2148,N_2418);
or U2659 (N_2659,N_2338,N_2374);
or U2660 (N_2660,N_2063,N_2405);
and U2661 (N_2661,N_2051,N_2352);
and U2662 (N_2662,N_2236,N_2320);
nor U2663 (N_2663,N_2081,N_2191);
and U2664 (N_2664,N_2330,N_2435);
nor U2665 (N_2665,N_2463,N_2136);
and U2666 (N_2666,N_2095,N_2458);
or U2667 (N_2667,N_2291,N_2461);
or U2668 (N_2668,N_2168,N_2068);
xnor U2669 (N_2669,N_2013,N_2175);
and U2670 (N_2670,N_2400,N_2472);
nor U2671 (N_2671,N_2248,N_2432);
and U2672 (N_2672,N_2487,N_2321);
nor U2673 (N_2673,N_2422,N_2140);
nand U2674 (N_2674,N_2470,N_2373);
xor U2675 (N_2675,N_2202,N_2311);
nor U2676 (N_2676,N_2080,N_2174);
and U2677 (N_2677,N_2037,N_2383);
nand U2678 (N_2678,N_2286,N_2323);
nor U2679 (N_2679,N_2442,N_2130);
nand U2680 (N_2680,N_2239,N_2155);
nor U2681 (N_2681,N_2324,N_2376);
nor U2682 (N_2682,N_2399,N_2445);
or U2683 (N_2683,N_2375,N_2349);
nand U2684 (N_2684,N_2427,N_2016);
or U2685 (N_2685,N_2053,N_2108);
or U2686 (N_2686,N_2303,N_2271);
nor U2687 (N_2687,N_2319,N_2218);
or U2688 (N_2688,N_2449,N_2079);
or U2689 (N_2689,N_2305,N_2379);
nor U2690 (N_2690,N_2208,N_2335);
nor U2691 (N_2691,N_2231,N_2365);
and U2692 (N_2692,N_2141,N_2105);
nor U2693 (N_2693,N_2170,N_2314);
and U2694 (N_2694,N_2433,N_2275);
xnor U2695 (N_2695,N_2110,N_2192);
nand U2696 (N_2696,N_2229,N_2183);
nor U2697 (N_2697,N_2073,N_2182);
or U2698 (N_2698,N_2045,N_2107);
and U2699 (N_2699,N_2026,N_2193);
nand U2700 (N_2700,N_2392,N_2028);
and U2701 (N_2701,N_2200,N_2090);
nand U2702 (N_2702,N_2217,N_2380);
nor U2703 (N_2703,N_2022,N_2447);
nor U2704 (N_2704,N_2350,N_2366);
nand U2705 (N_2705,N_2046,N_2056);
nor U2706 (N_2706,N_2361,N_2298);
or U2707 (N_2707,N_2186,N_2424);
and U2708 (N_2708,N_2404,N_2232);
or U2709 (N_2709,N_2389,N_2104);
and U2710 (N_2710,N_2216,N_2486);
nand U2711 (N_2711,N_2086,N_2417);
nor U2712 (N_2712,N_2301,N_2043);
and U2713 (N_2713,N_2154,N_2332);
nand U2714 (N_2714,N_2199,N_2278);
nand U2715 (N_2715,N_2452,N_2163);
nand U2716 (N_2716,N_2052,N_2475);
and U2717 (N_2717,N_2198,N_2018);
and U2718 (N_2718,N_2302,N_2059);
nand U2719 (N_2719,N_2103,N_2139);
or U2720 (N_2720,N_2004,N_2058);
or U2721 (N_2721,N_2044,N_2222);
xor U2722 (N_2722,N_2316,N_2025);
nor U2723 (N_2723,N_2181,N_2309);
or U2724 (N_2724,N_2023,N_2251);
nand U2725 (N_2725,N_2203,N_2304);
and U2726 (N_2726,N_2214,N_2243);
nor U2727 (N_2727,N_2370,N_2282);
or U2728 (N_2728,N_2091,N_2112);
or U2729 (N_2729,N_2178,N_2062);
nor U2730 (N_2730,N_2111,N_2210);
nand U2731 (N_2731,N_2211,N_2041);
or U2732 (N_2732,N_2205,N_2493);
nand U2733 (N_2733,N_2499,N_2171);
nor U2734 (N_2734,N_2457,N_2441);
nand U2735 (N_2735,N_2394,N_2017);
or U2736 (N_2736,N_2213,N_2115);
or U2737 (N_2737,N_2353,N_2228);
nand U2738 (N_2738,N_2212,N_2382);
nand U2739 (N_2739,N_2299,N_2343);
or U2740 (N_2740,N_2156,N_2358);
or U2741 (N_2741,N_2444,N_2122);
or U2742 (N_2742,N_2134,N_2333);
nand U2743 (N_2743,N_2084,N_2180);
nand U2744 (N_2744,N_2390,N_2254);
or U2745 (N_2745,N_2038,N_2478);
nand U2746 (N_2746,N_2477,N_2443);
nand U2747 (N_2747,N_2157,N_2152);
nor U2748 (N_2748,N_2295,N_2179);
nand U2749 (N_2749,N_2131,N_2050);
or U2750 (N_2750,N_2209,N_2499);
and U2751 (N_2751,N_2391,N_2136);
or U2752 (N_2752,N_2443,N_2434);
and U2753 (N_2753,N_2172,N_2101);
nor U2754 (N_2754,N_2324,N_2150);
nand U2755 (N_2755,N_2276,N_2428);
or U2756 (N_2756,N_2273,N_2257);
nor U2757 (N_2757,N_2435,N_2343);
nor U2758 (N_2758,N_2430,N_2115);
or U2759 (N_2759,N_2426,N_2402);
nand U2760 (N_2760,N_2207,N_2356);
or U2761 (N_2761,N_2122,N_2449);
and U2762 (N_2762,N_2386,N_2096);
nor U2763 (N_2763,N_2145,N_2033);
nor U2764 (N_2764,N_2016,N_2147);
nor U2765 (N_2765,N_2062,N_2478);
or U2766 (N_2766,N_2278,N_2052);
nand U2767 (N_2767,N_2371,N_2406);
or U2768 (N_2768,N_2318,N_2461);
or U2769 (N_2769,N_2133,N_2262);
nor U2770 (N_2770,N_2448,N_2332);
or U2771 (N_2771,N_2478,N_2041);
xor U2772 (N_2772,N_2255,N_2285);
nor U2773 (N_2773,N_2449,N_2093);
nand U2774 (N_2774,N_2347,N_2418);
nand U2775 (N_2775,N_2134,N_2137);
or U2776 (N_2776,N_2485,N_2258);
or U2777 (N_2777,N_2114,N_2303);
nor U2778 (N_2778,N_2375,N_2105);
or U2779 (N_2779,N_2132,N_2128);
and U2780 (N_2780,N_2128,N_2337);
and U2781 (N_2781,N_2242,N_2293);
nand U2782 (N_2782,N_2451,N_2056);
xnor U2783 (N_2783,N_2345,N_2066);
nand U2784 (N_2784,N_2204,N_2377);
and U2785 (N_2785,N_2170,N_2299);
or U2786 (N_2786,N_2098,N_2121);
or U2787 (N_2787,N_2391,N_2225);
and U2788 (N_2788,N_2196,N_2075);
nor U2789 (N_2789,N_2432,N_2257);
nor U2790 (N_2790,N_2314,N_2486);
or U2791 (N_2791,N_2433,N_2235);
nor U2792 (N_2792,N_2390,N_2022);
nor U2793 (N_2793,N_2129,N_2163);
or U2794 (N_2794,N_2201,N_2391);
nand U2795 (N_2795,N_2489,N_2311);
nor U2796 (N_2796,N_2493,N_2334);
or U2797 (N_2797,N_2172,N_2421);
and U2798 (N_2798,N_2091,N_2074);
nand U2799 (N_2799,N_2194,N_2260);
and U2800 (N_2800,N_2119,N_2285);
or U2801 (N_2801,N_2036,N_2210);
nand U2802 (N_2802,N_2252,N_2067);
nand U2803 (N_2803,N_2147,N_2443);
nor U2804 (N_2804,N_2132,N_2349);
nand U2805 (N_2805,N_2422,N_2324);
nor U2806 (N_2806,N_2431,N_2421);
nand U2807 (N_2807,N_2120,N_2331);
nand U2808 (N_2808,N_2072,N_2467);
nor U2809 (N_2809,N_2445,N_2240);
nor U2810 (N_2810,N_2022,N_2149);
and U2811 (N_2811,N_2163,N_2382);
or U2812 (N_2812,N_2145,N_2082);
or U2813 (N_2813,N_2034,N_2274);
and U2814 (N_2814,N_2425,N_2197);
or U2815 (N_2815,N_2069,N_2420);
and U2816 (N_2816,N_2422,N_2117);
and U2817 (N_2817,N_2477,N_2499);
and U2818 (N_2818,N_2046,N_2173);
and U2819 (N_2819,N_2379,N_2412);
nor U2820 (N_2820,N_2435,N_2206);
and U2821 (N_2821,N_2088,N_2218);
or U2822 (N_2822,N_2254,N_2475);
or U2823 (N_2823,N_2034,N_2083);
nand U2824 (N_2824,N_2134,N_2033);
or U2825 (N_2825,N_2286,N_2121);
or U2826 (N_2826,N_2257,N_2242);
nand U2827 (N_2827,N_2420,N_2208);
and U2828 (N_2828,N_2351,N_2338);
and U2829 (N_2829,N_2424,N_2063);
nor U2830 (N_2830,N_2017,N_2282);
or U2831 (N_2831,N_2140,N_2352);
and U2832 (N_2832,N_2401,N_2001);
nand U2833 (N_2833,N_2424,N_2411);
and U2834 (N_2834,N_2071,N_2280);
and U2835 (N_2835,N_2242,N_2230);
nor U2836 (N_2836,N_2246,N_2147);
nor U2837 (N_2837,N_2158,N_2174);
nand U2838 (N_2838,N_2496,N_2054);
and U2839 (N_2839,N_2428,N_2489);
nor U2840 (N_2840,N_2338,N_2429);
nor U2841 (N_2841,N_2226,N_2461);
nand U2842 (N_2842,N_2252,N_2458);
nor U2843 (N_2843,N_2089,N_2221);
or U2844 (N_2844,N_2184,N_2124);
nand U2845 (N_2845,N_2409,N_2032);
nor U2846 (N_2846,N_2322,N_2369);
nand U2847 (N_2847,N_2104,N_2296);
and U2848 (N_2848,N_2488,N_2064);
or U2849 (N_2849,N_2197,N_2343);
or U2850 (N_2850,N_2386,N_2466);
and U2851 (N_2851,N_2288,N_2061);
nand U2852 (N_2852,N_2241,N_2456);
nand U2853 (N_2853,N_2493,N_2251);
nor U2854 (N_2854,N_2244,N_2417);
nor U2855 (N_2855,N_2428,N_2246);
and U2856 (N_2856,N_2360,N_2175);
and U2857 (N_2857,N_2179,N_2236);
nand U2858 (N_2858,N_2349,N_2225);
or U2859 (N_2859,N_2371,N_2237);
or U2860 (N_2860,N_2099,N_2369);
nor U2861 (N_2861,N_2274,N_2058);
nor U2862 (N_2862,N_2298,N_2006);
or U2863 (N_2863,N_2154,N_2404);
or U2864 (N_2864,N_2418,N_2231);
and U2865 (N_2865,N_2084,N_2233);
nand U2866 (N_2866,N_2272,N_2294);
and U2867 (N_2867,N_2444,N_2072);
nor U2868 (N_2868,N_2413,N_2389);
xor U2869 (N_2869,N_2312,N_2359);
or U2870 (N_2870,N_2392,N_2352);
nand U2871 (N_2871,N_2319,N_2246);
nand U2872 (N_2872,N_2491,N_2424);
or U2873 (N_2873,N_2441,N_2027);
and U2874 (N_2874,N_2018,N_2273);
or U2875 (N_2875,N_2393,N_2085);
nor U2876 (N_2876,N_2296,N_2447);
and U2877 (N_2877,N_2348,N_2471);
and U2878 (N_2878,N_2155,N_2337);
or U2879 (N_2879,N_2158,N_2364);
nor U2880 (N_2880,N_2287,N_2401);
and U2881 (N_2881,N_2470,N_2434);
and U2882 (N_2882,N_2314,N_2163);
nor U2883 (N_2883,N_2292,N_2461);
nor U2884 (N_2884,N_2277,N_2442);
or U2885 (N_2885,N_2040,N_2332);
nor U2886 (N_2886,N_2335,N_2223);
and U2887 (N_2887,N_2204,N_2125);
nand U2888 (N_2888,N_2313,N_2104);
or U2889 (N_2889,N_2421,N_2215);
or U2890 (N_2890,N_2187,N_2219);
and U2891 (N_2891,N_2427,N_2004);
nor U2892 (N_2892,N_2309,N_2111);
and U2893 (N_2893,N_2296,N_2370);
or U2894 (N_2894,N_2300,N_2271);
or U2895 (N_2895,N_2400,N_2431);
and U2896 (N_2896,N_2385,N_2284);
and U2897 (N_2897,N_2437,N_2118);
or U2898 (N_2898,N_2037,N_2409);
and U2899 (N_2899,N_2494,N_2041);
and U2900 (N_2900,N_2335,N_2164);
or U2901 (N_2901,N_2220,N_2277);
and U2902 (N_2902,N_2175,N_2338);
nor U2903 (N_2903,N_2196,N_2171);
nand U2904 (N_2904,N_2111,N_2473);
nand U2905 (N_2905,N_2294,N_2276);
nand U2906 (N_2906,N_2201,N_2337);
and U2907 (N_2907,N_2289,N_2168);
nor U2908 (N_2908,N_2165,N_2121);
nand U2909 (N_2909,N_2025,N_2010);
or U2910 (N_2910,N_2283,N_2240);
nand U2911 (N_2911,N_2440,N_2418);
nand U2912 (N_2912,N_2140,N_2117);
and U2913 (N_2913,N_2268,N_2099);
or U2914 (N_2914,N_2270,N_2298);
nor U2915 (N_2915,N_2449,N_2454);
and U2916 (N_2916,N_2403,N_2399);
nor U2917 (N_2917,N_2155,N_2277);
or U2918 (N_2918,N_2269,N_2181);
nor U2919 (N_2919,N_2458,N_2283);
nor U2920 (N_2920,N_2153,N_2290);
or U2921 (N_2921,N_2162,N_2279);
and U2922 (N_2922,N_2361,N_2121);
and U2923 (N_2923,N_2236,N_2281);
or U2924 (N_2924,N_2383,N_2353);
xnor U2925 (N_2925,N_2365,N_2270);
and U2926 (N_2926,N_2210,N_2192);
nor U2927 (N_2927,N_2015,N_2066);
nand U2928 (N_2928,N_2118,N_2076);
and U2929 (N_2929,N_2487,N_2257);
and U2930 (N_2930,N_2263,N_2402);
or U2931 (N_2931,N_2286,N_2209);
nand U2932 (N_2932,N_2057,N_2465);
nand U2933 (N_2933,N_2441,N_2110);
and U2934 (N_2934,N_2285,N_2393);
nand U2935 (N_2935,N_2346,N_2415);
or U2936 (N_2936,N_2480,N_2238);
nor U2937 (N_2937,N_2062,N_2002);
and U2938 (N_2938,N_2106,N_2144);
nand U2939 (N_2939,N_2021,N_2435);
or U2940 (N_2940,N_2112,N_2130);
nand U2941 (N_2941,N_2459,N_2249);
and U2942 (N_2942,N_2061,N_2444);
nand U2943 (N_2943,N_2336,N_2470);
or U2944 (N_2944,N_2478,N_2250);
nand U2945 (N_2945,N_2076,N_2165);
nor U2946 (N_2946,N_2189,N_2353);
or U2947 (N_2947,N_2425,N_2227);
nand U2948 (N_2948,N_2312,N_2295);
nand U2949 (N_2949,N_2326,N_2010);
nor U2950 (N_2950,N_2039,N_2091);
nor U2951 (N_2951,N_2096,N_2469);
nor U2952 (N_2952,N_2134,N_2133);
and U2953 (N_2953,N_2375,N_2427);
or U2954 (N_2954,N_2098,N_2298);
and U2955 (N_2955,N_2353,N_2100);
nand U2956 (N_2956,N_2137,N_2099);
nor U2957 (N_2957,N_2071,N_2458);
or U2958 (N_2958,N_2212,N_2345);
and U2959 (N_2959,N_2302,N_2327);
nor U2960 (N_2960,N_2092,N_2427);
or U2961 (N_2961,N_2105,N_2351);
and U2962 (N_2962,N_2326,N_2334);
xnor U2963 (N_2963,N_2105,N_2178);
nand U2964 (N_2964,N_2451,N_2139);
xnor U2965 (N_2965,N_2315,N_2162);
nor U2966 (N_2966,N_2461,N_2254);
nand U2967 (N_2967,N_2450,N_2339);
nand U2968 (N_2968,N_2391,N_2435);
or U2969 (N_2969,N_2484,N_2421);
or U2970 (N_2970,N_2479,N_2458);
nor U2971 (N_2971,N_2330,N_2260);
and U2972 (N_2972,N_2117,N_2402);
nand U2973 (N_2973,N_2381,N_2180);
or U2974 (N_2974,N_2242,N_2310);
nand U2975 (N_2975,N_2046,N_2114);
nor U2976 (N_2976,N_2313,N_2176);
nor U2977 (N_2977,N_2003,N_2471);
nand U2978 (N_2978,N_2381,N_2179);
or U2979 (N_2979,N_2040,N_2213);
or U2980 (N_2980,N_2342,N_2300);
nand U2981 (N_2981,N_2101,N_2152);
nand U2982 (N_2982,N_2103,N_2255);
nand U2983 (N_2983,N_2441,N_2416);
nor U2984 (N_2984,N_2159,N_2053);
or U2985 (N_2985,N_2268,N_2495);
and U2986 (N_2986,N_2389,N_2294);
nand U2987 (N_2987,N_2301,N_2482);
nand U2988 (N_2988,N_2192,N_2416);
or U2989 (N_2989,N_2240,N_2474);
or U2990 (N_2990,N_2047,N_2340);
and U2991 (N_2991,N_2339,N_2277);
and U2992 (N_2992,N_2252,N_2092);
nor U2993 (N_2993,N_2393,N_2103);
or U2994 (N_2994,N_2490,N_2402);
and U2995 (N_2995,N_2249,N_2055);
or U2996 (N_2996,N_2464,N_2012);
nor U2997 (N_2997,N_2263,N_2431);
nand U2998 (N_2998,N_2431,N_2323);
or U2999 (N_2999,N_2381,N_2068);
nor UO_0 (O_0,N_2855,N_2973);
or UO_1 (O_1,N_2746,N_2588);
nand UO_2 (O_2,N_2529,N_2596);
or UO_3 (O_3,N_2925,N_2770);
nor UO_4 (O_4,N_2501,N_2920);
and UO_5 (O_5,N_2649,N_2790);
nand UO_6 (O_6,N_2924,N_2890);
nor UO_7 (O_7,N_2758,N_2764);
and UO_8 (O_8,N_2927,N_2772);
and UO_9 (O_9,N_2805,N_2697);
xor UO_10 (O_10,N_2503,N_2537);
nor UO_11 (O_11,N_2504,N_2775);
nor UO_12 (O_12,N_2765,N_2762);
nand UO_13 (O_13,N_2648,N_2892);
and UO_14 (O_14,N_2753,N_2943);
or UO_15 (O_15,N_2789,N_2827);
and UO_16 (O_16,N_2713,N_2558);
nor UO_17 (O_17,N_2694,N_2923);
or UO_18 (O_18,N_2657,N_2963);
and UO_19 (O_19,N_2593,N_2941);
and UO_20 (O_20,N_2771,N_2675);
and UO_21 (O_21,N_2612,N_2910);
nand UO_22 (O_22,N_2644,N_2954);
and UO_23 (O_23,N_2777,N_2806);
nand UO_24 (O_24,N_2922,N_2740);
nand UO_25 (O_25,N_2897,N_2522);
and UO_26 (O_26,N_2990,N_2718);
nor UO_27 (O_27,N_2668,N_2677);
or UO_28 (O_28,N_2662,N_2614);
nand UO_29 (O_29,N_2533,N_2549);
and UO_30 (O_30,N_2637,N_2751);
or UO_31 (O_31,N_2514,N_2725);
and UO_32 (O_32,N_2824,N_2802);
or UO_33 (O_33,N_2902,N_2717);
or UO_34 (O_34,N_2660,N_2520);
nand UO_35 (O_35,N_2800,N_2961);
or UO_36 (O_36,N_2951,N_2622);
or UO_37 (O_37,N_2987,N_2976);
or UO_38 (O_38,N_2926,N_2877);
nor UO_39 (O_39,N_2982,N_2852);
and UO_40 (O_40,N_2932,N_2761);
or UO_41 (O_41,N_2911,N_2848);
and UO_42 (O_42,N_2969,N_2566);
and UO_43 (O_43,N_2804,N_2613);
or UO_44 (O_44,N_2868,N_2842);
or UO_45 (O_45,N_2989,N_2913);
xor UO_46 (O_46,N_2864,N_2843);
nand UO_47 (O_47,N_2580,N_2985);
xnor UO_48 (O_48,N_2567,N_2665);
nor UO_49 (O_49,N_2658,N_2707);
and UO_50 (O_50,N_2791,N_2607);
nand UO_51 (O_51,N_2768,N_2659);
nor UO_52 (O_52,N_2543,N_2541);
xnor UO_53 (O_53,N_2851,N_2500);
nor UO_54 (O_54,N_2840,N_2507);
and UO_55 (O_55,N_2605,N_2524);
nor UO_56 (O_56,N_2623,N_2841);
and UO_57 (O_57,N_2886,N_2916);
and UO_58 (O_58,N_2896,N_2834);
or UO_59 (O_59,N_2914,N_2741);
xnor UO_60 (O_60,N_2749,N_2627);
and UO_61 (O_61,N_2516,N_2595);
and UO_62 (O_62,N_2705,N_2893);
xnor UO_63 (O_63,N_2819,N_2846);
and UO_64 (O_64,N_2950,N_2814);
or UO_65 (O_65,N_2933,N_2685);
or UO_66 (O_66,N_2517,N_2826);
and UO_67 (O_67,N_2722,N_2830);
and UO_68 (O_68,N_2590,N_2869);
nand UO_69 (O_69,N_2742,N_2734);
and UO_70 (O_70,N_2621,N_2945);
nand UO_71 (O_71,N_2988,N_2604);
and UO_72 (O_72,N_2701,N_2530);
or UO_73 (O_73,N_2519,N_2822);
nand UO_74 (O_74,N_2801,N_2652);
nand UO_75 (O_75,N_2872,N_2708);
nor UO_76 (O_76,N_2592,N_2556);
or UO_77 (O_77,N_2763,N_2617);
or UO_78 (O_78,N_2728,N_2774);
xor UO_79 (O_79,N_2818,N_2684);
nand UO_80 (O_80,N_2526,N_2642);
or UO_81 (O_81,N_2570,N_2527);
and UO_82 (O_82,N_2957,N_2981);
nand UO_83 (O_83,N_2545,N_2676);
or UO_84 (O_84,N_2720,N_2643);
or UO_85 (O_85,N_2629,N_2569);
nor UO_86 (O_86,N_2909,N_2636);
nor UO_87 (O_87,N_2810,N_2866);
and UO_88 (O_88,N_2798,N_2854);
or UO_89 (O_89,N_2631,N_2978);
nand UO_90 (O_90,N_2502,N_2583);
or UO_91 (O_91,N_2887,N_2993);
and UO_92 (O_92,N_2744,N_2823);
or UO_93 (O_93,N_2624,N_2906);
and UO_94 (O_94,N_2656,N_2626);
nor UO_95 (O_95,N_2881,N_2849);
nor UO_96 (O_96,N_2857,N_2863);
or UO_97 (O_97,N_2599,N_2862);
nor UO_98 (O_98,N_2784,N_2584);
nand UO_99 (O_99,N_2816,N_2650);
and UO_100 (O_100,N_2874,N_2555);
or UO_101 (O_101,N_2958,N_2853);
or UO_102 (O_102,N_2953,N_2528);
nor UO_103 (O_103,N_2921,N_2550);
or UO_104 (O_104,N_2609,N_2616);
xor UO_105 (O_105,N_2546,N_2664);
nor UO_106 (O_106,N_2692,N_2747);
or UO_107 (O_107,N_2535,N_2603);
or UO_108 (O_108,N_2714,N_2748);
or UO_109 (O_109,N_2571,N_2796);
and UO_110 (O_110,N_2554,N_2912);
and UO_111 (O_111,N_2547,N_2733);
nor UO_112 (O_112,N_2871,N_2776);
or UO_113 (O_113,N_2690,N_2878);
nor UO_114 (O_114,N_2700,N_2564);
nand UO_115 (O_115,N_2559,N_2946);
nor UO_116 (O_116,N_2999,N_2552);
nor UO_117 (O_117,N_2888,N_2671);
nor UO_118 (O_118,N_2991,N_2712);
and UO_119 (O_119,N_2817,N_2977);
and UO_120 (O_120,N_2769,N_2884);
nand UO_121 (O_121,N_2578,N_2667);
and UO_122 (O_122,N_2935,N_2688);
nand UO_123 (O_123,N_2778,N_2915);
nand UO_124 (O_124,N_2608,N_2828);
nor UO_125 (O_125,N_2577,N_2845);
and UO_126 (O_126,N_2880,N_2856);
nand UO_127 (O_127,N_2971,N_2727);
xnor UO_128 (O_128,N_2645,N_2719);
nor UO_129 (O_129,N_2674,N_2936);
nor UO_130 (O_130,N_2782,N_2579);
and UO_131 (O_131,N_2975,N_2581);
and UO_132 (O_132,N_2885,N_2736);
nand UO_133 (O_133,N_2792,N_2563);
nor UO_134 (O_134,N_2797,N_2610);
or UO_135 (O_135,N_2630,N_2506);
nor UO_136 (O_136,N_2898,N_2955);
nor UO_137 (O_137,N_2738,N_2956);
nor UO_138 (O_138,N_2542,N_2539);
nor UO_139 (O_139,N_2829,N_2825);
nor UO_140 (O_140,N_2757,N_2965);
and UO_141 (O_141,N_2861,N_2900);
and UO_142 (O_142,N_2974,N_2572);
nand UO_143 (O_143,N_2983,N_2998);
nor UO_144 (O_144,N_2587,N_2995);
nor UO_145 (O_145,N_2591,N_2760);
or UO_146 (O_146,N_2788,N_2634);
or UO_147 (O_147,N_2585,N_2695);
and UO_148 (O_148,N_2532,N_2870);
or UO_149 (O_149,N_2680,N_2598);
nor UO_150 (O_150,N_2619,N_2715);
nand UO_151 (O_151,N_2931,N_2689);
nor UO_152 (O_152,N_2628,N_2534);
nand UO_153 (O_153,N_2754,N_2794);
nor UO_154 (O_154,N_2850,N_2752);
and UO_155 (O_155,N_2908,N_2937);
nand UO_156 (O_156,N_2693,N_2837);
nor UO_157 (O_157,N_2709,N_2639);
nand UO_158 (O_158,N_2831,N_2858);
or UO_159 (O_159,N_2808,N_2726);
and UO_160 (O_160,N_2739,N_2602);
nor UO_161 (O_161,N_2544,N_2787);
nand UO_162 (O_162,N_2589,N_2980);
or UO_163 (O_163,N_2618,N_2723);
and UO_164 (O_164,N_2949,N_2551);
nand UO_165 (O_165,N_2836,N_2640);
nand UO_166 (O_166,N_2795,N_2565);
nor UO_167 (O_167,N_2879,N_2781);
and UO_168 (O_168,N_2929,N_2682);
nor UO_169 (O_169,N_2859,N_2560);
xnor UO_170 (O_170,N_2653,N_2681);
xnor UO_171 (O_171,N_2655,N_2745);
and UO_172 (O_172,N_2780,N_2638);
nand UO_173 (O_173,N_2773,N_2508);
nand UO_174 (O_174,N_2620,N_2821);
nand UO_175 (O_175,N_2905,N_2521);
nor UO_176 (O_176,N_2928,N_2786);
nor UO_177 (O_177,N_2641,N_2952);
and UO_178 (O_178,N_2679,N_2574);
nor UO_179 (O_179,N_2716,N_2686);
nand UO_180 (O_180,N_2901,N_2807);
and UO_181 (O_181,N_2767,N_2703);
nor UO_182 (O_182,N_2511,N_2594);
or UO_183 (O_183,N_2997,N_2510);
or UO_184 (O_184,N_2934,N_2597);
and UO_185 (O_185,N_2882,N_2730);
nand UO_186 (O_186,N_2515,N_2557);
or UO_187 (O_187,N_2672,N_2702);
and UO_188 (O_188,N_2779,N_2669);
or UO_189 (O_189,N_2553,N_2832);
or UO_190 (O_190,N_2972,N_2918);
or UO_191 (O_191,N_2996,N_2756);
nor UO_192 (O_192,N_2683,N_2970);
and UO_193 (O_193,N_2513,N_2860);
nor UO_194 (O_194,N_2729,N_2813);
nor UO_195 (O_195,N_2799,N_2663);
or UO_196 (O_196,N_2737,N_2959);
and UO_197 (O_197,N_2635,N_2839);
nand UO_198 (O_198,N_2670,N_2835);
and UO_199 (O_199,N_2711,N_2743);
nor UO_200 (O_200,N_2704,N_2948);
and UO_201 (O_201,N_2548,N_2576);
nor UO_202 (O_202,N_2633,N_2755);
nor UO_203 (O_203,N_2803,N_2994);
or UO_204 (O_204,N_2865,N_2942);
and UO_205 (O_205,N_2651,N_2531);
nor UO_206 (O_206,N_2809,N_2986);
nand UO_207 (O_207,N_2731,N_2568);
or UO_208 (O_208,N_2615,N_2600);
nor UO_209 (O_209,N_2759,N_2691);
nor UO_210 (O_210,N_2903,N_2966);
nor UO_211 (O_211,N_2876,N_2919);
nand UO_212 (O_212,N_2575,N_2509);
nand UO_213 (O_213,N_2930,N_2647);
or UO_214 (O_214,N_2646,N_2833);
xnor UO_215 (O_215,N_2632,N_2783);
nand UO_216 (O_216,N_2992,N_2873);
or UO_217 (O_217,N_2793,N_2939);
and UO_218 (O_218,N_2696,N_2891);
or UO_219 (O_219,N_2960,N_2766);
or UO_220 (O_220,N_2968,N_2875);
and UO_221 (O_221,N_2710,N_2732);
nor UO_222 (O_222,N_2847,N_2706);
and UO_223 (O_223,N_2586,N_2562);
and UO_224 (O_224,N_2938,N_2940);
nor UO_225 (O_225,N_2944,N_2889);
and UO_226 (O_226,N_2899,N_2536);
nor UO_227 (O_227,N_2666,N_2505);
nand UO_228 (O_228,N_2540,N_2735);
and UO_229 (O_229,N_2512,N_2917);
and UO_230 (O_230,N_2538,N_2625);
and UO_231 (O_231,N_2518,N_2661);
and UO_232 (O_232,N_2687,N_2964);
or UO_233 (O_233,N_2673,N_2844);
nor UO_234 (O_234,N_2812,N_2606);
and UO_235 (O_235,N_2979,N_2582);
nand UO_236 (O_236,N_2523,N_2947);
nor UO_237 (O_237,N_2678,N_2724);
nor UO_238 (O_238,N_2883,N_2699);
or UO_239 (O_239,N_2904,N_2967);
nand UO_240 (O_240,N_2894,N_2698);
nor UO_241 (O_241,N_2815,N_2895);
and UO_242 (O_242,N_2561,N_2611);
or UO_243 (O_243,N_2820,N_2750);
and UO_244 (O_244,N_2962,N_2867);
nor UO_245 (O_245,N_2785,N_2573);
and UO_246 (O_246,N_2721,N_2907);
xor UO_247 (O_247,N_2654,N_2984);
or UO_248 (O_248,N_2601,N_2811);
and UO_249 (O_249,N_2838,N_2525);
and UO_250 (O_250,N_2867,N_2595);
or UO_251 (O_251,N_2900,N_2977);
or UO_252 (O_252,N_2708,N_2584);
nor UO_253 (O_253,N_2704,N_2946);
or UO_254 (O_254,N_2542,N_2685);
nor UO_255 (O_255,N_2886,N_2866);
and UO_256 (O_256,N_2685,N_2622);
nand UO_257 (O_257,N_2966,N_2641);
nor UO_258 (O_258,N_2627,N_2540);
nor UO_259 (O_259,N_2670,N_2594);
or UO_260 (O_260,N_2921,N_2829);
xnor UO_261 (O_261,N_2514,N_2505);
or UO_262 (O_262,N_2584,N_2842);
and UO_263 (O_263,N_2681,N_2598);
nand UO_264 (O_264,N_2564,N_2715);
xnor UO_265 (O_265,N_2598,N_2630);
nor UO_266 (O_266,N_2673,N_2612);
nor UO_267 (O_267,N_2813,N_2799);
or UO_268 (O_268,N_2915,N_2590);
nor UO_269 (O_269,N_2856,N_2930);
nor UO_270 (O_270,N_2662,N_2562);
and UO_271 (O_271,N_2566,N_2925);
nand UO_272 (O_272,N_2552,N_2859);
or UO_273 (O_273,N_2644,N_2653);
and UO_274 (O_274,N_2801,N_2789);
or UO_275 (O_275,N_2784,N_2975);
nand UO_276 (O_276,N_2681,N_2900);
xnor UO_277 (O_277,N_2820,N_2735);
and UO_278 (O_278,N_2539,N_2648);
nor UO_279 (O_279,N_2504,N_2979);
nor UO_280 (O_280,N_2930,N_2996);
and UO_281 (O_281,N_2560,N_2855);
nand UO_282 (O_282,N_2946,N_2639);
or UO_283 (O_283,N_2649,N_2831);
nor UO_284 (O_284,N_2745,N_2998);
nor UO_285 (O_285,N_2535,N_2583);
and UO_286 (O_286,N_2817,N_2898);
nand UO_287 (O_287,N_2752,N_2909);
nand UO_288 (O_288,N_2642,N_2515);
and UO_289 (O_289,N_2816,N_2749);
and UO_290 (O_290,N_2596,N_2751);
nand UO_291 (O_291,N_2541,N_2708);
nand UO_292 (O_292,N_2923,N_2708);
and UO_293 (O_293,N_2690,N_2842);
nor UO_294 (O_294,N_2817,N_2768);
or UO_295 (O_295,N_2571,N_2944);
nand UO_296 (O_296,N_2606,N_2738);
nor UO_297 (O_297,N_2796,N_2875);
and UO_298 (O_298,N_2920,N_2927);
nand UO_299 (O_299,N_2594,N_2915);
nor UO_300 (O_300,N_2596,N_2787);
xor UO_301 (O_301,N_2598,N_2679);
nand UO_302 (O_302,N_2572,N_2839);
and UO_303 (O_303,N_2529,N_2603);
and UO_304 (O_304,N_2876,N_2817);
nand UO_305 (O_305,N_2817,N_2696);
nor UO_306 (O_306,N_2861,N_2656);
nand UO_307 (O_307,N_2836,N_2624);
and UO_308 (O_308,N_2603,N_2677);
or UO_309 (O_309,N_2553,N_2724);
and UO_310 (O_310,N_2791,N_2582);
or UO_311 (O_311,N_2821,N_2649);
nor UO_312 (O_312,N_2620,N_2662);
or UO_313 (O_313,N_2782,N_2990);
nor UO_314 (O_314,N_2614,N_2634);
nor UO_315 (O_315,N_2866,N_2755);
nand UO_316 (O_316,N_2882,N_2515);
or UO_317 (O_317,N_2796,N_2704);
and UO_318 (O_318,N_2774,N_2939);
or UO_319 (O_319,N_2965,N_2959);
xor UO_320 (O_320,N_2844,N_2613);
or UO_321 (O_321,N_2841,N_2948);
or UO_322 (O_322,N_2958,N_2978);
and UO_323 (O_323,N_2731,N_2911);
or UO_324 (O_324,N_2551,N_2715);
nand UO_325 (O_325,N_2743,N_2642);
and UO_326 (O_326,N_2660,N_2922);
nand UO_327 (O_327,N_2679,N_2519);
nor UO_328 (O_328,N_2900,N_2987);
and UO_329 (O_329,N_2885,N_2987);
nand UO_330 (O_330,N_2762,N_2920);
nand UO_331 (O_331,N_2791,N_2801);
or UO_332 (O_332,N_2823,N_2601);
and UO_333 (O_333,N_2641,N_2795);
nand UO_334 (O_334,N_2920,N_2588);
nand UO_335 (O_335,N_2835,N_2814);
nand UO_336 (O_336,N_2957,N_2685);
or UO_337 (O_337,N_2961,N_2630);
nor UO_338 (O_338,N_2855,N_2825);
and UO_339 (O_339,N_2651,N_2882);
and UO_340 (O_340,N_2765,N_2697);
nand UO_341 (O_341,N_2516,N_2611);
nand UO_342 (O_342,N_2773,N_2957);
nand UO_343 (O_343,N_2762,N_2773);
and UO_344 (O_344,N_2731,N_2827);
nor UO_345 (O_345,N_2733,N_2807);
nor UO_346 (O_346,N_2529,N_2826);
or UO_347 (O_347,N_2560,N_2696);
or UO_348 (O_348,N_2820,N_2543);
or UO_349 (O_349,N_2986,N_2859);
or UO_350 (O_350,N_2759,N_2628);
nor UO_351 (O_351,N_2697,N_2792);
and UO_352 (O_352,N_2536,N_2601);
or UO_353 (O_353,N_2938,N_2561);
or UO_354 (O_354,N_2763,N_2515);
nand UO_355 (O_355,N_2795,N_2878);
nand UO_356 (O_356,N_2568,N_2721);
or UO_357 (O_357,N_2752,N_2705);
and UO_358 (O_358,N_2561,N_2941);
and UO_359 (O_359,N_2739,N_2812);
nor UO_360 (O_360,N_2888,N_2769);
and UO_361 (O_361,N_2784,N_2892);
nor UO_362 (O_362,N_2727,N_2822);
nor UO_363 (O_363,N_2845,N_2721);
and UO_364 (O_364,N_2987,N_2665);
nor UO_365 (O_365,N_2797,N_2976);
and UO_366 (O_366,N_2792,N_2628);
nand UO_367 (O_367,N_2738,N_2848);
or UO_368 (O_368,N_2757,N_2877);
or UO_369 (O_369,N_2739,N_2598);
nor UO_370 (O_370,N_2796,N_2924);
or UO_371 (O_371,N_2882,N_2811);
or UO_372 (O_372,N_2713,N_2837);
or UO_373 (O_373,N_2841,N_2910);
or UO_374 (O_374,N_2747,N_2665);
xor UO_375 (O_375,N_2813,N_2572);
nor UO_376 (O_376,N_2887,N_2857);
and UO_377 (O_377,N_2695,N_2972);
nand UO_378 (O_378,N_2616,N_2543);
nor UO_379 (O_379,N_2655,N_2682);
or UO_380 (O_380,N_2738,N_2650);
nand UO_381 (O_381,N_2903,N_2676);
nor UO_382 (O_382,N_2842,N_2953);
and UO_383 (O_383,N_2743,N_2705);
nand UO_384 (O_384,N_2644,N_2791);
nand UO_385 (O_385,N_2745,N_2577);
and UO_386 (O_386,N_2555,N_2865);
or UO_387 (O_387,N_2791,N_2777);
xnor UO_388 (O_388,N_2709,N_2713);
or UO_389 (O_389,N_2970,N_2940);
nand UO_390 (O_390,N_2554,N_2784);
nand UO_391 (O_391,N_2639,N_2581);
and UO_392 (O_392,N_2978,N_2959);
nor UO_393 (O_393,N_2709,N_2996);
and UO_394 (O_394,N_2789,N_2894);
or UO_395 (O_395,N_2791,N_2686);
or UO_396 (O_396,N_2831,N_2711);
and UO_397 (O_397,N_2735,N_2509);
or UO_398 (O_398,N_2892,N_2803);
nand UO_399 (O_399,N_2542,N_2504);
nor UO_400 (O_400,N_2542,N_2725);
nand UO_401 (O_401,N_2780,N_2811);
and UO_402 (O_402,N_2992,N_2537);
nor UO_403 (O_403,N_2734,N_2643);
and UO_404 (O_404,N_2635,N_2637);
nand UO_405 (O_405,N_2863,N_2507);
nor UO_406 (O_406,N_2983,N_2990);
nor UO_407 (O_407,N_2679,N_2615);
nor UO_408 (O_408,N_2947,N_2609);
and UO_409 (O_409,N_2972,N_2810);
nor UO_410 (O_410,N_2796,N_2702);
xnor UO_411 (O_411,N_2519,N_2773);
and UO_412 (O_412,N_2507,N_2747);
nor UO_413 (O_413,N_2950,N_2638);
or UO_414 (O_414,N_2644,N_2972);
and UO_415 (O_415,N_2753,N_2709);
nand UO_416 (O_416,N_2849,N_2823);
or UO_417 (O_417,N_2873,N_2689);
and UO_418 (O_418,N_2847,N_2746);
and UO_419 (O_419,N_2675,N_2545);
or UO_420 (O_420,N_2924,N_2647);
and UO_421 (O_421,N_2839,N_2521);
or UO_422 (O_422,N_2961,N_2691);
nand UO_423 (O_423,N_2653,N_2887);
and UO_424 (O_424,N_2659,N_2865);
or UO_425 (O_425,N_2610,N_2898);
nand UO_426 (O_426,N_2930,N_2639);
nor UO_427 (O_427,N_2935,N_2945);
nand UO_428 (O_428,N_2956,N_2924);
nor UO_429 (O_429,N_2801,N_2783);
and UO_430 (O_430,N_2513,N_2560);
and UO_431 (O_431,N_2684,N_2836);
nand UO_432 (O_432,N_2561,N_2919);
or UO_433 (O_433,N_2778,N_2767);
nand UO_434 (O_434,N_2591,N_2571);
nor UO_435 (O_435,N_2541,N_2638);
or UO_436 (O_436,N_2650,N_2795);
nor UO_437 (O_437,N_2839,N_2815);
nor UO_438 (O_438,N_2944,N_2621);
nor UO_439 (O_439,N_2993,N_2741);
and UO_440 (O_440,N_2787,N_2839);
and UO_441 (O_441,N_2731,N_2975);
or UO_442 (O_442,N_2637,N_2574);
nand UO_443 (O_443,N_2679,N_2945);
and UO_444 (O_444,N_2654,N_2588);
nand UO_445 (O_445,N_2622,N_2693);
nor UO_446 (O_446,N_2774,N_2529);
nand UO_447 (O_447,N_2896,N_2918);
or UO_448 (O_448,N_2945,N_2916);
nand UO_449 (O_449,N_2697,N_2524);
nor UO_450 (O_450,N_2609,N_2506);
and UO_451 (O_451,N_2512,N_2757);
and UO_452 (O_452,N_2738,N_2540);
and UO_453 (O_453,N_2783,N_2673);
nand UO_454 (O_454,N_2942,N_2788);
or UO_455 (O_455,N_2669,N_2972);
and UO_456 (O_456,N_2562,N_2998);
nand UO_457 (O_457,N_2580,N_2791);
and UO_458 (O_458,N_2718,N_2715);
nand UO_459 (O_459,N_2664,N_2824);
and UO_460 (O_460,N_2687,N_2771);
xor UO_461 (O_461,N_2745,N_2672);
or UO_462 (O_462,N_2703,N_2903);
xnor UO_463 (O_463,N_2670,N_2812);
nor UO_464 (O_464,N_2564,N_2960);
nor UO_465 (O_465,N_2690,N_2519);
and UO_466 (O_466,N_2892,N_2635);
or UO_467 (O_467,N_2796,N_2676);
or UO_468 (O_468,N_2893,N_2501);
or UO_469 (O_469,N_2623,N_2724);
and UO_470 (O_470,N_2502,N_2537);
nand UO_471 (O_471,N_2944,N_2670);
nand UO_472 (O_472,N_2649,N_2876);
and UO_473 (O_473,N_2835,N_2594);
and UO_474 (O_474,N_2515,N_2869);
nand UO_475 (O_475,N_2548,N_2880);
and UO_476 (O_476,N_2675,N_2552);
xnor UO_477 (O_477,N_2791,N_2603);
nor UO_478 (O_478,N_2988,N_2587);
or UO_479 (O_479,N_2873,N_2669);
and UO_480 (O_480,N_2781,N_2941);
nand UO_481 (O_481,N_2929,N_2523);
and UO_482 (O_482,N_2942,N_2672);
nand UO_483 (O_483,N_2797,N_2700);
or UO_484 (O_484,N_2851,N_2800);
and UO_485 (O_485,N_2510,N_2525);
nand UO_486 (O_486,N_2730,N_2756);
or UO_487 (O_487,N_2845,N_2557);
or UO_488 (O_488,N_2732,N_2853);
nand UO_489 (O_489,N_2557,N_2801);
and UO_490 (O_490,N_2576,N_2970);
and UO_491 (O_491,N_2676,N_2571);
nor UO_492 (O_492,N_2978,N_2591);
nor UO_493 (O_493,N_2670,N_2656);
and UO_494 (O_494,N_2577,N_2564);
or UO_495 (O_495,N_2617,N_2705);
and UO_496 (O_496,N_2709,N_2943);
nand UO_497 (O_497,N_2563,N_2540);
or UO_498 (O_498,N_2531,N_2705);
nand UO_499 (O_499,N_2788,N_2989);
endmodule