module basic_500_3000_500_40_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_155,In_434);
nor U1 (N_1,In_387,In_143);
nor U2 (N_2,In_248,In_210);
or U3 (N_3,In_343,In_372);
or U4 (N_4,In_48,In_429);
xor U5 (N_5,In_162,In_287);
nor U6 (N_6,In_132,In_39);
nor U7 (N_7,In_190,In_94);
and U8 (N_8,In_67,In_159);
and U9 (N_9,In_208,In_167);
or U10 (N_10,In_425,In_64);
nor U11 (N_11,In_329,In_482);
or U12 (N_12,In_483,In_313);
nand U13 (N_13,In_129,In_395);
xnor U14 (N_14,In_336,In_135);
nor U15 (N_15,In_169,In_422);
and U16 (N_16,In_59,In_109);
or U17 (N_17,In_402,In_416);
nand U18 (N_18,In_203,In_23);
and U19 (N_19,In_347,In_229);
nor U20 (N_20,In_414,In_382);
xor U21 (N_21,In_195,In_78);
and U22 (N_22,In_241,In_199);
and U23 (N_23,In_16,In_152);
or U24 (N_24,In_185,In_219);
and U25 (N_25,In_421,In_89);
and U26 (N_26,In_456,In_243);
nand U27 (N_27,In_2,In_371);
and U28 (N_28,In_112,In_328);
xor U29 (N_29,In_299,In_377);
or U30 (N_30,In_242,In_289);
nor U31 (N_31,In_136,In_472);
or U32 (N_32,In_12,In_452);
nand U33 (N_33,In_388,In_270);
nor U34 (N_34,In_339,In_192);
xnor U35 (N_35,In_3,In_68);
nand U36 (N_36,In_357,In_80);
nand U37 (N_37,In_255,In_401);
or U38 (N_38,In_450,In_288);
xor U39 (N_39,In_120,In_107);
and U40 (N_40,In_378,In_217);
and U41 (N_41,In_392,In_22);
or U42 (N_42,In_367,In_330);
or U43 (N_43,In_295,In_264);
or U44 (N_44,In_433,In_471);
xor U45 (N_45,In_184,In_114);
nand U46 (N_46,In_305,In_215);
nor U47 (N_47,In_108,In_247);
or U48 (N_48,In_118,In_445);
nand U49 (N_49,In_117,In_87);
and U50 (N_50,In_53,In_276);
nor U51 (N_51,In_397,In_102);
and U52 (N_52,In_423,In_236);
nand U53 (N_53,In_494,In_447);
nand U54 (N_54,In_115,In_17);
and U55 (N_55,In_467,In_282);
and U56 (N_56,In_213,In_444);
or U57 (N_57,In_20,In_307);
nor U58 (N_58,In_426,In_491);
nand U59 (N_59,In_260,In_96);
and U60 (N_60,In_173,In_441);
or U61 (N_61,In_437,In_358);
nand U62 (N_62,In_151,In_325);
nand U63 (N_63,In_244,In_420);
or U64 (N_64,In_24,In_250);
nor U65 (N_65,In_498,In_5);
and U66 (N_66,In_331,In_386);
or U67 (N_67,In_166,In_235);
or U68 (N_68,In_262,In_363);
nor U69 (N_69,In_82,In_239);
nor U70 (N_70,In_227,In_431);
and U71 (N_71,In_301,In_340);
or U72 (N_72,In_318,In_15);
nand U73 (N_73,In_315,In_405);
nand U74 (N_74,In_476,In_480);
nand U75 (N_75,N_71,In_303);
nor U76 (N_76,In_164,In_19);
nand U77 (N_77,In_50,In_45);
nor U78 (N_78,In_338,N_70);
nand U79 (N_79,N_54,N_74);
or U80 (N_80,In_369,In_119);
and U81 (N_81,In_116,N_47);
or U82 (N_82,N_57,In_36);
and U83 (N_83,In_57,In_11);
nand U84 (N_84,In_179,In_234);
nor U85 (N_85,N_53,In_93);
and U86 (N_86,In_430,In_394);
nor U87 (N_87,In_281,N_32);
nand U88 (N_88,In_458,In_337);
nand U89 (N_89,In_317,N_64);
nand U90 (N_90,In_6,N_69);
nand U91 (N_91,In_165,In_137);
nand U92 (N_92,In_373,In_311);
or U93 (N_93,In_438,N_30);
nand U94 (N_94,N_55,In_261);
or U95 (N_95,N_27,N_48);
nand U96 (N_96,N_6,In_333);
nor U97 (N_97,In_150,In_344);
and U98 (N_98,N_50,In_202);
nand U99 (N_99,In_364,In_359);
and U100 (N_100,In_493,In_302);
nand U101 (N_101,In_345,N_39);
nand U102 (N_102,In_380,In_284);
and U103 (N_103,N_62,In_188);
and U104 (N_104,In_266,In_174);
nor U105 (N_105,In_322,In_465);
nor U106 (N_106,In_14,In_101);
and U107 (N_107,N_58,In_176);
or U108 (N_108,In_478,In_254);
nor U109 (N_109,In_157,In_7);
nand U110 (N_110,In_417,In_74);
nand U111 (N_111,In_449,In_454);
or U112 (N_112,In_470,In_40);
or U113 (N_113,In_198,In_273);
nor U114 (N_114,In_237,N_61);
and U115 (N_115,In_139,In_265);
or U116 (N_116,In_154,In_324);
xnor U117 (N_117,In_464,In_245);
or U118 (N_118,In_97,N_16);
nand U119 (N_119,N_45,In_221);
or U120 (N_120,In_413,In_473);
nor U121 (N_121,In_218,In_481);
nand U122 (N_122,In_246,N_2);
or U123 (N_123,In_308,In_418);
and U124 (N_124,In_396,In_0);
and U125 (N_125,N_51,In_293);
nand U126 (N_126,In_375,N_19);
or U127 (N_127,In_207,In_205);
or U128 (N_128,In_443,In_193);
nor U129 (N_129,In_403,In_103);
nor U130 (N_130,In_38,In_277);
or U131 (N_131,In_362,In_309);
or U132 (N_132,In_121,In_469);
or U133 (N_133,N_3,In_130);
nand U134 (N_134,In_495,In_9);
nand U135 (N_135,In_257,In_468);
and U136 (N_136,In_125,In_455);
and U137 (N_137,In_56,In_283);
nor U138 (N_138,In_28,In_79);
xor U139 (N_139,In_175,In_280);
nor U140 (N_140,In_335,In_351);
or U141 (N_141,N_13,In_61);
nor U142 (N_142,In_113,In_484);
and U143 (N_143,In_222,In_172);
and U144 (N_144,In_256,In_49);
nor U145 (N_145,In_487,In_342);
nor U146 (N_146,In_488,In_76);
and U147 (N_147,N_72,In_181);
nor U148 (N_148,In_85,In_326);
or U149 (N_149,N_5,In_225);
nor U150 (N_150,N_24,In_404);
nand U151 (N_151,In_408,N_100);
or U152 (N_152,In_439,In_407);
nand U153 (N_153,In_106,N_43);
and U154 (N_154,N_97,In_381);
or U155 (N_155,In_499,N_111);
nand U156 (N_156,In_354,In_486);
nand U157 (N_157,N_85,N_49);
nor U158 (N_158,N_109,N_119);
and U159 (N_159,In_156,N_67);
nor U160 (N_160,In_231,In_58);
or U161 (N_161,N_20,N_11);
and U162 (N_162,In_69,In_212);
nor U163 (N_163,In_95,In_191);
and U164 (N_164,N_141,In_238);
nand U165 (N_165,In_446,In_409);
or U166 (N_166,N_145,In_285);
nand U167 (N_167,N_137,N_91);
nand U168 (N_168,In_62,In_35);
nor U169 (N_169,In_126,In_182);
or U170 (N_170,N_84,In_83);
nand U171 (N_171,N_52,In_140);
and U172 (N_172,In_379,N_129);
nor U173 (N_173,In_389,N_14);
nand U174 (N_174,N_10,N_0);
or U175 (N_175,In_332,N_125);
nor U176 (N_176,N_138,In_296);
xor U177 (N_177,In_122,In_224);
nand U178 (N_178,N_44,In_268);
or U179 (N_179,In_63,In_314);
or U180 (N_180,N_107,In_361);
and U181 (N_181,In_91,In_310);
and U182 (N_182,N_132,N_41);
nand U183 (N_183,N_139,In_100);
nand U184 (N_184,In_460,In_42);
and U185 (N_185,In_160,N_116);
nand U186 (N_186,N_15,N_60);
nand U187 (N_187,In_233,In_13);
nand U188 (N_188,In_462,N_76);
nor U189 (N_189,In_46,N_81);
xnor U190 (N_190,N_140,In_355);
and U191 (N_191,In_259,N_143);
or U192 (N_192,N_127,In_497);
nor U193 (N_193,In_300,N_17);
or U194 (N_194,N_95,In_384);
nor U195 (N_195,In_30,In_400);
nor U196 (N_196,N_7,N_73);
nand U197 (N_197,In_75,N_128);
or U198 (N_198,In_406,In_274);
nor U199 (N_199,N_87,In_204);
and U200 (N_200,In_4,In_275);
or U201 (N_201,N_21,In_269);
nand U202 (N_202,In_294,In_70);
nand U203 (N_203,In_360,In_25);
nand U204 (N_204,In_144,In_147);
nor U205 (N_205,In_34,In_448);
and U206 (N_206,In_398,In_263);
or U207 (N_207,N_115,N_98);
nand U208 (N_208,In_327,In_319);
or U209 (N_209,In_183,In_124);
or U210 (N_210,N_103,In_290);
or U211 (N_211,In_411,N_92);
or U212 (N_212,In_435,N_123);
nand U213 (N_213,N_38,N_82);
or U214 (N_214,N_59,In_349);
nor U215 (N_215,In_92,In_211);
and U216 (N_216,N_105,In_228);
and U217 (N_217,N_136,N_68);
nor U218 (N_218,In_146,In_390);
or U219 (N_219,In_31,In_8);
nor U220 (N_220,In_393,N_89);
or U221 (N_221,In_158,In_223);
nor U222 (N_222,In_148,In_477);
or U223 (N_223,N_146,In_194);
nor U224 (N_224,In_178,In_252);
nor U225 (N_225,N_46,N_156);
or U226 (N_226,N_164,N_113);
or U227 (N_227,N_112,In_133);
nor U228 (N_228,N_65,In_312);
nor U229 (N_229,N_187,N_135);
and U230 (N_230,N_177,In_153);
or U231 (N_231,N_190,In_54);
xor U232 (N_232,N_22,N_28);
nand U233 (N_233,N_218,N_176);
and U234 (N_234,N_155,N_201);
nor U235 (N_235,N_124,In_492);
or U236 (N_236,In_86,In_321);
and U237 (N_237,In_90,N_184);
nand U238 (N_238,N_169,In_253);
nand U239 (N_239,In_127,N_161);
and U240 (N_240,In_196,In_98);
or U241 (N_241,N_86,In_415);
nor U242 (N_242,N_96,In_131);
nor U243 (N_243,N_56,N_217);
and U244 (N_244,N_178,N_206);
nor U245 (N_245,In_428,N_195);
and U246 (N_246,In_123,In_436);
and U247 (N_247,In_88,N_12);
nor U248 (N_248,N_36,In_1);
nand U249 (N_249,N_158,N_88);
or U250 (N_250,N_182,N_102);
or U251 (N_251,In_206,In_249);
and U252 (N_252,In_168,N_209);
xnor U253 (N_253,In_72,N_223);
and U254 (N_254,In_230,N_189);
nand U255 (N_255,In_99,N_34);
nor U256 (N_256,N_131,In_474);
or U257 (N_257,N_93,In_10);
and U258 (N_258,In_278,In_149);
and U259 (N_259,In_323,N_99);
nand U260 (N_260,N_200,N_142);
nand U261 (N_261,In_279,N_90);
nand U262 (N_262,N_18,N_202);
nor U263 (N_263,N_170,N_25);
and U264 (N_264,N_35,In_424);
nand U265 (N_265,N_213,N_167);
nor U266 (N_266,In_32,N_9);
or U267 (N_267,In_306,N_183);
or U268 (N_268,In_232,In_180);
nor U269 (N_269,In_316,N_29);
and U270 (N_270,In_81,In_451);
nor U271 (N_271,In_138,N_144);
and U272 (N_272,N_173,In_18);
nor U273 (N_273,In_334,In_44);
nand U274 (N_274,In_297,In_440);
nand U275 (N_275,In_356,N_151);
or U276 (N_276,In_442,N_118);
nor U277 (N_277,N_80,In_209);
nor U278 (N_278,N_4,N_207);
or U279 (N_279,N_31,In_374);
nor U280 (N_280,N_120,In_186);
nor U281 (N_281,N_211,N_175);
or U282 (N_282,N_215,In_341);
or U283 (N_283,In_128,In_427);
nor U284 (N_284,In_134,N_193);
and U285 (N_285,In_399,In_52);
or U286 (N_286,In_177,N_134);
and U287 (N_287,In_163,In_171);
xor U288 (N_288,N_185,N_122);
or U289 (N_289,N_23,In_27);
nor U290 (N_290,N_160,In_71);
or U291 (N_291,In_453,N_162);
or U292 (N_292,N_152,In_105);
and U293 (N_293,N_126,In_463);
or U294 (N_294,In_60,In_485);
nor U295 (N_295,N_174,N_165);
xnor U296 (N_296,In_33,N_33);
and U297 (N_297,N_149,N_133);
nor U298 (N_298,In_383,N_110);
or U299 (N_299,N_101,In_189);
nand U300 (N_300,In_346,In_466);
and U301 (N_301,N_299,N_150);
and U302 (N_302,In_479,N_194);
and U303 (N_303,N_83,N_292);
and U304 (N_304,In_370,N_220);
or U305 (N_305,In_286,In_197);
or U306 (N_306,N_256,N_280);
and U307 (N_307,N_245,N_216);
nand U308 (N_308,N_237,N_233);
or U309 (N_309,N_269,N_232);
nor U310 (N_310,N_186,N_121);
nor U311 (N_311,N_171,N_261);
xor U312 (N_312,N_253,N_226);
nor U313 (N_313,N_264,N_208);
or U314 (N_314,N_108,In_170);
nor U315 (N_315,N_249,In_366);
and U316 (N_316,N_204,N_288);
nor U317 (N_317,N_130,N_147);
nand U318 (N_318,In_368,N_242);
nor U319 (N_319,N_248,N_77);
nor U320 (N_320,N_63,In_489);
nand U321 (N_321,N_244,In_240);
or U322 (N_322,N_172,In_267);
and U323 (N_323,N_279,N_66);
nor U324 (N_324,N_234,In_187);
and U325 (N_325,N_79,In_55);
and U326 (N_326,In_141,N_205);
nor U327 (N_327,N_236,In_21);
and U328 (N_328,N_210,In_110);
or U329 (N_329,In_461,N_168);
nand U330 (N_330,N_262,N_243);
and U331 (N_331,In_73,N_94);
and U332 (N_332,N_114,In_200);
nor U333 (N_333,N_106,In_272);
and U334 (N_334,N_228,In_216);
or U335 (N_335,N_286,In_41);
and U336 (N_336,N_276,N_199);
nand U337 (N_337,In_271,N_8);
nor U338 (N_338,In_490,N_37);
or U339 (N_339,N_247,In_419);
xnor U340 (N_340,N_297,In_251);
nor U341 (N_341,N_246,In_385);
nand U342 (N_342,In_142,N_278);
and U343 (N_343,N_273,N_296);
xnor U344 (N_344,N_231,In_47);
xnor U345 (N_345,N_153,In_459);
or U346 (N_346,In_432,N_75);
nand U347 (N_347,N_267,N_42);
nor U348 (N_348,N_166,N_1);
and U349 (N_349,N_212,In_26);
or U350 (N_350,N_257,In_292);
nand U351 (N_351,N_157,N_260);
and U352 (N_352,N_241,In_77);
and U353 (N_353,N_289,N_203);
nand U354 (N_354,N_192,N_274);
nor U355 (N_355,N_290,N_258);
and U356 (N_356,N_117,N_293);
nand U357 (N_357,In_353,In_226);
or U358 (N_358,N_40,In_475);
nor U359 (N_359,In_84,In_29);
nand U360 (N_360,N_298,N_263);
and U361 (N_361,N_285,In_304);
and U362 (N_362,In_258,N_282);
nor U363 (N_363,N_271,N_287);
and U364 (N_364,N_188,N_214);
nor U365 (N_365,In_320,N_222);
xnor U366 (N_366,N_180,In_412);
or U367 (N_367,In_220,N_224);
or U368 (N_368,N_148,N_230);
and U369 (N_369,In_365,In_111);
nand U370 (N_370,N_191,N_238);
nand U371 (N_371,In_410,N_219);
and U372 (N_372,In_51,In_145);
nor U373 (N_373,N_259,In_37);
nand U374 (N_374,N_179,In_350);
and U375 (N_375,N_304,N_357);
or U376 (N_376,N_338,N_359);
and U377 (N_377,N_348,N_342);
and U378 (N_378,N_368,N_239);
nor U379 (N_379,N_333,N_104);
or U380 (N_380,N_198,N_369);
and U381 (N_381,N_154,N_331);
nor U382 (N_382,N_309,N_307);
and U383 (N_383,N_318,N_374);
and U384 (N_384,N_163,N_328);
nor U385 (N_385,In_496,N_302);
and U386 (N_386,N_353,N_330);
nor U387 (N_387,N_364,In_298);
and U388 (N_388,N_347,In_43);
or U389 (N_389,N_326,N_345);
and U390 (N_390,N_365,N_324);
nand U391 (N_391,N_341,N_314);
nor U392 (N_392,N_337,In_376);
or U393 (N_393,N_306,N_356);
nor U394 (N_394,N_350,N_362);
nor U395 (N_395,N_294,N_277);
and U396 (N_396,N_336,N_311);
or U397 (N_397,N_308,N_367);
nor U398 (N_398,N_315,N_251);
and U399 (N_399,N_295,N_358);
or U400 (N_400,N_339,N_351);
and U401 (N_401,N_361,N_275);
or U402 (N_402,In_104,N_235);
nand U403 (N_403,N_363,N_229);
or U404 (N_404,N_227,N_323);
and U405 (N_405,N_252,N_312);
nor U406 (N_406,N_319,N_334);
and U407 (N_407,N_321,N_250);
and U408 (N_408,N_343,N_197);
nor U409 (N_409,In_391,N_320);
nand U410 (N_410,N_329,N_322);
nor U411 (N_411,N_300,N_281);
and U412 (N_412,N_355,N_372);
or U413 (N_413,N_332,N_316);
nor U414 (N_414,In_214,N_268);
or U415 (N_415,N_283,N_327);
and U416 (N_416,N_346,N_284);
or U417 (N_417,N_225,N_317);
and U418 (N_418,In_352,In_65);
or U419 (N_419,N_373,In_66);
nor U420 (N_420,In_348,N_255);
nand U421 (N_421,N_310,N_266);
and U422 (N_422,N_240,N_371);
nor U423 (N_423,N_272,N_196);
or U424 (N_424,N_344,N_360);
nor U425 (N_425,N_335,In_457);
nand U426 (N_426,N_305,N_352);
nor U427 (N_427,N_340,N_291);
or U428 (N_428,N_254,In_161);
nor U429 (N_429,In_291,N_78);
and U430 (N_430,N_26,N_349);
nor U431 (N_431,N_265,N_370);
or U432 (N_432,N_313,N_303);
nand U433 (N_433,N_221,N_366);
or U434 (N_434,N_181,N_159);
nor U435 (N_435,N_301,N_270);
xor U436 (N_436,N_325,In_201);
and U437 (N_437,N_354,N_311);
nand U438 (N_438,In_496,N_314);
nor U439 (N_439,N_26,N_347);
nand U440 (N_440,N_356,N_335);
nand U441 (N_441,N_181,N_250);
and U442 (N_442,N_227,N_311);
and U443 (N_443,N_368,N_284);
and U444 (N_444,N_360,In_391);
nand U445 (N_445,In_201,N_181);
nand U446 (N_446,N_268,N_354);
xor U447 (N_447,N_159,N_330);
xnor U448 (N_448,In_214,N_334);
or U449 (N_449,N_331,N_250);
or U450 (N_450,N_434,N_411);
nor U451 (N_451,N_391,N_415);
or U452 (N_452,N_412,N_389);
xnor U453 (N_453,N_390,N_438);
nand U454 (N_454,N_429,N_413);
nor U455 (N_455,N_401,N_435);
nand U456 (N_456,N_442,N_376);
or U457 (N_457,N_430,N_431);
and U458 (N_458,N_439,N_449);
and U459 (N_459,N_395,N_425);
nand U460 (N_460,N_433,N_398);
nor U461 (N_461,N_407,N_375);
nand U462 (N_462,N_381,N_419);
and U463 (N_463,N_383,N_378);
and U464 (N_464,N_394,N_443);
nand U465 (N_465,N_416,N_428);
and U466 (N_466,N_446,N_385);
nor U467 (N_467,N_377,N_393);
nand U468 (N_468,N_423,N_382);
nand U469 (N_469,N_399,N_386);
nand U470 (N_470,N_400,N_380);
or U471 (N_471,N_422,N_440);
nand U472 (N_472,N_404,N_437);
or U473 (N_473,N_445,N_426);
and U474 (N_474,N_387,N_432);
or U475 (N_475,N_441,N_410);
nor U476 (N_476,N_420,N_392);
or U477 (N_477,N_421,N_397);
xnor U478 (N_478,N_414,N_448);
nor U479 (N_479,N_436,N_447);
and U480 (N_480,N_402,N_417);
nand U481 (N_481,N_409,N_396);
and U482 (N_482,N_379,N_405);
xnor U483 (N_483,N_408,N_427);
nand U484 (N_484,N_418,N_403);
or U485 (N_485,N_384,N_406);
nand U486 (N_486,N_388,N_444);
nand U487 (N_487,N_424,N_440);
and U488 (N_488,N_394,N_408);
or U489 (N_489,N_416,N_440);
and U490 (N_490,N_389,N_434);
nor U491 (N_491,N_449,N_444);
and U492 (N_492,N_400,N_390);
nor U493 (N_493,N_386,N_411);
nand U494 (N_494,N_387,N_437);
or U495 (N_495,N_416,N_433);
or U496 (N_496,N_434,N_383);
and U497 (N_497,N_425,N_391);
or U498 (N_498,N_432,N_404);
nand U499 (N_499,N_381,N_440);
nor U500 (N_500,N_443,N_400);
nand U501 (N_501,N_429,N_410);
nor U502 (N_502,N_382,N_399);
nor U503 (N_503,N_407,N_390);
nand U504 (N_504,N_397,N_381);
and U505 (N_505,N_396,N_406);
or U506 (N_506,N_448,N_400);
and U507 (N_507,N_442,N_426);
and U508 (N_508,N_381,N_411);
nor U509 (N_509,N_419,N_436);
nor U510 (N_510,N_411,N_379);
nand U511 (N_511,N_397,N_425);
nand U512 (N_512,N_435,N_394);
nand U513 (N_513,N_385,N_380);
or U514 (N_514,N_432,N_376);
and U515 (N_515,N_449,N_417);
xor U516 (N_516,N_402,N_446);
or U517 (N_517,N_388,N_439);
and U518 (N_518,N_388,N_420);
nand U519 (N_519,N_404,N_398);
or U520 (N_520,N_404,N_382);
or U521 (N_521,N_421,N_401);
nand U522 (N_522,N_377,N_426);
nor U523 (N_523,N_385,N_429);
and U524 (N_524,N_411,N_433);
or U525 (N_525,N_518,N_504);
and U526 (N_526,N_485,N_500);
or U527 (N_527,N_490,N_495);
or U528 (N_528,N_510,N_469);
and U529 (N_529,N_522,N_466);
nor U530 (N_530,N_521,N_515);
and U531 (N_531,N_451,N_452);
and U532 (N_532,N_472,N_476);
and U533 (N_533,N_470,N_458);
or U534 (N_534,N_475,N_491);
and U535 (N_535,N_511,N_507);
nor U536 (N_536,N_487,N_513);
xnor U537 (N_537,N_523,N_497);
or U538 (N_538,N_514,N_508);
nand U539 (N_539,N_498,N_501);
nand U540 (N_540,N_492,N_474);
nand U541 (N_541,N_496,N_465);
nand U542 (N_542,N_489,N_471);
or U543 (N_543,N_524,N_479);
or U544 (N_544,N_506,N_482);
nand U545 (N_545,N_464,N_454);
nand U546 (N_546,N_459,N_509);
or U547 (N_547,N_462,N_486);
or U548 (N_548,N_457,N_519);
nand U549 (N_549,N_480,N_481);
nor U550 (N_550,N_512,N_484);
or U551 (N_551,N_463,N_468);
or U552 (N_552,N_450,N_494);
and U553 (N_553,N_520,N_516);
and U554 (N_554,N_517,N_493);
and U555 (N_555,N_502,N_455);
nand U556 (N_556,N_478,N_453);
nand U557 (N_557,N_488,N_503);
nand U558 (N_558,N_499,N_460);
nand U559 (N_559,N_483,N_467);
nand U560 (N_560,N_477,N_461);
and U561 (N_561,N_505,N_456);
nor U562 (N_562,N_473,N_455);
and U563 (N_563,N_511,N_477);
and U564 (N_564,N_486,N_475);
xor U565 (N_565,N_455,N_462);
or U566 (N_566,N_453,N_500);
nor U567 (N_567,N_466,N_523);
and U568 (N_568,N_474,N_464);
xor U569 (N_569,N_470,N_520);
nor U570 (N_570,N_473,N_523);
nor U571 (N_571,N_475,N_492);
or U572 (N_572,N_473,N_487);
nor U573 (N_573,N_488,N_523);
and U574 (N_574,N_489,N_524);
and U575 (N_575,N_513,N_507);
or U576 (N_576,N_499,N_482);
nor U577 (N_577,N_458,N_492);
xor U578 (N_578,N_473,N_515);
nor U579 (N_579,N_486,N_468);
nand U580 (N_580,N_515,N_498);
or U581 (N_581,N_478,N_524);
nand U582 (N_582,N_520,N_478);
nor U583 (N_583,N_477,N_485);
and U584 (N_584,N_469,N_471);
or U585 (N_585,N_460,N_477);
and U586 (N_586,N_466,N_455);
nor U587 (N_587,N_523,N_505);
xnor U588 (N_588,N_488,N_485);
nor U589 (N_589,N_524,N_493);
or U590 (N_590,N_480,N_494);
and U591 (N_591,N_491,N_476);
nand U592 (N_592,N_492,N_520);
xnor U593 (N_593,N_517,N_472);
and U594 (N_594,N_451,N_502);
and U595 (N_595,N_497,N_463);
or U596 (N_596,N_496,N_497);
or U597 (N_597,N_494,N_451);
or U598 (N_598,N_507,N_519);
nand U599 (N_599,N_472,N_501);
and U600 (N_600,N_577,N_548);
and U601 (N_601,N_535,N_543);
nor U602 (N_602,N_573,N_594);
nor U603 (N_603,N_539,N_590);
nand U604 (N_604,N_560,N_588);
nand U605 (N_605,N_586,N_528);
or U606 (N_606,N_592,N_547);
and U607 (N_607,N_584,N_558);
nand U608 (N_608,N_541,N_553);
or U609 (N_609,N_538,N_589);
nand U610 (N_610,N_565,N_574);
or U611 (N_611,N_531,N_559);
nand U612 (N_612,N_537,N_575);
nand U613 (N_613,N_578,N_534);
or U614 (N_614,N_568,N_566);
nand U615 (N_615,N_597,N_525);
and U616 (N_616,N_598,N_576);
and U617 (N_617,N_540,N_582);
nand U618 (N_618,N_571,N_587);
nand U619 (N_619,N_529,N_536);
and U620 (N_620,N_533,N_555);
nor U621 (N_621,N_549,N_561);
and U622 (N_622,N_550,N_572);
or U623 (N_623,N_581,N_593);
nand U624 (N_624,N_532,N_526);
nor U625 (N_625,N_564,N_580);
and U626 (N_626,N_579,N_552);
nor U627 (N_627,N_546,N_591);
nand U628 (N_628,N_562,N_567);
or U629 (N_629,N_595,N_542);
nand U630 (N_630,N_556,N_557);
nor U631 (N_631,N_569,N_545);
xnor U632 (N_632,N_544,N_527);
nand U633 (N_633,N_554,N_585);
nand U634 (N_634,N_551,N_596);
and U635 (N_635,N_570,N_583);
and U636 (N_636,N_530,N_563);
nor U637 (N_637,N_599,N_565);
or U638 (N_638,N_591,N_530);
and U639 (N_639,N_530,N_537);
nor U640 (N_640,N_566,N_569);
nand U641 (N_641,N_580,N_544);
nand U642 (N_642,N_534,N_555);
nand U643 (N_643,N_548,N_531);
nand U644 (N_644,N_569,N_529);
nor U645 (N_645,N_556,N_584);
nand U646 (N_646,N_557,N_567);
or U647 (N_647,N_575,N_540);
nor U648 (N_648,N_542,N_583);
nor U649 (N_649,N_565,N_533);
nor U650 (N_650,N_585,N_532);
nor U651 (N_651,N_583,N_557);
and U652 (N_652,N_542,N_528);
or U653 (N_653,N_597,N_579);
nand U654 (N_654,N_588,N_535);
or U655 (N_655,N_535,N_571);
and U656 (N_656,N_569,N_543);
nand U657 (N_657,N_574,N_586);
or U658 (N_658,N_545,N_535);
or U659 (N_659,N_543,N_544);
nor U660 (N_660,N_548,N_584);
or U661 (N_661,N_551,N_582);
or U662 (N_662,N_584,N_572);
nand U663 (N_663,N_572,N_592);
nand U664 (N_664,N_554,N_541);
nor U665 (N_665,N_545,N_565);
nand U666 (N_666,N_538,N_561);
nor U667 (N_667,N_598,N_549);
or U668 (N_668,N_564,N_542);
or U669 (N_669,N_593,N_552);
and U670 (N_670,N_567,N_548);
or U671 (N_671,N_533,N_553);
and U672 (N_672,N_590,N_576);
nand U673 (N_673,N_527,N_535);
nor U674 (N_674,N_597,N_560);
nand U675 (N_675,N_619,N_647);
nor U676 (N_676,N_636,N_614);
or U677 (N_677,N_602,N_643);
and U678 (N_678,N_651,N_655);
and U679 (N_679,N_609,N_673);
and U680 (N_680,N_633,N_670);
or U681 (N_681,N_665,N_601);
nor U682 (N_682,N_634,N_659);
nor U683 (N_683,N_626,N_657);
and U684 (N_684,N_621,N_666);
xnor U685 (N_685,N_623,N_644);
or U686 (N_686,N_654,N_606);
or U687 (N_687,N_618,N_630);
or U688 (N_688,N_620,N_664);
or U689 (N_689,N_650,N_611);
nand U690 (N_690,N_638,N_635);
and U691 (N_691,N_669,N_607);
nand U692 (N_692,N_649,N_631);
or U693 (N_693,N_674,N_604);
or U694 (N_694,N_615,N_622);
and U695 (N_695,N_629,N_616);
nor U696 (N_696,N_662,N_656);
or U697 (N_697,N_668,N_642);
and U698 (N_698,N_608,N_667);
nand U699 (N_699,N_660,N_640);
nor U700 (N_700,N_627,N_603);
nand U701 (N_701,N_645,N_652);
nor U702 (N_702,N_639,N_605);
xor U703 (N_703,N_637,N_612);
nand U704 (N_704,N_641,N_671);
and U705 (N_705,N_600,N_613);
or U706 (N_706,N_610,N_663);
or U707 (N_707,N_672,N_632);
or U708 (N_708,N_617,N_661);
nor U709 (N_709,N_648,N_625);
or U710 (N_710,N_658,N_646);
and U711 (N_711,N_653,N_624);
nor U712 (N_712,N_628,N_609);
nor U713 (N_713,N_604,N_601);
or U714 (N_714,N_632,N_641);
nor U715 (N_715,N_671,N_626);
nand U716 (N_716,N_673,N_643);
and U717 (N_717,N_603,N_640);
nand U718 (N_718,N_649,N_635);
nor U719 (N_719,N_611,N_662);
nor U720 (N_720,N_607,N_605);
or U721 (N_721,N_652,N_651);
and U722 (N_722,N_623,N_645);
nor U723 (N_723,N_611,N_601);
or U724 (N_724,N_613,N_648);
nand U725 (N_725,N_651,N_663);
or U726 (N_726,N_601,N_620);
nand U727 (N_727,N_661,N_626);
and U728 (N_728,N_657,N_618);
nand U729 (N_729,N_615,N_614);
nand U730 (N_730,N_662,N_623);
and U731 (N_731,N_643,N_669);
or U732 (N_732,N_660,N_644);
or U733 (N_733,N_610,N_646);
nand U734 (N_734,N_631,N_602);
and U735 (N_735,N_621,N_606);
and U736 (N_736,N_639,N_632);
and U737 (N_737,N_614,N_648);
xor U738 (N_738,N_670,N_610);
nand U739 (N_739,N_600,N_624);
nor U740 (N_740,N_663,N_630);
nand U741 (N_741,N_652,N_620);
and U742 (N_742,N_648,N_607);
and U743 (N_743,N_629,N_651);
xor U744 (N_744,N_618,N_606);
and U745 (N_745,N_636,N_631);
or U746 (N_746,N_600,N_637);
nor U747 (N_747,N_660,N_670);
nor U748 (N_748,N_656,N_668);
and U749 (N_749,N_609,N_674);
or U750 (N_750,N_686,N_688);
xnor U751 (N_751,N_685,N_749);
nor U752 (N_752,N_713,N_690);
or U753 (N_753,N_716,N_687);
xnor U754 (N_754,N_703,N_731);
nand U755 (N_755,N_724,N_683);
and U756 (N_756,N_745,N_719);
xor U757 (N_757,N_722,N_725);
nand U758 (N_758,N_698,N_741);
nand U759 (N_759,N_693,N_718);
nand U760 (N_760,N_721,N_677);
nor U761 (N_761,N_712,N_699);
or U762 (N_762,N_729,N_696);
nand U763 (N_763,N_678,N_694);
nor U764 (N_764,N_710,N_675);
nor U765 (N_765,N_744,N_717);
and U766 (N_766,N_684,N_730);
or U767 (N_767,N_702,N_746);
nand U768 (N_768,N_707,N_728);
nor U769 (N_769,N_680,N_735);
or U770 (N_770,N_739,N_708);
or U771 (N_771,N_727,N_692);
nand U772 (N_772,N_711,N_679);
nor U773 (N_773,N_714,N_709);
xor U774 (N_774,N_732,N_697);
nor U775 (N_775,N_691,N_736);
nor U776 (N_776,N_747,N_700);
and U777 (N_777,N_742,N_734);
nor U778 (N_778,N_715,N_733);
nand U779 (N_779,N_705,N_704);
or U780 (N_780,N_681,N_720);
and U781 (N_781,N_726,N_738);
nand U782 (N_782,N_706,N_748);
nor U783 (N_783,N_701,N_682);
or U784 (N_784,N_689,N_743);
nand U785 (N_785,N_723,N_737);
xor U786 (N_786,N_676,N_695);
or U787 (N_787,N_740,N_697);
nor U788 (N_788,N_678,N_711);
and U789 (N_789,N_693,N_741);
or U790 (N_790,N_694,N_747);
and U791 (N_791,N_677,N_740);
or U792 (N_792,N_702,N_686);
or U793 (N_793,N_680,N_679);
or U794 (N_794,N_710,N_697);
nand U795 (N_795,N_677,N_718);
nand U796 (N_796,N_694,N_679);
nor U797 (N_797,N_726,N_682);
and U798 (N_798,N_713,N_675);
and U799 (N_799,N_676,N_715);
and U800 (N_800,N_712,N_749);
or U801 (N_801,N_725,N_721);
and U802 (N_802,N_689,N_747);
or U803 (N_803,N_741,N_737);
or U804 (N_804,N_703,N_736);
or U805 (N_805,N_710,N_690);
or U806 (N_806,N_695,N_720);
or U807 (N_807,N_705,N_699);
nand U808 (N_808,N_699,N_743);
and U809 (N_809,N_732,N_694);
nand U810 (N_810,N_696,N_705);
nand U811 (N_811,N_731,N_707);
nor U812 (N_812,N_718,N_733);
or U813 (N_813,N_744,N_689);
and U814 (N_814,N_675,N_677);
and U815 (N_815,N_706,N_685);
nor U816 (N_816,N_688,N_720);
or U817 (N_817,N_728,N_745);
nor U818 (N_818,N_703,N_713);
or U819 (N_819,N_678,N_698);
xor U820 (N_820,N_715,N_731);
nor U821 (N_821,N_687,N_728);
nand U822 (N_822,N_692,N_690);
or U823 (N_823,N_707,N_732);
and U824 (N_824,N_707,N_681);
and U825 (N_825,N_815,N_808);
nand U826 (N_826,N_759,N_804);
nor U827 (N_827,N_807,N_810);
or U828 (N_828,N_820,N_764);
or U829 (N_829,N_781,N_770);
nor U830 (N_830,N_774,N_814);
and U831 (N_831,N_762,N_803);
nand U832 (N_832,N_809,N_817);
xnor U833 (N_833,N_824,N_750);
and U834 (N_834,N_812,N_822);
nor U835 (N_835,N_773,N_772);
and U836 (N_836,N_768,N_763);
nor U837 (N_837,N_754,N_811);
and U838 (N_838,N_771,N_756);
and U839 (N_839,N_752,N_823);
and U840 (N_840,N_799,N_805);
nand U841 (N_841,N_813,N_775);
nand U842 (N_842,N_789,N_816);
and U843 (N_843,N_751,N_765);
or U844 (N_844,N_821,N_802);
and U845 (N_845,N_787,N_794);
nor U846 (N_846,N_798,N_753);
nand U847 (N_847,N_778,N_806);
and U848 (N_848,N_790,N_797);
nand U849 (N_849,N_791,N_755);
or U850 (N_850,N_780,N_819);
or U851 (N_851,N_796,N_788);
or U852 (N_852,N_795,N_784);
nand U853 (N_853,N_769,N_779);
xor U854 (N_854,N_757,N_786);
or U855 (N_855,N_818,N_761);
xor U856 (N_856,N_758,N_760);
and U857 (N_857,N_783,N_776);
or U858 (N_858,N_782,N_785);
and U859 (N_859,N_793,N_800);
and U860 (N_860,N_777,N_792);
nand U861 (N_861,N_801,N_766);
nand U862 (N_862,N_767,N_820);
or U863 (N_863,N_773,N_808);
xor U864 (N_864,N_797,N_803);
nor U865 (N_865,N_792,N_819);
and U866 (N_866,N_820,N_754);
xnor U867 (N_867,N_805,N_792);
or U868 (N_868,N_793,N_750);
nand U869 (N_869,N_790,N_800);
nor U870 (N_870,N_808,N_754);
nand U871 (N_871,N_763,N_800);
nor U872 (N_872,N_773,N_792);
or U873 (N_873,N_816,N_762);
nor U874 (N_874,N_798,N_795);
nor U875 (N_875,N_784,N_807);
or U876 (N_876,N_760,N_805);
and U877 (N_877,N_805,N_783);
nand U878 (N_878,N_806,N_784);
and U879 (N_879,N_750,N_803);
or U880 (N_880,N_802,N_771);
nor U881 (N_881,N_787,N_795);
nor U882 (N_882,N_772,N_818);
or U883 (N_883,N_755,N_773);
and U884 (N_884,N_823,N_765);
nand U885 (N_885,N_783,N_770);
nor U886 (N_886,N_764,N_757);
xor U887 (N_887,N_798,N_804);
nor U888 (N_888,N_812,N_771);
and U889 (N_889,N_809,N_794);
or U890 (N_890,N_803,N_784);
and U891 (N_891,N_822,N_767);
nor U892 (N_892,N_803,N_824);
nor U893 (N_893,N_809,N_757);
or U894 (N_894,N_792,N_764);
nand U895 (N_895,N_766,N_771);
and U896 (N_896,N_776,N_821);
and U897 (N_897,N_759,N_755);
nand U898 (N_898,N_767,N_766);
or U899 (N_899,N_755,N_785);
or U900 (N_900,N_864,N_832);
nand U901 (N_901,N_835,N_855);
nand U902 (N_902,N_860,N_841);
and U903 (N_903,N_880,N_872);
and U904 (N_904,N_838,N_857);
and U905 (N_905,N_851,N_863);
nor U906 (N_906,N_874,N_856);
nand U907 (N_907,N_870,N_848);
nand U908 (N_908,N_891,N_879);
nand U909 (N_909,N_825,N_829);
xnor U910 (N_910,N_868,N_887);
and U911 (N_911,N_896,N_840);
or U912 (N_912,N_850,N_865);
nand U913 (N_913,N_888,N_826);
nand U914 (N_914,N_845,N_852);
nand U915 (N_915,N_861,N_889);
nand U916 (N_916,N_831,N_828);
or U917 (N_917,N_847,N_859);
nand U918 (N_918,N_843,N_890);
nand U919 (N_919,N_882,N_899);
xor U920 (N_920,N_892,N_886);
or U921 (N_921,N_877,N_869);
or U922 (N_922,N_834,N_883);
nor U923 (N_923,N_895,N_875);
or U924 (N_924,N_878,N_884);
nor U925 (N_925,N_839,N_894);
or U926 (N_926,N_871,N_862);
nand U927 (N_927,N_897,N_842);
xor U928 (N_928,N_866,N_836);
nor U929 (N_929,N_849,N_853);
or U930 (N_930,N_867,N_854);
nor U931 (N_931,N_830,N_873);
and U932 (N_932,N_893,N_876);
nor U933 (N_933,N_885,N_827);
nor U934 (N_934,N_881,N_833);
nor U935 (N_935,N_858,N_844);
nand U936 (N_936,N_898,N_846);
nor U937 (N_937,N_837,N_870);
and U938 (N_938,N_839,N_860);
or U939 (N_939,N_893,N_883);
or U940 (N_940,N_841,N_858);
or U941 (N_941,N_829,N_863);
or U942 (N_942,N_849,N_829);
xor U943 (N_943,N_892,N_838);
nor U944 (N_944,N_848,N_893);
nor U945 (N_945,N_876,N_859);
nor U946 (N_946,N_844,N_825);
and U947 (N_947,N_830,N_827);
nor U948 (N_948,N_857,N_886);
or U949 (N_949,N_851,N_886);
nor U950 (N_950,N_840,N_878);
nand U951 (N_951,N_880,N_843);
nand U952 (N_952,N_862,N_835);
nand U953 (N_953,N_842,N_838);
nand U954 (N_954,N_848,N_857);
and U955 (N_955,N_836,N_885);
nand U956 (N_956,N_836,N_877);
nor U957 (N_957,N_885,N_879);
and U958 (N_958,N_854,N_889);
or U959 (N_959,N_840,N_860);
nand U960 (N_960,N_859,N_870);
nor U961 (N_961,N_892,N_836);
and U962 (N_962,N_877,N_850);
nor U963 (N_963,N_825,N_863);
nand U964 (N_964,N_864,N_865);
and U965 (N_965,N_837,N_896);
and U966 (N_966,N_889,N_836);
nor U967 (N_967,N_876,N_849);
nand U968 (N_968,N_892,N_827);
and U969 (N_969,N_879,N_871);
or U970 (N_970,N_852,N_853);
nor U971 (N_971,N_874,N_891);
or U972 (N_972,N_834,N_884);
or U973 (N_973,N_875,N_834);
or U974 (N_974,N_842,N_899);
nand U975 (N_975,N_953,N_906);
nor U976 (N_976,N_973,N_964);
or U977 (N_977,N_928,N_969);
nand U978 (N_978,N_901,N_929);
nor U979 (N_979,N_965,N_954);
or U980 (N_980,N_956,N_925);
or U981 (N_981,N_900,N_907);
or U982 (N_982,N_947,N_912);
xor U983 (N_983,N_948,N_968);
nor U984 (N_984,N_904,N_913);
or U985 (N_985,N_905,N_974);
or U986 (N_986,N_917,N_916);
or U987 (N_987,N_932,N_931);
and U988 (N_988,N_940,N_911);
and U989 (N_989,N_927,N_923);
nor U990 (N_990,N_937,N_920);
and U991 (N_991,N_955,N_935);
or U992 (N_992,N_926,N_959);
or U993 (N_993,N_924,N_944);
and U994 (N_994,N_930,N_958);
nand U995 (N_995,N_952,N_949);
and U996 (N_996,N_941,N_942);
nor U997 (N_997,N_972,N_914);
xnor U998 (N_998,N_915,N_963);
or U999 (N_999,N_943,N_903);
nand U1000 (N_1000,N_962,N_967);
or U1001 (N_1001,N_936,N_946);
or U1002 (N_1002,N_957,N_909);
or U1003 (N_1003,N_939,N_966);
or U1004 (N_1004,N_908,N_938);
or U1005 (N_1005,N_921,N_933);
nand U1006 (N_1006,N_950,N_961);
and U1007 (N_1007,N_970,N_945);
nor U1008 (N_1008,N_960,N_910);
and U1009 (N_1009,N_918,N_971);
nor U1010 (N_1010,N_919,N_951);
nand U1011 (N_1011,N_902,N_922);
and U1012 (N_1012,N_934,N_919);
and U1013 (N_1013,N_939,N_968);
nand U1014 (N_1014,N_921,N_922);
nand U1015 (N_1015,N_932,N_968);
xor U1016 (N_1016,N_946,N_970);
nor U1017 (N_1017,N_919,N_928);
nor U1018 (N_1018,N_911,N_948);
xnor U1019 (N_1019,N_974,N_934);
and U1020 (N_1020,N_939,N_928);
or U1021 (N_1021,N_950,N_911);
and U1022 (N_1022,N_923,N_961);
nor U1023 (N_1023,N_921,N_957);
or U1024 (N_1024,N_950,N_944);
or U1025 (N_1025,N_911,N_942);
and U1026 (N_1026,N_906,N_939);
nor U1027 (N_1027,N_908,N_931);
nor U1028 (N_1028,N_973,N_904);
or U1029 (N_1029,N_956,N_906);
nand U1030 (N_1030,N_928,N_904);
or U1031 (N_1031,N_917,N_973);
and U1032 (N_1032,N_934,N_964);
and U1033 (N_1033,N_930,N_913);
or U1034 (N_1034,N_921,N_910);
nor U1035 (N_1035,N_948,N_963);
nor U1036 (N_1036,N_955,N_948);
or U1037 (N_1037,N_942,N_954);
nor U1038 (N_1038,N_956,N_930);
nand U1039 (N_1039,N_913,N_946);
nor U1040 (N_1040,N_953,N_962);
and U1041 (N_1041,N_917,N_957);
or U1042 (N_1042,N_927,N_931);
nand U1043 (N_1043,N_911,N_932);
nor U1044 (N_1044,N_958,N_919);
and U1045 (N_1045,N_913,N_909);
or U1046 (N_1046,N_938,N_953);
nor U1047 (N_1047,N_901,N_963);
nand U1048 (N_1048,N_947,N_940);
or U1049 (N_1049,N_910,N_919);
and U1050 (N_1050,N_1030,N_975);
and U1051 (N_1051,N_1000,N_1038);
or U1052 (N_1052,N_1039,N_1033);
nor U1053 (N_1053,N_1008,N_985);
or U1054 (N_1054,N_1017,N_1028);
and U1055 (N_1055,N_1025,N_1009);
nand U1056 (N_1056,N_980,N_1010);
and U1057 (N_1057,N_1029,N_988);
or U1058 (N_1058,N_1031,N_1004);
and U1059 (N_1059,N_1023,N_976);
nor U1060 (N_1060,N_986,N_996);
nor U1061 (N_1061,N_1007,N_1001);
nor U1062 (N_1062,N_1014,N_992);
nor U1063 (N_1063,N_995,N_1013);
and U1064 (N_1064,N_1040,N_1042);
and U1065 (N_1065,N_990,N_1021);
and U1066 (N_1066,N_1045,N_998);
nand U1067 (N_1067,N_1026,N_982);
nor U1068 (N_1068,N_1036,N_1044);
nor U1069 (N_1069,N_1002,N_1018);
nor U1070 (N_1070,N_983,N_1041);
nor U1071 (N_1071,N_1024,N_1046);
nand U1072 (N_1072,N_1047,N_981);
and U1073 (N_1073,N_989,N_1035);
or U1074 (N_1074,N_1027,N_1019);
or U1075 (N_1075,N_994,N_1006);
or U1076 (N_1076,N_1043,N_1015);
or U1077 (N_1077,N_1037,N_1020);
or U1078 (N_1078,N_993,N_1016);
or U1079 (N_1079,N_1022,N_1032);
and U1080 (N_1080,N_977,N_999);
or U1081 (N_1081,N_1003,N_1034);
and U1082 (N_1082,N_1012,N_1005);
nand U1083 (N_1083,N_1048,N_1011);
and U1084 (N_1084,N_978,N_1049);
nand U1085 (N_1085,N_991,N_979);
and U1086 (N_1086,N_984,N_997);
or U1087 (N_1087,N_987,N_1014);
xnor U1088 (N_1088,N_1003,N_994);
and U1089 (N_1089,N_1039,N_1024);
nand U1090 (N_1090,N_1033,N_988);
and U1091 (N_1091,N_994,N_1019);
or U1092 (N_1092,N_990,N_979);
or U1093 (N_1093,N_1011,N_987);
and U1094 (N_1094,N_1000,N_1002);
nand U1095 (N_1095,N_987,N_1049);
nand U1096 (N_1096,N_1028,N_1023);
and U1097 (N_1097,N_1016,N_1033);
nand U1098 (N_1098,N_985,N_1004);
or U1099 (N_1099,N_1039,N_1011);
nand U1100 (N_1100,N_1034,N_1032);
or U1101 (N_1101,N_1016,N_1006);
or U1102 (N_1102,N_979,N_1009);
nor U1103 (N_1103,N_1023,N_983);
nor U1104 (N_1104,N_1013,N_1044);
or U1105 (N_1105,N_1027,N_1047);
nor U1106 (N_1106,N_1017,N_1048);
or U1107 (N_1107,N_980,N_987);
nor U1108 (N_1108,N_982,N_994);
nor U1109 (N_1109,N_1015,N_999);
nor U1110 (N_1110,N_1023,N_1005);
nor U1111 (N_1111,N_983,N_1002);
and U1112 (N_1112,N_997,N_980);
and U1113 (N_1113,N_1012,N_1029);
and U1114 (N_1114,N_1029,N_996);
nor U1115 (N_1115,N_1032,N_985);
nand U1116 (N_1116,N_983,N_1015);
nor U1117 (N_1117,N_991,N_982);
nand U1118 (N_1118,N_1024,N_991);
nor U1119 (N_1119,N_1025,N_998);
and U1120 (N_1120,N_985,N_997);
or U1121 (N_1121,N_1005,N_1025);
nand U1122 (N_1122,N_1022,N_987);
nand U1123 (N_1123,N_1030,N_1020);
nand U1124 (N_1124,N_1032,N_1007);
or U1125 (N_1125,N_1112,N_1077);
nor U1126 (N_1126,N_1097,N_1064);
nand U1127 (N_1127,N_1072,N_1076);
or U1128 (N_1128,N_1115,N_1096);
or U1129 (N_1129,N_1056,N_1114);
nand U1130 (N_1130,N_1071,N_1050);
nand U1131 (N_1131,N_1082,N_1120);
nor U1132 (N_1132,N_1055,N_1058);
or U1133 (N_1133,N_1123,N_1078);
or U1134 (N_1134,N_1104,N_1070);
nand U1135 (N_1135,N_1074,N_1113);
nor U1136 (N_1136,N_1110,N_1060);
and U1137 (N_1137,N_1105,N_1117);
nand U1138 (N_1138,N_1116,N_1106);
nor U1139 (N_1139,N_1054,N_1081);
nor U1140 (N_1140,N_1088,N_1108);
xor U1141 (N_1141,N_1069,N_1092);
nand U1142 (N_1142,N_1086,N_1073);
nor U1143 (N_1143,N_1059,N_1068);
nor U1144 (N_1144,N_1063,N_1102);
nand U1145 (N_1145,N_1065,N_1099);
nand U1146 (N_1146,N_1122,N_1101);
nand U1147 (N_1147,N_1109,N_1118);
nand U1148 (N_1148,N_1080,N_1079);
nand U1149 (N_1149,N_1103,N_1094);
and U1150 (N_1150,N_1107,N_1090);
or U1151 (N_1151,N_1124,N_1053);
and U1152 (N_1152,N_1057,N_1066);
or U1153 (N_1153,N_1084,N_1075);
nor U1154 (N_1154,N_1083,N_1087);
or U1155 (N_1155,N_1121,N_1067);
and U1156 (N_1156,N_1085,N_1098);
nand U1157 (N_1157,N_1093,N_1052);
and U1158 (N_1158,N_1100,N_1051);
and U1159 (N_1159,N_1091,N_1062);
nand U1160 (N_1160,N_1061,N_1095);
and U1161 (N_1161,N_1119,N_1089);
nor U1162 (N_1162,N_1111,N_1056);
and U1163 (N_1163,N_1091,N_1089);
nand U1164 (N_1164,N_1060,N_1101);
nand U1165 (N_1165,N_1121,N_1112);
nor U1166 (N_1166,N_1114,N_1110);
nor U1167 (N_1167,N_1117,N_1118);
nor U1168 (N_1168,N_1084,N_1052);
nand U1169 (N_1169,N_1122,N_1068);
and U1170 (N_1170,N_1087,N_1061);
or U1171 (N_1171,N_1100,N_1109);
nor U1172 (N_1172,N_1106,N_1066);
and U1173 (N_1173,N_1060,N_1116);
xnor U1174 (N_1174,N_1079,N_1061);
and U1175 (N_1175,N_1093,N_1098);
nor U1176 (N_1176,N_1106,N_1067);
nand U1177 (N_1177,N_1068,N_1078);
nand U1178 (N_1178,N_1050,N_1073);
nor U1179 (N_1179,N_1058,N_1084);
nand U1180 (N_1180,N_1080,N_1087);
nor U1181 (N_1181,N_1089,N_1108);
nor U1182 (N_1182,N_1124,N_1085);
and U1183 (N_1183,N_1064,N_1102);
nand U1184 (N_1184,N_1054,N_1053);
or U1185 (N_1185,N_1065,N_1075);
nand U1186 (N_1186,N_1051,N_1086);
xnor U1187 (N_1187,N_1051,N_1117);
and U1188 (N_1188,N_1069,N_1083);
nand U1189 (N_1189,N_1080,N_1051);
and U1190 (N_1190,N_1122,N_1075);
and U1191 (N_1191,N_1082,N_1094);
xnor U1192 (N_1192,N_1078,N_1100);
and U1193 (N_1193,N_1058,N_1113);
or U1194 (N_1194,N_1050,N_1103);
nor U1195 (N_1195,N_1093,N_1067);
nand U1196 (N_1196,N_1068,N_1067);
and U1197 (N_1197,N_1117,N_1052);
xor U1198 (N_1198,N_1055,N_1051);
and U1199 (N_1199,N_1124,N_1057);
nor U1200 (N_1200,N_1143,N_1146);
and U1201 (N_1201,N_1159,N_1154);
nand U1202 (N_1202,N_1166,N_1178);
and U1203 (N_1203,N_1139,N_1187);
and U1204 (N_1204,N_1184,N_1163);
nand U1205 (N_1205,N_1130,N_1155);
nor U1206 (N_1206,N_1129,N_1175);
nand U1207 (N_1207,N_1198,N_1160);
or U1208 (N_1208,N_1161,N_1162);
nor U1209 (N_1209,N_1179,N_1181);
and U1210 (N_1210,N_1194,N_1172);
nand U1211 (N_1211,N_1134,N_1168);
and U1212 (N_1212,N_1137,N_1193);
and U1213 (N_1213,N_1141,N_1151);
nand U1214 (N_1214,N_1138,N_1167);
and U1215 (N_1215,N_1133,N_1192);
and U1216 (N_1216,N_1140,N_1136);
or U1217 (N_1217,N_1195,N_1183);
or U1218 (N_1218,N_1126,N_1132);
nand U1219 (N_1219,N_1156,N_1147);
nand U1220 (N_1220,N_1145,N_1171);
or U1221 (N_1221,N_1197,N_1169);
and U1222 (N_1222,N_1180,N_1191);
nor U1223 (N_1223,N_1164,N_1158);
nand U1224 (N_1224,N_1165,N_1131);
and U1225 (N_1225,N_1125,N_1152);
nand U1226 (N_1226,N_1142,N_1186);
nor U1227 (N_1227,N_1153,N_1190);
nand U1228 (N_1228,N_1173,N_1149);
nor U1229 (N_1229,N_1185,N_1157);
nand U1230 (N_1230,N_1199,N_1176);
or U1231 (N_1231,N_1177,N_1188);
and U1232 (N_1232,N_1170,N_1189);
nand U1233 (N_1233,N_1127,N_1174);
and U1234 (N_1234,N_1135,N_1148);
nand U1235 (N_1235,N_1182,N_1196);
nand U1236 (N_1236,N_1150,N_1128);
and U1237 (N_1237,N_1144,N_1178);
and U1238 (N_1238,N_1165,N_1148);
xor U1239 (N_1239,N_1176,N_1129);
and U1240 (N_1240,N_1138,N_1147);
nand U1241 (N_1241,N_1171,N_1134);
or U1242 (N_1242,N_1177,N_1162);
nand U1243 (N_1243,N_1151,N_1133);
nand U1244 (N_1244,N_1146,N_1188);
and U1245 (N_1245,N_1171,N_1135);
nand U1246 (N_1246,N_1128,N_1147);
nand U1247 (N_1247,N_1145,N_1195);
xor U1248 (N_1248,N_1166,N_1156);
nand U1249 (N_1249,N_1152,N_1179);
xor U1250 (N_1250,N_1194,N_1183);
nor U1251 (N_1251,N_1160,N_1177);
and U1252 (N_1252,N_1143,N_1132);
nand U1253 (N_1253,N_1173,N_1151);
nor U1254 (N_1254,N_1176,N_1169);
or U1255 (N_1255,N_1151,N_1139);
or U1256 (N_1256,N_1183,N_1145);
nor U1257 (N_1257,N_1130,N_1129);
nor U1258 (N_1258,N_1131,N_1127);
nand U1259 (N_1259,N_1179,N_1132);
and U1260 (N_1260,N_1183,N_1188);
or U1261 (N_1261,N_1192,N_1144);
nor U1262 (N_1262,N_1127,N_1126);
nand U1263 (N_1263,N_1197,N_1190);
or U1264 (N_1264,N_1139,N_1172);
nand U1265 (N_1265,N_1127,N_1187);
nand U1266 (N_1266,N_1187,N_1165);
and U1267 (N_1267,N_1128,N_1158);
and U1268 (N_1268,N_1192,N_1137);
or U1269 (N_1269,N_1173,N_1139);
nor U1270 (N_1270,N_1162,N_1135);
xor U1271 (N_1271,N_1199,N_1127);
and U1272 (N_1272,N_1168,N_1140);
nand U1273 (N_1273,N_1183,N_1138);
nor U1274 (N_1274,N_1192,N_1129);
nor U1275 (N_1275,N_1266,N_1226);
nor U1276 (N_1276,N_1208,N_1243);
nand U1277 (N_1277,N_1268,N_1230);
nand U1278 (N_1278,N_1245,N_1213);
and U1279 (N_1279,N_1250,N_1224);
and U1280 (N_1280,N_1248,N_1220);
nand U1281 (N_1281,N_1225,N_1204);
nor U1282 (N_1282,N_1252,N_1214);
or U1283 (N_1283,N_1264,N_1201);
nand U1284 (N_1284,N_1256,N_1265);
and U1285 (N_1285,N_1203,N_1257);
nand U1286 (N_1286,N_1255,N_1270);
nand U1287 (N_1287,N_1253,N_1216);
and U1288 (N_1288,N_1240,N_1227);
nor U1289 (N_1289,N_1211,N_1237);
or U1290 (N_1290,N_1260,N_1274);
nand U1291 (N_1291,N_1200,N_1206);
and U1292 (N_1292,N_1205,N_1261);
nor U1293 (N_1293,N_1222,N_1221);
nand U1294 (N_1294,N_1241,N_1263);
and U1295 (N_1295,N_1249,N_1269);
nand U1296 (N_1296,N_1219,N_1262);
nor U1297 (N_1297,N_1233,N_1272);
nand U1298 (N_1298,N_1239,N_1217);
nand U1299 (N_1299,N_1258,N_1209);
nand U1300 (N_1300,N_1271,N_1254);
or U1301 (N_1301,N_1238,N_1212);
nand U1302 (N_1302,N_1207,N_1223);
or U1303 (N_1303,N_1259,N_1236);
and U1304 (N_1304,N_1273,N_1231);
nor U1305 (N_1305,N_1246,N_1210);
or U1306 (N_1306,N_1218,N_1215);
nand U1307 (N_1307,N_1247,N_1228);
nor U1308 (N_1308,N_1242,N_1235);
or U1309 (N_1309,N_1202,N_1229);
and U1310 (N_1310,N_1234,N_1232);
nand U1311 (N_1311,N_1267,N_1251);
and U1312 (N_1312,N_1244,N_1203);
nand U1313 (N_1313,N_1226,N_1257);
nor U1314 (N_1314,N_1274,N_1246);
nand U1315 (N_1315,N_1241,N_1200);
and U1316 (N_1316,N_1227,N_1247);
and U1317 (N_1317,N_1236,N_1235);
nand U1318 (N_1318,N_1229,N_1243);
or U1319 (N_1319,N_1266,N_1241);
nor U1320 (N_1320,N_1273,N_1226);
or U1321 (N_1321,N_1245,N_1242);
and U1322 (N_1322,N_1231,N_1247);
and U1323 (N_1323,N_1212,N_1220);
and U1324 (N_1324,N_1267,N_1225);
nor U1325 (N_1325,N_1252,N_1250);
or U1326 (N_1326,N_1274,N_1253);
and U1327 (N_1327,N_1205,N_1264);
or U1328 (N_1328,N_1237,N_1236);
nand U1329 (N_1329,N_1246,N_1242);
nand U1330 (N_1330,N_1209,N_1238);
nor U1331 (N_1331,N_1221,N_1250);
and U1332 (N_1332,N_1272,N_1237);
nand U1333 (N_1333,N_1236,N_1242);
and U1334 (N_1334,N_1264,N_1229);
and U1335 (N_1335,N_1263,N_1273);
nor U1336 (N_1336,N_1233,N_1268);
or U1337 (N_1337,N_1274,N_1204);
and U1338 (N_1338,N_1246,N_1212);
and U1339 (N_1339,N_1219,N_1267);
or U1340 (N_1340,N_1204,N_1206);
nor U1341 (N_1341,N_1203,N_1245);
and U1342 (N_1342,N_1259,N_1213);
or U1343 (N_1343,N_1203,N_1248);
nand U1344 (N_1344,N_1252,N_1269);
and U1345 (N_1345,N_1208,N_1226);
and U1346 (N_1346,N_1265,N_1260);
nand U1347 (N_1347,N_1229,N_1242);
or U1348 (N_1348,N_1202,N_1230);
nor U1349 (N_1349,N_1264,N_1252);
or U1350 (N_1350,N_1348,N_1317);
and U1351 (N_1351,N_1312,N_1297);
or U1352 (N_1352,N_1333,N_1278);
and U1353 (N_1353,N_1329,N_1302);
nand U1354 (N_1354,N_1316,N_1275);
nand U1355 (N_1355,N_1346,N_1347);
and U1356 (N_1356,N_1307,N_1337);
nand U1357 (N_1357,N_1292,N_1305);
and U1358 (N_1358,N_1282,N_1344);
and U1359 (N_1359,N_1325,N_1334);
or U1360 (N_1360,N_1308,N_1281);
nor U1361 (N_1361,N_1306,N_1338);
and U1362 (N_1362,N_1330,N_1341);
nand U1363 (N_1363,N_1318,N_1310);
nand U1364 (N_1364,N_1286,N_1299);
and U1365 (N_1365,N_1342,N_1322);
nand U1366 (N_1366,N_1343,N_1340);
and U1367 (N_1367,N_1314,N_1320);
nor U1368 (N_1368,N_1313,N_1323);
nand U1369 (N_1369,N_1283,N_1335);
or U1370 (N_1370,N_1315,N_1332);
nor U1371 (N_1371,N_1296,N_1345);
nor U1372 (N_1372,N_1309,N_1303);
nor U1373 (N_1373,N_1295,N_1276);
nor U1374 (N_1374,N_1298,N_1326);
or U1375 (N_1375,N_1280,N_1304);
and U1376 (N_1376,N_1284,N_1301);
nor U1377 (N_1377,N_1327,N_1311);
nor U1378 (N_1378,N_1290,N_1287);
and U1379 (N_1379,N_1300,N_1339);
nand U1380 (N_1380,N_1321,N_1291);
nor U1381 (N_1381,N_1277,N_1279);
and U1382 (N_1382,N_1349,N_1293);
or U1383 (N_1383,N_1288,N_1328);
and U1384 (N_1384,N_1294,N_1336);
or U1385 (N_1385,N_1331,N_1319);
nor U1386 (N_1386,N_1285,N_1324);
nor U1387 (N_1387,N_1289,N_1275);
nand U1388 (N_1388,N_1324,N_1340);
and U1389 (N_1389,N_1288,N_1276);
and U1390 (N_1390,N_1286,N_1343);
or U1391 (N_1391,N_1312,N_1332);
or U1392 (N_1392,N_1290,N_1306);
nand U1393 (N_1393,N_1334,N_1285);
nand U1394 (N_1394,N_1346,N_1333);
or U1395 (N_1395,N_1289,N_1345);
xnor U1396 (N_1396,N_1319,N_1295);
nand U1397 (N_1397,N_1330,N_1327);
or U1398 (N_1398,N_1320,N_1298);
xor U1399 (N_1399,N_1291,N_1315);
nand U1400 (N_1400,N_1349,N_1341);
and U1401 (N_1401,N_1295,N_1300);
and U1402 (N_1402,N_1294,N_1306);
and U1403 (N_1403,N_1298,N_1331);
nand U1404 (N_1404,N_1277,N_1275);
and U1405 (N_1405,N_1303,N_1310);
nor U1406 (N_1406,N_1337,N_1289);
nand U1407 (N_1407,N_1341,N_1297);
and U1408 (N_1408,N_1332,N_1330);
xor U1409 (N_1409,N_1327,N_1284);
nand U1410 (N_1410,N_1323,N_1286);
nor U1411 (N_1411,N_1324,N_1320);
xor U1412 (N_1412,N_1285,N_1313);
nor U1413 (N_1413,N_1289,N_1305);
nand U1414 (N_1414,N_1279,N_1349);
or U1415 (N_1415,N_1306,N_1309);
nand U1416 (N_1416,N_1308,N_1339);
xor U1417 (N_1417,N_1311,N_1318);
or U1418 (N_1418,N_1299,N_1349);
and U1419 (N_1419,N_1323,N_1302);
and U1420 (N_1420,N_1348,N_1349);
and U1421 (N_1421,N_1315,N_1290);
and U1422 (N_1422,N_1334,N_1345);
and U1423 (N_1423,N_1335,N_1282);
nor U1424 (N_1424,N_1313,N_1322);
or U1425 (N_1425,N_1412,N_1385);
nor U1426 (N_1426,N_1413,N_1364);
and U1427 (N_1427,N_1417,N_1384);
and U1428 (N_1428,N_1418,N_1397);
and U1429 (N_1429,N_1419,N_1372);
and U1430 (N_1430,N_1362,N_1369);
nand U1431 (N_1431,N_1377,N_1354);
nand U1432 (N_1432,N_1368,N_1394);
or U1433 (N_1433,N_1366,N_1395);
nor U1434 (N_1434,N_1422,N_1406);
nor U1435 (N_1435,N_1371,N_1400);
or U1436 (N_1436,N_1410,N_1367);
or U1437 (N_1437,N_1389,N_1365);
nand U1438 (N_1438,N_1363,N_1396);
nor U1439 (N_1439,N_1420,N_1393);
or U1440 (N_1440,N_1390,N_1379);
or U1441 (N_1441,N_1381,N_1415);
nand U1442 (N_1442,N_1352,N_1388);
or U1443 (N_1443,N_1401,N_1399);
nor U1444 (N_1444,N_1414,N_1375);
nor U1445 (N_1445,N_1353,N_1361);
nand U1446 (N_1446,N_1392,N_1376);
nor U1447 (N_1447,N_1391,N_1402);
or U1448 (N_1448,N_1398,N_1416);
nand U1449 (N_1449,N_1421,N_1380);
nor U1450 (N_1450,N_1373,N_1382);
and U1451 (N_1451,N_1407,N_1387);
nor U1452 (N_1452,N_1351,N_1403);
and U1453 (N_1453,N_1408,N_1357);
nor U1454 (N_1454,N_1409,N_1404);
and U1455 (N_1455,N_1358,N_1370);
or U1456 (N_1456,N_1405,N_1359);
or U1457 (N_1457,N_1424,N_1386);
and U1458 (N_1458,N_1355,N_1378);
xnor U1459 (N_1459,N_1374,N_1423);
or U1460 (N_1460,N_1350,N_1356);
or U1461 (N_1461,N_1411,N_1360);
nor U1462 (N_1462,N_1383,N_1411);
or U1463 (N_1463,N_1386,N_1400);
nor U1464 (N_1464,N_1375,N_1374);
and U1465 (N_1465,N_1379,N_1360);
xor U1466 (N_1466,N_1398,N_1369);
nand U1467 (N_1467,N_1376,N_1410);
or U1468 (N_1468,N_1391,N_1371);
nor U1469 (N_1469,N_1395,N_1414);
or U1470 (N_1470,N_1364,N_1353);
nand U1471 (N_1471,N_1364,N_1363);
nor U1472 (N_1472,N_1395,N_1408);
and U1473 (N_1473,N_1369,N_1410);
or U1474 (N_1474,N_1377,N_1356);
or U1475 (N_1475,N_1391,N_1363);
nand U1476 (N_1476,N_1424,N_1412);
xnor U1477 (N_1477,N_1397,N_1412);
and U1478 (N_1478,N_1416,N_1410);
nand U1479 (N_1479,N_1404,N_1400);
nor U1480 (N_1480,N_1424,N_1392);
and U1481 (N_1481,N_1399,N_1418);
nand U1482 (N_1482,N_1406,N_1351);
nor U1483 (N_1483,N_1407,N_1384);
or U1484 (N_1484,N_1350,N_1406);
nor U1485 (N_1485,N_1393,N_1389);
or U1486 (N_1486,N_1383,N_1375);
and U1487 (N_1487,N_1386,N_1382);
or U1488 (N_1488,N_1415,N_1351);
nand U1489 (N_1489,N_1394,N_1372);
or U1490 (N_1490,N_1370,N_1381);
xnor U1491 (N_1491,N_1374,N_1418);
or U1492 (N_1492,N_1393,N_1396);
or U1493 (N_1493,N_1394,N_1379);
xor U1494 (N_1494,N_1395,N_1351);
nor U1495 (N_1495,N_1394,N_1403);
or U1496 (N_1496,N_1415,N_1393);
and U1497 (N_1497,N_1387,N_1372);
or U1498 (N_1498,N_1409,N_1359);
nor U1499 (N_1499,N_1376,N_1363);
nor U1500 (N_1500,N_1470,N_1446);
nand U1501 (N_1501,N_1496,N_1491);
or U1502 (N_1502,N_1467,N_1479);
nor U1503 (N_1503,N_1474,N_1444);
and U1504 (N_1504,N_1445,N_1462);
nand U1505 (N_1505,N_1468,N_1458);
nand U1506 (N_1506,N_1494,N_1429);
nand U1507 (N_1507,N_1435,N_1490);
nand U1508 (N_1508,N_1492,N_1485);
and U1509 (N_1509,N_1466,N_1436);
nor U1510 (N_1510,N_1495,N_1487);
xor U1511 (N_1511,N_1498,N_1438);
nor U1512 (N_1512,N_1427,N_1450);
nand U1513 (N_1513,N_1447,N_1426);
nand U1514 (N_1514,N_1463,N_1449);
and U1515 (N_1515,N_1433,N_1453);
xnor U1516 (N_1516,N_1471,N_1431);
nand U1517 (N_1517,N_1434,N_1493);
nor U1518 (N_1518,N_1483,N_1477);
or U1519 (N_1519,N_1489,N_1499);
or U1520 (N_1520,N_1497,N_1480);
nand U1521 (N_1521,N_1482,N_1473);
and U1522 (N_1522,N_1442,N_1451);
or U1523 (N_1523,N_1461,N_1465);
and U1524 (N_1524,N_1432,N_1437);
and U1525 (N_1525,N_1475,N_1425);
nand U1526 (N_1526,N_1440,N_1457);
and U1527 (N_1527,N_1452,N_1443);
nor U1528 (N_1528,N_1441,N_1464);
and U1529 (N_1529,N_1454,N_1428);
xnor U1530 (N_1530,N_1486,N_1439);
nand U1531 (N_1531,N_1448,N_1460);
nor U1532 (N_1532,N_1430,N_1456);
and U1533 (N_1533,N_1455,N_1472);
nor U1534 (N_1534,N_1476,N_1469);
or U1535 (N_1535,N_1488,N_1484);
and U1536 (N_1536,N_1459,N_1481);
xnor U1537 (N_1537,N_1478,N_1490);
or U1538 (N_1538,N_1498,N_1474);
and U1539 (N_1539,N_1468,N_1497);
and U1540 (N_1540,N_1458,N_1432);
or U1541 (N_1541,N_1494,N_1475);
nand U1542 (N_1542,N_1493,N_1425);
nor U1543 (N_1543,N_1434,N_1471);
nand U1544 (N_1544,N_1496,N_1435);
or U1545 (N_1545,N_1462,N_1432);
nand U1546 (N_1546,N_1487,N_1477);
or U1547 (N_1547,N_1465,N_1475);
nand U1548 (N_1548,N_1462,N_1468);
and U1549 (N_1549,N_1426,N_1480);
and U1550 (N_1550,N_1462,N_1450);
or U1551 (N_1551,N_1446,N_1451);
nor U1552 (N_1552,N_1451,N_1427);
xnor U1553 (N_1553,N_1496,N_1446);
nand U1554 (N_1554,N_1498,N_1433);
and U1555 (N_1555,N_1487,N_1437);
nor U1556 (N_1556,N_1429,N_1489);
or U1557 (N_1557,N_1455,N_1444);
and U1558 (N_1558,N_1481,N_1471);
or U1559 (N_1559,N_1478,N_1477);
and U1560 (N_1560,N_1460,N_1489);
or U1561 (N_1561,N_1429,N_1488);
nand U1562 (N_1562,N_1498,N_1477);
or U1563 (N_1563,N_1463,N_1489);
and U1564 (N_1564,N_1461,N_1457);
nor U1565 (N_1565,N_1460,N_1478);
nor U1566 (N_1566,N_1441,N_1490);
or U1567 (N_1567,N_1439,N_1458);
nand U1568 (N_1568,N_1427,N_1494);
nand U1569 (N_1569,N_1453,N_1470);
nand U1570 (N_1570,N_1436,N_1491);
or U1571 (N_1571,N_1429,N_1456);
and U1572 (N_1572,N_1431,N_1469);
nand U1573 (N_1573,N_1430,N_1432);
and U1574 (N_1574,N_1498,N_1470);
and U1575 (N_1575,N_1530,N_1522);
and U1576 (N_1576,N_1536,N_1568);
and U1577 (N_1577,N_1535,N_1505);
and U1578 (N_1578,N_1541,N_1549);
xor U1579 (N_1579,N_1540,N_1544);
and U1580 (N_1580,N_1550,N_1552);
nand U1581 (N_1581,N_1546,N_1560);
and U1582 (N_1582,N_1501,N_1565);
or U1583 (N_1583,N_1545,N_1500);
or U1584 (N_1584,N_1524,N_1521);
nor U1585 (N_1585,N_1564,N_1555);
nand U1586 (N_1586,N_1561,N_1515);
and U1587 (N_1587,N_1573,N_1502);
nor U1588 (N_1588,N_1572,N_1523);
xor U1589 (N_1589,N_1562,N_1542);
or U1590 (N_1590,N_1504,N_1569);
nor U1591 (N_1591,N_1506,N_1517);
nor U1592 (N_1592,N_1529,N_1528);
and U1593 (N_1593,N_1557,N_1559);
nor U1594 (N_1594,N_1512,N_1526);
nor U1595 (N_1595,N_1543,N_1539);
nor U1596 (N_1596,N_1507,N_1556);
and U1597 (N_1597,N_1566,N_1547);
and U1598 (N_1598,N_1567,N_1534);
nand U1599 (N_1599,N_1532,N_1520);
and U1600 (N_1600,N_1518,N_1551);
and U1601 (N_1601,N_1511,N_1571);
nand U1602 (N_1602,N_1553,N_1516);
nor U1603 (N_1603,N_1533,N_1554);
nor U1604 (N_1604,N_1570,N_1510);
nand U1605 (N_1605,N_1525,N_1531);
or U1606 (N_1606,N_1548,N_1503);
or U1607 (N_1607,N_1558,N_1563);
xor U1608 (N_1608,N_1527,N_1514);
nand U1609 (N_1609,N_1509,N_1537);
or U1610 (N_1610,N_1519,N_1574);
or U1611 (N_1611,N_1508,N_1513);
nand U1612 (N_1612,N_1538,N_1564);
nor U1613 (N_1613,N_1547,N_1543);
nand U1614 (N_1614,N_1568,N_1550);
and U1615 (N_1615,N_1546,N_1543);
or U1616 (N_1616,N_1564,N_1537);
or U1617 (N_1617,N_1507,N_1515);
nor U1618 (N_1618,N_1569,N_1531);
or U1619 (N_1619,N_1528,N_1541);
and U1620 (N_1620,N_1541,N_1564);
and U1621 (N_1621,N_1540,N_1519);
nor U1622 (N_1622,N_1502,N_1574);
xor U1623 (N_1623,N_1527,N_1557);
nand U1624 (N_1624,N_1566,N_1543);
nor U1625 (N_1625,N_1523,N_1503);
and U1626 (N_1626,N_1571,N_1548);
or U1627 (N_1627,N_1528,N_1501);
or U1628 (N_1628,N_1550,N_1500);
or U1629 (N_1629,N_1560,N_1533);
and U1630 (N_1630,N_1501,N_1514);
or U1631 (N_1631,N_1529,N_1563);
and U1632 (N_1632,N_1555,N_1520);
nand U1633 (N_1633,N_1536,N_1534);
and U1634 (N_1634,N_1518,N_1570);
nor U1635 (N_1635,N_1502,N_1523);
and U1636 (N_1636,N_1507,N_1561);
nor U1637 (N_1637,N_1537,N_1526);
or U1638 (N_1638,N_1544,N_1501);
nand U1639 (N_1639,N_1563,N_1546);
nand U1640 (N_1640,N_1538,N_1534);
nor U1641 (N_1641,N_1513,N_1504);
and U1642 (N_1642,N_1548,N_1547);
nand U1643 (N_1643,N_1560,N_1509);
and U1644 (N_1644,N_1545,N_1567);
nor U1645 (N_1645,N_1541,N_1544);
or U1646 (N_1646,N_1516,N_1562);
and U1647 (N_1647,N_1521,N_1535);
or U1648 (N_1648,N_1565,N_1504);
or U1649 (N_1649,N_1570,N_1571);
nand U1650 (N_1650,N_1578,N_1606);
or U1651 (N_1651,N_1577,N_1640);
nand U1652 (N_1652,N_1641,N_1613);
nor U1653 (N_1653,N_1603,N_1637);
nor U1654 (N_1654,N_1610,N_1607);
nor U1655 (N_1655,N_1580,N_1630);
nand U1656 (N_1656,N_1625,N_1627);
and U1657 (N_1657,N_1621,N_1593);
xor U1658 (N_1658,N_1647,N_1584);
or U1659 (N_1659,N_1588,N_1599);
nand U1660 (N_1660,N_1623,N_1631);
or U1661 (N_1661,N_1632,N_1608);
nand U1662 (N_1662,N_1642,N_1635);
xnor U1663 (N_1663,N_1620,N_1628);
and U1664 (N_1664,N_1600,N_1585);
nand U1665 (N_1665,N_1586,N_1649);
or U1666 (N_1666,N_1597,N_1643);
and U1667 (N_1667,N_1622,N_1594);
xnor U1668 (N_1668,N_1591,N_1582);
or U1669 (N_1669,N_1614,N_1583);
nand U1670 (N_1670,N_1575,N_1618);
nand U1671 (N_1671,N_1612,N_1601);
or U1672 (N_1672,N_1636,N_1589);
nor U1673 (N_1673,N_1579,N_1633);
and U1674 (N_1674,N_1646,N_1605);
or U1675 (N_1675,N_1639,N_1587);
and U1676 (N_1676,N_1645,N_1648);
or U1677 (N_1677,N_1644,N_1604);
nand U1678 (N_1678,N_1596,N_1617);
nand U1679 (N_1679,N_1634,N_1595);
or U1680 (N_1680,N_1619,N_1590);
and U1681 (N_1681,N_1615,N_1611);
nor U1682 (N_1682,N_1581,N_1626);
and U1683 (N_1683,N_1602,N_1616);
or U1684 (N_1684,N_1629,N_1576);
nor U1685 (N_1685,N_1592,N_1609);
nand U1686 (N_1686,N_1638,N_1624);
nand U1687 (N_1687,N_1598,N_1596);
nand U1688 (N_1688,N_1616,N_1608);
and U1689 (N_1689,N_1614,N_1632);
and U1690 (N_1690,N_1628,N_1644);
or U1691 (N_1691,N_1647,N_1579);
nand U1692 (N_1692,N_1645,N_1596);
and U1693 (N_1693,N_1612,N_1595);
and U1694 (N_1694,N_1594,N_1608);
or U1695 (N_1695,N_1642,N_1631);
nand U1696 (N_1696,N_1623,N_1595);
and U1697 (N_1697,N_1580,N_1585);
nor U1698 (N_1698,N_1619,N_1585);
and U1699 (N_1699,N_1626,N_1596);
and U1700 (N_1700,N_1584,N_1630);
nand U1701 (N_1701,N_1647,N_1630);
nand U1702 (N_1702,N_1597,N_1642);
nand U1703 (N_1703,N_1639,N_1591);
nand U1704 (N_1704,N_1626,N_1625);
or U1705 (N_1705,N_1589,N_1587);
and U1706 (N_1706,N_1605,N_1609);
nor U1707 (N_1707,N_1591,N_1578);
or U1708 (N_1708,N_1615,N_1608);
and U1709 (N_1709,N_1609,N_1619);
nand U1710 (N_1710,N_1599,N_1643);
nor U1711 (N_1711,N_1624,N_1629);
nor U1712 (N_1712,N_1649,N_1626);
or U1713 (N_1713,N_1593,N_1639);
nand U1714 (N_1714,N_1590,N_1638);
nor U1715 (N_1715,N_1579,N_1589);
nor U1716 (N_1716,N_1606,N_1635);
and U1717 (N_1717,N_1644,N_1591);
or U1718 (N_1718,N_1614,N_1628);
nand U1719 (N_1719,N_1590,N_1603);
nand U1720 (N_1720,N_1587,N_1590);
nor U1721 (N_1721,N_1630,N_1610);
and U1722 (N_1722,N_1589,N_1607);
and U1723 (N_1723,N_1647,N_1576);
nor U1724 (N_1724,N_1638,N_1600);
nand U1725 (N_1725,N_1715,N_1671);
or U1726 (N_1726,N_1669,N_1720);
nor U1727 (N_1727,N_1677,N_1654);
or U1728 (N_1728,N_1716,N_1699);
and U1729 (N_1729,N_1659,N_1724);
or U1730 (N_1730,N_1667,N_1660);
nor U1731 (N_1731,N_1655,N_1678);
nand U1732 (N_1732,N_1687,N_1714);
xnor U1733 (N_1733,N_1657,N_1708);
or U1734 (N_1734,N_1718,N_1702);
nor U1735 (N_1735,N_1695,N_1682);
or U1736 (N_1736,N_1652,N_1665);
xnor U1737 (N_1737,N_1661,N_1653);
and U1738 (N_1738,N_1686,N_1656);
or U1739 (N_1739,N_1697,N_1675);
and U1740 (N_1740,N_1706,N_1670);
nor U1741 (N_1741,N_1722,N_1711);
and U1742 (N_1742,N_1723,N_1679);
nor U1743 (N_1743,N_1701,N_1666);
and U1744 (N_1744,N_1692,N_1710);
nand U1745 (N_1745,N_1681,N_1683);
and U1746 (N_1746,N_1673,N_1690);
xor U1747 (N_1747,N_1685,N_1703);
nand U1748 (N_1748,N_1698,N_1719);
nand U1749 (N_1749,N_1664,N_1650);
nor U1750 (N_1750,N_1668,N_1684);
xnor U1751 (N_1751,N_1662,N_1676);
and U1752 (N_1752,N_1700,N_1688);
or U1753 (N_1753,N_1696,N_1704);
nand U1754 (N_1754,N_1709,N_1680);
nor U1755 (N_1755,N_1663,N_1705);
and U1756 (N_1756,N_1717,N_1674);
nand U1757 (N_1757,N_1694,N_1672);
nand U1758 (N_1758,N_1658,N_1651);
nor U1759 (N_1759,N_1712,N_1713);
nor U1760 (N_1760,N_1707,N_1691);
or U1761 (N_1761,N_1693,N_1689);
nor U1762 (N_1762,N_1721,N_1665);
or U1763 (N_1763,N_1656,N_1675);
nor U1764 (N_1764,N_1664,N_1689);
nand U1765 (N_1765,N_1695,N_1668);
and U1766 (N_1766,N_1713,N_1707);
and U1767 (N_1767,N_1656,N_1650);
nand U1768 (N_1768,N_1696,N_1717);
nand U1769 (N_1769,N_1700,N_1691);
and U1770 (N_1770,N_1717,N_1660);
nor U1771 (N_1771,N_1717,N_1668);
and U1772 (N_1772,N_1710,N_1679);
nor U1773 (N_1773,N_1711,N_1656);
xor U1774 (N_1774,N_1718,N_1665);
or U1775 (N_1775,N_1701,N_1683);
and U1776 (N_1776,N_1678,N_1690);
nand U1777 (N_1777,N_1716,N_1721);
nand U1778 (N_1778,N_1655,N_1651);
nor U1779 (N_1779,N_1664,N_1678);
nand U1780 (N_1780,N_1720,N_1674);
nor U1781 (N_1781,N_1691,N_1682);
and U1782 (N_1782,N_1716,N_1687);
and U1783 (N_1783,N_1663,N_1664);
nor U1784 (N_1784,N_1661,N_1693);
nor U1785 (N_1785,N_1661,N_1662);
nor U1786 (N_1786,N_1720,N_1666);
and U1787 (N_1787,N_1712,N_1669);
and U1788 (N_1788,N_1720,N_1714);
and U1789 (N_1789,N_1693,N_1721);
nor U1790 (N_1790,N_1713,N_1701);
or U1791 (N_1791,N_1723,N_1714);
and U1792 (N_1792,N_1683,N_1654);
nand U1793 (N_1793,N_1706,N_1661);
and U1794 (N_1794,N_1679,N_1672);
or U1795 (N_1795,N_1656,N_1655);
or U1796 (N_1796,N_1678,N_1696);
and U1797 (N_1797,N_1673,N_1717);
and U1798 (N_1798,N_1662,N_1682);
and U1799 (N_1799,N_1662,N_1675);
nor U1800 (N_1800,N_1750,N_1790);
nor U1801 (N_1801,N_1782,N_1776);
or U1802 (N_1802,N_1771,N_1795);
and U1803 (N_1803,N_1738,N_1765);
nand U1804 (N_1804,N_1729,N_1777);
and U1805 (N_1805,N_1766,N_1780);
or U1806 (N_1806,N_1784,N_1751);
or U1807 (N_1807,N_1728,N_1792);
nor U1808 (N_1808,N_1791,N_1725);
xnor U1809 (N_1809,N_1785,N_1734);
nor U1810 (N_1810,N_1778,N_1786);
nand U1811 (N_1811,N_1769,N_1797);
nand U1812 (N_1812,N_1740,N_1753);
nor U1813 (N_1813,N_1748,N_1744);
nor U1814 (N_1814,N_1794,N_1745);
xnor U1815 (N_1815,N_1798,N_1739);
and U1816 (N_1816,N_1742,N_1767);
or U1817 (N_1817,N_1736,N_1787);
and U1818 (N_1818,N_1779,N_1773);
nor U1819 (N_1819,N_1741,N_1783);
nand U1820 (N_1820,N_1747,N_1756);
nand U1821 (N_1821,N_1761,N_1746);
or U1822 (N_1822,N_1757,N_1732);
xnor U1823 (N_1823,N_1759,N_1762);
nand U1824 (N_1824,N_1793,N_1730);
nor U1825 (N_1825,N_1781,N_1799);
or U1826 (N_1826,N_1796,N_1755);
nand U1827 (N_1827,N_1763,N_1735);
nor U1828 (N_1828,N_1731,N_1752);
nand U1829 (N_1829,N_1789,N_1726);
and U1830 (N_1830,N_1768,N_1760);
or U1831 (N_1831,N_1758,N_1764);
or U1832 (N_1832,N_1749,N_1754);
and U1833 (N_1833,N_1737,N_1772);
nor U1834 (N_1834,N_1770,N_1727);
nor U1835 (N_1835,N_1743,N_1775);
nor U1836 (N_1836,N_1788,N_1774);
or U1837 (N_1837,N_1733,N_1734);
nand U1838 (N_1838,N_1775,N_1752);
and U1839 (N_1839,N_1751,N_1769);
and U1840 (N_1840,N_1781,N_1748);
nand U1841 (N_1841,N_1734,N_1726);
or U1842 (N_1842,N_1795,N_1792);
or U1843 (N_1843,N_1725,N_1775);
and U1844 (N_1844,N_1787,N_1774);
nor U1845 (N_1845,N_1779,N_1742);
or U1846 (N_1846,N_1761,N_1745);
nor U1847 (N_1847,N_1731,N_1767);
or U1848 (N_1848,N_1757,N_1746);
nand U1849 (N_1849,N_1769,N_1749);
and U1850 (N_1850,N_1785,N_1758);
nor U1851 (N_1851,N_1736,N_1727);
and U1852 (N_1852,N_1755,N_1788);
nand U1853 (N_1853,N_1739,N_1773);
nor U1854 (N_1854,N_1750,N_1746);
nor U1855 (N_1855,N_1796,N_1754);
nor U1856 (N_1856,N_1768,N_1782);
or U1857 (N_1857,N_1758,N_1727);
nand U1858 (N_1858,N_1726,N_1794);
nand U1859 (N_1859,N_1735,N_1784);
xnor U1860 (N_1860,N_1754,N_1791);
nand U1861 (N_1861,N_1766,N_1744);
nor U1862 (N_1862,N_1749,N_1789);
or U1863 (N_1863,N_1754,N_1767);
nor U1864 (N_1864,N_1795,N_1733);
and U1865 (N_1865,N_1791,N_1795);
nand U1866 (N_1866,N_1789,N_1750);
nand U1867 (N_1867,N_1784,N_1754);
nand U1868 (N_1868,N_1799,N_1796);
or U1869 (N_1869,N_1774,N_1744);
nand U1870 (N_1870,N_1741,N_1787);
nor U1871 (N_1871,N_1754,N_1774);
nand U1872 (N_1872,N_1763,N_1790);
or U1873 (N_1873,N_1792,N_1751);
and U1874 (N_1874,N_1785,N_1779);
and U1875 (N_1875,N_1802,N_1824);
or U1876 (N_1876,N_1846,N_1854);
nand U1877 (N_1877,N_1867,N_1829);
nand U1878 (N_1878,N_1869,N_1860);
and U1879 (N_1879,N_1864,N_1816);
and U1880 (N_1880,N_1808,N_1805);
xnor U1881 (N_1881,N_1803,N_1850);
or U1882 (N_1882,N_1843,N_1856);
nor U1883 (N_1883,N_1800,N_1818);
and U1884 (N_1884,N_1863,N_1872);
or U1885 (N_1885,N_1813,N_1840);
or U1886 (N_1886,N_1842,N_1873);
or U1887 (N_1887,N_1819,N_1801);
or U1888 (N_1888,N_1871,N_1835);
nor U1889 (N_1889,N_1821,N_1852);
and U1890 (N_1890,N_1834,N_1838);
xnor U1891 (N_1891,N_1809,N_1823);
nand U1892 (N_1892,N_1857,N_1844);
and U1893 (N_1893,N_1848,N_1851);
nor U1894 (N_1894,N_1849,N_1855);
xor U1895 (N_1895,N_1862,N_1866);
or U1896 (N_1896,N_1858,N_1837);
or U1897 (N_1897,N_1810,N_1868);
nand U1898 (N_1898,N_1836,N_1826);
or U1899 (N_1899,N_1827,N_1822);
and U1900 (N_1900,N_1833,N_1817);
nand U1901 (N_1901,N_1874,N_1839);
nand U1902 (N_1902,N_1830,N_1853);
or U1903 (N_1903,N_1811,N_1841);
nor U1904 (N_1904,N_1847,N_1820);
nand U1905 (N_1905,N_1828,N_1807);
nand U1906 (N_1906,N_1832,N_1814);
nor U1907 (N_1907,N_1815,N_1806);
nand U1908 (N_1908,N_1804,N_1825);
or U1909 (N_1909,N_1845,N_1859);
nor U1910 (N_1910,N_1870,N_1861);
nand U1911 (N_1911,N_1831,N_1865);
nand U1912 (N_1912,N_1812,N_1821);
or U1913 (N_1913,N_1833,N_1866);
or U1914 (N_1914,N_1816,N_1857);
nand U1915 (N_1915,N_1865,N_1825);
nand U1916 (N_1916,N_1845,N_1807);
and U1917 (N_1917,N_1830,N_1812);
or U1918 (N_1918,N_1817,N_1821);
or U1919 (N_1919,N_1814,N_1808);
xor U1920 (N_1920,N_1811,N_1872);
or U1921 (N_1921,N_1861,N_1856);
nor U1922 (N_1922,N_1852,N_1862);
nor U1923 (N_1923,N_1820,N_1848);
nor U1924 (N_1924,N_1814,N_1839);
and U1925 (N_1925,N_1862,N_1851);
nor U1926 (N_1926,N_1864,N_1840);
nor U1927 (N_1927,N_1825,N_1859);
nor U1928 (N_1928,N_1809,N_1848);
nand U1929 (N_1929,N_1806,N_1818);
or U1930 (N_1930,N_1870,N_1845);
nand U1931 (N_1931,N_1867,N_1827);
or U1932 (N_1932,N_1873,N_1840);
nor U1933 (N_1933,N_1847,N_1815);
nand U1934 (N_1934,N_1831,N_1803);
nand U1935 (N_1935,N_1862,N_1820);
nand U1936 (N_1936,N_1872,N_1873);
nor U1937 (N_1937,N_1821,N_1834);
nor U1938 (N_1938,N_1829,N_1826);
nand U1939 (N_1939,N_1827,N_1818);
nor U1940 (N_1940,N_1841,N_1852);
nor U1941 (N_1941,N_1804,N_1869);
nor U1942 (N_1942,N_1835,N_1858);
nor U1943 (N_1943,N_1826,N_1821);
and U1944 (N_1944,N_1830,N_1823);
nand U1945 (N_1945,N_1811,N_1856);
and U1946 (N_1946,N_1809,N_1859);
and U1947 (N_1947,N_1873,N_1816);
or U1948 (N_1948,N_1849,N_1862);
or U1949 (N_1949,N_1842,N_1864);
or U1950 (N_1950,N_1919,N_1923);
nand U1951 (N_1951,N_1877,N_1927);
and U1952 (N_1952,N_1914,N_1916);
nand U1953 (N_1953,N_1886,N_1915);
nand U1954 (N_1954,N_1924,N_1887);
nand U1955 (N_1955,N_1875,N_1880);
and U1956 (N_1956,N_1932,N_1900);
nor U1957 (N_1957,N_1878,N_1894);
nor U1958 (N_1958,N_1940,N_1903);
xnor U1959 (N_1959,N_1926,N_1884);
nor U1960 (N_1960,N_1892,N_1902);
and U1961 (N_1961,N_1943,N_1942);
or U1962 (N_1962,N_1947,N_1938);
and U1963 (N_1963,N_1920,N_1945);
nor U1964 (N_1964,N_1883,N_1917);
nand U1965 (N_1965,N_1904,N_1948);
nor U1966 (N_1966,N_1934,N_1899);
nor U1967 (N_1967,N_1937,N_1944);
or U1968 (N_1968,N_1896,N_1918);
nor U1969 (N_1969,N_1906,N_1930);
nor U1970 (N_1970,N_1928,N_1898);
nor U1971 (N_1971,N_1895,N_1910);
nand U1972 (N_1972,N_1931,N_1925);
and U1973 (N_1973,N_1879,N_1888);
nand U1974 (N_1974,N_1908,N_1933);
nand U1975 (N_1975,N_1936,N_1929);
or U1976 (N_1976,N_1893,N_1946);
and U1977 (N_1977,N_1881,N_1890);
or U1978 (N_1978,N_1882,N_1913);
nor U1979 (N_1979,N_1935,N_1911);
or U1980 (N_1980,N_1885,N_1876);
and U1981 (N_1981,N_1905,N_1922);
nand U1982 (N_1982,N_1889,N_1941);
nor U1983 (N_1983,N_1912,N_1939);
nor U1984 (N_1984,N_1921,N_1907);
nand U1985 (N_1985,N_1909,N_1901);
nor U1986 (N_1986,N_1891,N_1949);
and U1987 (N_1987,N_1897,N_1887);
nor U1988 (N_1988,N_1886,N_1945);
or U1989 (N_1989,N_1946,N_1926);
or U1990 (N_1990,N_1923,N_1943);
nand U1991 (N_1991,N_1903,N_1942);
nor U1992 (N_1992,N_1879,N_1937);
nand U1993 (N_1993,N_1895,N_1886);
nand U1994 (N_1994,N_1919,N_1887);
nand U1995 (N_1995,N_1897,N_1902);
xor U1996 (N_1996,N_1938,N_1925);
nand U1997 (N_1997,N_1918,N_1898);
nor U1998 (N_1998,N_1923,N_1928);
or U1999 (N_1999,N_1933,N_1937);
xor U2000 (N_2000,N_1941,N_1933);
nand U2001 (N_2001,N_1939,N_1887);
and U2002 (N_2002,N_1886,N_1885);
or U2003 (N_2003,N_1891,N_1937);
or U2004 (N_2004,N_1889,N_1885);
nand U2005 (N_2005,N_1890,N_1876);
and U2006 (N_2006,N_1891,N_1927);
or U2007 (N_2007,N_1930,N_1927);
or U2008 (N_2008,N_1924,N_1892);
and U2009 (N_2009,N_1899,N_1920);
nand U2010 (N_2010,N_1897,N_1913);
nor U2011 (N_2011,N_1881,N_1906);
xnor U2012 (N_2012,N_1925,N_1898);
nor U2013 (N_2013,N_1878,N_1939);
nor U2014 (N_2014,N_1906,N_1918);
nor U2015 (N_2015,N_1929,N_1883);
nor U2016 (N_2016,N_1889,N_1949);
or U2017 (N_2017,N_1885,N_1915);
xor U2018 (N_2018,N_1949,N_1923);
or U2019 (N_2019,N_1936,N_1930);
or U2020 (N_2020,N_1941,N_1898);
xnor U2021 (N_2021,N_1900,N_1946);
or U2022 (N_2022,N_1933,N_1879);
and U2023 (N_2023,N_1911,N_1946);
and U2024 (N_2024,N_1906,N_1902);
or U2025 (N_2025,N_1986,N_2020);
and U2026 (N_2026,N_1994,N_2011);
or U2027 (N_2027,N_1966,N_1970);
and U2028 (N_2028,N_2008,N_2002);
nor U2029 (N_2029,N_2012,N_1995);
and U2030 (N_2030,N_1999,N_1991);
and U2031 (N_2031,N_1971,N_1982);
and U2032 (N_2032,N_1984,N_1960);
nand U2033 (N_2033,N_2017,N_2019);
nor U2034 (N_2034,N_1987,N_2004);
and U2035 (N_2035,N_1955,N_1989);
or U2036 (N_2036,N_2014,N_1977);
nor U2037 (N_2037,N_1964,N_1956);
nand U2038 (N_2038,N_1990,N_1958);
or U2039 (N_2039,N_1954,N_1965);
and U2040 (N_2040,N_1957,N_1951);
nor U2041 (N_2041,N_1998,N_1976);
nor U2042 (N_2042,N_2023,N_1996);
nor U2043 (N_2043,N_2005,N_2013);
nand U2044 (N_2044,N_1981,N_1993);
and U2045 (N_2045,N_1973,N_1988);
or U2046 (N_2046,N_2000,N_1969);
nand U2047 (N_2047,N_1992,N_1950);
or U2048 (N_2048,N_1959,N_1962);
nor U2049 (N_2049,N_1997,N_2018);
nand U2050 (N_2050,N_1974,N_2006);
and U2051 (N_2051,N_2021,N_1985);
or U2052 (N_2052,N_2001,N_1952);
and U2053 (N_2053,N_1963,N_1953);
nor U2054 (N_2054,N_2007,N_1961);
nand U2055 (N_2055,N_1980,N_1978);
nor U2056 (N_2056,N_2015,N_1968);
nor U2057 (N_2057,N_2024,N_1975);
nand U2058 (N_2058,N_1979,N_1967);
and U2059 (N_2059,N_2009,N_2022);
or U2060 (N_2060,N_2003,N_2010);
and U2061 (N_2061,N_1983,N_2016);
nand U2062 (N_2062,N_1972,N_1963);
xnor U2063 (N_2063,N_2008,N_1995);
or U2064 (N_2064,N_2019,N_1960);
and U2065 (N_2065,N_2017,N_1961);
nand U2066 (N_2066,N_1999,N_1964);
and U2067 (N_2067,N_1978,N_1950);
and U2068 (N_2068,N_2014,N_1951);
or U2069 (N_2069,N_1966,N_2001);
and U2070 (N_2070,N_1986,N_1996);
nor U2071 (N_2071,N_2011,N_1975);
and U2072 (N_2072,N_1976,N_1983);
nand U2073 (N_2073,N_1984,N_1978);
nor U2074 (N_2074,N_1980,N_2016);
or U2075 (N_2075,N_1975,N_1953);
nand U2076 (N_2076,N_2005,N_2024);
nor U2077 (N_2077,N_2001,N_1980);
or U2078 (N_2078,N_2014,N_2005);
xor U2079 (N_2079,N_2019,N_1972);
nor U2080 (N_2080,N_1965,N_1986);
or U2081 (N_2081,N_1963,N_2000);
nor U2082 (N_2082,N_1995,N_1968);
or U2083 (N_2083,N_1991,N_1988);
nor U2084 (N_2084,N_1967,N_2017);
and U2085 (N_2085,N_1962,N_1964);
or U2086 (N_2086,N_1986,N_1968);
and U2087 (N_2087,N_1981,N_1997);
or U2088 (N_2088,N_1992,N_1979);
xnor U2089 (N_2089,N_1991,N_1958);
nor U2090 (N_2090,N_2015,N_1987);
nor U2091 (N_2091,N_1985,N_2005);
and U2092 (N_2092,N_2008,N_1985);
nand U2093 (N_2093,N_1971,N_2011);
or U2094 (N_2094,N_2021,N_1972);
or U2095 (N_2095,N_1987,N_1968);
or U2096 (N_2096,N_1954,N_1973);
or U2097 (N_2097,N_2005,N_1957);
and U2098 (N_2098,N_2010,N_1987);
and U2099 (N_2099,N_2012,N_1960);
nor U2100 (N_2100,N_2037,N_2074);
nand U2101 (N_2101,N_2080,N_2058);
nor U2102 (N_2102,N_2078,N_2066);
nand U2103 (N_2103,N_2044,N_2030);
nand U2104 (N_2104,N_2051,N_2060);
nor U2105 (N_2105,N_2049,N_2027);
nand U2106 (N_2106,N_2055,N_2072);
or U2107 (N_2107,N_2068,N_2029);
or U2108 (N_2108,N_2031,N_2036);
or U2109 (N_2109,N_2077,N_2098);
nand U2110 (N_2110,N_2088,N_2057);
nor U2111 (N_2111,N_2048,N_2025);
and U2112 (N_2112,N_2033,N_2097);
and U2113 (N_2113,N_2092,N_2026);
and U2114 (N_2114,N_2040,N_2087);
nand U2115 (N_2115,N_2065,N_2071);
nor U2116 (N_2116,N_2038,N_2083);
or U2117 (N_2117,N_2089,N_2093);
nor U2118 (N_2118,N_2082,N_2042);
and U2119 (N_2119,N_2064,N_2073);
and U2120 (N_2120,N_2047,N_2032);
or U2121 (N_2121,N_2062,N_2053);
or U2122 (N_2122,N_2099,N_2035);
nand U2123 (N_2123,N_2069,N_2086);
nor U2124 (N_2124,N_2046,N_2067);
nand U2125 (N_2125,N_2070,N_2084);
or U2126 (N_2126,N_2045,N_2061);
nor U2127 (N_2127,N_2063,N_2050);
and U2128 (N_2128,N_2091,N_2034);
and U2129 (N_2129,N_2056,N_2094);
or U2130 (N_2130,N_2052,N_2076);
and U2131 (N_2131,N_2059,N_2096);
xnor U2132 (N_2132,N_2081,N_2075);
and U2133 (N_2133,N_2090,N_2095);
nor U2134 (N_2134,N_2039,N_2079);
or U2135 (N_2135,N_2028,N_2041);
nand U2136 (N_2136,N_2043,N_2054);
nor U2137 (N_2137,N_2085,N_2071);
nor U2138 (N_2138,N_2059,N_2054);
nor U2139 (N_2139,N_2091,N_2054);
xnor U2140 (N_2140,N_2052,N_2042);
and U2141 (N_2141,N_2088,N_2048);
and U2142 (N_2142,N_2048,N_2081);
nor U2143 (N_2143,N_2067,N_2096);
nor U2144 (N_2144,N_2077,N_2047);
and U2145 (N_2145,N_2032,N_2064);
nand U2146 (N_2146,N_2051,N_2056);
nor U2147 (N_2147,N_2078,N_2054);
nor U2148 (N_2148,N_2039,N_2065);
nand U2149 (N_2149,N_2070,N_2053);
or U2150 (N_2150,N_2044,N_2082);
xnor U2151 (N_2151,N_2080,N_2034);
or U2152 (N_2152,N_2098,N_2087);
and U2153 (N_2153,N_2026,N_2034);
nor U2154 (N_2154,N_2068,N_2033);
nor U2155 (N_2155,N_2068,N_2032);
nor U2156 (N_2156,N_2053,N_2049);
or U2157 (N_2157,N_2084,N_2048);
nand U2158 (N_2158,N_2090,N_2030);
and U2159 (N_2159,N_2078,N_2088);
nand U2160 (N_2160,N_2085,N_2093);
or U2161 (N_2161,N_2076,N_2093);
nand U2162 (N_2162,N_2071,N_2048);
nor U2163 (N_2163,N_2058,N_2040);
nand U2164 (N_2164,N_2051,N_2071);
and U2165 (N_2165,N_2090,N_2098);
nor U2166 (N_2166,N_2095,N_2045);
nor U2167 (N_2167,N_2032,N_2034);
or U2168 (N_2168,N_2075,N_2048);
nor U2169 (N_2169,N_2037,N_2040);
nor U2170 (N_2170,N_2055,N_2098);
nand U2171 (N_2171,N_2048,N_2079);
nor U2172 (N_2172,N_2064,N_2031);
nor U2173 (N_2173,N_2065,N_2069);
nor U2174 (N_2174,N_2079,N_2081);
nand U2175 (N_2175,N_2119,N_2169);
nor U2176 (N_2176,N_2154,N_2149);
and U2177 (N_2177,N_2144,N_2153);
nor U2178 (N_2178,N_2129,N_2114);
nand U2179 (N_2179,N_2107,N_2132);
or U2180 (N_2180,N_2142,N_2171);
or U2181 (N_2181,N_2159,N_2137);
nand U2182 (N_2182,N_2150,N_2160);
nor U2183 (N_2183,N_2115,N_2166);
nor U2184 (N_2184,N_2148,N_2124);
nand U2185 (N_2185,N_2157,N_2128);
xnor U2186 (N_2186,N_2111,N_2109);
or U2187 (N_2187,N_2112,N_2162);
nor U2188 (N_2188,N_2102,N_2131);
and U2189 (N_2189,N_2127,N_2161);
or U2190 (N_2190,N_2134,N_2126);
nand U2191 (N_2191,N_2172,N_2151);
and U2192 (N_2192,N_2135,N_2106);
nor U2193 (N_2193,N_2141,N_2100);
and U2194 (N_2194,N_2167,N_2123);
and U2195 (N_2195,N_2113,N_2139);
nand U2196 (N_2196,N_2147,N_2140);
or U2197 (N_2197,N_2103,N_2163);
nand U2198 (N_2198,N_2122,N_2105);
nor U2199 (N_2199,N_2133,N_2143);
and U2200 (N_2200,N_2138,N_2125);
nand U2201 (N_2201,N_2104,N_2145);
nand U2202 (N_2202,N_2174,N_2121);
or U2203 (N_2203,N_2146,N_2118);
and U2204 (N_2204,N_2120,N_2155);
nand U2205 (N_2205,N_2158,N_2136);
and U2206 (N_2206,N_2173,N_2108);
xor U2207 (N_2207,N_2164,N_2130);
nand U2208 (N_2208,N_2116,N_2156);
or U2209 (N_2209,N_2152,N_2110);
or U2210 (N_2210,N_2168,N_2170);
nand U2211 (N_2211,N_2165,N_2117);
or U2212 (N_2212,N_2101,N_2112);
or U2213 (N_2213,N_2166,N_2153);
nor U2214 (N_2214,N_2114,N_2103);
nand U2215 (N_2215,N_2134,N_2157);
or U2216 (N_2216,N_2105,N_2144);
nand U2217 (N_2217,N_2103,N_2128);
or U2218 (N_2218,N_2119,N_2132);
nor U2219 (N_2219,N_2158,N_2107);
or U2220 (N_2220,N_2172,N_2116);
nor U2221 (N_2221,N_2147,N_2145);
nand U2222 (N_2222,N_2112,N_2146);
nor U2223 (N_2223,N_2117,N_2160);
and U2224 (N_2224,N_2152,N_2102);
and U2225 (N_2225,N_2160,N_2143);
or U2226 (N_2226,N_2120,N_2100);
nand U2227 (N_2227,N_2123,N_2160);
and U2228 (N_2228,N_2103,N_2126);
and U2229 (N_2229,N_2165,N_2137);
or U2230 (N_2230,N_2145,N_2114);
and U2231 (N_2231,N_2118,N_2100);
nor U2232 (N_2232,N_2141,N_2164);
nor U2233 (N_2233,N_2106,N_2121);
nand U2234 (N_2234,N_2160,N_2130);
and U2235 (N_2235,N_2169,N_2113);
nand U2236 (N_2236,N_2160,N_2135);
or U2237 (N_2237,N_2172,N_2141);
and U2238 (N_2238,N_2150,N_2161);
nand U2239 (N_2239,N_2155,N_2115);
or U2240 (N_2240,N_2123,N_2151);
and U2241 (N_2241,N_2129,N_2149);
or U2242 (N_2242,N_2118,N_2110);
nor U2243 (N_2243,N_2113,N_2164);
or U2244 (N_2244,N_2109,N_2103);
nor U2245 (N_2245,N_2167,N_2128);
nand U2246 (N_2246,N_2139,N_2126);
and U2247 (N_2247,N_2111,N_2158);
and U2248 (N_2248,N_2111,N_2168);
xnor U2249 (N_2249,N_2102,N_2167);
nand U2250 (N_2250,N_2236,N_2207);
or U2251 (N_2251,N_2239,N_2249);
nand U2252 (N_2252,N_2196,N_2213);
nand U2253 (N_2253,N_2218,N_2188);
nand U2254 (N_2254,N_2220,N_2203);
or U2255 (N_2255,N_2202,N_2198);
xor U2256 (N_2256,N_2215,N_2238);
and U2257 (N_2257,N_2235,N_2176);
xor U2258 (N_2258,N_2241,N_2180);
nor U2259 (N_2259,N_2248,N_2204);
or U2260 (N_2260,N_2191,N_2222);
xor U2261 (N_2261,N_2209,N_2178);
or U2262 (N_2262,N_2217,N_2190);
or U2263 (N_2263,N_2189,N_2184);
nand U2264 (N_2264,N_2185,N_2197);
nor U2265 (N_2265,N_2186,N_2234);
nor U2266 (N_2266,N_2247,N_2230);
nand U2267 (N_2267,N_2245,N_2175);
or U2268 (N_2268,N_2226,N_2242);
or U2269 (N_2269,N_2246,N_2206);
nor U2270 (N_2270,N_2221,N_2182);
or U2271 (N_2271,N_2199,N_2179);
nor U2272 (N_2272,N_2211,N_2240);
nand U2273 (N_2273,N_2212,N_2229);
nand U2274 (N_2274,N_2194,N_2223);
nor U2275 (N_2275,N_2231,N_2214);
nor U2276 (N_2276,N_2193,N_2244);
nand U2277 (N_2277,N_2225,N_2227);
nor U2278 (N_2278,N_2243,N_2210);
nor U2279 (N_2279,N_2219,N_2201);
and U2280 (N_2280,N_2228,N_2195);
nor U2281 (N_2281,N_2181,N_2233);
or U2282 (N_2282,N_2200,N_2205);
nor U2283 (N_2283,N_2216,N_2183);
and U2284 (N_2284,N_2177,N_2232);
and U2285 (N_2285,N_2208,N_2237);
nor U2286 (N_2286,N_2187,N_2224);
nand U2287 (N_2287,N_2192,N_2236);
nor U2288 (N_2288,N_2189,N_2223);
and U2289 (N_2289,N_2203,N_2179);
xnor U2290 (N_2290,N_2220,N_2196);
and U2291 (N_2291,N_2239,N_2209);
nand U2292 (N_2292,N_2183,N_2236);
nor U2293 (N_2293,N_2233,N_2176);
and U2294 (N_2294,N_2200,N_2201);
nor U2295 (N_2295,N_2206,N_2182);
nand U2296 (N_2296,N_2243,N_2197);
and U2297 (N_2297,N_2228,N_2194);
and U2298 (N_2298,N_2189,N_2227);
and U2299 (N_2299,N_2191,N_2175);
and U2300 (N_2300,N_2241,N_2184);
and U2301 (N_2301,N_2184,N_2201);
or U2302 (N_2302,N_2229,N_2243);
nand U2303 (N_2303,N_2186,N_2192);
nand U2304 (N_2304,N_2207,N_2226);
and U2305 (N_2305,N_2209,N_2197);
or U2306 (N_2306,N_2230,N_2248);
nor U2307 (N_2307,N_2189,N_2245);
or U2308 (N_2308,N_2229,N_2192);
nand U2309 (N_2309,N_2176,N_2215);
or U2310 (N_2310,N_2178,N_2222);
or U2311 (N_2311,N_2216,N_2235);
nand U2312 (N_2312,N_2204,N_2234);
nor U2313 (N_2313,N_2183,N_2239);
nor U2314 (N_2314,N_2224,N_2183);
nor U2315 (N_2315,N_2197,N_2232);
nand U2316 (N_2316,N_2185,N_2230);
xnor U2317 (N_2317,N_2231,N_2208);
or U2318 (N_2318,N_2232,N_2204);
or U2319 (N_2319,N_2197,N_2244);
nand U2320 (N_2320,N_2238,N_2245);
and U2321 (N_2321,N_2212,N_2184);
and U2322 (N_2322,N_2175,N_2240);
nor U2323 (N_2323,N_2212,N_2211);
and U2324 (N_2324,N_2175,N_2212);
nand U2325 (N_2325,N_2258,N_2278);
or U2326 (N_2326,N_2321,N_2299);
or U2327 (N_2327,N_2314,N_2269);
or U2328 (N_2328,N_2271,N_2276);
nor U2329 (N_2329,N_2302,N_2265);
or U2330 (N_2330,N_2261,N_2290);
and U2331 (N_2331,N_2316,N_2268);
or U2332 (N_2332,N_2295,N_2280);
nor U2333 (N_2333,N_2311,N_2272);
xor U2334 (N_2334,N_2294,N_2322);
or U2335 (N_2335,N_2293,N_2313);
and U2336 (N_2336,N_2323,N_2301);
nand U2337 (N_2337,N_2250,N_2273);
nand U2338 (N_2338,N_2285,N_2281);
nand U2339 (N_2339,N_2267,N_2309);
and U2340 (N_2340,N_2312,N_2318);
and U2341 (N_2341,N_2296,N_2315);
and U2342 (N_2342,N_2270,N_2298);
nor U2343 (N_2343,N_2308,N_2279);
or U2344 (N_2344,N_2304,N_2300);
or U2345 (N_2345,N_2266,N_2254);
or U2346 (N_2346,N_2287,N_2324);
nand U2347 (N_2347,N_2277,N_2310);
and U2348 (N_2348,N_2259,N_2256);
nor U2349 (N_2349,N_2255,N_2284);
nor U2350 (N_2350,N_2307,N_2289);
and U2351 (N_2351,N_2317,N_2292);
nor U2352 (N_2352,N_2260,N_2291);
or U2353 (N_2353,N_2288,N_2320);
nor U2354 (N_2354,N_2257,N_2297);
nor U2355 (N_2355,N_2319,N_2282);
xnor U2356 (N_2356,N_2275,N_2306);
nor U2357 (N_2357,N_2303,N_2274);
and U2358 (N_2358,N_2305,N_2263);
nor U2359 (N_2359,N_2253,N_2262);
nor U2360 (N_2360,N_2252,N_2251);
xor U2361 (N_2361,N_2264,N_2283);
or U2362 (N_2362,N_2286,N_2273);
nor U2363 (N_2363,N_2258,N_2274);
nand U2364 (N_2364,N_2270,N_2312);
or U2365 (N_2365,N_2280,N_2261);
nand U2366 (N_2366,N_2314,N_2288);
nand U2367 (N_2367,N_2285,N_2293);
and U2368 (N_2368,N_2281,N_2260);
nand U2369 (N_2369,N_2324,N_2263);
and U2370 (N_2370,N_2308,N_2307);
nor U2371 (N_2371,N_2295,N_2307);
nor U2372 (N_2372,N_2307,N_2320);
nand U2373 (N_2373,N_2291,N_2294);
and U2374 (N_2374,N_2271,N_2253);
nor U2375 (N_2375,N_2285,N_2296);
or U2376 (N_2376,N_2252,N_2313);
nor U2377 (N_2377,N_2269,N_2276);
nand U2378 (N_2378,N_2301,N_2290);
or U2379 (N_2379,N_2255,N_2315);
nand U2380 (N_2380,N_2250,N_2324);
or U2381 (N_2381,N_2265,N_2251);
nor U2382 (N_2382,N_2313,N_2322);
or U2383 (N_2383,N_2279,N_2258);
or U2384 (N_2384,N_2312,N_2267);
nor U2385 (N_2385,N_2258,N_2308);
nand U2386 (N_2386,N_2269,N_2287);
nand U2387 (N_2387,N_2275,N_2250);
nor U2388 (N_2388,N_2271,N_2307);
nand U2389 (N_2389,N_2289,N_2291);
nor U2390 (N_2390,N_2256,N_2307);
nor U2391 (N_2391,N_2291,N_2252);
and U2392 (N_2392,N_2258,N_2266);
and U2393 (N_2393,N_2318,N_2252);
xor U2394 (N_2394,N_2279,N_2273);
and U2395 (N_2395,N_2258,N_2252);
nor U2396 (N_2396,N_2284,N_2256);
xnor U2397 (N_2397,N_2276,N_2314);
or U2398 (N_2398,N_2297,N_2296);
xnor U2399 (N_2399,N_2294,N_2263);
or U2400 (N_2400,N_2342,N_2372);
or U2401 (N_2401,N_2382,N_2358);
nand U2402 (N_2402,N_2356,N_2352);
and U2403 (N_2403,N_2350,N_2349);
or U2404 (N_2404,N_2376,N_2345);
and U2405 (N_2405,N_2395,N_2346);
nor U2406 (N_2406,N_2326,N_2369);
nand U2407 (N_2407,N_2393,N_2386);
and U2408 (N_2408,N_2370,N_2387);
or U2409 (N_2409,N_2399,N_2366);
nor U2410 (N_2410,N_2353,N_2340);
nor U2411 (N_2411,N_2341,N_2329);
and U2412 (N_2412,N_2359,N_2368);
nor U2413 (N_2413,N_2365,N_2347);
and U2414 (N_2414,N_2357,N_2383);
nor U2415 (N_2415,N_2379,N_2396);
and U2416 (N_2416,N_2333,N_2392);
nor U2417 (N_2417,N_2331,N_2348);
nand U2418 (N_2418,N_2330,N_2385);
nand U2419 (N_2419,N_2328,N_2390);
or U2420 (N_2420,N_2375,N_2384);
and U2421 (N_2421,N_2327,N_2371);
nand U2422 (N_2422,N_2363,N_2374);
xnor U2423 (N_2423,N_2391,N_2380);
and U2424 (N_2424,N_2373,N_2360);
nor U2425 (N_2425,N_2377,N_2337);
and U2426 (N_2426,N_2378,N_2351);
and U2427 (N_2427,N_2394,N_2398);
nand U2428 (N_2428,N_2335,N_2397);
and U2429 (N_2429,N_2336,N_2388);
or U2430 (N_2430,N_2332,N_2362);
nor U2431 (N_2431,N_2389,N_2344);
nand U2432 (N_2432,N_2334,N_2361);
nor U2433 (N_2433,N_2343,N_2338);
and U2434 (N_2434,N_2364,N_2354);
or U2435 (N_2435,N_2339,N_2381);
xnor U2436 (N_2436,N_2355,N_2325);
xnor U2437 (N_2437,N_2367,N_2332);
and U2438 (N_2438,N_2362,N_2395);
or U2439 (N_2439,N_2383,N_2372);
and U2440 (N_2440,N_2348,N_2369);
and U2441 (N_2441,N_2325,N_2384);
and U2442 (N_2442,N_2368,N_2386);
and U2443 (N_2443,N_2340,N_2376);
nor U2444 (N_2444,N_2330,N_2381);
nor U2445 (N_2445,N_2340,N_2360);
nor U2446 (N_2446,N_2339,N_2335);
nand U2447 (N_2447,N_2350,N_2386);
or U2448 (N_2448,N_2380,N_2352);
or U2449 (N_2449,N_2349,N_2373);
or U2450 (N_2450,N_2383,N_2381);
or U2451 (N_2451,N_2362,N_2388);
and U2452 (N_2452,N_2331,N_2361);
nor U2453 (N_2453,N_2351,N_2360);
and U2454 (N_2454,N_2347,N_2383);
and U2455 (N_2455,N_2393,N_2345);
nand U2456 (N_2456,N_2397,N_2399);
or U2457 (N_2457,N_2339,N_2329);
or U2458 (N_2458,N_2332,N_2385);
or U2459 (N_2459,N_2358,N_2356);
and U2460 (N_2460,N_2356,N_2340);
nor U2461 (N_2461,N_2336,N_2364);
nand U2462 (N_2462,N_2354,N_2334);
nand U2463 (N_2463,N_2372,N_2398);
nor U2464 (N_2464,N_2356,N_2330);
and U2465 (N_2465,N_2386,N_2362);
and U2466 (N_2466,N_2334,N_2332);
and U2467 (N_2467,N_2368,N_2329);
and U2468 (N_2468,N_2350,N_2371);
nor U2469 (N_2469,N_2325,N_2386);
or U2470 (N_2470,N_2395,N_2393);
or U2471 (N_2471,N_2344,N_2399);
and U2472 (N_2472,N_2358,N_2377);
nand U2473 (N_2473,N_2384,N_2386);
nand U2474 (N_2474,N_2337,N_2384);
nand U2475 (N_2475,N_2428,N_2418);
or U2476 (N_2476,N_2446,N_2461);
and U2477 (N_2477,N_2450,N_2470);
nand U2478 (N_2478,N_2406,N_2465);
nor U2479 (N_2479,N_2429,N_2443);
and U2480 (N_2480,N_2468,N_2441);
or U2481 (N_2481,N_2456,N_2473);
or U2482 (N_2482,N_2436,N_2411);
nand U2483 (N_2483,N_2474,N_2449);
or U2484 (N_2484,N_2419,N_2434);
and U2485 (N_2485,N_2405,N_2422);
and U2486 (N_2486,N_2442,N_2431);
nor U2487 (N_2487,N_2464,N_2439);
or U2488 (N_2488,N_2421,N_2467);
xor U2489 (N_2489,N_2425,N_2471);
and U2490 (N_2490,N_2432,N_2417);
and U2491 (N_2491,N_2435,N_2433);
nand U2492 (N_2492,N_2407,N_2451);
or U2493 (N_2493,N_2424,N_2440);
or U2494 (N_2494,N_2454,N_2415);
nand U2495 (N_2495,N_2472,N_2402);
nand U2496 (N_2496,N_2408,N_2469);
or U2497 (N_2497,N_2409,N_2448);
xnor U2498 (N_2498,N_2414,N_2430);
nor U2499 (N_2499,N_2452,N_2457);
or U2500 (N_2500,N_2412,N_2410);
and U2501 (N_2501,N_2458,N_2413);
and U2502 (N_2502,N_2466,N_2453);
and U2503 (N_2503,N_2437,N_2462);
xnor U2504 (N_2504,N_2416,N_2438);
and U2505 (N_2505,N_2447,N_2460);
or U2506 (N_2506,N_2403,N_2426);
or U2507 (N_2507,N_2420,N_2444);
nand U2508 (N_2508,N_2423,N_2401);
nor U2509 (N_2509,N_2455,N_2459);
nor U2510 (N_2510,N_2404,N_2463);
nor U2511 (N_2511,N_2445,N_2400);
nand U2512 (N_2512,N_2427,N_2441);
or U2513 (N_2513,N_2447,N_2406);
and U2514 (N_2514,N_2430,N_2434);
and U2515 (N_2515,N_2410,N_2451);
nand U2516 (N_2516,N_2410,N_2471);
or U2517 (N_2517,N_2417,N_2413);
xnor U2518 (N_2518,N_2434,N_2435);
nor U2519 (N_2519,N_2444,N_2428);
and U2520 (N_2520,N_2434,N_2463);
or U2521 (N_2521,N_2452,N_2424);
and U2522 (N_2522,N_2460,N_2469);
and U2523 (N_2523,N_2466,N_2407);
or U2524 (N_2524,N_2460,N_2408);
nand U2525 (N_2525,N_2457,N_2437);
and U2526 (N_2526,N_2439,N_2457);
nand U2527 (N_2527,N_2441,N_2444);
and U2528 (N_2528,N_2400,N_2451);
and U2529 (N_2529,N_2472,N_2474);
nor U2530 (N_2530,N_2400,N_2438);
and U2531 (N_2531,N_2453,N_2414);
or U2532 (N_2532,N_2469,N_2429);
and U2533 (N_2533,N_2419,N_2455);
or U2534 (N_2534,N_2424,N_2469);
nand U2535 (N_2535,N_2412,N_2446);
nor U2536 (N_2536,N_2406,N_2454);
nor U2537 (N_2537,N_2452,N_2449);
and U2538 (N_2538,N_2426,N_2462);
nor U2539 (N_2539,N_2412,N_2454);
nand U2540 (N_2540,N_2472,N_2451);
and U2541 (N_2541,N_2459,N_2437);
xor U2542 (N_2542,N_2411,N_2417);
nand U2543 (N_2543,N_2464,N_2407);
nor U2544 (N_2544,N_2438,N_2423);
and U2545 (N_2545,N_2458,N_2407);
nor U2546 (N_2546,N_2450,N_2414);
xor U2547 (N_2547,N_2429,N_2400);
or U2548 (N_2548,N_2451,N_2465);
nand U2549 (N_2549,N_2408,N_2429);
or U2550 (N_2550,N_2525,N_2476);
and U2551 (N_2551,N_2549,N_2516);
nor U2552 (N_2552,N_2539,N_2508);
nor U2553 (N_2553,N_2523,N_2510);
and U2554 (N_2554,N_2520,N_2493);
nor U2555 (N_2555,N_2489,N_2500);
nand U2556 (N_2556,N_2530,N_2488);
nor U2557 (N_2557,N_2502,N_2546);
or U2558 (N_2558,N_2513,N_2548);
and U2559 (N_2559,N_2533,N_2487);
and U2560 (N_2560,N_2521,N_2529);
nor U2561 (N_2561,N_2503,N_2496);
and U2562 (N_2562,N_2486,N_2532);
nand U2563 (N_2563,N_2538,N_2505);
nor U2564 (N_2564,N_2535,N_2477);
and U2565 (N_2565,N_2483,N_2484);
or U2566 (N_2566,N_2542,N_2515);
nand U2567 (N_2567,N_2544,N_2537);
or U2568 (N_2568,N_2527,N_2495);
or U2569 (N_2569,N_2545,N_2501);
nor U2570 (N_2570,N_2517,N_2482);
or U2571 (N_2571,N_2512,N_2481);
xnor U2572 (N_2572,N_2524,N_2504);
nand U2573 (N_2573,N_2509,N_2531);
and U2574 (N_2574,N_2528,N_2511);
nand U2575 (N_2575,N_2547,N_2506);
nor U2576 (N_2576,N_2499,N_2494);
or U2577 (N_2577,N_2479,N_2507);
or U2578 (N_2578,N_2480,N_2478);
nand U2579 (N_2579,N_2518,N_2540);
nor U2580 (N_2580,N_2492,N_2522);
nand U2581 (N_2581,N_2497,N_2519);
nand U2582 (N_2582,N_2526,N_2543);
or U2583 (N_2583,N_2475,N_2485);
nand U2584 (N_2584,N_2498,N_2514);
and U2585 (N_2585,N_2490,N_2491);
nand U2586 (N_2586,N_2536,N_2534);
nor U2587 (N_2587,N_2541,N_2529);
and U2588 (N_2588,N_2514,N_2528);
nor U2589 (N_2589,N_2520,N_2488);
nand U2590 (N_2590,N_2502,N_2503);
nor U2591 (N_2591,N_2540,N_2535);
nand U2592 (N_2592,N_2515,N_2499);
nand U2593 (N_2593,N_2540,N_2502);
or U2594 (N_2594,N_2483,N_2478);
nor U2595 (N_2595,N_2540,N_2507);
nand U2596 (N_2596,N_2526,N_2519);
or U2597 (N_2597,N_2490,N_2519);
or U2598 (N_2598,N_2539,N_2511);
nand U2599 (N_2599,N_2501,N_2520);
or U2600 (N_2600,N_2480,N_2522);
or U2601 (N_2601,N_2500,N_2509);
and U2602 (N_2602,N_2523,N_2518);
or U2603 (N_2603,N_2485,N_2519);
or U2604 (N_2604,N_2526,N_2522);
nor U2605 (N_2605,N_2502,N_2535);
and U2606 (N_2606,N_2488,N_2484);
or U2607 (N_2607,N_2519,N_2488);
or U2608 (N_2608,N_2490,N_2547);
nand U2609 (N_2609,N_2530,N_2516);
or U2610 (N_2610,N_2541,N_2511);
nand U2611 (N_2611,N_2499,N_2534);
and U2612 (N_2612,N_2487,N_2480);
or U2613 (N_2613,N_2547,N_2521);
nor U2614 (N_2614,N_2507,N_2526);
or U2615 (N_2615,N_2543,N_2482);
nor U2616 (N_2616,N_2530,N_2535);
nor U2617 (N_2617,N_2478,N_2531);
or U2618 (N_2618,N_2537,N_2475);
and U2619 (N_2619,N_2488,N_2487);
and U2620 (N_2620,N_2520,N_2532);
nor U2621 (N_2621,N_2500,N_2504);
and U2622 (N_2622,N_2501,N_2536);
or U2623 (N_2623,N_2480,N_2511);
or U2624 (N_2624,N_2516,N_2528);
xor U2625 (N_2625,N_2597,N_2621);
nor U2626 (N_2626,N_2578,N_2592);
and U2627 (N_2627,N_2573,N_2618);
nor U2628 (N_2628,N_2607,N_2622);
or U2629 (N_2629,N_2594,N_2577);
and U2630 (N_2630,N_2611,N_2596);
nor U2631 (N_2631,N_2609,N_2563);
nand U2632 (N_2632,N_2608,N_2600);
nand U2633 (N_2633,N_2624,N_2613);
nand U2634 (N_2634,N_2620,N_2583);
or U2635 (N_2635,N_2561,N_2551);
nand U2636 (N_2636,N_2555,N_2554);
and U2637 (N_2637,N_2623,N_2605);
nor U2638 (N_2638,N_2556,N_2567);
nor U2639 (N_2639,N_2616,N_2590);
nor U2640 (N_2640,N_2598,N_2619);
nor U2641 (N_2641,N_2581,N_2585);
nand U2642 (N_2642,N_2569,N_2574);
xor U2643 (N_2643,N_2571,N_2593);
and U2644 (N_2644,N_2553,N_2566);
nor U2645 (N_2645,N_2617,N_2599);
and U2646 (N_2646,N_2601,N_2612);
or U2647 (N_2647,N_2564,N_2557);
or U2648 (N_2648,N_2602,N_2575);
nand U2649 (N_2649,N_2588,N_2604);
and U2650 (N_2650,N_2603,N_2582);
and U2651 (N_2651,N_2559,N_2589);
or U2652 (N_2652,N_2610,N_2562);
nand U2653 (N_2653,N_2552,N_2572);
or U2654 (N_2654,N_2576,N_2565);
or U2655 (N_2655,N_2579,N_2615);
and U2656 (N_2656,N_2606,N_2584);
or U2657 (N_2657,N_2614,N_2595);
or U2658 (N_2658,N_2591,N_2560);
or U2659 (N_2659,N_2558,N_2570);
and U2660 (N_2660,N_2568,N_2550);
nor U2661 (N_2661,N_2587,N_2580);
nor U2662 (N_2662,N_2586,N_2596);
nor U2663 (N_2663,N_2561,N_2600);
nand U2664 (N_2664,N_2577,N_2598);
nor U2665 (N_2665,N_2582,N_2618);
nor U2666 (N_2666,N_2581,N_2567);
and U2667 (N_2667,N_2553,N_2594);
nor U2668 (N_2668,N_2604,N_2590);
or U2669 (N_2669,N_2581,N_2572);
and U2670 (N_2670,N_2574,N_2602);
or U2671 (N_2671,N_2614,N_2552);
and U2672 (N_2672,N_2586,N_2579);
nor U2673 (N_2673,N_2616,N_2600);
nand U2674 (N_2674,N_2606,N_2564);
nor U2675 (N_2675,N_2609,N_2586);
and U2676 (N_2676,N_2620,N_2567);
or U2677 (N_2677,N_2619,N_2590);
or U2678 (N_2678,N_2613,N_2578);
or U2679 (N_2679,N_2622,N_2614);
nor U2680 (N_2680,N_2555,N_2613);
and U2681 (N_2681,N_2579,N_2552);
or U2682 (N_2682,N_2578,N_2603);
or U2683 (N_2683,N_2607,N_2551);
and U2684 (N_2684,N_2623,N_2587);
or U2685 (N_2685,N_2551,N_2564);
nand U2686 (N_2686,N_2620,N_2572);
nand U2687 (N_2687,N_2621,N_2587);
nor U2688 (N_2688,N_2585,N_2587);
and U2689 (N_2689,N_2595,N_2575);
nor U2690 (N_2690,N_2563,N_2619);
nor U2691 (N_2691,N_2599,N_2622);
and U2692 (N_2692,N_2616,N_2581);
and U2693 (N_2693,N_2573,N_2593);
or U2694 (N_2694,N_2621,N_2569);
nand U2695 (N_2695,N_2603,N_2606);
or U2696 (N_2696,N_2614,N_2617);
or U2697 (N_2697,N_2553,N_2589);
and U2698 (N_2698,N_2614,N_2577);
nor U2699 (N_2699,N_2623,N_2552);
nor U2700 (N_2700,N_2655,N_2645);
nor U2701 (N_2701,N_2652,N_2659);
or U2702 (N_2702,N_2666,N_2634);
or U2703 (N_2703,N_2693,N_2653);
and U2704 (N_2704,N_2632,N_2680);
nor U2705 (N_2705,N_2674,N_2679);
nand U2706 (N_2706,N_2638,N_2644);
nor U2707 (N_2707,N_2654,N_2629);
nor U2708 (N_2708,N_2665,N_2688);
xor U2709 (N_2709,N_2663,N_2656);
xnor U2710 (N_2710,N_2668,N_2628);
nand U2711 (N_2711,N_2643,N_2677);
and U2712 (N_2712,N_2670,N_2630);
nand U2713 (N_2713,N_2687,N_2646);
nor U2714 (N_2714,N_2637,N_2691);
nand U2715 (N_2715,N_2694,N_2698);
or U2716 (N_2716,N_2633,N_2650);
nor U2717 (N_2717,N_2642,N_2641);
nor U2718 (N_2718,N_2664,N_2673);
nor U2719 (N_2719,N_2627,N_2626);
and U2720 (N_2720,N_2675,N_2636);
nor U2721 (N_2721,N_2671,N_2696);
and U2722 (N_2722,N_2662,N_2635);
xnor U2723 (N_2723,N_2686,N_2661);
nand U2724 (N_2724,N_2648,N_2682);
and U2725 (N_2725,N_2651,N_2690);
nand U2726 (N_2726,N_2685,N_2678);
or U2727 (N_2727,N_2689,N_2699);
nand U2728 (N_2728,N_2695,N_2660);
nand U2729 (N_2729,N_2658,N_2639);
and U2730 (N_2730,N_2647,N_2657);
or U2731 (N_2731,N_2684,N_2631);
nor U2732 (N_2732,N_2640,N_2692);
nor U2733 (N_2733,N_2697,N_2681);
or U2734 (N_2734,N_2672,N_2683);
xor U2735 (N_2735,N_2625,N_2676);
or U2736 (N_2736,N_2649,N_2667);
xor U2737 (N_2737,N_2669,N_2648);
or U2738 (N_2738,N_2637,N_2678);
or U2739 (N_2739,N_2693,N_2668);
nor U2740 (N_2740,N_2659,N_2647);
or U2741 (N_2741,N_2688,N_2684);
or U2742 (N_2742,N_2656,N_2699);
or U2743 (N_2743,N_2636,N_2641);
nand U2744 (N_2744,N_2640,N_2642);
nand U2745 (N_2745,N_2642,N_2693);
xor U2746 (N_2746,N_2697,N_2694);
nor U2747 (N_2747,N_2642,N_2645);
nand U2748 (N_2748,N_2698,N_2640);
or U2749 (N_2749,N_2694,N_2680);
xor U2750 (N_2750,N_2649,N_2690);
nor U2751 (N_2751,N_2652,N_2657);
or U2752 (N_2752,N_2655,N_2682);
or U2753 (N_2753,N_2687,N_2660);
nand U2754 (N_2754,N_2664,N_2631);
nand U2755 (N_2755,N_2671,N_2667);
nor U2756 (N_2756,N_2660,N_2663);
or U2757 (N_2757,N_2688,N_2657);
and U2758 (N_2758,N_2671,N_2694);
or U2759 (N_2759,N_2695,N_2639);
nor U2760 (N_2760,N_2685,N_2636);
nand U2761 (N_2761,N_2651,N_2682);
or U2762 (N_2762,N_2635,N_2686);
nand U2763 (N_2763,N_2650,N_2636);
nand U2764 (N_2764,N_2664,N_2663);
and U2765 (N_2765,N_2687,N_2629);
nand U2766 (N_2766,N_2638,N_2627);
or U2767 (N_2767,N_2661,N_2690);
or U2768 (N_2768,N_2652,N_2664);
nand U2769 (N_2769,N_2689,N_2675);
and U2770 (N_2770,N_2658,N_2699);
nand U2771 (N_2771,N_2658,N_2694);
or U2772 (N_2772,N_2638,N_2628);
nand U2773 (N_2773,N_2652,N_2699);
or U2774 (N_2774,N_2681,N_2666);
and U2775 (N_2775,N_2709,N_2713);
nor U2776 (N_2776,N_2758,N_2768);
nand U2777 (N_2777,N_2773,N_2718);
nand U2778 (N_2778,N_2763,N_2741);
and U2779 (N_2779,N_2737,N_2700);
and U2780 (N_2780,N_2717,N_2732);
nor U2781 (N_2781,N_2712,N_2749);
or U2782 (N_2782,N_2747,N_2769);
nand U2783 (N_2783,N_2754,N_2743);
nor U2784 (N_2784,N_2745,N_2727);
and U2785 (N_2785,N_2735,N_2711);
nand U2786 (N_2786,N_2724,N_2723);
nand U2787 (N_2787,N_2729,N_2707);
or U2788 (N_2788,N_2719,N_2703);
or U2789 (N_2789,N_2744,N_2752);
nor U2790 (N_2790,N_2725,N_2731);
and U2791 (N_2791,N_2738,N_2757);
nand U2792 (N_2792,N_2753,N_2755);
or U2793 (N_2793,N_2739,N_2726);
and U2794 (N_2794,N_2760,N_2736);
nand U2795 (N_2795,N_2710,N_2733);
nor U2796 (N_2796,N_2748,N_2730);
nor U2797 (N_2797,N_2746,N_2764);
and U2798 (N_2798,N_2721,N_2720);
nand U2799 (N_2799,N_2759,N_2716);
or U2800 (N_2800,N_2770,N_2742);
xor U2801 (N_2801,N_2772,N_2722);
nand U2802 (N_2802,N_2715,N_2762);
and U2803 (N_2803,N_2701,N_2756);
nor U2804 (N_2804,N_2728,N_2771);
nor U2805 (N_2805,N_2702,N_2767);
nor U2806 (N_2806,N_2766,N_2765);
and U2807 (N_2807,N_2751,N_2704);
and U2808 (N_2808,N_2774,N_2740);
nand U2809 (N_2809,N_2750,N_2705);
and U2810 (N_2810,N_2714,N_2708);
nor U2811 (N_2811,N_2706,N_2734);
or U2812 (N_2812,N_2761,N_2773);
nand U2813 (N_2813,N_2705,N_2719);
and U2814 (N_2814,N_2747,N_2771);
or U2815 (N_2815,N_2707,N_2709);
nor U2816 (N_2816,N_2745,N_2761);
xnor U2817 (N_2817,N_2756,N_2702);
or U2818 (N_2818,N_2769,N_2731);
nor U2819 (N_2819,N_2751,N_2764);
and U2820 (N_2820,N_2770,N_2740);
nor U2821 (N_2821,N_2725,N_2736);
nand U2822 (N_2822,N_2736,N_2716);
nor U2823 (N_2823,N_2700,N_2716);
or U2824 (N_2824,N_2710,N_2736);
or U2825 (N_2825,N_2744,N_2750);
nor U2826 (N_2826,N_2707,N_2754);
or U2827 (N_2827,N_2752,N_2700);
nor U2828 (N_2828,N_2703,N_2742);
and U2829 (N_2829,N_2715,N_2736);
and U2830 (N_2830,N_2732,N_2765);
xnor U2831 (N_2831,N_2731,N_2743);
nor U2832 (N_2832,N_2774,N_2750);
and U2833 (N_2833,N_2740,N_2711);
nor U2834 (N_2834,N_2701,N_2762);
or U2835 (N_2835,N_2742,N_2734);
or U2836 (N_2836,N_2746,N_2768);
and U2837 (N_2837,N_2740,N_2771);
or U2838 (N_2838,N_2764,N_2723);
and U2839 (N_2839,N_2702,N_2733);
nand U2840 (N_2840,N_2713,N_2753);
nand U2841 (N_2841,N_2739,N_2736);
nor U2842 (N_2842,N_2759,N_2711);
nor U2843 (N_2843,N_2739,N_2710);
or U2844 (N_2844,N_2747,N_2706);
and U2845 (N_2845,N_2731,N_2765);
and U2846 (N_2846,N_2772,N_2718);
nand U2847 (N_2847,N_2739,N_2728);
nand U2848 (N_2848,N_2743,N_2726);
or U2849 (N_2849,N_2729,N_2750);
nor U2850 (N_2850,N_2818,N_2800);
nor U2851 (N_2851,N_2806,N_2839);
and U2852 (N_2852,N_2777,N_2799);
nand U2853 (N_2853,N_2819,N_2816);
and U2854 (N_2854,N_2785,N_2823);
and U2855 (N_2855,N_2848,N_2822);
or U2856 (N_2856,N_2807,N_2824);
or U2857 (N_2857,N_2805,N_2847);
and U2858 (N_2858,N_2843,N_2815);
nor U2859 (N_2859,N_2828,N_2825);
nor U2860 (N_2860,N_2817,N_2846);
or U2861 (N_2861,N_2827,N_2793);
nand U2862 (N_2862,N_2830,N_2836);
or U2863 (N_2863,N_2781,N_2832);
xnor U2864 (N_2864,N_2776,N_2842);
or U2865 (N_2865,N_2787,N_2831);
nor U2866 (N_2866,N_2789,N_2795);
xnor U2867 (N_2867,N_2797,N_2821);
and U2868 (N_2868,N_2838,N_2790);
or U2869 (N_2869,N_2784,N_2810);
nor U2870 (N_2870,N_2798,N_2845);
nor U2871 (N_2871,N_2791,N_2794);
nor U2872 (N_2872,N_2812,N_2820);
nand U2873 (N_2873,N_2786,N_2803);
or U2874 (N_2874,N_2809,N_2796);
nand U2875 (N_2875,N_2782,N_2829);
and U2876 (N_2876,N_2844,N_2833);
or U2877 (N_2877,N_2840,N_2849);
nor U2878 (N_2878,N_2835,N_2808);
nor U2879 (N_2879,N_2783,N_2826);
or U2880 (N_2880,N_2780,N_2801);
nor U2881 (N_2881,N_2788,N_2837);
nor U2882 (N_2882,N_2778,N_2841);
or U2883 (N_2883,N_2792,N_2814);
nand U2884 (N_2884,N_2779,N_2804);
or U2885 (N_2885,N_2834,N_2813);
nor U2886 (N_2886,N_2775,N_2811);
nand U2887 (N_2887,N_2802,N_2808);
or U2888 (N_2888,N_2811,N_2836);
or U2889 (N_2889,N_2781,N_2836);
and U2890 (N_2890,N_2806,N_2821);
and U2891 (N_2891,N_2823,N_2816);
or U2892 (N_2892,N_2845,N_2812);
nand U2893 (N_2893,N_2842,N_2839);
nor U2894 (N_2894,N_2814,N_2845);
nand U2895 (N_2895,N_2838,N_2822);
or U2896 (N_2896,N_2847,N_2813);
nor U2897 (N_2897,N_2811,N_2796);
nand U2898 (N_2898,N_2812,N_2786);
or U2899 (N_2899,N_2842,N_2779);
xor U2900 (N_2900,N_2803,N_2794);
and U2901 (N_2901,N_2823,N_2814);
or U2902 (N_2902,N_2787,N_2812);
nand U2903 (N_2903,N_2818,N_2815);
or U2904 (N_2904,N_2797,N_2794);
and U2905 (N_2905,N_2775,N_2802);
or U2906 (N_2906,N_2792,N_2830);
nand U2907 (N_2907,N_2783,N_2818);
and U2908 (N_2908,N_2792,N_2835);
and U2909 (N_2909,N_2844,N_2823);
or U2910 (N_2910,N_2827,N_2807);
nand U2911 (N_2911,N_2839,N_2812);
nand U2912 (N_2912,N_2833,N_2822);
nor U2913 (N_2913,N_2806,N_2833);
nor U2914 (N_2914,N_2786,N_2809);
or U2915 (N_2915,N_2804,N_2839);
nor U2916 (N_2916,N_2781,N_2783);
nor U2917 (N_2917,N_2786,N_2807);
nand U2918 (N_2918,N_2781,N_2844);
nand U2919 (N_2919,N_2803,N_2846);
or U2920 (N_2920,N_2782,N_2826);
and U2921 (N_2921,N_2808,N_2843);
nand U2922 (N_2922,N_2779,N_2824);
nor U2923 (N_2923,N_2781,N_2777);
or U2924 (N_2924,N_2842,N_2781);
or U2925 (N_2925,N_2892,N_2909);
and U2926 (N_2926,N_2883,N_2866);
nand U2927 (N_2927,N_2901,N_2904);
and U2928 (N_2928,N_2911,N_2872);
and U2929 (N_2929,N_2868,N_2903);
or U2930 (N_2930,N_2888,N_2918);
nor U2931 (N_2931,N_2863,N_2862);
nor U2932 (N_2932,N_2922,N_2907);
and U2933 (N_2933,N_2882,N_2915);
nand U2934 (N_2934,N_2890,N_2908);
nand U2935 (N_2935,N_2870,N_2884);
and U2936 (N_2936,N_2891,N_2864);
nor U2937 (N_2937,N_2865,N_2858);
or U2938 (N_2938,N_2920,N_2854);
or U2939 (N_2939,N_2924,N_2889);
nand U2940 (N_2940,N_2902,N_2861);
and U2941 (N_2941,N_2855,N_2857);
nand U2942 (N_2942,N_2887,N_2885);
or U2943 (N_2943,N_2921,N_2874);
nand U2944 (N_2944,N_2894,N_2856);
and U2945 (N_2945,N_2871,N_2913);
nor U2946 (N_2946,N_2897,N_2880);
and U2947 (N_2947,N_2879,N_2916);
nor U2948 (N_2948,N_2886,N_2869);
and U2949 (N_2949,N_2859,N_2910);
and U2950 (N_2950,N_2873,N_2906);
nand U2951 (N_2951,N_2895,N_2919);
nand U2952 (N_2952,N_2900,N_2852);
and U2953 (N_2953,N_2893,N_2860);
nand U2954 (N_2954,N_2850,N_2905);
nand U2955 (N_2955,N_2914,N_2851);
nor U2956 (N_2956,N_2896,N_2917);
xnor U2957 (N_2957,N_2899,N_2875);
or U2958 (N_2958,N_2878,N_2912);
nor U2959 (N_2959,N_2876,N_2881);
nand U2960 (N_2960,N_2898,N_2853);
or U2961 (N_2961,N_2923,N_2877);
nand U2962 (N_2962,N_2867,N_2915);
or U2963 (N_2963,N_2878,N_2922);
nor U2964 (N_2964,N_2902,N_2882);
nand U2965 (N_2965,N_2916,N_2891);
nand U2966 (N_2966,N_2874,N_2884);
and U2967 (N_2967,N_2868,N_2859);
nor U2968 (N_2968,N_2883,N_2916);
or U2969 (N_2969,N_2868,N_2882);
nand U2970 (N_2970,N_2881,N_2889);
and U2971 (N_2971,N_2922,N_2900);
nand U2972 (N_2972,N_2910,N_2860);
and U2973 (N_2973,N_2865,N_2898);
and U2974 (N_2974,N_2863,N_2899);
nand U2975 (N_2975,N_2908,N_2861);
nor U2976 (N_2976,N_2856,N_2887);
and U2977 (N_2977,N_2858,N_2892);
and U2978 (N_2978,N_2902,N_2913);
nor U2979 (N_2979,N_2866,N_2860);
nor U2980 (N_2980,N_2864,N_2882);
and U2981 (N_2981,N_2862,N_2912);
or U2982 (N_2982,N_2912,N_2867);
or U2983 (N_2983,N_2896,N_2923);
and U2984 (N_2984,N_2902,N_2885);
nand U2985 (N_2985,N_2868,N_2904);
nor U2986 (N_2986,N_2867,N_2880);
and U2987 (N_2987,N_2852,N_2893);
nand U2988 (N_2988,N_2886,N_2904);
and U2989 (N_2989,N_2917,N_2894);
xnor U2990 (N_2990,N_2923,N_2887);
and U2991 (N_2991,N_2862,N_2874);
nor U2992 (N_2992,N_2883,N_2872);
nor U2993 (N_2993,N_2858,N_2884);
and U2994 (N_2994,N_2894,N_2879);
or U2995 (N_2995,N_2868,N_2855);
or U2996 (N_2996,N_2904,N_2919);
or U2997 (N_2997,N_2913,N_2919);
nand U2998 (N_2998,N_2915,N_2894);
nand U2999 (N_2999,N_2905,N_2877);
or UO_0 (O_0,N_2952,N_2980);
and UO_1 (O_1,N_2964,N_2936);
nor UO_2 (O_2,N_2973,N_2928);
nor UO_3 (O_3,N_2946,N_2983);
nand UO_4 (O_4,N_2996,N_2959);
or UO_5 (O_5,N_2966,N_2997);
and UO_6 (O_6,N_2944,N_2970);
nand UO_7 (O_7,N_2942,N_2950);
nor UO_8 (O_8,N_2977,N_2953);
xor UO_9 (O_9,N_2963,N_2937);
nand UO_10 (O_10,N_2929,N_2969);
nor UO_11 (O_11,N_2926,N_2978);
nor UO_12 (O_12,N_2954,N_2976);
nand UO_13 (O_13,N_2994,N_2938);
nand UO_14 (O_14,N_2975,N_2930);
or UO_15 (O_15,N_2951,N_2956);
nand UO_16 (O_16,N_2987,N_2990);
or UO_17 (O_17,N_2925,N_2974);
or UO_18 (O_18,N_2968,N_2941);
nor UO_19 (O_19,N_2999,N_2947);
nand UO_20 (O_20,N_2949,N_2931);
and UO_21 (O_21,N_2939,N_2934);
nand UO_22 (O_22,N_2988,N_2927);
nand UO_23 (O_23,N_2960,N_2955);
nand UO_24 (O_24,N_2933,N_2957);
nand UO_25 (O_25,N_2961,N_2998);
and UO_26 (O_26,N_2981,N_2948);
nand UO_27 (O_27,N_2991,N_2993);
nand UO_28 (O_28,N_2985,N_2945);
and UO_29 (O_29,N_2958,N_2971);
or UO_30 (O_30,N_2979,N_2940);
or UO_31 (O_31,N_2995,N_2935);
and UO_32 (O_32,N_2986,N_2984);
nor UO_33 (O_33,N_2982,N_2992);
nand UO_34 (O_34,N_2932,N_2965);
nand UO_35 (O_35,N_2943,N_2962);
nor UO_36 (O_36,N_2967,N_2989);
or UO_37 (O_37,N_2972,N_2935);
nor UO_38 (O_38,N_2934,N_2943);
and UO_39 (O_39,N_2935,N_2984);
or UO_40 (O_40,N_2933,N_2976);
nor UO_41 (O_41,N_2943,N_2996);
nor UO_42 (O_42,N_2987,N_2998);
or UO_43 (O_43,N_2958,N_2955);
nand UO_44 (O_44,N_2976,N_2950);
or UO_45 (O_45,N_2925,N_2939);
nor UO_46 (O_46,N_2987,N_2992);
nor UO_47 (O_47,N_2950,N_2955);
and UO_48 (O_48,N_2955,N_2926);
or UO_49 (O_49,N_2944,N_2969);
nor UO_50 (O_50,N_2928,N_2970);
and UO_51 (O_51,N_2975,N_2997);
or UO_52 (O_52,N_2996,N_2958);
and UO_53 (O_53,N_2952,N_2968);
or UO_54 (O_54,N_2973,N_2961);
nand UO_55 (O_55,N_2999,N_2980);
or UO_56 (O_56,N_2991,N_2933);
and UO_57 (O_57,N_2985,N_2935);
nor UO_58 (O_58,N_2991,N_2929);
xnor UO_59 (O_59,N_2942,N_2946);
nand UO_60 (O_60,N_2962,N_2945);
and UO_61 (O_61,N_2952,N_2994);
or UO_62 (O_62,N_2975,N_2986);
nand UO_63 (O_63,N_2967,N_2937);
or UO_64 (O_64,N_2943,N_2950);
nand UO_65 (O_65,N_2975,N_2956);
nand UO_66 (O_66,N_2969,N_2948);
nor UO_67 (O_67,N_2986,N_2932);
and UO_68 (O_68,N_2989,N_2933);
nor UO_69 (O_69,N_2986,N_2998);
or UO_70 (O_70,N_2946,N_2987);
nor UO_71 (O_71,N_2995,N_2966);
nand UO_72 (O_72,N_2983,N_2949);
and UO_73 (O_73,N_2950,N_2969);
nand UO_74 (O_74,N_2989,N_2930);
nor UO_75 (O_75,N_2929,N_2987);
nand UO_76 (O_76,N_2964,N_2977);
nor UO_77 (O_77,N_2959,N_2951);
nor UO_78 (O_78,N_2940,N_2945);
nor UO_79 (O_79,N_2999,N_2961);
or UO_80 (O_80,N_2996,N_2949);
nor UO_81 (O_81,N_2961,N_2945);
nor UO_82 (O_82,N_2978,N_2973);
and UO_83 (O_83,N_2982,N_2960);
nand UO_84 (O_84,N_2938,N_2925);
and UO_85 (O_85,N_2988,N_2998);
and UO_86 (O_86,N_2952,N_2950);
nor UO_87 (O_87,N_2937,N_2972);
nand UO_88 (O_88,N_2992,N_2959);
and UO_89 (O_89,N_2952,N_2985);
and UO_90 (O_90,N_2968,N_2962);
nor UO_91 (O_91,N_2982,N_2966);
or UO_92 (O_92,N_2930,N_2940);
nand UO_93 (O_93,N_2991,N_2987);
or UO_94 (O_94,N_2954,N_2944);
or UO_95 (O_95,N_2975,N_2977);
or UO_96 (O_96,N_2961,N_2960);
nor UO_97 (O_97,N_2931,N_2998);
and UO_98 (O_98,N_2985,N_2966);
and UO_99 (O_99,N_2942,N_2975);
or UO_100 (O_100,N_2956,N_2930);
nand UO_101 (O_101,N_2941,N_2944);
and UO_102 (O_102,N_2962,N_2978);
and UO_103 (O_103,N_2965,N_2945);
nand UO_104 (O_104,N_2979,N_2960);
xnor UO_105 (O_105,N_2982,N_2976);
and UO_106 (O_106,N_2937,N_2981);
nor UO_107 (O_107,N_2932,N_2979);
nand UO_108 (O_108,N_2934,N_2979);
nor UO_109 (O_109,N_2951,N_2931);
nor UO_110 (O_110,N_2937,N_2926);
nor UO_111 (O_111,N_2934,N_2938);
or UO_112 (O_112,N_2939,N_2987);
and UO_113 (O_113,N_2946,N_2934);
and UO_114 (O_114,N_2981,N_2952);
nor UO_115 (O_115,N_2966,N_2974);
nand UO_116 (O_116,N_2984,N_2959);
nand UO_117 (O_117,N_2985,N_2980);
nor UO_118 (O_118,N_2951,N_2927);
nor UO_119 (O_119,N_2998,N_2951);
nand UO_120 (O_120,N_2981,N_2944);
nand UO_121 (O_121,N_2957,N_2968);
nor UO_122 (O_122,N_2933,N_2972);
nor UO_123 (O_123,N_2932,N_2937);
nor UO_124 (O_124,N_2961,N_2976);
nand UO_125 (O_125,N_2988,N_2979);
and UO_126 (O_126,N_2963,N_2934);
and UO_127 (O_127,N_2960,N_2967);
nand UO_128 (O_128,N_2957,N_2982);
nor UO_129 (O_129,N_2997,N_2942);
or UO_130 (O_130,N_2982,N_2963);
and UO_131 (O_131,N_2989,N_2949);
and UO_132 (O_132,N_2941,N_2925);
nand UO_133 (O_133,N_2934,N_2961);
nor UO_134 (O_134,N_2968,N_2997);
nor UO_135 (O_135,N_2946,N_2937);
nor UO_136 (O_136,N_2955,N_2937);
and UO_137 (O_137,N_2974,N_2938);
nand UO_138 (O_138,N_2973,N_2996);
or UO_139 (O_139,N_2926,N_2935);
or UO_140 (O_140,N_2978,N_2986);
nor UO_141 (O_141,N_2989,N_2996);
nor UO_142 (O_142,N_2981,N_2961);
and UO_143 (O_143,N_2949,N_2954);
and UO_144 (O_144,N_2994,N_2968);
or UO_145 (O_145,N_2940,N_2927);
xnor UO_146 (O_146,N_2957,N_2997);
nor UO_147 (O_147,N_2930,N_2928);
nor UO_148 (O_148,N_2933,N_2959);
or UO_149 (O_149,N_2974,N_2967);
and UO_150 (O_150,N_2936,N_2993);
nand UO_151 (O_151,N_2996,N_2941);
and UO_152 (O_152,N_2928,N_2994);
and UO_153 (O_153,N_2982,N_2987);
and UO_154 (O_154,N_2952,N_2953);
and UO_155 (O_155,N_2928,N_2982);
or UO_156 (O_156,N_2951,N_2967);
nand UO_157 (O_157,N_2982,N_2946);
and UO_158 (O_158,N_2933,N_2946);
or UO_159 (O_159,N_2938,N_2927);
nor UO_160 (O_160,N_2929,N_2927);
nand UO_161 (O_161,N_2947,N_2989);
nand UO_162 (O_162,N_2929,N_2949);
nor UO_163 (O_163,N_2969,N_2934);
and UO_164 (O_164,N_2927,N_2970);
nor UO_165 (O_165,N_2986,N_2926);
nor UO_166 (O_166,N_2965,N_2993);
nor UO_167 (O_167,N_2975,N_2995);
or UO_168 (O_168,N_2932,N_2926);
nand UO_169 (O_169,N_2992,N_2957);
or UO_170 (O_170,N_2996,N_2952);
nor UO_171 (O_171,N_2952,N_2931);
nand UO_172 (O_172,N_2933,N_2963);
and UO_173 (O_173,N_2958,N_2925);
and UO_174 (O_174,N_2969,N_2985);
nand UO_175 (O_175,N_2967,N_2971);
nor UO_176 (O_176,N_2966,N_2935);
and UO_177 (O_177,N_2973,N_2987);
nor UO_178 (O_178,N_2996,N_2947);
xnor UO_179 (O_179,N_2981,N_2957);
and UO_180 (O_180,N_2934,N_2984);
and UO_181 (O_181,N_2931,N_2995);
nand UO_182 (O_182,N_2971,N_2943);
or UO_183 (O_183,N_2978,N_2951);
nand UO_184 (O_184,N_2953,N_2976);
and UO_185 (O_185,N_2935,N_2937);
nor UO_186 (O_186,N_2958,N_2951);
or UO_187 (O_187,N_2957,N_2935);
nor UO_188 (O_188,N_2956,N_2943);
nor UO_189 (O_189,N_2944,N_2987);
or UO_190 (O_190,N_2955,N_2941);
or UO_191 (O_191,N_2997,N_2987);
nor UO_192 (O_192,N_2950,N_2945);
or UO_193 (O_193,N_2970,N_2978);
and UO_194 (O_194,N_2944,N_2963);
nand UO_195 (O_195,N_2988,N_2941);
nand UO_196 (O_196,N_2988,N_2964);
and UO_197 (O_197,N_2979,N_2958);
nand UO_198 (O_198,N_2969,N_2995);
nand UO_199 (O_199,N_2998,N_2935);
xor UO_200 (O_200,N_2961,N_2970);
nand UO_201 (O_201,N_2982,N_2950);
nand UO_202 (O_202,N_2982,N_2956);
nor UO_203 (O_203,N_2991,N_2930);
or UO_204 (O_204,N_2948,N_2935);
or UO_205 (O_205,N_2974,N_2997);
or UO_206 (O_206,N_2984,N_2983);
xnor UO_207 (O_207,N_2993,N_2959);
nor UO_208 (O_208,N_2995,N_2939);
and UO_209 (O_209,N_2932,N_2972);
nor UO_210 (O_210,N_2947,N_2946);
nand UO_211 (O_211,N_2941,N_2978);
and UO_212 (O_212,N_2941,N_2967);
nor UO_213 (O_213,N_2933,N_2993);
or UO_214 (O_214,N_2969,N_2994);
nand UO_215 (O_215,N_2984,N_2982);
or UO_216 (O_216,N_2983,N_2959);
and UO_217 (O_217,N_2980,N_2941);
nand UO_218 (O_218,N_2953,N_2936);
or UO_219 (O_219,N_2940,N_2966);
and UO_220 (O_220,N_2963,N_2993);
or UO_221 (O_221,N_2971,N_2998);
nor UO_222 (O_222,N_2974,N_2981);
xnor UO_223 (O_223,N_2940,N_2983);
nor UO_224 (O_224,N_2970,N_2940);
nand UO_225 (O_225,N_2980,N_2930);
or UO_226 (O_226,N_2940,N_2972);
nor UO_227 (O_227,N_2988,N_2960);
nand UO_228 (O_228,N_2935,N_2974);
and UO_229 (O_229,N_2948,N_2980);
and UO_230 (O_230,N_2990,N_2951);
and UO_231 (O_231,N_2978,N_2952);
and UO_232 (O_232,N_2929,N_2953);
nor UO_233 (O_233,N_2950,N_2956);
or UO_234 (O_234,N_2934,N_2973);
and UO_235 (O_235,N_2934,N_2945);
nor UO_236 (O_236,N_2943,N_2952);
nand UO_237 (O_237,N_2993,N_2951);
or UO_238 (O_238,N_2976,N_2996);
nand UO_239 (O_239,N_2987,N_2925);
nor UO_240 (O_240,N_2932,N_2995);
nand UO_241 (O_241,N_2963,N_2979);
nor UO_242 (O_242,N_2994,N_2992);
nor UO_243 (O_243,N_2948,N_2931);
and UO_244 (O_244,N_2944,N_2953);
nor UO_245 (O_245,N_2960,N_2985);
and UO_246 (O_246,N_2994,N_2949);
and UO_247 (O_247,N_2946,N_2969);
or UO_248 (O_248,N_2954,N_2986);
nor UO_249 (O_249,N_2994,N_2926);
and UO_250 (O_250,N_2949,N_2962);
and UO_251 (O_251,N_2945,N_2956);
nand UO_252 (O_252,N_2984,N_2929);
nor UO_253 (O_253,N_2978,N_2960);
nand UO_254 (O_254,N_2963,N_2948);
and UO_255 (O_255,N_2972,N_2991);
and UO_256 (O_256,N_2927,N_2960);
and UO_257 (O_257,N_2925,N_2948);
xor UO_258 (O_258,N_2992,N_2989);
or UO_259 (O_259,N_2951,N_2965);
or UO_260 (O_260,N_2988,N_2929);
nand UO_261 (O_261,N_2973,N_2972);
or UO_262 (O_262,N_2994,N_2982);
nor UO_263 (O_263,N_2967,N_2950);
nor UO_264 (O_264,N_2997,N_2980);
nor UO_265 (O_265,N_2938,N_2955);
or UO_266 (O_266,N_2936,N_2975);
nor UO_267 (O_267,N_2933,N_2978);
nand UO_268 (O_268,N_2932,N_2934);
nand UO_269 (O_269,N_2928,N_2986);
or UO_270 (O_270,N_2965,N_2971);
nand UO_271 (O_271,N_2952,N_2955);
and UO_272 (O_272,N_2972,N_2954);
or UO_273 (O_273,N_2988,N_2956);
nor UO_274 (O_274,N_2972,N_2998);
or UO_275 (O_275,N_2976,N_2967);
or UO_276 (O_276,N_2929,N_2942);
and UO_277 (O_277,N_2929,N_2928);
and UO_278 (O_278,N_2951,N_2986);
nor UO_279 (O_279,N_2952,N_2945);
and UO_280 (O_280,N_2966,N_2946);
nor UO_281 (O_281,N_2968,N_2967);
and UO_282 (O_282,N_2947,N_2925);
or UO_283 (O_283,N_2956,N_2949);
or UO_284 (O_284,N_2961,N_2946);
and UO_285 (O_285,N_2980,N_2962);
nand UO_286 (O_286,N_2949,N_2977);
or UO_287 (O_287,N_2948,N_2975);
or UO_288 (O_288,N_2932,N_2991);
nand UO_289 (O_289,N_2944,N_2984);
or UO_290 (O_290,N_2962,N_2957);
nand UO_291 (O_291,N_2962,N_2938);
and UO_292 (O_292,N_2978,N_2964);
and UO_293 (O_293,N_2982,N_2967);
nand UO_294 (O_294,N_2993,N_2942);
or UO_295 (O_295,N_2934,N_2935);
or UO_296 (O_296,N_2957,N_2937);
nand UO_297 (O_297,N_2943,N_2984);
and UO_298 (O_298,N_2951,N_2972);
and UO_299 (O_299,N_2958,N_2987);
nor UO_300 (O_300,N_2952,N_2983);
nor UO_301 (O_301,N_2979,N_2989);
and UO_302 (O_302,N_2976,N_2965);
or UO_303 (O_303,N_2992,N_2996);
or UO_304 (O_304,N_2953,N_2978);
or UO_305 (O_305,N_2985,N_2965);
nand UO_306 (O_306,N_2975,N_2929);
or UO_307 (O_307,N_2991,N_2990);
nor UO_308 (O_308,N_2944,N_2996);
and UO_309 (O_309,N_2933,N_2958);
or UO_310 (O_310,N_2997,N_2960);
nor UO_311 (O_311,N_2961,N_2966);
nor UO_312 (O_312,N_2931,N_2992);
and UO_313 (O_313,N_2976,N_2934);
nand UO_314 (O_314,N_2939,N_2950);
nand UO_315 (O_315,N_2983,N_2939);
or UO_316 (O_316,N_2976,N_2948);
nor UO_317 (O_317,N_2970,N_2967);
nand UO_318 (O_318,N_2977,N_2938);
and UO_319 (O_319,N_2938,N_2971);
nor UO_320 (O_320,N_2942,N_2947);
nor UO_321 (O_321,N_2972,N_2997);
nor UO_322 (O_322,N_2934,N_2960);
and UO_323 (O_323,N_2951,N_2948);
nor UO_324 (O_324,N_2956,N_2932);
and UO_325 (O_325,N_2968,N_2990);
or UO_326 (O_326,N_2994,N_2964);
nand UO_327 (O_327,N_2970,N_2986);
and UO_328 (O_328,N_2975,N_2952);
and UO_329 (O_329,N_2993,N_2989);
and UO_330 (O_330,N_2987,N_2930);
nor UO_331 (O_331,N_2977,N_2929);
and UO_332 (O_332,N_2954,N_2942);
or UO_333 (O_333,N_2960,N_2986);
and UO_334 (O_334,N_2985,N_2928);
or UO_335 (O_335,N_2963,N_2936);
or UO_336 (O_336,N_2987,N_2931);
and UO_337 (O_337,N_2959,N_2953);
or UO_338 (O_338,N_2995,N_2973);
and UO_339 (O_339,N_2955,N_2972);
nand UO_340 (O_340,N_2956,N_2977);
or UO_341 (O_341,N_2938,N_2988);
nand UO_342 (O_342,N_2965,N_2930);
and UO_343 (O_343,N_2930,N_2958);
nand UO_344 (O_344,N_2954,N_2997);
nor UO_345 (O_345,N_2992,N_2999);
nor UO_346 (O_346,N_2945,N_2993);
or UO_347 (O_347,N_2989,N_2965);
xor UO_348 (O_348,N_2968,N_2975);
or UO_349 (O_349,N_2951,N_2994);
or UO_350 (O_350,N_2953,N_2987);
nand UO_351 (O_351,N_2958,N_2929);
xor UO_352 (O_352,N_2929,N_2947);
and UO_353 (O_353,N_2978,N_2948);
or UO_354 (O_354,N_2925,N_2990);
and UO_355 (O_355,N_2939,N_2929);
or UO_356 (O_356,N_2954,N_2940);
and UO_357 (O_357,N_2954,N_2991);
or UO_358 (O_358,N_2941,N_2952);
or UO_359 (O_359,N_2965,N_2939);
nor UO_360 (O_360,N_2981,N_2942);
or UO_361 (O_361,N_2934,N_2957);
nor UO_362 (O_362,N_2982,N_2972);
or UO_363 (O_363,N_2944,N_2932);
and UO_364 (O_364,N_2982,N_2986);
nand UO_365 (O_365,N_2990,N_2972);
or UO_366 (O_366,N_2925,N_2973);
nand UO_367 (O_367,N_2966,N_2970);
nor UO_368 (O_368,N_2940,N_2944);
or UO_369 (O_369,N_2983,N_2977);
or UO_370 (O_370,N_2927,N_2995);
or UO_371 (O_371,N_2936,N_2992);
nand UO_372 (O_372,N_2983,N_2967);
nand UO_373 (O_373,N_2961,N_2991);
nand UO_374 (O_374,N_2929,N_2935);
nor UO_375 (O_375,N_2985,N_2970);
or UO_376 (O_376,N_2932,N_2951);
or UO_377 (O_377,N_2931,N_2958);
nand UO_378 (O_378,N_2936,N_2997);
nor UO_379 (O_379,N_2991,N_2937);
nand UO_380 (O_380,N_2959,N_2935);
nor UO_381 (O_381,N_2952,N_2928);
or UO_382 (O_382,N_2947,N_2964);
or UO_383 (O_383,N_2953,N_2943);
xor UO_384 (O_384,N_2960,N_2928);
nor UO_385 (O_385,N_2988,N_2931);
nand UO_386 (O_386,N_2961,N_2969);
or UO_387 (O_387,N_2930,N_2997);
and UO_388 (O_388,N_2980,N_2933);
and UO_389 (O_389,N_2935,N_2983);
and UO_390 (O_390,N_2958,N_2967);
or UO_391 (O_391,N_2964,N_2998);
nor UO_392 (O_392,N_2985,N_2944);
nor UO_393 (O_393,N_2933,N_2961);
and UO_394 (O_394,N_2985,N_2973);
nor UO_395 (O_395,N_2940,N_2958);
nor UO_396 (O_396,N_2939,N_2959);
or UO_397 (O_397,N_2994,N_2931);
and UO_398 (O_398,N_2981,N_2995);
nor UO_399 (O_399,N_2929,N_2998);
nand UO_400 (O_400,N_2986,N_2955);
nor UO_401 (O_401,N_2955,N_2939);
nor UO_402 (O_402,N_2974,N_2948);
and UO_403 (O_403,N_2982,N_2947);
and UO_404 (O_404,N_2942,N_2988);
nor UO_405 (O_405,N_2938,N_2933);
and UO_406 (O_406,N_2938,N_2940);
nor UO_407 (O_407,N_2974,N_2941);
nor UO_408 (O_408,N_2931,N_2925);
xor UO_409 (O_409,N_2944,N_2948);
and UO_410 (O_410,N_2969,N_2938);
and UO_411 (O_411,N_2950,N_2959);
nand UO_412 (O_412,N_2956,N_2962);
or UO_413 (O_413,N_2995,N_2930);
nand UO_414 (O_414,N_2975,N_2928);
nor UO_415 (O_415,N_2945,N_2957);
xor UO_416 (O_416,N_2980,N_2939);
nand UO_417 (O_417,N_2970,N_2991);
nand UO_418 (O_418,N_2984,N_2997);
nand UO_419 (O_419,N_2991,N_2948);
nor UO_420 (O_420,N_2997,N_2940);
or UO_421 (O_421,N_2929,N_2931);
and UO_422 (O_422,N_2942,N_2971);
nand UO_423 (O_423,N_2962,N_2979);
nand UO_424 (O_424,N_2930,N_2968);
nand UO_425 (O_425,N_2964,N_2958);
and UO_426 (O_426,N_2982,N_2925);
nor UO_427 (O_427,N_2981,N_2986);
nand UO_428 (O_428,N_2961,N_2931);
nand UO_429 (O_429,N_2985,N_2971);
and UO_430 (O_430,N_2983,N_2964);
nand UO_431 (O_431,N_2977,N_2943);
nor UO_432 (O_432,N_2978,N_2931);
or UO_433 (O_433,N_2934,N_2931);
or UO_434 (O_434,N_2972,N_2969);
and UO_435 (O_435,N_2977,N_2981);
nor UO_436 (O_436,N_2948,N_2954);
and UO_437 (O_437,N_2994,N_2988);
nor UO_438 (O_438,N_2961,N_2971);
nor UO_439 (O_439,N_2977,N_2934);
nor UO_440 (O_440,N_2982,N_2958);
nand UO_441 (O_441,N_2968,N_2939);
or UO_442 (O_442,N_2989,N_2994);
and UO_443 (O_443,N_2987,N_2970);
and UO_444 (O_444,N_2936,N_2987);
or UO_445 (O_445,N_2969,N_2953);
nand UO_446 (O_446,N_2970,N_2988);
and UO_447 (O_447,N_2934,N_2951);
nand UO_448 (O_448,N_2968,N_2995);
nand UO_449 (O_449,N_2966,N_2960);
nor UO_450 (O_450,N_2928,N_2948);
nor UO_451 (O_451,N_2992,N_2926);
and UO_452 (O_452,N_2969,N_2951);
nor UO_453 (O_453,N_2993,N_2928);
and UO_454 (O_454,N_2997,N_2969);
nor UO_455 (O_455,N_2941,N_2985);
and UO_456 (O_456,N_2932,N_2975);
and UO_457 (O_457,N_2999,N_2967);
and UO_458 (O_458,N_2942,N_2952);
nand UO_459 (O_459,N_2993,N_2925);
or UO_460 (O_460,N_2933,N_2943);
and UO_461 (O_461,N_2968,N_2942);
and UO_462 (O_462,N_2974,N_2937);
nand UO_463 (O_463,N_2926,N_2942);
nand UO_464 (O_464,N_2933,N_2997);
and UO_465 (O_465,N_2976,N_2986);
nor UO_466 (O_466,N_2998,N_2941);
xnor UO_467 (O_467,N_2976,N_2959);
and UO_468 (O_468,N_2963,N_2994);
and UO_469 (O_469,N_2970,N_2998);
nand UO_470 (O_470,N_2973,N_2999);
or UO_471 (O_471,N_2939,N_2932);
nand UO_472 (O_472,N_2955,N_2948);
xnor UO_473 (O_473,N_2955,N_2945);
nand UO_474 (O_474,N_2985,N_2933);
nand UO_475 (O_475,N_2991,N_2960);
nor UO_476 (O_476,N_2945,N_2967);
nor UO_477 (O_477,N_2942,N_2991);
nor UO_478 (O_478,N_2941,N_2987);
and UO_479 (O_479,N_2949,N_2950);
nor UO_480 (O_480,N_2985,N_2938);
or UO_481 (O_481,N_2985,N_2979);
and UO_482 (O_482,N_2955,N_2994);
nand UO_483 (O_483,N_2999,N_2988);
and UO_484 (O_484,N_2977,N_2927);
nor UO_485 (O_485,N_2946,N_2938);
xor UO_486 (O_486,N_2993,N_2985);
nand UO_487 (O_487,N_2927,N_2932);
nor UO_488 (O_488,N_2994,N_2986);
or UO_489 (O_489,N_2928,N_2996);
or UO_490 (O_490,N_2930,N_2979);
or UO_491 (O_491,N_2992,N_2939);
nand UO_492 (O_492,N_2966,N_2932);
nor UO_493 (O_493,N_2967,N_2963);
nand UO_494 (O_494,N_2993,N_2956);
and UO_495 (O_495,N_2975,N_2958);
nor UO_496 (O_496,N_2991,N_2957);
nand UO_497 (O_497,N_2956,N_2928);
or UO_498 (O_498,N_2951,N_2942);
nor UO_499 (O_499,N_2935,N_2939);
endmodule