module basic_750_5000_1000_2_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2504,N_2505,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2552,N_2553,N_2554,N_2555,N_2557,N_2558,N_2559,N_2561,N_2562,N_2564,N_2565,N_2566,N_2567,N_2568,N_2570,N_2571,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2591,N_2593,N_2594,N_2595,N_2596,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2616,N_2618,N_2621,N_2622,N_2623,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2653,N_2655,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2673,N_2674,N_2675,N_2677,N_2678,N_2679,N_2680,N_2682,N_2684,N_2688,N_2689,N_2690,N_2692,N_2695,N_2696,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2716,N_2718,N_2719,N_2721,N_2722,N_2726,N_2727,N_2728,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2747,N_2748,N_2749,N_2751,N_2752,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2770,N_2771,N_2772,N_2773,N_2774,N_2776,N_2777,N_2779,N_2780,N_2782,N_2783,N_2784,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2807,N_2808,N_2809,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2818,N_2819,N_2821,N_2822,N_2823,N_2824,N_2826,N_2827,N_2828,N_2830,N_2831,N_2832,N_2834,N_2837,N_2838,N_2839,N_2840,N_2841,N_2843,N_2844,N_2845,N_2846,N_2848,N_2849,N_2851,N_2852,N_2854,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2865,N_2866,N_2867,N_2868,N_2870,N_2873,N_2874,N_2876,N_2877,N_2878,N_2879,N_2880,N_2883,N_2884,N_2885,N_2887,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2945,N_2946,N_2947,N_2948,N_2949,N_2951,N_2952,N_2953,N_2954,N_2955,N_2957,N_2958,N_2959,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2977,N_2978,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2987,N_2989,N_2990,N_2991,N_2993,N_2994,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3003,N_3004,N_3005,N_3009,N_3010,N_3011,N_3012,N_3013,N_3017,N_3019,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3029,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3068,N_3070,N_3071,N_3075,N_3076,N_3078,N_3079,N_3080,N_3081,N_3082,N_3084,N_3085,N_3086,N_3088,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3098,N_3101,N_3103,N_3104,N_3105,N_3106,N_3107,N_3109,N_3111,N_3112,N_3114,N_3115,N_3116,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3138,N_3139,N_3140,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3151,N_3152,N_3153,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3185,N_3186,N_3187,N_3189,N_3190,N_3191,N_3194,N_3197,N_3199,N_3200,N_3201,N_3202,N_3203,N_3206,N_3207,N_3208,N_3209,N_3210,N_3212,N_3214,N_3216,N_3217,N_3218,N_3219,N_3220,N_3223,N_3224,N_3225,N_3227,N_3228,N_3229,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3241,N_3242,N_3243,N_3245,N_3246,N_3247,N_3248,N_3249,N_3251,N_3252,N_3253,N_3255,N_3257,N_3259,N_3260,N_3261,N_3263,N_3264,N_3265,N_3266,N_3267,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3284,N_3285,N_3286,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3300,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3311,N_3312,N_3313,N_3314,N_3317,N_3319,N_3320,N_3321,N_3322,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3359,N_3360,N_3361,N_3363,N_3364,N_3365,N_3366,N_3367,N_3369,N_3371,N_3373,N_3374,N_3375,N_3376,N_3377,N_3379,N_3381,N_3382,N_3383,N_3384,N_3385,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3398,N_3401,N_3403,N_3404,N_3405,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3416,N_3417,N_3418,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3440,N_3441,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3460,N_3461,N_3462,N_3463,N_3465,N_3466,N_3467,N_3471,N_3473,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3495,N_3496,N_3497,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3511,N_3513,N_3514,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3547,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3587,N_3588,N_3589,N_3590,N_3592,N_3593,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3607,N_3609,N_3610,N_3611,N_3612,N_3613,N_3615,N_3616,N_3617,N_3618,N_3619,N_3621,N_3623,N_3624,N_3627,N_3628,N_3629,N_3630,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3641,N_3642,N_3643,N_3644,N_3646,N_3648,N_3649,N_3653,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3672,N_3674,N_3675,N_3677,N_3679,N_3680,N_3681,N_3682,N_3684,N_3685,N_3686,N_3687,N_3690,N_3692,N_3693,N_3695,N_3696,N_3697,N_3698,N_3700,N_3702,N_3703,N_3704,N_3706,N_3707,N_3708,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3744,N_3746,N_3747,N_3748,N_3754,N_3756,N_3757,N_3758,N_3760,N_3761,N_3762,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3775,N_3776,N_3777,N_3778,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3789,N_3791,N_3792,N_3793,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3804,N_3805,N_3806,N_3807,N_3808,N_3810,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3828,N_3829,N_3830,N_3831,N_3832,N_3834,N_3835,N_3836,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3852,N_3854,N_3855,N_3856,N_3859,N_3860,N_3861,N_3862,N_3863,N_3865,N_3866,N_3867,N_3870,N_3871,N_3872,N_3873,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3882,N_3883,N_3884,N_3886,N_3887,N_3888,N_3889,N_3890,N_3892,N_3893,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3907,N_3908,N_3909,N_3913,N_3917,N_3918,N_3919,N_3920,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3932,N_3933,N_3935,N_3937,N_3939,N_3940,N_3941,N_3942,N_3943,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3954,N_3955,N_3956,N_3957,N_3958,N_3961,N_3962,N_3964,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3984,N_3985,N_3986,N_3987,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3996,N_3997,N_3998,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4018,N_4019,N_4021,N_4023,N_4025,N_4026,N_4027,N_4028,N_4030,N_4032,N_4033,N_4035,N_4036,N_4037,N_4038,N_4040,N_4041,N_4043,N_4044,N_4046,N_4048,N_4049,N_4050,N_4052,N_4053,N_4054,N_4055,N_4057,N_4058,N_4059,N_4061,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4083,N_4084,N_4085,N_4088,N_4089,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4100,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4113,N_4114,N_4116,N_4117,N_4118,N_4119,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4148,N_4149,N_4150,N_4151,N_4152,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4163,N_4164,N_4165,N_4167,N_4168,N_4169,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4191,N_4192,N_4194,N_4195,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4207,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4218,N_4219,N_4220,N_4222,N_4223,N_4224,N_4225,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4235,N_4237,N_4238,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4272,N_4273,N_4275,N_4276,N_4277,N_4278,N_4279,N_4282,N_4283,N_4284,N_4285,N_4286,N_4288,N_4289,N_4290,N_4291,N_4292,N_4295,N_4296,N_4297,N_4299,N_4301,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4319,N_4321,N_4322,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4337,N_4339,N_4340,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4369,N_4370,N_4371,N_4373,N_4374,N_4376,N_4377,N_4379,N_4380,N_4382,N_4383,N_4384,N_4385,N_4386,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4423,N_4424,N_4425,N_4427,N_4428,N_4429,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4466,N_4467,N_4468,N_4469,N_4470,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4521,N_4522,N_4523,N_4524,N_4525,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4541,N_4542,N_4543,N_4545,N_4546,N_4548,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4559,N_4561,N_4566,N_4567,N_4569,N_4570,N_4571,N_4572,N_4573,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4583,N_4584,N_4585,N_4589,N_4590,N_4592,N_4594,N_4595,N_4596,N_4597,N_4598,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4613,N_4614,N_4615,N_4616,N_4618,N_4619,N_4620,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4631,N_4632,N_4634,N_4635,N_4636,N_4637,N_4639,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4656,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4679,N_4681,N_4682,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4705,N_4706,N_4708,N_4709,N_4712,N_4713,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4742,N_4743,N_4745,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4755,N_4756,N_4757,N_4758,N_4759,N_4763,N_4764,N_4768,N_4770,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4829,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4840,N_4841,N_4842,N_4843,N_4845,N_4846,N_4847,N_4849,N_4851,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4869,N_4871,N_4872,N_4873,N_4874,N_4875,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4887,N_4888,N_4889,N_4890,N_4891,N_4894,N_4895,N_4896,N_4898,N_4900,N_4901,N_4902,N_4903,N_4904,N_4907,N_4908,N_4909,N_4911,N_4912,N_4913,N_4914,N_4915,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4946,N_4947,N_4948,N_4949,N_4950,N_4952,N_4953,N_4954,N_4955,N_4956,N_4958,N_4959,N_4960,N_4962,N_4963,N_4964,N_4966,N_4967,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4986,N_4988,N_4989,N_4991,N_4992,N_4993,N_4996,N_4999;
nand U0 (N_0,In_278,In_52);
or U1 (N_1,In_200,In_638);
nor U2 (N_2,In_169,In_241);
xnor U3 (N_3,In_458,In_701);
nand U4 (N_4,In_694,In_743);
nor U5 (N_5,In_575,In_56);
xor U6 (N_6,In_530,In_6);
or U7 (N_7,In_389,In_528);
nand U8 (N_8,In_565,In_550);
and U9 (N_9,In_246,In_218);
nand U10 (N_10,In_716,In_454);
nand U11 (N_11,In_370,In_196);
nor U12 (N_12,In_579,In_117);
or U13 (N_13,In_734,In_708);
nand U14 (N_14,In_372,In_234);
nand U15 (N_15,In_461,In_36);
nor U16 (N_16,In_340,In_676);
nand U17 (N_17,In_192,In_67);
and U18 (N_18,In_490,In_586);
nor U19 (N_19,In_651,In_189);
and U20 (N_20,In_713,In_705);
and U21 (N_21,In_96,In_308);
or U22 (N_22,In_236,In_548);
nand U23 (N_23,In_437,In_726);
nor U24 (N_24,In_210,In_466);
nand U25 (N_25,In_97,In_741);
nand U26 (N_26,In_347,In_478);
or U27 (N_27,In_686,In_628);
and U28 (N_28,In_401,In_589);
nand U29 (N_29,In_43,In_13);
or U30 (N_30,In_300,In_604);
and U31 (N_31,In_105,In_2);
and U32 (N_32,In_733,In_400);
nor U33 (N_33,In_615,In_76);
nand U34 (N_34,In_568,In_115);
and U35 (N_35,In_298,In_260);
nand U36 (N_36,In_573,In_744);
nor U37 (N_37,In_470,In_516);
and U38 (N_38,In_309,In_227);
or U39 (N_39,In_731,In_109);
or U40 (N_40,In_46,In_337);
nor U41 (N_41,In_381,In_620);
xnor U42 (N_42,In_165,In_358);
nor U43 (N_43,In_555,In_139);
nor U44 (N_44,In_406,In_39);
and U45 (N_45,In_584,In_313);
or U46 (N_46,In_275,In_271);
nor U47 (N_47,In_197,In_63);
or U48 (N_48,In_679,In_459);
nand U49 (N_49,In_344,In_425);
and U50 (N_50,In_545,In_322);
nand U51 (N_51,In_511,In_75);
nor U52 (N_52,In_678,In_525);
or U53 (N_53,In_420,In_728);
nand U54 (N_54,In_131,In_449);
or U55 (N_55,In_26,In_147);
and U56 (N_56,In_282,In_623);
nor U57 (N_57,In_710,In_352);
nor U58 (N_58,In_50,In_605);
or U59 (N_59,In_320,In_281);
nor U60 (N_60,In_630,In_92);
nand U61 (N_61,In_94,In_262);
nor U62 (N_62,In_132,In_637);
nand U63 (N_63,In_42,In_252);
and U64 (N_64,In_356,In_700);
nor U65 (N_65,In_225,In_29);
nand U66 (N_66,In_680,In_738);
or U67 (N_67,In_727,In_622);
and U68 (N_68,In_664,In_178);
nand U69 (N_69,In_89,In_632);
nor U70 (N_70,In_500,In_624);
nor U71 (N_71,In_243,In_314);
nand U72 (N_72,In_464,In_532);
nand U73 (N_73,In_317,In_672);
or U74 (N_74,In_606,In_283);
nand U75 (N_75,In_539,In_148);
nor U76 (N_76,In_704,In_412);
nand U77 (N_77,In_190,In_287);
or U78 (N_78,In_621,In_489);
or U79 (N_79,In_167,In_455);
nor U80 (N_80,In_219,In_725);
nor U81 (N_81,In_659,In_581);
nor U82 (N_82,In_611,In_11);
nand U83 (N_83,In_506,In_533);
or U84 (N_84,In_657,In_480);
or U85 (N_85,In_41,In_587);
nand U86 (N_86,In_557,In_614);
or U87 (N_87,In_285,In_286);
nand U88 (N_88,In_502,In_327);
nand U89 (N_89,In_334,In_576);
or U90 (N_90,In_158,In_336);
nand U91 (N_91,In_343,In_712);
nor U92 (N_92,In_631,In_86);
and U93 (N_93,In_421,In_510);
nor U94 (N_94,In_215,In_114);
nand U95 (N_95,In_193,In_325);
and U96 (N_96,In_452,In_536);
and U97 (N_97,In_492,In_173);
nand U98 (N_98,In_121,In_475);
or U99 (N_99,In_16,In_293);
nor U100 (N_100,In_27,In_209);
and U101 (N_101,In_143,In_18);
or U102 (N_102,In_479,In_463);
or U103 (N_103,In_693,In_681);
and U104 (N_104,In_140,In_745);
or U105 (N_105,In_491,In_164);
or U106 (N_106,In_261,In_88);
and U107 (N_107,In_485,In_721);
or U108 (N_108,In_265,In_328);
and U109 (N_109,In_64,In_494);
and U110 (N_110,In_608,In_682);
or U111 (N_111,In_438,In_134);
nand U112 (N_112,In_656,In_229);
nor U113 (N_113,In_626,In_501);
or U114 (N_114,In_467,In_645);
nor U115 (N_115,In_527,In_155);
and U116 (N_116,In_288,In_504);
or U117 (N_117,In_17,In_351);
and U118 (N_118,In_570,In_345);
and U119 (N_119,In_577,In_719);
and U120 (N_120,In_411,In_652);
nor U121 (N_121,In_222,In_216);
nor U122 (N_122,In_7,In_152);
or U123 (N_123,In_49,In_208);
nor U124 (N_124,In_71,In_112);
or U125 (N_125,In_8,In_714);
nand U126 (N_126,In_474,In_161);
and U127 (N_127,In_667,In_204);
nand U128 (N_128,In_85,In_302);
or U129 (N_129,In_537,In_684);
and U130 (N_130,In_20,In_87);
or U131 (N_131,In_590,In_177);
nor U132 (N_132,In_446,In_562);
nand U133 (N_133,In_543,In_15);
nand U134 (N_134,In_303,In_199);
nor U135 (N_135,In_670,In_19);
nor U136 (N_136,In_166,In_440);
nor U137 (N_137,In_141,In_366);
nor U138 (N_138,In_697,In_129);
and U139 (N_139,In_277,In_360);
nor U140 (N_140,In_609,In_619);
and U141 (N_141,In_448,In_498);
nor U142 (N_142,In_72,In_299);
or U143 (N_143,In_397,In_186);
or U144 (N_144,In_28,In_331);
nor U145 (N_145,In_297,In_593);
nand U146 (N_146,In_578,In_654);
and U147 (N_147,In_332,In_258);
and U148 (N_148,In_142,In_385);
nand U149 (N_149,In_206,In_171);
nor U150 (N_150,In_558,In_183);
nand U151 (N_151,In_487,In_24);
or U152 (N_152,In_301,In_698);
nor U153 (N_153,In_130,In_191);
and U154 (N_154,In_696,In_40);
nand U155 (N_155,In_124,In_290);
or U156 (N_156,In_378,In_635);
nor U157 (N_157,In_321,In_515);
nand U158 (N_158,In_53,In_413);
nor U159 (N_159,In_482,In_172);
and U160 (N_160,In_217,In_595);
and U161 (N_161,In_429,In_497);
nand U162 (N_162,In_47,In_692);
and U163 (N_163,In_503,In_245);
or U164 (N_164,In_460,In_364);
nand U165 (N_165,In_445,In_5);
nor U166 (N_166,In_666,In_108);
nor U167 (N_167,In_407,In_405);
or U168 (N_168,In_214,In_116);
or U169 (N_169,In_711,In_444);
or U170 (N_170,In_57,In_368);
and U171 (N_171,In_122,In_599);
nand U172 (N_172,In_235,In_507);
nor U173 (N_173,In_333,In_508);
and U174 (N_174,In_136,In_184);
and U175 (N_175,In_230,In_125);
nor U176 (N_176,In_371,In_82);
nor U177 (N_177,In_12,In_594);
or U178 (N_178,In_648,In_379);
xnor U179 (N_179,In_735,In_365);
and U180 (N_180,In_1,In_556);
nor U181 (N_181,In_231,In_729);
nor U182 (N_182,In_38,In_382);
and U183 (N_183,In_484,In_384);
or U184 (N_184,In_205,In_30);
or U185 (N_185,In_468,In_644);
or U186 (N_186,In_483,In_677);
or U187 (N_187,In_709,In_153);
nor U188 (N_188,In_529,In_629);
nor U189 (N_189,In_362,In_95);
nor U190 (N_190,In_395,In_391);
or U191 (N_191,In_585,In_566);
and U192 (N_192,In_549,In_119);
nand U193 (N_193,In_553,In_603);
nor U194 (N_194,In_22,In_341);
nor U195 (N_195,In_607,In_251);
and U196 (N_196,In_10,In_403);
or U197 (N_197,In_23,In_514);
or U198 (N_198,In_610,In_394);
nor U199 (N_199,In_408,In_274);
nand U200 (N_200,In_737,In_432);
and U201 (N_201,In_418,In_633);
and U202 (N_202,In_58,In_509);
nand U203 (N_203,In_361,In_613);
nor U204 (N_204,In_32,In_228);
nand U205 (N_205,In_272,In_718);
and U206 (N_206,In_393,In_383);
and U207 (N_207,In_357,In_242);
and U208 (N_208,In_339,In_685);
or U209 (N_209,In_748,In_653);
or U210 (N_210,In_106,In_588);
nand U211 (N_211,In_640,In_98);
and U212 (N_212,In_239,In_233);
nor U213 (N_213,In_427,In_390);
nor U214 (N_214,In_538,In_226);
or U215 (N_215,In_146,In_447);
and U216 (N_216,In_306,In_127);
or U217 (N_217,In_133,In_583);
nor U218 (N_218,In_722,In_240);
and U219 (N_219,In_723,In_304);
and U220 (N_220,In_699,In_33);
and U221 (N_221,In_673,In_62);
nand U222 (N_222,In_668,In_329);
nor U223 (N_223,In_582,In_195);
or U224 (N_224,In_359,In_707);
and U225 (N_225,In_675,In_31);
and U226 (N_226,In_0,In_469);
nor U227 (N_227,In_574,In_691);
nor U228 (N_228,In_443,In_663);
and U229 (N_229,In_292,In_59);
nand U230 (N_230,In_221,In_749);
nor U231 (N_231,In_149,In_316);
or U232 (N_232,In_601,In_662);
and U233 (N_233,In_561,In_102);
or U234 (N_234,In_353,In_103);
or U235 (N_235,In_179,In_441);
nor U236 (N_236,In_717,In_456);
and U237 (N_237,In_83,In_695);
and U238 (N_238,In_355,In_690);
nor U239 (N_239,In_477,In_706);
nand U240 (N_240,In_254,In_380);
and U241 (N_241,In_616,In_720);
nand U242 (N_242,In_263,In_79);
and U243 (N_243,In_688,In_296);
nor U244 (N_244,In_66,In_202);
and U245 (N_245,In_513,In_182);
nor U246 (N_246,In_736,In_415);
nor U247 (N_247,In_433,In_517);
or U248 (N_248,In_289,In_111);
or U249 (N_249,In_534,In_37);
nor U250 (N_250,In_521,In_118);
nand U251 (N_251,In_213,In_671);
nand U252 (N_252,In_247,In_255);
and U253 (N_253,In_212,In_476);
and U254 (N_254,In_732,In_157);
nor U255 (N_255,In_658,In_571);
and U256 (N_256,In_646,In_373);
nor U257 (N_257,In_250,In_104);
or U258 (N_258,In_416,In_665);
and U259 (N_259,In_74,In_244);
nor U260 (N_260,In_617,In_311);
and U261 (N_261,In_392,In_3);
nor U262 (N_262,In_518,In_669);
nor U263 (N_263,In_291,In_546);
and U264 (N_264,In_367,In_175);
nand U265 (N_265,In_560,In_715);
nor U266 (N_266,In_439,In_404);
nor U267 (N_267,In_377,In_423);
or U268 (N_268,In_35,In_151);
nor U269 (N_269,In_375,In_598);
and U270 (N_270,In_535,In_551);
nor U271 (N_271,In_279,In_48);
or U272 (N_272,In_541,In_564);
or U273 (N_273,In_326,In_481);
nand U274 (N_274,In_627,In_493);
and U275 (N_275,In_55,In_524);
and U276 (N_276,In_323,In_597);
xnor U277 (N_277,In_386,In_702);
xor U278 (N_278,In_91,In_376);
or U279 (N_279,In_324,In_642);
or U280 (N_280,In_128,In_315);
or U281 (N_281,In_268,In_451);
or U282 (N_282,In_232,In_519);
or U283 (N_283,In_442,In_544);
or U284 (N_284,In_264,In_248);
nand U285 (N_285,In_180,In_267);
or U286 (N_286,In_526,In_223);
and U287 (N_287,In_295,In_428);
nand U288 (N_288,In_73,In_65);
nor U289 (N_289,In_68,In_211);
nand U290 (N_290,In_661,In_409);
nor U291 (N_291,In_572,In_655);
or U292 (N_292,In_249,In_496);
nor U293 (N_293,In_144,In_256);
nand U294 (N_294,In_338,In_54);
nor U295 (N_295,In_69,In_137);
and U296 (N_296,In_531,In_387);
or U297 (N_297,In_307,In_703);
and U298 (N_298,In_457,In_194);
or U299 (N_299,In_660,In_101);
or U300 (N_300,In_330,In_253);
nand U301 (N_301,In_554,In_224);
nor U302 (N_302,In_625,In_634);
nand U303 (N_303,In_374,In_540);
nand U304 (N_304,In_99,In_145);
nand U305 (N_305,In_643,In_45);
nor U306 (N_306,In_419,In_563);
nor U307 (N_307,In_399,In_520);
and U308 (N_308,In_542,In_284);
nand U309 (N_309,In_276,In_350);
and U310 (N_310,In_110,In_237);
nand U311 (N_311,In_649,In_417);
and U312 (N_312,In_348,In_473);
or U313 (N_313,In_472,In_505);
nand U314 (N_314,In_126,In_77);
and U315 (N_315,In_569,In_60);
and U316 (N_316,In_93,In_294);
nor U317 (N_317,In_414,In_641);
nand U318 (N_318,In_107,In_522);
nand U319 (N_319,In_159,In_14);
nand U320 (N_320,In_259,In_591);
and U321 (N_321,In_689,In_747);
or U322 (N_322,In_739,In_740);
nand U323 (N_323,In_523,In_154);
or U324 (N_324,In_176,In_185);
and U325 (N_325,In_170,In_305);
and U326 (N_326,In_51,In_201);
or U327 (N_327,In_430,In_270);
nor U328 (N_328,In_388,In_410);
nand U329 (N_329,In_471,In_552);
and U330 (N_330,In_160,In_465);
or U331 (N_331,In_4,In_547);
or U332 (N_332,In_369,In_319);
nor U333 (N_333,In_612,In_312);
xnor U334 (N_334,In_724,In_495);
or U335 (N_335,In_349,In_600);
and U336 (N_336,In_402,In_318);
or U337 (N_337,In_434,In_163);
nand U338 (N_338,In_120,In_450);
nand U339 (N_339,In_435,In_257);
nand U340 (N_340,In_592,In_462);
nand U341 (N_341,In_44,In_310);
nand U342 (N_342,In_138,In_687);
and U343 (N_343,In_78,In_266);
and U344 (N_344,In_61,In_123);
nand U345 (N_345,In_363,In_34);
and U346 (N_346,In_84,In_90);
xor U347 (N_347,In_207,In_280);
xnor U348 (N_348,In_436,In_512);
nor U349 (N_349,In_168,In_426);
or U350 (N_350,In_488,In_618);
and U351 (N_351,In_431,In_198);
and U352 (N_352,In_188,In_650);
xor U353 (N_353,In_187,In_203);
and U354 (N_354,In_220,In_396);
xnor U355 (N_355,In_181,In_21);
and U356 (N_356,In_100,In_746);
nand U357 (N_357,In_499,In_422);
or U358 (N_358,In_150,In_113);
or U359 (N_359,In_269,In_238);
and U360 (N_360,In_162,In_453);
and U361 (N_361,In_273,In_80);
nor U362 (N_362,In_25,In_647);
and U363 (N_363,In_156,In_335);
or U364 (N_364,In_135,In_486);
nand U365 (N_365,In_346,In_424);
nor U366 (N_366,In_81,In_639);
and U367 (N_367,In_398,In_70);
nor U368 (N_368,In_674,In_580);
and U369 (N_369,In_602,In_636);
and U370 (N_370,In_567,In_683);
or U371 (N_371,In_559,In_354);
or U372 (N_372,In_730,In_596);
nand U373 (N_373,In_342,In_9);
nand U374 (N_374,In_742,In_174);
or U375 (N_375,In_241,In_147);
nor U376 (N_376,In_48,In_380);
nand U377 (N_377,In_133,In_185);
or U378 (N_378,In_680,In_2);
nand U379 (N_379,In_240,In_289);
nand U380 (N_380,In_609,In_565);
and U381 (N_381,In_5,In_733);
nor U382 (N_382,In_614,In_109);
or U383 (N_383,In_697,In_343);
nor U384 (N_384,In_472,In_305);
nand U385 (N_385,In_729,In_583);
or U386 (N_386,In_720,In_365);
nor U387 (N_387,In_53,In_472);
and U388 (N_388,In_641,In_422);
nor U389 (N_389,In_73,In_731);
or U390 (N_390,In_546,In_537);
nand U391 (N_391,In_426,In_40);
and U392 (N_392,In_506,In_589);
xor U393 (N_393,In_669,In_476);
nand U394 (N_394,In_264,In_354);
nor U395 (N_395,In_345,In_119);
and U396 (N_396,In_87,In_662);
or U397 (N_397,In_390,In_408);
nor U398 (N_398,In_292,In_645);
nor U399 (N_399,In_223,In_325);
or U400 (N_400,In_702,In_359);
or U401 (N_401,In_384,In_235);
or U402 (N_402,In_543,In_749);
or U403 (N_403,In_719,In_258);
nor U404 (N_404,In_53,In_329);
nor U405 (N_405,In_65,In_262);
and U406 (N_406,In_435,In_341);
and U407 (N_407,In_270,In_626);
or U408 (N_408,In_45,In_477);
nor U409 (N_409,In_286,In_651);
nand U410 (N_410,In_39,In_143);
or U411 (N_411,In_171,In_608);
nor U412 (N_412,In_324,In_58);
nor U413 (N_413,In_632,In_153);
nand U414 (N_414,In_712,In_547);
nor U415 (N_415,In_355,In_499);
nand U416 (N_416,In_164,In_97);
and U417 (N_417,In_539,In_99);
nand U418 (N_418,In_24,In_502);
or U419 (N_419,In_402,In_243);
nor U420 (N_420,In_18,In_65);
nand U421 (N_421,In_418,In_590);
nand U422 (N_422,In_613,In_581);
or U423 (N_423,In_682,In_739);
nor U424 (N_424,In_645,In_406);
and U425 (N_425,In_74,In_29);
nand U426 (N_426,In_420,In_62);
nor U427 (N_427,In_46,In_491);
nor U428 (N_428,In_180,In_197);
and U429 (N_429,In_651,In_104);
and U430 (N_430,In_11,In_141);
and U431 (N_431,In_407,In_619);
nor U432 (N_432,In_282,In_551);
or U433 (N_433,In_450,In_707);
nand U434 (N_434,In_679,In_462);
and U435 (N_435,In_239,In_91);
nand U436 (N_436,In_272,In_413);
nor U437 (N_437,In_335,In_298);
nor U438 (N_438,In_446,In_545);
and U439 (N_439,In_216,In_668);
nor U440 (N_440,In_389,In_242);
nor U441 (N_441,In_612,In_632);
nor U442 (N_442,In_11,In_576);
nand U443 (N_443,In_589,In_230);
nor U444 (N_444,In_210,In_337);
nor U445 (N_445,In_312,In_114);
or U446 (N_446,In_686,In_437);
or U447 (N_447,In_727,In_712);
and U448 (N_448,In_166,In_1);
and U449 (N_449,In_350,In_283);
and U450 (N_450,In_140,In_90);
or U451 (N_451,In_220,In_565);
or U452 (N_452,In_183,In_544);
nand U453 (N_453,In_102,In_242);
or U454 (N_454,In_328,In_567);
nor U455 (N_455,In_183,In_334);
and U456 (N_456,In_372,In_278);
nand U457 (N_457,In_280,In_735);
and U458 (N_458,In_243,In_104);
nor U459 (N_459,In_409,In_509);
or U460 (N_460,In_663,In_57);
nor U461 (N_461,In_528,In_424);
nand U462 (N_462,In_448,In_501);
nor U463 (N_463,In_165,In_209);
and U464 (N_464,In_167,In_119);
and U465 (N_465,In_124,In_64);
and U466 (N_466,In_334,In_164);
nand U467 (N_467,In_106,In_60);
and U468 (N_468,In_36,In_143);
nand U469 (N_469,In_84,In_497);
or U470 (N_470,In_308,In_293);
or U471 (N_471,In_694,In_744);
nand U472 (N_472,In_719,In_361);
nor U473 (N_473,In_410,In_375);
or U474 (N_474,In_219,In_372);
and U475 (N_475,In_401,In_508);
or U476 (N_476,In_548,In_384);
nor U477 (N_477,In_34,In_744);
nor U478 (N_478,In_393,In_422);
nand U479 (N_479,In_720,In_320);
or U480 (N_480,In_644,In_303);
and U481 (N_481,In_615,In_251);
or U482 (N_482,In_38,In_23);
nand U483 (N_483,In_292,In_404);
nor U484 (N_484,In_60,In_466);
or U485 (N_485,In_487,In_37);
nor U486 (N_486,In_612,In_407);
and U487 (N_487,In_191,In_226);
nor U488 (N_488,In_214,In_644);
or U489 (N_489,In_148,In_174);
and U490 (N_490,In_685,In_513);
or U491 (N_491,In_188,In_388);
and U492 (N_492,In_412,In_273);
nor U493 (N_493,In_203,In_365);
or U494 (N_494,In_478,In_582);
or U495 (N_495,In_24,In_85);
xnor U496 (N_496,In_619,In_22);
nand U497 (N_497,In_233,In_460);
or U498 (N_498,In_302,In_218);
nor U499 (N_499,In_240,In_75);
nand U500 (N_500,In_630,In_52);
nor U501 (N_501,In_179,In_527);
and U502 (N_502,In_414,In_468);
nand U503 (N_503,In_372,In_743);
and U504 (N_504,In_541,In_652);
nor U505 (N_505,In_262,In_605);
nor U506 (N_506,In_686,In_618);
nor U507 (N_507,In_115,In_398);
nor U508 (N_508,In_470,In_205);
or U509 (N_509,In_210,In_45);
or U510 (N_510,In_540,In_586);
nor U511 (N_511,In_234,In_613);
or U512 (N_512,In_432,In_279);
nand U513 (N_513,In_166,In_370);
nor U514 (N_514,In_374,In_472);
and U515 (N_515,In_639,In_407);
nand U516 (N_516,In_713,In_193);
and U517 (N_517,In_170,In_658);
xor U518 (N_518,In_432,In_742);
xnor U519 (N_519,In_87,In_584);
and U520 (N_520,In_47,In_30);
nand U521 (N_521,In_217,In_198);
and U522 (N_522,In_264,In_574);
and U523 (N_523,In_37,In_610);
nand U524 (N_524,In_298,In_150);
or U525 (N_525,In_315,In_563);
and U526 (N_526,In_162,In_221);
nor U527 (N_527,In_176,In_282);
nor U528 (N_528,In_540,In_669);
nand U529 (N_529,In_151,In_351);
nand U530 (N_530,In_12,In_336);
or U531 (N_531,In_320,In_188);
and U532 (N_532,In_662,In_68);
nor U533 (N_533,In_489,In_493);
or U534 (N_534,In_121,In_581);
nand U535 (N_535,In_158,In_403);
and U536 (N_536,In_672,In_89);
nand U537 (N_537,In_491,In_290);
nand U538 (N_538,In_297,In_81);
and U539 (N_539,In_576,In_641);
xnor U540 (N_540,In_181,In_589);
nor U541 (N_541,In_288,In_303);
and U542 (N_542,In_374,In_101);
and U543 (N_543,In_335,In_700);
nor U544 (N_544,In_525,In_282);
nand U545 (N_545,In_105,In_742);
or U546 (N_546,In_455,In_457);
or U547 (N_547,In_352,In_395);
nor U548 (N_548,In_82,In_214);
and U549 (N_549,In_218,In_614);
and U550 (N_550,In_252,In_53);
nor U551 (N_551,In_707,In_260);
nor U552 (N_552,In_59,In_50);
or U553 (N_553,In_115,In_334);
and U554 (N_554,In_552,In_509);
or U555 (N_555,In_259,In_601);
nand U556 (N_556,In_140,In_559);
nor U557 (N_557,In_725,In_419);
nand U558 (N_558,In_631,In_294);
nor U559 (N_559,In_73,In_224);
nor U560 (N_560,In_645,In_589);
nand U561 (N_561,In_225,In_459);
nor U562 (N_562,In_457,In_375);
and U563 (N_563,In_268,In_286);
nand U564 (N_564,In_347,In_485);
nor U565 (N_565,In_490,In_658);
nand U566 (N_566,In_405,In_138);
nand U567 (N_567,In_478,In_166);
nor U568 (N_568,In_319,In_190);
nand U569 (N_569,In_185,In_72);
nand U570 (N_570,In_401,In_563);
nand U571 (N_571,In_61,In_591);
nand U572 (N_572,In_721,In_592);
nor U573 (N_573,In_382,In_69);
nand U574 (N_574,In_663,In_420);
or U575 (N_575,In_583,In_39);
or U576 (N_576,In_547,In_694);
nor U577 (N_577,In_744,In_191);
nor U578 (N_578,In_685,In_381);
or U579 (N_579,In_508,In_725);
nor U580 (N_580,In_391,In_458);
nand U581 (N_581,In_537,In_268);
nand U582 (N_582,In_353,In_618);
and U583 (N_583,In_389,In_39);
or U584 (N_584,In_42,In_194);
or U585 (N_585,In_127,In_478);
or U586 (N_586,In_332,In_202);
nor U587 (N_587,In_447,In_129);
and U588 (N_588,In_510,In_355);
and U589 (N_589,In_8,In_27);
nand U590 (N_590,In_190,In_307);
or U591 (N_591,In_591,In_653);
nor U592 (N_592,In_30,In_650);
nand U593 (N_593,In_342,In_428);
and U594 (N_594,In_191,In_397);
nand U595 (N_595,In_256,In_455);
nor U596 (N_596,In_673,In_9);
and U597 (N_597,In_202,In_368);
nor U598 (N_598,In_697,In_516);
and U599 (N_599,In_333,In_314);
or U600 (N_600,In_399,In_382);
and U601 (N_601,In_53,In_107);
and U602 (N_602,In_262,In_41);
nor U603 (N_603,In_193,In_424);
nor U604 (N_604,In_497,In_347);
or U605 (N_605,In_472,In_159);
and U606 (N_606,In_26,In_447);
nand U607 (N_607,In_86,In_164);
or U608 (N_608,In_446,In_203);
and U609 (N_609,In_743,In_574);
nand U610 (N_610,In_174,In_364);
and U611 (N_611,In_144,In_725);
nor U612 (N_612,In_645,In_476);
and U613 (N_613,In_621,In_711);
or U614 (N_614,In_150,In_205);
or U615 (N_615,In_553,In_606);
nand U616 (N_616,In_696,In_240);
nor U617 (N_617,In_216,In_693);
and U618 (N_618,In_360,In_675);
and U619 (N_619,In_270,In_115);
or U620 (N_620,In_353,In_535);
or U621 (N_621,In_160,In_44);
nand U622 (N_622,In_87,In_267);
or U623 (N_623,In_99,In_749);
and U624 (N_624,In_500,In_335);
or U625 (N_625,In_186,In_235);
nor U626 (N_626,In_457,In_402);
or U627 (N_627,In_737,In_310);
and U628 (N_628,In_576,In_492);
and U629 (N_629,In_332,In_75);
or U630 (N_630,In_532,In_499);
and U631 (N_631,In_682,In_66);
nand U632 (N_632,In_653,In_179);
nor U633 (N_633,In_143,In_352);
or U634 (N_634,In_574,In_217);
nor U635 (N_635,In_38,In_246);
nor U636 (N_636,In_1,In_506);
nand U637 (N_637,In_212,In_618);
nor U638 (N_638,In_12,In_232);
nand U639 (N_639,In_693,In_94);
and U640 (N_640,In_654,In_64);
or U641 (N_641,In_296,In_416);
and U642 (N_642,In_445,In_291);
or U643 (N_643,In_217,In_188);
or U644 (N_644,In_493,In_8);
or U645 (N_645,In_89,In_10);
or U646 (N_646,In_279,In_475);
or U647 (N_647,In_74,In_25);
and U648 (N_648,In_446,In_501);
nor U649 (N_649,In_738,In_443);
or U650 (N_650,In_720,In_201);
or U651 (N_651,In_273,In_625);
nand U652 (N_652,In_535,In_561);
or U653 (N_653,In_441,In_595);
and U654 (N_654,In_489,In_629);
and U655 (N_655,In_197,In_31);
nand U656 (N_656,In_121,In_20);
nand U657 (N_657,In_180,In_458);
and U658 (N_658,In_488,In_748);
nand U659 (N_659,In_53,In_212);
and U660 (N_660,In_309,In_436);
nand U661 (N_661,In_423,In_695);
and U662 (N_662,In_50,In_704);
nor U663 (N_663,In_608,In_519);
nand U664 (N_664,In_667,In_33);
nand U665 (N_665,In_115,In_731);
nand U666 (N_666,In_166,In_720);
nor U667 (N_667,In_656,In_348);
nor U668 (N_668,In_673,In_264);
or U669 (N_669,In_229,In_272);
nand U670 (N_670,In_191,In_540);
nand U671 (N_671,In_689,In_525);
nor U672 (N_672,In_164,In_254);
or U673 (N_673,In_452,In_144);
nand U674 (N_674,In_250,In_602);
nand U675 (N_675,In_200,In_625);
or U676 (N_676,In_237,In_511);
nor U677 (N_677,In_26,In_133);
nand U678 (N_678,In_42,In_550);
and U679 (N_679,In_312,In_68);
nor U680 (N_680,In_275,In_365);
nor U681 (N_681,In_195,In_511);
or U682 (N_682,In_425,In_491);
nand U683 (N_683,In_268,In_533);
or U684 (N_684,In_459,In_175);
nor U685 (N_685,In_336,In_317);
nand U686 (N_686,In_70,In_120);
and U687 (N_687,In_212,In_515);
nand U688 (N_688,In_476,In_689);
and U689 (N_689,In_448,In_399);
nor U690 (N_690,In_499,In_272);
nor U691 (N_691,In_429,In_593);
nand U692 (N_692,In_743,In_131);
and U693 (N_693,In_597,In_604);
or U694 (N_694,In_235,In_359);
nand U695 (N_695,In_571,In_34);
nand U696 (N_696,In_727,In_584);
nor U697 (N_697,In_105,In_67);
nand U698 (N_698,In_503,In_387);
nor U699 (N_699,In_252,In_570);
nand U700 (N_700,In_678,In_722);
nor U701 (N_701,In_713,In_434);
nor U702 (N_702,In_599,In_395);
and U703 (N_703,In_324,In_709);
nand U704 (N_704,In_558,In_24);
nor U705 (N_705,In_106,In_710);
or U706 (N_706,In_505,In_302);
nor U707 (N_707,In_283,In_522);
or U708 (N_708,In_162,In_462);
and U709 (N_709,In_519,In_658);
or U710 (N_710,In_547,In_128);
nand U711 (N_711,In_720,In_690);
and U712 (N_712,In_670,In_95);
nand U713 (N_713,In_546,In_245);
nor U714 (N_714,In_9,In_544);
and U715 (N_715,In_399,In_583);
nor U716 (N_716,In_665,In_97);
xnor U717 (N_717,In_15,In_527);
xnor U718 (N_718,In_228,In_656);
and U719 (N_719,In_488,In_41);
nand U720 (N_720,In_347,In_588);
and U721 (N_721,In_422,In_330);
and U722 (N_722,In_596,In_604);
nand U723 (N_723,In_117,In_460);
nor U724 (N_724,In_367,In_392);
or U725 (N_725,In_305,In_313);
and U726 (N_726,In_210,In_183);
nand U727 (N_727,In_226,In_568);
and U728 (N_728,In_328,In_77);
nor U729 (N_729,In_485,In_681);
and U730 (N_730,In_541,In_233);
nor U731 (N_731,In_616,In_652);
and U732 (N_732,In_213,In_643);
and U733 (N_733,In_653,In_364);
or U734 (N_734,In_7,In_561);
and U735 (N_735,In_152,In_257);
nand U736 (N_736,In_603,In_84);
and U737 (N_737,In_237,In_725);
and U738 (N_738,In_37,In_633);
nand U739 (N_739,In_594,In_636);
or U740 (N_740,In_237,In_528);
nand U741 (N_741,In_670,In_41);
nand U742 (N_742,In_71,In_624);
or U743 (N_743,In_41,In_216);
or U744 (N_744,In_107,In_28);
and U745 (N_745,In_74,In_638);
or U746 (N_746,In_16,In_158);
nor U747 (N_747,In_19,In_173);
nand U748 (N_748,In_518,In_690);
and U749 (N_749,In_497,In_53);
and U750 (N_750,In_126,In_548);
nor U751 (N_751,In_18,In_654);
nand U752 (N_752,In_390,In_557);
nor U753 (N_753,In_32,In_114);
and U754 (N_754,In_173,In_627);
nand U755 (N_755,In_0,In_495);
and U756 (N_756,In_319,In_501);
and U757 (N_757,In_302,In_119);
nand U758 (N_758,In_220,In_699);
nor U759 (N_759,In_333,In_446);
or U760 (N_760,In_477,In_641);
nor U761 (N_761,In_331,In_212);
nand U762 (N_762,In_738,In_702);
or U763 (N_763,In_74,In_631);
and U764 (N_764,In_408,In_595);
nand U765 (N_765,In_48,In_547);
nand U766 (N_766,In_127,In_324);
or U767 (N_767,In_100,In_426);
or U768 (N_768,In_625,In_189);
nand U769 (N_769,In_347,In_395);
or U770 (N_770,In_706,In_715);
or U771 (N_771,In_33,In_98);
or U772 (N_772,In_627,In_734);
nand U773 (N_773,In_629,In_646);
or U774 (N_774,In_323,In_462);
xor U775 (N_775,In_105,In_731);
nor U776 (N_776,In_20,In_192);
or U777 (N_777,In_199,In_238);
and U778 (N_778,In_352,In_609);
and U779 (N_779,In_656,In_710);
nor U780 (N_780,In_289,In_613);
nor U781 (N_781,In_483,In_212);
or U782 (N_782,In_666,In_619);
and U783 (N_783,In_84,In_563);
nor U784 (N_784,In_178,In_589);
xnor U785 (N_785,In_348,In_378);
or U786 (N_786,In_389,In_122);
and U787 (N_787,In_634,In_461);
and U788 (N_788,In_435,In_748);
and U789 (N_789,In_105,In_465);
nand U790 (N_790,In_688,In_674);
nor U791 (N_791,In_728,In_603);
nand U792 (N_792,In_734,In_584);
and U793 (N_793,In_463,In_713);
nor U794 (N_794,In_386,In_457);
nand U795 (N_795,In_533,In_382);
nand U796 (N_796,In_425,In_336);
nor U797 (N_797,In_635,In_115);
nand U798 (N_798,In_296,In_248);
and U799 (N_799,In_231,In_161);
nor U800 (N_800,In_51,In_571);
or U801 (N_801,In_253,In_410);
and U802 (N_802,In_749,In_591);
nor U803 (N_803,In_251,In_287);
and U804 (N_804,In_44,In_263);
and U805 (N_805,In_424,In_151);
or U806 (N_806,In_689,In_86);
and U807 (N_807,In_235,In_140);
nand U808 (N_808,In_509,In_525);
nand U809 (N_809,In_667,In_133);
or U810 (N_810,In_593,In_24);
nand U811 (N_811,In_199,In_316);
nand U812 (N_812,In_605,In_209);
and U813 (N_813,In_44,In_380);
and U814 (N_814,In_691,In_305);
nand U815 (N_815,In_597,In_735);
or U816 (N_816,In_377,In_518);
nand U817 (N_817,In_575,In_143);
or U818 (N_818,In_324,In_100);
nand U819 (N_819,In_650,In_238);
nor U820 (N_820,In_23,In_10);
and U821 (N_821,In_275,In_111);
nor U822 (N_822,In_574,In_674);
nand U823 (N_823,In_688,In_126);
and U824 (N_824,In_597,In_570);
and U825 (N_825,In_532,In_485);
nor U826 (N_826,In_380,In_111);
or U827 (N_827,In_106,In_24);
or U828 (N_828,In_379,In_248);
nand U829 (N_829,In_389,In_349);
nand U830 (N_830,In_429,In_75);
or U831 (N_831,In_9,In_405);
or U832 (N_832,In_18,In_618);
nor U833 (N_833,In_716,In_593);
nor U834 (N_834,In_568,In_19);
nor U835 (N_835,In_531,In_380);
nand U836 (N_836,In_667,In_389);
and U837 (N_837,In_560,In_498);
and U838 (N_838,In_744,In_311);
nand U839 (N_839,In_299,In_286);
or U840 (N_840,In_386,In_694);
and U841 (N_841,In_8,In_382);
and U842 (N_842,In_699,In_671);
and U843 (N_843,In_622,In_274);
or U844 (N_844,In_200,In_106);
or U845 (N_845,In_736,In_117);
or U846 (N_846,In_25,In_547);
nand U847 (N_847,In_295,In_63);
nor U848 (N_848,In_541,In_502);
or U849 (N_849,In_391,In_24);
and U850 (N_850,In_536,In_613);
nor U851 (N_851,In_389,In_459);
or U852 (N_852,In_284,In_493);
or U853 (N_853,In_17,In_308);
and U854 (N_854,In_7,In_304);
nor U855 (N_855,In_683,In_122);
or U856 (N_856,In_453,In_81);
and U857 (N_857,In_643,In_655);
and U858 (N_858,In_179,In_725);
or U859 (N_859,In_457,In_586);
and U860 (N_860,In_593,In_636);
and U861 (N_861,In_65,In_684);
nor U862 (N_862,In_441,In_649);
and U863 (N_863,In_139,In_361);
or U864 (N_864,In_188,In_464);
and U865 (N_865,In_133,In_266);
nor U866 (N_866,In_169,In_264);
or U867 (N_867,In_61,In_644);
or U868 (N_868,In_24,In_652);
nor U869 (N_869,In_8,In_177);
nor U870 (N_870,In_627,In_192);
or U871 (N_871,In_588,In_244);
and U872 (N_872,In_656,In_458);
nor U873 (N_873,In_683,In_95);
nand U874 (N_874,In_435,In_510);
and U875 (N_875,In_440,In_239);
nand U876 (N_876,In_377,In_459);
and U877 (N_877,In_695,In_542);
nor U878 (N_878,In_615,In_254);
or U879 (N_879,In_153,In_555);
or U880 (N_880,In_399,In_421);
or U881 (N_881,In_406,In_316);
nor U882 (N_882,In_589,In_428);
or U883 (N_883,In_91,In_396);
nor U884 (N_884,In_722,In_689);
and U885 (N_885,In_33,In_83);
or U886 (N_886,In_198,In_147);
nand U887 (N_887,In_398,In_337);
nor U888 (N_888,In_409,In_575);
or U889 (N_889,In_690,In_183);
and U890 (N_890,In_377,In_694);
nor U891 (N_891,In_426,In_613);
or U892 (N_892,In_118,In_100);
or U893 (N_893,In_78,In_598);
or U894 (N_894,In_230,In_454);
and U895 (N_895,In_280,In_724);
nand U896 (N_896,In_390,In_255);
xor U897 (N_897,In_516,In_521);
nand U898 (N_898,In_90,In_500);
nor U899 (N_899,In_460,In_687);
nor U900 (N_900,In_616,In_497);
or U901 (N_901,In_515,In_732);
or U902 (N_902,In_202,In_576);
and U903 (N_903,In_692,In_127);
nand U904 (N_904,In_407,In_347);
nor U905 (N_905,In_577,In_344);
and U906 (N_906,In_724,In_576);
or U907 (N_907,In_309,In_315);
or U908 (N_908,In_103,In_584);
and U909 (N_909,In_191,In_147);
and U910 (N_910,In_292,In_719);
nand U911 (N_911,In_737,In_356);
or U912 (N_912,In_607,In_372);
nor U913 (N_913,In_548,In_2);
nand U914 (N_914,In_462,In_19);
and U915 (N_915,In_96,In_59);
and U916 (N_916,In_153,In_507);
and U917 (N_917,In_551,In_626);
or U918 (N_918,In_104,In_301);
or U919 (N_919,In_348,In_452);
or U920 (N_920,In_460,In_699);
nand U921 (N_921,In_585,In_478);
or U922 (N_922,In_232,In_335);
and U923 (N_923,In_123,In_556);
nor U924 (N_924,In_203,In_195);
and U925 (N_925,In_728,In_669);
or U926 (N_926,In_83,In_657);
and U927 (N_927,In_314,In_143);
or U928 (N_928,In_699,In_388);
nand U929 (N_929,In_49,In_402);
or U930 (N_930,In_182,In_237);
nor U931 (N_931,In_369,In_87);
nand U932 (N_932,In_493,In_299);
and U933 (N_933,In_49,In_185);
nor U934 (N_934,In_288,In_347);
or U935 (N_935,In_64,In_681);
nand U936 (N_936,In_331,In_655);
nor U937 (N_937,In_744,In_95);
and U938 (N_938,In_128,In_409);
or U939 (N_939,In_714,In_677);
nand U940 (N_940,In_341,In_196);
nand U941 (N_941,In_65,In_696);
xor U942 (N_942,In_25,In_158);
and U943 (N_943,In_502,In_43);
or U944 (N_944,In_112,In_475);
nor U945 (N_945,In_299,In_199);
and U946 (N_946,In_704,In_546);
nor U947 (N_947,In_120,In_514);
and U948 (N_948,In_65,In_679);
and U949 (N_949,In_254,In_394);
or U950 (N_950,In_576,In_165);
or U951 (N_951,In_253,In_415);
or U952 (N_952,In_150,In_681);
nand U953 (N_953,In_68,In_160);
nor U954 (N_954,In_627,In_704);
and U955 (N_955,In_723,In_183);
or U956 (N_956,In_170,In_624);
nor U957 (N_957,In_48,In_77);
or U958 (N_958,In_13,In_568);
and U959 (N_959,In_296,In_139);
or U960 (N_960,In_422,In_540);
nor U961 (N_961,In_179,In_538);
nand U962 (N_962,In_255,In_170);
nand U963 (N_963,In_609,In_560);
or U964 (N_964,In_152,In_245);
and U965 (N_965,In_384,In_321);
or U966 (N_966,In_553,In_646);
and U967 (N_967,In_259,In_585);
or U968 (N_968,In_179,In_576);
nand U969 (N_969,In_288,In_503);
nand U970 (N_970,In_646,In_271);
or U971 (N_971,In_203,In_285);
or U972 (N_972,In_588,In_284);
or U973 (N_973,In_612,In_332);
nor U974 (N_974,In_277,In_150);
or U975 (N_975,In_391,In_488);
nor U976 (N_976,In_51,In_348);
and U977 (N_977,In_152,In_158);
and U978 (N_978,In_659,In_311);
nor U979 (N_979,In_141,In_45);
nand U980 (N_980,In_193,In_603);
and U981 (N_981,In_349,In_0);
nand U982 (N_982,In_214,In_710);
nor U983 (N_983,In_458,In_222);
nor U984 (N_984,In_297,In_514);
and U985 (N_985,In_731,In_740);
or U986 (N_986,In_189,In_594);
and U987 (N_987,In_728,In_670);
nand U988 (N_988,In_203,In_144);
nand U989 (N_989,In_62,In_27);
and U990 (N_990,In_677,In_105);
nor U991 (N_991,In_441,In_588);
and U992 (N_992,In_400,In_465);
or U993 (N_993,In_253,In_1);
or U994 (N_994,In_457,In_281);
nand U995 (N_995,In_49,In_600);
or U996 (N_996,In_387,In_326);
and U997 (N_997,In_124,In_68);
or U998 (N_998,In_13,In_580);
nand U999 (N_999,In_713,In_436);
or U1000 (N_1000,In_9,In_272);
nor U1001 (N_1001,In_743,In_167);
and U1002 (N_1002,In_14,In_296);
or U1003 (N_1003,In_137,In_623);
nor U1004 (N_1004,In_476,In_466);
or U1005 (N_1005,In_637,In_61);
nor U1006 (N_1006,In_383,In_531);
or U1007 (N_1007,In_709,In_209);
nor U1008 (N_1008,In_742,In_508);
and U1009 (N_1009,In_441,In_637);
and U1010 (N_1010,In_227,In_236);
nand U1011 (N_1011,In_644,In_487);
nand U1012 (N_1012,In_652,In_585);
and U1013 (N_1013,In_354,In_742);
or U1014 (N_1014,In_280,In_598);
nand U1015 (N_1015,In_250,In_146);
or U1016 (N_1016,In_232,In_258);
nand U1017 (N_1017,In_683,In_123);
nor U1018 (N_1018,In_566,In_454);
nand U1019 (N_1019,In_654,In_89);
and U1020 (N_1020,In_184,In_614);
and U1021 (N_1021,In_290,In_485);
and U1022 (N_1022,In_442,In_726);
or U1023 (N_1023,In_148,In_373);
and U1024 (N_1024,In_278,In_158);
nand U1025 (N_1025,In_20,In_35);
nor U1026 (N_1026,In_465,In_430);
nor U1027 (N_1027,In_71,In_630);
and U1028 (N_1028,In_687,In_192);
nand U1029 (N_1029,In_265,In_746);
nand U1030 (N_1030,In_141,In_429);
nand U1031 (N_1031,In_445,In_564);
or U1032 (N_1032,In_405,In_140);
nand U1033 (N_1033,In_42,In_649);
and U1034 (N_1034,In_356,In_580);
and U1035 (N_1035,In_434,In_466);
and U1036 (N_1036,In_254,In_578);
and U1037 (N_1037,In_247,In_163);
nor U1038 (N_1038,In_233,In_556);
and U1039 (N_1039,In_297,In_557);
nor U1040 (N_1040,In_233,In_183);
or U1041 (N_1041,In_449,In_474);
nor U1042 (N_1042,In_646,In_483);
nand U1043 (N_1043,In_607,In_81);
or U1044 (N_1044,In_314,In_42);
nor U1045 (N_1045,In_218,In_736);
nand U1046 (N_1046,In_75,In_286);
and U1047 (N_1047,In_318,In_286);
nand U1048 (N_1048,In_375,In_29);
or U1049 (N_1049,In_490,In_318);
nand U1050 (N_1050,In_47,In_499);
or U1051 (N_1051,In_690,In_560);
nand U1052 (N_1052,In_312,In_151);
nand U1053 (N_1053,In_362,In_545);
nand U1054 (N_1054,In_372,In_66);
nand U1055 (N_1055,In_309,In_13);
nor U1056 (N_1056,In_210,In_18);
or U1057 (N_1057,In_405,In_360);
and U1058 (N_1058,In_636,In_403);
nor U1059 (N_1059,In_287,In_722);
nor U1060 (N_1060,In_21,In_495);
or U1061 (N_1061,In_534,In_536);
and U1062 (N_1062,In_677,In_348);
or U1063 (N_1063,In_531,In_118);
nor U1064 (N_1064,In_113,In_626);
nor U1065 (N_1065,In_130,In_656);
nor U1066 (N_1066,In_224,In_470);
nor U1067 (N_1067,In_107,In_216);
and U1068 (N_1068,In_578,In_0);
nor U1069 (N_1069,In_405,In_118);
or U1070 (N_1070,In_447,In_39);
or U1071 (N_1071,In_326,In_544);
and U1072 (N_1072,In_607,In_359);
or U1073 (N_1073,In_83,In_621);
nor U1074 (N_1074,In_227,In_622);
or U1075 (N_1075,In_575,In_531);
or U1076 (N_1076,In_381,In_408);
nand U1077 (N_1077,In_495,In_520);
nor U1078 (N_1078,In_537,In_656);
xor U1079 (N_1079,In_557,In_188);
or U1080 (N_1080,In_749,In_155);
nor U1081 (N_1081,In_291,In_183);
nor U1082 (N_1082,In_733,In_344);
nor U1083 (N_1083,In_480,In_537);
nor U1084 (N_1084,In_640,In_53);
or U1085 (N_1085,In_468,In_349);
nand U1086 (N_1086,In_41,In_699);
nor U1087 (N_1087,In_744,In_338);
nand U1088 (N_1088,In_582,In_586);
and U1089 (N_1089,In_320,In_143);
or U1090 (N_1090,In_637,In_97);
nor U1091 (N_1091,In_115,In_205);
or U1092 (N_1092,In_632,In_415);
nand U1093 (N_1093,In_115,In_534);
nor U1094 (N_1094,In_561,In_314);
nand U1095 (N_1095,In_180,In_355);
nand U1096 (N_1096,In_280,In_579);
or U1097 (N_1097,In_644,In_342);
and U1098 (N_1098,In_550,In_173);
nor U1099 (N_1099,In_694,In_327);
and U1100 (N_1100,In_516,In_186);
nor U1101 (N_1101,In_362,In_578);
and U1102 (N_1102,In_691,In_233);
nand U1103 (N_1103,In_165,In_436);
and U1104 (N_1104,In_463,In_409);
or U1105 (N_1105,In_73,In_338);
or U1106 (N_1106,In_209,In_97);
nand U1107 (N_1107,In_1,In_157);
nor U1108 (N_1108,In_364,In_316);
and U1109 (N_1109,In_629,In_430);
or U1110 (N_1110,In_474,In_261);
and U1111 (N_1111,In_391,In_541);
and U1112 (N_1112,In_329,In_508);
nand U1113 (N_1113,In_38,In_576);
and U1114 (N_1114,In_47,In_508);
and U1115 (N_1115,In_175,In_390);
and U1116 (N_1116,In_548,In_191);
nand U1117 (N_1117,In_277,In_181);
and U1118 (N_1118,In_374,In_408);
nand U1119 (N_1119,In_175,In_517);
or U1120 (N_1120,In_0,In_429);
and U1121 (N_1121,In_532,In_414);
or U1122 (N_1122,In_41,In_462);
nor U1123 (N_1123,In_534,In_716);
or U1124 (N_1124,In_366,In_412);
nand U1125 (N_1125,In_128,In_575);
or U1126 (N_1126,In_587,In_201);
nor U1127 (N_1127,In_253,In_44);
nor U1128 (N_1128,In_169,In_127);
nand U1129 (N_1129,In_161,In_138);
nand U1130 (N_1130,In_725,In_493);
or U1131 (N_1131,In_374,In_16);
xnor U1132 (N_1132,In_435,In_468);
nand U1133 (N_1133,In_93,In_26);
nor U1134 (N_1134,In_742,In_583);
nor U1135 (N_1135,In_464,In_333);
and U1136 (N_1136,In_445,In_582);
and U1137 (N_1137,In_38,In_677);
nor U1138 (N_1138,In_332,In_271);
and U1139 (N_1139,In_400,In_439);
and U1140 (N_1140,In_173,In_518);
or U1141 (N_1141,In_646,In_129);
nand U1142 (N_1142,In_103,In_382);
nor U1143 (N_1143,In_173,In_165);
nor U1144 (N_1144,In_227,In_36);
nand U1145 (N_1145,In_75,In_315);
nand U1146 (N_1146,In_29,In_711);
or U1147 (N_1147,In_743,In_427);
nor U1148 (N_1148,In_11,In_493);
nor U1149 (N_1149,In_671,In_623);
nand U1150 (N_1150,In_337,In_190);
nand U1151 (N_1151,In_182,In_31);
or U1152 (N_1152,In_263,In_189);
and U1153 (N_1153,In_338,In_66);
and U1154 (N_1154,In_65,In_665);
nand U1155 (N_1155,In_248,In_617);
or U1156 (N_1156,In_189,In_429);
nor U1157 (N_1157,In_449,In_378);
or U1158 (N_1158,In_574,In_269);
nor U1159 (N_1159,In_232,In_552);
nand U1160 (N_1160,In_519,In_174);
and U1161 (N_1161,In_404,In_29);
and U1162 (N_1162,In_707,In_370);
and U1163 (N_1163,In_198,In_587);
nand U1164 (N_1164,In_604,In_27);
nor U1165 (N_1165,In_300,In_267);
nand U1166 (N_1166,In_69,In_570);
nand U1167 (N_1167,In_567,In_703);
and U1168 (N_1168,In_116,In_128);
nand U1169 (N_1169,In_527,In_683);
or U1170 (N_1170,In_526,In_83);
or U1171 (N_1171,In_211,In_96);
and U1172 (N_1172,In_197,In_177);
and U1173 (N_1173,In_735,In_221);
and U1174 (N_1174,In_270,In_91);
nand U1175 (N_1175,In_610,In_358);
or U1176 (N_1176,In_438,In_502);
nor U1177 (N_1177,In_657,In_710);
and U1178 (N_1178,In_615,In_72);
nor U1179 (N_1179,In_603,In_638);
and U1180 (N_1180,In_320,In_2);
nor U1181 (N_1181,In_28,In_529);
and U1182 (N_1182,In_146,In_611);
nand U1183 (N_1183,In_558,In_17);
and U1184 (N_1184,In_168,In_476);
nor U1185 (N_1185,In_587,In_44);
and U1186 (N_1186,In_366,In_533);
nand U1187 (N_1187,In_570,In_644);
nor U1188 (N_1188,In_194,In_119);
nor U1189 (N_1189,In_282,In_708);
and U1190 (N_1190,In_561,In_609);
nand U1191 (N_1191,In_256,In_89);
nand U1192 (N_1192,In_404,In_443);
or U1193 (N_1193,In_115,In_603);
nor U1194 (N_1194,In_191,In_713);
and U1195 (N_1195,In_687,In_684);
nand U1196 (N_1196,In_162,In_377);
or U1197 (N_1197,In_474,In_349);
nand U1198 (N_1198,In_172,In_202);
or U1199 (N_1199,In_301,In_71);
nor U1200 (N_1200,In_19,In_336);
nand U1201 (N_1201,In_601,In_626);
nor U1202 (N_1202,In_535,In_332);
and U1203 (N_1203,In_469,In_255);
nand U1204 (N_1204,In_109,In_575);
nand U1205 (N_1205,In_639,In_514);
nand U1206 (N_1206,In_692,In_639);
nand U1207 (N_1207,In_546,In_577);
nand U1208 (N_1208,In_290,In_747);
and U1209 (N_1209,In_100,In_716);
and U1210 (N_1210,In_211,In_45);
nand U1211 (N_1211,In_75,In_64);
and U1212 (N_1212,In_630,In_250);
or U1213 (N_1213,In_470,In_63);
and U1214 (N_1214,In_320,In_510);
or U1215 (N_1215,In_400,In_637);
nand U1216 (N_1216,In_236,In_538);
nor U1217 (N_1217,In_594,In_461);
xnor U1218 (N_1218,In_253,In_73);
nor U1219 (N_1219,In_256,In_635);
nor U1220 (N_1220,In_737,In_605);
or U1221 (N_1221,In_305,In_702);
nor U1222 (N_1222,In_72,In_697);
nor U1223 (N_1223,In_577,In_607);
nor U1224 (N_1224,In_399,In_298);
and U1225 (N_1225,In_43,In_185);
or U1226 (N_1226,In_301,In_154);
or U1227 (N_1227,In_608,In_55);
and U1228 (N_1228,In_424,In_546);
and U1229 (N_1229,In_166,In_630);
nand U1230 (N_1230,In_77,In_690);
or U1231 (N_1231,In_136,In_137);
nor U1232 (N_1232,In_481,In_230);
xor U1233 (N_1233,In_261,In_224);
and U1234 (N_1234,In_681,In_625);
and U1235 (N_1235,In_42,In_665);
nand U1236 (N_1236,In_393,In_577);
nor U1237 (N_1237,In_306,In_505);
nor U1238 (N_1238,In_125,In_133);
nand U1239 (N_1239,In_453,In_2);
nor U1240 (N_1240,In_686,In_221);
and U1241 (N_1241,In_517,In_488);
or U1242 (N_1242,In_541,In_180);
nor U1243 (N_1243,In_86,In_96);
xor U1244 (N_1244,In_130,In_94);
or U1245 (N_1245,In_447,In_488);
nand U1246 (N_1246,In_196,In_303);
or U1247 (N_1247,In_163,In_323);
nor U1248 (N_1248,In_496,In_475);
or U1249 (N_1249,In_405,In_426);
nor U1250 (N_1250,In_608,In_189);
nand U1251 (N_1251,In_544,In_359);
nand U1252 (N_1252,In_742,In_601);
nor U1253 (N_1253,In_738,In_82);
and U1254 (N_1254,In_749,In_248);
nor U1255 (N_1255,In_251,In_740);
or U1256 (N_1256,In_587,In_241);
nand U1257 (N_1257,In_452,In_22);
or U1258 (N_1258,In_177,In_110);
and U1259 (N_1259,In_79,In_561);
nor U1260 (N_1260,In_20,In_191);
and U1261 (N_1261,In_332,In_446);
nor U1262 (N_1262,In_484,In_743);
nand U1263 (N_1263,In_379,In_314);
or U1264 (N_1264,In_540,In_75);
or U1265 (N_1265,In_636,In_268);
nor U1266 (N_1266,In_658,In_25);
and U1267 (N_1267,In_233,In_630);
or U1268 (N_1268,In_578,In_736);
or U1269 (N_1269,In_703,In_84);
nor U1270 (N_1270,In_95,In_368);
nand U1271 (N_1271,In_253,In_450);
nor U1272 (N_1272,In_420,In_630);
or U1273 (N_1273,In_423,In_256);
or U1274 (N_1274,In_25,In_443);
and U1275 (N_1275,In_146,In_615);
and U1276 (N_1276,In_697,In_356);
or U1277 (N_1277,In_478,In_295);
or U1278 (N_1278,In_700,In_552);
and U1279 (N_1279,In_655,In_379);
and U1280 (N_1280,In_135,In_251);
and U1281 (N_1281,In_132,In_661);
nor U1282 (N_1282,In_514,In_58);
nand U1283 (N_1283,In_479,In_222);
or U1284 (N_1284,In_405,In_610);
nor U1285 (N_1285,In_86,In_198);
and U1286 (N_1286,In_495,In_395);
or U1287 (N_1287,In_621,In_563);
or U1288 (N_1288,In_417,In_168);
nor U1289 (N_1289,In_597,In_243);
or U1290 (N_1290,In_415,In_193);
and U1291 (N_1291,In_746,In_282);
nand U1292 (N_1292,In_150,In_474);
xnor U1293 (N_1293,In_257,In_220);
and U1294 (N_1294,In_576,In_325);
nor U1295 (N_1295,In_630,In_676);
and U1296 (N_1296,In_262,In_739);
and U1297 (N_1297,In_55,In_117);
nor U1298 (N_1298,In_206,In_661);
nor U1299 (N_1299,In_352,In_677);
or U1300 (N_1300,In_141,In_215);
nand U1301 (N_1301,In_165,In_356);
or U1302 (N_1302,In_698,In_743);
nor U1303 (N_1303,In_288,In_386);
nor U1304 (N_1304,In_410,In_94);
or U1305 (N_1305,In_323,In_431);
or U1306 (N_1306,In_466,In_601);
or U1307 (N_1307,In_19,In_538);
or U1308 (N_1308,In_321,In_450);
nor U1309 (N_1309,In_432,In_405);
and U1310 (N_1310,In_387,In_92);
and U1311 (N_1311,In_387,In_230);
nand U1312 (N_1312,In_678,In_494);
and U1313 (N_1313,In_496,In_399);
nand U1314 (N_1314,In_123,In_260);
nor U1315 (N_1315,In_499,In_309);
nand U1316 (N_1316,In_719,In_224);
nand U1317 (N_1317,In_127,In_690);
nand U1318 (N_1318,In_50,In_573);
nand U1319 (N_1319,In_743,In_91);
and U1320 (N_1320,In_717,In_491);
xor U1321 (N_1321,In_258,In_645);
nand U1322 (N_1322,In_318,In_101);
or U1323 (N_1323,In_257,In_82);
nand U1324 (N_1324,In_104,In_573);
and U1325 (N_1325,In_220,In_176);
nand U1326 (N_1326,In_18,In_103);
nand U1327 (N_1327,In_307,In_203);
nand U1328 (N_1328,In_331,In_713);
or U1329 (N_1329,In_273,In_534);
nor U1330 (N_1330,In_95,In_13);
nor U1331 (N_1331,In_494,In_639);
or U1332 (N_1332,In_610,In_148);
nor U1333 (N_1333,In_728,In_509);
nand U1334 (N_1334,In_742,In_200);
and U1335 (N_1335,In_668,In_684);
nor U1336 (N_1336,In_302,In_238);
nor U1337 (N_1337,In_228,In_528);
or U1338 (N_1338,In_3,In_661);
nor U1339 (N_1339,In_4,In_472);
and U1340 (N_1340,In_158,In_7);
or U1341 (N_1341,In_375,In_507);
nand U1342 (N_1342,In_293,In_20);
nand U1343 (N_1343,In_664,In_424);
nand U1344 (N_1344,In_337,In_674);
or U1345 (N_1345,In_56,In_420);
nor U1346 (N_1346,In_272,In_58);
nand U1347 (N_1347,In_195,In_236);
nor U1348 (N_1348,In_394,In_607);
or U1349 (N_1349,In_639,In_379);
or U1350 (N_1350,In_143,In_239);
and U1351 (N_1351,In_201,In_74);
nor U1352 (N_1352,In_4,In_197);
nor U1353 (N_1353,In_90,In_203);
nand U1354 (N_1354,In_73,In_479);
and U1355 (N_1355,In_508,In_679);
or U1356 (N_1356,In_561,In_268);
nand U1357 (N_1357,In_533,In_263);
and U1358 (N_1358,In_333,In_136);
or U1359 (N_1359,In_559,In_580);
nor U1360 (N_1360,In_431,In_584);
and U1361 (N_1361,In_306,In_204);
nor U1362 (N_1362,In_429,In_605);
or U1363 (N_1363,In_68,In_167);
nor U1364 (N_1364,In_14,In_452);
nand U1365 (N_1365,In_454,In_519);
or U1366 (N_1366,In_728,In_269);
nand U1367 (N_1367,In_501,In_741);
nor U1368 (N_1368,In_538,In_241);
nand U1369 (N_1369,In_414,In_101);
nand U1370 (N_1370,In_603,In_521);
and U1371 (N_1371,In_356,In_685);
nor U1372 (N_1372,In_573,In_243);
nand U1373 (N_1373,In_588,In_472);
nor U1374 (N_1374,In_246,In_348);
nor U1375 (N_1375,In_58,In_313);
and U1376 (N_1376,In_376,In_349);
and U1377 (N_1377,In_719,In_238);
nor U1378 (N_1378,In_262,In_101);
or U1379 (N_1379,In_82,In_477);
nor U1380 (N_1380,In_253,In_104);
nor U1381 (N_1381,In_89,In_123);
or U1382 (N_1382,In_522,In_222);
nand U1383 (N_1383,In_567,In_380);
and U1384 (N_1384,In_348,In_620);
nand U1385 (N_1385,In_423,In_492);
nand U1386 (N_1386,In_663,In_408);
nand U1387 (N_1387,In_728,In_75);
or U1388 (N_1388,In_565,In_430);
and U1389 (N_1389,In_232,In_162);
nand U1390 (N_1390,In_150,In_395);
nor U1391 (N_1391,In_28,In_363);
nand U1392 (N_1392,In_187,In_499);
or U1393 (N_1393,In_224,In_147);
and U1394 (N_1394,In_513,In_483);
nor U1395 (N_1395,In_602,In_119);
nor U1396 (N_1396,In_490,In_480);
nand U1397 (N_1397,In_219,In_413);
and U1398 (N_1398,In_157,In_597);
or U1399 (N_1399,In_25,In_316);
or U1400 (N_1400,In_44,In_642);
nor U1401 (N_1401,In_562,In_335);
nor U1402 (N_1402,In_602,In_65);
and U1403 (N_1403,In_631,In_449);
and U1404 (N_1404,In_253,In_209);
nor U1405 (N_1405,In_431,In_506);
and U1406 (N_1406,In_698,In_359);
nand U1407 (N_1407,In_315,In_709);
and U1408 (N_1408,In_540,In_99);
nor U1409 (N_1409,In_79,In_607);
nor U1410 (N_1410,In_502,In_324);
or U1411 (N_1411,In_509,In_125);
or U1412 (N_1412,In_213,In_729);
and U1413 (N_1413,In_41,In_379);
or U1414 (N_1414,In_21,In_211);
nor U1415 (N_1415,In_243,In_248);
nor U1416 (N_1416,In_121,In_744);
and U1417 (N_1417,In_292,In_473);
nand U1418 (N_1418,In_45,In_719);
and U1419 (N_1419,In_2,In_325);
or U1420 (N_1420,In_463,In_737);
and U1421 (N_1421,In_449,In_173);
nor U1422 (N_1422,In_590,In_651);
or U1423 (N_1423,In_417,In_326);
or U1424 (N_1424,In_456,In_213);
or U1425 (N_1425,In_711,In_641);
and U1426 (N_1426,In_356,In_145);
and U1427 (N_1427,In_228,In_222);
nor U1428 (N_1428,In_336,In_741);
or U1429 (N_1429,In_79,In_374);
and U1430 (N_1430,In_262,In_205);
or U1431 (N_1431,In_485,In_733);
and U1432 (N_1432,In_142,In_134);
nand U1433 (N_1433,In_320,In_460);
nor U1434 (N_1434,In_620,In_669);
nand U1435 (N_1435,In_92,In_165);
nand U1436 (N_1436,In_633,In_721);
nor U1437 (N_1437,In_532,In_561);
or U1438 (N_1438,In_115,In_152);
nand U1439 (N_1439,In_694,In_636);
and U1440 (N_1440,In_67,In_87);
nand U1441 (N_1441,In_726,In_35);
nand U1442 (N_1442,In_120,In_122);
nand U1443 (N_1443,In_408,In_180);
nand U1444 (N_1444,In_220,In_695);
nand U1445 (N_1445,In_120,In_552);
and U1446 (N_1446,In_146,In_487);
and U1447 (N_1447,In_487,In_624);
nand U1448 (N_1448,In_257,In_639);
and U1449 (N_1449,In_411,In_78);
and U1450 (N_1450,In_341,In_400);
xor U1451 (N_1451,In_153,In_254);
or U1452 (N_1452,In_465,In_526);
and U1453 (N_1453,In_375,In_333);
nand U1454 (N_1454,In_504,In_21);
nor U1455 (N_1455,In_132,In_317);
xnor U1456 (N_1456,In_542,In_674);
nand U1457 (N_1457,In_165,In_503);
nor U1458 (N_1458,In_369,In_586);
nor U1459 (N_1459,In_697,In_83);
nor U1460 (N_1460,In_213,In_579);
or U1461 (N_1461,In_409,In_340);
nand U1462 (N_1462,In_681,In_115);
nand U1463 (N_1463,In_706,In_210);
and U1464 (N_1464,In_448,In_659);
or U1465 (N_1465,In_168,In_210);
nand U1466 (N_1466,In_12,In_448);
and U1467 (N_1467,In_176,In_724);
and U1468 (N_1468,In_659,In_367);
nand U1469 (N_1469,In_703,In_579);
and U1470 (N_1470,In_401,In_34);
nand U1471 (N_1471,In_609,In_728);
or U1472 (N_1472,In_433,In_408);
and U1473 (N_1473,In_153,In_702);
and U1474 (N_1474,In_412,In_317);
nand U1475 (N_1475,In_24,In_356);
nor U1476 (N_1476,In_9,In_63);
and U1477 (N_1477,In_236,In_606);
nor U1478 (N_1478,In_581,In_460);
nor U1479 (N_1479,In_710,In_345);
nor U1480 (N_1480,In_96,In_227);
and U1481 (N_1481,In_45,In_579);
or U1482 (N_1482,In_423,In_227);
nor U1483 (N_1483,In_403,In_19);
and U1484 (N_1484,In_89,In_141);
nand U1485 (N_1485,In_95,In_237);
and U1486 (N_1486,In_70,In_305);
and U1487 (N_1487,In_323,In_86);
or U1488 (N_1488,In_103,In_439);
and U1489 (N_1489,In_188,In_246);
or U1490 (N_1490,In_400,In_723);
nand U1491 (N_1491,In_57,In_551);
nand U1492 (N_1492,In_712,In_637);
nand U1493 (N_1493,In_667,In_281);
and U1494 (N_1494,In_21,In_53);
nor U1495 (N_1495,In_266,In_112);
nand U1496 (N_1496,In_481,In_573);
or U1497 (N_1497,In_10,In_688);
nor U1498 (N_1498,In_87,In_748);
nand U1499 (N_1499,In_684,In_529);
nor U1500 (N_1500,In_99,In_571);
nand U1501 (N_1501,In_447,In_737);
nand U1502 (N_1502,In_296,In_640);
nor U1503 (N_1503,In_69,In_122);
and U1504 (N_1504,In_72,In_354);
nor U1505 (N_1505,In_17,In_312);
or U1506 (N_1506,In_202,In_310);
or U1507 (N_1507,In_411,In_52);
nand U1508 (N_1508,In_500,In_685);
nand U1509 (N_1509,In_252,In_552);
nand U1510 (N_1510,In_120,In_501);
nor U1511 (N_1511,In_148,In_166);
nand U1512 (N_1512,In_21,In_533);
and U1513 (N_1513,In_427,In_535);
nand U1514 (N_1514,In_97,In_118);
nor U1515 (N_1515,In_225,In_527);
or U1516 (N_1516,In_406,In_367);
and U1517 (N_1517,In_643,In_257);
nor U1518 (N_1518,In_247,In_279);
nand U1519 (N_1519,In_595,In_678);
and U1520 (N_1520,In_222,In_484);
nand U1521 (N_1521,In_9,In_735);
nor U1522 (N_1522,In_260,In_574);
nor U1523 (N_1523,In_252,In_715);
and U1524 (N_1524,In_224,In_515);
nand U1525 (N_1525,In_624,In_195);
and U1526 (N_1526,In_650,In_509);
nor U1527 (N_1527,In_515,In_602);
nand U1528 (N_1528,In_185,In_117);
and U1529 (N_1529,In_346,In_522);
nand U1530 (N_1530,In_452,In_705);
or U1531 (N_1531,In_11,In_537);
and U1532 (N_1532,In_83,In_309);
nand U1533 (N_1533,In_427,In_183);
nor U1534 (N_1534,In_354,In_211);
or U1535 (N_1535,In_388,In_494);
and U1536 (N_1536,In_174,In_27);
nand U1537 (N_1537,In_664,In_537);
and U1538 (N_1538,In_358,In_306);
nand U1539 (N_1539,In_107,In_51);
or U1540 (N_1540,In_298,In_14);
and U1541 (N_1541,In_513,In_489);
nor U1542 (N_1542,In_208,In_294);
nand U1543 (N_1543,In_654,In_243);
or U1544 (N_1544,In_701,In_554);
and U1545 (N_1545,In_360,In_447);
nand U1546 (N_1546,In_345,In_245);
nand U1547 (N_1547,In_298,In_371);
and U1548 (N_1548,In_579,In_50);
nor U1549 (N_1549,In_457,In_666);
and U1550 (N_1550,In_390,In_539);
and U1551 (N_1551,In_150,In_316);
and U1552 (N_1552,In_295,In_242);
and U1553 (N_1553,In_182,In_582);
nor U1554 (N_1554,In_134,In_111);
nand U1555 (N_1555,In_271,In_478);
or U1556 (N_1556,In_533,In_282);
nand U1557 (N_1557,In_236,In_419);
nor U1558 (N_1558,In_138,In_607);
nor U1559 (N_1559,In_220,In_743);
or U1560 (N_1560,In_288,In_86);
and U1561 (N_1561,In_627,In_684);
and U1562 (N_1562,In_76,In_664);
or U1563 (N_1563,In_590,In_39);
xor U1564 (N_1564,In_429,In_123);
nor U1565 (N_1565,In_560,In_579);
nor U1566 (N_1566,In_678,In_261);
nand U1567 (N_1567,In_600,In_603);
xor U1568 (N_1568,In_103,In_101);
or U1569 (N_1569,In_98,In_34);
and U1570 (N_1570,In_210,In_280);
nand U1571 (N_1571,In_215,In_228);
and U1572 (N_1572,In_668,In_294);
nor U1573 (N_1573,In_664,In_732);
and U1574 (N_1574,In_409,In_691);
or U1575 (N_1575,In_50,In_128);
and U1576 (N_1576,In_21,In_693);
nand U1577 (N_1577,In_175,In_297);
and U1578 (N_1578,In_147,In_583);
nand U1579 (N_1579,In_680,In_395);
or U1580 (N_1580,In_400,In_639);
and U1581 (N_1581,In_688,In_227);
and U1582 (N_1582,In_401,In_464);
and U1583 (N_1583,In_178,In_713);
and U1584 (N_1584,In_343,In_136);
nor U1585 (N_1585,In_432,In_444);
nor U1586 (N_1586,In_406,In_674);
nand U1587 (N_1587,In_58,In_630);
or U1588 (N_1588,In_736,In_646);
or U1589 (N_1589,In_344,In_41);
nand U1590 (N_1590,In_342,In_676);
or U1591 (N_1591,In_91,In_246);
and U1592 (N_1592,In_40,In_604);
nor U1593 (N_1593,In_608,In_128);
nand U1594 (N_1594,In_474,In_345);
or U1595 (N_1595,In_360,In_476);
nand U1596 (N_1596,In_75,In_303);
nand U1597 (N_1597,In_133,In_168);
nand U1598 (N_1598,In_288,In_445);
or U1599 (N_1599,In_398,In_644);
or U1600 (N_1600,In_144,In_115);
and U1601 (N_1601,In_442,In_425);
nand U1602 (N_1602,In_737,In_291);
nand U1603 (N_1603,In_33,In_682);
nor U1604 (N_1604,In_444,In_89);
and U1605 (N_1605,In_287,In_230);
nand U1606 (N_1606,In_514,In_171);
and U1607 (N_1607,In_158,In_39);
nand U1608 (N_1608,In_661,In_657);
or U1609 (N_1609,In_448,In_176);
nand U1610 (N_1610,In_171,In_561);
or U1611 (N_1611,In_416,In_304);
or U1612 (N_1612,In_144,In_367);
nand U1613 (N_1613,In_430,In_0);
or U1614 (N_1614,In_707,In_668);
nor U1615 (N_1615,In_506,In_99);
or U1616 (N_1616,In_116,In_78);
nand U1617 (N_1617,In_201,In_478);
and U1618 (N_1618,In_727,In_153);
nor U1619 (N_1619,In_372,In_718);
or U1620 (N_1620,In_153,In_543);
nor U1621 (N_1621,In_656,In_340);
or U1622 (N_1622,In_702,In_707);
or U1623 (N_1623,In_367,In_323);
nor U1624 (N_1624,In_520,In_663);
nor U1625 (N_1625,In_457,In_573);
nor U1626 (N_1626,In_468,In_239);
or U1627 (N_1627,In_684,In_261);
nor U1628 (N_1628,In_85,In_218);
nand U1629 (N_1629,In_546,In_242);
nand U1630 (N_1630,In_707,In_138);
nor U1631 (N_1631,In_538,In_459);
or U1632 (N_1632,In_372,In_378);
nor U1633 (N_1633,In_718,In_69);
nand U1634 (N_1634,In_257,In_500);
and U1635 (N_1635,In_152,In_74);
nor U1636 (N_1636,In_239,In_357);
and U1637 (N_1637,In_36,In_142);
nand U1638 (N_1638,In_241,In_353);
and U1639 (N_1639,In_714,In_264);
nand U1640 (N_1640,In_651,In_553);
nand U1641 (N_1641,In_94,In_393);
nor U1642 (N_1642,In_561,In_748);
nor U1643 (N_1643,In_32,In_457);
nor U1644 (N_1644,In_306,In_697);
nand U1645 (N_1645,In_72,In_172);
or U1646 (N_1646,In_7,In_8);
or U1647 (N_1647,In_170,In_340);
or U1648 (N_1648,In_282,In_127);
nand U1649 (N_1649,In_605,In_308);
or U1650 (N_1650,In_500,In_38);
or U1651 (N_1651,In_443,In_703);
nand U1652 (N_1652,In_545,In_330);
nor U1653 (N_1653,In_401,In_635);
or U1654 (N_1654,In_522,In_313);
nand U1655 (N_1655,In_321,In_293);
nor U1656 (N_1656,In_159,In_223);
nor U1657 (N_1657,In_527,In_389);
or U1658 (N_1658,In_633,In_90);
nand U1659 (N_1659,In_702,In_81);
or U1660 (N_1660,In_198,In_665);
or U1661 (N_1661,In_358,In_61);
nor U1662 (N_1662,In_399,In_552);
nand U1663 (N_1663,In_472,In_571);
and U1664 (N_1664,In_335,In_689);
and U1665 (N_1665,In_614,In_565);
and U1666 (N_1666,In_446,In_23);
nand U1667 (N_1667,In_150,In_602);
or U1668 (N_1668,In_482,In_65);
and U1669 (N_1669,In_322,In_645);
or U1670 (N_1670,In_273,In_409);
nor U1671 (N_1671,In_212,In_482);
and U1672 (N_1672,In_459,In_528);
nand U1673 (N_1673,In_500,In_610);
and U1674 (N_1674,In_346,In_85);
nand U1675 (N_1675,In_138,In_240);
xor U1676 (N_1676,In_548,In_605);
or U1677 (N_1677,In_178,In_63);
nor U1678 (N_1678,In_448,In_156);
and U1679 (N_1679,In_610,In_209);
and U1680 (N_1680,In_305,In_466);
or U1681 (N_1681,In_717,In_9);
or U1682 (N_1682,In_334,In_220);
or U1683 (N_1683,In_461,In_142);
nor U1684 (N_1684,In_31,In_611);
nand U1685 (N_1685,In_153,In_49);
nand U1686 (N_1686,In_664,In_731);
nor U1687 (N_1687,In_474,In_600);
nand U1688 (N_1688,In_298,In_580);
and U1689 (N_1689,In_469,In_387);
nor U1690 (N_1690,In_372,In_251);
and U1691 (N_1691,In_730,In_9);
or U1692 (N_1692,In_294,In_360);
or U1693 (N_1693,In_373,In_106);
nor U1694 (N_1694,In_35,In_59);
nand U1695 (N_1695,In_280,In_191);
xnor U1696 (N_1696,In_53,In_2);
nor U1697 (N_1697,In_101,In_47);
nor U1698 (N_1698,In_106,In_356);
nor U1699 (N_1699,In_419,In_537);
or U1700 (N_1700,In_172,In_59);
or U1701 (N_1701,In_210,In_429);
nand U1702 (N_1702,In_320,In_248);
nor U1703 (N_1703,In_100,In_431);
nand U1704 (N_1704,In_528,In_345);
and U1705 (N_1705,In_512,In_2);
or U1706 (N_1706,In_178,In_525);
nor U1707 (N_1707,In_403,In_33);
nor U1708 (N_1708,In_745,In_340);
and U1709 (N_1709,In_739,In_610);
nand U1710 (N_1710,In_164,In_351);
or U1711 (N_1711,In_351,In_150);
and U1712 (N_1712,In_287,In_494);
nand U1713 (N_1713,In_332,In_359);
nand U1714 (N_1714,In_268,In_152);
and U1715 (N_1715,In_560,In_706);
nor U1716 (N_1716,In_223,In_509);
nor U1717 (N_1717,In_670,In_493);
or U1718 (N_1718,In_469,In_65);
nor U1719 (N_1719,In_404,In_249);
and U1720 (N_1720,In_325,In_407);
nand U1721 (N_1721,In_81,In_696);
or U1722 (N_1722,In_663,In_352);
nand U1723 (N_1723,In_275,In_429);
and U1724 (N_1724,In_190,In_77);
xnor U1725 (N_1725,In_478,In_695);
nand U1726 (N_1726,In_506,In_202);
nand U1727 (N_1727,In_517,In_95);
or U1728 (N_1728,In_148,In_236);
or U1729 (N_1729,In_23,In_451);
or U1730 (N_1730,In_21,In_379);
or U1731 (N_1731,In_497,In_717);
or U1732 (N_1732,In_693,In_363);
and U1733 (N_1733,In_78,In_335);
nor U1734 (N_1734,In_308,In_523);
nor U1735 (N_1735,In_227,In_94);
and U1736 (N_1736,In_633,In_12);
nor U1737 (N_1737,In_532,In_264);
nand U1738 (N_1738,In_659,In_463);
and U1739 (N_1739,In_337,In_18);
or U1740 (N_1740,In_520,In_379);
or U1741 (N_1741,In_678,In_245);
or U1742 (N_1742,In_359,In_220);
nor U1743 (N_1743,In_526,In_229);
nor U1744 (N_1744,In_612,In_156);
nand U1745 (N_1745,In_619,In_419);
nor U1746 (N_1746,In_133,In_260);
and U1747 (N_1747,In_704,In_684);
or U1748 (N_1748,In_245,In_2);
nand U1749 (N_1749,In_653,In_674);
nand U1750 (N_1750,In_473,In_731);
and U1751 (N_1751,In_414,In_170);
nand U1752 (N_1752,In_197,In_453);
nor U1753 (N_1753,In_443,In_422);
or U1754 (N_1754,In_710,In_417);
nor U1755 (N_1755,In_539,In_267);
or U1756 (N_1756,In_130,In_34);
nand U1757 (N_1757,In_654,In_347);
nor U1758 (N_1758,In_19,In_116);
nor U1759 (N_1759,In_723,In_420);
nor U1760 (N_1760,In_21,In_498);
or U1761 (N_1761,In_100,In_438);
xor U1762 (N_1762,In_719,In_215);
or U1763 (N_1763,In_232,In_571);
and U1764 (N_1764,In_6,In_180);
nor U1765 (N_1765,In_651,In_695);
nand U1766 (N_1766,In_14,In_293);
nor U1767 (N_1767,In_9,In_643);
and U1768 (N_1768,In_128,In_233);
and U1769 (N_1769,In_749,In_599);
or U1770 (N_1770,In_602,In_574);
or U1771 (N_1771,In_256,In_291);
nand U1772 (N_1772,In_294,In_737);
and U1773 (N_1773,In_336,In_416);
and U1774 (N_1774,In_453,In_527);
xnor U1775 (N_1775,In_508,In_25);
nor U1776 (N_1776,In_655,In_328);
nor U1777 (N_1777,In_470,In_135);
nand U1778 (N_1778,In_414,In_686);
nand U1779 (N_1779,In_443,In_623);
and U1780 (N_1780,In_64,In_246);
nand U1781 (N_1781,In_246,In_380);
nand U1782 (N_1782,In_733,In_741);
or U1783 (N_1783,In_656,In_499);
nor U1784 (N_1784,In_408,In_181);
nor U1785 (N_1785,In_401,In_522);
nor U1786 (N_1786,In_189,In_381);
nand U1787 (N_1787,In_262,In_290);
and U1788 (N_1788,In_37,In_593);
nand U1789 (N_1789,In_527,In_565);
nand U1790 (N_1790,In_658,In_445);
nand U1791 (N_1791,In_201,In_191);
or U1792 (N_1792,In_89,In_703);
or U1793 (N_1793,In_523,In_132);
or U1794 (N_1794,In_646,In_559);
nor U1795 (N_1795,In_101,In_299);
nand U1796 (N_1796,In_240,In_144);
and U1797 (N_1797,In_493,In_288);
or U1798 (N_1798,In_638,In_506);
nand U1799 (N_1799,In_137,In_108);
and U1800 (N_1800,In_11,In_748);
nor U1801 (N_1801,In_385,In_107);
nand U1802 (N_1802,In_208,In_97);
nand U1803 (N_1803,In_424,In_399);
nor U1804 (N_1804,In_153,In_650);
nor U1805 (N_1805,In_192,In_740);
nand U1806 (N_1806,In_274,In_367);
and U1807 (N_1807,In_30,In_193);
nor U1808 (N_1808,In_337,In_331);
nor U1809 (N_1809,In_406,In_489);
nand U1810 (N_1810,In_47,In_62);
or U1811 (N_1811,In_630,In_289);
nor U1812 (N_1812,In_9,In_86);
nor U1813 (N_1813,In_482,In_3);
nand U1814 (N_1814,In_726,In_65);
nor U1815 (N_1815,In_661,In_706);
or U1816 (N_1816,In_572,In_71);
or U1817 (N_1817,In_91,In_667);
or U1818 (N_1818,In_225,In_363);
nor U1819 (N_1819,In_249,In_525);
nand U1820 (N_1820,In_97,In_626);
nand U1821 (N_1821,In_566,In_225);
or U1822 (N_1822,In_640,In_357);
nor U1823 (N_1823,In_263,In_370);
nor U1824 (N_1824,In_448,In_254);
or U1825 (N_1825,In_156,In_570);
nor U1826 (N_1826,In_225,In_84);
and U1827 (N_1827,In_273,In_693);
or U1828 (N_1828,In_361,In_707);
or U1829 (N_1829,In_645,In_439);
nor U1830 (N_1830,In_65,In_348);
nand U1831 (N_1831,In_651,In_392);
or U1832 (N_1832,In_478,In_592);
nor U1833 (N_1833,In_657,In_359);
nor U1834 (N_1834,In_503,In_390);
or U1835 (N_1835,In_738,In_504);
nand U1836 (N_1836,In_84,In_38);
and U1837 (N_1837,In_283,In_558);
nand U1838 (N_1838,In_487,In_147);
and U1839 (N_1839,In_278,In_629);
or U1840 (N_1840,In_54,In_175);
nor U1841 (N_1841,In_324,In_460);
nor U1842 (N_1842,In_424,In_224);
nor U1843 (N_1843,In_713,In_742);
and U1844 (N_1844,In_186,In_517);
xor U1845 (N_1845,In_395,In_576);
nand U1846 (N_1846,In_141,In_665);
or U1847 (N_1847,In_337,In_694);
or U1848 (N_1848,In_615,In_416);
nand U1849 (N_1849,In_28,In_413);
or U1850 (N_1850,In_100,In_339);
nand U1851 (N_1851,In_7,In_274);
nor U1852 (N_1852,In_574,In_327);
and U1853 (N_1853,In_586,In_318);
nand U1854 (N_1854,In_8,In_319);
or U1855 (N_1855,In_317,In_298);
nor U1856 (N_1856,In_470,In_198);
or U1857 (N_1857,In_739,In_384);
or U1858 (N_1858,In_225,In_139);
nand U1859 (N_1859,In_530,In_141);
and U1860 (N_1860,In_421,In_546);
nand U1861 (N_1861,In_267,In_278);
nor U1862 (N_1862,In_669,In_378);
and U1863 (N_1863,In_554,In_436);
nand U1864 (N_1864,In_410,In_432);
nor U1865 (N_1865,In_627,In_633);
nor U1866 (N_1866,In_2,In_183);
and U1867 (N_1867,In_713,In_440);
nor U1868 (N_1868,In_114,In_279);
or U1869 (N_1869,In_275,In_457);
nor U1870 (N_1870,In_82,In_574);
or U1871 (N_1871,In_729,In_686);
nor U1872 (N_1872,In_182,In_741);
nand U1873 (N_1873,In_525,In_698);
and U1874 (N_1874,In_654,In_319);
and U1875 (N_1875,In_506,In_378);
nor U1876 (N_1876,In_102,In_181);
nor U1877 (N_1877,In_606,In_300);
nor U1878 (N_1878,In_360,In_686);
nand U1879 (N_1879,In_66,In_236);
nor U1880 (N_1880,In_443,In_223);
nand U1881 (N_1881,In_688,In_705);
nand U1882 (N_1882,In_102,In_580);
nor U1883 (N_1883,In_574,In_383);
or U1884 (N_1884,In_520,In_25);
nand U1885 (N_1885,In_617,In_739);
and U1886 (N_1886,In_497,In_307);
nand U1887 (N_1887,In_62,In_13);
nand U1888 (N_1888,In_498,In_414);
nand U1889 (N_1889,In_732,In_603);
xor U1890 (N_1890,In_670,In_36);
nand U1891 (N_1891,In_242,In_97);
nor U1892 (N_1892,In_454,In_472);
or U1893 (N_1893,In_715,In_506);
and U1894 (N_1894,In_171,In_225);
and U1895 (N_1895,In_330,In_327);
nand U1896 (N_1896,In_640,In_534);
nor U1897 (N_1897,In_525,In_216);
nor U1898 (N_1898,In_140,In_146);
and U1899 (N_1899,In_744,In_640);
and U1900 (N_1900,In_229,In_61);
or U1901 (N_1901,In_104,In_322);
or U1902 (N_1902,In_731,In_307);
nor U1903 (N_1903,In_371,In_542);
nand U1904 (N_1904,In_97,In_213);
or U1905 (N_1905,In_500,In_520);
nor U1906 (N_1906,In_140,In_636);
nand U1907 (N_1907,In_142,In_163);
and U1908 (N_1908,In_221,In_459);
or U1909 (N_1909,In_593,In_638);
or U1910 (N_1910,In_567,In_23);
nor U1911 (N_1911,In_305,In_49);
or U1912 (N_1912,In_496,In_305);
or U1913 (N_1913,In_700,In_577);
nor U1914 (N_1914,In_227,In_132);
and U1915 (N_1915,In_245,In_285);
or U1916 (N_1916,In_594,In_593);
and U1917 (N_1917,In_552,In_158);
nand U1918 (N_1918,In_20,In_54);
nor U1919 (N_1919,In_479,In_717);
nor U1920 (N_1920,In_267,In_429);
nand U1921 (N_1921,In_546,In_160);
nand U1922 (N_1922,In_250,In_167);
or U1923 (N_1923,In_424,In_578);
and U1924 (N_1924,In_734,In_674);
and U1925 (N_1925,In_14,In_404);
nand U1926 (N_1926,In_20,In_46);
and U1927 (N_1927,In_48,In_364);
nand U1928 (N_1928,In_131,In_27);
nand U1929 (N_1929,In_490,In_416);
or U1930 (N_1930,In_606,In_196);
and U1931 (N_1931,In_634,In_166);
nand U1932 (N_1932,In_294,In_219);
nor U1933 (N_1933,In_640,In_629);
nor U1934 (N_1934,In_198,In_120);
nand U1935 (N_1935,In_212,In_233);
and U1936 (N_1936,In_182,In_129);
or U1937 (N_1937,In_113,In_643);
xor U1938 (N_1938,In_184,In_467);
and U1939 (N_1939,In_461,In_481);
nor U1940 (N_1940,In_388,In_181);
and U1941 (N_1941,In_659,In_33);
or U1942 (N_1942,In_392,In_419);
and U1943 (N_1943,In_118,In_194);
nand U1944 (N_1944,In_352,In_489);
and U1945 (N_1945,In_61,In_620);
or U1946 (N_1946,In_378,In_241);
and U1947 (N_1947,In_116,In_556);
nand U1948 (N_1948,In_98,In_7);
and U1949 (N_1949,In_399,In_147);
and U1950 (N_1950,In_447,In_115);
nand U1951 (N_1951,In_682,In_542);
and U1952 (N_1952,In_699,In_708);
or U1953 (N_1953,In_559,In_198);
nand U1954 (N_1954,In_275,In_528);
or U1955 (N_1955,In_313,In_0);
nand U1956 (N_1956,In_307,In_670);
nand U1957 (N_1957,In_427,In_584);
or U1958 (N_1958,In_253,In_356);
and U1959 (N_1959,In_546,In_615);
and U1960 (N_1960,In_386,In_201);
nor U1961 (N_1961,In_432,In_95);
and U1962 (N_1962,In_683,In_633);
or U1963 (N_1963,In_614,In_349);
nor U1964 (N_1964,In_265,In_687);
nand U1965 (N_1965,In_291,In_109);
and U1966 (N_1966,In_120,In_277);
nor U1967 (N_1967,In_25,In_304);
and U1968 (N_1968,In_48,In_537);
nor U1969 (N_1969,In_345,In_479);
and U1970 (N_1970,In_21,In_679);
nand U1971 (N_1971,In_585,In_62);
and U1972 (N_1972,In_433,In_51);
or U1973 (N_1973,In_571,In_594);
or U1974 (N_1974,In_57,In_404);
nor U1975 (N_1975,In_230,In_297);
or U1976 (N_1976,In_574,In_37);
nand U1977 (N_1977,In_352,In_747);
nor U1978 (N_1978,In_258,In_100);
nand U1979 (N_1979,In_159,In_157);
and U1980 (N_1980,In_722,In_234);
nor U1981 (N_1981,In_618,In_401);
and U1982 (N_1982,In_556,In_467);
or U1983 (N_1983,In_748,In_608);
or U1984 (N_1984,In_477,In_690);
nor U1985 (N_1985,In_540,In_671);
and U1986 (N_1986,In_262,In_170);
or U1987 (N_1987,In_7,In_715);
nor U1988 (N_1988,In_556,In_544);
or U1989 (N_1989,In_186,In_438);
nand U1990 (N_1990,In_31,In_271);
or U1991 (N_1991,In_585,In_56);
or U1992 (N_1992,In_663,In_444);
nor U1993 (N_1993,In_21,In_682);
and U1994 (N_1994,In_567,In_198);
nand U1995 (N_1995,In_606,In_52);
nand U1996 (N_1996,In_235,In_517);
nor U1997 (N_1997,In_640,In_122);
nor U1998 (N_1998,In_592,In_686);
nor U1999 (N_1999,In_325,In_507);
nor U2000 (N_2000,In_53,In_108);
nor U2001 (N_2001,In_37,In_421);
or U2002 (N_2002,In_150,In_248);
nand U2003 (N_2003,In_370,In_21);
nand U2004 (N_2004,In_107,In_34);
or U2005 (N_2005,In_286,In_705);
and U2006 (N_2006,In_145,In_371);
or U2007 (N_2007,In_93,In_283);
or U2008 (N_2008,In_293,In_198);
nand U2009 (N_2009,In_265,In_730);
nand U2010 (N_2010,In_586,In_296);
and U2011 (N_2011,In_89,In_522);
and U2012 (N_2012,In_454,In_548);
or U2013 (N_2013,In_597,In_728);
or U2014 (N_2014,In_604,In_269);
nand U2015 (N_2015,In_383,In_632);
nand U2016 (N_2016,In_687,In_663);
or U2017 (N_2017,In_4,In_327);
nand U2018 (N_2018,In_660,In_126);
nor U2019 (N_2019,In_150,In_704);
or U2020 (N_2020,In_672,In_322);
or U2021 (N_2021,In_726,In_532);
or U2022 (N_2022,In_223,In_455);
and U2023 (N_2023,In_571,In_312);
nand U2024 (N_2024,In_580,In_228);
or U2025 (N_2025,In_69,In_466);
nand U2026 (N_2026,In_612,In_336);
nor U2027 (N_2027,In_170,In_696);
or U2028 (N_2028,In_226,In_81);
nor U2029 (N_2029,In_405,In_630);
nand U2030 (N_2030,In_540,In_295);
and U2031 (N_2031,In_738,In_277);
or U2032 (N_2032,In_347,In_458);
nor U2033 (N_2033,In_717,In_365);
and U2034 (N_2034,In_283,In_75);
and U2035 (N_2035,In_694,In_644);
and U2036 (N_2036,In_72,In_537);
or U2037 (N_2037,In_93,In_659);
or U2038 (N_2038,In_123,In_463);
nand U2039 (N_2039,In_65,In_213);
or U2040 (N_2040,In_261,In_29);
nor U2041 (N_2041,In_575,In_659);
and U2042 (N_2042,In_277,In_114);
nor U2043 (N_2043,In_686,In_212);
or U2044 (N_2044,In_123,In_281);
and U2045 (N_2045,In_455,In_586);
and U2046 (N_2046,In_106,In_321);
or U2047 (N_2047,In_59,In_597);
and U2048 (N_2048,In_80,In_324);
nand U2049 (N_2049,In_665,In_748);
nand U2050 (N_2050,In_20,In_542);
and U2051 (N_2051,In_646,In_267);
and U2052 (N_2052,In_362,In_277);
nand U2053 (N_2053,In_656,In_134);
and U2054 (N_2054,In_52,In_353);
or U2055 (N_2055,In_720,In_692);
and U2056 (N_2056,In_484,In_726);
and U2057 (N_2057,In_20,In_16);
and U2058 (N_2058,In_227,In_394);
and U2059 (N_2059,In_66,In_530);
nor U2060 (N_2060,In_213,In_423);
or U2061 (N_2061,In_546,In_476);
and U2062 (N_2062,In_604,In_309);
nor U2063 (N_2063,In_454,In_414);
and U2064 (N_2064,In_21,In_444);
xnor U2065 (N_2065,In_58,In_438);
nand U2066 (N_2066,In_677,In_640);
nor U2067 (N_2067,In_183,In_360);
or U2068 (N_2068,In_49,In_184);
nor U2069 (N_2069,In_395,In_730);
and U2070 (N_2070,In_149,In_704);
or U2071 (N_2071,In_57,In_618);
nor U2072 (N_2072,In_57,In_43);
or U2073 (N_2073,In_145,In_699);
nand U2074 (N_2074,In_82,In_561);
and U2075 (N_2075,In_567,In_177);
or U2076 (N_2076,In_493,In_465);
and U2077 (N_2077,In_570,In_507);
nor U2078 (N_2078,In_489,In_619);
or U2079 (N_2079,In_611,In_339);
and U2080 (N_2080,In_519,In_130);
nor U2081 (N_2081,In_218,In_157);
or U2082 (N_2082,In_334,In_337);
nand U2083 (N_2083,In_405,In_591);
nor U2084 (N_2084,In_627,In_569);
nor U2085 (N_2085,In_125,In_75);
nand U2086 (N_2086,In_66,In_493);
nand U2087 (N_2087,In_589,In_326);
or U2088 (N_2088,In_118,In_381);
and U2089 (N_2089,In_629,In_198);
nand U2090 (N_2090,In_388,In_473);
or U2091 (N_2091,In_68,In_141);
and U2092 (N_2092,In_736,In_271);
nand U2093 (N_2093,In_393,In_330);
nand U2094 (N_2094,In_108,In_139);
nor U2095 (N_2095,In_567,In_46);
or U2096 (N_2096,In_512,In_459);
nand U2097 (N_2097,In_442,In_55);
nor U2098 (N_2098,In_418,In_358);
and U2099 (N_2099,In_618,In_660);
nand U2100 (N_2100,In_19,In_607);
or U2101 (N_2101,In_383,In_382);
or U2102 (N_2102,In_216,In_501);
and U2103 (N_2103,In_436,In_26);
nand U2104 (N_2104,In_385,In_624);
or U2105 (N_2105,In_374,In_92);
and U2106 (N_2106,In_744,In_474);
nor U2107 (N_2107,In_313,In_20);
nand U2108 (N_2108,In_73,In_443);
nand U2109 (N_2109,In_241,In_635);
and U2110 (N_2110,In_339,In_465);
xor U2111 (N_2111,In_259,In_467);
or U2112 (N_2112,In_624,In_726);
nand U2113 (N_2113,In_257,In_511);
nand U2114 (N_2114,In_220,In_619);
or U2115 (N_2115,In_738,In_92);
or U2116 (N_2116,In_582,In_525);
nand U2117 (N_2117,In_112,In_543);
and U2118 (N_2118,In_496,In_37);
nor U2119 (N_2119,In_673,In_165);
or U2120 (N_2120,In_516,In_463);
or U2121 (N_2121,In_186,In_346);
or U2122 (N_2122,In_173,In_695);
nor U2123 (N_2123,In_589,In_500);
and U2124 (N_2124,In_235,In_584);
or U2125 (N_2125,In_446,In_526);
nor U2126 (N_2126,In_521,In_35);
nand U2127 (N_2127,In_466,In_518);
or U2128 (N_2128,In_396,In_698);
nor U2129 (N_2129,In_528,In_282);
or U2130 (N_2130,In_440,In_495);
nand U2131 (N_2131,In_492,In_291);
nand U2132 (N_2132,In_395,In_482);
and U2133 (N_2133,In_733,In_24);
nor U2134 (N_2134,In_640,In_390);
and U2135 (N_2135,In_280,In_165);
or U2136 (N_2136,In_161,In_177);
or U2137 (N_2137,In_649,In_461);
nor U2138 (N_2138,In_650,In_633);
nand U2139 (N_2139,In_367,In_503);
nor U2140 (N_2140,In_593,In_540);
or U2141 (N_2141,In_306,In_555);
or U2142 (N_2142,In_302,In_351);
nor U2143 (N_2143,In_688,In_87);
and U2144 (N_2144,In_273,In_593);
or U2145 (N_2145,In_598,In_470);
or U2146 (N_2146,In_561,In_36);
nor U2147 (N_2147,In_451,In_294);
nor U2148 (N_2148,In_656,In_273);
or U2149 (N_2149,In_629,In_235);
or U2150 (N_2150,In_741,In_247);
and U2151 (N_2151,In_317,In_3);
nor U2152 (N_2152,In_478,In_444);
nand U2153 (N_2153,In_95,In_158);
nor U2154 (N_2154,In_151,In_139);
and U2155 (N_2155,In_276,In_618);
nor U2156 (N_2156,In_667,In_549);
nand U2157 (N_2157,In_3,In_343);
nor U2158 (N_2158,In_219,In_344);
or U2159 (N_2159,In_570,In_9);
nor U2160 (N_2160,In_409,In_665);
nand U2161 (N_2161,In_174,In_189);
or U2162 (N_2162,In_78,In_485);
and U2163 (N_2163,In_62,In_389);
or U2164 (N_2164,In_298,In_182);
and U2165 (N_2165,In_574,In_241);
nand U2166 (N_2166,In_163,In_46);
nor U2167 (N_2167,In_113,In_186);
nor U2168 (N_2168,In_283,In_444);
nor U2169 (N_2169,In_2,In_715);
nor U2170 (N_2170,In_303,In_624);
or U2171 (N_2171,In_675,In_743);
and U2172 (N_2172,In_612,In_379);
nor U2173 (N_2173,In_634,In_188);
nand U2174 (N_2174,In_170,In_473);
nor U2175 (N_2175,In_128,In_683);
nor U2176 (N_2176,In_580,In_629);
and U2177 (N_2177,In_432,In_303);
and U2178 (N_2178,In_511,In_501);
nand U2179 (N_2179,In_184,In_650);
nor U2180 (N_2180,In_672,In_245);
nor U2181 (N_2181,In_622,In_492);
nor U2182 (N_2182,In_115,In_381);
nand U2183 (N_2183,In_539,In_492);
nand U2184 (N_2184,In_631,In_439);
nand U2185 (N_2185,In_497,In_146);
nand U2186 (N_2186,In_301,In_489);
and U2187 (N_2187,In_323,In_233);
or U2188 (N_2188,In_352,In_407);
or U2189 (N_2189,In_479,In_462);
or U2190 (N_2190,In_77,In_514);
nand U2191 (N_2191,In_517,In_513);
and U2192 (N_2192,In_116,In_315);
and U2193 (N_2193,In_354,In_76);
nor U2194 (N_2194,In_321,In_652);
nor U2195 (N_2195,In_393,In_601);
or U2196 (N_2196,In_681,In_248);
and U2197 (N_2197,In_249,In_403);
and U2198 (N_2198,In_486,In_110);
nand U2199 (N_2199,In_335,In_103);
nand U2200 (N_2200,In_39,In_306);
nor U2201 (N_2201,In_212,In_256);
or U2202 (N_2202,In_545,In_289);
and U2203 (N_2203,In_280,In_197);
and U2204 (N_2204,In_223,In_65);
and U2205 (N_2205,In_264,In_390);
nand U2206 (N_2206,In_475,In_176);
or U2207 (N_2207,In_564,In_486);
or U2208 (N_2208,In_378,In_170);
nor U2209 (N_2209,In_23,In_128);
or U2210 (N_2210,In_1,In_481);
nor U2211 (N_2211,In_12,In_92);
or U2212 (N_2212,In_211,In_291);
nand U2213 (N_2213,In_363,In_39);
or U2214 (N_2214,In_82,In_596);
nor U2215 (N_2215,In_747,In_590);
nand U2216 (N_2216,In_275,In_706);
nand U2217 (N_2217,In_52,In_584);
nor U2218 (N_2218,In_616,In_656);
nor U2219 (N_2219,In_600,In_583);
and U2220 (N_2220,In_374,In_524);
nor U2221 (N_2221,In_371,In_534);
nand U2222 (N_2222,In_740,In_221);
nand U2223 (N_2223,In_8,In_738);
and U2224 (N_2224,In_321,In_219);
or U2225 (N_2225,In_115,In_181);
and U2226 (N_2226,In_128,In_466);
or U2227 (N_2227,In_727,In_81);
nand U2228 (N_2228,In_655,In_721);
nor U2229 (N_2229,In_365,In_320);
or U2230 (N_2230,In_357,In_211);
nand U2231 (N_2231,In_251,In_59);
nor U2232 (N_2232,In_61,In_604);
nand U2233 (N_2233,In_573,In_148);
xor U2234 (N_2234,In_282,In_229);
nand U2235 (N_2235,In_240,In_206);
and U2236 (N_2236,In_91,In_403);
and U2237 (N_2237,In_472,In_618);
or U2238 (N_2238,In_177,In_167);
nor U2239 (N_2239,In_143,In_652);
or U2240 (N_2240,In_413,In_150);
nand U2241 (N_2241,In_369,In_403);
or U2242 (N_2242,In_591,In_64);
xnor U2243 (N_2243,In_700,In_528);
and U2244 (N_2244,In_289,In_371);
nor U2245 (N_2245,In_574,In_471);
nor U2246 (N_2246,In_13,In_659);
nand U2247 (N_2247,In_366,In_97);
nand U2248 (N_2248,In_481,In_168);
and U2249 (N_2249,In_478,In_619);
nand U2250 (N_2250,In_442,In_294);
nor U2251 (N_2251,In_611,In_596);
nand U2252 (N_2252,In_518,In_743);
or U2253 (N_2253,In_254,In_517);
nand U2254 (N_2254,In_88,In_80);
nand U2255 (N_2255,In_145,In_258);
xor U2256 (N_2256,In_9,In_187);
and U2257 (N_2257,In_128,In_415);
nand U2258 (N_2258,In_125,In_674);
and U2259 (N_2259,In_247,In_208);
nand U2260 (N_2260,In_215,In_164);
or U2261 (N_2261,In_526,In_215);
nand U2262 (N_2262,In_628,In_55);
and U2263 (N_2263,In_38,In_386);
and U2264 (N_2264,In_36,In_32);
nand U2265 (N_2265,In_745,In_43);
and U2266 (N_2266,In_209,In_590);
or U2267 (N_2267,In_44,In_284);
nor U2268 (N_2268,In_718,In_155);
and U2269 (N_2269,In_720,In_1);
nand U2270 (N_2270,In_401,In_345);
nand U2271 (N_2271,In_377,In_255);
nor U2272 (N_2272,In_352,In_563);
nand U2273 (N_2273,In_333,In_86);
nor U2274 (N_2274,In_380,In_630);
or U2275 (N_2275,In_294,In_175);
nand U2276 (N_2276,In_520,In_43);
nand U2277 (N_2277,In_306,In_625);
and U2278 (N_2278,In_741,In_320);
nand U2279 (N_2279,In_69,In_320);
and U2280 (N_2280,In_210,In_380);
or U2281 (N_2281,In_637,In_573);
nor U2282 (N_2282,In_133,In_30);
and U2283 (N_2283,In_191,In_268);
or U2284 (N_2284,In_437,In_592);
or U2285 (N_2285,In_288,In_170);
or U2286 (N_2286,In_361,In_694);
nand U2287 (N_2287,In_529,In_293);
and U2288 (N_2288,In_123,In_140);
nand U2289 (N_2289,In_557,In_223);
and U2290 (N_2290,In_212,In_569);
and U2291 (N_2291,In_430,In_706);
and U2292 (N_2292,In_303,In_151);
nand U2293 (N_2293,In_466,In_309);
or U2294 (N_2294,In_548,In_91);
or U2295 (N_2295,In_333,In_565);
nor U2296 (N_2296,In_464,In_438);
nand U2297 (N_2297,In_573,In_737);
or U2298 (N_2298,In_383,In_54);
or U2299 (N_2299,In_451,In_544);
nor U2300 (N_2300,In_582,In_237);
nand U2301 (N_2301,In_293,In_328);
or U2302 (N_2302,In_65,In_720);
nand U2303 (N_2303,In_476,In_390);
nor U2304 (N_2304,In_158,In_184);
nor U2305 (N_2305,In_314,In_632);
or U2306 (N_2306,In_414,In_387);
nor U2307 (N_2307,In_478,In_446);
or U2308 (N_2308,In_178,In_563);
nand U2309 (N_2309,In_101,In_408);
and U2310 (N_2310,In_517,In_130);
nor U2311 (N_2311,In_546,In_708);
or U2312 (N_2312,In_391,In_440);
or U2313 (N_2313,In_139,In_221);
nor U2314 (N_2314,In_118,In_173);
nor U2315 (N_2315,In_510,In_551);
and U2316 (N_2316,In_163,In_108);
and U2317 (N_2317,In_181,In_28);
or U2318 (N_2318,In_345,In_690);
nor U2319 (N_2319,In_21,In_72);
nor U2320 (N_2320,In_559,In_564);
and U2321 (N_2321,In_603,In_316);
nor U2322 (N_2322,In_615,In_685);
and U2323 (N_2323,In_134,In_24);
or U2324 (N_2324,In_656,In_590);
or U2325 (N_2325,In_569,In_308);
nor U2326 (N_2326,In_385,In_464);
or U2327 (N_2327,In_576,In_150);
or U2328 (N_2328,In_341,In_44);
nand U2329 (N_2329,In_39,In_356);
nor U2330 (N_2330,In_361,In_455);
nor U2331 (N_2331,In_14,In_345);
and U2332 (N_2332,In_588,In_173);
and U2333 (N_2333,In_587,In_73);
nand U2334 (N_2334,In_451,In_701);
or U2335 (N_2335,In_396,In_611);
nand U2336 (N_2336,In_163,In_44);
nand U2337 (N_2337,In_81,In_227);
or U2338 (N_2338,In_706,In_227);
nor U2339 (N_2339,In_62,In_473);
and U2340 (N_2340,In_461,In_165);
and U2341 (N_2341,In_536,In_677);
nor U2342 (N_2342,In_446,In_13);
nor U2343 (N_2343,In_683,In_576);
and U2344 (N_2344,In_574,In_623);
nand U2345 (N_2345,In_317,In_372);
nand U2346 (N_2346,In_604,In_351);
and U2347 (N_2347,In_571,In_592);
and U2348 (N_2348,In_742,In_709);
nand U2349 (N_2349,In_92,In_147);
nor U2350 (N_2350,In_152,In_439);
nor U2351 (N_2351,In_661,In_27);
nand U2352 (N_2352,In_572,In_520);
nor U2353 (N_2353,In_101,In_748);
and U2354 (N_2354,In_504,In_164);
or U2355 (N_2355,In_18,In_562);
nand U2356 (N_2356,In_501,In_127);
nand U2357 (N_2357,In_150,In_451);
nor U2358 (N_2358,In_203,In_221);
nor U2359 (N_2359,In_414,In_116);
and U2360 (N_2360,In_386,In_649);
nand U2361 (N_2361,In_69,In_236);
and U2362 (N_2362,In_474,In_266);
and U2363 (N_2363,In_580,In_20);
or U2364 (N_2364,In_132,In_564);
or U2365 (N_2365,In_551,In_177);
or U2366 (N_2366,In_50,In_476);
or U2367 (N_2367,In_171,In_583);
nand U2368 (N_2368,In_687,In_604);
or U2369 (N_2369,In_470,In_524);
nand U2370 (N_2370,In_53,In_654);
nand U2371 (N_2371,In_431,In_335);
nor U2372 (N_2372,In_168,In_737);
or U2373 (N_2373,In_584,In_161);
nand U2374 (N_2374,In_615,In_39);
nand U2375 (N_2375,In_33,In_599);
and U2376 (N_2376,In_409,In_525);
nand U2377 (N_2377,In_513,In_390);
nand U2378 (N_2378,In_187,In_545);
or U2379 (N_2379,In_489,In_379);
nor U2380 (N_2380,In_699,In_9);
and U2381 (N_2381,In_326,In_445);
nand U2382 (N_2382,In_210,In_109);
or U2383 (N_2383,In_402,In_441);
nor U2384 (N_2384,In_325,In_298);
nor U2385 (N_2385,In_656,In_272);
nor U2386 (N_2386,In_88,In_134);
nor U2387 (N_2387,In_95,In_90);
or U2388 (N_2388,In_28,In_564);
or U2389 (N_2389,In_138,In_639);
nor U2390 (N_2390,In_345,In_104);
and U2391 (N_2391,In_9,In_373);
or U2392 (N_2392,In_539,In_259);
nand U2393 (N_2393,In_660,In_120);
nor U2394 (N_2394,In_647,In_575);
nand U2395 (N_2395,In_430,In_122);
or U2396 (N_2396,In_66,In_95);
or U2397 (N_2397,In_180,In_718);
or U2398 (N_2398,In_421,In_189);
and U2399 (N_2399,In_60,In_183);
nand U2400 (N_2400,In_566,In_569);
and U2401 (N_2401,In_12,In_66);
and U2402 (N_2402,In_215,In_439);
nand U2403 (N_2403,In_149,In_559);
and U2404 (N_2404,In_282,In_81);
nor U2405 (N_2405,In_229,In_344);
nor U2406 (N_2406,In_495,In_481);
or U2407 (N_2407,In_285,In_382);
and U2408 (N_2408,In_583,In_221);
or U2409 (N_2409,In_390,In_327);
nor U2410 (N_2410,In_692,In_534);
and U2411 (N_2411,In_720,In_309);
nor U2412 (N_2412,In_556,In_335);
nand U2413 (N_2413,In_740,In_614);
or U2414 (N_2414,In_456,In_294);
nor U2415 (N_2415,In_128,In_274);
or U2416 (N_2416,In_304,In_541);
nor U2417 (N_2417,In_641,In_540);
nor U2418 (N_2418,In_667,In_70);
or U2419 (N_2419,In_536,In_707);
nor U2420 (N_2420,In_713,In_503);
and U2421 (N_2421,In_341,In_607);
nand U2422 (N_2422,In_53,In_650);
nand U2423 (N_2423,In_121,In_47);
or U2424 (N_2424,In_321,In_126);
nand U2425 (N_2425,In_216,In_464);
or U2426 (N_2426,In_316,In_524);
nand U2427 (N_2427,In_87,In_527);
or U2428 (N_2428,In_482,In_438);
nand U2429 (N_2429,In_218,In_365);
and U2430 (N_2430,In_548,In_566);
nor U2431 (N_2431,In_167,In_620);
xor U2432 (N_2432,In_542,In_202);
or U2433 (N_2433,In_324,In_365);
or U2434 (N_2434,In_144,In_342);
or U2435 (N_2435,In_279,In_156);
nand U2436 (N_2436,In_726,In_490);
nand U2437 (N_2437,In_233,In_207);
and U2438 (N_2438,In_484,In_644);
nor U2439 (N_2439,In_703,In_446);
xnor U2440 (N_2440,In_90,In_201);
nand U2441 (N_2441,In_87,In_472);
or U2442 (N_2442,In_341,In_333);
or U2443 (N_2443,In_733,In_504);
nand U2444 (N_2444,In_671,In_422);
or U2445 (N_2445,In_666,In_321);
nor U2446 (N_2446,In_14,In_174);
nand U2447 (N_2447,In_611,In_587);
nand U2448 (N_2448,In_632,In_27);
nand U2449 (N_2449,In_124,In_493);
nand U2450 (N_2450,In_146,In_201);
nand U2451 (N_2451,In_192,In_586);
nor U2452 (N_2452,In_398,In_28);
nor U2453 (N_2453,In_299,In_421);
nand U2454 (N_2454,In_48,In_419);
nor U2455 (N_2455,In_12,In_69);
nor U2456 (N_2456,In_525,In_348);
or U2457 (N_2457,In_128,In_326);
nor U2458 (N_2458,In_678,In_218);
nand U2459 (N_2459,In_712,In_653);
nand U2460 (N_2460,In_383,In_10);
and U2461 (N_2461,In_676,In_243);
and U2462 (N_2462,In_116,In_425);
nor U2463 (N_2463,In_602,In_748);
nor U2464 (N_2464,In_674,In_749);
and U2465 (N_2465,In_170,In_679);
nand U2466 (N_2466,In_475,In_515);
and U2467 (N_2467,In_499,In_79);
or U2468 (N_2468,In_522,In_707);
nor U2469 (N_2469,In_704,In_207);
and U2470 (N_2470,In_544,In_434);
nor U2471 (N_2471,In_248,In_141);
and U2472 (N_2472,In_362,In_630);
or U2473 (N_2473,In_551,In_236);
or U2474 (N_2474,In_249,In_437);
xor U2475 (N_2475,In_442,In_54);
nand U2476 (N_2476,In_196,In_695);
nor U2477 (N_2477,In_289,In_697);
nand U2478 (N_2478,In_709,In_537);
nor U2479 (N_2479,In_482,In_648);
or U2480 (N_2480,In_430,In_625);
and U2481 (N_2481,In_282,In_338);
nor U2482 (N_2482,In_405,In_396);
nand U2483 (N_2483,In_452,In_316);
or U2484 (N_2484,In_293,In_74);
and U2485 (N_2485,In_739,In_277);
and U2486 (N_2486,In_157,In_705);
or U2487 (N_2487,In_338,In_181);
nor U2488 (N_2488,In_709,In_632);
nand U2489 (N_2489,In_148,In_313);
nand U2490 (N_2490,In_366,In_623);
nor U2491 (N_2491,In_693,In_31);
and U2492 (N_2492,In_115,In_650);
and U2493 (N_2493,In_716,In_123);
nor U2494 (N_2494,In_283,In_159);
or U2495 (N_2495,In_164,In_318);
nor U2496 (N_2496,In_746,In_263);
or U2497 (N_2497,In_551,In_295);
and U2498 (N_2498,In_271,In_507);
or U2499 (N_2499,In_391,In_718);
or U2500 (N_2500,N_2454,N_2285);
or U2501 (N_2501,N_527,N_1867);
and U2502 (N_2502,N_2365,N_156);
nor U2503 (N_2503,N_2460,N_166);
or U2504 (N_2504,N_2081,N_1734);
or U2505 (N_2505,N_1958,N_1011);
nor U2506 (N_2506,N_994,N_1648);
nand U2507 (N_2507,N_217,N_1082);
xnor U2508 (N_2508,N_332,N_1807);
or U2509 (N_2509,N_2304,N_1111);
nor U2510 (N_2510,N_1293,N_719);
nand U2511 (N_2511,N_292,N_1411);
nand U2512 (N_2512,N_2261,N_2348);
nor U2513 (N_2513,N_1093,N_259);
nand U2514 (N_2514,N_1189,N_1072);
nor U2515 (N_2515,N_1501,N_1);
and U2516 (N_2516,N_1581,N_790);
and U2517 (N_2517,N_91,N_1757);
or U2518 (N_2518,N_1039,N_782);
nand U2519 (N_2519,N_2376,N_10);
or U2520 (N_2520,N_1809,N_2406);
nor U2521 (N_2521,N_557,N_767);
nand U2522 (N_2522,N_184,N_729);
or U2523 (N_2523,N_670,N_1570);
nor U2524 (N_2524,N_1963,N_243);
nor U2525 (N_2525,N_1362,N_569);
nand U2526 (N_2526,N_1972,N_1413);
and U2527 (N_2527,N_1657,N_1296);
nor U2528 (N_2528,N_1669,N_662);
nor U2529 (N_2529,N_1140,N_515);
nand U2530 (N_2530,N_815,N_741);
nor U2531 (N_2531,N_21,N_82);
nand U2532 (N_2532,N_2145,N_412);
or U2533 (N_2533,N_1000,N_1044);
nor U2534 (N_2534,N_1046,N_1444);
or U2535 (N_2535,N_1801,N_483);
or U2536 (N_2536,N_2154,N_11);
nor U2537 (N_2537,N_1965,N_1373);
or U2538 (N_2538,N_297,N_1136);
and U2539 (N_2539,N_299,N_2186);
nor U2540 (N_2540,N_2357,N_2192);
nand U2541 (N_2541,N_2216,N_567);
nand U2542 (N_2542,N_1765,N_737);
or U2543 (N_2543,N_857,N_824);
nand U2544 (N_2544,N_227,N_971);
nor U2545 (N_2545,N_566,N_471);
nor U2546 (N_2546,N_2046,N_117);
nor U2547 (N_2547,N_360,N_923);
and U2548 (N_2548,N_890,N_214);
or U2549 (N_2549,N_749,N_1130);
nor U2550 (N_2550,N_2243,N_387);
or U2551 (N_2551,N_2245,N_2003);
or U2552 (N_2552,N_1675,N_1896);
and U2553 (N_2553,N_850,N_552);
nand U2554 (N_2554,N_1421,N_2188);
nand U2555 (N_2555,N_1107,N_931);
and U2556 (N_2556,N_2112,N_1608);
nor U2557 (N_2557,N_1232,N_592);
nand U2558 (N_2558,N_1528,N_2409);
nand U2559 (N_2559,N_880,N_1694);
or U2560 (N_2560,N_634,N_1917);
and U2561 (N_2561,N_1493,N_549);
and U2562 (N_2562,N_2461,N_2108);
nand U2563 (N_2563,N_2339,N_530);
nand U2564 (N_2564,N_1885,N_1695);
nand U2565 (N_2565,N_1230,N_1805);
nand U2566 (N_2566,N_1062,N_2280);
nor U2567 (N_2567,N_950,N_734);
or U2568 (N_2568,N_173,N_1558);
or U2569 (N_2569,N_1895,N_1204);
and U2570 (N_2570,N_591,N_1886);
nor U2571 (N_2571,N_798,N_2318);
nor U2572 (N_2572,N_980,N_2143);
or U2573 (N_2573,N_377,N_153);
xor U2574 (N_2574,N_1873,N_2259);
and U2575 (N_2575,N_98,N_2041);
and U2576 (N_2576,N_2465,N_498);
xor U2577 (N_2577,N_150,N_1894);
nand U2578 (N_2578,N_1970,N_2250);
nor U2579 (N_2579,N_1193,N_619);
and U2580 (N_2580,N_2341,N_1168);
nand U2581 (N_2581,N_2386,N_1556);
nor U2582 (N_2582,N_608,N_2097);
nand U2583 (N_2583,N_1430,N_460);
nand U2584 (N_2584,N_1290,N_1016);
nand U2585 (N_2585,N_305,N_240);
and U2586 (N_2586,N_462,N_1384);
nor U2587 (N_2587,N_1103,N_758);
nor U2588 (N_2588,N_45,N_255);
or U2589 (N_2589,N_1153,N_241);
and U2590 (N_2590,N_943,N_625);
nand U2591 (N_2591,N_945,N_1147);
nand U2592 (N_2592,N_2126,N_2313);
or U2593 (N_2593,N_553,N_492);
and U2594 (N_2594,N_2347,N_126);
nand U2595 (N_2595,N_842,N_2099);
nor U2596 (N_2596,N_1739,N_1235);
or U2597 (N_2597,N_2173,N_1018);
or U2598 (N_2598,N_773,N_159);
and U2599 (N_2599,N_1334,N_446);
nor U2600 (N_2600,N_1910,N_1364);
or U2601 (N_2601,N_143,N_274);
nand U2602 (N_2602,N_1745,N_2423);
nand U2603 (N_2603,N_1706,N_92);
and U2604 (N_2604,N_2019,N_67);
nor U2605 (N_2605,N_2310,N_2262);
or U2606 (N_2606,N_2105,N_746);
or U2607 (N_2607,N_167,N_939);
or U2608 (N_2608,N_638,N_1877);
nor U2609 (N_2609,N_1670,N_723);
nand U2610 (N_2610,N_1918,N_1735);
or U2611 (N_2611,N_2148,N_1664);
nand U2612 (N_2612,N_1741,N_65);
and U2613 (N_2613,N_147,N_72);
nor U2614 (N_2614,N_2078,N_148);
and U2615 (N_2615,N_1248,N_2276);
or U2616 (N_2616,N_328,N_1174);
nand U2617 (N_2617,N_742,N_1366);
nor U2618 (N_2618,N_1118,N_655);
nand U2619 (N_2619,N_928,N_1627);
nor U2620 (N_2620,N_2147,N_1157);
and U2621 (N_2621,N_171,N_1665);
and U2622 (N_2622,N_2361,N_195);
or U2623 (N_2623,N_1621,N_1844);
or U2624 (N_2624,N_1418,N_2151);
nor U2625 (N_2625,N_2211,N_2416);
nand U2626 (N_2626,N_36,N_87);
or U2627 (N_2627,N_1119,N_2462);
nand U2628 (N_2628,N_1388,N_2054);
and U2629 (N_2629,N_1173,N_2433);
nor U2630 (N_2630,N_1547,N_104);
nor U2631 (N_2631,N_432,N_1791);
or U2632 (N_2632,N_812,N_334);
nor U2633 (N_2633,N_1236,N_142);
and U2634 (N_2634,N_541,N_315);
nand U2635 (N_2635,N_1860,N_122);
nor U2636 (N_2636,N_1078,N_189);
nand U2637 (N_2637,N_1994,N_2420);
and U2638 (N_2638,N_1061,N_290);
and U2639 (N_2639,N_312,N_1169);
nand U2640 (N_2640,N_2152,N_2484);
nor U2641 (N_2641,N_2066,N_2084);
or U2642 (N_2642,N_2297,N_37);
or U2643 (N_2643,N_694,N_1412);
and U2644 (N_2644,N_338,N_1969);
and U2645 (N_2645,N_60,N_579);
nand U2646 (N_2646,N_69,N_791);
and U2647 (N_2647,N_1112,N_2056);
and U2648 (N_2648,N_2294,N_1081);
and U2649 (N_2649,N_56,N_1749);
or U2650 (N_2650,N_1470,N_411);
nor U2651 (N_2651,N_2422,N_2174);
nand U2652 (N_2652,N_1442,N_771);
nor U2653 (N_2653,N_2346,N_947);
and U2654 (N_2654,N_852,N_1800);
nor U2655 (N_2655,N_1568,N_897);
nand U2656 (N_2656,N_847,N_985);
or U2657 (N_2657,N_1224,N_2375);
and U2658 (N_2658,N_2384,N_960);
and U2659 (N_2659,N_1312,N_846);
nand U2660 (N_2660,N_1035,N_250);
and U2661 (N_2661,N_1121,N_477);
nor U2662 (N_2662,N_2263,N_1602);
or U2663 (N_2663,N_891,N_2236);
and U2664 (N_2664,N_2426,N_1100);
and U2665 (N_2665,N_1966,N_337);
and U2666 (N_2666,N_2475,N_494);
nor U2667 (N_2667,N_649,N_293);
or U2668 (N_2668,N_1409,N_2010);
and U2669 (N_2669,N_1606,N_1604);
nor U2670 (N_2670,N_9,N_1616);
nor U2671 (N_2671,N_1273,N_970);
nor U2672 (N_2672,N_2176,N_2324);
or U2673 (N_2673,N_2150,N_1689);
or U2674 (N_2674,N_520,N_1848);
nor U2675 (N_2675,N_1510,N_1831);
and U2676 (N_2676,N_1787,N_1600);
nor U2677 (N_2677,N_2129,N_978);
and U2678 (N_2678,N_1998,N_1923);
nand U2679 (N_2679,N_796,N_1681);
or U2680 (N_2680,N_1251,N_1359);
nand U2681 (N_2681,N_2366,N_705);
and U2682 (N_2682,N_487,N_626);
nand U2683 (N_2683,N_1518,N_1474);
nor U2684 (N_2684,N_457,N_849);
and U2685 (N_2685,N_1012,N_1048);
nand U2686 (N_2686,N_306,N_1197);
nand U2687 (N_2687,N_28,N_1261);
nor U2688 (N_2688,N_2074,N_2079);
or U2689 (N_2689,N_1387,N_309);
nor U2690 (N_2690,N_405,N_743);
nand U2691 (N_2691,N_1552,N_2328);
or U2692 (N_2692,N_63,N_1904);
and U2693 (N_2693,N_883,N_197);
nor U2694 (N_2694,N_631,N_598);
nand U2695 (N_2695,N_1098,N_33);
xnor U2696 (N_2696,N_1661,N_1819);
nor U2697 (N_2697,N_1068,N_2215);
and U2698 (N_2698,N_2298,N_1794);
nor U2699 (N_2699,N_208,N_2269);
nand U2700 (N_2700,N_2302,N_588);
or U2701 (N_2701,N_268,N_1983);
or U2702 (N_2702,N_1882,N_859);
and U2703 (N_2703,N_2479,N_1386);
or U2704 (N_2704,N_2073,N_1357);
nand U2705 (N_2705,N_1677,N_1530);
or U2706 (N_2706,N_445,N_822);
nor U2707 (N_2707,N_1915,N_1924);
nand U2708 (N_2708,N_1069,N_327);
nor U2709 (N_2709,N_523,N_1815);
nand U2710 (N_2710,N_1065,N_775);
or U2711 (N_2711,N_2193,N_1203);
or U2712 (N_2712,N_593,N_1881);
or U2713 (N_2713,N_2400,N_1651);
nor U2714 (N_2714,N_1973,N_681);
and U2715 (N_2715,N_49,N_401);
nand U2716 (N_2716,N_999,N_1370);
or U2717 (N_2717,N_2213,N_1252);
nor U2718 (N_2718,N_1215,N_1128);
and U2719 (N_2719,N_1188,N_2160);
nand U2720 (N_2720,N_2277,N_394);
nand U2721 (N_2721,N_1300,N_1986);
nor U2722 (N_2722,N_2155,N_1862);
nand U2723 (N_2723,N_1846,N_1243);
or U2724 (N_2724,N_270,N_2195);
and U2725 (N_2725,N_839,N_34);
nor U2726 (N_2726,N_1700,N_835);
nand U2727 (N_2727,N_1453,N_232);
nand U2728 (N_2728,N_100,N_1978);
or U2729 (N_2729,N_2453,N_1186);
nand U2730 (N_2730,N_1467,N_428);
and U2731 (N_2731,N_2352,N_584);
nor U2732 (N_2732,N_1671,N_144);
or U2733 (N_2733,N_281,N_777);
nand U2734 (N_2734,N_5,N_478);
and U2735 (N_2735,N_1821,N_1541);
nand U2736 (N_2736,N_121,N_1397);
nor U2737 (N_2737,N_1223,N_2325);
nor U2738 (N_2738,N_689,N_525);
and U2739 (N_2739,N_19,N_1875);
and U2740 (N_2740,N_1521,N_786);
nand U2741 (N_2741,N_2349,N_864);
and U2742 (N_2742,N_213,N_2229);
or U2743 (N_2743,N_785,N_2024);
nand U2744 (N_2744,N_1812,N_418);
and U2745 (N_2745,N_2271,N_886);
or U2746 (N_2746,N_1240,N_2440);
and U2747 (N_2747,N_559,N_2093);
nand U2748 (N_2748,N_1287,N_212);
nor U2749 (N_2749,N_888,N_695);
nor U2750 (N_2750,N_853,N_2106);
nand U2751 (N_2751,N_2225,N_533);
nand U2752 (N_2752,N_2191,N_1902);
nand U2753 (N_2753,N_909,N_797);
nand U2754 (N_2754,N_399,N_180);
and U2755 (N_2755,N_2025,N_112);
or U2756 (N_2756,N_1133,N_802);
or U2757 (N_2757,N_651,N_384);
nand U2758 (N_2758,N_823,N_644);
and U2759 (N_2759,N_501,N_1201);
nor U2760 (N_2760,N_339,N_2090);
or U2761 (N_2761,N_1916,N_479);
and U2762 (N_2762,N_1043,N_1869);
nand U2763 (N_2763,N_1380,N_365);
nor U2764 (N_2764,N_187,N_1624);
nor U2765 (N_2765,N_1355,N_613);
nor U2766 (N_2766,N_903,N_621);
nand U2767 (N_2767,N_969,N_1485);
nor U2768 (N_2768,N_1054,N_226);
and U2769 (N_2769,N_2335,N_1676);
nor U2770 (N_2770,N_1907,N_1714);
nor U2771 (N_2771,N_2134,N_2094);
nor U2772 (N_2772,N_490,N_560);
nand U2773 (N_2773,N_977,N_1784);
and U2774 (N_2774,N_996,N_683);
or U2775 (N_2775,N_2464,N_1826);
and U2776 (N_2776,N_2166,N_635);
and U2777 (N_2777,N_753,N_336);
nand U2778 (N_2778,N_1152,N_2083);
nand U2779 (N_2779,N_673,N_1631);
and U2780 (N_2780,N_562,N_510);
or U2781 (N_2781,N_661,N_1834);
nand U2782 (N_2782,N_807,N_415);
nand U2783 (N_2783,N_2385,N_1320);
nand U2784 (N_2784,N_2477,N_1257);
nand U2785 (N_2785,N_1900,N_1277);
and U2786 (N_2786,N_1170,N_787);
nor U2787 (N_2787,N_587,N_1284);
and U2788 (N_2788,N_1336,N_1414);
or U2789 (N_2789,N_89,N_1160);
and U2790 (N_2790,N_979,N_1613);
nand U2791 (N_2791,N_2063,N_1959);
or U2792 (N_2792,N_1259,N_1849);
nand U2793 (N_2793,N_1233,N_423);
nand U2794 (N_2794,N_717,N_1306);
and U2795 (N_2795,N_160,N_764);
nand U2796 (N_2796,N_335,N_910);
and U2797 (N_2797,N_2457,N_825);
or U2798 (N_2798,N_2340,N_1859);
nor U2799 (N_2799,N_276,N_1225);
nor U2800 (N_2800,N_1864,N_1066);
or U2801 (N_2801,N_42,N_1806);
nor U2802 (N_2802,N_732,N_1297);
and U2803 (N_2803,N_434,N_652);
or U2804 (N_2804,N_2431,N_654);
nor U2805 (N_2805,N_194,N_1574);
or U2806 (N_2806,N_2042,N_351);
nor U2807 (N_2807,N_145,N_2473);
and U2808 (N_2808,N_547,N_1632);
nand U2809 (N_2809,N_1008,N_2203);
and U2810 (N_2810,N_192,N_905);
or U2811 (N_2811,N_2,N_1148);
or U2812 (N_2812,N_107,N_865);
or U2813 (N_2813,N_304,N_1544);
nor U2814 (N_2814,N_1449,N_1294);
nor U2815 (N_2815,N_946,N_2059);
and U2816 (N_2816,N_813,N_2432);
and U2817 (N_2817,N_2159,N_2396);
nor U2818 (N_2818,N_2255,N_2264);
and U2819 (N_2819,N_216,N_2164);
nor U2820 (N_2820,N_368,N_275);
nor U2821 (N_2821,N_313,N_200);
and U2822 (N_2822,N_2028,N_1206);
nand U2823 (N_2823,N_2436,N_877);
nor U2824 (N_2824,N_2049,N_783);
or U2825 (N_2825,N_1537,N_778);
or U2826 (N_2826,N_794,N_1578);
nor U2827 (N_2827,N_311,N_1723);
and U2828 (N_2828,N_288,N_738);
and U2829 (N_2829,N_185,N_1949);
nand U2830 (N_2830,N_2095,N_990);
nand U2831 (N_2831,N_934,N_314);
or U2832 (N_2832,N_1356,N_781);
nand U2833 (N_2833,N_1995,N_1597);
and U2834 (N_2834,N_1381,N_2096);
or U2835 (N_2835,N_1692,N_325);
nor U2836 (N_2836,N_1617,N_74);
and U2837 (N_2837,N_1484,N_1721);
nor U2838 (N_2838,N_589,N_927);
and U2839 (N_2839,N_1351,N_2233);
and U2840 (N_2840,N_953,N_417);
nand U2841 (N_2841,N_1562,N_516);
or U2842 (N_2842,N_1473,N_1222);
and U2843 (N_2843,N_2198,N_389);
nor U2844 (N_2844,N_1956,N_1780);
nor U2845 (N_2845,N_899,N_1813);
or U2846 (N_2846,N_324,N_1643);
and U2847 (N_2847,N_2362,N_426);
or U2848 (N_2848,N_1595,N_289);
and U2849 (N_2849,N_2419,N_2004);
and U2850 (N_2850,N_642,N_172);
and U2851 (N_2851,N_2201,N_1984);
nor U2852 (N_2852,N_2169,N_935);
and U2853 (N_2853,N_1579,N_1253);
nor U2854 (N_2854,N_951,N_341);
and U2855 (N_2855,N_1580,N_2135);
and U2856 (N_2856,N_1181,N_1064);
nor U2857 (N_2857,N_131,N_1938);
and U2858 (N_2858,N_271,N_982);
or U2859 (N_2859,N_1854,N_1847);
nand U2860 (N_2860,N_1154,N_2012);
or U2861 (N_2861,N_1271,N_948);
nor U2862 (N_2862,N_1930,N_278);
or U2863 (N_2863,N_273,N_1256);
nor U2864 (N_2864,N_885,N_2451);
nor U2865 (N_2865,N_1023,N_1625);
and U2866 (N_2866,N_1802,N_941);
or U2867 (N_2867,N_287,N_508);
and U2868 (N_2868,N_1029,N_2387);
nand U2869 (N_2869,N_114,N_7);
and U2870 (N_2870,N_1063,N_1731);
nand U2871 (N_2871,N_47,N_572);
nand U2872 (N_2872,N_410,N_1853);
nor U2873 (N_2873,N_1109,N_601);
nand U2874 (N_2874,N_1454,N_1102);
nand U2875 (N_2875,N_998,N_537);
nor U2876 (N_2876,N_519,N_1987);
or U2877 (N_2877,N_2102,N_920);
nand U2878 (N_2878,N_132,N_1520);
xnor U2879 (N_2879,N_382,N_1716);
xor U2880 (N_2880,N_406,N_2364);
or U2881 (N_2881,N_1006,N_2301);
nand U2882 (N_2882,N_2249,N_2140);
and U2883 (N_2883,N_1754,N_643);
nand U2884 (N_2884,N_427,N_52);
and U2885 (N_2885,N_369,N_1099);
nand U2886 (N_2886,N_1056,N_2359);
and U2887 (N_2887,N_2478,N_1175);
nand U2888 (N_2888,N_1177,N_663);
nand U2889 (N_2889,N_115,N_1990);
and U2890 (N_2890,N_162,N_2246);
or U2891 (N_2891,N_1495,N_1360);
and U2892 (N_2892,N_514,N_603);
nand U2893 (N_2893,N_1673,N_1946);
nand U2894 (N_2894,N_140,N_1941);
and U2895 (N_2895,N_1639,N_1298);
or U2896 (N_2896,N_660,N_2332);
nand U2897 (N_2897,N_1605,N_1811);
nand U2898 (N_2898,N_1220,N_364);
or U2899 (N_2899,N_2446,N_668);
or U2900 (N_2900,N_2343,N_1561);
and U2901 (N_2901,N_1909,N_2070);
and U2902 (N_2902,N_2214,N_1863);
nand U2903 (N_2903,N_628,N_656);
and U2904 (N_2904,N_1303,N_1115);
and U2905 (N_2905,N_1372,N_757);
nand U2906 (N_2906,N_680,N_1030);
or U2907 (N_2907,N_205,N_1905);
and U2908 (N_2908,N_1034,N_1289);
nor U2909 (N_2909,N_2077,N_0);
or U2910 (N_2910,N_1553,N_930);
and U2911 (N_2911,N_1926,N_1650);
nand U2912 (N_2912,N_793,N_321);
and U2913 (N_2913,N_2330,N_455);
and U2914 (N_2914,N_29,N_123);
nand U2915 (N_2915,N_2487,N_473);
and U2916 (N_2916,N_1536,N_2165);
and U2917 (N_2917,N_1378,N_728);
nand U2918 (N_2918,N_395,N_1962);
or U2919 (N_2919,N_354,N_811);
nand U2920 (N_2920,N_357,N_1509);
nand U2921 (N_2921,N_2170,N_263);
nand U2922 (N_2922,N_53,N_1656);
and U2923 (N_2923,N_2020,N_1117);
nor U2924 (N_2924,N_641,N_1855);
and U2925 (N_2925,N_375,N_1382);
and U2926 (N_2926,N_407,N_1090);
or U2927 (N_2927,N_340,N_1105);
xnor U2928 (N_2928,N_1266,N_2064);
nand U2929 (N_2929,N_913,N_2043);
nand U2930 (N_2930,N_983,N_1728);
nor U2931 (N_2931,N_609,N_88);
and U2932 (N_2932,N_1050,N_24);
nand U2933 (N_2933,N_1968,N_1051);
and U2934 (N_2934,N_1891,N_2469);
and U2935 (N_2935,N_1960,N_1055);
nor U2936 (N_2936,N_2336,N_667);
nand U2937 (N_2937,N_687,N_2239);
nand U2938 (N_2938,N_1270,N_1301);
nor U2939 (N_2939,N_1328,N_711);
nor U2940 (N_2940,N_1392,N_2086);
nor U2941 (N_2941,N_1437,N_671);
or U2942 (N_2942,N_1479,N_348);
nor U2943 (N_2943,N_1324,N_186);
or U2944 (N_2944,N_1207,N_1014);
or U2945 (N_2945,N_1316,N_898);
nand U2946 (N_2946,N_1234,N_714);
nand U2947 (N_2947,N_538,N_932);
nand U2948 (N_2948,N_1250,N_23);
and U2949 (N_2949,N_1150,N_1653);
nor U2950 (N_2950,N_2481,N_1868);
or U2951 (N_2951,N_1954,N_1151);
or U2952 (N_2952,N_464,N_1329);
nand U2953 (N_2953,N_1007,N_2380);
nand U2954 (N_2954,N_2013,N_1049);
nor U2955 (N_2955,N_684,N_182);
nor U2956 (N_2956,N_373,N_1337);
nor U2957 (N_2957,N_2224,N_1948);
or U2958 (N_2958,N_469,N_1438);
or U2959 (N_2959,N_1443,N_511);
nand U2960 (N_2960,N_2065,N_1194);
and U2961 (N_2961,N_1679,N_1113);
nand U2962 (N_2962,N_1461,N_678);
and U2963 (N_2963,N_1654,N_247);
or U2964 (N_2964,N_1655,N_1045);
nand U2965 (N_2965,N_349,N_874);
nor U2966 (N_2966,N_959,N_2312);
nand U2967 (N_2967,N_356,N_837);
nor U2968 (N_2968,N_421,N_2207);
and U2969 (N_2969,N_1619,N_2008);
nand U2970 (N_2970,N_1519,N_1892);
or U2971 (N_2971,N_27,N_1040);
and U2972 (N_2972,N_209,N_1139);
or U2973 (N_2973,N_2403,N_1260);
or U2974 (N_2974,N_582,N_699);
nor U2975 (N_2975,N_1319,N_316);
and U2976 (N_2976,N_1401,N_257);
nand U2977 (N_2977,N_1545,N_997);
nor U2978 (N_2978,N_1460,N_2153);
and U2979 (N_2979,N_843,N_1772);
and U2980 (N_2980,N_2300,N_70);
or U2981 (N_2981,N_1718,N_721);
nand U2982 (N_2982,N_1084,N_736);
and U2983 (N_2983,N_1901,N_868);
nor U2984 (N_2984,N_2425,N_2017);
nand U2985 (N_2985,N_1101,N_2394);
nand U2986 (N_2986,N_1943,N_2128);
and U2987 (N_2987,N_2091,N_2226);
and U2988 (N_2988,N_1208,N_1793);
and U2989 (N_2989,N_2044,N_300);
nand U2990 (N_2990,N_733,N_2142);
nor U2991 (N_2991,N_1183,N_1024);
nor U2992 (N_2992,N_2001,N_279);
nor U2993 (N_2993,N_810,N_15);
or U2994 (N_2994,N_25,N_2368);
or U2995 (N_2995,N_2321,N_2061);
and U2996 (N_2996,N_914,N_1612);
and U2997 (N_2997,N_1952,N_2204);
nand U2998 (N_2998,N_575,N_1588);
or U2999 (N_2999,N_1285,N_2303);
nor U3000 (N_3000,N_2466,N_1214);
or U3001 (N_3001,N_1707,N_342);
nand U3002 (N_3002,N_1032,N_302);
or U3003 (N_3003,N_1583,N_1164);
or U3004 (N_3004,N_383,N_294);
nor U3005 (N_3005,N_607,N_392);
nor U3006 (N_3006,N_1264,N_2060);
and U3007 (N_3007,N_1094,N_1999);
and U3008 (N_3008,N_1379,N_1908);
and U3009 (N_3009,N_2130,N_441);
nand U3010 (N_3010,N_1982,N_1587);
nor U3011 (N_3011,N_1988,N_376);
or U3012 (N_3012,N_430,N_1142);
nand U3013 (N_3013,N_1766,N_1638);
and U3014 (N_3014,N_2272,N_1229);
nor U3015 (N_3015,N_989,N_966);
or U3016 (N_3016,N_911,N_14);
nand U3017 (N_3017,N_236,N_1540);
nor U3018 (N_3018,N_1861,N_916);
nor U3019 (N_3019,N_1705,N_747);
nor U3020 (N_3020,N_1709,N_1897);
or U3021 (N_3021,N_249,N_1088);
nand U3022 (N_3022,N_177,N_95);
or U3023 (N_3023,N_2467,N_242);
or U3024 (N_3024,N_789,N_1404);
nor U3025 (N_3025,N_22,N_1196);
and U3026 (N_3026,N_2048,N_1693);
and U3027 (N_3027,N_677,N_2181);
or U3028 (N_3028,N_1845,N_1526);
and U3029 (N_3029,N_1363,N_2463);
and U3030 (N_3030,N_1469,N_1857);
and U3031 (N_3031,N_2278,N_1981);
and U3032 (N_3032,N_539,N_500);
nor U3033 (N_3033,N_679,N_1953);
nand U3034 (N_3034,N_809,N_564);
or U3035 (N_3035,N_915,N_2018);
nand U3036 (N_3036,N_2144,N_1614);
and U3037 (N_3037,N_925,N_1975);
nor U3038 (N_3038,N_2401,N_1126);
nand U3039 (N_3039,N_378,N_1347);
nor U3040 (N_3040,N_2326,N_2038);
xnor U3041 (N_3041,N_1125,N_2444);
nand U3042 (N_3042,N_178,N_895);
or U3043 (N_3043,N_2222,N_438);
nor U3044 (N_3044,N_1365,N_2327);
and U3045 (N_3045,N_1795,N_1827);
or U3046 (N_3046,N_2237,N_470);
and U3047 (N_3047,N_254,N_266);
nand U3048 (N_3048,N_762,N_750);
or U3049 (N_3049,N_230,N_139);
nand U3050 (N_3050,N_1172,N_1647);
and U3051 (N_3051,N_2005,N_151);
nand U3052 (N_3052,N_1083,N_1955);
and U3053 (N_3053,N_1571,N_2219);
nor U3054 (N_3054,N_206,N_1792);
and U3055 (N_3055,N_1920,N_2089);
nor U3056 (N_3056,N_1013,N_2363);
nor U3057 (N_3057,N_924,N_2241);
nor U3058 (N_3058,N_2449,N_957);
nor U3059 (N_3059,N_1808,N_1028);
or U3060 (N_3060,N_1361,N_2293);
and U3061 (N_3061,N_1796,N_727);
or U3062 (N_3062,N_995,N_1017);
nor U3063 (N_3063,N_2316,N_792);
nand U3064 (N_3064,N_2209,N_573);
nor U3065 (N_3065,N_2162,N_1674);
nor U3066 (N_3066,N_77,N_1763);
or U3067 (N_3067,N_18,N_1010);
nor U3068 (N_3068,N_2404,N_1368);
and U3069 (N_3069,N_1097,N_1508);
nor U3070 (N_3070,N_554,N_944);
and U3071 (N_3071,N_179,N_956);
nand U3072 (N_3072,N_2057,N_497);
nand U3073 (N_3073,N_1506,N_2337);
and U3074 (N_3074,N_393,N_1500);
nand U3075 (N_3075,N_2288,N_2485);
nand U3076 (N_3076,N_372,N_1841);
nand U3077 (N_3077,N_648,N_2260);
and U3078 (N_3078,N_2286,N_265);
or U3079 (N_3079,N_988,N_2103);
or U3080 (N_3080,N_2163,N_2405);
nor U3081 (N_3081,N_1037,N_2491);
and U3082 (N_3082,N_964,N_461);
nand U3083 (N_3083,N_2411,N_1748);
or U3084 (N_3084,N_532,N_2323);
or U3085 (N_3085,N_992,N_1344);
nand U3086 (N_3086,N_907,N_900);
or U3087 (N_3087,N_929,N_215);
or U3088 (N_3088,N_618,N_1426);
nor U3089 (N_3089,N_1992,N_2482);
and U3090 (N_3090,N_84,N_1991);
or U3091 (N_3091,N_2266,N_2124);
and U3092 (N_3092,N_1790,N_2415);
and U3093 (N_3093,N_366,N_146);
or U3094 (N_3094,N_1996,N_283);
nor U3095 (N_3095,N_225,N_1543);
nor U3096 (N_3096,N_805,N_522);
and U3097 (N_3097,N_1354,N_467);
and U3098 (N_3098,N_872,N_766);
nor U3099 (N_3099,N_135,N_1529);
and U3100 (N_3100,N_922,N_1993);
nor U3101 (N_3101,N_1464,N_2014);
or U3102 (N_3102,N_2408,N_1838);
nor U3103 (N_3103,N_596,N_420);
nand U3104 (N_3104,N_2468,N_1440);
or U3105 (N_3105,N_1549,N_1132);
nor U3106 (N_3106,N_1209,N_2418);
nor U3107 (N_3107,N_908,N_774);
and U3108 (N_3108,N_1471,N_343);
nand U3109 (N_3109,N_1166,N_1195);
nand U3110 (N_3110,N_647,N_2254);
or U3111 (N_3111,N_119,N_1830);
nand U3112 (N_3112,N_2299,N_1202);
nand U3113 (N_3113,N_1699,N_2398);
or U3114 (N_3114,N_2053,N_2493);
nand U3115 (N_3115,N_1459,N_2251);
nor U3116 (N_3116,N_1925,N_1237);
and U3117 (N_3117,N_277,N_93);
or U3118 (N_3118,N_149,N_1980);
or U3119 (N_3119,N_2305,N_109);
nand U3120 (N_3120,N_1345,N_1199);
or U3121 (N_3121,N_1783,N_2287);
and U3122 (N_3122,N_509,N_1342);
or U3123 (N_3123,N_2062,N_2306);
or U3124 (N_3124,N_1431,N_99);
and U3125 (N_3125,N_1660,N_505);
or U3126 (N_3126,N_1879,N_2334);
nor U3127 (N_3127,N_1021,N_1933);
or U3128 (N_3128,N_1009,N_1513);
xnor U3129 (N_3129,N_202,N_1108);
nor U3130 (N_3130,N_120,N_105);
and U3131 (N_3131,N_840,N_2047);
nor U3132 (N_3132,N_949,N_529);
nor U3133 (N_3133,N_2034,N_50);
nor U3134 (N_3134,N_414,N_484);
nand U3135 (N_3135,N_1001,N_1906);
nor U3136 (N_3136,N_1913,N_1928);
nand U3137 (N_3137,N_1488,N_229);
and U3138 (N_3138,N_40,N_952);
and U3139 (N_3139,N_218,N_1644);
xor U3140 (N_3140,N_912,N_1465);
and U3141 (N_3141,N_544,N_1163);
nand U3142 (N_3142,N_1592,N_2317);
and U3143 (N_3143,N_1546,N_1180);
nor U3144 (N_3144,N_2372,N_1123);
or U3145 (N_3145,N_2499,N_2315);
and U3146 (N_3146,N_2448,N_754);
nand U3147 (N_3147,N_861,N_2413);
or U3148 (N_3148,N_284,N_698);
and U3149 (N_3149,N_355,N_1004);
xnor U3150 (N_3150,N_474,N_513);
and U3151 (N_3151,N_237,N_1523);
nand U3152 (N_3152,N_118,N_380);
nor U3153 (N_3153,N_730,N_1434);
and U3154 (N_3154,N_2441,N_188);
nand U3155 (N_3155,N_1832,N_506);
xor U3156 (N_3156,N_260,N_1590);
xor U3157 (N_3157,N_2345,N_1778);
or U3158 (N_3158,N_739,N_2027);
or U3159 (N_3159,N_2210,N_1607);
and U3160 (N_3160,N_152,N_1522);
or U3161 (N_3161,N_425,N_1810);
or U3162 (N_3162,N_286,N_2109);
or U3163 (N_3163,N_1872,N_2437);
nand U3164 (N_3164,N_2098,N_1652);
nand U3165 (N_3165,N_2421,N_1462);
and U3166 (N_3166,N_2033,N_1307);
or U3167 (N_3167,N_1353,N_940);
nand U3168 (N_3168,N_1358,N_2279);
and U3169 (N_3169,N_106,N_157);
nand U3170 (N_3170,N_1769,N_1335);
nor U3171 (N_3171,N_526,N_561);
nor U3172 (N_3172,N_975,N_1106);
nand U3173 (N_3173,N_2427,N_333);
and U3174 (N_3174,N_1331,N_1268);
nand U3175 (N_3175,N_1515,N_876);
and U3176 (N_3176,N_2189,N_623);
or U3177 (N_3177,N_2068,N_2360);
and U3178 (N_3178,N_1446,N_658);
nor U3179 (N_3179,N_599,N_301);
nand U3180 (N_3180,N_1756,N_1025);
and U3181 (N_3181,N_1369,N_616);
and U3182 (N_3182,N_2227,N_622);
nor U3183 (N_3183,N_543,N_1701);
nor U3184 (N_3184,N_1408,N_258);
and U3185 (N_3185,N_1346,N_2088);
or U3186 (N_3186,N_396,N_884);
nor U3187 (N_3187,N_1489,N_2050);
nand U3188 (N_3188,N_451,N_1416);
or U3189 (N_3189,N_124,N_307);
or U3190 (N_3190,N_855,N_163);
and U3191 (N_3191,N_1075,N_101);
or U3192 (N_3192,N_1087,N_51);
nor U3193 (N_3193,N_204,N_454);
nor U3194 (N_3194,N_1348,N_2447);
nand U3195 (N_3195,N_1280,N_1771);
nand U3196 (N_3196,N_1263,N_1124);
or U3197 (N_3197,N_2497,N_704);
nand U3198 (N_3198,N_2132,N_1478);
nand U3199 (N_3199,N_71,N_2080);
or U3200 (N_3200,N_1406,N_1687);
nor U3201 (N_3201,N_745,N_1599);
nand U3202 (N_3202,N_540,N_1971);
nor U3203 (N_3203,N_1659,N_1314);
nand U3204 (N_3204,N_317,N_605);
or U3205 (N_3205,N_653,N_2494);
or U3206 (N_3206,N_1551,N_708);
nand U3207 (N_3207,N_1569,N_2149);
and U3208 (N_3208,N_1743,N_556);
nand U3209 (N_3209,N_2356,N_1929);
or U3210 (N_3210,N_1542,N_674);
nand U3211 (N_3211,N_385,N_2021);
or U3212 (N_3212,N_1468,N_665);
nand U3213 (N_3213,N_2127,N_765);
and U3214 (N_3214,N_2185,N_235);
nand U3215 (N_3215,N_2072,N_1292);
nor U3216 (N_3216,N_581,N_450);
or U3217 (N_3217,N_1274,N_1742);
and U3218 (N_3218,N_1629,N_326);
nand U3219 (N_3219,N_1496,N_1751);
nor U3220 (N_3220,N_66,N_1730);
nand U3221 (N_3221,N_2388,N_1376);
or U3222 (N_3222,N_893,N_594);
nand U3223 (N_3223,N_986,N_1598);
nor U3224 (N_3224,N_1685,N_1502);
or U3225 (N_3225,N_1927,N_1275);
or U3226 (N_3226,N_1487,N_615);
nand U3227 (N_3227,N_480,N_1759);
and U3228 (N_3228,N_1452,N_1278);
nand U3229 (N_3229,N_756,N_1635);
and U3230 (N_3230,N_1410,N_239);
nor U3231 (N_3231,N_1622,N_2085);
nand U3232 (N_3232,N_2338,N_1903);
or U3233 (N_3233,N_2350,N_1708);
or U3234 (N_3234,N_1403,N_391);
nor U3235 (N_3235,N_322,N_2382);
or U3236 (N_3236,N_475,N_906);
nor U3237 (N_3237,N_1753,N_331);
nand U3238 (N_3238,N_604,N_967);
or U3239 (N_3239,N_1752,N_1114);
and U3240 (N_3240,N_2082,N_1340);
or U3241 (N_3241,N_2353,N_1727);
nor U3242 (N_3242,N_2157,N_234);
and U3243 (N_3243,N_894,N_1283);
and U3244 (N_3244,N_1057,N_1424);
or U3245 (N_3245,N_1429,N_2265);
and U3246 (N_3246,N_489,N_1750);
nand U3247 (N_3247,N_2314,N_2231);
nand U3248 (N_3248,N_1394,N_817);
nand U3249 (N_3249,N_436,N_1603);
nor U3250 (N_3250,N_1936,N_449);
or U3251 (N_3251,N_1947,N_1371);
nor U3252 (N_3252,N_770,N_2307);
and U3253 (N_3253,N_374,N_1441);
or U3254 (N_3254,N_136,N_844);
nand U3255 (N_3255,N_2311,N_1433);
nor U3256 (N_3256,N_921,N_2490);
or U3257 (N_3257,N_1836,N_2414);
nor U3258 (N_3258,N_675,N_1171);
nand U3259 (N_3259,N_1499,N_2417);
nor U3260 (N_3260,N_2399,N_2424);
or U3261 (N_3261,N_1589,N_856);
nor U3262 (N_3262,N_1305,N_1038);
nor U3263 (N_3263,N_2342,N_46);
and U3264 (N_3264,N_1258,N_129);
nor U3265 (N_3265,N_452,N_826);
or U3266 (N_3266,N_1666,N_576);
nand U3267 (N_3267,N_1804,N_419);
and U3268 (N_3268,N_2410,N_1961);
or U3269 (N_3269,N_2367,N_1782);
nor U3270 (N_3270,N_1724,N_2092);
nand U3271 (N_3271,N_1550,N_1490);
nor U3272 (N_3272,N_578,N_1668);
nor U3273 (N_3273,N_1129,N_1702);
and U3274 (N_3274,N_1717,N_2187);
and U3275 (N_3275,N_1737,N_600);
xnor U3276 (N_3276,N_2110,N_1565);
and U3277 (N_3277,N_1833,N_413);
nand U3278 (N_3278,N_2052,N_251);
and U3279 (N_3279,N_918,N_2371);
and U3280 (N_3280,N_1187,N_1554);
and U3281 (N_3281,N_1179,N_1976);
or U3282 (N_3282,N_676,N_851);
or U3283 (N_3283,N_650,N_2498);
and U3284 (N_3284,N_1476,N_2455);
and U3285 (N_3285,N_1400,N_1422);
nand U3286 (N_3286,N_402,N_585);
and U3287 (N_3287,N_433,N_252);
and U3288 (N_3288,N_710,N_2223);
nand U3289 (N_3289,N_201,N_1146);
nor U3290 (N_3290,N_1041,N_38);
nand U3291 (N_3291,N_531,N_690);
or U3292 (N_3292,N_1939,N_1219);
and U3293 (N_3293,N_2267,N_1803);
or U3294 (N_3294,N_353,N_495);
or U3295 (N_3295,N_1074,N_1053);
nand U3296 (N_3296,N_1732,N_1758);
and U3297 (N_3297,N_1633,N_1144);
and U3298 (N_3298,N_1596,N_1740);
and U3299 (N_3299,N_1427,N_1874);
and U3300 (N_3300,N_463,N_712);
nor U3301 (N_3301,N_2218,N_1843);
nor U3302 (N_3302,N_1713,N_32);
and U3303 (N_3303,N_108,N_1110);
nor U3304 (N_3304,N_1858,N_1390);
nand U3305 (N_3305,N_546,N_1711);
and U3306 (N_3306,N_1839,N_691);
and U3307 (N_3307,N_503,N_657);
and U3308 (N_3308,N_1079,N_1878);
or U3309 (N_3309,N_1391,N_308);
or U3310 (N_3310,N_1672,N_1385);
or U3311 (N_3311,N_845,N_808);
and U3312 (N_3312,N_1626,N_1350);
or U3313 (N_3313,N_1310,N_1585);
xnor U3314 (N_3314,N_2087,N_1463);
nand U3315 (N_3315,N_437,N_30);
or U3316 (N_3316,N_2039,N_496);
or U3317 (N_3317,N_2442,N_1407);
or U3318 (N_3318,N_1814,N_2194);
nand U3319 (N_3319,N_58,N_1785);
nor U3320 (N_3320,N_1480,N_1377);
nor U3321 (N_3321,N_1198,N_1774);
and U3322 (N_3322,N_1974,N_361);
or U3323 (N_3323,N_1491,N_863);
nor U3324 (N_3324,N_2196,N_134);
and U3325 (N_3325,N_1582,N_2071);
or U3326 (N_3326,N_1267,N_85);
nand U3327 (N_3327,N_666,N_233);
nand U3328 (N_3328,N_1835,N_1323);
nor U3329 (N_3329,N_2333,N_379);
nand U3330 (N_3330,N_468,N_2274);
and U3331 (N_3331,N_1919,N_1871);
nor U3332 (N_3332,N_1073,N_1033);
nor U3333 (N_3333,N_2055,N_1281);
nand U3334 (N_3334,N_570,N_1884);
or U3335 (N_3335,N_1228,N_211);
nand U3336 (N_3336,N_2331,N_1985);
nor U3337 (N_3337,N_183,N_170);
nor U3338 (N_3338,N_1667,N_748);
nand U3339 (N_3339,N_528,N_203);
or U3340 (N_3340,N_344,N_1182);
and U3341 (N_3341,N_1686,N_1779);
or U3342 (N_3342,N_1497,N_130);
nand U3343 (N_3343,N_238,N_456);
nor U3344 (N_3344,N_493,N_550);
nand U3345 (N_3345,N_2075,N_1077);
and U3346 (N_3346,N_688,N_1269);
nor U3347 (N_3347,N_1089,N_44);
nand U3348 (N_3348,N_2476,N_435);
nor U3349 (N_3349,N_833,N_1483);
nand U3350 (N_3350,N_984,N_1031);
or U3351 (N_3351,N_1591,N_1498);
and U3352 (N_3352,N_1899,N_1797);
or U3353 (N_3353,N_860,N_2197);
and U3354 (N_3354,N_804,N_97);
nor U3355 (N_3355,N_954,N_1192);
nor U3356 (N_3356,N_2480,N_1036);
nand U3357 (N_3357,N_2161,N_466);
nor U3358 (N_3358,N_693,N_2067);
and U3359 (N_3359,N_784,N_1457);
nand U3360 (N_3360,N_267,N_772);
and U3361 (N_3361,N_1451,N_720);
nor U3362 (N_3362,N_1276,N_3);
nor U3363 (N_3363,N_169,N_367);
nand U3364 (N_3364,N_62,N_761);
or U3365 (N_3365,N_1254,N_1680);
nor U3366 (N_3366,N_2016,N_113);
nand U3367 (N_3367,N_1967,N_1052);
or U3368 (N_3368,N_1122,N_1159);
nor U3369 (N_3369,N_974,N_1576);
nor U3370 (N_3370,N_386,N_2496);
and U3371 (N_3371,N_453,N_2177);
or U3372 (N_3372,N_1816,N_16);
nand U3373 (N_3373,N_882,N_534);
and U3374 (N_3374,N_154,N_1524);
and U3375 (N_3375,N_878,N_610);
or U3376 (N_3376,N_1481,N_1116);
nand U3377 (N_3377,N_261,N_1466);
or U3378 (N_3378,N_190,N_2354);
nand U3379 (N_3379,N_827,N_1733);
nand U3380 (N_3380,N_2117,N_858);
nor U3381 (N_3381,N_917,N_2030);
xnor U3382 (N_3382,N_191,N_1231);
and U3383 (N_3383,N_73,N_1279);
nand U3384 (N_3384,N_1213,N_2474);
nor U3385 (N_3385,N_2136,N_2257);
nor U3386 (N_3386,N_697,N_2175);
nand U3387 (N_3387,N_174,N_59);
nor U3388 (N_3388,N_1352,N_424);
nor U3389 (N_3389,N_2045,N_196);
nand U3390 (N_3390,N_352,N_848);
or U3391 (N_3391,N_1047,N_2492);
or U3392 (N_3392,N_2115,N_760);
and U3393 (N_3393,N_2015,N_1876);
and U3394 (N_3394,N_1776,N_889);
or U3395 (N_3395,N_1719,N_219);
nand U3396 (N_3396,N_2146,N_1092);
and U3397 (N_3397,N_2172,N_244);
nor U3398 (N_3398,N_61,N_222);
or U3399 (N_3399,N_2495,N_81);
nor U3400 (N_3400,N_1856,N_2428);
or U3401 (N_3401,N_2370,N_2202);
and U3402 (N_3402,N_485,N_2320);
nor U3403 (N_3403,N_1837,N_871);
nor U3404 (N_3404,N_1134,N_1770);
nand U3405 (N_3405,N_1226,N_1997);
or U3406 (N_3406,N_31,N_2430);
nand U3407 (N_3407,N_2270,N_1768);
nand U3408 (N_3408,N_1914,N_403);
nand U3409 (N_3409,N_1852,N_1889);
and U3410 (N_3410,N_2379,N_1472);
nor U3411 (N_3411,N_1678,N_1822);
or U3412 (N_3412,N_512,N_2358);
nand U3413 (N_3413,N_1249,N_887);
and U3414 (N_3414,N_870,N_595);
or U3415 (N_3415,N_580,N_535);
nand U3416 (N_3416,N_1825,N_1637);
or U3417 (N_3417,N_524,N_981);
and U3418 (N_3418,N_221,N_323);
nand U3419 (N_3419,N_958,N_854);
and U3420 (N_3420,N_1567,N_1559);
nor U3421 (N_3421,N_933,N_1725);
nor U3422 (N_3422,N_1977,N_1851);
nand U3423 (N_3423,N_1746,N_1691);
nor U3424 (N_3424,N_867,N_2439);
nor U3425 (N_3425,N_536,N_1091);
and U3426 (N_3426,N_751,N_488);
and U3427 (N_3427,N_976,N_2412);
and U3428 (N_3428,N_2292,N_2378);
xor U3429 (N_3429,N_2104,N_199);
nor U3430 (N_3430,N_818,N_20);
or U3431 (N_3431,N_165,N_329);
nor U3432 (N_3432,N_1555,N_901);
nor U3433 (N_3433,N_1210,N_398);
nand U3434 (N_3434,N_2006,N_814);
and U3435 (N_3435,N_1773,N_2168);
and U3436 (N_3436,N_245,N_2011);
nand U3437 (N_3437,N_448,N_1247);
nand U3438 (N_3438,N_1615,N_2121);
nor U3439 (N_3439,N_700,N_1636);
nor U3440 (N_3440,N_936,N_2283);
or U3441 (N_3441,N_2248,N_502);
or U3442 (N_3442,N_795,N_1517);
nor U3443 (N_3443,N_2205,N_1238);
and U3444 (N_3444,N_1242,N_1942);
or U3445 (N_3445,N_1447,N_602);
or U3446 (N_3446,N_2051,N_1218);
or U3447 (N_3447,N_1789,N_875);
nor U3448 (N_3448,N_1722,N_1842);
nor U3449 (N_3449,N_2178,N_207);
or U3450 (N_3450,N_879,N_2190);
nand U3451 (N_3451,N_1070,N_1321);
or U3452 (N_3452,N_350,N_716);
or U3453 (N_3453,N_2171,N_2100);
nor U3454 (N_3454,N_1934,N_696);
nor U3455 (N_3455,N_2023,N_111);
or U3456 (N_3456,N_2247,N_2456);
nand U3457 (N_3457,N_722,N_1317);
or U3458 (N_3458,N_1548,N_1343);
nand U3459 (N_3459,N_1145,N_2206);
nand U3460 (N_3460,N_1628,N_1937);
nand U3461 (N_3461,N_1682,N_320);
and U3462 (N_3462,N_836,N_2141);
nand U3463 (N_3463,N_2101,N_388);
nor U3464 (N_3464,N_2167,N_1911);
xnor U3465 (N_3465,N_639,N_2291);
nand U3466 (N_3466,N_1593,N_1456);
or U3467 (N_3467,N_1866,N_2397);
nand U3468 (N_3468,N_1432,N_869);
nand U3469 (N_3469,N_1535,N_1532);
xnor U3470 (N_3470,N_718,N_1200);
nand U3471 (N_3471,N_346,N_2374);
nand U3472 (N_3472,N_1211,N_1720);
or U3473 (N_3473,N_1494,N_1840);
or U3474 (N_3474,N_1747,N_1375);
nor U3475 (N_3475,N_517,N_264);
and U3476 (N_3476,N_1311,N_1155);
or U3477 (N_3477,N_1205,N_1684);
nand U3478 (N_3478,N_2268,N_735);
or U3479 (N_3479,N_2009,N_55);
nand U3480 (N_3480,N_703,N_1295);
nor U3481 (N_3481,N_586,N_499);
or U3482 (N_3482,N_54,N_759);
and U3483 (N_3483,N_955,N_2289);
nor U3484 (N_3484,N_669,N_1601);
and U3485 (N_3485,N_1662,N_347);
nand U3486 (N_3486,N_993,N_1396);
nor U3487 (N_3487,N_2282,N_1663);
nand U3488 (N_3488,N_991,N_1245);
nor U3489 (N_3489,N_518,N_2199);
nor U3490 (N_3490,N_2007,N_624);
nor U3491 (N_3491,N_2000,N_2182);
or U3492 (N_3492,N_1019,N_246);
and U3493 (N_3493,N_1104,N_1533);
nor U3494 (N_3494,N_486,N_545);
or U3495 (N_3495,N_1888,N_779);
and U3496 (N_3496,N_752,N_1272);
and U3497 (N_3497,N_1964,N_319);
and U3498 (N_3498,N_345,N_1244);
nand U3499 (N_3499,N_2122,N_57);
nand U3500 (N_3500,N_2381,N_612);
or U3501 (N_3501,N_1330,N_2238);
nor U3502 (N_3502,N_439,N_1338);
or U3503 (N_3503,N_659,N_2309);
nor U3504 (N_3504,N_1085,N_881);
xnor U3505 (N_3505,N_1255,N_1744);
nor U3506 (N_3506,N_1932,N_731);
and U3507 (N_3507,N_555,N_1922);
nor U3508 (N_3508,N_2434,N_801);
and U3509 (N_3509,N_2351,N_1420);
nand U3510 (N_3510,N_1492,N_431);
or U3511 (N_3511,N_2308,N_1823);
and U3512 (N_3512,N_1393,N_298);
and U3513 (N_3513,N_1349,N_1096);
or U3514 (N_3514,N_1799,N_1308);
nand U3515 (N_3515,N_1060,N_800);
nor U3516 (N_3516,N_35,N_409);
and U3517 (N_3517,N_86,N_713);
nor U3518 (N_3518,N_763,N_1291);
nand U3519 (N_3519,N_2230,N_39);
or U3520 (N_3520,N_1940,N_2450);
nand U3521 (N_3521,N_2452,N_838);
or U3522 (N_3522,N_2138,N_1095);
nand U3523 (N_3523,N_1005,N_1399);
nor U3524 (N_3524,N_458,N_155);
or U3525 (N_3525,N_1658,N_2253);
nor U3526 (N_3526,N_2158,N_829);
and U3527 (N_3527,N_2032,N_2179);
xor U3528 (N_3528,N_1127,N_1436);
nor U3529 (N_3529,N_1696,N_1042);
and U3530 (N_3530,N_1641,N_491);
and U3531 (N_3531,N_2252,N_125);
nor U3532 (N_3532,N_1313,N_2228);
and U3533 (N_3533,N_973,N_740);
nand U3534 (N_3534,N_285,N_1880);
nand U3535 (N_3535,N_632,N_590);
or U3536 (N_3536,N_1594,N_1557);
or U3537 (N_3537,N_1241,N_2107);
nor U3538 (N_3538,N_1630,N_2383);
nand U3539 (N_3539,N_571,N_1820);
nor U3540 (N_3540,N_443,N_2002);
and U3541 (N_3541,N_429,N_1341);
nor U3542 (N_3542,N_2137,N_444);
and U3543 (N_3543,N_1445,N_231);
or U3544 (N_3544,N_709,N_2488);
nor U3545 (N_3545,N_726,N_138);
or U3546 (N_3546,N_1697,N_633);
nand U3547 (N_3547,N_2040,N_2390);
nand U3548 (N_3548,N_390,N_1149);
nand U3549 (N_3549,N_2443,N_2184);
or U3550 (N_3550,N_158,N_937);
or U3551 (N_3551,N_1262,N_542);
nor U3552 (N_3552,N_397,N_2036);
nor U3553 (N_3553,N_1419,N_1318);
xnor U3554 (N_3554,N_701,N_303);
nor U3555 (N_3555,N_702,N_1762);
nor U3556 (N_3556,N_2438,N_862);
nor U3557 (N_3557,N_780,N_210);
nand U3558 (N_3558,N_359,N_2391);
nand U3559 (N_3559,N_558,N_942);
nand U3560 (N_3560,N_2029,N_1538);
nor U3561 (N_3561,N_1246,N_1755);
nor U3562 (N_3562,N_1398,N_2483);
and U3563 (N_3563,N_282,N_2429);
or U3564 (N_3564,N_1764,N_1086);
nor U3565 (N_3565,N_1282,N_362);
nand U3566 (N_3566,N_2118,N_79);
or U3567 (N_3567,N_164,N_1325);
and U3568 (N_3568,N_2133,N_1883);
nand U3569 (N_3569,N_1921,N_2472);
and U3570 (N_3570,N_1649,N_1767);
or U3571 (N_3571,N_43,N_1634);
nand U3572 (N_3572,N_1131,N_1458);
and U3573 (N_3573,N_968,N_1137);
and U3574 (N_3574,N_2212,N_2026);
nand U3575 (N_3575,N_1738,N_1989);
nor U3576 (N_3576,N_1850,N_2131);
and U3577 (N_3577,N_828,N_1002);
nand U3578 (N_3578,N_2373,N_253);
or U3579 (N_3579,N_1216,N_1584);
nor U3580 (N_3580,N_280,N_2273);
nand U3581 (N_3581,N_551,N_2393);
nor U3582 (N_3582,N_269,N_2058);
nand U3583 (N_3583,N_1712,N_318);
and U3584 (N_3584,N_12,N_2119);
nand U3585 (N_3585,N_1435,N_1870);
nand U3586 (N_3586,N_1286,N_892);
nor U3587 (N_3587,N_707,N_645);
nor U3588 (N_3588,N_1950,N_2220);
or U3589 (N_3589,N_820,N_193);
and U3590 (N_3590,N_2295,N_1688);
nand U3591 (N_3591,N_1304,N_26);
nand U3592 (N_3592,N_1315,N_358);
nand U3593 (N_3593,N_2322,N_1945);
nand U3594 (N_3594,N_2113,N_965);
nor U3595 (N_3595,N_2235,N_96);
and U3596 (N_3596,N_629,N_755);
nor U3597 (N_3597,N_583,N_2183);
or U3598 (N_3598,N_819,N_1893);
nor U3599 (N_3599,N_1761,N_776);
and U3600 (N_3600,N_248,N_1566);
and U3601 (N_3601,N_2319,N_481);
or U3602 (N_3602,N_1736,N_1322);
nand U3603 (N_3603,N_1572,N_161);
nand U3604 (N_3604,N_1405,N_1327);
nor U3605 (N_3605,N_834,N_1309);
and U3606 (N_3606,N_682,N_1527);
or U3607 (N_3607,N_371,N_1143);
nor U3608 (N_3608,N_41,N_2123);
nor U3609 (N_3609,N_110,N_363);
nor U3610 (N_3610,N_76,N_408);
and U3611 (N_3611,N_1560,N_2234);
nand U3612 (N_3612,N_1339,N_1931);
or U3613 (N_3613,N_176,N_2458);
and U3614 (N_3614,N_422,N_548);
or U3615 (N_3615,N_1979,N_672);
and U3616 (N_3616,N_563,N_78);
nor U3617 (N_3617,N_2344,N_476);
and U3618 (N_3618,N_1227,N_1239);
or U3619 (N_3619,N_1775,N_68);
or U3620 (N_3620,N_806,N_2389);
or U3621 (N_3621,N_2445,N_1610);
nor U3622 (N_3622,N_1190,N_1178);
and U3623 (N_3623,N_896,N_2120);
or U3624 (N_3624,N_1503,N_816);
or U3625 (N_3625,N_2329,N_400);
nand U3626 (N_3626,N_2240,N_1026);
nor U3627 (N_3627,N_1015,N_568);
xnor U3628 (N_3628,N_1167,N_295);
and U3629 (N_3629,N_90,N_48);
and U3630 (N_3630,N_2180,N_1703);
nand U3631 (N_3631,N_2471,N_2035);
nor U3632 (N_3632,N_664,N_1951);
or U3633 (N_3633,N_1071,N_1477);
nor U3634 (N_3634,N_725,N_1176);
nor U3635 (N_3635,N_1710,N_597);
or U3636 (N_3636,N_620,N_646);
or U3637 (N_3637,N_1486,N_75);
nor U3638 (N_3638,N_1786,N_1623);
nor U3639 (N_3639,N_1586,N_103);
or U3640 (N_3640,N_291,N_440);
and U3641 (N_3641,N_1161,N_133);
nand U3642 (N_3642,N_1425,N_1788);
or U3643 (N_3643,N_1781,N_1138);
nand U3644 (N_3644,N_310,N_1577);
nor U3645 (N_3645,N_220,N_1698);
nand U3646 (N_3646,N_1020,N_102);
and U3647 (N_3647,N_2435,N_1428);
or U3648 (N_3648,N_2395,N_521);
xor U3649 (N_3649,N_2296,N_507);
or U3650 (N_3650,N_228,N_2369);
or U3651 (N_3651,N_80,N_2076);
or U3652 (N_3652,N_1265,N_2290);
nand U3653 (N_3653,N_2407,N_692);
nand U3654 (N_3654,N_1450,N_2242);
or U3655 (N_3655,N_1058,N_724);
or U3656 (N_3656,N_1505,N_482);
or U3657 (N_3657,N_1165,N_175);
nor U3658 (N_3658,N_447,N_1482);
nand U3659 (N_3659,N_1003,N_2200);
nand U3660 (N_3660,N_1887,N_2031);
nand U3661 (N_3661,N_1185,N_2355);
nand U3662 (N_3662,N_8,N_128);
or U3663 (N_3663,N_6,N_1642);
nor U3664 (N_3664,N_404,N_961);
nor U3665 (N_3665,N_627,N_686);
or U3666 (N_3666,N_13,N_1534);
and U3667 (N_3667,N_137,N_198);
or U3668 (N_3668,N_873,N_1059);
and U3669 (N_3669,N_370,N_1067);
nand U3670 (N_3670,N_636,N_1645);
and U3671 (N_3671,N_1828,N_465);
nor U3672 (N_3672,N_904,N_2402);
or U3673 (N_3673,N_1212,N_962);
nor U3674 (N_3674,N_2232,N_841);
nor U3675 (N_3675,N_4,N_1890);
nor U3676 (N_3676,N_1221,N_1158);
nand U3677 (N_3677,N_1935,N_902);
nor U3678 (N_3678,N_2139,N_1288);
nor U3679 (N_3679,N_1760,N_1704);
nand U3680 (N_3680,N_459,N_2221);
nor U3681 (N_3681,N_1076,N_1646);
or U3682 (N_3682,N_2069,N_919);
or U3683 (N_3683,N_1504,N_821);
nor U3684 (N_3684,N_1729,N_1726);
and U3685 (N_3685,N_2377,N_442);
and U3686 (N_3686,N_2281,N_2284);
and U3687 (N_3687,N_926,N_1439);
nor U3688 (N_3688,N_1184,N_2111);
nand U3689 (N_3689,N_416,N_617);
and U3690 (N_3690,N_963,N_2037);
nor U3691 (N_3691,N_2156,N_1514);
and U3692 (N_3692,N_1080,N_256);
nor U3693 (N_3693,N_1818,N_799);
or U3694 (N_3694,N_1326,N_1798);
and U3695 (N_3695,N_1191,N_1162);
or U3696 (N_3696,N_938,N_1332);
nor U3697 (N_3697,N_1423,N_2022);
and U3698 (N_3698,N_1898,N_1573);
or U3699 (N_3699,N_574,N_141);
xor U3700 (N_3700,N_2208,N_1383);
nor U3701 (N_3701,N_2459,N_224);
nand U3702 (N_3702,N_1563,N_1120);
or U3703 (N_3703,N_1539,N_83);
nor U3704 (N_3704,N_614,N_1507);
and U3705 (N_3705,N_1824,N_832);
and U3706 (N_3706,N_1302,N_1865);
and U3707 (N_3707,N_637,N_577);
nand U3708 (N_3708,N_381,N_1620);
nor U3709 (N_3709,N_2486,N_1575);
nand U3710 (N_3710,N_606,N_1455);
and U3711 (N_3711,N_64,N_1618);
or U3712 (N_3712,N_1022,N_1715);
and U3713 (N_3713,N_1135,N_94);
and U3714 (N_3714,N_272,N_472);
nand U3715 (N_3715,N_972,N_116);
or U3716 (N_3716,N_2217,N_2470);
nor U3717 (N_3717,N_1957,N_127);
and U3718 (N_3718,N_1299,N_611);
nor U3719 (N_3719,N_2275,N_1475);
nand U3720 (N_3720,N_565,N_2114);
or U3721 (N_3721,N_2116,N_1448);
and U3722 (N_3722,N_1525,N_744);
and U3723 (N_3723,N_504,N_1829);
and U3724 (N_3724,N_1817,N_1402);
or U3725 (N_3725,N_803,N_2258);
and U3726 (N_3726,N_1417,N_1027);
or U3727 (N_3727,N_1611,N_1333);
nor U3728 (N_3728,N_1415,N_630);
nand U3729 (N_3729,N_640,N_788);
nand U3730 (N_3730,N_706,N_2489);
and U3731 (N_3731,N_1389,N_1141);
nor U3732 (N_3732,N_1217,N_1395);
and U3733 (N_3733,N_685,N_181);
and U3734 (N_3734,N_296,N_1367);
nor U3735 (N_3735,N_1511,N_768);
and U3736 (N_3736,N_1156,N_1640);
or U3737 (N_3737,N_1777,N_769);
and U3738 (N_3738,N_2256,N_1531);
and U3739 (N_3739,N_262,N_987);
nand U3740 (N_3740,N_1683,N_831);
or U3741 (N_3741,N_2244,N_168);
nor U3742 (N_3742,N_1564,N_1512);
nor U3743 (N_3743,N_715,N_866);
nand U3744 (N_3744,N_1912,N_1944);
or U3745 (N_3745,N_2125,N_830);
nand U3746 (N_3746,N_1374,N_2392);
nand U3747 (N_3747,N_1690,N_1609);
nor U3748 (N_3748,N_223,N_330);
nand U3749 (N_3749,N_1516,N_17);
or U3750 (N_3750,N_659,N_1535);
nor U3751 (N_3751,N_1331,N_1909);
nand U3752 (N_3752,N_1116,N_870);
or U3753 (N_3753,N_576,N_63);
and U3754 (N_3754,N_1928,N_2156);
or U3755 (N_3755,N_1873,N_1922);
or U3756 (N_3756,N_1774,N_1256);
nor U3757 (N_3757,N_1959,N_487);
or U3758 (N_3758,N_2020,N_1253);
or U3759 (N_3759,N_1061,N_216);
nor U3760 (N_3760,N_849,N_804);
nor U3761 (N_3761,N_749,N_876);
nand U3762 (N_3762,N_2142,N_865);
or U3763 (N_3763,N_517,N_2409);
and U3764 (N_3764,N_1807,N_2071);
xnor U3765 (N_3765,N_1421,N_800);
nor U3766 (N_3766,N_924,N_1536);
nor U3767 (N_3767,N_1713,N_664);
or U3768 (N_3768,N_424,N_1330);
nor U3769 (N_3769,N_1364,N_256);
and U3770 (N_3770,N_1444,N_72);
nand U3771 (N_3771,N_738,N_2402);
or U3772 (N_3772,N_2082,N_538);
nor U3773 (N_3773,N_860,N_2175);
and U3774 (N_3774,N_2093,N_1844);
and U3775 (N_3775,N_2289,N_341);
and U3776 (N_3776,N_582,N_152);
nand U3777 (N_3777,N_1270,N_1669);
nor U3778 (N_3778,N_1434,N_2158);
nor U3779 (N_3779,N_1210,N_833);
or U3780 (N_3780,N_1340,N_2432);
nor U3781 (N_3781,N_256,N_1124);
xor U3782 (N_3782,N_1931,N_2446);
nor U3783 (N_3783,N_1140,N_1100);
nand U3784 (N_3784,N_1196,N_1665);
nand U3785 (N_3785,N_2040,N_2426);
and U3786 (N_3786,N_628,N_49);
nor U3787 (N_3787,N_1501,N_899);
and U3788 (N_3788,N_1688,N_1252);
or U3789 (N_3789,N_246,N_2267);
or U3790 (N_3790,N_2178,N_1256);
and U3791 (N_3791,N_2310,N_259);
nor U3792 (N_3792,N_124,N_2375);
nand U3793 (N_3793,N_1997,N_1244);
and U3794 (N_3794,N_1865,N_2456);
or U3795 (N_3795,N_2096,N_842);
nor U3796 (N_3796,N_867,N_1599);
nor U3797 (N_3797,N_622,N_2268);
nor U3798 (N_3798,N_339,N_2021);
nand U3799 (N_3799,N_2400,N_2461);
or U3800 (N_3800,N_478,N_927);
nor U3801 (N_3801,N_2242,N_359);
nor U3802 (N_3802,N_1639,N_2408);
and U3803 (N_3803,N_1215,N_487);
or U3804 (N_3804,N_2391,N_586);
and U3805 (N_3805,N_353,N_1369);
nand U3806 (N_3806,N_1873,N_2431);
nor U3807 (N_3807,N_2498,N_2133);
or U3808 (N_3808,N_626,N_2331);
nor U3809 (N_3809,N_1305,N_543);
nand U3810 (N_3810,N_712,N_2086);
nand U3811 (N_3811,N_827,N_670);
and U3812 (N_3812,N_1121,N_178);
and U3813 (N_3813,N_1376,N_263);
nand U3814 (N_3814,N_1865,N_2015);
and U3815 (N_3815,N_292,N_192);
nand U3816 (N_3816,N_1069,N_912);
and U3817 (N_3817,N_958,N_588);
nor U3818 (N_3818,N_1494,N_169);
and U3819 (N_3819,N_708,N_370);
nand U3820 (N_3820,N_359,N_2270);
and U3821 (N_3821,N_10,N_810);
and U3822 (N_3822,N_72,N_1205);
or U3823 (N_3823,N_632,N_364);
nor U3824 (N_3824,N_2131,N_2061);
and U3825 (N_3825,N_121,N_1607);
nor U3826 (N_3826,N_1412,N_1595);
nand U3827 (N_3827,N_1787,N_1211);
nor U3828 (N_3828,N_2297,N_1982);
and U3829 (N_3829,N_1991,N_1526);
nand U3830 (N_3830,N_451,N_337);
nand U3831 (N_3831,N_196,N_569);
or U3832 (N_3832,N_553,N_965);
nand U3833 (N_3833,N_1888,N_1581);
and U3834 (N_3834,N_2261,N_1014);
or U3835 (N_3835,N_420,N_1702);
nand U3836 (N_3836,N_2065,N_1031);
or U3837 (N_3837,N_1583,N_1345);
and U3838 (N_3838,N_1199,N_160);
or U3839 (N_3839,N_1323,N_808);
and U3840 (N_3840,N_860,N_712);
and U3841 (N_3841,N_2227,N_1308);
nand U3842 (N_3842,N_1902,N_209);
or U3843 (N_3843,N_647,N_1007);
or U3844 (N_3844,N_1303,N_1182);
and U3845 (N_3845,N_151,N_522);
nor U3846 (N_3846,N_518,N_73);
or U3847 (N_3847,N_1740,N_2055);
nor U3848 (N_3848,N_94,N_2061);
nand U3849 (N_3849,N_1615,N_1667);
and U3850 (N_3850,N_490,N_1651);
and U3851 (N_3851,N_1629,N_1633);
or U3852 (N_3852,N_1866,N_571);
nand U3853 (N_3853,N_1478,N_2209);
xor U3854 (N_3854,N_2123,N_2169);
or U3855 (N_3855,N_2082,N_2145);
nand U3856 (N_3856,N_1033,N_215);
nand U3857 (N_3857,N_1292,N_1830);
or U3858 (N_3858,N_2387,N_1228);
and U3859 (N_3859,N_1797,N_570);
and U3860 (N_3860,N_1052,N_2259);
nand U3861 (N_3861,N_652,N_2294);
nor U3862 (N_3862,N_838,N_716);
or U3863 (N_3863,N_1407,N_344);
nand U3864 (N_3864,N_991,N_857);
nor U3865 (N_3865,N_343,N_2408);
nand U3866 (N_3866,N_2332,N_1315);
nor U3867 (N_3867,N_93,N_2485);
or U3868 (N_3868,N_122,N_1671);
and U3869 (N_3869,N_25,N_1225);
or U3870 (N_3870,N_2269,N_1552);
or U3871 (N_3871,N_370,N_633);
or U3872 (N_3872,N_339,N_3);
nand U3873 (N_3873,N_140,N_1986);
nor U3874 (N_3874,N_0,N_1090);
nor U3875 (N_3875,N_2282,N_330);
nand U3876 (N_3876,N_1224,N_2431);
and U3877 (N_3877,N_570,N_891);
nand U3878 (N_3878,N_316,N_1245);
nand U3879 (N_3879,N_1172,N_1393);
and U3880 (N_3880,N_437,N_1909);
and U3881 (N_3881,N_1200,N_1506);
nor U3882 (N_3882,N_934,N_1926);
nand U3883 (N_3883,N_2423,N_1402);
xor U3884 (N_3884,N_1389,N_79);
or U3885 (N_3885,N_1421,N_1730);
nor U3886 (N_3886,N_2406,N_1657);
or U3887 (N_3887,N_1967,N_1471);
nor U3888 (N_3888,N_2477,N_1772);
and U3889 (N_3889,N_1563,N_690);
nand U3890 (N_3890,N_1816,N_105);
nor U3891 (N_3891,N_1978,N_834);
xnor U3892 (N_3892,N_1760,N_2098);
nand U3893 (N_3893,N_2310,N_174);
nand U3894 (N_3894,N_1576,N_696);
and U3895 (N_3895,N_364,N_23);
or U3896 (N_3896,N_1355,N_832);
and U3897 (N_3897,N_409,N_2214);
nand U3898 (N_3898,N_569,N_1670);
and U3899 (N_3899,N_2014,N_835);
nor U3900 (N_3900,N_1130,N_2352);
or U3901 (N_3901,N_838,N_2226);
nor U3902 (N_3902,N_1382,N_1540);
or U3903 (N_3903,N_343,N_752);
nand U3904 (N_3904,N_1382,N_877);
nor U3905 (N_3905,N_2319,N_306);
and U3906 (N_3906,N_15,N_2166);
or U3907 (N_3907,N_1371,N_2132);
nand U3908 (N_3908,N_964,N_2409);
nor U3909 (N_3909,N_1236,N_2081);
and U3910 (N_3910,N_2010,N_1511);
nand U3911 (N_3911,N_318,N_738);
nand U3912 (N_3912,N_677,N_1432);
nor U3913 (N_3913,N_1763,N_353);
nand U3914 (N_3914,N_2452,N_1370);
nand U3915 (N_3915,N_1509,N_949);
nand U3916 (N_3916,N_1399,N_819);
nand U3917 (N_3917,N_865,N_1550);
nand U3918 (N_3918,N_701,N_894);
and U3919 (N_3919,N_979,N_2371);
or U3920 (N_3920,N_979,N_896);
or U3921 (N_3921,N_1527,N_1724);
xor U3922 (N_3922,N_711,N_1909);
nor U3923 (N_3923,N_874,N_1967);
nand U3924 (N_3924,N_1276,N_2275);
or U3925 (N_3925,N_338,N_2140);
or U3926 (N_3926,N_2386,N_1349);
or U3927 (N_3927,N_2214,N_2114);
and U3928 (N_3928,N_1568,N_1564);
and U3929 (N_3929,N_2132,N_432);
or U3930 (N_3930,N_2243,N_1559);
and U3931 (N_3931,N_2374,N_1961);
nor U3932 (N_3932,N_483,N_1481);
and U3933 (N_3933,N_2119,N_2146);
nor U3934 (N_3934,N_2187,N_591);
nor U3935 (N_3935,N_2053,N_1353);
and U3936 (N_3936,N_1092,N_861);
nor U3937 (N_3937,N_901,N_1346);
and U3938 (N_3938,N_2219,N_1645);
and U3939 (N_3939,N_1194,N_994);
nor U3940 (N_3940,N_569,N_2404);
or U3941 (N_3941,N_1806,N_1443);
nor U3942 (N_3942,N_1577,N_2227);
or U3943 (N_3943,N_825,N_822);
and U3944 (N_3944,N_39,N_709);
or U3945 (N_3945,N_1294,N_1334);
nand U3946 (N_3946,N_1022,N_2435);
nor U3947 (N_3947,N_1552,N_1115);
nor U3948 (N_3948,N_1391,N_1243);
or U3949 (N_3949,N_2481,N_1936);
nand U3950 (N_3950,N_939,N_952);
and U3951 (N_3951,N_700,N_189);
nand U3952 (N_3952,N_597,N_2100);
nor U3953 (N_3953,N_1533,N_149);
and U3954 (N_3954,N_537,N_113);
and U3955 (N_3955,N_897,N_1182);
or U3956 (N_3956,N_1152,N_441);
nand U3957 (N_3957,N_77,N_61);
nor U3958 (N_3958,N_1532,N_887);
and U3959 (N_3959,N_1835,N_763);
or U3960 (N_3960,N_233,N_1040);
nand U3961 (N_3961,N_1151,N_606);
nor U3962 (N_3962,N_460,N_1609);
nand U3963 (N_3963,N_1434,N_1911);
or U3964 (N_3964,N_1567,N_1875);
or U3965 (N_3965,N_1942,N_513);
nor U3966 (N_3966,N_1772,N_364);
or U3967 (N_3967,N_2045,N_2490);
and U3968 (N_3968,N_1837,N_1097);
or U3969 (N_3969,N_2057,N_1778);
nor U3970 (N_3970,N_180,N_1081);
or U3971 (N_3971,N_2054,N_1621);
or U3972 (N_3972,N_1275,N_1426);
or U3973 (N_3973,N_1805,N_774);
and U3974 (N_3974,N_1237,N_299);
nor U3975 (N_3975,N_2139,N_1813);
nor U3976 (N_3976,N_2136,N_2054);
nor U3977 (N_3977,N_1260,N_865);
or U3978 (N_3978,N_842,N_2063);
or U3979 (N_3979,N_1535,N_1805);
or U3980 (N_3980,N_998,N_2153);
or U3981 (N_3981,N_2081,N_1263);
or U3982 (N_3982,N_1739,N_492);
nor U3983 (N_3983,N_34,N_1060);
nor U3984 (N_3984,N_2371,N_1727);
or U3985 (N_3985,N_106,N_668);
xor U3986 (N_3986,N_572,N_2350);
or U3987 (N_3987,N_264,N_1264);
nand U3988 (N_3988,N_37,N_1514);
nand U3989 (N_3989,N_283,N_1483);
and U3990 (N_3990,N_1887,N_1274);
and U3991 (N_3991,N_2451,N_1217);
or U3992 (N_3992,N_75,N_959);
nand U3993 (N_3993,N_39,N_2452);
or U3994 (N_3994,N_2426,N_1447);
or U3995 (N_3995,N_1079,N_609);
and U3996 (N_3996,N_1125,N_2315);
and U3997 (N_3997,N_2265,N_1052);
nor U3998 (N_3998,N_2216,N_391);
nand U3999 (N_3999,N_163,N_2161);
and U4000 (N_4000,N_2278,N_2091);
or U4001 (N_4001,N_1782,N_2302);
and U4002 (N_4002,N_234,N_664);
xor U4003 (N_4003,N_457,N_205);
or U4004 (N_4004,N_2243,N_1536);
nor U4005 (N_4005,N_2118,N_264);
nor U4006 (N_4006,N_1747,N_1867);
nor U4007 (N_4007,N_95,N_639);
or U4008 (N_4008,N_1792,N_794);
nand U4009 (N_4009,N_1215,N_902);
and U4010 (N_4010,N_1476,N_1171);
and U4011 (N_4011,N_301,N_1166);
and U4012 (N_4012,N_1026,N_1053);
nand U4013 (N_4013,N_451,N_2376);
or U4014 (N_4014,N_1510,N_1149);
or U4015 (N_4015,N_937,N_1398);
nor U4016 (N_4016,N_223,N_1686);
or U4017 (N_4017,N_1666,N_1356);
and U4018 (N_4018,N_1832,N_483);
or U4019 (N_4019,N_1953,N_297);
or U4020 (N_4020,N_375,N_955);
nor U4021 (N_4021,N_1626,N_480);
nand U4022 (N_4022,N_1766,N_2384);
nand U4023 (N_4023,N_1851,N_1370);
nand U4024 (N_4024,N_744,N_872);
nand U4025 (N_4025,N_1250,N_491);
and U4026 (N_4026,N_345,N_2195);
or U4027 (N_4027,N_459,N_553);
nand U4028 (N_4028,N_610,N_706);
or U4029 (N_4029,N_1758,N_487);
nor U4030 (N_4030,N_1868,N_2333);
nor U4031 (N_4031,N_275,N_129);
or U4032 (N_4032,N_1015,N_1029);
and U4033 (N_4033,N_750,N_840);
nor U4034 (N_4034,N_2381,N_1948);
or U4035 (N_4035,N_1412,N_1778);
and U4036 (N_4036,N_455,N_710);
and U4037 (N_4037,N_1922,N_16);
nand U4038 (N_4038,N_898,N_154);
nor U4039 (N_4039,N_410,N_176);
nor U4040 (N_4040,N_185,N_2065);
or U4041 (N_4041,N_388,N_340);
nand U4042 (N_4042,N_1093,N_138);
nand U4043 (N_4043,N_313,N_345);
or U4044 (N_4044,N_1921,N_2381);
nor U4045 (N_4045,N_2324,N_2444);
or U4046 (N_4046,N_1482,N_1517);
nor U4047 (N_4047,N_1317,N_1390);
and U4048 (N_4048,N_1564,N_2449);
nand U4049 (N_4049,N_336,N_370);
nor U4050 (N_4050,N_488,N_1896);
or U4051 (N_4051,N_829,N_2118);
and U4052 (N_4052,N_1399,N_2012);
or U4053 (N_4053,N_268,N_1252);
nor U4054 (N_4054,N_524,N_447);
nor U4055 (N_4055,N_1645,N_2246);
nor U4056 (N_4056,N_1261,N_663);
nor U4057 (N_4057,N_2363,N_1399);
or U4058 (N_4058,N_1535,N_1019);
or U4059 (N_4059,N_968,N_1715);
nand U4060 (N_4060,N_1849,N_729);
nand U4061 (N_4061,N_548,N_201);
xor U4062 (N_4062,N_142,N_1454);
nand U4063 (N_4063,N_478,N_2498);
or U4064 (N_4064,N_1864,N_507);
or U4065 (N_4065,N_771,N_766);
or U4066 (N_4066,N_1218,N_746);
and U4067 (N_4067,N_2163,N_1715);
nor U4068 (N_4068,N_2199,N_1923);
nor U4069 (N_4069,N_877,N_1047);
or U4070 (N_4070,N_956,N_1492);
nand U4071 (N_4071,N_880,N_1827);
or U4072 (N_4072,N_2227,N_1147);
and U4073 (N_4073,N_592,N_1110);
or U4074 (N_4074,N_1132,N_1123);
and U4075 (N_4075,N_1754,N_322);
nor U4076 (N_4076,N_243,N_1077);
or U4077 (N_4077,N_2002,N_1556);
and U4078 (N_4078,N_522,N_102);
nand U4079 (N_4079,N_1209,N_2490);
and U4080 (N_4080,N_1611,N_1049);
nand U4081 (N_4081,N_1268,N_1695);
nand U4082 (N_4082,N_381,N_1516);
nand U4083 (N_4083,N_1912,N_2100);
nand U4084 (N_4084,N_2029,N_1300);
nor U4085 (N_4085,N_1249,N_1611);
or U4086 (N_4086,N_2406,N_1214);
and U4087 (N_4087,N_2050,N_399);
nor U4088 (N_4088,N_796,N_1910);
nand U4089 (N_4089,N_1812,N_479);
and U4090 (N_4090,N_596,N_2014);
or U4091 (N_4091,N_517,N_1120);
nor U4092 (N_4092,N_1336,N_996);
and U4093 (N_4093,N_1283,N_2208);
and U4094 (N_4094,N_621,N_700);
or U4095 (N_4095,N_1193,N_697);
nor U4096 (N_4096,N_370,N_95);
and U4097 (N_4097,N_124,N_980);
nand U4098 (N_4098,N_83,N_2149);
nor U4099 (N_4099,N_873,N_1946);
xnor U4100 (N_4100,N_2113,N_919);
nor U4101 (N_4101,N_2272,N_2441);
or U4102 (N_4102,N_1368,N_1320);
and U4103 (N_4103,N_2452,N_1440);
and U4104 (N_4104,N_2486,N_2060);
and U4105 (N_4105,N_488,N_1925);
nor U4106 (N_4106,N_770,N_1189);
nor U4107 (N_4107,N_1500,N_1088);
nor U4108 (N_4108,N_1407,N_940);
nor U4109 (N_4109,N_2005,N_182);
or U4110 (N_4110,N_311,N_1799);
or U4111 (N_4111,N_1091,N_1086);
nor U4112 (N_4112,N_942,N_165);
xor U4113 (N_4113,N_1277,N_1191);
nand U4114 (N_4114,N_118,N_1860);
nor U4115 (N_4115,N_1787,N_2408);
and U4116 (N_4116,N_705,N_44);
or U4117 (N_4117,N_1896,N_2185);
nor U4118 (N_4118,N_773,N_1955);
nand U4119 (N_4119,N_2014,N_215);
or U4120 (N_4120,N_2332,N_1908);
nor U4121 (N_4121,N_1999,N_1911);
nor U4122 (N_4122,N_110,N_1308);
and U4123 (N_4123,N_740,N_1932);
or U4124 (N_4124,N_2126,N_1744);
nor U4125 (N_4125,N_2469,N_2169);
or U4126 (N_4126,N_288,N_1627);
nor U4127 (N_4127,N_1604,N_31);
nor U4128 (N_4128,N_2241,N_2395);
nand U4129 (N_4129,N_2481,N_2270);
nand U4130 (N_4130,N_1261,N_1832);
and U4131 (N_4131,N_1930,N_457);
or U4132 (N_4132,N_287,N_2156);
and U4133 (N_4133,N_1548,N_1532);
nor U4134 (N_4134,N_1428,N_842);
nor U4135 (N_4135,N_1816,N_1544);
or U4136 (N_4136,N_1857,N_149);
and U4137 (N_4137,N_1495,N_231);
nor U4138 (N_4138,N_421,N_2166);
and U4139 (N_4139,N_299,N_115);
nor U4140 (N_4140,N_1914,N_2354);
and U4141 (N_4141,N_749,N_2128);
nand U4142 (N_4142,N_1615,N_2147);
or U4143 (N_4143,N_531,N_454);
nor U4144 (N_4144,N_791,N_457);
and U4145 (N_4145,N_2155,N_2356);
nor U4146 (N_4146,N_1556,N_165);
nor U4147 (N_4147,N_2165,N_1150);
or U4148 (N_4148,N_75,N_1143);
nor U4149 (N_4149,N_294,N_467);
nand U4150 (N_4150,N_102,N_1181);
xnor U4151 (N_4151,N_1439,N_573);
nor U4152 (N_4152,N_2171,N_1717);
nor U4153 (N_4153,N_1834,N_1236);
xor U4154 (N_4154,N_1638,N_1328);
or U4155 (N_4155,N_406,N_2374);
or U4156 (N_4156,N_751,N_2425);
or U4157 (N_4157,N_2374,N_506);
or U4158 (N_4158,N_1493,N_1371);
and U4159 (N_4159,N_729,N_2455);
and U4160 (N_4160,N_1009,N_2189);
nand U4161 (N_4161,N_1901,N_683);
or U4162 (N_4162,N_1142,N_2003);
nor U4163 (N_4163,N_1751,N_984);
or U4164 (N_4164,N_1370,N_968);
nand U4165 (N_4165,N_1970,N_808);
nand U4166 (N_4166,N_1366,N_1039);
and U4167 (N_4167,N_1831,N_1319);
or U4168 (N_4168,N_130,N_2455);
or U4169 (N_4169,N_999,N_1525);
and U4170 (N_4170,N_181,N_1254);
nand U4171 (N_4171,N_1052,N_361);
nand U4172 (N_4172,N_520,N_296);
nor U4173 (N_4173,N_2220,N_1008);
and U4174 (N_4174,N_2309,N_1291);
xnor U4175 (N_4175,N_669,N_353);
and U4176 (N_4176,N_20,N_1);
nand U4177 (N_4177,N_372,N_825);
nand U4178 (N_4178,N_817,N_988);
nor U4179 (N_4179,N_1318,N_640);
or U4180 (N_4180,N_202,N_423);
nand U4181 (N_4181,N_1135,N_666);
nand U4182 (N_4182,N_1527,N_845);
and U4183 (N_4183,N_901,N_2049);
or U4184 (N_4184,N_816,N_2101);
xor U4185 (N_4185,N_1760,N_328);
or U4186 (N_4186,N_2202,N_187);
nand U4187 (N_4187,N_1133,N_2135);
or U4188 (N_4188,N_1252,N_2282);
nand U4189 (N_4189,N_224,N_1269);
nand U4190 (N_4190,N_2224,N_797);
or U4191 (N_4191,N_1064,N_1691);
or U4192 (N_4192,N_233,N_2317);
and U4193 (N_4193,N_119,N_1679);
and U4194 (N_4194,N_1908,N_128);
or U4195 (N_4195,N_1254,N_944);
or U4196 (N_4196,N_1499,N_430);
or U4197 (N_4197,N_457,N_792);
or U4198 (N_4198,N_2479,N_1187);
and U4199 (N_4199,N_1367,N_2415);
and U4200 (N_4200,N_21,N_1718);
or U4201 (N_4201,N_908,N_1612);
or U4202 (N_4202,N_497,N_58);
or U4203 (N_4203,N_2157,N_369);
nand U4204 (N_4204,N_113,N_2076);
and U4205 (N_4205,N_1932,N_872);
and U4206 (N_4206,N_1329,N_1747);
nor U4207 (N_4207,N_2491,N_464);
nand U4208 (N_4208,N_1973,N_58);
nor U4209 (N_4209,N_2030,N_1554);
and U4210 (N_4210,N_2256,N_37);
nand U4211 (N_4211,N_2013,N_1690);
or U4212 (N_4212,N_45,N_188);
nor U4213 (N_4213,N_874,N_1959);
nor U4214 (N_4214,N_1503,N_478);
nor U4215 (N_4215,N_1193,N_1408);
or U4216 (N_4216,N_843,N_317);
or U4217 (N_4217,N_1019,N_2378);
or U4218 (N_4218,N_1176,N_500);
nand U4219 (N_4219,N_494,N_2488);
or U4220 (N_4220,N_764,N_72);
nor U4221 (N_4221,N_1013,N_2392);
nor U4222 (N_4222,N_2308,N_624);
nor U4223 (N_4223,N_573,N_517);
nor U4224 (N_4224,N_321,N_1436);
and U4225 (N_4225,N_2187,N_328);
nor U4226 (N_4226,N_2125,N_351);
or U4227 (N_4227,N_1324,N_1427);
nor U4228 (N_4228,N_1441,N_1517);
nand U4229 (N_4229,N_429,N_547);
and U4230 (N_4230,N_410,N_488);
and U4231 (N_4231,N_773,N_291);
nand U4232 (N_4232,N_1286,N_2272);
or U4233 (N_4233,N_2041,N_1386);
or U4234 (N_4234,N_1307,N_2486);
or U4235 (N_4235,N_472,N_2494);
and U4236 (N_4236,N_280,N_515);
nand U4237 (N_4237,N_2428,N_159);
or U4238 (N_4238,N_696,N_1590);
nor U4239 (N_4239,N_2043,N_644);
nand U4240 (N_4240,N_247,N_1352);
nand U4241 (N_4241,N_1718,N_1498);
nor U4242 (N_4242,N_1516,N_1073);
nand U4243 (N_4243,N_326,N_2467);
nor U4244 (N_4244,N_67,N_1101);
nor U4245 (N_4245,N_839,N_1222);
nand U4246 (N_4246,N_571,N_1537);
and U4247 (N_4247,N_2152,N_491);
nand U4248 (N_4248,N_1659,N_1546);
nor U4249 (N_4249,N_1256,N_331);
nand U4250 (N_4250,N_2278,N_2049);
nor U4251 (N_4251,N_1409,N_1946);
nor U4252 (N_4252,N_1260,N_1489);
and U4253 (N_4253,N_1545,N_1636);
nor U4254 (N_4254,N_812,N_62);
or U4255 (N_4255,N_843,N_1876);
nor U4256 (N_4256,N_2329,N_2116);
or U4257 (N_4257,N_293,N_1381);
nor U4258 (N_4258,N_764,N_429);
or U4259 (N_4259,N_1704,N_1201);
nor U4260 (N_4260,N_1457,N_2399);
nor U4261 (N_4261,N_184,N_2356);
nand U4262 (N_4262,N_2019,N_1399);
and U4263 (N_4263,N_74,N_2292);
or U4264 (N_4264,N_2179,N_2214);
nand U4265 (N_4265,N_865,N_155);
and U4266 (N_4266,N_1066,N_53);
nor U4267 (N_4267,N_870,N_1499);
nor U4268 (N_4268,N_310,N_556);
or U4269 (N_4269,N_1794,N_212);
or U4270 (N_4270,N_1179,N_2023);
nand U4271 (N_4271,N_51,N_1026);
and U4272 (N_4272,N_603,N_127);
and U4273 (N_4273,N_1803,N_1519);
and U4274 (N_4274,N_1603,N_1385);
nand U4275 (N_4275,N_470,N_2181);
or U4276 (N_4276,N_2099,N_1510);
nor U4277 (N_4277,N_436,N_1927);
nand U4278 (N_4278,N_2455,N_1774);
nand U4279 (N_4279,N_1477,N_1247);
nand U4280 (N_4280,N_1646,N_2178);
nand U4281 (N_4281,N_1340,N_2352);
or U4282 (N_4282,N_1766,N_2415);
or U4283 (N_4283,N_1443,N_2071);
nand U4284 (N_4284,N_2329,N_1989);
nand U4285 (N_4285,N_825,N_209);
nor U4286 (N_4286,N_229,N_1769);
nor U4287 (N_4287,N_1586,N_893);
nor U4288 (N_4288,N_2373,N_1746);
and U4289 (N_4289,N_674,N_270);
or U4290 (N_4290,N_1260,N_692);
and U4291 (N_4291,N_2264,N_105);
nor U4292 (N_4292,N_517,N_1260);
nand U4293 (N_4293,N_1149,N_90);
nor U4294 (N_4294,N_1959,N_2182);
nor U4295 (N_4295,N_301,N_11);
and U4296 (N_4296,N_2464,N_1343);
or U4297 (N_4297,N_1364,N_1861);
and U4298 (N_4298,N_591,N_509);
and U4299 (N_4299,N_1069,N_2110);
or U4300 (N_4300,N_1170,N_14);
nor U4301 (N_4301,N_1450,N_2343);
xor U4302 (N_4302,N_1732,N_318);
or U4303 (N_4303,N_1429,N_216);
or U4304 (N_4304,N_2446,N_2498);
nor U4305 (N_4305,N_1498,N_2265);
and U4306 (N_4306,N_2351,N_1128);
nand U4307 (N_4307,N_33,N_2080);
and U4308 (N_4308,N_232,N_608);
nand U4309 (N_4309,N_1691,N_1072);
nor U4310 (N_4310,N_2349,N_777);
nor U4311 (N_4311,N_635,N_579);
nor U4312 (N_4312,N_1480,N_1164);
or U4313 (N_4313,N_1833,N_220);
or U4314 (N_4314,N_144,N_468);
nand U4315 (N_4315,N_876,N_1329);
and U4316 (N_4316,N_2387,N_752);
nor U4317 (N_4317,N_1180,N_1814);
nor U4318 (N_4318,N_436,N_421);
or U4319 (N_4319,N_1907,N_2483);
or U4320 (N_4320,N_347,N_524);
and U4321 (N_4321,N_1036,N_283);
and U4322 (N_4322,N_1232,N_2367);
or U4323 (N_4323,N_700,N_1062);
or U4324 (N_4324,N_711,N_616);
nor U4325 (N_4325,N_478,N_1544);
and U4326 (N_4326,N_409,N_2373);
nand U4327 (N_4327,N_1032,N_2363);
and U4328 (N_4328,N_1736,N_2417);
and U4329 (N_4329,N_1487,N_1512);
and U4330 (N_4330,N_1365,N_1255);
or U4331 (N_4331,N_403,N_2099);
or U4332 (N_4332,N_2425,N_1180);
and U4333 (N_4333,N_1822,N_112);
or U4334 (N_4334,N_220,N_2279);
and U4335 (N_4335,N_893,N_2407);
nor U4336 (N_4336,N_207,N_64);
nand U4337 (N_4337,N_230,N_1870);
nand U4338 (N_4338,N_1693,N_1319);
or U4339 (N_4339,N_2358,N_1128);
or U4340 (N_4340,N_1570,N_490);
nand U4341 (N_4341,N_1587,N_2424);
and U4342 (N_4342,N_1766,N_625);
nor U4343 (N_4343,N_2007,N_2287);
and U4344 (N_4344,N_1698,N_533);
nor U4345 (N_4345,N_1506,N_638);
and U4346 (N_4346,N_1747,N_1669);
nand U4347 (N_4347,N_4,N_1256);
and U4348 (N_4348,N_2387,N_2140);
nor U4349 (N_4349,N_1419,N_917);
and U4350 (N_4350,N_1385,N_2480);
nor U4351 (N_4351,N_1876,N_1490);
and U4352 (N_4352,N_1898,N_1726);
and U4353 (N_4353,N_1513,N_210);
or U4354 (N_4354,N_536,N_202);
nand U4355 (N_4355,N_59,N_772);
and U4356 (N_4356,N_556,N_877);
nor U4357 (N_4357,N_1188,N_186);
nor U4358 (N_4358,N_448,N_1647);
or U4359 (N_4359,N_1136,N_1237);
nand U4360 (N_4360,N_576,N_1045);
nor U4361 (N_4361,N_1286,N_2187);
nand U4362 (N_4362,N_770,N_328);
nand U4363 (N_4363,N_1031,N_748);
or U4364 (N_4364,N_107,N_25);
or U4365 (N_4365,N_2062,N_1150);
and U4366 (N_4366,N_1459,N_901);
or U4367 (N_4367,N_695,N_215);
and U4368 (N_4368,N_1955,N_2110);
nand U4369 (N_4369,N_12,N_426);
nand U4370 (N_4370,N_748,N_605);
nor U4371 (N_4371,N_1371,N_2085);
nor U4372 (N_4372,N_796,N_552);
or U4373 (N_4373,N_1788,N_640);
nand U4374 (N_4374,N_1762,N_1787);
or U4375 (N_4375,N_428,N_2312);
nor U4376 (N_4376,N_2252,N_2238);
nor U4377 (N_4377,N_738,N_2121);
or U4378 (N_4378,N_2337,N_1120);
nand U4379 (N_4379,N_76,N_1526);
and U4380 (N_4380,N_1925,N_114);
nor U4381 (N_4381,N_1750,N_225);
nor U4382 (N_4382,N_1462,N_1461);
nor U4383 (N_4383,N_1910,N_25);
nand U4384 (N_4384,N_458,N_1944);
and U4385 (N_4385,N_114,N_2337);
nor U4386 (N_4386,N_907,N_559);
nor U4387 (N_4387,N_2062,N_277);
and U4388 (N_4388,N_946,N_1333);
and U4389 (N_4389,N_2160,N_1986);
or U4390 (N_4390,N_137,N_931);
nor U4391 (N_4391,N_2301,N_1797);
and U4392 (N_4392,N_818,N_424);
nor U4393 (N_4393,N_141,N_298);
or U4394 (N_4394,N_1092,N_2474);
and U4395 (N_4395,N_2297,N_670);
nor U4396 (N_4396,N_274,N_1997);
nand U4397 (N_4397,N_1382,N_1133);
or U4398 (N_4398,N_1218,N_1090);
or U4399 (N_4399,N_976,N_1869);
nand U4400 (N_4400,N_685,N_1529);
nor U4401 (N_4401,N_89,N_1149);
or U4402 (N_4402,N_539,N_1236);
and U4403 (N_4403,N_567,N_2455);
and U4404 (N_4404,N_2289,N_794);
nand U4405 (N_4405,N_1849,N_1131);
nor U4406 (N_4406,N_2196,N_794);
nor U4407 (N_4407,N_493,N_1599);
or U4408 (N_4408,N_1727,N_225);
nand U4409 (N_4409,N_1682,N_492);
or U4410 (N_4410,N_1598,N_413);
or U4411 (N_4411,N_1077,N_1911);
nand U4412 (N_4412,N_2468,N_172);
nand U4413 (N_4413,N_1241,N_33);
or U4414 (N_4414,N_378,N_2004);
nor U4415 (N_4415,N_1172,N_1056);
nor U4416 (N_4416,N_1794,N_760);
nor U4417 (N_4417,N_855,N_371);
or U4418 (N_4418,N_392,N_1130);
or U4419 (N_4419,N_1353,N_456);
xor U4420 (N_4420,N_503,N_432);
nor U4421 (N_4421,N_185,N_602);
nand U4422 (N_4422,N_1771,N_495);
or U4423 (N_4423,N_1320,N_1610);
nor U4424 (N_4424,N_804,N_716);
nor U4425 (N_4425,N_2490,N_2461);
or U4426 (N_4426,N_1245,N_2374);
or U4427 (N_4427,N_1897,N_840);
and U4428 (N_4428,N_762,N_687);
nor U4429 (N_4429,N_86,N_1112);
or U4430 (N_4430,N_965,N_703);
nand U4431 (N_4431,N_933,N_1939);
or U4432 (N_4432,N_1788,N_1624);
or U4433 (N_4433,N_1755,N_1668);
nand U4434 (N_4434,N_1418,N_2328);
nor U4435 (N_4435,N_664,N_1044);
nand U4436 (N_4436,N_357,N_7);
or U4437 (N_4437,N_1434,N_1760);
nand U4438 (N_4438,N_173,N_2490);
and U4439 (N_4439,N_495,N_615);
nor U4440 (N_4440,N_141,N_2311);
or U4441 (N_4441,N_2411,N_2202);
nand U4442 (N_4442,N_1847,N_499);
xnor U4443 (N_4443,N_664,N_2487);
nor U4444 (N_4444,N_511,N_1639);
nand U4445 (N_4445,N_2497,N_1067);
nand U4446 (N_4446,N_415,N_1161);
nand U4447 (N_4447,N_95,N_2239);
and U4448 (N_4448,N_378,N_661);
or U4449 (N_4449,N_2352,N_932);
nand U4450 (N_4450,N_883,N_1534);
and U4451 (N_4451,N_2410,N_1792);
and U4452 (N_4452,N_1180,N_1001);
nand U4453 (N_4453,N_1285,N_1225);
and U4454 (N_4454,N_1310,N_49);
nand U4455 (N_4455,N_776,N_364);
or U4456 (N_4456,N_930,N_667);
or U4457 (N_4457,N_1578,N_2387);
xnor U4458 (N_4458,N_1410,N_1398);
nor U4459 (N_4459,N_1321,N_1807);
or U4460 (N_4460,N_1300,N_1354);
or U4461 (N_4461,N_781,N_2308);
and U4462 (N_4462,N_353,N_1917);
or U4463 (N_4463,N_301,N_2303);
nand U4464 (N_4464,N_1256,N_2151);
nand U4465 (N_4465,N_1329,N_499);
and U4466 (N_4466,N_1536,N_1889);
nor U4467 (N_4467,N_2310,N_1701);
or U4468 (N_4468,N_1546,N_1489);
nand U4469 (N_4469,N_1791,N_1561);
or U4470 (N_4470,N_1948,N_1172);
xor U4471 (N_4471,N_1728,N_1309);
nand U4472 (N_4472,N_1151,N_398);
and U4473 (N_4473,N_987,N_1972);
or U4474 (N_4474,N_2402,N_1413);
nor U4475 (N_4475,N_1006,N_262);
or U4476 (N_4476,N_1731,N_2444);
or U4477 (N_4477,N_1732,N_548);
and U4478 (N_4478,N_2151,N_220);
and U4479 (N_4479,N_1854,N_502);
and U4480 (N_4480,N_654,N_1711);
nor U4481 (N_4481,N_722,N_1664);
nor U4482 (N_4482,N_1442,N_1474);
or U4483 (N_4483,N_227,N_2357);
nand U4484 (N_4484,N_2106,N_2149);
and U4485 (N_4485,N_1563,N_294);
and U4486 (N_4486,N_219,N_1530);
nor U4487 (N_4487,N_2118,N_2219);
nand U4488 (N_4488,N_349,N_1060);
nor U4489 (N_4489,N_189,N_2271);
and U4490 (N_4490,N_763,N_665);
nand U4491 (N_4491,N_1833,N_2296);
or U4492 (N_4492,N_2334,N_337);
and U4493 (N_4493,N_159,N_2393);
nand U4494 (N_4494,N_1820,N_2374);
or U4495 (N_4495,N_1779,N_2164);
and U4496 (N_4496,N_60,N_621);
nand U4497 (N_4497,N_1052,N_342);
or U4498 (N_4498,N_1513,N_2024);
nor U4499 (N_4499,N_530,N_668);
nor U4500 (N_4500,N_845,N_301);
and U4501 (N_4501,N_612,N_656);
nand U4502 (N_4502,N_64,N_397);
nor U4503 (N_4503,N_1868,N_2494);
or U4504 (N_4504,N_1803,N_2251);
nand U4505 (N_4505,N_578,N_399);
or U4506 (N_4506,N_2132,N_966);
or U4507 (N_4507,N_1951,N_1692);
nor U4508 (N_4508,N_1428,N_1222);
or U4509 (N_4509,N_199,N_1992);
nor U4510 (N_4510,N_1349,N_749);
or U4511 (N_4511,N_976,N_1947);
and U4512 (N_4512,N_2077,N_1309);
nor U4513 (N_4513,N_683,N_1216);
or U4514 (N_4514,N_1324,N_1154);
or U4515 (N_4515,N_1265,N_1513);
or U4516 (N_4516,N_509,N_1443);
and U4517 (N_4517,N_1568,N_473);
nand U4518 (N_4518,N_1059,N_1430);
and U4519 (N_4519,N_1143,N_2147);
and U4520 (N_4520,N_104,N_516);
xor U4521 (N_4521,N_1077,N_1392);
or U4522 (N_4522,N_1103,N_1086);
or U4523 (N_4523,N_253,N_1210);
and U4524 (N_4524,N_146,N_1502);
nand U4525 (N_4525,N_2415,N_1090);
nor U4526 (N_4526,N_20,N_1438);
nand U4527 (N_4527,N_1727,N_1306);
or U4528 (N_4528,N_1456,N_135);
and U4529 (N_4529,N_440,N_967);
or U4530 (N_4530,N_478,N_2112);
nand U4531 (N_4531,N_2406,N_744);
or U4532 (N_4532,N_2079,N_1403);
nand U4533 (N_4533,N_1061,N_1218);
and U4534 (N_4534,N_964,N_1251);
nor U4535 (N_4535,N_1596,N_1758);
nand U4536 (N_4536,N_317,N_115);
and U4537 (N_4537,N_812,N_793);
nand U4538 (N_4538,N_915,N_1754);
or U4539 (N_4539,N_536,N_344);
nor U4540 (N_4540,N_333,N_1159);
xor U4541 (N_4541,N_1490,N_680);
and U4542 (N_4542,N_40,N_1389);
or U4543 (N_4543,N_2397,N_650);
nor U4544 (N_4544,N_1620,N_1007);
and U4545 (N_4545,N_1976,N_1988);
or U4546 (N_4546,N_181,N_2013);
and U4547 (N_4547,N_479,N_1167);
or U4548 (N_4548,N_300,N_1496);
or U4549 (N_4549,N_1799,N_227);
nor U4550 (N_4550,N_1920,N_1495);
or U4551 (N_4551,N_75,N_2348);
nor U4552 (N_4552,N_441,N_1920);
nand U4553 (N_4553,N_1794,N_1597);
nor U4554 (N_4554,N_2144,N_906);
nor U4555 (N_4555,N_981,N_1721);
nor U4556 (N_4556,N_1547,N_1371);
nor U4557 (N_4557,N_96,N_1370);
nand U4558 (N_4558,N_1835,N_2315);
and U4559 (N_4559,N_2121,N_70);
nor U4560 (N_4560,N_803,N_276);
nand U4561 (N_4561,N_722,N_899);
or U4562 (N_4562,N_1965,N_915);
nand U4563 (N_4563,N_231,N_2244);
or U4564 (N_4564,N_1774,N_150);
or U4565 (N_4565,N_109,N_1139);
nand U4566 (N_4566,N_774,N_4);
nand U4567 (N_4567,N_444,N_350);
nand U4568 (N_4568,N_389,N_2300);
and U4569 (N_4569,N_112,N_673);
and U4570 (N_4570,N_1808,N_1774);
or U4571 (N_4571,N_2298,N_67);
and U4572 (N_4572,N_1308,N_457);
nor U4573 (N_4573,N_1005,N_1420);
and U4574 (N_4574,N_50,N_861);
or U4575 (N_4575,N_2180,N_1729);
and U4576 (N_4576,N_54,N_2241);
nor U4577 (N_4577,N_1903,N_205);
nand U4578 (N_4578,N_1734,N_1011);
and U4579 (N_4579,N_1283,N_441);
nand U4580 (N_4580,N_1422,N_294);
or U4581 (N_4581,N_716,N_340);
nor U4582 (N_4582,N_2030,N_2035);
and U4583 (N_4583,N_2426,N_1456);
or U4584 (N_4584,N_664,N_211);
or U4585 (N_4585,N_543,N_475);
or U4586 (N_4586,N_999,N_1122);
or U4587 (N_4587,N_452,N_2271);
or U4588 (N_4588,N_2457,N_1453);
or U4589 (N_4589,N_1089,N_1053);
nor U4590 (N_4590,N_40,N_2314);
nand U4591 (N_4591,N_1079,N_1666);
or U4592 (N_4592,N_262,N_173);
and U4593 (N_4593,N_677,N_1203);
and U4594 (N_4594,N_324,N_2210);
xor U4595 (N_4595,N_1783,N_1832);
nand U4596 (N_4596,N_882,N_2363);
or U4597 (N_4597,N_1905,N_940);
and U4598 (N_4598,N_102,N_744);
nand U4599 (N_4599,N_1269,N_1907);
nand U4600 (N_4600,N_479,N_2325);
nand U4601 (N_4601,N_2268,N_1196);
nor U4602 (N_4602,N_218,N_482);
nor U4603 (N_4603,N_2156,N_2145);
nor U4604 (N_4604,N_15,N_1809);
and U4605 (N_4605,N_2369,N_685);
and U4606 (N_4606,N_2123,N_1017);
nand U4607 (N_4607,N_2494,N_1804);
nand U4608 (N_4608,N_2065,N_2284);
nand U4609 (N_4609,N_2119,N_1379);
or U4610 (N_4610,N_1014,N_757);
xnor U4611 (N_4611,N_1842,N_1833);
nand U4612 (N_4612,N_2059,N_857);
nand U4613 (N_4613,N_2265,N_413);
and U4614 (N_4614,N_1622,N_2040);
and U4615 (N_4615,N_777,N_39);
or U4616 (N_4616,N_721,N_395);
nand U4617 (N_4617,N_611,N_646);
or U4618 (N_4618,N_1499,N_1930);
nand U4619 (N_4619,N_1934,N_1391);
nand U4620 (N_4620,N_2075,N_1075);
or U4621 (N_4621,N_1413,N_163);
xnor U4622 (N_4622,N_1542,N_184);
nor U4623 (N_4623,N_2028,N_1734);
nand U4624 (N_4624,N_534,N_685);
and U4625 (N_4625,N_1167,N_892);
or U4626 (N_4626,N_1939,N_1400);
nand U4627 (N_4627,N_1507,N_126);
or U4628 (N_4628,N_1465,N_1800);
and U4629 (N_4629,N_2246,N_2429);
and U4630 (N_4630,N_2038,N_2312);
or U4631 (N_4631,N_239,N_584);
nand U4632 (N_4632,N_413,N_1775);
nor U4633 (N_4633,N_1305,N_1382);
nand U4634 (N_4634,N_1161,N_1226);
and U4635 (N_4635,N_1099,N_2060);
or U4636 (N_4636,N_1608,N_199);
and U4637 (N_4637,N_21,N_2333);
or U4638 (N_4638,N_2038,N_879);
nor U4639 (N_4639,N_945,N_2132);
and U4640 (N_4640,N_1407,N_549);
nor U4641 (N_4641,N_1708,N_461);
nand U4642 (N_4642,N_2492,N_1240);
or U4643 (N_4643,N_1577,N_2257);
or U4644 (N_4644,N_497,N_575);
nor U4645 (N_4645,N_1786,N_413);
or U4646 (N_4646,N_992,N_2179);
and U4647 (N_4647,N_1912,N_2064);
nor U4648 (N_4648,N_1889,N_2128);
nor U4649 (N_4649,N_1143,N_19);
and U4650 (N_4650,N_2272,N_1650);
nand U4651 (N_4651,N_213,N_881);
or U4652 (N_4652,N_1306,N_778);
nor U4653 (N_4653,N_2158,N_1536);
and U4654 (N_4654,N_79,N_27);
or U4655 (N_4655,N_1194,N_239);
nand U4656 (N_4656,N_324,N_1544);
nand U4657 (N_4657,N_261,N_1332);
nand U4658 (N_4658,N_2314,N_930);
nand U4659 (N_4659,N_2424,N_1498);
nand U4660 (N_4660,N_1139,N_1871);
and U4661 (N_4661,N_2283,N_410);
xor U4662 (N_4662,N_452,N_1073);
nor U4663 (N_4663,N_433,N_1263);
xor U4664 (N_4664,N_2405,N_1456);
or U4665 (N_4665,N_1262,N_1852);
nor U4666 (N_4666,N_2009,N_1844);
and U4667 (N_4667,N_511,N_2456);
nand U4668 (N_4668,N_788,N_1135);
xor U4669 (N_4669,N_1121,N_600);
nor U4670 (N_4670,N_1872,N_860);
nor U4671 (N_4671,N_112,N_1464);
and U4672 (N_4672,N_2299,N_863);
nor U4673 (N_4673,N_1144,N_770);
nand U4674 (N_4674,N_1762,N_2215);
and U4675 (N_4675,N_856,N_1841);
nor U4676 (N_4676,N_755,N_966);
or U4677 (N_4677,N_1342,N_1502);
nor U4678 (N_4678,N_1591,N_613);
or U4679 (N_4679,N_1083,N_1051);
nor U4680 (N_4680,N_2375,N_66);
and U4681 (N_4681,N_324,N_1705);
and U4682 (N_4682,N_2426,N_2109);
nor U4683 (N_4683,N_731,N_123);
or U4684 (N_4684,N_471,N_937);
xor U4685 (N_4685,N_1380,N_238);
or U4686 (N_4686,N_28,N_660);
or U4687 (N_4687,N_2145,N_186);
and U4688 (N_4688,N_1183,N_677);
and U4689 (N_4689,N_159,N_1485);
and U4690 (N_4690,N_1816,N_1695);
and U4691 (N_4691,N_2071,N_1730);
or U4692 (N_4692,N_369,N_1465);
nand U4693 (N_4693,N_2306,N_1991);
or U4694 (N_4694,N_1280,N_382);
nand U4695 (N_4695,N_111,N_434);
nand U4696 (N_4696,N_297,N_1220);
or U4697 (N_4697,N_2401,N_958);
nand U4698 (N_4698,N_1005,N_696);
nand U4699 (N_4699,N_2168,N_1421);
nor U4700 (N_4700,N_104,N_535);
nor U4701 (N_4701,N_59,N_98);
nor U4702 (N_4702,N_1838,N_1400);
nor U4703 (N_4703,N_2005,N_1146);
xor U4704 (N_4704,N_455,N_247);
and U4705 (N_4705,N_22,N_2291);
or U4706 (N_4706,N_78,N_2000);
nand U4707 (N_4707,N_2387,N_1053);
nand U4708 (N_4708,N_172,N_2084);
nor U4709 (N_4709,N_639,N_1590);
and U4710 (N_4710,N_2136,N_2293);
nand U4711 (N_4711,N_806,N_1405);
nand U4712 (N_4712,N_1957,N_1457);
and U4713 (N_4713,N_2389,N_1989);
or U4714 (N_4714,N_74,N_508);
or U4715 (N_4715,N_1490,N_1723);
nor U4716 (N_4716,N_1327,N_1522);
nor U4717 (N_4717,N_88,N_1293);
nand U4718 (N_4718,N_1579,N_414);
and U4719 (N_4719,N_1680,N_2427);
nand U4720 (N_4720,N_849,N_946);
and U4721 (N_4721,N_1497,N_2458);
nor U4722 (N_4722,N_2256,N_761);
nand U4723 (N_4723,N_475,N_1912);
nor U4724 (N_4724,N_749,N_1855);
nor U4725 (N_4725,N_1852,N_571);
and U4726 (N_4726,N_1701,N_509);
and U4727 (N_4727,N_1947,N_1864);
and U4728 (N_4728,N_519,N_820);
nor U4729 (N_4729,N_122,N_254);
nor U4730 (N_4730,N_2167,N_1575);
and U4731 (N_4731,N_1128,N_1116);
and U4732 (N_4732,N_717,N_2010);
nand U4733 (N_4733,N_1084,N_2346);
nand U4734 (N_4734,N_1813,N_446);
nor U4735 (N_4735,N_1101,N_2370);
nor U4736 (N_4736,N_989,N_129);
nor U4737 (N_4737,N_723,N_2155);
or U4738 (N_4738,N_742,N_2130);
and U4739 (N_4739,N_1361,N_1817);
or U4740 (N_4740,N_2350,N_1532);
nand U4741 (N_4741,N_1788,N_1010);
and U4742 (N_4742,N_957,N_830);
or U4743 (N_4743,N_130,N_1616);
and U4744 (N_4744,N_99,N_2005);
nand U4745 (N_4745,N_1032,N_1049);
or U4746 (N_4746,N_157,N_348);
and U4747 (N_4747,N_1019,N_1813);
or U4748 (N_4748,N_1395,N_2236);
nand U4749 (N_4749,N_408,N_949);
nor U4750 (N_4750,N_1842,N_2317);
and U4751 (N_4751,N_214,N_1456);
or U4752 (N_4752,N_1231,N_529);
nand U4753 (N_4753,N_843,N_21);
nor U4754 (N_4754,N_2172,N_1829);
or U4755 (N_4755,N_1535,N_1898);
or U4756 (N_4756,N_287,N_179);
xor U4757 (N_4757,N_332,N_839);
or U4758 (N_4758,N_2148,N_2003);
and U4759 (N_4759,N_1004,N_1726);
or U4760 (N_4760,N_1987,N_1644);
or U4761 (N_4761,N_2169,N_1224);
or U4762 (N_4762,N_1716,N_2491);
nor U4763 (N_4763,N_1064,N_823);
nor U4764 (N_4764,N_1346,N_247);
nand U4765 (N_4765,N_2011,N_1091);
and U4766 (N_4766,N_511,N_1060);
nand U4767 (N_4767,N_2263,N_36);
nor U4768 (N_4768,N_336,N_529);
nor U4769 (N_4769,N_968,N_1509);
and U4770 (N_4770,N_1228,N_1399);
nand U4771 (N_4771,N_769,N_1044);
nand U4772 (N_4772,N_2122,N_514);
nand U4773 (N_4773,N_577,N_1094);
and U4774 (N_4774,N_2362,N_706);
or U4775 (N_4775,N_2163,N_1020);
or U4776 (N_4776,N_1044,N_965);
or U4777 (N_4777,N_1493,N_2191);
nor U4778 (N_4778,N_318,N_380);
and U4779 (N_4779,N_2358,N_494);
or U4780 (N_4780,N_136,N_1740);
nor U4781 (N_4781,N_1002,N_1159);
nor U4782 (N_4782,N_1830,N_257);
nand U4783 (N_4783,N_2469,N_1336);
nor U4784 (N_4784,N_159,N_1966);
and U4785 (N_4785,N_277,N_53);
and U4786 (N_4786,N_1880,N_726);
and U4787 (N_4787,N_1018,N_762);
and U4788 (N_4788,N_1769,N_2146);
nor U4789 (N_4789,N_1788,N_2002);
nor U4790 (N_4790,N_556,N_1435);
or U4791 (N_4791,N_902,N_1756);
or U4792 (N_4792,N_1602,N_2294);
and U4793 (N_4793,N_1425,N_330);
and U4794 (N_4794,N_275,N_2231);
nor U4795 (N_4795,N_1069,N_2498);
or U4796 (N_4796,N_676,N_1977);
and U4797 (N_4797,N_698,N_831);
nor U4798 (N_4798,N_182,N_297);
xor U4799 (N_4799,N_1924,N_2356);
nor U4800 (N_4800,N_2335,N_1745);
or U4801 (N_4801,N_2273,N_1379);
xnor U4802 (N_4802,N_1416,N_18);
nor U4803 (N_4803,N_831,N_1486);
and U4804 (N_4804,N_1369,N_2150);
and U4805 (N_4805,N_2377,N_750);
or U4806 (N_4806,N_58,N_1845);
nor U4807 (N_4807,N_687,N_2094);
nor U4808 (N_4808,N_2157,N_2146);
nor U4809 (N_4809,N_575,N_611);
and U4810 (N_4810,N_1894,N_1164);
nand U4811 (N_4811,N_862,N_1586);
nand U4812 (N_4812,N_575,N_2154);
nand U4813 (N_4813,N_1022,N_1631);
nor U4814 (N_4814,N_964,N_2185);
nand U4815 (N_4815,N_2197,N_2260);
and U4816 (N_4816,N_2172,N_374);
nand U4817 (N_4817,N_704,N_1494);
and U4818 (N_4818,N_1070,N_439);
nand U4819 (N_4819,N_690,N_961);
nor U4820 (N_4820,N_1562,N_458);
nand U4821 (N_4821,N_2398,N_489);
and U4822 (N_4822,N_1683,N_745);
nand U4823 (N_4823,N_2200,N_1860);
and U4824 (N_4824,N_2299,N_1974);
nor U4825 (N_4825,N_20,N_1947);
and U4826 (N_4826,N_114,N_2446);
and U4827 (N_4827,N_695,N_765);
nand U4828 (N_4828,N_969,N_350);
and U4829 (N_4829,N_2079,N_1952);
or U4830 (N_4830,N_1735,N_195);
nand U4831 (N_4831,N_1047,N_198);
nand U4832 (N_4832,N_2421,N_1490);
nor U4833 (N_4833,N_1663,N_1727);
nand U4834 (N_4834,N_885,N_1187);
nand U4835 (N_4835,N_1031,N_2311);
nand U4836 (N_4836,N_1752,N_239);
nor U4837 (N_4837,N_225,N_848);
nor U4838 (N_4838,N_2007,N_641);
nand U4839 (N_4839,N_1429,N_1161);
nand U4840 (N_4840,N_1562,N_1807);
nor U4841 (N_4841,N_1500,N_1875);
or U4842 (N_4842,N_1419,N_1121);
and U4843 (N_4843,N_1558,N_336);
and U4844 (N_4844,N_911,N_313);
nand U4845 (N_4845,N_2423,N_2243);
nand U4846 (N_4846,N_1096,N_366);
nor U4847 (N_4847,N_1051,N_1232);
nand U4848 (N_4848,N_1324,N_2468);
or U4849 (N_4849,N_1806,N_1868);
nor U4850 (N_4850,N_2389,N_7);
and U4851 (N_4851,N_1608,N_2499);
nor U4852 (N_4852,N_662,N_113);
nor U4853 (N_4853,N_1673,N_921);
nor U4854 (N_4854,N_84,N_2433);
nand U4855 (N_4855,N_79,N_1602);
and U4856 (N_4856,N_1175,N_1113);
or U4857 (N_4857,N_1237,N_1549);
and U4858 (N_4858,N_149,N_2240);
nor U4859 (N_4859,N_261,N_612);
nand U4860 (N_4860,N_31,N_1042);
and U4861 (N_4861,N_2235,N_624);
nand U4862 (N_4862,N_1257,N_1003);
xnor U4863 (N_4863,N_2033,N_1777);
nor U4864 (N_4864,N_1922,N_1289);
nand U4865 (N_4865,N_1899,N_1401);
nand U4866 (N_4866,N_1365,N_820);
nor U4867 (N_4867,N_12,N_619);
and U4868 (N_4868,N_1700,N_1887);
nand U4869 (N_4869,N_1501,N_1939);
nor U4870 (N_4870,N_550,N_963);
and U4871 (N_4871,N_2437,N_847);
nand U4872 (N_4872,N_2201,N_1831);
and U4873 (N_4873,N_1521,N_35);
or U4874 (N_4874,N_621,N_1295);
or U4875 (N_4875,N_903,N_24);
and U4876 (N_4876,N_2371,N_345);
nor U4877 (N_4877,N_1406,N_46);
and U4878 (N_4878,N_993,N_1197);
nand U4879 (N_4879,N_699,N_1247);
nand U4880 (N_4880,N_44,N_793);
nand U4881 (N_4881,N_1767,N_2);
or U4882 (N_4882,N_2472,N_1804);
nand U4883 (N_4883,N_219,N_1969);
nand U4884 (N_4884,N_1321,N_2040);
nand U4885 (N_4885,N_247,N_1232);
nor U4886 (N_4886,N_2426,N_319);
nor U4887 (N_4887,N_516,N_409);
nor U4888 (N_4888,N_759,N_2457);
or U4889 (N_4889,N_1150,N_1738);
nand U4890 (N_4890,N_417,N_1109);
or U4891 (N_4891,N_386,N_2300);
nand U4892 (N_4892,N_2142,N_378);
or U4893 (N_4893,N_164,N_287);
nor U4894 (N_4894,N_1265,N_2269);
or U4895 (N_4895,N_697,N_404);
or U4896 (N_4896,N_844,N_502);
nor U4897 (N_4897,N_1889,N_1497);
or U4898 (N_4898,N_24,N_889);
and U4899 (N_4899,N_2067,N_1361);
nand U4900 (N_4900,N_678,N_829);
nand U4901 (N_4901,N_265,N_880);
or U4902 (N_4902,N_1389,N_815);
or U4903 (N_4903,N_1252,N_27);
or U4904 (N_4904,N_1359,N_458);
and U4905 (N_4905,N_1555,N_2415);
nand U4906 (N_4906,N_1432,N_1108);
or U4907 (N_4907,N_1191,N_1075);
and U4908 (N_4908,N_534,N_1912);
nand U4909 (N_4909,N_1464,N_9);
and U4910 (N_4910,N_2400,N_535);
nand U4911 (N_4911,N_330,N_1201);
and U4912 (N_4912,N_178,N_146);
or U4913 (N_4913,N_1745,N_1671);
nor U4914 (N_4914,N_795,N_290);
and U4915 (N_4915,N_1747,N_1270);
or U4916 (N_4916,N_1583,N_1106);
or U4917 (N_4917,N_429,N_2136);
and U4918 (N_4918,N_2321,N_503);
or U4919 (N_4919,N_998,N_18);
nand U4920 (N_4920,N_554,N_2318);
and U4921 (N_4921,N_538,N_1036);
nand U4922 (N_4922,N_709,N_896);
nand U4923 (N_4923,N_965,N_12);
or U4924 (N_4924,N_331,N_2019);
nor U4925 (N_4925,N_931,N_731);
nand U4926 (N_4926,N_1975,N_1793);
or U4927 (N_4927,N_2011,N_1591);
and U4928 (N_4928,N_1026,N_1214);
xnor U4929 (N_4929,N_148,N_2274);
nand U4930 (N_4930,N_1009,N_2257);
and U4931 (N_4931,N_1520,N_1698);
and U4932 (N_4932,N_2199,N_147);
nor U4933 (N_4933,N_914,N_2431);
nor U4934 (N_4934,N_2254,N_1831);
and U4935 (N_4935,N_830,N_820);
or U4936 (N_4936,N_1440,N_916);
and U4937 (N_4937,N_1512,N_1238);
nor U4938 (N_4938,N_367,N_260);
or U4939 (N_4939,N_2452,N_1682);
or U4940 (N_4940,N_2440,N_15);
and U4941 (N_4941,N_29,N_1547);
nand U4942 (N_4942,N_1795,N_184);
or U4943 (N_4943,N_1997,N_2287);
nor U4944 (N_4944,N_888,N_925);
or U4945 (N_4945,N_1059,N_1621);
nor U4946 (N_4946,N_679,N_834);
nand U4947 (N_4947,N_1426,N_650);
xnor U4948 (N_4948,N_601,N_809);
nand U4949 (N_4949,N_2170,N_2468);
nor U4950 (N_4950,N_833,N_632);
nor U4951 (N_4951,N_406,N_1883);
or U4952 (N_4952,N_1369,N_1009);
or U4953 (N_4953,N_605,N_1968);
nand U4954 (N_4954,N_1767,N_2428);
nand U4955 (N_4955,N_2420,N_2395);
nor U4956 (N_4956,N_1413,N_246);
and U4957 (N_4957,N_1781,N_1069);
or U4958 (N_4958,N_2215,N_2150);
or U4959 (N_4959,N_1202,N_325);
nand U4960 (N_4960,N_2111,N_579);
nor U4961 (N_4961,N_2044,N_1507);
nand U4962 (N_4962,N_1440,N_951);
or U4963 (N_4963,N_854,N_535);
nor U4964 (N_4964,N_2402,N_1367);
nand U4965 (N_4965,N_343,N_1203);
and U4966 (N_4966,N_416,N_182);
nor U4967 (N_4967,N_1316,N_2319);
and U4968 (N_4968,N_2070,N_21);
and U4969 (N_4969,N_1216,N_920);
or U4970 (N_4970,N_1851,N_1712);
nand U4971 (N_4971,N_258,N_2355);
or U4972 (N_4972,N_2048,N_998);
and U4973 (N_4973,N_1188,N_45);
nor U4974 (N_4974,N_975,N_621);
nor U4975 (N_4975,N_2069,N_18);
or U4976 (N_4976,N_2260,N_275);
nor U4977 (N_4977,N_793,N_1143);
or U4978 (N_4978,N_945,N_1576);
nand U4979 (N_4979,N_130,N_1331);
nor U4980 (N_4980,N_2470,N_681);
or U4981 (N_4981,N_1074,N_1929);
nor U4982 (N_4982,N_1958,N_970);
or U4983 (N_4983,N_1956,N_2101);
nor U4984 (N_4984,N_126,N_1538);
and U4985 (N_4985,N_956,N_1993);
nand U4986 (N_4986,N_1093,N_2369);
and U4987 (N_4987,N_1914,N_1852);
nand U4988 (N_4988,N_751,N_1962);
or U4989 (N_4989,N_1714,N_2211);
nor U4990 (N_4990,N_1658,N_1094);
nand U4991 (N_4991,N_680,N_1929);
nor U4992 (N_4992,N_1441,N_1563);
nor U4993 (N_4993,N_645,N_67);
and U4994 (N_4994,N_2337,N_124);
nand U4995 (N_4995,N_1094,N_1333);
or U4996 (N_4996,N_2354,N_708);
nand U4997 (N_4997,N_681,N_2454);
and U4998 (N_4998,N_1595,N_283);
and U4999 (N_4999,N_2006,N_199);
nand UO_0 (O_0,N_3171,N_4596);
nand UO_1 (O_1,N_3945,N_3091);
nand UO_2 (O_2,N_3514,N_3050);
and UO_3 (O_3,N_4049,N_4822);
or UO_4 (O_4,N_3541,N_3684);
nand UO_5 (O_5,N_3276,N_3734);
nor UO_6 (O_6,N_2640,N_4437);
and UO_7 (O_7,N_4329,N_3052);
or UO_8 (O_8,N_3495,N_2958);
xnor UO_9 (O_9,N_4074,N_2939);
nand UO_10 (O_10,N_4245,N_2604);
or UO_11 (O_11,N_2669,N_4498);
nor UO_12 (O_12,N_4382,N_3367);
and UO_13 (O_13,N_3706,N_3278);
and UO_14 (O_14,N_3529,N_3836);
or UO_15 (O_15,N_3969,N_3326);
nand UO_16 (O_16,N_2605,N_3831);
nand UO_17 (O_17,N_3697,N_3731);
nand UO_18 (O_18,N_4628,N_4584);
nand UO_19 (O_19,N_4018,N_4722);
nand UO_20 (O_20,N_2530,N_4930);
nand UO_21 (O_21,N_3334,N_3329);
or UO_22 (O_22,N_2700,N_4423);
or UO_23 (O_23,N_2534,N_2914);
xor UO_24 (O_24,N_4903,N_3949);
nor UO_25 (O_25,N_3019,N_3549);
or UO_26 (O_26,N_3436,N_3428);
nand UO_27 (O_27,N_2525,N_2957);
and UO_28 (O_28,N_2591,N_4269);
or UO_29 (O_29,N_3375,N_3333);
nand UO_30 (O_30,N_3736,N_4823);
nand UO_31 (O_31,N_2754,N_4631);
nand UO_32 (O_32,N_3711,N_2661);
nand UO_33 (O_33,N_3958,N_4270);
nand UO_34 (O_34,N_4360,N_3552);
nor UO_35 (O_35,N_3109,N_4614);
and UO_36 (O_36,N_2675,N_2711);
nor UO_37 (O_37,N_4192,N_4812);
nor UO_38 (O_38,N_4072,N_3092);
and UO_39 (O_39,N_3628,N_4237);
and UO_40 (O_40,N_3718,N_3497);
nand UO_41 (O_41,N_4629,N_2730);
and UO_42 (O_42,N_3556,N_4779);
or UO_43 (O_43,N_4483,N_2896);
nor UO_44 (O_44,N_3064,N_4493);
nand UO_45 (O_45,N_4447,N_4386);
nor UO_46 (O_46,N_3173,N_3139);
or UO_47 (O_47,N_3806,N_2653);
nand UO_48 (O_48,N_3111,N_3685);
or UO_49 (O_49,N_2856,N_3328);
nor UO_50 (O_50,N_3744,N_4817);
nand UO_51 (O_51,N_2523,N_3284);
nor UO_52 (O_52,N_3304,N_4457);
nand UO_53 (O_53,N_3939,N_2616);
nor UO_54 (O_54,N_3724,N_3924);
or UO_55 (O_55,N_3838,N_2581);
or UO_56 (O_56,N_3441,N_2571);
and UO_57 (O_57,N_2943,N_2876);
and UO_58 (O_58,N_3670,N_3872);
and UO_59 (O_59,N_3272,N_3601);
nor UO_60 (O_60,N_4992,N_2909);
or UO_61 (O_61,N_4525,N_3805);
nor UO_62 (O_62,N_4798,N_3702);
and UO_63 (O_63,N_2771,N_3383);
nor UO_64 (O_64,N_2644,N_3423);
nand UO_65 (O_65,N_4069,N_3876);
or UO_66 (O_66,N_4485,N_3964);
nor UO_67 (O_67,N_3235,N_3767);
and UO_68 (O_68,N_4233,N_3770);
nor UO_69 (O_69,N_3237,N_4376);
nor UO_70 (O_70,N_4653,N_3330);
or UO_71 (O_71,N_3327,N_3879);
nand UO_72 (O_72,N_4199,N_2748);
and UO_73 (O_73,N_4334,N_4809);
and UO_74 (O_74,N_2972,N_3234);
and UO_75 (O_75,N_4048,N_2728);
and UO_76 (O_76,N_3152,N_4212);
and UO_77 (O_77,N_3444,N_4124);
or UO_78 (O_78,N_3520,N_3022);
and UO_79 (O_79,N_2994,N_3786);
nand UO_80 (O_80,N_2531,N_3277);
nor UO_81 (O_81,N_4396,N_4730);
nor UO_82 (O_82,N_2965,N_3615);
nand UO_83 (O_83,N_4040,N_3506);
or UO_84 (O_84,N_3970,N_4324);
nor UO_85 (O_85,N_3438,N_4636);
or UO_86 (O_86,N_4164,N_4339);
and UO_87 (O_87,N_3322,N_3792);
nor UO_88 (O_88,N_4102,N_3430);
nand UO_89 (O_89,N_4751,N_3909);
nor UO_90 (O_90,N_3151,N_4935);
or UO_91 (O_91,N_2982,N_4658);
and UO_92 (O_92,N_3259,N_2809);
nand UO_93 (O_93,N_4737,N_3948);
nand UO_94 (O_94,N_3848,N_4435);
and UO_95 (O_95,N_4073,N_3509);
nand UO_96 (O_96,N_3940,N_4469);
and UO_97 (O_97,N_4926,N_4666);
and UO_98 (O_98,N_4466,N_2774);
nand UO_99 (O_99,N_2920,N_3955);
and UO_100 (O_100,N_4977,N_2814);
nand UO_101 (O_101,N_3693,N_3485);
nor UO_102 (O_102,N_3369,N_2794);
nor UO_103 (O_103,N_3599,N_4937);
nor UO_104 (O_104,N_4108,N_4782);
or UO_105 (O_105,N_2567,N_2826);
nor UO_106 (O_106,N_3493,N_4076);
and UO_107 (O_107,N_4696,N_3500);
nand UO_108 (O_108,N_2803,N_4180);
or UO_109 (O_109,N_3976,N_3289);
nand UO_110 (O_110,N_3522,N_4016);
nand UO_111 (O_111,N_3737,N_4825);
nor UO_112 (O_112,N_4125,N_4727);
and UO_113 (O_113,N_4492,N_2975);
and UO_114 (O_114,N_4515,N_4802);
or UO_115 (O_115,N_2690,N_4384);
nor UO_116 (O_116,N_4537,N_3385);
or UO_117 (O_117,N_3070,N_4609);
nor UO_118 (O_118,N_4445,N_4008);
nor UO_119 (O_119,N_3584,N_4624);
nor UO_120 (O_120,N_4030,N_3563);
nand UO_121 (O_121,N_4577,N_3721);
or UO_122 (O_122,N_2541,N_2659);
nor UO_123 (O_123,N_3892,N_4507);
or UO_124 (O_124,N_3621,N_4479);
xnor UO_125 (O_125,N_2772,N_4972);
nor UO_126 (O_126,N_3210,N_2879);
nand UO_127 (O_127,N_2938,N_3672);
or UO_128 (O_128,N_4551,N_4309);
and UO_129 (O_129,N_2822,N_4229);
and UO_130 (O_130,N_3465,N_2764);
or UO_131 (O_131,N_4708,N_3480);
or UO_132 (O_132,N_2688,N_3148);
or UO_133 (O_133,N_3147,N_2658);
nor UO_134 (O_134,N_3695,N_3413);
nor UO_135 (O_135,N_2786,N_4605);
nand UO_136 (O_136,N_4758,N_4379);
nand UO_137 (O_137,N_4784,N_4228);
nor UO_138 (O_138,N_2519,N_4442);
nor UO_139 (O_139,N_3888,N_4406);
nand UO_140 (O_140,N_4713,N_3987);
nor UO_141 (O_141,N_3103,N_4869);
or UO_142 (O_142,N_2766,N_4209);
nand UO_143 (O_143,N_4512,N_3985);
nand UO_144 (O_144,N_3454,N_3227);
and UO_145 (O_145,N_3997,N_3342);
and UO_146 (O_146,N_4807,N_4385);
nand UO_147 (O_147,N_2716,N_4800);
nor UO_148 (O_148,N_3132,N_3477);
nand UO_149 (O_149,N_4095,N_4213);
nand UO_150 (O_150,N_3098,N_2639);
nand UO_151 (O_151,N_3352,N_3280);
or UO_152 (O_152,N_4509,N_4219);
nand UO_153 (O_153,N_4189,N_4319);
nand UO_154 (O_154,N_4390,N_3439);
or UO_155 (O_155,N_4436,N_3686);
nor UO_156 (O_156,N_2736,N_4608);
nor UO_157 (O_157,N_3817,N_3081);
nand UO_158 (O_158,N_2626,N_3143);
and UO_159 (O_159,N_4548,N_4855);
and UO_160 (O_160,N_3396,N_2955);
or UO_161 (O_161,N_3828,N_3663);
or UO_162 (O_162,N_4725,N_4909);
nand UO_163 (O_163,N_4726,N_3411);
and UO_164 (O_164,N_3101,N_4299);
nor UO_165 (O_165,N_3800,N_2870);
nor UO_166 (O_166,N_2990,N_4461);
or UO_167 (O_167,N_2635,N_4671);
nand UO_168 (O_168,N_3133,N_4304);
or UO_169 (O_169,N_2598,N_4585);
and UO_170 (O_170,N_3978,N_2970);
and UO_171 (O_171,N_4752,N_4399);
and UO_172 (O_172,N_3209,N_3742);
or UO_173 (O_173,N_2783,N_3798);
or UO_174 (O_174,N_3971,N_4982);
and UO_175 (O_175,N_4721,N_4889);
or UO_176 (O_176,N_2756,N_3638);
or UO_177 (O_177,N_2599,N_4787);
or UO_178 (O_178,N_4774,N_2801);
or UO_179 (O_179,N_2731,N_2699);
nor UO_180 (O_180,N_4337,N_4128);
or UO_181 (O_181,N_4011,N_3636);
nor UO_182 (O_182,N_3521,N_3899);
or UO_183 (O_183,N_4613,N_4026);
and UO_184 (O_184,N_4500,N_3114);
or UO_185 (O_185,N_2828,N_3409);
nand UO_186 (O_186,N_4149,N_4842);
or UO_187 (O_187,N_3633,N_3725);
and UO_188 (O_188,N_4964,N_4733);
and UO_189 (O_189,N_2632,N_3799);
or UO_190 (O_190,N_2735,N_4181);
nor UO_191 (O_191,N_3292,N_2692);
nand UO_192 (O_192,N_4312,N_4815);
and UO_193 (O_193,N_2670,N_4388);
nand UO_194 (O_194,N_2703,N_4021);
nand UO_195 (O_195,N_3168,N_2586);
or UO_196 (O_196,N_4345,N_3476);
and UO_197 (O_197,N_3285,N_4068);
nor UO_198 (O_198,N_4531,N_4646);
or UO_199 (O_199,N_3629,N_4600);
nand UO_200 (O_200,N_3710,N_3311);
nand UO_201 (O_201,N_3657,N_2877);
or UO_202 (O_202,N_2695,N_4250);
or UO_203 (O_203,N_2974,N_3565);
or UO_204 (O_204,N_3947,N_4610);
or UO_205 (O_205,N_3667,N_4182);
nor UO_206 (O_206,N_4452,N_3534);
nand UO_207 (O_207,N_4351,N_4174);
or UO_208 (O_208,N_3804,N_3242);
and UO_209 (O_209,N_4491,N_2588);
nor UO_210 (O_210,N_3550,N_3401);
and UO_211 (O_211,N_4732,N_3808);
nor UO_212 (O_212,N_2536,N_3716);
nand UO_213 (O_213,N_3769,N_2682);
nor UO_214 (O_214,N_4620,N_3747);
nor UO_215 (O_215,N_3275,N_3540);
or UO_216 (O_216,N_3780,N_3075);
nor UO_217 (O_217,N_3248,N_4326);
nand UO_218 (O_218,N_3190,N_4583);
nor UO_219 (O_219,N_3037,N_4983);
nor UO_220 (O_220,N_4440,N_2839);
nand UO_221 (O_221,N_4023,N_3232);
and UO_222 (O_222,N_3475,N_3124);
nand UO_223 (O_223,N_4427,N_4845);
nor UO_224 (O_224,N_3491,N_3172);
or UO_225 (O_225,N_4973,N_3354);
and UO_226 (O_226,N_2945,N_3632);
nor UO_227 (O_227,N_3001,N_3612);
or UO_228 (O_228,N_4041,N_2899);
or UO_229 (O_229,N_4874,N_3863);
nor UO_230 (O_230,N_3160,N_4619);
nor UO_231 (O_231,N_4790,N_3031);
and UO_232 (O_232,N_3451,N_2935);
nor UO_233 (O_233,N_2627,N_2951);
nor UO_234 (O_234,N_4006,N_3047);
nor UO_235 (O_235,N_4718,N_4882);
and UO_236 (O_236,N_3392,N_3739);
nor UO_237 (O_237,N_4739,N_3505);
nor UO_238 (O_238,N_3252,N_4070);
xnor UO_239 (O_239,N_4913,N_3363);
and UO_240 (O_240,N_4521,N_4719);
and UO_241 (O_241,N_4321,N_2953);
or UO_242 (O_242,N_3538,N_3816);
and UO_243 (O_243,N_3347,N_2643);
nor UO_244 (O_244,N_3366,N_4301);
nor UO_245 (O_245,N_4150,N_2727);
or UO_246 (O_246,N_3754,N_4888);
or UO_247 (O_247,N_2807,N_3034);
nand UO_248 (O_248,N_3027,N_3373);
or UO_249 (O_249,N_4954,N_3426);
or UO_250 (O_250,N_2966,N_2552);
and UO_251 (O_251,N_3417,N_3776);
nor UO_252 (O_252,N_4433,N_4091);
nor UO_253 (O_253,N_2816,N_4644);
nand UO_254 (O_254,N_3349,N_4996);
nand UO_255 (O_255,N_3241,N_3291);
nand UO_256 (O_256,N_3331,N_4706);
nor UO_257 (O_257,N_3680,N_4821);
nand UO_258 (O_258,N_2800,N_4539);
or UO_259 (O_259,N_4035,N_3025);
and UO_260 (O_260,N_2777,N_2765);
and UO_261 (O_261,N_3040,N_4603);
and UO_262 (O_262,N_4872,N_2743);
nor UO_263 (O_263,N_4772,N_3975);
and UO_264 (O_264,N_2768,N_3518);
and UO_265 (O_265,N_4463,N_4311);
xor UO_266 (O_266,N_4488,N_4538);
nand UO_267 (O_267,N_2933,N_3033);
or UO_268 (O_268,N_3170,N_3704);
nand UO_269 (O_269,N_2508,N_4728);
xor UO_270 (O_270,N_3182,N_2740);
nand UO_271 (O_271,N_2824,N_3611);
and UO_272 (O_272,N_4879,N_2845);
nand UO_273 (O_273,N_4357,N_4478);
nand UO_274 (O_274,N_2621,N_2949);
and UO_275 (O_275,N_4847,N_2517);
and UO_276 (O_276,N_3760,N_2901);
nor UO_277 (O_277,N_2742,N_2647);
nor UO_278 (O_278,N_4931,N_4867);
xor UO_279 (O_279,N_4940,N_4673);
and UO_280 (O_280,N_4327,N_4484);
or UO_281 (O_281,N_3183,N_3698);
nand UO_282 (O_282,N_2893,N_4716);
xor UO_283 (O_283,N_3462,N_2545);
or UO_284 (O_284,N_3346,N_2645);
nand UO_285 (O_285,N_4118,N_4681);
or UO_286 (O_286,N_2996,N_3935);
and UO_287 (O_287,N_2813,N_3532);
and UO_288 (O_288,N_2606,N_4434);
and UO_289 (O_289,N_3307,N_4459);
and UO_290 (O_290,N_3335,N_3957);
nor UO_291 (O_291,N_2533,N_4777);
and UO_292 (O_292,N_4261,N_2865);
nor UO_293 (O_293,N_2565,N_4204);
or UO_294 (O_294,N_3951,N_2846);
or UO_295 (O_295,N_3913,N_4276);
and UO_296 (O_296,N_4296,N_3178);
nand UO_297 (O_297,N_2747,N_2638);
and UO_298 (O_298,N_3977,N_3893);
nor UO_299 (O_299,N_3577,N_2821);
nor UO_300 (O_300,N_3842,N_4195);
or UO_301 (O_301,N_2782,N_3448);
and UO_302 (O_302,N_4141,N_4402);
nand UO_303 (O_303,N_2827,N_2880);
nand UO_304 (O_304,N_4896,N_3690);
nand UO_305 (O_305,N_2612,N_4598);
xor UO_306 (O_306,N_3791,N_3847);
nand UO_307 (O_307,N_4542,N_4829);
and UO_308 (O_308,N_4841,N_3627);
or UO_309 (O_309,N_2584,N_3492);
or UO_310 (O_310,N_3048,N_4064);
nand UO_311 (O_311,N_2954,N_4883);
nor UO_312 (O_312,N_4093,N_2564);
and UO_313 (O_313,N_4138,N_4205);
and UO_314 (O_314,N_4639,N_2890);
nand UO_315 (O_315,N_3758,N_4650);
and UO_316 (O_316,N_3581,N_4578);
nor UO_317 (O_317,N_3635,N_4374);
or UO_318 (O_318,N_3717,N_4832);
or UO_319 (O_319,N_2734,N_3282);
and UO_320 (O_320,N_3823,N_4453);
nand UO_321 (O_321,N_4944,N_4203);
or UO_322 (O_322,N_3059,N_2998);
nand UO_323 (O_323,N_4114,N_3416);
and UO_324 (O_324,N_3539,N_2762);
and UO_325 (O_325,N_4306,N_4098);
nand UO_326 (O_326,N_3887,N_4796);
and UO_327 (O_327,N_3658,N_3554);
or UO_328 (O_328,N_3772,N_3267);
nor UO_329 (O_329,N_2857,N_4688);
nand UO_330 (O_330,N_3169,N_4545);
or UO_331 (O_331,N_4316,N_4924);
nor UO_332 (O_332,N_3517,N_3993);
nor UO_333 (O_333,N_3202,N_2712);
or UO_334 (O_334,N_4687,N_2662);
nor UO_335 (O_335,N_3513,N_4272);
nand UO_336 (O_336,N_4770,N_4172);
and UO_337 (O_337,N_4569,N_4559);
and UO_338 (O_338,N_3785,N_4103);
or UO_339 (O_339,N_3136,N_4571);
nor UO_340 (O_340,N_3525,N_3239);
nor UO_341 (O_341,N_3231,N_4450);
and UO_342 (O_342,N_4389,N_3371);
nor UO_343 (O_343,N_4377,N_3162);
and UO_344 (O_344,N_4470,N_4277);
and UO_345 (O_345,N_4604,N_3345);
nand UO_346 (O_346,N_3605,N_4891);
and UO_347 (O_347,N_4046,N_4028);
or UO_348 (O_348,N_3021,N_3986);
xnor UO_349 (O_349,N_3078,N_4135);
nand UO_350 (O_350,N_4952,N_3212);
or UO_351 (O_351,N_4259,N_2554);
and UO_352 (O_352,N_2528,N_3972);
nor UO_353 (O_353,N_3286,N_4503);
and UO_354 (O_354,N_2710,N_3967);
nor UO_355 (O_355,N_3261,N_4519);
nand UO_356 (O_356,N_3138,N_2843);
nand UO_357 (O_357,N_2634,N_2529);
and UO_358 (O_358,N_4425,N_3720);
nand UO_359 (O_359,N_3603,N_2849);
and UO_360 (O_360,N_4414,N_4499);
or UO_361 (O_361,N_2925,N_4273);
nand UO_362 (O_362,N_3589,N_2904);
nor UO_363 (O_363,N_4993,N_2737);
nand UO_364 (O_364,N_3236,N_4282);
nand UO_365 (O_365,N_3377,N_2684);
nand UO_366 (O_366,N_2929,N_4731);
and UO_367 (O_367,N_3167,N_4200);
and UO_368 (O_368,N_4980,N_4567);
and UO_369 (O_369,N_2641,N_4570);
nor UO_370 (O_370,N_4179,N_4133);
nand UO_371 (O_371,N_3533,N_3526);
or UO_372 (O_372,N_3898,N_2580);
nand UO_373 (O_373,N_3901,N_3507);
and UO_374 (O_374,N_3499,N_2964);
and UO_375 (O_375,N_4085,N_4970);
and UO_376 (O_376,N_2576,N_3422);
and UO_377 (O_377,N_3719,N_3889);
nand UO_378 (O_378,N_4201,N_2946);
and UO_379 (O_379,N_2568,N_2993);
or UO_380 (O_380,N_4533,N_2997);
or UO_381 (O_381,N_4094,N_4136);
nand UO_382 (O_382,N_2991,N_2798);
nand UO_383 (O_383,N_4249,N_2587);
nor UO_384 (O_384,N_3314,N_4058);
nand UO_385 (O_385,N_3131,N_2713);
nand UO_386 (O_386,N_3826,N_4840);
nand UO_387 (O_387,N_2574,N_4220);
or UO_388 (O_388,N_3145,N_4256);
nand UO_389 (O_389,N_4831,N_3260);
nand UO_390 (O_390,N_3648,N_3157);
nand UO_391 (O_391,N_3896,N_4053);
and UO_392 (O_392,N_4348,N_3994);
or UO_393 (O_393,N_3923,N_3664);
or UO_394 (O_394,N_4335,N_4347);
or UO_395 (O_395,N_2570,N_4514);
nand UO_396 (O_396,N_4984,N_3279);
and UO_397 (O_397,N_4080,N_2931);
nand UO_398 (O_398,N_2757,N_3624);
or UO_399 (O_399,N_4919,N_2971);
nand UO_400 (O_400,N_2791,N_3460);
nor UO_401 (O_401,N_3966,N_2898);
or UO_402 (O_402,N_2646,N_3176);
nand UO_403 (O_403,N_3156,N_3435);
nand UO_404 (O_404,N_4362,N_2511);
nor UO_405 (O_405,N_4057,N_4218);
nor UO_406 (O_406,N_2524,N_4543);
nor UO_407 (O_407,N_4419,N_4670);
and UO_408 (O_408,N_4079,N_4071);
nor UO_409 (O_409,N_2749,N_4750);
nand UO_410 (O_410,N_4285,N_2793);
or UO_411 (O_411,N_3812,N_4353);
nor UO_412 (O_412,N_4735,N_4227);
nand UO_413 (O_413,N_3308,N_3223);
nand UO_414 (O_414,N_2797,N_2614);
or UO_415 (O_415,N_4900,N_4960);
and UO_416 (O_416,N_3208,N_3412);
nor UO_417 (O_417,N_4412,N_4432);
and UO_418 (O_418,N_3445,N_3274);
nand UO_419 (O_419,N_4936,N_3634);
nor UO_420 (O_420,N_4856,N_3447);
nor UO_421 (O_421,N_4594,N_3273);
or UO_422 (O_422,N_4691,N_4467);
or UO_423 (O_423,N_4404,N_2751);
nand UO_424 (O_424,N_3829,N_2752);
nand UO_425 (O_425,N_3787,N_3989);
or UO_426 (O_426,N_4859,N_4176);
nand UO_427 (O_427,N_4592,N_3035);
or UO_428 (O_428,N_3897,N_4003);
nand UO_429 (O_429,N_4651,N_3946);
nor UO_430 (O_430,N_2812,N_3933);
and UO_431 (O_431,N_3655,N_4611);
nor UO_432 (O_432,N_2891,N_3580);
nor UO_433 (O_433,N_2940,N_2858);
or UO_434 (O_434,N_2582,N_4037);
nor UO_435 (O_435,N_2522,N_3922);
nand UO_436 (O_436,N_2947,N_3123);
nand UO_437 (O_437,N_4814,N_4283);
and UO_438 (O_438,N_3247,N_4660);
or UO_439 (O_439,N_2607,N_2629);
or UO_440 (O_440,N_2981,N_2932);
xor UO_441 (O_441,N_4151,N_2948);
nor UO_442 (O_442,N_3567,N_4460);
nand UO_443 (O_443,N_4065,N_4866);
nor UO_444 (O_444,N_3457,N_2985);
and UO_445 (O_445,N_4067,N_3609);
nand UO_446 (O_446,N_3159,N_3708);
nor UO_447 (O_447,N_3974,N_3061);
nand UO_448 (O_448,N_3194,N_3877);
and UO_449 (O_449,N_4210,N_4169);
and UO_450 (O_450,N_3668,N_3305);
or UO_451 (O_451,N_3535,N_3592);
nor UO_452 (O_452,N_3613,N_3918);
or UO_453 (O_453,N_4284,N_4589);
or UO_454 (O_454,N_3574,N_3116);
nand UO_455 (O_455,N_4838,N_3659);
nor UO_456 (O_456,N_4966,N_4949);
and UO_457 (O_457,N_3783,N_3961);
nor UO_458 (O_458,N_2916,N_4107);
nand UO_459 (O_459,N_2770,N_4043);
nand UO_460 (O_460,N_3134,N_3727);
nor UO_461 (O_461,N_4749,N_4981);
and UO_462 (O_462,N_3729,N_3590);
and UO_463 (O_463,N_3343,N_3559);
or UO_464 (O_464,N_3784,N_4242);
nand UO_465 (O_465,N_3819,N_3246);
nor UO_466 (O_466,N_3009,N_4723);
xor UO_467 (O_467,N_2611,N_2962);
nor UO_468 (O_468,N_4933,N_2815);
nand UO_469 (O_469,N_3297,N_3295);
nor UO_470 (O_470,N_3937,N_3496);
nor UO_471 (O_471,N_4595,N_3980);
nor UO_472 (O_472,N_4623,N_3391);
nand UO_473 (O_473,N_4986,N_2830);
nand UO_474 (O_474,N_3288,N_3068);
and UO_475 (O_475,N_4950,N_4894);
nor UO_476 (O_476,N_3104,N_3527);
and UO_477 (O_477,N_4975,N_3867);
and UO_478 (O_478,N_4305,N_4476);
and UO_479 (O_479,N_3748,N_4532);
nand UO_480 (O_480,N_3233,N_3861);
and UO_481 (O_481,N_4474,N_4364);
and UO_482 (O_482,N_3900,N_4702);
and UO_483 (O_483,N_3757,N_4363);
or UO_484 (O_484,N_3516,N_4914);
nor UO_485 (O_485,N_4078,N_3703);
nand UO_486 (O_486,N_3467,N_3607);
and UO_487 (O_487,N_2521,N_4689);
nand UO_488 (O_488,N_4475,N_4487);
nor UO_489 (O_489,N_2504,N_3920);
or UO_490 (O_490,N_3389,N_3979);
and UO_491 (O_491,N_4446,N_4325);
nor UO_492 (O_492,N_4116,N_4618);
nor UO_493 (O_493,N_4553,N_4763);
nor UO_494 (O_494,N_3884,N_3835);
or UO_495 (O_495,N_2701,N_3573);
nor UO_496 (O_496,N_3395,N_3618);
nand UO_497 (O_497,N_2874,N_2557);
nor UO_498 (O_498,N_2633,N_2883);
and UO_499 (O_499,N_3337,N_4123);
nor UO_500 (O_500,N_2719,N_4747);
and UO_501 (O_501,N_4052,N_4775);
and UO_502 (O_502,N_3929,N_4505);
and UO_503 (O_503,N_4835,N_4441);
or UO_504 (O_504,N_4186,N_4171);
and UO_505 (O_505,N_2601,N_4917);
and UO_506 (O_506,N_3818,N_4111);
and UO_507 (O_507,N_3562,N_4607);
and UO_508 (O_508,N_3281,N_4698);
nand UO_509 (O_509,N_3000,N_4254);
or UO_510 (O_510,N_4232,N_3524);
or UO_511 (O_511,N_4907,N_3917);
nand UO_512 (O_512,N_2745,N_4428);
nor UO_513 (O_513,N_4398,N_3038);
nand UO_514 (O_514,N_4554,N_4871);
nor UO_515 (O_515,N_4014,N_4808);
nor UO_516 (O_516,N_3866,N_4417);
nand UO_517 (O_517,N_3859,N_4050);
and UO_518 (O_518,N_4664,N_2868);
nand UO_519 (O_519,N_2767,N_2831);
and UO_520 (O_520,N_4806,N_4144);
or UO_521 (O_521,N_2510,N_4255);
and UO_522 (O_522,N_4648,N_2763);
or UO_523 (O_523,N_4634,N_3225);
nand UO_524 (O_524,N_4632,N_4185);
and UO_525 (O_525,N_4579,N_4511);
nand UO_526 (O_526,N_4240,N_3270);
nor UO_527 (O_527,N_2577,N_4580);
nor UO_528 (O_528,N_3403,N_4911);
or UO_529 (O_529,N_3017,N_4679);
nor UO_530 (O_530,N_3365,N_3135);
nor UO_531 (O_531,N_4686,N_3560);
or UO_532 (O_532,N_2912,N_2895);
and UO_533 (O_533,N_4694,N_3732);
and UO_534 (O_534,N_2622,N_4313);
nand UO_535 (O_535,N_2844,N_3666);
and UO_536 (O_536,N_3582,N_3355);
or UO_537 (O_537,N_2671,N_2718);
nor UO_538 (O_538,N_3478,N_4015);
nand UO_539 (O_539,N_3243,N_2702);
or UO_540 (O_540,N_4797,N_3661);
nand UO_541 (O_541,N_3121,N_3046);
nor UO_542 (O_542,N_4925,N_2885);
or UO_543 (O_543,N_3086,N_2631);
and UO_544 (O_544,N_3179,N_4408);
nor UO_545 (O_545,N_4295,N_3825);
or UO_546 (O_546,N_4877,N_4659);
nand UO_547 (O_547,N_4194,N_3338);
and UO_548 (O_548,N_4109,N_3481);
or UO_549 (O_549,N_3376,N_3740);
nand UO_550 (O_550,N_3427,N_4497);
nand UO_551 (O_551,N_4581,N_4699);
or UO_552 (O_552,N_4358,N_2566);
and UO_553 (O_553,N_2894,N_4451);
nand UO_554 (O_554,N_3537,N_3768);
nand UO_555 (O_555,N_3630,N_3880);
or UO_556 (O_556,N_4576,N_2823);
nand UO_557 (O_557,N_4675,N_3393);
and UO_558 (O_558,N_2575,N_4154);
nand UO_559 (O_559,N_3862,N_4134);
nand UO_560 (O_560,N_4516,N_2501);
nor UO_561 (O_561,N_2760,N_3255);
or UO_562 (O_562,N_4333,N_3158);
nand UO_563 (O_563,N_4110,N_4780);
and UO_564 (O_564,N_2759,N_4566);
nand UO_565 (O_565,N_4701,N_3332);
and UO_566 (O_566,N_4370,N_3029);
nor UO_567 (O_567,N_2705,N_4705);
nand UO_568 (O_568,N_2788,N_3814);
nand UO_569 (O_569,N_3186,N_3700);
nor UO_570 (O_570,N_4529,N_4012);
nand UO_571 (O_571,N_4405,N_4536);
nor UO_572 (O_572,N_3303,N_2538);
xor UO_573 (O_573,N_4690,N_3106);
nor UO_574 (O_574,N_4991,N_3339);
or UO_575 (O_575,N_4837,N_3681);
nand UO_576 (O_576,N_4202,N_2999);
and UO_577 (O_577,N_4674,N_4669);
nor UO_578 (O_578,N_3992,N_3723);
or UO_579 (O_579,N_3569,N_4524);
nor UO_580 (O_580,N_3165,N_2561);
nand UO_581 (O_581,N_4089,N_3878);
nor UO_582 (O_582,N_3504,N_2903);
nand UO_583 (O_583,N_4759,N_4458);
nand UO_584 (O_584,N_2583,N_3065);
or UO_585 (O_585,N_4504,N_4518);
nor UO_586 (O_586,N_4947,N_4361);
and UO_587 (O_587,N_2867,N_2532);
or UO_588 (O_588,N_3361,N_3320);
and UO_589 (O_589,N_4346,N_3619);
nand UO_590 (O_590,N_3583,N_4635);
nor UO_591 (O_591,N_3649,N_2978);
nor UO_592 (O_592,N_3404,N_4117);
nand UO_593 (O_593,N_3713,N_4622);
and UO_594 (O_594,N_3984,N_2923);
nor UO_595 (O_595,N_3542,N_3503);
nor UO_596 (O_596,N_4097,N_2679);
nor UO_597 (O_597,N_3841,N_4693);
nand UO_598 (O_598,N_2550,N_4148);
and UO_599 (O_599,N_2623,N_3296);
xnor UO_600 (O_600,N_2650,N_4303);
nand UO_601 (O_601,N_4315,N_2733);
or UO_602 (O_602,N_3585,N_3023);
nand UO_603 (O_603,N_3290,N_4942);
nor UO_604 (O_604,N_2941,N_3856);
or UO_605 (O_605,N_3782,N_3714);
and UO_606 (O_606,N_4380,N_3875);
or UO_607 (O_607,N_2673,N_2841);
nand UO_608 (O_608,N_3797,N_3991);
nand UO_609 (O_609,N_2663,N_3801);
and UO_610 (O_610,N_4416,N_4394);
and UO_611 (O_611,N_3128,N_4601);
nand UO_612 (O_612,N_2787,N_3843);
nand UO_613 (O_613,N_3140,N_2969);
nand UO_614 (O_614,N_2526,N_2698);
nand UO_615 (O_615,N_2512,N_2595);
nor UO_616 (O_616,N_4756,N_3746);
nand UO_617 (O_617,N_3802,N_2696);
nand UO_618 (O_618,N_3677,N_3218);
and UO_619 (O_619,N_4999,N_3741);
nor UO_620 (O_620,N_3107,N_2539);
or UO_621 (O_621,N_4873,N_2795);
nand UO_622 (O_622,N_2789,N_3351);
nand UO_623 (O_623,N_3458,N_3637);
nand UO_624 (O_624,N_4988,N_4354);
or UO_625 (O_625,N_4158,N_3090);
and UO_626 (O_626,N_4007,N_4941);
nand UO_627 (O_627,N_4004,N_3410);
and UO_628 (O_628,N_3854,N_4168);
nor UO_629 (O_629,N_2618,N_4243);
nand UO_630 (O_630,N_4159,N_3293);
or UO_631 (O_631,N_2802,N_2900);
nand UO_632 (O_632,N_3011,N_3095);
and UO_633 (O_633,N_3452,N_4449);
nand UO_634 (O_634,N_4343,N_3079);
and UO_635 (O_635,N_2732,N_4395);
or UO_636 (O_636,N_4652,N_4508);
nor UO_637 (O_637,N_4075,N_3076);
nor UO_638 (O_638,N_4956,N_3105);
or UO_639 (O_639,N_3398,N_3547);
nor UO_640 (O_640,N_3005,N_4510);
or UO_641 (O_641,N_4495,N_4409);
or UO_642 (O_642,N_4264,N_3200);
nand UO_643 (O_643,N_4501,N_4647);
or UO_644 (O_644,N_4685,N_3431);
and UO_645 (O_645,N_2677,N_4244);
and UO_646 (O_646,N_3870,N_2930);
or UO_647 (O_647,N_3166,N_4643);
and UO_648 (O_648,N_4191,N_2884);
and UO_649 (O_649,N_4921,N_4454);
and UO_650 (O_650,N_3982,N_4262);
and UO_651 (O_651,N_4978,N_4263);
and UO_652 (O_652,N_4677,N_3350);
nor UO_653 (O_653,N_2834,N_4745);
or UO_654 (O_654,N_4009,N_2509);
nor UO_655 (O_655,N_4627,N_3587);
nand UO_656 (O_656,N_2738,N_4005);
nand UO_657 (O_657,N_3115,N_4369);
nor UO_658 (O_658,N_3187,N_3463);
nor UO_659 (O_659,N_2667,N_4902);
nand UO_660 (O_660,N_2555,N_4279);
nor UO_661 (O_661,N_4989,N_3778);
and UO_662 (O_662,N_4527,N_4715);
nor UO_663 (O_663,N_4645,N_3144);
nor UO_664 (O_664,N_3789,N_4849);
or UO_665 (O_665,N_4371,N_3712);
nor UO_666 (O_666,N_3418,N_4943);
or UO_667 (O_667,N_4616,N_3660);
nor UO_668 (O_668,N_3579,N_4895);
or UO_669 (O_669,N_2910,N_3094);
or UO_670 (O_670,N_4625,N_3189);
or UO_671 (O_671,N_3588,N_3653);
and UO_672 (O_672,N_3730,N_4286);
nand UO_673 (O_673,N_3319,N_4288);
nor UO_674 (O_674,N_3312,N_3206);
nor UO_675 (O_675,N_4113,N_4858);
or UO_676 (O_676,N_3558,N_4602);
and UO_677 (O_677,N_3214,N_3265);
nor UO_678 (O_678,N_3566,N_3855);
xnor UO_679 (O_679,N_3266,N_3381);
or UO_680 (O_680,N_4291,N_4448);
or UO_681 (O_681,N_3928,N_2989);
and UO_682 (O_682,N_4267,N_2784);
or UO_683 (O_683,N_4036,N_2926);
nor UO_684 (O_684,N_4001,N_3907);
nand UO_685 (O_685,N_4979,N_2603);
or UO_686 (O_686,N_3530,N_3348);
nand UO_687 (O_687,N_4383,N_3771);
and UO_688 (O_688,N_3483,N_4359);
or UO_689 (O_689,N_3298,N_4462);
nand UO_690 (O_690,N_4755,N_3224);
xnor UO_691 (O_691,N_4207,N_4260);
and UO_692 (O_692,N_4122,N_4177);
or UO_693 (O_693,N_4923,N_4641);
nand UO_694 (O_694,N_4494,N_2585);
nand UO_695 (O_695,N_3815,N_3489);
nor UO_696 (O_696,N_3926,N_3057);
nor UO_697 (O_697,N_3932,N_3860);
nand UO_698 (O_698,N_3707,N_4438);
nand UO_699 (O_699,N_2648,N_4055);
and UO_700 (O_700,N_3013,N_2911);
nand UO_701 (O_701,N_4880,N_3249);
nor UO_702 (O_702,N_4799,N_3341);
nand UO_703 (O_703,N_4126,N_4477);
nor UO_704 (O_704,N_2537,N_4642);
nand UO_705 (O_705,N_2928,N_3570);
nand UO_706 (O_706,N_3294,N_4908);
nor UO_707 (O_707,N_4424,N_3865);
and UO_708 (O_708,N_2922,N_4915);
and UO_709 (O_709,N_3807,N_3682);
nand UO_710 (O_710,N_3271,N_2721);
and UO_711 (O_711,N_3082,N_4332);
and UO_712 (O_712,N_2838,N_3643);
nand UO_713 (O_713,N_4918,N_4502);
nor UO_714 (O_714,N_2878,N_3353);
and UO_715 (O_715,N_4969,N_3238);
nand UO_716 (O_716,N_3088,N_2937);
nor UO_717 (O_717,N_4757,N_4953);
nor UO_718 (O_718,N_3919,N_3557);
xor UO_719 (O_719,N_2515,N_4513);
nor UO_720 (O_720,N_2804,N_3461);
nand UO_721 (O_721,N_2963,N_2739);
xor UO_722 (O_722,N_4974,N_4331);
or UO_723 (O_723,N_4920,N_3773);
nor UO_724 (O_724,N_4092,N_3129);
and UO_725 (O_725,N_4178,N_3163);
nor UO_726 (O_726,N_4344,N_4257);
nand UO_727 (O_727,N_3434,N_2959);
and UO_728 (O_728,N_3313,N_3656);
and UO_729 (O_729,N_3696,N_4901);
or UO_730 (O_730,N_2722,N_4729);
nand UO_731 (O_731,N_2558,N_3161);
nor UO_732 (O_732,N_4314,N_2707);
nor UO_733 (O_733,N_3679,N_4373);
or UO_734 (O_734,N_3623,N_4038);
nand UO_735 (O_735,N_4865,N_3471);
nand UO_736 (O_736,N_3055,N_4742);
nor UO_737 (O_737,N_3336,N_3665);
or UO_738 (O_738,N_4971,N_3641);
nor UO_739 (O_739,N_4672,N_4963);
nor UO_740 (O_740,N_4682,N_3728);
or UO_741 (O_741,N_3766,N_3142);
or UO_742 (O_742,N_2602,N_4676);
or UO_743 (O_743,N_4163,N_2840);
or UO_744 (O_744,N_4139,N_4393);
nor UO_745 (O_745,N_4224,N_3886);
and UO_746 (O_746,N_4356,N_2889);
nand UO_747 (O_747,N_3572,N_2505);
and UO_748 (O_748,N_2917,N_4557);
nand UO_749 (O_749,N_4473,N_2578);
or UO_750 (O_750,N_3394,N_3321);
or UO_751 (O_751,N_4397,N_4027);
and UO_752 (O_752,N_2608,N_3216);
nand UO_753 (O_753,N_3421,N_3617);
and UO_754 (O_754,N_4552,N_4225);
nor UO_755 (O_755,N_2779,N_3733);
and UO_756 (O_756,N_3775,N_2919);
and UO_757 (O_757,N_3127,N_3646);
and UO_758 (O_758,N_3125,N_2934);
or UO_759 (O_759,N_3219,N_3850);
or UO_760 (O_760,N_3388,N_4401);
or UO_761 (O_761,N_2848,N_2805);
and UO_762 (O_762,N_3600,N_3382);
nand UO_763 (O_763,N_4222,N_3026);
nor UO_764 (O_764,N_3735,N_4668);
and UO_765 (O_765,N_3344,N_2579);
nand UO_766 (O_766,N_3146,N_2758);
or UO_767 (O_767,N_4597,N_4976);
or UO_768 (O_768,N_4044,N_2549);
nand UO_769 (O_769,N_2924,N_2559);
and UO_770 (O_770,N_3071,N_4938);
and UO_771 (O_771,N_2547,N_3981);
and UO_772 (O_772,N_3080,N_4875);
and UO_773 (O_773,N_3390,N_4033);
or UO_774 (O_774,N_4861,N_4773);
or UO_775 (O_775,N_4084,N_3902);
and UO_776 (O_776,N_3455,N_3844);
nor UO_777 (O_777,N_4482,N_2755);
nor UO_778 (O_778,N_3130,N_4857);
nor UO_779 (O_779,N_4308,N_2819);
nand UO_780 (O_780,N_4887,N_3642);
or UO_781 (O_781,N_4932,N_4322);
nand UO_782 (O_782,N_4748,N_4740);
nor UO_783 (O_783,N_2741,N_4088);
and UO_784 (O_784,N_3486,N_3761);
xnor UO_785 (O_785,N_4898,N_2655);
and UO_786 (O_786,N_3793,N_3927);
nor UO_787 (O_787,N_2832,N_4137);
or UO_788 (O_788,N_4367,N_3824);
nor UO_789 (O_789,N_4805,N_4127);
or UO_790 (O_790,N_4066,N_3220);
nand UO_791 (O_791,N_2678,N_3908);
nor UO_792 (O_792,N_2674,N_3466);
and UO_793 (O_793,N_4187,N_2507);
or UO_794 (O_794,N_3364,N_4967);
nand UO_795 (O_795,N_4884,N_4692);
or UO_796 (O_796,N_4946,N_3245);
nand UO_797 (O_797,N_4573,N_3153);
and UO_798 (O_798,N_3199,N_3045);
nor UO_799 (O_799,N_3251,N_4167);
nor UO_800 (O_800,N_2776,N_4738);
or UO_801 (O_801,N_2613,N_4211);
nor UO_802 (O_802,N_3895,N_3201);
nand UO_803 (O_803,N_4188,N_4251);
nor UO_804 (O_804,N_3738,N_2637);
nor UO_805 (O_805,N_3536,N_4851);
or UO_806 (O_806,N_2811,N_2548);
and UO_807 (O_807,N_2596,N_3122);
nand UO_808 (O_808,N_4156,N_2859);
nand UO_809 (O_809,N_3012,N_2860);
nand UO_810 (O_810,N_4241,N_2862);
and UO_811 (O_811,N_4794,N_4366);
nor UO_812 (O_812,N_3593,N_2636);
nor UO_813 (O_813,N_2744,N_3956);
nand UO_814 (O_814,N_2902,N_3453);
nor UO_815 (O_815,N_3765,N_4958);
nand UO_816 (O_816,N_4792,N_4266);
nand UO_817 (O_817,N_3950,N_3781);
or UO_818 (O_818,N_3930,N_4522);
nand UO_819 (O_819,N_4328,N_4927);
nand UO_820 (O_820,N_3309,N_3669);
and UO_821 (O_821,N_4420,N_3840);
or UO_822 (O_822,N_3482,N_4129);
nor UO_823 (O_823,N_3356,N_4890);
or UO_824 (O_824,N_4535,N_4928);
nand UO_825 (O_825,N_2649,N_3715);
nor UO_826 (O_826,N_3845,N_3578);
nor UO_827 (O_827,N_3085,N_4541);
nor UO_828 (O_828,N_3384,N_3905);
or UO_829 (O_829,N_4439,N_4275);
nand UO_830 (O_830,N_2866,N_4816);
and UO_831 (O_831,N_4864,N_4788);
nand UO_832 (O_832,N_4155,N_4662);
nand UO_833 (O_833,N_2780,N_2927);
or UO_834 (O_834,N_3692,N_3849);
nor UO_835 (O_835,N_3024,N_4590);
nor UO_836 (O_836,N_3839,N_3990);
nor UO_837 (O_837,N_4791,N_4736);
nor UO_838 (O_838,N_2792,N_3954);
or UO_839 (O_839,N_4813,N_3762);
nand UO_840 (O_840,N_3968,N_3228);
or UO_841 (O_841,N_4862,N_3852);
and UO_842 (O_842,N_2593,N_3180);
or UO_843 (O_843,N_4231,N_2513);
nand UO_844 (O_844,N_2714,N_4297);
nor UO_845 (O_845,N_2952,N_3796);
nand UO_846 (O_846,N_2518,N_4743);
nand UO_847 (O_847,N_3177,N_4061);
nor UO_848 (O_848,N_4649,N_4783);
or UO_849 (O_849,N_3473,N_2915);
nor UO_850 (O_850,N_3598,N_2887);
and UO_851 (O_851,N_3973,N_4081);
xnor UO_852 (O_852,N_4606,N_4863);
and UO_853 (O_853,N_3511,N_4962);
nand UO_854 (O_854,N_4833,N_3359);
or UO_855 (O_855,N_4214,N_3056);
and UO_856 (O_856,N_4789,N_3822);
or UO_857 (O_857,N_4836,N_4054);
nor UO_858 (O_858,N_3726,N_2520);
nand UO_859 (O_859,N_3264,N_2796);
or UO_860 (O_860,N_3508,N_4656);
nor UO_861 (O_861,N_2708,N_2562);
or UO_862 (O_862,N_3528,N_2892);
nand UO_863 (O_863,N_4881,N_3543);
and UO_864 (O_864,N_2628,N_3644);
or UO_865 (O_865,N_4059,N_2664);
nand UO_866 (O_866,N_2983,N_3821);
and UO_867 (O_867,N_4768,N_4215);
nor UO_868 (O_868,N_4216,N_3440);
or UO_869 (O_869,N_2535,N_4104);
nor UO_870 (O_870,N_4468,N_4292);
nand UO_871 (O_871,N_4258,N_4352);
or UO_872 (O_872,N_2861,N_3306);
nor UO_873 (O_873,N_4140,N_4904);
or UO_874 (O_874,N_2610,N_4801);
and UO_875 (O_875,N_3207,N_4247);
nand UO_876 (O_876,N_3551,N_2942);
or UO_877 (O_877,N_4922,N_2918);
and UO_878 (O_878,N_4939,N_4278);
nor UO_879 (O_879,N_2908,N_3253);
or UO_880 (O_880,N_4720,N_3191);
nand UO_881 (O_881,N_4846,N_4100);
nand UO_882 (O_882,N_4142,N_4912);
nor UO_883 (O_883,N_4400,N_3904);
nor UO_884 (O_884,N_3903,N_3604);
or UO_885 (O_885,N_3043,N_2790);
nand UO_886 (O_886,N_4096,N_2873);
or UO_887 (O_887,N_3032,N_4843);
and UO_888 (O_888,N_3996,N_4695);
and UO_889 (O_889,N_3203,N_2600);
nor UO_890 (O_890,N_2980,N_4700);
nand UO_891 (O_891,N_4697,N_4105);
or UO_892 (O_892,N_2913,N_3810);
nor UO_893 (O_893,N_4703,N_4340);
nand UO_894 (O_894,N_3998,N_4002);
nor UO_895 (O_895,N_4753,N_3357);
xnor UO_896 (O_896,N_4290,N_3424);
nor UO_897 (O_897,N_2773,N_4661);
nor UO_898 (O_898,N_3830,N_3058);
or UO_899 (O_899,N_2609,N_4077);
nor UO_900 (O_900,N_3360,N_3943);
and UO_901 (O_901,N_3501,N_4032);
and UO_902 (O_902,N_4878,N_3519);
nor UO_903 (O_903,N_3181,N_4330);
xnor UO_904 (O_904,N_2630,N_2514);
or UO_905 (O_905,N_4764,N_3687);
nor UO_906 (O_906,N_3197,N_4413);
nand UO_907 (O_907,N_4013,N_3084);
nand UO_908 (O_908,N_3039,N_3576);
and UO_909 (O_909,N_2854,N_3722);
and UO_910 (O_910,N_4342,N_3112);
or UO_911 (O_911,N_2851,N_3325);
or UO_912 (O_912,N_3317,N_2516);
or UO_913 (O_913,N_3942,N_3387);
and UO_914 (O_914,N_3882,N_4528);
nor UO_915 (O_915,N_2589,N_4365);
or UO_916 (O_916,N_4106,N_2660);
or UO_917 (O_917,N_4948,N_3834);
nor UO_918 (O_918,N_3302,N_3616);
nand UO_919 (O_919,N_4173,N_3174);
and UO_920 (O_920,N_3484,N_2936);
nand UO_921 (O_921,N_4709,N_4546);
or UO_922 (O_922,N_4834,N_3004);
or UO_923 (O_923,N_3479,N_2818);
nand UO_924 (O_924,N_2984,N_4184);
nor UO_925 (O_925,N_4025,N_3675);
nor UO_926 (O_926,N_4019,N_3777);
nand UO_927 (O_927,N_4523,N_2973);
or UO_928 (O_928,N_4246,N_4248);
or UO_929 (O_929,N_4143,N_4555);
nor UO_930 (O_930,N_3003,N_4083);
nand UO_931 (O_931,N_4854,N_4230);
and UO_932 (O_932,N_3229,N_4268);
nor UO_933 (O_933,N_3126,N_4421);
or UO_934 (O_934,N_3502,N_3062);
nor UO_935 (O_935,N_2704,N_3185);
and UO_936 (O_936,N_3257,N_4407);
or UO_937 (O_937,N_4615,N_3813);
and UO_938 (O_938,N_2852,N_3925);
and UO_939 (O_939,N_4350,N_2837);
nand UO_940 (O_940,N_4490,N_3010);
nor UO_941 (O_941,N_3054,N_3405);
and UO_942 (O_942,N_3873,N_3597);
and UO_943 (O_943,N_2897,N_4934);
nor UO_944 (O_944,N_4391,N_3846);
or UO_945 (O_945,N_3433,N_3553);
nor UO_946 (O_946,N_3456,N_4556);
nor UO_947 (O_947,N_2502,N_4152);
nand UO_948 (O_948,N_4119,N_4786);
nand UO_949 (O_949,N_4355,N_3053);
nand UO_950 (O_950,N_4955,N_4637);
nor UO_951 (O_951,N_3044,N_3883);
or UO_952 (O_952,N_2665,N_3175);
nor UO_953 (O_953,N_4146,N_2500);
or UO_954 (O_954,N_2657,N_2540);
nand UO_955 (O_955,N_4403,N_3871);
nor UO_956 (O_956,N_4712,N_3555);
and UO_957 (O_957,N_3379,N_3036);
nor UO_958 (O_958,N_4486,N_4253);
nor UO_959 (O_959,N_4415,N_4265);
and UO_960 (O_960,N_4165,N_2905);
nand UO_961 (O_961,N_4429,N_3443);
nand UO_962 (O_962,N_3063,N_2689);
and UO_963 (O_963,N_3674,N_3408);
nand UO_964 (O_964,N_3066,N_3832);
and UO_965 (O_965,N_4517,N_4223);
and UO_966 (O_966,N_4157,N_2987);
and UO_967 (O_967,N_3602,N_3449);
or UO_968 (O_968,N_3446,N_3217);
or UO_969 (O_969,N_2961,N_2553);
or UO_970 (O_970,N_3425,N_3561);
or UO_971 (O_971,N_3488,N_4781);
nor UO_972 (O_972,N_3941,N_3820);
nand UO_973 (O_973,N_3432,N_2666);
nor UO_974 (O_974,N_4776,N_2680);
nor UO_975 (O_975,N_4443,N_2546);
or UO_976 (O_976,N_4132,N_4131);
or UO_977 (O_977,N_2808,N_4289);
nand UO_978 (O_978,N_3610,N_3756);
nor UO_979 (O_979,N_3571,N_4235);
and UO_980 (O_980,N_3093,N_4795);
nor UO_981 (O_981,N_3639,N_4824);
nand UO_982 (O_982,N_3890,N_3407);
or UO_983 (O_983,N_2726,N_4480);
nand UO_984 (O_984,N_4667,N_4572);
nor UO_985 (O_985,N_3487,N_4626);
and UO_986 (O_986,N_3764,N_4663);
or UO_987 (O_987,N_4717,N_4534);
nand UO_988 (O_988,N_4145,N_4826);
nand UO_989 (O_989,N_4804,N_4959);
nor UO_990 (O_990,N_3962,N_4530);
nor UO_991 (O_991,N_4238,N_2709);
or UO_992 (O_992,N_4175,N_2977);
and UO_993 (O_993,N_4418,N_3568);
nand UO_994 (O_994,N_3429,N_3263);
or UO_995 (O_995,N_3049,N_4307);
nor UO_996 (O_996,N_3564,N_4392);
and UO_997 (O_997,N_3374,N_3490);
and UO_998 (O_998,N_3300,N_2668);
nand UO_999 (O_999,N_4561,N_2594);
endmodule