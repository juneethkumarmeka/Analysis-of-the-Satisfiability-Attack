module basic_2000_20000_2500_125_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_1680,In_1688);
nand U1 (N_1,In_212,In_1077);
xor U2 (N_2,In_1586,In_136);
and U3 (N_3,In_871,In_1461);
or U4 (N_4,In_859,In_1233);
xor U5 (N_5,In_1321,In_1611);
or U6 (N_6,In_745,In_603);
xnor U7 (N_7,In_1027,In_63);
xnor U8 (N_8,In_467,In_100);
and U9 (N_9,In_1698,In_1516);
nand U10 (N_10,In_1115,In_1080);
or U11 (N_11,In_504,In_303);
xnor U12 (N_12,In_98,In_1898);
nor U13 (N_13,In_450,In_1226);
xnor U14 (N_14,In_1736,In_509);
and U15 (N_15,In_374,In_667);
xnor U16 (N_16,In_644,In_1220);
nor U17 (N_17,In_388,In_329);
nor U18 (N_18,In_1776,In_1687);
xor U19 (N_19,In_1913,In_201);
or U20 (N_20,In_1616,In_80);
and U21 (N_21,In_1967,In_559);
xnor U22 (N_22,In_576,In_1392);
nor U23 (N_23,In_247,In_769);
nor U24 (N_24,In_1256,In_1710);
and U25 (N_25,In_969,In_736);
nand U26 (N_26,In_1525,In_456);
and U27 (N_27,In_1530,In_645);
nor U28 (N_28,In_6,In_739);
nor U29 (N_29,In_1757,In_673);
nor U30 (N_30,In_1519,In_453);
nor U31 (N_31,In_596,In_485);
xnor U32 (N_32,In_1935,In_1492);
xor U33 (N_33,In_213,In_638);
nand U34 (N_34,In_1417,In_491);
or U35 (N_35,In_1914,In_1154);
and U36 (N_36,In_1265,In_1369);
xor U37 (N_37,In_397,In_698);
and U38 (N_38,In_1542,In_454);
and U39 (N_39,In_909,In_686);
and U40 (N_40,In_1416,In_95);
nor U41 (N_41,In_417,In_110);
xor U42 (N_42,In_305,In_1775);
and U43 (N_43,In_1524,In_1310);
or U44 (N_44,In_1756,In_55);
or U45 (N_45,In_330,In_197);
nor U46 (N_46,In_127,In_1635);
xor U47 (N_47,In_1028,In_279);
nand U48 (N_48,In_549,In_1090);
xor U49 (N_49,In_1514,In_1925);
or U50 (N_50,In_1699,In_0);
nor U51 (N_51,In_1856,In_782);
nor U52 (N_52,In_1789,In_662);
and U53 (N_53,In_1062,In_1668);
or U54 (N_54,In_1407,In_135);
or U55 (N_55,In_1634,In_17);
and U56 (N_56,In_1061,In_1085);
nor U57 (N_57,In_1239,In_1665);
or U58 (N_58,In_10,In_394);
or U59 (N_59,In_1401,In_1866);
xor U60 (N_60,In_142,In_1653);
and U61 (N_61,In_412,In_799);
and U62 (N_62,In_1372,In_392);
xor U63 (N_63,In_1550,In_524);
xnor U64 (N_64,In_1351,In_1997);
nand U65 (N_65,In_477,In_66);
and U66 (N_66,In_1165,In_1870);
and U67 (N_67,In_1670,In_1303);
nor U68 (N_68,In_1112,In_1485);
xor U69 (N_69,In_500,In_1628);
nor U70 (N_70,In_1824,In_387);
xor U71 (N_71,In_1273,In_992);
xor U72 (N_72,In_1329,In_1672);
nor U73 (N_73,In_1383,In_921);
or U74 (N_74,In_1053,In_101);
and U75 (N_75,In_1119,In_368);
nor U76 (N_76,In_78,In_1049);
or U77 (N_77,In_836,In_902);
nand U78 (N_78,In_382,In_125);
xor U79 (N_79,In_1228,In_344);
or U80 (N_80,In_821,In_1174);
nor U81 (N_81,In_1229,In_233);
and U82 (N_82,In_128,In_109);
xor U83 (N_83,In_1686,In_946);
and U84 (N_84,In_705,In_660);
xor U85 (N_85,In_1703,In_1422);
nand U86 (N_86,In_1939,In_1252);
and U87 (N_87,In_187,In_123);
nor U88 (N_88,In_1325,In_883);
xnor U89 (N_89,In_196,In_1350);
and U90 (N_90,In_1095,In_360);
nor U91 (N_91,In_1158,In_238);
or U92 (N_92,In_1359,In_484);
nor U93 (N_93,In_1716,In_929);
nor U94 (N_94,In_376,In_200);
or U95 (N_95,In_270,In_1783);
or U96 (N_96,In_928,In_246);
nor U97 (N_97,In_428,In_255);
nand U98 (N_98,In_832,In_1786);
nor U99 (N_99,In_361,In_1352);
or U100 (N_100,In_1784,In_297);
nor U101 (N_101,In_138,In_882);
xor U102 (N_102,In_1551,In_399);
nand U103 (N_103,In_1780,In_1408);
nand U104 (N_104,In_1510,In_1613);
nor U105 (N_105,In_906,In_1587);
and U106 (N_106,In_1732,In_1627);
and U107 (N_107,In_35,In_1978);
or U108 (N_108,In_1526,In_1943);
or U109 (N_109,In_966,In_150);
nor U110 (N_110,In_1884,In_824);
nand U111 (N_111,In_370,In_106);
nor U112 (N_112,In_391,In_621);
nor U113 (N_113,In_770,In_7);
nand U114 (N_114,In_1639,In_301);
xnor U115 (N_115,In_1176,In_577);
xnor U116 (N_116,In_521,In_758);
and U117 (N_117,In_1,In_1218);
nand U118 (N_118,In_1646,In_1840);
nand U119 (N_119,In_1110,In_157);
nor U120 (N_120,In_126,In_1597);
nand U121 (N_121,In_444,In_111);
or U122 (N_122,In_77,In_272);
and U123 (N_123,In_515,In_99);
nand U124 (N_124,In_1098,In_221);
or U125 (N_125,In_403,In_217);
nor U126 (N_126,In_476,In_1696);
or U127 (N_127,In_846,In_520);
nand U128 (N_128,In_1952,In_1950);
and U129 (N_129,In_597,In_557);
nor U130 (N_130,In_1755,In_1508);
or U131 (N_131,In_265,In_292);
or U132 (N_132,In_1173,In_240);
or U133 (N_133,In_1035,In_1196);
nor U134 (N_134,In_1205,In_1560);
and U135 (N_135,In_845,In_658);
xnor U136 (N_136,In_993,In_566);
nor U137 (N_137,In_203,In_1466);
and U138 (N_138,In_1652,In_923);
xnor U139 (N_139,In_593,In_937);
or U140 (N_140,In_1713,In_1367);
nor U141 (N_141,In_1896,In_812);
nor U142 (N_142,In_314,In_919);
nor U143 (N_143,In_85,In_271);
and U144 (N_144,In_877,In_1827);
nand U145 (N_145,In_1153,In_766);
nand U146 (N_146,In_1195,In_1497);
and U147 (N_147,In_525,In_588);
xnor U148 (N_148,In_1963,In_1293);
nor U149 (N_149,In_1382,In_1880);
or U150 (N_150,In_345,In_1754);
nand U151 (N_151,In_1415,In_1473);
nor U152 (N_152,In_974,In_897);
nor U153 (N_153,In_1948,In_1442);
or U154 (N_154,In_1395,In_1370);
xor U155 (N_155,In_62,In_88);
nor U156 (N_156,In_1503,In_1316);
or U157 (N_157,In_1488,In_180);
or U158 (N_158,In_1044,In_1905);
or U159 (N_159,In_340,In_1720);
xor U160 (N_160,In_1447,In_129);
or U161 (N_161,In_619,In_818);
nand U162 (N_162,In_1179,In_552);
xnor U163 (N_163,In_837,In_1828);
and U164 (N_164,In_1439,In_1254);
and U165 (N_165,In_1332,In_730);
nand U166 (N_166,In_1163,In_390);
nand U167 (N_167,In_1093,In_1983);
or U168 (N_168,In_1452,In_231);
or U169 (N_169,In_1976,In_1043);
xor U170 (N_170,In_1770,In_1830);
and U171 (N_171,In_1617,In_19);
xor U172 (N_172,In_1929,In_1225);
nor U173 (N_173,In_888,In_398);
or U174 (N_174,In_1462,In_961);
and U175 (N_175,In_1106,In_1603);
nor U176 (N_176,In_1150,In_1326);
or U177 (N_177,In_634,In_37);
and U178 (N_178,In_317,In_1025);
and U179 (N_179,In_190,In_594);
and U180 (N_180,In_267,In_995);
nor U181 (N_181,In_1660,N_125);
nor U182 (N_182,In_924,In_1607);
or U183 (N_183,In_1164,In_1638);
xnor U184 (N_184,In_1109,In_1796);
nand U185 (N_185,In_1299,In_636);
and U186 (N_186,In_1219,N_70);
nand U187 (N_187,In_1702,N_123);
nor U188 (N_188,In_1450,In_179);
or U189 (N_189,In_115,In_1663);
nand U190 (N_190,In_1190,In_965);
nand U191 (N_191,In_1869,In_696);
xnor U192 (N_192,In_1889,In_1169);
or U193 (N_193,In_9,In_1216);
xnor U194 (N_194,In_1436,In_1868);
xor U195 (N_195,In_304,In_1835);
nor U196 (N_196,In_1811,In_905);
nor U197 (N_197,In_1182,In_1527);
and U198 (N_198,In_872,In_733);
nor U199 (N_199,In_1575,In_373);
nand U200 (N_200,In_280,In_1867);
or U201 (N_201,In_1120,N_20);
or U202 (N_202,In_1599,N_146);
xor U203 (N_203,In_1002,N_94);
and U204 (N_204,In_1026,In_1353);
nor U205 (N_205,In_1418,In_1319);
and U206 (N_206,In_1297,N_72);
nor U207 (N_207,In_1821,In_413);
and U208 (N_208,In_12,In_1556);
xnor U209 (N_209,In_1727,In_439);
xnor U210 (N_210,In_16,In_1381);
xor U211 (N_211,In_797,In_1760);
nand U212 (N_212,In_589,In_1344);
nor U213 (N_213,In_1269,In_757);
nor U214 (N_214,In_1096,In_1537);
or U215 (N_215,In_659,In_1358);
nand U216 (N_216,In_1052,In_1191);
and U217 (N_217,In_1576,In_257);
nand U218 (N_218,In_162,In_1301);
or U219 (N_219,In_438,In_618);
or U220 (N_220,In_606,In_1640);
xnor U221 (N_221,In_1136,In_1454);
and U222 (N_222,In_1743,In_516);
nor U223 (N_223,In_1393,In_1151);
nand U224 (N_224,In_754,In_1340);
xor U225 (N_225,In_73,In_1006);
nand U226 (N_226,In_1388,In_1572);
xnor U227 (N_227,In_79,In_1773);
nand U228 (N_228,In_496,N_140);
or U229 (N_229,In_748,In_497);
xnor U230 (N_230,In_1435,In_418);
nand U231 (N_231,In_1232,In_436);
nand U232 (N_232,In_389,In_1331);
nor U233 (N_233,In_1570,In_1446);
nor U234 (N_234,In_868,In_568);
nor U235 (N_235,In_273,In_1504);
or U236 (N_236,In_911,In_982);
and U237 (N_237,In_176,In_1464);
or U238 (N_238,In_224,In_1569);
nor U239 (N_239,In_1557,In_1936);
and U240 (N_240,In_1546,In_774);
xnor U241 (N_241,In_781,In_464);
nand U242 (N_242,In_721,In_259);
xnor U243 (N_243,N_122,In_651);
nand U244 (N_244,In_457,In_1031);
nand U245 (N_245,In_184,In_410);
nand U246 (N_246,In_564,In_1612);
and U247 (N_247,In_1582,In_1295);
xor U248 (N_248,In_808,In_790);
xor U249 (N_249,In_1246,In_86);
and U250 (N_250,In_1449,N_131);
and U251 (N_251,In_994,In_321);
or U252 (N_252,In_141,In_1354);
and U253 (N_253,In_1521,In_599);
xnor U254 (N_254,In_1791,N_99);
nor U255 (N_255,In_1045,In_396);
and U256 (N_256,In_843,In_964);
nor U257 (N_257,In_433,In_121);
nor U258 (N_258,In_1724,In_1723);
nand U259 (N_259,In_1910,In_296);
xnor U260 (N_260,In_627,In_1932);
or U261 (N_261,N_156,In_1363);
or U262 (N_262,In_1604,In_1021);
nand U263 (N_263,In_237,In_1260);
nor U264 (N_264,In_1583,In_546);
nor U265 (N_265,In_1101,In_737);
xor U266 (N_266,In_1865,In_1956);
or U267 (N_267,In_849,In_1066);
nor U268 (N_268,In_1955,In_980);
nand U269 (N_269,In_1281,In_498);
xor U270 (N_270,In_1306,In_1036);
nor U271 (N_271,In_1730,In_1498);
or U272 (N_272,In_186,In_230);
nor U273 (N_273,In_1313,In_1270);
or U274 (N_274,In_199,In_865);
nand U275 (N_275,In_744,In_1651);
or U276 (N_276,In_1209,In_989);
and U277 (N_277,In_894,In_510);
xor U278 (N_278,In_851,In_567);
nor U279 (N_279,In_407,In_1506);
nor U280 (N_280,In_1289,N_27);
nand U281 (N_281,In_117,In_1079);
nand U282 (N_282,In_1368,In_1779);
and U283 (N_283,In_1901,N_67);
nor U284 (N_284,In_1788,N_109);
nor U285 (N_285,In_1142,In_1704);
nand U286 (N_286,In_1494,In_74);
nand U287 (N_287,In_879,In_786);
nor U288 (N_288,In_1923,In_1500);
and U289 (N_289,N_63,In_487);
nor U290 (N_290,In_1130,In_1425);
nor U291 (N_291,In_1945,In_421);
and U292 (N_292,In_94,In_1734);
nand U293 (N_293,In_1211,In_1648);
nor U294 (N_294,In_343,In_538);
or U295 (N_295,N_6,In_572);
or U296 (N_296,In_14,In_302);
xnor U297 (N_297,In_278,In_963);
xnor U298 (N_298,In_558,In_772);
nand U299 (N_299,In_1701,In_1960);
nor U300 (N_300,In_1481,In_1197);
and U301 (N_301,In_540,In_967);
and U302 (N_302,N_16,In_1596);
or U303 (N_303,In_656,In_1903);
nor U304 (N_304,In_1738,N_136);
xnor U305 (N_305,In_1404,N_141);
or U306 (N_306,N_103,In_1991);
and U307 (N_307,In_1808,In_1157);
nor U308 (N_308,In_380,In_1421);
and U309 (N_309,In_424,In_1831);
nor U310 (N_310,In_641,N_119);
nand U311 (N_311,In_1041,In_161);
nand U312 (N_312,In_1857,In_530);
and U313 (N_313,In_1394,In_1279);
nand U314 (N_314,In_352,In_1694);
nand U315 (N_315,In_1377,In_1102);
xor U316 (N_316,N_2,In_420);
and U317 (N_317,In_1201,In_910);
nor U318 (N_318,In_218,In_1739);
or U319 (N_319,In_1785,N_148);
or U320 (N_320,In_1592,In_1558);
nand U321 (N_321,In_550,In_976);
xnor U322 (N_322,In_1700,In_695);
and U323 (N_323,In_935,In_1740);
nor U324 (N_324,In_1222,In_72);
or U325 (N_325,In_1735,In_326);
nand U326 (N_326,In_1308,In_1148);
or U327 (N_327,In_828,N_158);
and U328 (N_328,In_1000,In_778);
nand U329 (N_329,N_126,In_985);
xor U330 (N_330,N_7,In_622);
and U331 (N_331,In_1916,In_1056);
and U332 (N_332,In_1766,In_36);
nand U333 (N_333,In_5,In_1479);
or U334 (N_334,In_1207,In_60);
nor U335 (N_335,In_1986,In_1682);
xor U336 (N_336,In_1237,In_152);
nand U337 (N_337,In_1515,In_1975);
nor U338 (N_338,In_1145,In_1656);
or U339 (N_339,N_160,In_1227);
xnor U340 (N_340,In_1387,In_1649);
nand U341 (N_341,N_279,N_280);
nor U342 (N_342,In_105,In_473);
or U343 (N_343,In_999,N_101);
or U344 (N_344,In_853,N_261);
nand U345 (N_345,In_245,In_1873);
or U346 (N_346,In_277,In_291);
nand U347 (N_347,In_283,In_1834);
or U348 (N_348,In_1444,In_1501);
nor U349 (N_349,In_1584,N_310);
nand U350 (N_350,N_175,In_248);
or U351 (N_351,N_128,N_57);
xor U352 (N_352,In_1888,N_32);
nor U353 (N_353,In_1750,In_1841);
xnor U354 (N_354,In_2,In_50);
nand U355 (N_355,In_1618,N_78);
nand U356 (N_356,In_1549,In_1328);
and U357 (N_357,In_258,N_145);
and U358 (N_358,In_971,N_264);
xnor U359 (N_359,In_1919,In_53);
nor U360 (N_360,In_1589,N_177);
and U361 (N_361,In_1793,In_518);
xor U362 (N_362,In_263,N_69);
nor U363 (N_363,In_648,In_735);
or U364 (N_364,In_167,In_1129);
or U365 (N_365,In_83,In_235);
nor U366 (N_366,In_81,In_1075);
nor U367 (N_367,In_850,In_652);
xnor U368 (N_368,In_502,In_1305);
and U369 (N_369,In_1374,N_306);
or U370 (N_370,In_1330,In_182);
or U371 (N_371,In_563,N_164);
xor U372 (N_372,In_1259,In_1250);
and U373 (N_373,N_55,In_598);
or U374 (N_374,In_674,In_1941);
nor U375 (N_375,In_132,In_427);
and U376 (N_376,In_202,In_1470);
nor U377 (N_377,In_383,In_541);
nor U378 (N_378,In_1568,In_810);
or U379 (N_379,In_873,In_1008);
and U380 (N_380,In_466,N_237);
nand U381 (N_381,In_249,In_1807);
nor U382 (N_382,In_372,In_1661);
or U383 (N_383,In_188,In_1317);
or U384 (N_384,In_844,In_1143);
nand U385 (N_385,N_302,In_1046);
and U386 (N_386,In_350,N_24);
or U387 (N_387,In_1161,In_1091);
or U388 (N_388,In_1675,In_404);
and U389 (N_389,In_90,In_814);
or U390 (N_390,In_1768,In_1994);
nand U391 (N_391,In_975,In_813);
nand U392 (N_392,In_1794,In_896);
nand U393 (N_393,In_932,In_801);
nor U394 (N_394,In_1141,In_346);
nand U395 (N_395,In_171,In_997);
xnor U396 (N_396,In_1223,In_458);
or U397 (N_397,In_1862,In_1647);
nor U398 (N_398,In_691,In_1455);
and U399 (N_399,In_118,In_998);
nor U400 (N_400,In_144,In_722);
nand U401 (N_401,In_571,In_710);
nand U402 (N_402,In_779,In_1839);
or U403 (N_403,In_855,In_59);
or U404 (N_404,In_1541,In_762);
nor U405 (N_405,N_77,In_1972);
nand U406 (N_406,N_170,In_44);
or U407 (N_407,In_1030,In_205);
nand U408 (N_408,In_983,In_825);
nor U409 (N_409,N_19,In_1619);
nand U410 (N_410,In_131,In_941);
xor U411 (N_411,In_1745,In_944);
and U412 (N_412,In_1581,In_1263);
or U413 (N_413,In_889,N_165);
xnor U414 (N_414,In_1988,N_193);
xor U415 (N_415,In_429,In_1765);
xor U416 (N_416,In_1610,In_988);
or U417 (N_417,In_1078,In_1114);
and U418 (N_418,In_285,In_834);
xnor U419 (N_419,In_1457,N_102);
nand U420 (N_420,In_1721,N_257);
or U421 (N_421,In_1128,In_465);
xor U422 (N_422,N_41,In_1626);
nand U423 (N_423,In_1005,In_338);
and U424 (N_424,In_1014,In_1189);
nand U425 (N_425,In_945,In_827);
nand U426 (N_426,In_806,In_1790);
and U427 (N_427,In_917,N_272);
nand U428 (N_428,In_1763,In_1480);
nor U429 (N_429,In_1375,In_1762);
nor U430 (N_430,In_1210,N_120);
nor U431 (N_431,In_1645,In_1904);
xor U432 (N_432,N_179,N_86);
nor U433 (N_433,In_140,In_22);
and U434 (N_434,N_89,In_445);
or U435 (N_435,In_1644,In_907);
or U436 (N_436,In_1906,N_311);
or U437 (N_437,In_1202,In_1341);
and U438 (N_438,In_82,In_1468);
or U439 (N_439,N_112,N_276);
and U440 (N_440,N_144,In_1371);
or U441 (N_441,In_69,In_1257);
or U442 (N_442,In_1314,In_1453);
or U443 (N_443,In_887,In_539);
nand U444 (N_444,In_401,In_1007);
or U445 (N_445,In_1787,N_45);
nor U446 (N_446,N_196,In_1116);
nor U447 (N_447,In_954,In_359);
or U448 (N_448,In_435,In_462);
or U449 (N_449,In_1463,In_1437);
or U450 (N_450,In_743,In_1380);
nor U451 (N_451,In_616,In_193);
nand U452 (N_452,In_1117,In_300);
or U453 (N_453,N_107,In_318);
nand U454 (N_454,In_1961,In_1926);
nor U455 (N_455,In_590,In_613);
or U456 (N_456,In_363,N_298);
xnor U457 (N_457,In_1726,In_1336);
nand U458 (N_458,In_1288,In_1029);
and U459 (N_459,In_1100,N_251);
and U460 (N_460,In_1574,In_1047);
nand U461 (N_461,In_1822,In_1188);
xor U462 (N_462,N_299,In_1826);
nand U463 (N_463,N_252,In_717);
or U464 (N_464,In_908,In_522);
xor U465 (N_465,In_1039,In_565);
or U466 (N_466,In_712,In_791);
or U467 (N_467,N_8,In_1915);
nand U468 (N_468,In_324,N_73);
nor U469 (N_469,In_319,In_1864);
nand U470 (N_470,N_300,N_296);
and U471 (N_471,In_513,In_1034);
nor U472 (N_472,In_1854,In_1108);
and U473 (N_473,N_43,In_1302);
xnor U474 (N_474,In_1015,N_15);
and U475 (N_475,In_24,In_92);
or U476 (N_476,In_1771,In_31);
nor U477 (N_477,In_649,In_96);
xnor U478 (N_478,In_1609,In_1271);
or U479 (N_479,In_901,In_1709);
nor U480 (N_480,In_1654,N_233);
and U481 (N_481,In_684,N_475);
nand U482 (N_482,In_1140,In_312);
and U483 (N_483,In_1998,In_933);
or U484 (N_484,In_1063,In_1089);
xnor U485 (N_485,In_269,In_847);
nand U486 (N_486,In_1683,In_411);
nand U487 (N_487,In_243,In_236);
nand U488 (N_488,In_1725,N_361);
xnor U489 (N_489,In_1817,N_267);
nand U490 (N_490,N_387,In_752);
nand U491 (N_491,In_451,N_12);
nand U492 (N_492,In_728,N_21);
xnor U493 (N_493,N_396,In_1477);
nand U494 (N_494,In_867,In_671);
xnor U495 (N_495,In_723,N_418);
or U496 (N_496,N_203,In_569);
nand U497 (N_497,In_449,In_1206);
and U498 (N_498,In_1171,N_368);
and U499 (N_499,N_462,In_1718);
nor U500 (N_500,N_275,In_173);
nand U501 (N_501,In_1083,In_543);
xnor U502 (N_502,N_255,In_145);
nand U503 (N_503,N_304,In_1722);
nand U504 (N_504,In_1249,N_98);
nor U505 (N_505,In_289,N_402);
or U506 (N_506,In_339,In_1010);
nor U507 (N_507,In_1475,N_96);
xor U508 (N_508,In_226,N_256);
xnor U509 (N_509,In_623,In_893);
and U510 (N_510,N_408,In_629);
nand U511 (N_511,In_1139,N_208);
and U512 (N_512,N_357,In_1474);
nand U513 (N_513,In_750,In_996);
nand U514 (N_514,N_465,N_87);
or U515 (N_515,N_364,In_430);
xnor U516 (N_516,N_31,In_393);
or U517 (N_517,N_392,In_523);
nand U518 (N_518,In_137,N_91);
and U519 (N_519,In_32,In_195);
or U520 (N_520,In_783,In_1097);
xor U521 (N_521,N_312,In_1928);
nand U522 (N_522,In_211,N_190);
or U523 (N_523,In_679,In_1386);
and U524 (N_524,In_1087,In_1378);
nor U525 (N_525,N_22,In_1594);
nor U526 (N_526,In_1184,In_1567);
and U527 (N_527,In_1962,In_809);
nand U528 (N_528,N_149,In_1215);
nor U529 (N_529,N_371,In_642);
nand U530 (N_530,In_841,In_1887);
and U531 (N_531,In_1847,In_1520);
nand U532 (N_532,In_1135,In_1275);
or U533 (N_533,In_1517,In_731);
and U534 (N_534,In_1992,In_562);
nand U535 (N_535,In_1606,In_1471);
nand U536 (N_536,In_716,In_1547);
nor U537 (N_537,N_84,In_489);
or U538 (N_538,In_1798,In_1534);
or U539 (N_539,N_200,N_192);
xor U540 (N_540,In_777,N_297);
nand U541 (N_541,In_46,N_260);
and U542 (N_542,In_507,N_48);
xnor U543 (N_543,In_612,In_1213);
or U544 (N_544,In_536,N_332);
or U545 (N_545,In_337,N_295);
xnor U546 (N_546,N_211,In_688);
nand U547 (N_547,N_79,In_1655);
xnor U548 (N_548,In_64,N_29);
nor U549 (N_549,In_286,In_1057);
xor U550 (N_550,N_404,In_103);
nand U551 (N_551,In_1071,In_1253);
nand U552 (N_552,In_1650,N_314);
xnor U553 (N_553,In_1286,In_817);
and U554 (N_554,N_258,In_1861);
xnor U555 (N_555,In_1819,In_517);
xor U556 (N_556,In_1614,In_288);
and U557 (N_557,In_1199,In_624);
or U558 (N_558,In_253,N_181);
nand U559 (N_559,In_335,In_1658);
or U560 (N_560,N_452,In_1020);
nor U561 (N_561,In_657,In_1883);
and U562 (N_562,N_245,N_25);
nor U563 (N_563,In_470,N_320);
xnor U564 (N_564,In_1748,In_1484);
xor U565 (N_565,In_811,In_1620);
or U566 (N_566,In_1185,In_463);
nand U567 (N_567,In_1685,N_61);
or U568 (N_568,N_301,N_82);
and U569 (N_569,In_1054,In_1989);
or U570 (N_570,N_75,In_1280);
or U571 (N_571,In_1348,In_1958);
and U572 (N_572,In_1432,In_708);
nand U573 (N_573,In_1879,In_1664);
nor U574 (N_574,N_472,N_307);
xnor U575 (N_575,N_97,In_362);
or U576 (N_576,In_268,In_108);
nand U577 (N_577,In_198,In_842);
xnor U578 (N_578,N_278,In_93);
xor U579 (N_579,In_1907,In_1893);
nor U580 (N_580,In_1832,In_900);
or U581 (N_581,In_1347,In_574);
and U582 (N_582,In_665,In_1287);
nor U583 (N_583,In_431,N_173);
or U584 (N_584,In_1337,N_425);
nand U585 (N_585,In_1881,In_1290);
or U586 (N_586,In_669,N_342);
nor U587 (N_587,In_1908,N_132);
nand U588 (N_588,In_1152,In_165);
xor U589 (N_589,In_1897,In_931);
or U590 (N_590,In_802,N_228);
and U591 (N_591,In_1621,In_1134);
and U592 (N_592,In_1282,N_340);
or U593 (N_593,N_427,In_1133);
xnor U594 (N_594,In_794,N_157);
and U595 (N_595,In_1070,In_1759);
and U596 (N_596,In_687,In_863);
xor U597 (N_597,N_176,In_890);
and U598 (N_598,In_91,In_38);
or U599 (N_599,In_1706,In_461);
nor U600 (N_600,N_326,N_391);
and U601 (N_601,In_189,In_1899);
or U602 (N_602,In_1406,In_1274);
xnor U603 (N_603,In_1084,N_263);
or U604 (N_604,In_1565,N_60);
or U605 (N_605,In_322,In_903);
xor U606 (N_606,In_1334,In_1637);
nor U607 (N_607,N_108,In_369);
nor U608 (N_608,In_753,In_1985);
or U609 (N_609,In_1984,In_1930);
or U610 (N_610,In_789,In_1578);
and U611 (N_611,In_578,In_122);
nand U612 (N_612,In_1086,N_247);
and U613 (N_613,In_426,In_639);
nor U614 (N_614,In_987,In_1162);
nand U615 (N_615,In_1409,In_1823);
nor U616 (N_616,In_1124,N_174);
and U617 (N_617,N_414,N_370);
xor U618 (N_618,In_765,N_167);
xnor U619 (N_619,N_5,In_18);
xor U620 (N_620,In_215,In_1859);
and U621 (N_621,In_1561,In_720);
or U622 (N_622,In_1376,N_186);
nor U623 (N_623,In_628,In_1818);
nor U624 (N_624,In_1598,In_351);
or U625 (N_625,In_544,In_979);
nand U626 (N_626,In_1953,In_692);
or U627 (N_627,In_1693,In_1630);
and U628 (N_628,In_1060,N_283);
and U629 (N_629,In_114,N_321);
xnor U630 (N_630,In_1333,In_816);
nor U631 (N_631,In_42,In_822);
nor U632 (N_632,In_1632,In_1458);
xnor U633 (N_633,N_453,In_1366);
or U634 (N_634,In_796,In_1441);
xor U635 (N_635,In_776,In_156);
nand U636 (N_636,In_170,In_1933);
nand U637 (N_637,In_220,In_819);
and U638 (N_638,N_430,N_351);
or U639 (N_639,In_1924,In_1361);
or U640 (N_640,In_990,In_1615);
nor U641 (N_641,In_1429,In_1518);
xor U642 (N_642,N_106,N_480);
xnor U643 (N_643,N_474,In_742);
nor U644 (N_644,In_1591,In_1127);
and U645 (N_645,N_540,In_755);
or U646 (N_646,In_97,In_1251);
nand U647 (N_647,N_531,N_512);
nand U648 (N_648,In_342,N_339);
xor U649 (N_649,In_210,In_1741);
and U650 (N_650,In_1678,N_234);
xnor U651 (N_651,N_441,In_437);
nand U652 (N_652,In_27,N_23);
nor U653 (N_653,In_1815,In_1657);
and U654 (N_654,In_1631,In_481);
nor U655 (N_655,N_573,In_1126);
and U656 (N_656,N_603,In_1545);
and U657 (N_657,In_229,In_1585);
nor U658 (N_658,N_596,In_1243);
xnor U659 (N_659,N_529,In_334);
nor U660 (N_660,N_405,In_864);
xnor U661 (N_661,In_21,In_409);
xnor U662 (N_662,In_1911,In_275);
nand U663 (N_663,N_511,In_1717);
or U664 (N_664,N_217,In_354);
nor U665 (N_665,In_501,In_386);
xor U666 (N_666,N_248,In_1799);
or U667 (N_667,In_1430,In_820);
and U668 (N_668,In_925,In_719);
nor U669 (N_669,In_134,In_1731);
nand U670 (N_670,N_64,In_1947);
nand U671 (N_671,In_89,N_526);
xnor U672 (N_672,In_166,N_58);
or U673 (N_673,In_1405,In_299);
and U674 (N_674,N_114,In_1167);
xor U675 (N_675,N_493,N_305);
xor U676 (N_676,In_1338,In_678);
nand U677 (N_677,In_787,In_1431);
nor U678 (N_678,N_13,N_547);
nor U679 (N_679,In_348,N_49);
nor U680 (N_680,N_397,In_927);
or U681 (N_681,In_113,In_711);
nor U682 (N_682,N_551,N_277);
and U683 (N_683,In_1122,In_356);
nor U684 (N_684,In_1900,In_1487);
xor U685 (N_685,In_1999,In_1082);
and U686 (N_686,In_554,In_367);
or U687 (N_687,N_230,In_194);
nor U688 (N_688,N_555,In_1511);
or U689 (N_689,In_1318,In_124);
and U690 (N_690,In_1711,In_174);
nor U691 (N_691,In_654,In_840);
nor U692 (N_692,In_1312,In_130);
or U693 (N_693,In_579,N_409);
nand U694 (N_694,In_1094,In_1708);
nand U695 (N_695,In_1959,In_1820);
or U696 (N_696,In_1949,N_337);
nor U697 (N_697,N_598,In_1954);
or U698 (N_698,N_510,In_1067);
and U699 (N_699,In_29,In_1107);
nor U700 (N_700,In_1414,In_1284);
xor U701 (N_701,N_130,In_274);
and U702 (N_702,N_636,In_1878);
nor U703 (N_703,In_650,N_290);
nand U704 (N_704,N_62,In_1806);
nor U705 (N_705,N_490,In_47);
or U706 (N_706,In_379,N_600);
xnor U707 (N_707,In_1013,In_1742);
and U708 (N_708,In_1965,In_815);
nand U709 (N_709,In_630,In_1402);
nor U710 (N_710,In_1016,In_1848);
xnor U711 (N_711,N_259,In_1810);
or U712 (N_712,N_561,In_1797);
or U713 (N_713,In_1712,In_767);
nor U714 (N_714,In_34,In_1917);
nand U715 (N_715,In_377,In_551);
nor U716 (N_716,In_1037,N_169);
nand U717 (N_717,N_214,N_372);
xor U718 (N_718,In_1103,In_1800);
nor U719 (N_719,In_693,In_1691);
and U720 (N_720,In_492,In_1050);
or U721 (N_721,In_432,In_915);
nor U722 (N_722,In_1974,In_474);
nor U723 (N_723,In_874,In_1894);
xnor U724 (N_724,In_601,In_1902);
xnor U725 (N_725,In_1081,In_1507);
xor U726 (N_726,In_1751,In_1689);
or U727 (N_727,In_1573,In_1977);
or U728 (N_728,In_1968,In_916);
or U729 (N_729,In_155,N_253);
and U730 (N_730,N_243,N_574);
and U731 (N_731,In_1764,N_479);
xnor U732 (N_732,In_1580,In_177);
or U733 (N_733,In_287,N_489);
nand U734 (N_734,In_663,N_579);
nand U735 (N_735,In_1278,In_1781);
xnor U736 (N_736,In_1970,In_1113);
nand U737 (N_737,In_953,N_4);
or U738 (N_738,In_1496,In_561);
nand U739 (N_739,In_1230,N_168);
nand U740 (N_740,N_380,N_550);
nor U741 (N_741,In_697,N_617);
nor U742 (N_742,N_350,In_349);
or U743 (N_743,In_49,In_1844);
and U744 (N_744,In_899,In_582);
nor U745 (N_745,In_440,N_90);
or U746 (N_746,N_115,N_289);
nor U747 (N_747,N_552,In_441);
nand U748 (N_748,N_507,In_959);
xnor U749 (N_749,N_495,N_369);
nor U750 (N_750,N_100,N_587);
or U751 (N_751,In_1895,N_412);
or U752 (N_752,In_614,In_320);
nand U753 (N_753,In_1667,N_184);
or U754 (N_754,In_1579,In_870);
nor U755 (N_755,In_1662,N_590);
nand U756 (N_756,N_580,N_487);
xor U757 (N_757,N_469,N_486);
xnor U758 (N_758,In_1194,N_93);
and U759 (N_759,In_1231,In_308);
and U760 (N_760,In_353,In_1995);
and U761 (N_761,In_1105,In_1440);
nand U762 (N_762,In_1629,N_207);
or U763 (N_763,In_1753,N_0);
or U764 (N_764,N_143,In_570);
or U765 (N_765,N_265,N_390);
and U766 (N_766,In_580,In_1882);
or U767 (N_767,In_610,In_48);
or U768 (N_768,N_9,In_154);
and U769 (N_769,N_218,N_416);
or U770 (N_770,In_75,N_88);
and U771 (N_771,In_1149,In_1168);
nor U772 (N_772,In_447,In_972);
nand U773 (N_773,N_204,In_1069);
and U774 (N_774,N_113,N_627);
nand U775 (N_775,In_1170,In_1132);
or U776 (N_776,In_160,In_605);
or U777 (N_777,In_1390,N_225);
nor U778 (N_778,In_1761,In_207);
nand U779 (N_779,In_1940,N_324);
nor U780 (N_780,N_419,In_40);
or U781 (N_781,In_1004,In_1419);
xnor U782 (N_782,N_42,In_955);
or U783 (N_783,N_609,N_496);
or U784 (N_784,N_542,In_957);
nor U785 (N_785,In_1420,In_1801);
or U786 (N_786,N_595,N_51);
nor U787 (N_787,N_388,In_699);
nand U788 (N_788,N_348,In_1927);
xor U789 (N_789,N_394,N_481);
and U790 (N_790,N_400,N_437);
nand U791 (N_791,In_986,N_594);
nor U792 (N_792,N_544,In_260);
nor U793 (N_793,In_1944,In_228);
xor U794 (N_794,N_343,N_242);
or U795 (N_795,N_426,N_374);
and U796 (N_796,In_316,In_459);
or U797 (N_797,In_1123,N_583);
xor U798 (N_798,In_1495,In_646);
xnor U799 (N_799,In_493,N_520);
nor U800 (N_800,N_616,In_239);
xnor U801 (N_801,N_118,N_421);
nand U802 (N_802,In_1476,In_169);
nand U803 (N_803,In_1964,N_456);
nor U804 (N_804,In_378,N_334);
and U805 (N_805,In_478,In_922);
xnor U806 (N_806,N_375,N_652);
or U807 (N_807,In_1187,N_442);
nor U808 (N_808,In_1812,In_798);
xnor U809 (N_809,In_336,N_563);
xnor U810 (N_810,In_1072,In_1032);
and U811 (N_811,N_505,N_464);
xor U812 (N_812,In_1540,N_352);
or U813 (N_813,N_269,In_1493);
or U814 (N_814,N_379,In_771);
xor U815 (N_815,In_773,N_344);
nand U816 (N_816,N_459,N_782);
xnor U817 (N_817,In_39,N_776);
nand U818 (N_818,N_420,N_618);
or U819 (N_819,In_341,N_159);
and U820 (N_820,N_155,N_274);
nand U821 (N_821,N_711,N_605);
xnor U822 (N_822,N_517,In_643);
nand U823 (N_823,N_411,In_709);
or U824 (N_824,N_654,N_676);
nor U825 (N_825,N_212,In_1224);
nand U826 (N_826,In_51,In_3);
and U827 (N_827,In_1059,In_526);
and U828 (N_828,N_787,In_514);
xnor U829 (N_829,In_531,In_1593);
and U830 (N_830,N_443,In_13);
and U831 (N_831,N_680,In_707);
nand U832 (N_832,In_175,N_282);
nand U833 (N_833,N_732,N_788);
nor U834 (N_834,N_795,In_575);
and U835 (N_835,N_629,N_743);
or U836 (N_836,In_1982,In_446);
and U837 (N_837,N_694,In_581);
or U838 (N_838,In_1554,N_185);
xor U839 (N_839,In_252,N_549);
nor U840 (N_840,In_1885,In_1412);
nand U841 (N_841,N_440,In_1074);
or U842 (N_842,In_1838,In_1622);
xor U843 (N_843,N_503,N_539);
nor U844 (N_844,N_780,N_554);
xor U845 (N_845,N_50,N_525);
or U846 (N_846,N_95,N_198);
xor U847 (N_847,N_724,In_869);
xor U848 (N_848,In_609,In_333);
and U849 (N_849,In_823,N_37);
nand U850 (N_850,N_621,In_1659);
or U851 (N_851,N_725,In_977);
nor U852 (N_852,N_284,In_1144);
and U853 (N_853,N_556,In_866);
nand U854 (N_854,N_195,N_303);
or U855 (N_855,N_772,In_448);
or U856 (N_856,N_626,In_71);
and U857 (N_857,In_1373,N_422);
nor U858 (N_858,N_622,N_216);
and U859 (N_859,In_1728,In_1562);
and U860 (N_860,In_756,N_718);
nor U861 (N_861,In_1172,In_807);
and U862 (N_862,In_759,N_241);
and U863 (N_863,N_135,In_1389);
xor U864 (N_864,N_127,In_586);
or U865 (N_865,N_244,In_1469);
xnor U866 (N_866,N_133,N_401);
and U867 (N_867,In_54,N_449);
nor U868 (N_868,N_470,N_183);
xor U869 (N_869,N_154,N_641);
and U870 (N_870,In_1737,In_1758);
nand U871 (N_871,N_675,N_735);
xnor U872 (N_872,In_494,N_182);
and U873 (N_873,N_52,In_1238);
nor U874 (N_874,N_704,N_367);
or U875 (N_875,In_1357,In_1845);
nor U876 (N_876,In_26,In_943);
nand U877 (N_877,In_1509,In_795);
xnor U878 (N_878,N_435,In_227);
nor U879 (N_879,In_486,In_1624);
xnor U880 (N_880,N_484,N_18);
xnor U881 (N_881,In_1633,N_756);
nand U882 (N_882,In_852,In_560);
and U883 (N_883,N_407,N_74);
and U884 (N_884,N_706,In_1403);
and U885 (N_885,N_738,In_958);
xor U886 (N_886,In_365,N_393);
and U887 (N_887,In_804,In_978);
nor U888 (N_888,N_586,In_204);
or U889 (N_889,N_34,N_794);
or U890 (N_890,In_1486,In_585);
nand U891 (N_891,In_313,In_419);
nor U892 (N_892,In_375,In_617);
or U893 (N_893,N_766,In_729);
or U894 (N_894,N_785,In_1298);
xnor U895 (N_895,N_378,In_298);
nand U896 (N_896,In_556,In_1311);
and U897 (N_897,N_35,In_1602);
nand U898 (N_898,In_416,In_1264);
and U899 (N_899,N_572,N_463);
and U900 (N_900,N_530,In_1160);
and U901 (N_901,N_558,N_466);
xor U902 (N_902,In_1204,In_1362);
nor U903 (N_903,In_1795,In_680);
nand U904 (N_904,In_1891,N_398);
and U905 (N_905,In_480,In_968);
nand U906 (N_906,In_584,N_786);
nor U907 (N_907,In_876,In_1147);
and U908 (N_908,In_1192,In_683);
xor U909 (N_909,N_593,N_317);
nor U910 (N_910,In_1088,N_199);
nand U911 (N_911,In_912,In_219);
nor U912 (N_912,In_1156,In_761);
nand U913 (N_913,In_1842,In_23);
and U914 (N_914,In_1671,N_161);
xnor U915 (N_915,In_1384,In_251);
nand U916 (N_916,In_1772,In_1018);
xor U917 (N_917,N_429,N_335);
xor U918 (N_918,In_1513,In_1478);
or U919 (N_919,N_792,N_746);
xor U920 (N_920,In_1512,N_450);
and U921 (N_921,N_565,N_384);
and U922 (N_922,N_683,N_730);
xor U923 (N_923,N_645,In_443);
nor U924 (N_924,In_939,In_1398);
xor U925 (N_925,In_1555,In_1058);
nor U926 (N_926,In_408,In_43);
nand U927 (N_927,In_1465,N_653);
xnor U928 (N_928,In_532,In_172);
nor U929 (N_929,N_632,N_38);
and U930 (N_930,In_120,N_328);
xnor U931 (N_931,N_528,N_36);
xor U932 (N_932,In_1697,In_793);
nor U933 (N_933,In_675,In_1104);
and U934 (N_934,N_417,N_85);
and U935 (N_935,In_1460,N_3);
nand U936 (N_936,In_861,In_1489);
nor U937 (N_937,In_1990,N_266);
and U938 (N_938,N_221,N_790);
or U939 (N_939,In_1921,In_1296);
xnor U940 (N_940,In_1327,In_84);
xor U941 (N_941,In_482,N_562);
nand U942 (N_942,In_422,In_191);
xor U943 (N_943,In_1203,In_1595);
and U944 (N_944,In_962,In_892);
nor U945 (N_945,N_222,In_1068);
nor U946 (N_946,N_187,In_1491);
xnor U947 (N_947,In_1714,N_739);
nor U948 (N_948,N_288,In_1535);
xnor U949 (N_949,In_960,N_506);
or U950 (N_950,In_1566,In_1267);
and U951 (N_951,In_185,In_1410);
or U952 (N_952,N_650,N_642);
nand U953 (N_953,In_1769,N_532);
nand U954 (N_954,In_1217,N_753);
or U955 (N_955,N_250,N_634);
or U956 (N_956,In_1180,N_147);
nor U957 (N_957,N_751,N_403);
and U958 (N_958,In_1669,In_371);
xor U959 (N_959,In_1009,In_76);
nand U960 (N_960,In_1244,N_309);
xor U961 (N_961,N_823,N_468);
nor U962 (N_962,N_588,N_801);
and U963 (N_963,In_1502,In_402);
nand U964 (N_964,In_764,N_325);
or U965 (N_965,In_294,N_232);
nand U966 (N_966,N_607,N_721);
nand U967 (N_967,N_44,N_775);
xor U968 (N_968,In_1920,In_948);
or U969 (N_969,N_578,N_461);
and U970 (N_970,In_1399,N_602);
xnor U971 (N_971,In_1137,In_395);
or U972 (N_972,In_1852,N_950);
nor U973 (N_973,In_1532,N_919);
and U974 (N_974,N_818,N_498);
nor U975 (N_975,In_1522,In_1339);
or U976 (N_976,N_571,In_1467);
and U977 (N_977,N_830,In_1445);
nand U978 (N_978,In_1212,In_1851);
nor U979 (N_979,In_45,N_640);
xor U980 (N_980,N_707,In_455);
nand U981 (N_981,In_1849,N_536);
and U982 (N_982,N_614,In_1241);
xor U983 (N_983,In_749,N_852);
nand U984 (N_984,In_1825,In_1003);
nand U985 (N_985,N_327,N_604);
and U986 (N_986,In_854,N_271);
or U987 (N_987,N_191,In_548);
nor U988 (N_988,N_124,N_522);
xor U989 (N_989,In_637,N_737);
nand U990 (N_990,N_413,In_647);
nor U991 (N_991,N_434,N_769);
or U992 (N_992,In_1426,In_553);
nor U993 (N_993,In_1236,In_973);
and U994 (N_994,N_444,In_1483);
and U995 (N_995,N_799,In_61);
nor U996 (N_996,N_564,In_244);
nand U997 (N_997,N_651,N_847);
xnor U998 (N_998,N_537,In_1946);
xor U999 (N_999,N_872,In_685);
xor U1000 (N_1000,N_920,N_681);
or U1001 (N_1001,In_940,N_347);
nand U1002 (N_1002,In_58,N_770);
and U1003 (N_1003,In_1552,N_47);
and U1004 (N_1004,N_1,In_1673);
xnor U1005 (N_1005,N_194,N_30);
or U1006 (N_1006,In_768,In_545);
and U1007 (N_1007,In_831,In_1571);
and U1008 (N_1008,N_927,N_942);
xor U1009 (N_1009,In_358,N_906);
or U1010 (N_1010,In_499,N_699);
nand U1011 (N_1011,N_527,In_701);
nand U1012 (N_1012,In_1677,In_604);
nand U1013 (N_1013,N_220,In_891);
nand U1014 (N_1014,N_841,N_909);
and U1015 (N_1015,N_581,N_896);
or U1016 (N_1016,N_386,N_837);
nand U1017 (N_1017,In_895,N_773);
nand U1018 (N_1018,In_1605,N_389);
xor U1019 (N_1019,N_879,N_570);
nor U1020 (N_1020,In_1200,In_936);
or U1021 (N_1021,N_949,In_1996);
or U1022 (N_1022,In_1538,In_328);
nor U1023 (N_1023,In_8,N_861);
nand U1024 (N_1024,N_765,N_700);
nand U1025 (N_1025,In_1221,N_688);
or U1026 (N_1026,N_860,In_56);
xor U1027 (N_1027,N_709,In_1767);
and U1028 (N_1028,In_1863,In_1600);
or U1029 (N_1029,In_1804,N_668);
and U1030 (N_1030,In_690,N_494);
nor U1031 (N_1031,N_875,In_942);
or U1032 (N_1032,N_485,In_780);
nand U1033 (N_1033,In_632,N_501);
nand U1034 (N_1034,N_859,N_491);
xnor U1035 (N_1035,N_878,In_726);
nor U1036 (N_1036,N_933,In_537);
nor U1037 (N_1037,N_710,In_311);
xnor U1038 (N_1038,N_959,In_763);
nor U1039 (N_1039,N_727,N_39);
nand U1040 (N_1040,N_477,In_192);
or U1041 (N_1041,In_1909,N_797);
xnor U1042 (N_1042,In_661,N_870);
nor U1043 (N_1043,N_869,In_1177);
or U1044 (N_1044,In_595,N_867);
or U1045 (N_1045,In_178,In_1829);
or U1046 (N_1046,N_918,In_534);
nand U1047 (N_1047,N_907,N_291);
xnor U1048 (N_1048,In_1400,N_697);
nor U1049 (N_1049,N_832,N_834);
and U1050 (N_1050,N_197,In_591);
nand U1051 (N_1051,In_1855,In_183);
xor U1052 (N_1052,N_428,In_1146);
xor U1053 (N_1053,N_541,In_1017);
nand U1054 (N_1054,In_682,In_740);
or U1055 (N_1055,In_1690,In_1577);
xnor U1056 (N_1056,In_1877,N_366);
or U1057 (N_1057,In_880,In_938);
xnor U1058 (N_1058,In_1676,N_750);
nor U1059 (N_1059,N_720,N_665);
nand U1060 (N_1060,In_1092,N_483);
nor U1061 (N_1061,In_535,N_649);
nor U1062 (N_1062,N_455,N_900);
nor U1063 (N_1063,In_28,In_1642);
and U1064 (N_1064,In_1365,In_232);
and U1065 (N_1065,N_568,N_912);
and U1066 (N_1066,In_1183,N_383);
and U1067 (N_1067,N_105,N_210);
and U1068 (N_1068,In_1276,In_904);
nand U1069 (N_1069,N_755,In_519);
nor U1070 (N_1070,N_533,In_1777);
nor U1071 (N_1071,In_1428,N_757);
nor U1072 (N_1072,In_583,N_293);
xor U1073 (N_1073,In_587,In_785);
nor U1074 (N_1074,N_209,In_1774);
nand U1075 (N_1075,In_1749,N_273);
or U1076 (N_1076,N_858,In_1752);
and U1077 (N_1077,N_943,In_1186);
and U1078 (N_1078,In_1918,In_1258);
and U1079 (N_1079,N_935,In_490);
nand U1080 (N_1080,In_1981,N_423);
and U1081 (N_1081,In_602,In_1448);
or U1082 (N_1082,In_694,N_538);
xor U1083 (N_1083,In_139,N_701);
xor U1084 (N_1084,N_682,In_918);
and U1085 (N_1085,N_206,N_473);
nand U1086 (N_1086,In_143,N_373);
nor U1087 (N_1087,In_1272,N_921);
and U1088 (N_1088,In_11,N_882);
xor U1089 (N_1089,N_695,N_153);
nand U1090 (N_1090,N_885,N_945);
nor U1091 (N_1091,N_804,N_482);
nor U1092 (N_1092,N_415,In_702);
nor U1093 (N_1093,In_528,N_513);
xnor U1094 (N_1094,N_142,In_1666);
and U1095 (N_1095,In_615,In_159);
or U1096 (N_1096,In_608,In_805);
or U1097 (N_1097,N_877,N_758);
and U1098 (N_1098,N_354,In_1973);
nor U1099 (N_1099,N_763,In_366);
nor U1100 (N_1100,N_582,In_741);
xnor U1101 (N_1101,N_890,N_915);
or U1102 (N_1102,In_1360,N_445);
or U1103 (N_1103,In_282,N_355);
and U1104 (N_1104,In_146,N_178);
xor U1105 (N_1105,In_920,N_319);
xor U1106 (N_1106,N_798,N_851);
xor U1107 (N_1107,N_904,In_1692);
and U1108 (N_1108,N_612,N_10);
and U1109 (N_1109,N_956,N_722);
xor U1110 (N_1110,N_844,N_467);
xor U1111 (N_1111,N_68,In_835);
nand U1112 (N_1112,N_809,N_315);
xor U1113 (N_1113,N_914,In_1397);
nand U1114 (N_1114,In_15,In_4);
nand U1115 (N_1115,In_1969,N_729);
or U1116 (N_1116,N_613,In_881);
xor U1117 (N_1117,N_454,In_1456);
or U1118 (N_1118,N_623,In_1746);
and U1119 (N_1119,In_1833,N_65);
xor U1120 (N_1120,N_693,In_290);
and U1121 (N_1121,N_1063,N_666);
and U1122 (N_1122,In_1385,In_573);
and U1123 (N_1123,N_726,In_1459);
nor U1124 (N_1124,N_502,N_268);
nor U1125 (N_1125,N_171,N_1068);
xor U1126 (N_1126,In_1055,In_1355);
nand U1127 (N_1127,In_803,N_703);
nand U1128 (N_1128,In_991,N_898);
nand U1129 (N_1129,N_911,In_829);
nor U1130 (N_1130,N_1042,In_1245);
or U1131 (N_1131,In_1121,In_1411);
and U1132 (N_1132,N_638,In_423);
or U1133 (N_1133,In_357,In_1934);
nand U1134 (N_1134,N_759,In_1255);
nand U1135 (N_1135,N_643,N_987);
xor U1136 (N_1136,N_635,In_1747);
nor U1137 (N_1137,In_57,N_1036);
nand U1138 (N_1138,In_1892,N_329);
or U1139 (N_1139,In_1322,In_262);
or U1140 (N_1140,N_965,N_836);
and U1141 (N_1141,N_925,N_840);
nor U1142 (N_1142,N_1116,In_1553);
nor U1143 (N_1143,N_886,In_1871);
nand U1144 (N_1144,N_864,N_227);
or U1145 (N_1145,In_620,N_843);
xor U1146 (N_1146,In_1198,N_781);
xor U1147 (N_1147,N_356,In_885);
nand U1148 (N_1148,In_856,N_448);
and U1149 (N_1149,In_1294,In_1051);
or U1150 (N_1150,N_545,In_1744);
and U1151 (N_1151,N_808,In_133);
nor U1152 (N_1152,N_1034,N_1070);
nand U1153 (N_1153,N_137,N_671);
or U1154 (N_1154,In_788,N_940);
nand U1155 (N_1155,In_1563,N_1023);
xor U1156 (N_1156,In_1131,In_1531);
nand U1157 (N_1157,N_360,N_1067);
and U1158 (N_1158,N_1010,N_761);
and U1159 (N_1159,N_592,N_944);
and U1160 (N_1160,N_982,N_819);
or U1161 (N_1161,N_939,N_395);
nor U1162 (N_1162,N_553,N_1054);
nand U1163 (N_1163,In_655,N_1015);
xnor U1164 (N_1164,N_771,In_1038);
xor U1165 (N_1165,In_1181,N_985);
and U1166 (N_1166,N_767,N_916);
or U1167 (N_1167,N_341,N_1117);
or U1168 (N_1168,N_1009,N_1073);
or U1169 (N_1169,N_1077,In_405);
and U1170 (N_1170,In_1858,N_741);
nand U1171 (N_1171,N_76,N_504);
or U1172 (N_1172,N_560,In_434);
or U1173 (N_1173,N_917,In_1803);
and U1174 (N_1174,N_644,N_662);
and U1175 (N_1175,In_1309,In_1733);
nand U1176 (N_1176,N_460,N_11);
or U1177 (N_1177,N_262,N_803);
nor U1178 (N_1178,N_40,N_104);
nand U1179 (N_1179,In_1166,In_400);
and U1180 (N_1180,In_1291,In_310);
nor U1181 (N_1181,N_376,In_488);
or U1182 (N_1182,In_1443,N_236);
or U1183 (N_1183,In_860,N_1052);
nand U1184 (N_1184,In_1349,In_1809);
nand U1185 (N_1185,N_17,In_223);
xor U1186 (N_1186,In_956,In_1505);
nand U1187 (N_1187,N_365,N_323);
xor U1188 (N_1188,N_575,N_1097);
xnor U1189 (N_1189,N_224,N_1005);
xnor U1190 (N_1190,In_542,In_914);
and U1191 (N_1191,In_276,N_1114);
or U1192 (N_1192,N_1085,In_1012);
or U1193 (N_1193,N_692,In_715);
nor U1194 (N_1194,N_1019,N_796);
or U1195 (N_1195,In_1451,N_815);
xnor U1196 (N_1196,In_1886,In_164);
or U1197 (N_1197,N_53,N_1028);
nand U1198 (N_1198,In_479,In_1705);
nand U1199 (N_1199,In_1987,In_1022);
nand U1200 (N_1200,In_951,In_1641);
nor U1201 (N_1201,N_817,N_975);
and U1202 (N_1202,N_163,N_1024);
nand U1203 (N_1203,N_974,N_923);
xnor U1204 (N_1204,In_1413,N_239);
or U1205 (N_1205,In_1423,N_1086);
and U1206 (N_1206,N_762,N_121);
or U1207 (N_1207,N_1043,N_249);
xnor U1208 (N_1208,In_527,N_784);
and U1209 (N_1209,In_718,In_1472);
nor U1210 (N_1210,N_887,In_406);
xnor U1211 (N_1211,In_87,In_1346);
and U1212 (N_1212,N_313,In_261);
nand U1213 (N_1213,N_812,N_447);
and U1214 (N_1214,In_385,In_1019);
or U1215 (N_1215,In_112,N_1058);
nor U1216 (N_1216,N_597,In_672);
or U1217 (N_1217,N_521,N_1006);
and U1218 (N_1218,N_1105,In_25);
xnor U1219 (N_1219,N_807,In_1482);
nor U1220 (N_1220,N_1104,In_1277);
nand U1221 (N_1221,N_991,In_1805);
or U1222 (N_1222,In_20,In_1285);
xnor U1223 (N_1223,N_717,N_774);
and U1224 (N_1224,N_509,N_849);
nor U1225 (N_1225,N_857,N_92);
nand U1226 (N_1226,N_984,N_873);
or U1227 (N_1227,N_333,N_514);
nor U1228 (N_1228,In_1300,In_41);
and U1229 (N_1229,In_460,In_1283);
and U1230 (N_1230,N_745,In_1850);
nor U1231 (N_1231,In_884,N_231);
nand U1232 (N_1232,N_910,N_59);
and U1233 (N_1233,N_778,N_674);
nand U1234 (N_1234,In_1499,In_216);
and U1235 (N_1235,In_468,In_452);
and U1236 (N_1236,In_1528,In_1966);
or U1237 (N_1237,N_292,N_999);
nor U1238 (N_1238,N_213,N_677);
or U1239 (N_1239,In_666,N_1046);
and U1240 (N_1240,In_747,In_1490);
or U1241 (N_1241,N_791,N_1002);
xor U1242 (N_1242,N_793,N_648);
xor U1243 (N_1243,N_281,N_736);
or U1244 (N_1244,In_725,In_1813);
and U1245 (N_1245,N_749,N_689);
nor U1246 (N_1246,N_691,In_981);
xor U1247 (N_1247,In_181,In_1240);
or U1248 (N_1248,N_789,In_1262);
and U1249 (N_1249,N_1061,In_1023);
nand U1250 (N_1250,N_639,N_576);
and U1251 (N_1251,In_1427,In_148);
nand U1252 (N_1252,N_712,In_415);
xnor U1253 (N_1253,N_436,In_857);
or U1254 (N_1254,In_1715,In_676);
or U1255 (N_1255,In_1802,In_1155);
nand U1256 (N_1256,N_663,N_577);
nand U1257 (N_1257,N_56,In_1175);
nand U1258 (N_1258,N_219,In_677);
xor U1259 (N_1259,In_1099,In_1433);
and U1260 (N_1260,N_768,N_876);
xor U1261 (N_1261,N_862,N_500);
nand U1262 (N_1262,In_1874,N_270);
xor U1263 (N_1263,In_381,N_1111);
xor U1264 (N_1264,In_875,N_678);
nand U1265 (N_1265,In_930,N_33);
and U1266 (N_1266,In_1942,In_1042);
xor U1267 (N_1267,N_723,N_286);
or U1268 (N_1268,In_713,N_814);
and U1269 (N_1269,N_1090,N_802);
nor U1270 (N_1270,In_970,In_1307);
and U1271 (N_1271,In_355,N_977);
nand U1272 (N_1272,N_601,In_1292);
or U1273 (N_1273,In_68,In_1033);
or U1274 (N_1274,In_1890,N_1069);
and U1275 (N_1275,In_1234,N_535);
or U1276 (N_1276,In_984,N_1091);
and U1277 (N_1277,N_658,In_1922);
and U1278 (N_1278,N_215,In_1681);
and U1279 (N_1279,N_150,In_775);
nand U1280 (N_1280,N_1049,In_1559);
or U1281 (N_1281,N_888,N_1164);
and U1282 (N_1282,N_608,N_1135);
or U1283 (N_1283,In_347,In_511);
xor U1284 (N_1284,N_932,In_503);
nand U1285 (N_1285,N_752,N_1027);
xnor U1286 (N_1286,N_1098,N_138);
nand U1287 (N_1287,In_1073,N_546);
nand U1288 (N_1288,N_1025,In_1872);
nor U1289 (N_1289,N_705,In_934);
nor U1290 (N_1290,N_967,N_947);
xnor U1291 (N_1291,N_958,N_1158);
xnor U1292 (N_1292,In_104,N_1195);
or U1293 (N_1293,In_1315,In_1304);
and U1294 (N_1294,N_330,N_661);
nor U1295 (N_1295,N_80,N_567);
nor U1296 (N_1296,N_1250,N_359);
nor U1297 (N_1297,N_246,N_657);
xor U1298 (N_1298,N_471,N_1096);
nor U1299 (N_1299,N_172,N_1271);
xor U1300 (N_1300,N_1230,N_26);
nand U1301 (N_1301,N_83,In_1843);
nor U1302 (N_1302,In_1938,In_315);
and U1303 (N_1303,N_760,N_670);
or U1304 (N_1304,N_476,N_957);
or U1305 (N_1305,In_1931,N_805);
or U1306 (N_1306,In_1837,In_1533);
xnor U1307 (N_1307,In_242,N_1088);
xnor U1308 (N_1308,N_1139,N_871);
nand U1309 (N_1309,In_732,N_201);
xnor U1310 (N_1310,In_384,In_1836);
nand U1311 (N_1311,N_824,N_1269);
nand U1312 (N_1312,In_689,In_1957);
xnor U1313 (N_1313,N_557,In_913);
nand U1314 (N_1314,In_704,N_1132);
or U1315 (N_1315,N_1080,In_681);
xor U1316 (N_1316,N_1267,N_708);
and U1317 (N_1317,In_611,In_1118);
nor U1318 (N_1318,N_606,In_158);
nor U1319 (N_1319,N_1126,N_986);
xor U1320 (N_1320,N_1236,N_822);
and U1321 (N_1321,In_800,N_1197);
nor U1322 (N_1322,N_936,N_152);
and U1323 (N_1323,In_839,N_385);
xor U1324 (N_1324,N_1014,N_1194);
xnor U1325 (N_1325,N_1272,N_839);
nand U1326 (N_1326,N_1118,N_1044);
nor U1327 (N_1327,N_1153,N_783);
xor U1328 (N_1328,N_660,N_1039);
or U1329 (N_1329,In_1529,In_264);
or U1330 (N_1330,In_1548,In_635);
xor U1331 (N_1331,N_853,N_696);
or U1332 (N_1332,N_1225,In_1356);
nand U1333 (N_1333,N_981,N_591);
xnor U1334 (N_1334,N_929,N_1112);
nand U1335 (N_1335,N_318,N_1037);
and U1336 (N_1336,N_960,N_1262);
nand U1337 (N_1337,In_1590,In_1178);
and U1338 (N_1338,N_1166,N_1120);
or U1339 (N_1339,N_952,In_256);
nand U1340 (N_1340,N_1020,N_1242);
xor U1341 (N_1341,In_727,N_1013);
or U1342 (N_1342,N_81,In_1979);
nand U1343 (N_1343,N_744,N_1012);
nor U1344 (N_1344,N_410,N_1134);
nor U1345 (N_1345,N_1001,In_327);
and U1346 (N_1346,N_1065,N_838);
nor U1347 (N_1347,N_913,N_1254);
and U1348 (N_1348,In_153,N_1273);
or U1349 (N_1349,N_880,In_738);
nand U1350 (N_1350,In_1391,In_1846);
and U1351 (N_1351,N_363,N_1130);
xor U1352 (N_1352,N_180,In_208);
xor U1353 (N_1353,In_1342,N_1169);
or U1354 (N_1354,N_1220,N_1183);
or U1355 (N_1355,N_1182,N_338);
or U1356 (N_1356,N_1084,In_784);
and U1357 (N_1357,N_458,In_746);
or U1358 (N_1358,In_1001,N_731);
xor U1359 (N_1359,N_446,N_866);
nor U1360 (N_1360,N_679,N_139);
nor U1361 (N_1361,N_478,In_414);
or U1362 (N_1362,In_284,In_1434);
or U1363 (N_1363,N_931,In_425);
nor U1364 (N_1364,N_1011,N_1258);
xor U1365 (N_1365,In_1625,N_1179);
and U1366 (N_1366,N_656,In_1323);
and U1367 (N_1367,N_979,In_1543);
and U1368 (N_1368,In_1268,N_433);
or U1369 (N_1369,N_322,N_1201);
xor U1370 (N_1370,N_438,N_995);
nor U1371 (N_1371,N_990,N_1162);
and U1372 (N_1372,N_1055,N_1071);
nand U1373 (N_1373,In_107,N_1243);
or U1374 (N_1374,N_713,N_54);
nand U1375 (N_1375,N_1108,N_901);
nor U1376 (N_1376,N_1261,N_968);
nand U1377 (N_1377,N_1178,In_1674);
nand U1378 (N_1378,N_924,In_471);
nor U1379 (N_1379,N_1121,N_1032);
and U1380 (N_1380,N_1150,N_229);
nand U1381 (N_1381,N_611,N_1053);
nor U1382 (N_1382,N_892,N_294);
nor U1383 (N_1383,In_250,In_830);
nand U1384 (N_1384,N_1147,N_988);
nor U1385 (N_1385,In_1729,N_1137);
nor U1386 (N_1386,N_1141,N_166);
nor U1387 (N_1387,In_838,N_358);
nand U1388 (N_1388,N_1109,In_640);
xor U1389 (N_1389,N_684,In_149);
or U1390 (N_1390,N_1270,In_30);
nand U1391 (N_1391,N_972,N_345);
nand U1392 (N_1392,N_1040,In_508);
xnor U1393 (N_1393,N_46,In_792);
and U1394 (N_1394,N_1245,N_1207);
and U1395 (N_1395,N_1246,N_664);
nor U1396 (N_1396,In_1011,In_234);
nand U1397 (N_1397,N_1159,In_1695);
or U1398 (N_1398,In_147,N_1209);
nand U1399 (N_1399,In_1623,N_1205);
and U1400 (N_1400,N_14,N_28);
nand U1401 (N_1401,N_1101,N_976);
xor U1402 (N_1402,N_714,N_821);
nor U1403 (N_1403,N_1004,N_1155);
and U1404 (N_1404,N_1008,N_902);
nand U1405 (N_1405,In_475,N_800);
and U1406 (N_1406,In_714,N_1232);
nor U1407 (N_1407,In_506,N_903);
nand U1408 (N_1408,N_845,N_926);
or U1409 (N_1409,N_964,N_451);
nand U1410 (N_1410,In_102,N_116);
xnor U1411 (N_1411,N_728,N_1208);
nand U1412 (N_1412,In_1064,N_1075);
nor U1413 (N_1413,N_820,N_1184);
and U1414 (N_1414,N_955,In_1707);
nand U1415 (N_1415,N_969,N_518);
xnor U1416 (N_1416,N_754,N_1277);
and U1417 (N_1417,N_1268,N_1051);
nand U1418 (N_1418,In_1261,N_1022);
or U1419 (N_1419,In_512,N_1156);
and U1420 (N_1420,N_1196,In_826);
or U1421 (N_1421,In_254,N_1279);
nor U1422 (N_1422,In_555,N_1248);
nand U1423 (N_1423,N_589,N_631);
xor U1424 (N_1424,In_700,N_633);
nand U1425 (N_1425,N_1180,In_833);
and U1426 (N_1426,N_1172,N_1266);
xor U1427 (N_1427,N_584,N_953);
or U1428 (N_1428,N_1017,N_1095);
xor U1429 (N_1429,N_715,N_346);
or U1430 (N_1430,N_1237,N_240);
nor U1431 (N_1431,In_848,N_716);
xor U1432 (N_1432,N_874,N_1144);
and U1433 (N_1433,N_948,In_664);
xnor U1434 (N_1434,N_188,In_878);
nand U1435 (N_1435,In_505,In_1193);
nor U1436 (N_1436,N_1059,N_1218);
or U1437 (N_1437,N_826,N_1175);
xnor U1438 (N_1438,N_897,N_1226);
xnor U1439 (N_1439,N_189,N_1045);
or U1440 (N_1440,N_238,N_508);
nor U1441 (N_1441,In_1335,N_1211);
xor U1442 (N_1442,N_1347,N_1393);
nand U1443 (N_1443,N_1129,N_828);
and U1444 (N_1444,N_1124,In_1248);
nand U1445 (N_1445,N_1081,N_1078);
xnor U1446 (N_1446,In_119,N_1405);
or U1447 (N_1447,In_1424,In_898);
nand U1448 (N_1448,In_293,N_316);
xnor U1449 (N_1449,N_748,N_1186);
nor U1450 (N_1450,N_1388,N_1157);
xor U1451 (N_1451,In_952,N_1115);
or U1452 (N_1452,In_1247,N_1348);
nand U1453 (N_1453,In_1364,N_1328);
xor U1454 (N_1454,N_647,N_1021);
nand U1455 (N_1455,N_619,N_331);
or U1456 (N_1456,N_1173,N_381);
nor U1457 (N_1457,N_1033,N_863);
or U1458 (N_1458,N_1285,N_1312);
or U1459 (N_1459,N_1072,N_1185);
nor U1460 (N_1460,N_934,N_702);
nand U1461 (N_1461,N_1389,N_1386);
or U1462 (N_1462,In_1266,N_1333);
and U1463 (N_1463,N_1103,In_325);
nand U1464 (N_1464,In_668,N_881);
nor U1465 (N_1465,In_734,N_655);
and U1466 (N_1466,N_1133,In_1138);
nor U1467 (N_1467,N_202,N_1302);
and U1468 (N_1468,N_779,N_1231);
nand U1469 (N_1469,N_1062,N_764);
and U1470 (N_1470,N_524,In_1379);
and U1471 (N_1471,N_71,In_1993);
and U1472 (N_1472,N_1321,N_406);
nor U1473 (N_1473,In_1076,N_1311);
xor U1474 (N_1474,N_548,N_992);
nand U1475 (N_1475,N_1407,N_1341);
xnor U1476 (N_1476,In_1564,N_1047);
nand U1477 (N_1477,N_811,N_599);
xor U1478 (N_1478,N_399,N_1221);
xnor U1479 (N_1479,N_894,In_163);
and U1480 (N_1480,N_637,In_1980);
nor U1481 (N_1481,In_670,N_1355);
nor U1482 (N_1482,N_1235,N_1057);
and U1483 (N_1483,N_1368,N_895);
nand U1484 (N_1484,N_980,N_1359);
xnor U1485 (N_1485,In_1242,N_742);
nor U1486 (N_1486,N_1146,N_1434);
and U1487 (N_1487,N_1249,N_424);
xor U1488 (N_1488,In_364,N_1259);
nand U1489 (N_1489,N_1050,N_1357);
nor U1490 (N_1490,N_1190,N_1174);
nand U1491 (N_1491,In_625,N_1122);
nor U1492 (N_1492,N_1399,N_951);
and U1493 (N_1493,In_886,N_1413);
nand U1494 (N_1494,N_1131,N_1430);
xor U1495 (N_1495,In_1065,N_1056);
or U1496 (N_1496,N_1398,In_1912);
and U1497 (N_1497,N_1224,N_1374);
or U1498 (N_1498,N_1278,N_1344);
nand U1499 (N_1499,N_1257,In_703);
nor U1500 (N_1500,In_1814,N_1031);
xnor U1501 (N_1501,In_1111,N_1260);
xnor U1502 (N_1502,In_214,N_1038);
nand U1503 (N_1503,N_432,N_129);
or U1504 (N_1504,N_685,N_523);
xor U1505 (N_1505,N_1286,N_1330);
xnor U1506 (N_1506,N_983,N_686);
xor U1507 (N_1507,N_1030,N_1200);
or U1508 (N_1508,In_1601,N_962);
or U1509 (N_1509,N_497,N_1353);
or U1510 (N_1510,N_1240,N_1188);
or U1511 (N_1511,N_1187,N_733);
and U1512 (N_1512,In_626,In_1875);
xnor U1513 (N_1513,N_1106,N_1306);
xnor U1514 (N_1514,N_908,In_1816);
nor U1515 (N_1515,N_1265,N_846);
xnor U1516 (N_1516,N_646,N_1029);
nand U1517 (N_1517,N_1066,N_254);
nand U1518 (N_1518,N_884,In_1684);
and U1519 (N_1519,In_225,N_889);
nand U1520 (N_1520,In_266,N_777);
or U1521 (N_1521,N_1329,N_1064);
nor U1522 (N_1522,N_1154,N_1397);
or U1523 (N_1523,N_287,In_295);
xnor U1524 (N_1524,N_1391,N_1412);
and U1525 (N_1525,In_483,N_810);
nor U1526 (N_1526,N_1192,In_1937);
nor U1527 (N_1527,N_1214,N_1373);
or U1528 (N_1528,N_1234,N_625);
or U1529 (N_1529,N_993,N_734);
nor U1530 (N_1530,N_1408,N_1007);
or U1531 (N_1531,N_1151,In_331);
nor U1532 (N_1532,In_1876,N_439);
xnor U1533 (N_1533,N_672,N_1395);
nor U1534 (N_1534,N_1256,N_1315);
xor U1535 (N_1535,N_1228,N_1167);
or U1536 (N_1536,N_1251,N_1294);
and U1537 (N_1537,N_1079,N_1168);
xnor U1538 (N_1538,N_996,N_905);
nand U1539 (N_1539,N_1171,N_1410);
or U1540 (N_1540,N_1204,N_1216);
or U1541 (N_1541,N_1301,N_1283);
and U1542 (N_1542,N_1210,In_949);
xor U1543 (N_1543,N_1060,N_1018);
or U1544 (N_1544,N_1390,N_1100);
xor U1545 (N_1545,N_1354,N_223);
nor U1546 (N_1546,N_961,N_719);
or U1547 (N_1547,In_469,N_973);
or U1548 (N_1548,N_854,In_533);
or U1549 (N_1549,In_592,In_70);
and U1550 (N_1550,N_1381,N_1423);
nor U1551 (N_1551,In_1792,N_1418);
xnor U1552 (N_1552,In_1539,N_1000);
nand U1553 (N_1553,N_1202,N_1299);
or U1554 (N_1554,N_1316,N_488);
or U1555 (N_1555,N_1327,N_1140);
xnor U1556 (N_1556,N_1342,In_1040);
nor U1557 (N_1557,N_1119,N_519);
nor U1558 (N_1558,N_1439,In_222);
nor U1559 (N_1559,N_687,In_950);
or U1560 (N_1560,N_698,N_1343);
and U1561 (N_1561,N_1138,N_1244);
nand U1562 (N_1562,N_1366,N_1284);
xor U1563 (N_1563,N_1145,N_624);
nand U1564 (N_1564,N_1107,N_659);
nor U1565 (N_1565,In_633,N_941);
and U1566 (N_1566,N_349,N_1414);
or U1567 (N_1567,N_457,N_1350);
and U1568 (N_1568,N_1308,N_1349);
nor U1569 (N_1569,In_1214,N_1384);
or U1570 (N_1570,N_1361,N_1113);
xor U1571 (N_1571,N_1016,In_323);
or U1572 (N_1572,In_607,N_1199);
nand U1573 (N_1573,N_1370,N_1396);
and U1574 (N_1574,N_989,N_842);
and U1575 (N_1575,N_534,N_1403);
and U1576 (N_1576,N_1400,N_1035);
and U1577 (N_1577,N_1127,N_569);
nand U1578 (N_1578,N_1252,N_1337);
or U1579 (N_1579,N_954,N_1128);
nand U1580 (N_1580,In_168,In_1235);
xor U1581 (N_1581,N_1429,N_1345);
or U1582 (N_1582,N_1255,N_134);
xnor U1583 (N_1583,N_1143,N_1300);
or U1584 (N_1584,In_547,N_1048);
xor U1585 (N_1585,N_1305,In_209);
or U1586 (N_1586,N_1191,N_856);
nor U1587 (N_1587,N_1074,N_1287);
or U1588 (N_1588,N_1082,N_1417);
or U1589 (N_1589,N_1322,N_1142);
nor U1590 (N_1590,N_1189,N_928);
nor U1591 (N_1591,N_1026,In_307);
and U1592 (N_1592,N_1334,In_1320);
and U1593 (N_1593,N_1087,N_628);
xnor U1594 (N_1594,N_1379,In_653);
nor U1595 (N_1595,N_835,N_1281);
nand U1596 (N_1596,N_1339,N_1402);
or U1597 (N_1597,N_1416,N_946);
nand U1598 (N_1598,In_1636,N_516);
and U1599 (N_1599,N_1276,N_1365);
or U1600 (N_1600,N_1099,N_1471);
and U1601 (N_1601,N_1415,N_1093);
and U1602 (N_1602,N_1579,N_833);
nand U1603 (N_1603,N_937,N_1238);
or U1604 (N_1604,N_162,N_1488);
and U1605 (N_1605,N_978,N_1376);
xor U1606 (N_1606,N_1590,N_1161);
nand U1607 (N_1607,N_1222,N_806);
xor U1608 (N_1608,N_1452,N_1596);
nand U1609 (N_1609,N_1537,N_111);
nor U1610 (N_1610,N_994,N_1346);
nand U1611 (N_1611,N_1432,N_117);
and U1612 (N_1612,N_1292,N_1497);
xor U1613 (N_1613,N_1247,In_1588);
and U1614 (N_1614,N_1505,In_241);
and U1615 (N_1615,N_1371,N_1288);
nand U1616 (N_1616,N_1480,In_1024);
xor U1617 (N_1617,N_66,N_1123);
and U1618 (N_1618,N_1372,N_1485);
xor U1619 (N_1619,In_1345,N_1451);
nand U1620 (N_1620,N_1470,N_1148);
nand U1621 (N_1621,N_1521,N_492);
or U1622 (N_1622,In_529,In_281);
xor U1623 (N_1623,N_938,N_585);
and U1624 (N_1624,In_706,N_1431);
nor U1625 (N_1625,N_1385,N_1442);
and U1626 (N_1626,N_1003,N_1296);
or U1627 (N_1627,N_1102,N_831);
and U1628 (N_1628,N_1392,N_1176);
and U1629 (N_1629,N_1436,In_151);
xor U1630 (N_1630,N_1518,N_1572);
nor U1631 (N_1631,N_1465,In_926);
or U1632 (N_1632,N_1581,N_1571);
and U1633 (N_1633,N_1586,N_1110);
xnor U1634 (N_1634,N_1177,N_1464);
nor U1635 (N_1635,N_1457,N_1553);
xor U1636 (N_1636,N_1562,N_1549);
xnor U1637 (N_1637,N_1377,N_893);
xnor U1638 (N_1638,N_1543,N_1303);
or U1639 (N_1639,N_515,N_1420);
nor U1640 (N_1640,N_1203,In_1343);
and U1641 (N_1641,N_1421,In_1860);
or U1642 (N_1642,N_971,N_1263);
xor U1643 (N_1643,N_377,N_865);
nor U1644 (N_1644,N_1282,N_1486);
nor U1645 (N_1645,N_1483,N_855);
xnor U1646 (N_1646,N_1510,N_667);
nor U1647 (N_1647,N_1534,In_1719);
or U1648 (N_1648,In_1853,N_1599);
nor U1649 (N_1649,N_1498,N_1583);
and U1650 (N_1650,N_1472,N_922);
nor U1651 (N_1651,N_1484,N_1567);
nand U1652 (N_1652,N_1516,N_1219);
nand U1653 (N_1653,N_1360,N_1125);
nor U1654 (N_1654,N_1364,N_1489);
and U1655 (N_1655,N_1428,N_1519);
or U1656 (N_1656,N_1574,N_1542);
nand U1657 (N_1657,N_1499,N_1554);
xor U1658 (N_1658,N_1506,In_1208);
nand U1659 (N_1659,N_1314,N_336);
nor U1660 (N_1660,N_1493,N_1313);
and U1661 (N_1661,N_1476,N_1587);
xnor U1662 (N_1662,N_1383,N_1435);
nor U1663 (N_1663,N_1193,N_1356);
xnor U1664 (N_1664,N_1229,In_1778);
xor U1665 (N_1665,N_1475,N_1490);
xor U1666 (N_1666,N_1455,N_1495);
and U1667 (N_1667,N_1297,In_751);
xor U1668 (N_1668,N_1533,N_1411);
and U1669 (N_1669,N_1509,N_1541);
or U1670 (N_1670,N_1409,N_848);
and U1671 (N_1671,N_1181,N_1426);
or U1672 (N_1672,N_630,N_1367);
nand U1673 (N_1673,In_1438,N_1578);
or U1674 (N_1674,N_1500,N_1598);
nor U1675 (N_1675,N_1401,N_1478);
nor U1676 (N_1676,N_1441,N_1212);
nand U1677 (N_1677,N_1275,N_1338);
nor U1678 (N_1678,N_1589,N_1404);
nor U1679 (N_1679,N_963,In_1679);
nand U1680 (N_1680,N_930,In_309);
and U1681 (N_1681,N_1526,N_1592);
or U1682 (N_1682,N_1215,N_559);
nand U1683 (N_1683,N_1566,N_1570);
nand U1684 (N_1684,In_1396,N_1445);
and U1685 (N_1685,N_1515,N_353);
nand U1686 (N_1686,N_1425,In_442);
nor U1687 (N_1687,N_615,N_1468);
nor U1688 (N_1688,N_1380,N_1536);
nor U1689 (N_1689,In_1971,N_1461);
xor U1690 (N_1690,In_1782,In_1536);
xnor U1691 (N_1691,N_1595,N_1325);
or U1692 (N_1692,N_1459,N_1443);
xor U1693 (N_1693,N_1473,In_495);
and U1694 (N_1694,N_1508,N_816);
and U1695 (N_1695,N_1593,N_1513);
nand U1696 (N_1696,N_1503,N_1163);
or U1697 (N_1697,N_1565,N_1462);
nand U1698 (N_1698,N_850,In_862);
and U1699 (N_1699,N_1331,N_1076);
and U1700 (N_1700,N_1568,N_1479);
nand U1701 (N_1701,N_1469,N_1466);
nor U1702 (N_1702,N_1531,N_1547);
xor U1703 (N_1703,N_1501,N_1556);
or U1704 (N_1704,In_472,N_1363);
xnor U1705 (N_1705,N_1326,N_1213);
or U1706 (N_1706,N_1577,N_1290);
nor U1707 (N_1707,In_1608,N_1481);
xor U1708 (N_1708,N_1561,N_1540);
and U1709 (N_1709,N_1569,N_1433);
xor U1710 (N_1710,N_151,N_1233);
xnor U1711 (N_1711,N_1324,N_1546);
nor U1712 (N_1712,N_1149,N_673);
or U1713 (N_1713,In_1159,N_1575);
xor U1714 (N_1714,N_1422,In_306);
xnor U1715 (N_1715,N_1089,N_998);
nand U1716 (N_1716,N_226,N_1447);
nor U1717 (N_1717,N_1352,N_1438);
and U1718 (N_1718,N_1545,N_1482);
nor U1719 (N_1719,N_1559,N_1539);
nand U1720 (N_1720,N_1477,N_1467);
or U1721 (N_1721,N_827,N_1588);
and U1722 (N_1722,N_1557,N_1309);
and U1723 (N_1723,N_1585,N_1239);
nor U1724 (N_1724,N_1358,N_883);
xnor U1725 (N_1725,In_760,N_308);
xor U1726 (N_1726,N_1351,N_1576);
and U1727 (N_1727,In_1125,N_1323);
nor U1728 (N_1728,In_1643,N_1253);
xnor U1729 (N_1729,N_1440,N_543);
nand U1730 (N_1730,In_858,N_1584);
and U1731 (N_1731,N_110,N_1524);
and U1732 (N_1732,N_1563,In_332);
xnor U1733 (N_1733,N_1512,N_1504);
xnor U1734 (N_1734,N_1597,N_1591);
nor U1735 (N_1735,N_1544,N_1555);
xnor U1736 (N_1736,N_1552,In_206);
xor U1737 (N_1737,N_1487,In_52);
and U1738 (N_1738,N_1335,N_285);
or U1739 (N_1739,N_1444,N_1092);
or U1740 (N_1740,N_1295,N_1502);
or U1741 (N_1741,N_1454,In_1951);
xor U1742 (N_1742,N_1525,N_1560);
nand U1743 (N_1743,N_1319,N_1532);
xnor U1744 (N_1744,N_825,N_1528);
xor U1745 (N_1745,N_1291,N_1507);
or U1746 (N_1746,N_1582,N_1520);
nor U1747 (N_1747,N_966,N_566);
xnor U1748 (N_1748,N_1280,N_1514);
or U1749 (N_1749,N_1474,N_1463);
nand U1750 (N_1750,N_1427,N_1136);
nand U1751 (N_1751,N_1317,N_899);
xor U1752 (N_1752,N_1558,In_33);
or U1753 (N_1753,N_620,N_1538);
xor U1754 (N_1754,N_829,N_1550);
nand U1755 (N_1755,N_1448,N_1453);
and U1756 (N_1756,N_1458,N_1530);
and U1757 (N_1757,N_1320,N_1406);
nand U1758 (N_1758,N_1382,N_1094);
xnor U1759 (N_1759,N_1580,N_1394);
and U1760 (N_1760,N_1754,N_1644);
nor U1761 (N_1761,N_1664,In_65);
nor U1762 (N_1762,N_1749,N_1631);
and U1763 (N_1763,N_1170,N_1665);
nor U1764 (N_1764,N_1611,N_1692);
and U1765 (N_1765,N_1710,N_1437);
xor U1766 (N_1766,N_1223,N_1641);
nand U1767 (N_1767,N_1640,N_1449);
and U1768 (N_1768,N_1672,N_1696);
and U1769 (N_1769,N_1446,N_1728);
or U1770 (N_1770,N_1636,N_1491);
or U1771 (N_1771,In_724,N_1711);
nor U1772 (N_1772,N_1683,N_1609);
xor U1773 (N_1773,N_1548,N_1751);
xor U1774 (N_1774,N_1340,N_1733);
nor U1775 (N_1775,N_1699,In_1324);
or U1776 (N_1776,N_1617,N_499);
and U1777 (N_1777,N_1714,N_1707);
nor U1778 (N_1778,N_1635,N_362);
xor U1779 (N_1779,N_1613,N_1689);
nor U1780 (N_1780,N_1627,N_1667);
nand U1781 (N_1781,N_1731,N_1307);
or U1782 (N_1782,N_1669,N_1676);
nand U1783 (N_1783,In_631,N_1289);
nor U1784 (N_1784,N_1293,N_1713);
or U1785 (N_1785,N_1652,N_1573);
nor U1786 (N_1786,N_1628,N_1691);
xnor U1787 (N_1787,N_1725,N_1419);
nand U1788 (N_1788,N_1715,N_1626);
or U1789 (N_1789,N_1523,N_1621);
nor U1790 (N_1790,N_1601,N_1651);
or U1791 (N_1791,N_1511,N_1638);
and U1792 (N_1792,N_1647,N_1639);
nand U1793 (N_1793,N_1650,N_1670);
nand U1794 (N_1794,N_1310,N_1673);
nor U1795 (N_1795,N_1606,N_1758);
xor U1796 (N_1796,N_1722,N_1535);
and U1797 (N_1797,N_1494,N_1727);
or U1798 (N_1798,N_1732,N_1622);
nor U1799 (N_1799,N_1678,N_1083);
xor U1800 (N_1800,N_1736,N_1643);
and U1801 (N_1801,N_1619,In_1048);
nand U1802 (N_1802,N_1594,N_1706);
nor U1803 (N_1803,N_1752,N_1739);
nand U1804 (N_1804,N_1656,N_1757);
nand U1805 (N_1805,N_1682,N_1740);
nor U1806 (N_1806,N_1700,N_1608);
nand U1807 (N_1807,In_1523,N_1742);
xor U1808 (N_1808,N_1624,N_1694);
nor U1809 (N_1809,N_1658,N_1654);
nand U1810 (N_1810,N_1600,N_1735);
nand U1811 (N_1811,N_970,N_1375);
and U1812 (N_1812,N_1724,N_205);
nor U1813 (N_1813,N_610,N_1456);
and U1814 (N_1814,N_1274,N_1648);
or U1815 (N_1815,N_1618,N_1709);
or U1816 (N_1816,N_1637,N_1620);
and U1817 (N_1817,N_1745,N_1668);
and U1818 (N_1818,N_1527,N_1450);
nand U1819 (N_1819,N_1152,N_997);
xor U1820 (N_1820,N_1387,N_1655);
and U1821 (N_1821,N_1496,N_1708);
and U1822 (N_1822,N_1629,N_1759);
nand U1823 (N_1823,N_1649,N_1702);
nor U1824 (N_1824,N_1660,N_868);
nor U1825 (N_1825,N_1616,N_1424);
nor U1826 (N_1826,N_740,N_1615);
nor U1827 (N_1827,N_1517,N_1610);
nor U1828 (N_1828,N_1529,N_1378);
and U1829 (N_1829,N_1674,N_1755);
and U1830 (N_1830,N_382,N_1623);
and U1831 (N_1831,N_1747,N_1217);
nor U1832 (N_1832,N_1720,N_1684);
and U1833 (N_1833,N_1687,N_1750);
nand U1834 (N_1834,N_1675,N_1332);
nand U1835 (N_1835,N_1492,N_747);
nor U1836 (N_1836,N_1604,N_1041);
nor U1837 (N_1837,N_1522,N_1685);
xor U1838 (N_1838,N_1746,N_1730);
nand U1839 (N_1839,N_1756,N_1744);
nor U1840 (N_1840,N_1642,N_1646);
or U1841 (N_1841,N_1666,N_1369);
nor U1842 (N_1842,N_1634,N_1717);
or U1843 (N_1843,N_1362,N_1198);
nor U1844 (N_1844,N_1686,N_1716);
xnor U1845 (N_1845,N_1738,N_1661);
xnor U1846 (N_1846,N_1612,N_1614);
nor U1847 (N_1847,N_1645,N_1701);
xnor U1848 (N_1848,N_1241,N_1657);
nor U1849 (N_1849,N_1712,N_1607);
nand U1850 (N_1850,N_1726,N_1753);
or U1851 (N_1851,N_1721,N_1551);
nor U1852 (N_1852,N_1718,N_1705);
nand U1853 (N_1853,N_1719,N_1743);
or U1854 (N_1854,N_1704,N_1723);
nand U1855 (N_1855,N_1632,N_1688);
and U1856 (N_1856,N_1729,N_1741);
xnor U1857 (N_1857,In_947,N_891);
nor U1858 (N_1858,N_1160,N_1318);
or U1859 (N_1859,N_690,N_1603);
nor U1860 (N_1860,N_1564,N_1304);
nand U1861 (N_1861,N_1336,N_1663);
nor U1862 (N_1862,N_1680,N_1206);
nand U1863 (N_1863,N_1697,N_1602);
and U1864 (N_1864,N_1695,N_1298);
and U1865 (N_1865,N_1633,N_1662);
xnor U1866 (N_1866,N_1630,N_1460);
or U1867 (N_1867,N_235,N_1625);
or U1868 (N_1868,N_813,N_1659);
and U1869 (N_1869,N_1748,N_1703);
nand U1870 (N_1870,In_67,In_116);
nor U1871 (N_1871,In_600,N_669);
nor U1872 (N_1872,N_1681,N_1690);
and U1873 (N_1873,N_1693,N_1679);
nand U1874 (N_1874,N_1677,In_1544);
nand U1875 (N_1875,N_1264,N_1737);
nor U1876 (N_1876,N_1698,N_1734);
nor U1877 (N_1877,N_431,N_1653);
nor U1878 (N_1878,N_1671,N_1605);
nor U1879 (N_1879,N_1165,N_1227);
or U1880 (N_1880,N_1631,N_1340);
or U1881 (N_1881,N_1298,N_1640);
nor U1882 (N_1882,N_1702,N_970);
xnor U1883 (N_1883,N_1632,N_891);
nor U1884 (N_1884,N_1605,In_631);
nand U1885 (N_1885,N_1690,N_1603);
nand U1886 (N_1886,N_1632,N_1744);
nand U1887 (N_1887,N_1694,N_1206);
nor U1888 (N_1888,N_1336,N_1492);
nand U1889 (N_1889,N_1460,N_1594);
nand U1890 (N_1890,N_1739,N_1437);
and U1891 (N_1891,In_1048,In_947);
nor U1892 (N_1892,N_1647,N_1264);
xor U1893 (N_1893,N_1198,N_1681);
nand U1894 (N_1894,N_1642,N_1740);
and U1895 (N_1895,N_1744,N_1623);
nand U1896 (N_1896,N_1711,N_1624);
and U1897 (N_1897,N_1694,N_1743);
xnor U1898 (N_1898,N_1492,N_1728);
xnor U1899 (N_1899,N_1756,N_1750);
nor U1900 (N_1900,N_690,N_1668);
nor U1901 (N_1901,N_1605,N_1492);
xnor U1902 (N_1902,N_1600,N_1694);
nor U1903 (N_1903,N_1491,In_1048);
nor U1904 (N_1904,N_1387,N_1643);
xnor U1905 (N_1905,N_1340,N_1660);
or U1906 (N_1906,N_1625,N_610);
and U1907 (N_1907,N_970,N_235);
xor U1908 (N_1908,N_1362,N_1646);
nand U1909 (N_1909,N_1651,N_1727);
nand U1910 (N_1910,N_1494,N_1732);
nor U1911 (N_1911,N_1264,N_1607);
or U1912 (N_1912,N_1684,N_1741);
or U1913 (N_1913,N_1704,N_1622);
and U1914 (N_1914,N_1307,N_970);
nand U1915 (N_1915,N_1749,N_1744);
nand U1916 (N_1916,In_600,N_431);
nor U1917 (N_1917,N_813,N_1756);
nand U1918 (N_1918,N_1684,N_431);
nand U1919 (N_1919,N_1755,N_1749);
nor U1920 (N_1920,N_1824,N_1802);
nor U1921 (N_1921,N_1883,N_1913);
nor U1922 (N_1922,N_1864,N_1823);
xor U1923 (N_1923,N_1881,N_1818);
and U1924 (N_1924,N_1820,N_1885);
nand U1925 (N_1925,N_1816,N_1768);
nand U1926 (N_1926,N_1787,N_1833);
or U1927 (N_1927,N_1830,N_1867);
xor U1928 (N_1928,N_1813,N_1915);
and U1929 (N_1929,N_1880,N_1775);
nor U1930 (N_1930,N_1786,N_1774);
nand U1931 (N_1931,N_1840,N_1907);
nor U1932 (N_1932,N_1773,N_1834);
nand U1933 (N_1933,N_1844,N_1839);
and U1934 (N_1934,N_1767,N_1917);
or U1935 (N_1935,N_1868,N_1850);
and U1936 (N_1936,N_1899,N_1836);
xnor U1937 (N_1937,N_1795,N_1919);
and U1938 (N_1938,N_1819,N_1766);
and U1939 (N_1939,N_1879,N_1845);
or U1940 (N_1940,N_1769,N_1807);
nor U1941 (N_1941,N_1841,N_1870);
xnor U1942 (N_1942,N_1854,N_1863);
nand U1943 (N_1943,N_1911,N_1831);
xor U1944 (N_1944,N_1842,N_1893);
nor U1945 (N_1945,N_1875,N_1914);
xor U1946 (N_1946,N_1886,N_1825);
xnor U1947 (N_1947,N_1829,N_1905);
xnor U1948 (N_1948,N_1916,N_1791);
or U1949 (N_1949,N_1910,N_1869);
nand U1950 (N_1950,N_1770,N_1865);
nor U1951 (N_1951,N_1908,N_1884);
nand U1952 (N_1952,N_1792,N_1835);
and U1953 (N_1953,N_1873,N_1801);
nand U1954 (N_1954,N_1760,N_1871);
nand U1955 (N_1955,N_1855,N_1860);
nor U1956 (N_1956,N_1809,N_1892);
or U1957 (N_1957,N_1778,N_1782);
nand U1958 (N_1958,N_1797,N_1896);
and U1959 (N_1959,N_1812,N_1846);
or U1960 (N_1960,N_1800,N_1765);
xor U1961 (N_1961,N_1779,N_1866);
or U1962 (N_1962,N_1811,N_1882);
or U1963 (N_1963,N_1815,N_1861);
nand U1964 (N_1964,N_1826,N_1771);
nor U1965 (N_1965,N_1889,N_1858);
and U1966 (N_1966,N_1817,N_1906);
nor U1967 (N_1967,N_1859,N_1888);
nor U1968 (N_1968,N_1777,N_1862);
nor U1969 (N_1969,N_1890,N_1763);
xnor U1970 (N_1970,N_1843,N_1799);
xor U1971 (N_1971,N_1847,N_1793);
nor U1972 (N_1972,N_1805,N_1803);
and U1973 (N_1973,N_1832,N_1918);
nor U1974 (N_1974,N_1851,N_1772);
and U1975 (N_1975,N_1810,N_1838);
nand U1976 (N_1976,N_1814,N_1877);
and U1977 (N_1977,N_1872,N_1776);
and U1978 (N_1978,N_1806,N_1887);
or U1979 (N_1979,N_1794,N_1900);
nor U1980 (N_1980,N_1895,N_1852);
xnor U1981 (N_1981,N_1764,N_1761);
nand U1982 (N_1982,N_1848,N_1878);
nand U1983 (N_1983,N_1856,N_1897);
and U1984 (N_1984,N_1784,N_1804);
or U1985 (N_1985,N_1898,N_1849);
nor U1986 (N_1986,N_1853,N_1874);
nor U1987 (N_1987,N_1891,N_1780);
nand U1988 (N_1988,N_1902,N_1821);
and U1989 (N_1989,N_1796,N_1837);
nor U1990 (N_1990,N_1904,N_1903);
xor U1991 (N_1991,N_1762,N_1828);
nor U1992 (N_1992,N_1808,N_1790);
or U1993 (N_1993,N_1876,N_1788);
xnor U1994 (N_1994,N_1785,N_1857);
or U1995 (N_1995,N_1798,N_1822);
or U1996 (N_1996,N_1909,N_1912);
and U1997 (N_1997,N_1827,N_1783);
and U1998 (N_1998,N_1894,N_1901);
xnor U1999 (N_1999,N_1781,N_1789);
nor U2000 (N_2000,N_1827,N_1774);
nor U2001 (N_2001,N_1860,N_1871);
nor U2002 (N_2002,N_1848,N_1771);
nor U2003 (N_2003,N_1899,N_1860);
and U2004 (N_2004,N_1842,N_1863);
or U2005 (N_2005,N_1890,N_1914);
nand U2006 (N_2006,N_1834,N_1899);
nand U2007 (N_2007,N_1913,N_1799);
or U2008 (N_2008,N_1798,N_1825);
and U2009 (N_2009,N_1771,N_1820);
or U2010 (N_2010,N_1818,N_1776);
or U2011 (N_2011,N_1763,N_1910);
and U2012 (N_2012,N_1892,N_1804);
and U2013 (N_2013,N_1806,N_1779);
xor U2014 (N_2014,N_1797,N_1774);
xnor U2015 (N_2015,N_1785,N_1866);
nor U2016 (N_2016,N_1776,N_1898);
xor U2017 (N_2017,N_1873,N_1915);
nor U2018 (N_2018,N_1802,N_1908);
and U2019 (N_2019,N_1915,N_1897);
nor U2020 (N_2020,N_1769,N_1764);
or U2021 (N_2021,N_1822,N_1909);
nand U2022 (N_2022,N_1761,N_1787);
nand U2023 (N_2023,N_1838,N_1863);
xnor U2024 (N_2024,N_1848,N_1810);
or U2025 (N_2025,N_1806,N_1886);
nand U2026 (N_2026,N_1817,N_1873);
and U2027 (N_2027,N_1864,N_1812);
or U2028 (N_2028,N_1791,N_1820);
and U2029 (N_2029,N_1829,N_1765);
or U2030 (N_2030,N_1813,N_1802);
or U2031 (N_2031,N_1791,N_1857);
nor U2032 (N_2032,N_1894,N_1907);
or U2033 (N_2033,N_1810,N_1912);
nor U2034 (N_2034,N_1893,N_1814);
nor U2035 (N_2035,N_1764,N_1869);
nand U2036 (N_2036,N_1911,N_1875);
nand U2037 (N_2037,N_1911,N_1836);
or U2038 (N_2038,N_1888,N_1895);
and U2039 (N_2039,N_1900,N_1879);
or U2040 (N_2040,N_1761,N_1774);
or U2041 (N_2041,N_1804,N_1868);
nor U2042 (N_2042,N_1760,N_1883);
nand U2043 (N_2043,N_1888,N_1812);
xnor U2044 (N_2044,N_1917,N_1779);
nand U2045 (N_2045,N_1838,N_1917);
and U2046 (N_2046,N_1760,N_1804);
or U2047 (N_2047,N_1792,N_1841);
and U2048 (N_2048,N_1916,N_1870);
xnor U2049 (N_2049,N_1889,N_1888);
and U2050 (N_2050,N_1878,N_1804);
nor U2051 (N_2051,N_1849,N_1811);
or U2052 (N_2052,N_1809,N_1854);
xor U2053 (N_2053,N_1852,N_1815);
nor U2054 (N_2054,N_1863,N_1866);
nand U2055 (N_2055,N_1761,N_1854);
nand U2056 (N_2056,N_1803,N_1882);
or U2057 (N_2057,N_1802,N_1887);
and U2058 (N_2058,N_1905,N_1915);
nand U2059 (N_2059,N_1889,N_1867);
xnor U2060 (N_2060,N_1916,N_1847);
or U2061 (N_2061,N_1803,N_1781);
or U2062 (N_2062,N_1858,N_1891);
xnor U2063 (N_2063,N_1887,N_1865);
nor U2064 (N_2064,N_1894,N_1804);
xnor U2065 (N_2065,N_1780,N_1909);
or U2066 (N_2066,N_1784,N_1822);
nor U2067 (N_2067,N_1888,N_1844);
nor U2068 (N_2068,N_1799,N_1857);
and U2069 (N_2069,N_1794,N_1852);
nor U2070 (N_2070,N_1912,N_1846);
nand U2071 (N_2071,N_1855,N_1900);
and U2072 (N_2072,N_1809,N_1826);
nor U2073 (N_2073,N_1881,N_1782);
or U2074 (N_2074,N_1773,N_1821);
or U2075 (N_2075,N_1777,N_1906);
or U2076 (N_2076,N_1819,N_1833);
or U2077 (N_2077,N_1843,N_1779);
and U2078 (N_2078,N_1801,N_1902);
or U2079 (N_2079,N_1827,N_1764);
or U2080 (N_2080,N_1990,N_2031);
xor U2081 (N_2081,N_2040,N_2061);
xor U2082 (N_2082,N_1975,N_1944);
xnor U2083 (N_2083,N_1934,N_1970);
and U2084 (N_2084,N_2052,N_2034);
xor U2085 (N_2085,N_2066,N_2046);
xor U2086 (N_2086,N_2069,N_1983);
nor U2087 (N_2087,N_1997,N_2053);
or U2088 (N_2088,N_2001,N_2016);
nor U2089 (N_2089,N_2070,N_1957);
and U2090 (N_2090,N_2048,N_2023);
nor U2091 (N_2091,N_2018,N_1929);
xor U2092 (N_2092,N_1933,N_2059);
nand U2093 (N_2093,N_2027,N_2067);
or U2094 (N_2094,N_2062,N_2024);
or U2095 (N_2095,N_1930,N_2006);
nand U2096 (N_2096,N_1999,N_1927);
or U2097 (N_2097,N_1939,N_2043);
and U2098 (N_2098,N_1937,N_2054);
nor U2099 (N_2099,N_1985,N_2038);
nand U2100 (N_2100,N_2065,N_2026);
and U2101 (N_2101,N_2058,N_1921);
xor U2102 (N_2102,N_2028,N_1981);
xnor U2103 (N_2103,N_1953,N_2019);
nor U2104 (N_2104,N_2007,N_1977);
nand U2105 (N_2105,N_1935,N_2063);
nor U2106 (N_2106,N_1967,N_2025);
nor U2107 (N_2107,N_1984,N_2057);
and U2108 (N_2108,N_1956,N_1980);
nor U2109 (N_2109,N_1923,N_1973);
xor U2110 (N_2110,N_2017,N_1966);
nor U2111 (N_2111,N_1976,N_2032);
or U2112 (N_2112,N_1926,N_1949);
or U2113 (N_2113,N_2030,N_2005);
nor U2114 (N_2114,N_1987,N_1961);
or U2115 (N_2115,N_2015,N_2073);
nor U2116 (N_2116,N_2004,N_2068);
xnor U2117 (N_2117,N_1940,N_1946);
xor U2118 (N_2118,N_2042,N_2047);
nor U2119 (N_2119,N_2009,N_1938);
and U2120 (N_2120,N_1947,N_1978);
or U2121 (N_2121,N_1942,N_1991);
nor U2122 (N_2122,N_1945,N_1959);
nand U2123 (N_2123,N_2037,N_1920);
nor U2124 (N_2124,N_1992,N_1964);
or U2125 (N_2125,N_2039,N_1941);
nand U2126 (N_2126,N_1952,N_1950);
and U2127 (N_2127,N_2033,N_2003);
nand U2128 (N_2128,N_1974,N_2050);
or U2129 (N_2129,N_2060,N_1969);
or U2130 (N_2130,N_2041,N_2008);
nand U2131 (N_2131,N_2002,N_2035);
nor U2132 (N_2132,N_1996,N_2075);
and U2133 (N_2133,N_2014,N_1963);
or U2134 (N_2134,N_2029,N_1943);
nor U2135 (N_2135,N_1951,N_1962);
xnor U2136 (N_2136,N_1993,N_1960);
nand U2137 (N_2137,N_1971,N_2044);
xnor U2138 (N_2138,N_2012,N_2056);
and U2139 (N_2139,N_1994,N_1965);
and U2140 (N_2140,N_2077,N_2072);
nand U2141 (N_2141,N_1986,N_1998);
xor U2142 (N_2142,N_2049,N_1932);
nand U2143 (N_2143,N_2071,N_1922);
and U2144 (N_2144,N_1968,N_2022);
or U2145 (N_2145,N_1948,N_2076);
or U2146 (N_2146,N_1982,N_2013);
xnor U2147 (N_2147,N_1954,N_2074);
and U2148 (N_2148,N_2045,N_2079);
or U2149 (N_2149,N_1995,N_2078);
and U2150 (N_2150,N_2010,N_1955);
xor U2151 (N_2151,N_2064,N_2021);
xnor U2152 (N_2152,N_1988,N_1928);
or U2153 (N_2153,N_2051,N_1924);
nor U2154 (N_2154,N_2000,N_2020);
and U2155 (N_2155,N_2055,N_2036);
and U2156 (N_2156,N_1936,N_1931);
nand U2157 (N_2157,N_1979,N_1972);
or U2158 (N_2158,N_1958,N_2011);
nor U2159 (N_2159,N_1925,N_1989);
xor U2160 (N_2160,N_1945,N_1952);
nand U2161 (N_2161,N_2063,N_1947);
and U2162 (N_2162,N_2072,N_2038);
nand U2163 (N_2163,N_2006,N_1992);
xor U2164 (N_2164,N_2019,N_2076);
and U2165 (N_2165,N_2045,N_1993);
nor U2166 (N_2166,N_1999,N_1921);
xnor U2167 (N_2167,N_1967,N_1942);
xor U2168 (N_2168,N_2009,N_1977);
nor U2169 (N_2169,N_1986,N_2015);
nor U2170 (N_2170,N_1963,N_1957);
and U2171 (N_2171,N_1985,N_2062);
or U2172 (N_2172,N_2038,N_1983);
xor U2173 (N_2173,N_2058,N_2007);
nor U2174 (N_2174,N_1996,N_2002);
and U2175 (N_2175,N_1993,N_1952);
xnor U2176 (N_2176,N_2039,N_2036);
nor U2177 (N_2177,N_1948,N_1961);
and U2178 (N_2178,N_1929,N_1997);
nor U2179 (N_2179,N_2079,N_2054);
nor U2180 (N_2180,N_2063,N_1974);
and U2181 (N_2181,N_2023,N_1993);
nand U2182 (N_2182,N_2076,N_1985);
nor U2183 (N_2183,N_1945,N_2027);
xnor U2184 (N_2184,N_2008,N_1983);
nor U2185 (N_2185,N_1942,N_1989);
or U2186 (N_2186,N_2072,N_1974);
or U2187 (N_2187,N_1936,N_1967);
nand U2188 (N_2188,N_1982,N_1929);
xor U2189 (N_2189,N_2046,N_2006);
xnor U2190 (N_2190,N_2029,N_1970);
and U2191 (N_2191,N_2006,N_1955);
or U2192 (N_2192,N_1972,N_2022);
and U2193 (N_2193,N_2036,N_1938);
nand U2194 (N_2194,N_1976,N_2046);
and U2195 (N_2195,N_2021,N_1980);
xnor U2196 (N_2196,N_2018,N_2030);
or U2197 (N_2197,N_2025,N_1984);
nor U2198 (N_2198,N_1976,N_2064);
or U2199 (N_2199,N_1972,N_2077);
nand U2200 (N_2200,N_2027,N_1946);
and U2201 (N_2201,N_1938,N_2050);
nor U2202 (N_2202,N_1929,N_1935);
xor U2203 (N_2203,N_1984,N_1937);
xor U2204 (N_2204,N_1958,N_1922);
and U2205 (N_2205,N_1953,N_2023);
nand U2206 (N_2206,N_2034,N_2029);
or U2207 (N_2207,N_1931,N_2038);
and U2208 (N_2208,N_1987,N_1927);
and U2209 (N_2209,N_2025,N_1962);
and U2210 (N_2210,N_1941,N_1950);
and U2211 (N_2211,N_1924,N_2007);
nand U2212 (N_2212,N_2017,N_1997);
nand U2213 (N_2213,N_1950,N_1969);
xor U2214 (N_2214,N_2059,N_1934);
and U2215 (N_2215,N_2010,N_2023);
xnor U2216 (N_2216,N_2041,N_1969);
nor U2217 (N_2217,N_1984,N_1998);
nand U2218 (N_2218,N_1923,N_2032);
nor U2219 (N_2219,N_2044,N_2042);
and U2220 (N_2220,N_1942,N_1925);
and U2221 (N_2221,N_1986,N_1984);
nand U2222 (N_2222,N_1958,N_2054);
or U2223 (N_2223,N_1979,N_2078);
and U2224 (N_2224,N_1961,N_2034);
and U2225 (N_2225,N_1979,N_1974);
and U2226 (N_2226,N_2019,N_1926);
nand U2227 (N_2227,N_1925,N_2041);
xnor U2228 (N_2228,N_2016,N_2002);
xor U2229 (N_2229,N_1974,N_2020);
and U2230 (N_2230,N_2060,N_1989);
or U2231 (N_2231,N_1926,N_1991);
or U2232 (N_2232,N_2025,N_1996);
xnor U2233 (N_2233,N_1975,N_2004);
xor U2234 (N_2234,N_1970,N_1993);
xnor U2235 (N_2235,N_2061,N_1951);
xnor U2236 (N_2236,N_2051,N_1948);
or U2237 (N_2237,N_2002,N_1944);
or U2238 (N_2238,N_1963,N_2005);
nor U2239 (N_2239,N_1982,N_2039);
nor U2240 (N_2240,N_2121,N_2091);
nand U2241 (N_2241,N_2131,N_2200);
nor U2242 (N_2242,N_2125,N_2210);
and U2243 (N_2243,N_2123,N_2198);
or U2244 (N_2244,N_2165,N_2211);
and U2245 (N_2245,N_2133,N_2103);
xnor U2246 (N_2246,N_2151,N_2176);
or U2247 (N_2247,N_2107,N_2181);
xnor U2248 (N_2248,N_2137,N_2188);
nor U2249 (N_2249,N_2114,N_2206);
nor U2250 (N_2250,N_2179,N_2116);
or U2251 (N_2251,N_2204,N_2191);
nand U2252 (N_2252,N_2122,N_2111);
xor U2253 (N_2253,N_2108,N_2147);
or U2254 (N_2254,N_2175,N_2096);
nor U2255 (N_2255,N_2239,N_2219);
and U2256 (N_2256,N_2174,N_2120);
nor U2257 (N_2257,N_2232,N_2119);
or U2258 (N_2258,N_2201,N_2190);
nand U2259 (N_2259,N_2212,N_2118);
or U2260 (N_2260,N_2127,N_2230);
xor U2261 (N_2261,N_2154,N_2148);
xnor U2262 (N_2262,N_2162,N_2187);
xor U2263 (N_2263,N_2109,N_2089);
nor U2264 (N_2264,N_2215,N_2139);
xor U2265 (N_2265,N_2104,N_2196);
or U2266 (N_2266,N_2203,N_2140);
xnor U2267 (N_2267,N_2226,N_2189);
or U2268 (N_2268,N_2161,N_2234);
nor U2269 (N_2269,N_2153,N_2087);
nor U2270 (N_2270,N_2115,N_2138);
nand U2271 (N_2271,N_2086,N_2145);
nor U2272 (N_2272,N_2134,N_2142);
or U2273 (N_2273,N_2225,N_2157);
nor U2274 (N_2274,N_2135,N_2218);
xor U2275 (N_2275,N_2170,N_2081);
nor U2276 (N_2276,N_2186,N_2128);
and U2277 (N_2277,N_2169,N_2163);
xor U2278 (N_2278,N_2183,N_2236);
or U2279 (N_2279,N_2084,N_2152);
or U2280 (N_2280,N_2237,N_2223);
xor U2281 (N_2281,N_2159,N_2083);
nand U2282 (N_2282,N_2199,N_2150);
or U2283 (N_2283,N_2105,N_2224);
nand U2284 (N_2284,N_2090,N_2117);
or U2285 (N_2285,N_2233,N_2177);
and U2286 (N_2286,N_2209,N_2197);
nor U2287 (N_2287,N_2229,N_2102);
nor U2288 (N_2288,N_2222,N_2182);
nand U2289 (N_2289,N_2172,N_2214);
nor U2290 (N_2290,N_2155,N_2143);
nand U2291 (N_2291,N_2195,N_2213);
nand U2292 (N_2292,N_2101,N_2235);
or U2293 (N_2293,N_2171,N_2132);
and U2294 (N_2294,N_2180,N_2100);
or U2295 (N_2295,N_2217,N_2106);
nand U2296 (N_2296,N_2146,N_2095);
and U2297 (N_2297,N_2110,N_2166);
xnor U2298 (N_2298,N_2136,N_2093);
nand U2299 (N_2299,N_2124,N_2092);
and U2300 (N_2300,N_2160,N_2094);
and U2301 (N_2301,N_2099,N_2220);
or U2302 (N_2302,N_2130,N_2194);
nor U2303 (N_2303,N_2098,N_2168);
or U2304 (N_2304,N_2088,N_2173);
or U2305 (N_2305,N_2193,N_2202);
or U2306 (N_2306,N_2156,N_2227);
and U2307 (N_2307,N_2192,N_2208);
xor U2308 (N_2308,N_2112,N_2228);
or U2309 (N_2309,N_2097,N_2126);
nand U2310 (N_2310,N_2149,N_2082);
xnor U2311 (N_2311,N_2238,N_2221);
nor U2312 (N_2312,N_2113,N_2164);
and U2313 (N_2313,N_2205,N_2178);
nand U2314 (N_2314,N_2216,N_2080);
xnor U2315 (N_2315,N_2141,N_2085);
nor U2316 (N_2316,N_2129,N_2144);
or U2317 (N_2317,N_2184,N_2167);
nand U2318 (N_2318,N_2207,N_2158);
and U2319 (N_2319,N_2231,N_2185);
nand U2320 (N_2320,N_2174,N_2115);
nor U2321 (N_2321,N_2104,N_2152);
and U2322 (N_2322,N_2189,N_2184);
or U2323 (N_2323,N_2085,N_2092);
xor U2324 (N_2324,N_2112,N_2100);
nand U2325 (N_2325,N_2189,N_2223);
nor U2326 (N_2326,N_2142,N_2148);
xnor U2327 (N_2327,N_2166,N_2100);
or U2328 (N_2328,N_2100,N_2164);
xor U2329 (N_2329,N_2133,N_2194);
and U2330 (N_2330,N_2182,N_2219);
nor U2331 (N_2331,N_2200,N_2110);
nand U2332 (N_2332,N_2209,N_2214);
nor U2333 (N_2333,N_2222,N_2180);
or U2334 (N_2334,N_2098,N_2085);
nand U2335 (N_2335,N_2239,N_2113);
xor U2336 (N_2336,N_2107,N_2171);
xnor U2337 (N_2337,N_2105,N_2099);
nand U2338 (N_2338,N_2219,N_2196);
nor U2339 (N_2339,N_2106,N_2211);
or U2340 (N_2340,N_2213,N_2238);
xnor U2341 (N_2341,N_2093,N_2224);
nor U2342 (N_2342,N_2108,N_2099);
nand U2343 (N_2343,N_2142,N_2234);
nand U2344 (N_2344,N_2137,N_2197);
nand U2345 (N_2345,N_2200,N_2132);
xnor U2346 (N_2346,N_2084,N_2226);
nor U2347 (N_2347,N_2126,N_2152);
nor U2348 (N_2348,N_2221,N_2174);
and U2349 (N_2349,N_2081,N_2108);
nand U2350 (N_2350,N_2222,N_2147);
or U2351 (N_2351,N_2168,N_2217);
nand U2352 (N_2352,N_2137,N_2157);
xnor U2353 (N_2353,N_2125,N_2155);
nand U2354 (N_2354,N_2161,N_2111);
nand U2355 (N_2355,N_2108,N_2111);
nor U2356 (N_2356,N_2086,N_2166);
nand U2357 (N_2357,N_2141,N_2228);
nor U2358 (N_2358,N_2138,N_2127);
and U2359 (N_2359,N_2142,N_2125);
or U2360 (N_2360,N_2140,N_2189);
and U2361 (N_2361,N_2138,N_2195);
and U2362 (N_2362,N_2088,N_2179);
or U2363 (N_2363,N_2179,N_2182);
xor U2364 (N_2364,N_2214,N_2143);
or U2365 (N_2365,N_2157,N_2220);
and U2366 (N_2366,N_2123,N_2227);
nor U2367 (N_2367,N_2216,N_2117);
or U2368 (N_2368,N_2122,N_2141);
nand U2369 (N_2369,N_2097,N_2145);
xnor U2370 (N_2370,N_2234,N_2184);
or U2371 (N_2371,N_2167,N_2192);
or U2372 (N_2372,N_2230,N_2103);
nand U2373 (N_2373,N_2231,N_2222);
and U2374 (N_2374,N_2159,N_2178);
xor U2375 (N_2375,N_2191,N_2111);
nand U2376 (N_2376,N_2163,N_2203);
nand U2377 (N_2377,N_2185,N_2167);
xnor U2378 (N_2378,N_2176,N_2132);
nor U2379 (N_2379,N_2180,N_2136);
nand U2380 (N_2380,N_2142,N_2131);
and U2381 (N_2381,N_2081,N_2188);
or U2382 (N_2382,N_2156,N_2090);
nor U2383 (N_2383,N_2180,N_2137);
and U2384 (N_2384,N_2191,N_2167);
nor U2385 (N_2385,N_2231,N_2195);
nand U2386 (N_2386,N_2136,N_2112);
and U2387 (N_2387,N_2208,N_2161);
or U2388 (N_2388,N_2189,N_2115);
or U2389 (N_2389,N_2209,N_2164);
xnor U2390 (N_2390,N_2189,N_2229);
xnor U2391 (N_2391,N_2089,N_2147);
and U2392 (N_2392,N_2114,N_2105);
or U2393 (N_2393,N_2136,N_2164);
or U2394 (N_2394,N_2212,N_2084);
xnor U2395 (N_2395,N_2168,N_2162);
or U2396 (N_2396,N_2146,N_2128);
nor U2397 (N_2397,N_2206,N_2156);
or U2398 (N_2398,N_2181,N_2088);
and U2399 (N_2399,N_2227,N_2206);
and U2400 (N_2400,N_2383,N_2284);
nand U2401 (N_2401,N_2260,N_2262);
xnor U2402 (N_2402,N_2372,N_2302);
and U2403 (N_2403,N_2333,N_2252);
nand U2404 (N_2404,N_2396,N_2381);
and U2405 (N_2405,N_2392,N_2265);
xor U2406 (N_2406,N_2391,N_2388);
and U2407 (N_2407,N_2353,N_2294);
nor U2408 (N_2408,N_2393,N_2242);
or U2409 (N_2409,N_2269,N_2290);
nand U2410 (N_2410,N_2378,N_2325);
or U2411 (N_2411,N_2253,N_2272);
nand U2412 (N_2412,N_2307,N_2267);
nor U2413 (N_2413,N_2332,N_2334);
nor U2414 (N_2414,N_2329,N_2330);
and U2415 (N_2415,N_2326,N_2288);
or U2416 (N_2416,N_2286,N_2247);
xnor U2417 (N_2417,N_2338,N_2349);
nor U2418 (N_2418,N_2335,N_2375);
xor U2419 (N_2419,N_2310,N_2348);
xor U2420 (N_2420,N_2379,N_2314);
nor U2421 (N_2421,N_2240,N_2343);
nor U2422 (N_2422,N_2271,N_2398);
or U2423 (N_2423,N_2305,N_2281);
nor U2424 (N_2424,N_2358,N_2374);
or U2425 (N_2425,N_2357,N_2280);
xnor U2426 (N_2426,N_2251,N_2386);
or U2427 (N_2427,N_2370,N_2278);
nor U2428 (N_2428,N_2352,N_2243);
or U2429 (N_2429,N_2359,N_2395);
nor U2430 (N_2430,N_2316,N_2368);
nand U2431 (N_2431,N_2331,N_2342);
and U2432 (N_2432,N_2394,N_2360);
xor U2433 (N_2433,N_2373,N_2364);
nor U2434 (N_2434,N_2328,N_2276);
or U2435 (N_2435,N_2308,N_2293);
nor U2436 (N_2436,N_2248,N_2345);
and U2437 (N_2437,N_2351,N_2277);
xor U2438 (N_2438,N_2241,N_2275);
nor U2439 (N_2439,N_2289,N_2303);
nand U2440 (N_2440,N_2313,N_2350);
or U2441 (N_2441,N_2245,N_2244);
or U2442 (N_2442,N_2363,N_2336);
xnor U2443 (N_2443,N_2377,N_2309);
nand U2444 (N_2444,N_2259,N_2361);
or U2445 (N_2445,N_2323,N_2312);
nor U2446 (N_2446,N_2274,N_2257);
xor U2447 (N_2447,N_2315,N_2321);
nor U2448 (N_2448,N_2306,N_2376);
nand U2449 (N_2449,N_2268,N_2322);
and U2450 (N_2450,N_2297,N_2355);
xnor U2451 (N_2451,N_2273,N_2371);
nand U2452 (N_2452,N_2385,N_2347);
or U2453 (N_2453,N_2339,N_2263);
and U2454 (N_2454,N_2258,N_2387);
nor U2455 (N_2455,N_2344,N_2365);
xnor U2456 (N_2456,N_2324,N_2296);
and U2457 (N_2457,N_2380,N_2255);
xnor U2458 (N_2458,N_2337,N_2399);
nor U2459 (N_2459,N_2369,N_2304);
nor U2460 (N_2460,N_2264,N_2254);
and U2461 (N_2461,N_2382,N_2319);
or U2462 (N_2462,N_2282,N_2346);
nor U2463 (N_2463,N_2299,N_2341);
and U2464 (N_2464,N_2354,N_2397);
or U2465 (N_2465,N_2261,N_2246);
nor U2466 (N_2466,N_2317,N_2249);
and U2467 (N_2467,N_2362,N_2266);
and U2468 (N_2468,N_2356,N_2295);
nor U2469 (N_2469,N_2292,N_2285);
nor U2470 (N_2470,N_2390,N_2287);
xnor U2471 (N_2471,N_2320,N_2340);
nor U2472 (N_2472,N_2327,N_2311);
or U2473 (N_2473,N_2366,N_2279);
xnor U2474 (N_2474,N_2389,N_2298);
nor U2475 (N_2475,N_2300,N_2301);
nand U2476 (N_2476,N_2291,N_2283);
and U2477 (N_2477,N_2384,N_2318);
and U2478 (N_2478,N_2367,N_2250);
and U2479 (N_2479,N_2256,N_2270);
and U2480 (N_2480,N_2377,N_2246);
or U2481 (N_2481,N_2247,N_2367);
nand U2482 (N_2482,N_2356,N_2334);
nand U2483 (N_2483,N_2349,N_2385);
or U2484 (N_2484,N_2298,N_2371);
xnor U2485 (N_2485,N_2327,N_2322);
or U2486 (N_2486,N_2243,N_2319);
xnor U2487 (N_2487,N_2360,N_2319);
and U2488 (N_2488,N_2344,N_2262);
nand U2489 (N_2489,N_2366,N_2301);
or U2490 (N_2490,N_2259,N_2356);
nand U2491 (N_2491,N_2348,N_2247);
nand U2492 (N_2492,N_2300,N_2306);
nor U2493 (N_2493,N_2252,N_2332);
xor U2494 (N_2494,N_2259,N_2322);
or U2495 (N_2495,N_2353,N_2398);
nand U2496 (N_2496,N_2265,N_2348);
nand U2497 (N_2497,N_2278,N_2275);
nor U2498 (N_2498,N_2332,N_2260);
xor U2499 (N_2499,N_2374,N_2308);
nand U2500 (N_2500,N_2375,N_2358);
xor U2501 (N_2501,N_2307,N_2274);
xnor U2502 (N_2502,N_2252,N_2284);
xor U2503 (N_2503,N_2261,N_2299);
or U2504 (N_2504,N_2305,N_2315);
xor U2505 (N_2505,N_2258,N_2290);
nand U2506 (N_2506,N_2366,N_2273);
and U2507 (N_2507,N_2291,N_2282);
and U2508 (N_2508,N_2306,N_2286);
nand U2509 (N_2509,N_2351,N_2388);
or U2510 (N_2510,N_2328,N_2356);
xor U2511 (N_2511,N_2309,N_2315);
nor U2512 (N_2512,N_2333,N_2394);
or U2513 (N_2513,N_2387,N_2247);
or U2514 (N_2514,N_2374,N_2380);
nand U2515 (N_2515,N_2377,N_2331);
xnor U2516 (N_2516,N_2305,N_2372);
or U2517 (N_2517,N_2277,N_2361);
or U2518 (N_2518,N_2345,N_2342);
or U2519 (N_2519,N_2312,N_2243);
or U2520 (N_2520,N_2391,N_2268);
or U2521 (N_2521,N_2286,N_2387);
and U2522 (N_2522,N_2338,N_2278);
nor U2523 (N_2523,N_2374,N_2346);
or U2524 (N_2524,N_2353,N_2241);
xor U2525 (N_2525,N_2369,N_2243);
nor U2526 (N_2526,N_2320,N_2334);
nand U2527 (N_2527,N_2263,N_2264);
and U2528 (N_2528,N_2288,N_2386);
or U2529 (N_2529,N_2244,N_2266);
and U2530 (N_2530,N_2308,N_2344);
or U2531 (N_2531,N_2360,N_2261);
xor U2532 (N_2532,N_2355,N_2365);
or U2533 (N_2533,N_2366,N_2346);
and U2534 (N_2534,N_2275,N_2320);
or U2535 (N_2535,N_2356,N_2297);
xor U2536 (N_2536,N_2332,N_2391);
or U2537 (N_2537,N_2247,N_2336);
and U2538 (N_2538,N_2323,N_2354);
nand U2539 (N_2539,N_2264,N_2317);
nand U2540 (N_2540,N_2369,N_2371);
xnor U2541 (N_2541,N_2387,N_2254);
and U2542 (N_2542,N_2341,N_2371);
and U2543 (N_2543,N_2279,N_2392);
nor U2544 (N_2544,N_2393,N_2353);
nor U2545 (N_2545,N_2323,N_2263);
or U2546 (N_2546,N_2385,N_2322);
xnor U2547 (N_2547,N_2284,N_2288);
nor U2548 (N_2548,N_2373,N_2247);
nor U2549 (N_2549,N_2321,N_2285);
nand U2550 (N_2550,N_2277,N_2344);
nand U2551 (N_2551,N_2293,N_2243);
nor U2552 (N_2552,N_2348,N_2306);
nand U2553 (N_2553,N_2373,N_2281);
nor U2554 (N_2554,N_2254,N_2289);
and U2555 (N_2555,N_2294,N_2323);
and U2556 (N_2556,N_2243,N_2328);
nor U2557 (N_2557,N_2378,N_2250);
nor U2558 (N_2558,N_2342,N_2259);
and U2559 (N_2559,N_2340,N_2375);
and U2560 (N_2560,N_2446,N_2420);
or U2561 (N_2561,N_2418,N_2531);
and U2562 (N_2562,N_2436,N_2445);
nand U2563 (N_2563,N_2526,N_2517);
nor U2564 (N_2564,N_2492,N_2475);
and U2565 (N_2565,N_2441,N_2455);
nor U2566 (N_2566,N_2542,N_2433);
xor U2567 (N_2567,N_2488,N_2449);
nor U2568 (N_2568,N_2452,N_2514);
nor U2569 (N_2569,N_2413,N_2419);
nand U2570 (N_2570,N_2508,N_2505);
and U2571 (N_2571,N_2440,N_2536);
nor U2572 (N_2572,N_2443,N_2484);
and U2573 (N_2573,N_2550,N_2528);
and U2574 (N_2574,N_2558,N_2406);
nor U2575 (N_2575,N_2540,N_2557);
nor U2576 (N_2576,N_2479,N_2468);
nor U2577 (N_2577,N_2471,N_2489);
or U2578 (N_2578,N_2523,N_2426);
nor U2579 (N_2579,N_2423,N_2491);
xor U2580 (N_2580,N_2482,N_2400);
or U2581 (N_2581,N_2466,N_2506);
or U2582 (N_2582,N_2431,N_2555);
nand U2583 (N_2583,N_2453,N_2444);
nand U2584 (N_2584,N_2502,N_2416);
nor U2585 (N_2585,N_2545,N_2473);
nand U2586 (N_2586,N_2450,N_2497);
xor U2587 (N_2587,N_2403,N_2490);
nor U2588 (N_2588,N_2537,N_2507);
nand U2589 (N_2589,N_2401,N_2456);
or U2590 (N_2590,N_2414,N_2481);
nand U2591 (N_2591,N_2430,N_2457);
nor U2592 (N_2592,N_2415,N_2549);
xor U2593 (N_2593,N_2524,N_2422);
or U2594 (N_2594,N_2434,N_2432);
and U2595 (N_2595,N_2404,N_2509);
xor U2596 (N_2596,N_2500,N_2516);
or U2597 (N_2597,N_2554,N_2503);
nand U2598 (N_2598,N_2474,N_2409);
xor U2599 (N_2599,N_2438,N_2464);
and U2600 (N_2600,N_2527,N_2559);
nand U2601 (N_2601,N_2530,N_2510);
nor U2602 (N_2602,N_2535,N_2412);
or U2603 (N_2603,N_2551,N_2487);
or U2604 (N_2604,N_2448,N_2513);
nand U2605 (N_2605,N_2469,N_2520);
nand U2606 (N_2606,N_2511,N_2427);
nor U2607 (N_2607,N_2548,N_2518);
and U2608 (N_2608,N_2429,N_2437);
nor U2609 (N_2609,N_2477,N_2470);
xnor U2610 (N_2610,N_2408,N_2435);
xor U2611 (N_2611,N_2533,N_2447);
xor U2612 (N_2612,N_2467,N_2465);
or U2613 (N_2613,N_2411,N_2499);
or U2614 (N_2614,N_2424,N_2439);
xnor U2615 (N_2615,N_2534,N_2483);
nor U2616 (N_2616,N_2543,N_2493);
and U2617 (N_2617,N_2539,N_2472);
or U2618 (N_2618,N_2486,N_2512);
nor U2619 (N_2619,N_2405,N_2451);
xor U2620 (N_2620,N_2547,N_2478);
xnor U2621 (N_2621,N_2515,N_2556);
or U2622 (N_2622,N_2407,N_2496);
nand U2623 (N_2623,N_2460,N_2529);
or U2624 (N_2624,N_2463,N_2521);
nand U2625 (N_2625,N_2425,N_2454);
nand U2626 (N_2626,N_2519,N_2421);
and U2627 (N_2627,N_2476,N_2546);
nand U2628 (N_2628,N_2501,N_2498);
nor U2629 (N_2629,N_2458,N_2417);
nor U2630 (N_2630,N_2538,N_2504);
xor U2631 (N_2631,N_2525,N_2480);
and U2632 (N_2632,N_2428,N_2553);
or U2633 (N_2633,N_2552,N_2402);
nand U2634 (N_2634,N_2494,N_2459);
or U2635 (N_2635,N_2541,N_2485);
nor U2636 (N_2636,N_2522,N_2410);
xnor U2637 (N_2637,N_2461,N_2532);
nand U2638 (N_2638,N_2495,N_2544);
nor U2639 (N_2639,N_2442,N_2462);
and U2640 (N_2640,N_2435,N_2501);
and U2641 (N_2641,N_2407,N_2559);
or U2642 (N_2642,N_2437,N_2521);
or U2643 (N_2643,N_2492,N_2467);
nor U2644 (N_2644,N_2448,N_2414);
and U2645 (N_2645,N_2527,N_2450);
and U2646 (N_2646,N_2419,N_2535);
and U2647 (N_2647,N_2455,N_2444);
nor U2648 (N_2648,N_2540,N_2543);
xnor U2649 (N_2649,N_2448,N_2502);
or U2650 (N_2650,N_2526,N_2510);
nor U2651 (N_2651,N_2551,N_2533);
nor U2652 (N_2652,N_2555,N_2520);
and U2653 (N_2653,N_2559,N_2443);
nor U2654 (N_2654,N_2549,N_2508);
or U2655 (N_2655,N_2407,N_2415);
xnor U2656 (N_2656,N_2431,N_2482);
and U2657 (N_2657,N_2521,N_2522);
or U2658 (N_2658,N_2458,N_2420);
and U2659 (N_2659,N_2420,N_2461);
nand U2660 (N_2660,N_2413,N_2554);
nand U2661 (N_2661,N_2403,N_2556);
or U2662 (N_2662,N_2551,N_2473);
or U2663 (N_2663,N_2546,N_2495);
nor U2664 (N_2664,N_2524,N_2501);
xor U2665 (N_2665,N_2487,N_2471);
and U2666 (N_2666,N_2428,N_2495);
nor U2667 (N_2667,N_2495,N_2475);
nor U2668 (N_2668,N_2496,N_2525);
nand U2669 (N_2669,N_2548,N_2524);
and U2670 (N_2670,N_2451,N_2536);
and U2671 (N_2671,N_2416,N_2455);
xnor U2672 (N_2672,N_2530,N_2421);
xor U2673 (N_2673,N_2418,N_2505);
nand U2674 (N_2674,N_2412,N_2496);
or U2675 (N_2675,N_2454,N_2416);
and U2676 (N_2676,N_2500,N_2458);
xor U2677 (N_2677,N_2518,N_2439);
nor U2678 (N_2678,N_2524,N_2462);
nand U2679 (N_2679,N_2525,N_2402);
xnor U2680 (N_2680,N_2494,N_2432);
and U2681 (N_2681,N_2494,N_2502);
or U2682 (N_2682,N_2545,N_2500);
nand U2683 (N_2683,N_2533,N_2539);
nand U2684 (N_2684,N_2400,N_2437);
nor U2685 (N_2685,N_2521,N_2442);
or U2686 (N_2686,N_2475,N_2510);
xnor U2687 (N_2687,N_2544,N_2486);
and U2688 (N_2688,N_2446,N_2508);
or U2689 (N_2689,N_2419,N_2550);
nand U2690 (N_2690,N_2550,N_2400);
nand U2691 (N_2691,N_2506,N_2454);
nand U2692 (N_2692,N_2417,N_2436);
nor U2693 (N_2693,N_2508,N_2439);
nand U2694 (N_2694,N_2419,N_2472);
xor U2695 (N_2695,N_2494,N_2544);
nand U2696 (N_2696,N_2558,N_2522);
or U2697 (N_2697,N_2450,N_2517);
nand U2698 (N_2698,N_2544,N_2452);
or U2699 (N_2699,N_2480,N_2473);
nand U2700 (N_2700,N_2548,N_2500);
nor U2701 (N_2701,N_2437,N_2469);
nand U2702 (N_2702,N_2510,N_2424);
nor U2703 (N_2703,N_2558,N_2489);
xor U2704 (N_2704,N_2538,N_2513);
or U2705 (N_2705,N_2455,N_2457);
or U2706 (N_2706,N_2486,N_2472);
nand U2707 (N_2707,N_2400,N_2412);
nor U2708 (N_2708,N_2449,N_2475);
and U2709 (N_2709,N_2553,N_2471);
nand U2710 (N_2710,N_2428,N_2419);
and U2711 (N_2711,N_2459,N_2524);
xor U2712 (N_2712,N_2405,N_2503);
nor U2713 (N_2713,N_2521,N_2500);
and U2714 (N_2714,N_2416,N_2531);
nand U2715 (N_2715,N_2509,N_2557);
or U2716 (N_2716,N_2550,N_2479);
or U2717 (N_2717,N_2556,N_2519);
nor U2718 (N_2718,N_2527,N_2541);
nor U2719 (N_2719,N_2413,N_2495);
or U2720 (N_2720,N_2653,N_2693);
nor U2721 (N_2721,N_2658,N_2627);
or U2722 (N_2722,N_2686,N_2625);
or U2723 (N_2723,N_2675,N_2567);
and U2724 (N_2724,N_2704,N_2645);
nand U2725 (N_2725,N_2681,N_2650);
nor U2726 (N_2726,N_2697,N_2565);
nand U2727 (N_2727,N_2641,N_2608);
or U2728 (N_2728,N_2576,N_2589);
and U2729 (N_2729,N_2707,N_2668);
nor U2730 (N_2730,N_2581,N_2626);
or U2731 (N_2731,N_2630,N_2598);
or U2732 (N_2732,N_2660,N_2709);
xnor U2733 (N_2733,N_2579,N_2659);
and U2734 (N_2734,N_2666,N_2604);
nand U2735 (N_2735,N_2618,N_2570);
and U2736 (N_2736,N_2599,N_2710);
nand U2737 (N_2737,N_2602,N_2701);
nand U2738 (N_2738,N_2663,N_2575);
or U2739 (N_2739,N_2657,N_2612);
nor U2740 (N_2740,N_2560,N_2635);
or U2741 (N_2741,N_2673,N_2572);
nand U2742 (N_2742,N_2574,N_2689);
xor U2743 (N_2743,N_2718,N_2646);
and U2744 (N_2744,N_2703,N_2655);
xor U2745 (N_2745,N_2682,N_2593);
nor U2746 (N_2746,N_2617,N_2652);
nand U2747 (N_2747,N_2628,N_2597);
nor U2748 (N_2748,N_2620,N_2606);
nor U2749 (N_2749,N_2702,N_2588);
xnor U2750 (N_2750,N_2586,N_2562);
xor U2751 (N_2751,N_2680,N_2590);
nand U2752 (N_2752,N_2568,N_2661);
nor U2753 (N_2753,N_2610,N_2648);
nor U2754 (N_2754,N_2632,N_2684);
or U2755 (N_2755,N_2561,N_2600);
xor U2756 (N_2756,N_2669,N_2705);
xnor U2757 (N_2757,N_2584,N_2609);
nor U2758 (N_2758,N_2714,N_2613);
or U2759 (N_2759,N_2654,N_2638);
xnor U2760 (N_2760,N_2671,N_2629);
nor U2761 (N_2761,N_2582,N_2687);
or U2762 (N_2762,N_2717,N_2670);
and U2763 (N_2763,N_2677,N_2715);
or U2764 (N_2764,N_2691,N_2601);
and U2765 (N_2765,N_2685,N_2595);
and U2766 (N_2766,N_2719,N_2636);
xnor U2767 (N_2767,N_2577,N_2651);
and U2768 (N_2768,N_2591,N_2622);
or U2769 (N_2769,N_2564,N_2679);
xor U2770 (N_2770,N_2640,N_2642);
nor U2771 (N_2771,N_2605,N_2633);
nor U2772 (N_2772,N_2649,N_2643);
and U2773 (N_2773,N_2573,N_2656);
xnor U2774 (N_2774,N_2637,N_2690);
nor U2775 (N_2775,N_2611,N_2592);
nor U2776 (N_2776,N_2634,N_2712);
xor U2777 (N_2777,N_2614,N_2580);
nand U2778 (N_2778,N_2624,N_2700);
nand U2779 (N_2779,N_2688,N_2583);
nand U2780 (N_2780,N_2683,N_2706);
and U2781 (N_2781,N_2694,N_2711);
or U2782 (N_2782,N_2665,N_2698);
nor U2783 (N_2783,N_2603,N_2667);
or U2784 (N_2784,N_2692,N_2585);
nor U2785 (N_2785,N_2674,N_2713);
nand U2786 (N_2786,N_2672,N_2594);
xnor U2787 (N_2787,N_2623,N_2596);
xnor U2788 (N_2788,N_2621,N_2619);
or U2789 (N_2789,N_2566,N_2569);
xor U2790 (N_2790,N_2639,N_2664);
nor U2791 (N_2791,N_2563,N_2615);
nor U2792 (N_2792,N_2587,N_2647);
or U2793 (N_2793,N_2716,N_2676);
nand U2794 (N_2794,N_2699,N_2696);
nor U2795 (N_2795,N_2578,N_2607);
xor U2796 (N_2796,N_2631,N_2662);
xnor U2797 (N_2797,N_2644,N_2695);
xor U2798 (N_2798,N_2616,N_2571);
xor U2799 (N_2799,N_2708,N_2678);
nand U2800 (N_2800,N_2636,N_2563);
xnor U2801 (N_2801,N_2653,N_2698);
nand U2802 (N_2802,N_2681,N_2672);
nor U2803 (N_2803,N_2698,N_2662);
xnor U2804 (N_2804,N_2681,N_2685);
xnor U2805 (N_2805,N_2658,N_2694);
or U2806 (N_2806,N_2661,N_2637);
nor U2807 (N_2807,N_2671,N_2596);
and U2808 (N_2808,N_2569,N_2585);
xor U2809 (N_2809,N_2644,N_2608);
nand U2810 (N_2810,N_2697,N_2593);
xor U2811 (N_2811,N_2599,N_2567);
and U2812 (N_2812,N_2565,N_2715);
or U2813 (N_2813,N_2690,N_2706);
nor U2814 (N_2814,N_2629,N_2588);
and U2815 (N_2815,N_2563,N_2682);
or U2816 (N_2816,N_2601,N_2647);
nor U2817 (N_2817,N_2589,N_2564);
xnor U2818 (N_2818,N_2676,N_2615);
and U2819 (N_2819,N_2603,N_2632);
nand U2820 (N_2820,N_2675,N_2647);
and U2821 (N_2821,N_2699,N_2571);
nor U2822 (N_2822,N_2602,N_2678);
nor U2823 (N_2823,N_2657,N_2689);
or U2824 (N_2824,N_2714,N_2651);
nor U2825 (N_2825,N_2624,N_2609);
and U2826 (N_2826,N_2711,N_2574);
nor U2827 (N_2827,N_2685,N_2653);
nor U2828 (N_2828,N_2645,N_2606);
nor U2829 (N_2829,N_2561,N_2618);
nor U2830 (N_2830,N_2656,N_2653);
nand U2831 (N_2831,N_2605,N_2604);
nand U2832 (N_2832,N_2678,N_2649);
or U2833 (N_2833,N_2653,N_2568);
nor U2834 (N_2834,N_2654,N_2575);
and U2835 (N_2835,N_2697,N_2699);
xnor U2836 (N_2836,N_2619,N_2593);
or U2837 (N_2837,N_2614,N_2662);
xnor U2838 (N_2838,N_2617,N_2692);
xor U2839 (N_2839,N_2662,N_2589);
nor U2840 (N_2840,N_2682,N_2609);
nor U2841 (N_2841,N_2680,N_2585);
or U2842 (N_2842,N_2564,N_2603);
or U2843 (N_2843,N_2605,N_2681);
or U2844 (N_2844,N_2689,N_2663);
xnor U2845 (N_2845,N_2564,N_2639);
nand U2846 (N_2846,N_2708,N_2636);
or U2847 (N_2847,N_2678,N_2632);
xnor U2848 (N_2848,N_2586,N_2648);
or U2849 (N_2849,N_2718,N_2661);
xnor U2850 (N_2850,N_2700,N_2714);
nor U2851 (N_2851,N_2666,N_2681);
and U2852 (N_2852,N_2694,N_2623);
nand U2853 (N_2853,N_2669,N_2662);
nor U2854 (N_2854,N_2715,N_2681);
nor U2855 (N_2855,N_2658,N_2718);
nor U2856 (N_2856,N_2583,N_2563);
nand U2857 (N_2857,N_2590,N_2681);
or U2858 (N_2858,N_2697,N_2712);
or U2859 (N_2859,N_2620,N_2590);
nor U2860 (N_2860,N_2632,N_2611);
xnor U2861 (N_2861,N_2656,N_2618);
nand U2862 (N_2862,N_2683,N_2678);
and U2863 (N_2863,N_2712,N_2645);
and U2864 (N_2864,N_2695,N_2645);
nand U2865 (N_2865,N_2699,N_2642);
xor U2866 (N_2866,N_2666,N_2643);
and U2867 (N_2867,N_2658,N_2665);
nor U2868 (N_2868,N_2595,N_2677);
and U2869 (N_2869,N_2611,N_2614);
nand U2870 (N_2870,N_2599,N_2660);
xnor U2871 (N_2871,N_2682,N_2615);
and U2872 (N_2872,N_2659,N_2698);
or U2873 (N_2873,N_2581,N_2591);
or U2874 (N_2874,N_2607,N_2633);
or U2875 (N_2875,N_2683,N_2589);
xnor U2876 (N_2876,N_2582,N_2684);
and U2877 (N_2877,N_2634,N_2715);
nand U2878 (N_2878,N_2712,N_2571);
nor U2879 (N_2879,N_2675,N_2584);
nor U2880 (N_2880,N_2767,N_2780);
xor U2881 (N_2881,N_2776,N_2870);
nor U2882 (N_2882,N_2762,N_2813);
xnor U2883 (N_2883,N_2790,N_2832);
and U2884 (N_2884,N_2841,N_2738);
or U2885 (N_2885,N_2743,N_2733);
and U2886 (N_2886,N_2773,N_2839);
xor U2887 (N_2887,N_2864,N_2861);
and U2888 (N_2888,N_2745,N_2791);
xor U2889 (N_2889,N_2850,N_2855);
nor U2890 (N_2890,N_2748,N_2807);
nand U2891 (N_2891,N_2825,N_2835);
xnor U2892 (N_2892,N_2805,N_2866);
nor U2893 (N_2893,N_2799,N_2763);
xnor U2894 (N_2894,N_2721,N_2869);
and U2895 (N_2895,N_2831,N_2749);
or U2896 (N_2896,N_2865,N_2808);
or U2897 (N_2897,N_2766,N_2844);
and U2898 (N_2898,N_2859,N_2729);
nor U2899 (N_2899,N_2801,N_2877);
nand U2900 (N_2900,N_2827,N_2744);
nor U2901 (N_2901,N_2875,N_2803);
or U2902 (N_2902,N_2772,N_2830);
nand U2903 (N_2903,N_2802,N_2826);
nor U2904 (N_2904,N_2828,N_2775);
and U2905 (N_2905,N_2795,N_2874);
or U2906 (N_2906,N_2821,N_2731);
nand U2907 (N_2907,N_2812,N_2754);
nor U2908 (N_2908,N_2750,N_2817);
nand U2909 (N_2909,N_2756,N_2739);
or U2910 (N_2910,N_2737,N_2787);
or U2911 (N_2911,N_2783,N_2811);
and U2912 (N_2912,N_2768,N_2771);
or U2913 (N_2913,N_2760,N_2796);
nand U2914 (N_2914,N_2806,N_2845);
or U2915 (N_2915,N_2793,N_2823);
nor U2916 (N_2916,N_2818,N_2868);
xnor U2917 (N_2917,N_2819,N_2778);
xor U2918 (N_2918,N_2863,N_2798);
nor U2919 (N_2919,N_2860,N_2769);
nand U2920 (N_2920,N_2879,N_2837);
or U2921 (N_2921,N_2727,N_2854);
and U2922 (N_2922,N_2797,N_2872);
xnor U2923 (N_2923,N_2765,N_2840);
and U2924 (N_2924,N_2757,N_2842);
or U2925 (N_2925,N_2770,N_2809);
xor U2926 (N_2926,N_2758,N_2788);
nand U2927 (N_2927,N_2848,N_2764);
and U2928 (N_2928,N_2820,N_2736);
nor U2929 (N_2929,N_2836,N_2720);
xnor U2930 (N_2930,N_2735,N_2810);
nor U2931 (N_2931,N_2752,N_2824);
nor U2932 (N_2932,N_2838,N_2878);
and U2933 (N_2933,N_2779,N_2833);
or U2934 (N_2934,N_2774,N_2834);
nor U2935 (N_2935,N_2728,N_2829);
and U2936 (N_2936,N_2723,N_2746);
xnor U2937 (N_2937,N_2784,N_2724);
and U2938 (N_2938,N_2730,N_2871);
nand U2939 (N_2939,N_2755,N_2816);
xnor U2940 (N_2940,N_2725,N_2876);
or U2941 (N_2941,N_2786,N_2777);
xor U2942 (N_2942,N_2815,N_2740);
or U2943 (N_2943,N_2753,N_2847);
xor U2944 (N_2944,N_2853,N_2782);
and U2945 (N_2945,N_2732,N_2792);
or U2946 (N_2946,N_2873,N_2862);
nand U2947 (N_2947,N_2751,N_2843);
nor U2948 (N_2948,N_2761,N_2800);
nor U2949 (N_2949,N_2867,N_2789);
nand U2950 (N_2950,N_2849,N_2804);
nand U2951 (N_2951,N_2759,N_2846);
xnor U2952 (N_2952,N_2794,N_2814);
and U2953 (N_2953,N_2734,N_2722);
xnor U2954 (N_2954,N_2856,N_2857);
nor U2955 (N_2955,N_2781,N_2726);
and U2956 (N_2956,N_2747,N_2742);
and U2957 (N_2957,N_2851,N_2852);
xor U2958 (N_2958,N_2785,N_2858);
nor U2959 (N_2959,N_2822,N_2741);
xor U2960 (N_2960,N_2775,N_2843);
and U2961 (N_2961,N_2779,N_2867);
and U2962 (N_2962,N_2790,N_2799);
and U2963 (N_2963,N_2725,N_2804);
or U2964 (N_2964,N_2747,N_2848);
or U2965 (N_2965,N_2868,N_2822);
nor U2966 (N_2966,N_2778,N_2821);
nor U2967 (N_2967,N_2763,N_2737);
nor U2968 (N_2968,N_2758,N_2808);
and U2969 (N_2969,N_2771,N_2832);
xor U2970 (N_2970,N_2775,N_2821);
nand U2971 (N_2971,N_2762,N_2792);
and U2972 (N_2972,N_2872,N_2742);
and U2973 (N_2973,N_2823,N_2808);
or U2974 (N_2974,N_2792,N_2786);
and U2975 (N_2975,N_2738,N_2765);
nand U2976 (N_2976,N_2773,N_2804);
nand U2977 (N_2977,N_2758,N_2827);
xor U2978 (N_2978,N_2785,N_2796);
nor U2979 (N_2979,N_2784,N_2849);
xnor U2980 (N_2980,N_2772,N_2751);
and U2981 (N_2981,N_2730,N_2856);
or U2982 (N_2982,N_2758,N_2733);
nand U2983 (N_2983,N_2737,N_2725);
nor U2984 (N_2984,N_2781,N_2758);
nor U2985 (N_2985,N_2818,N_2791);
or U2986 (N_2986,N_2737,N_2870);
xor U2987 (N_2987,N_2832,N_2838);
nor U2988 (N_2988,N_2777,N_2782);
and U2989 (N_2989,N_2826,N_2813);
nand U2990 (N_2990,N_2745,N_2764);
or U2991 (N_2991,N_2812,N_2823);
nand U2992 (N_2992,N_2740,N_2844);
nor U2993 (N_2993,N_2793,N_2778);
and U2994 (N_2994,N_2733,N_2807);
nand U2995 (N_2995,N_2742,N_2869);
nor U2996 (N_2996,N_2792,N_2816);
nor U2997 (N_2997,N_2770,N_2870);
and U2998 (N_2998,N_2832,N_2859);
and U2999 (N_2999,N_2798,N_2729);
nand U3000 (N_3000,N_2784,N_2830);
nand U3001 (N_3001,N_2761,N_2851);
and U3002 (N_3002,N_2768,N_2749);
xnor U3003 (N_3003,N_2796,N_2786);
nor U3004 (N_3004,N_2821,N_2736);
nor U3005 (N_3005,N_2744,N_2869);
xor U3006 (N_3006,N_2878,N_2744);
xnor U3007 (N_3007,N_2734,N_2855);
and U3008 (N_3008,N_2851,N_2850);
nand U3009 (N_3009,N_2877,N_2740);
nor U3010 (N_3010,N_2835,N_2829);
xor U3011 (N_3011,N_2814,N_2787);
nor U3012 (N_3012,N_2780,N_2873);
xor U3013 (N_3013,N_2853,N_2874);
nand U3014 (N_3014,N_2726,N_2735);
nand U3015 (N_3015,N_2791,N_2870);
or U3016 (N_3016,N_2788,N_2725);
xnor U3017 (N_3017,N_2780,N_2851);
xnor U3018 (N_3018,N_2748,N_2795);
or U3019 (N_3019,N_2872,N_2784);
or U3020 (N_3020,N_2776,N_2812);
and U3021 (N_3021,N_2803,N_2799);
or U3022 (N_3022,N_2789,N_2845);
nand U3023 (N_3023,N_2844,N_2806);
nor U3024 (N_3024,N_2726,N_2863);
and U3025 (N_3025,N_2818,N_2843);
and U3026 (N_3026,N_2725,N_2853);
nand U3027 (N_3027,N_2817,N_2768);
xor U3028 (N_3028,N_2874,N_2827);
or U3029 (N_3029,N_2788,N_2827);
or U3030 (N_3030,N_2821,N_2806);
xor U3031 (N_3031,N_2842,N_2796);
nor U3032 (N_3032,N_2844,N_2808);
or U3033 (N_3033,N_2778,N_2859);
nand U3034 (N_3034,N_2787,N_2723);
xor U3035 (N_3035,N_2829,N_2774);
or U3036 (N_3036,N_2825,N_2773);
xnor U3037 (N_3037,N_2871,N_2724);
nand U3038 (N_3038,N_2812,N_2766);
nor U3039 (N_3039,N_2829,N_2767);
xor U3040 (N_3040,N_2987,N_2976);
xor U3041 (N_3041,N_2959,N_3017);
nor U3042 (N_3042,N_2978,N_3010);
and U3043 (N_3043,N_2958,N_2890);
or U3044 (N_3044,N_2885,N_2968);
or U3045 (N_3045,N_2886,N_2927);
nor U3046 (N_3046,N_2883,N_2992);
nor U3047 (N_3047,N_3018,N_3002);
and U3048 (N_3048,N_2980,N_2881);
nand U3049 (N_3049,N_2906,N_2953);
nor U3050 (N_3050,N_3012,N_2975);
xor U3051 (N_3051,N_3024,N_2913);
nor U3052 (N_3052,N_2941,N_3025);
and U3053 (N_3053,N_2994,N_2974);
or U3054 (N_3054,N_2923,N_2920);
xnor U3055 (N_3055,N_2967,N_2981);
nor U3056 (N_3056,N_2943,N_2986);
and U3057 (N_3057,N_3006,N_3030);
xnor U3058 (N_3058,N_2948,N_2955);
nand U3059 (N_3059,N_2991,N_3021);
or U3060 (N_3060,N_2888,N_2973);
xor U3061 (N_3061,N_2971,N_3014);
nand U3062 (N_3062,N_3034,N_3011);
nor U3063 (N_3063,N_3009,N_2999);
xnor U3064 (N_3064,N_2960,N_3015);
and U3065 (N_3065,N_2893,N_3023);
or U3066 (N_3066,N_3004,N_2964);
and U3067 (N_3067,N_3000,N_2965);
or U3068 (N_3068,N_2910,N_3031);
xor U3069 (N_3069,N_2954,N_2952);
nand U3070 (N_3070,N_2882,N_3003);
and U3071 (N_3071,N_2908,N_2984);
and U3072 (N_3072,N_3013,N_2897);
nand U3073 (N_3073,N_2937,N_2901);
xnor U3074 (N_3074,N_3020,N_3027);
and U3075 (N_3075,N_3037,N_2915);
nand U3076 (N_3076,N_2951,N_2938);
nor U3077 (N_3077,N_2903,N_2990);
nand U3078 (N_3078,N_2928,N_2925);
nor U3079 (N_3079,N_3028,N_2949);
xor U3080 (N_3080,N_2892,N_2929);
nand U3081 (N_3081,N_3008,N_2956);
or U3082 (N_3082,N_3036,N_2887);
xor U3083 (N_3083,N_2997,N_2889);
nor U3084 (N_3084,N_2966,N_2962);
nor U3085 (N_3085,N_2919,N_2902);
xnor U3086 (N_3086,N_2904,N_3001);
or U3087 (N_3087,N_2899,N_2880);
nor U3088 (N_3088,N_2905,N_3035);
and U3089 (N_3089,N_3026,N_2946);
nand U3090 (N_3090,N_2894,N_2944);
nor U3091 (N_3091,N_3032,N_2970);
nand U3092 (N_3092,N_2891,N_2983);
nor U3093 (N_3093,N_2895,N_2940);
xnor U3094 (N_3094,N_2996,N_2985);
nand U3095 (N_3095,N_2898,N_2931);
and U3096 (N_3096,N_2926,N_2998);
nand U3097 (N_3097,N_2977,N_2969);
nor U3098 (N_3098,N_2921,N_2912);
xnor U3099 (N_3099,N_2972,N_3007);
or U3100 (N_3100,N_2922,N_3033);
or U3101 (N_3101,N_2933,N_2989);
nand U3102 (N_3102,N_2939,N_2957);
xor U3103 (N_3103,N_2914,N_2930);
xor U3104 (N_3104,N_2924,N_3005);
or U3105 (N_3105,N_2934,N_3039);
and U3106 (N_3106,N_2993,N_3022);
nand U3107 (N_3107,N_2982,N_2907);
and U3108 (N_3108,N_2884,N_2896);
xor U3109 (N_3109,N_2963,N_3038);
and U3110 (N_3110,N_2979,N_2950);
xnor U3111 (N_3111,N_2900,N_2945);
or U3112 (N_3112,N_2911,N_2995);
nor U3113 (N_3113,N_2935,N_3019);
or U3114 (N_3114,N_2961,N_3016);
nand U3115 (N_3115,N_2909,N_2947);
xnor U3116 (N_3116,N_2918,N_2917);
nor U3117 (N_3117,N_2942,N_2936);
xnor U3118 (N_3118,N_2988,N_3029);
and U3119 (N_3119,N_2916,N_2932);
and U3120 (N_3120,N_2966,N_2938);
or U3121 (N_3121,N_3025,N_2933);
nor U3122 (N_3122,N_3035,N_3018);
xnor U3123 (N_3123,N_3032,N_3005);
or U3124 (N_3124,N_2986,N_3002);
xor U3125 (N_3125,N_2935,N_2938);
nor U3126 (N_3126,N_2914,N_3018);
and U3127 (N_3127,N_2918,N_2884);
nor U3128 (N_3128,N_2888,N_2943);
and U3129 (N_3129,N_2946,N_2985);
or U3130 (N_3130,N_3023,N_3020);
xnor U3131 (N_3131,N_2952,N_3004);
xnor U3132 (N_3132,N_3032,N_3029);
xor U3133 (N_3133,N_2975,N_2946);
xor U3134 (N_3134,N_2952,N_2961);
xnor U3135 (N_3135,N_2919,N_2884);
or U3136 (N_3136,N_2962,N_2910);
xor U3137 (N_3137,N_2904,N_2910);
xnor U3138 (N_3138,N_2962,N_2915);
or U3139 (N_3139,N_2886,N_2929);
nor U3140 (N_3140,N_2988,N_3030);
nor U3141 (N_3141,N_2927,N_2983);
xnor U3142 (N_3142,N_2972,N_2913);
and U3143 (N_3143,N_2932,N_2943);
or U3144 (N_3144,N_2982,N_2903);
nand U3145 (N_3145,N_2949,N_3039);
xor U3146 (N_3146,N_3020,N_2881);
nor U3147 (N_3147,N_2889,N_3024);
nand U3148 (N_3148,N_2975,N_2889);
nand U3149 (N_3149,N_3010,N_2947);
nand U3150 (N_3150,N_3000,N_2982);
and U3151 (N_3151,N_2982,N_3023);
and U3152 (N_3152,N_2982,N_3009);
or U3153 (N_3153,N_2963,N_3010);
nand U3154 (N_3154,N_3002,N_2924);
nor U3155 (N_3155,N_2979,N_2963);
nor U3156 (N_3156,N_2943,N_2980);
or U3157 (N_3157,N_2923,N_2891);
and U3158 (N_3158,N_2881,N_2922);
and U3159 (N_3159,N_2938,N_2891);
xnor U3160 (N_3160,N_2884,N_2965);
or U3161 (N_3161,N_3003,N_3004);
nor U3162 (N_3162,N_2982,N_2979);
xor U3163 (N_3163,N_2957,N_2934);
nand U3164 (N_3164,N_2994,N_3004);
or U3165 (N_3165,N_2961,N_3032);
and U3166 (N_3166,N_3012,N_2896);
and U3167 (N_3167,N_2970,N_2905);
and U3168 (N_3168,N_2991,N_3035);
or U3169 (N_3169,N_2994,N_2950);
or U3170 (N_3170,N_2965,N_2955);
and U3171 (N_3171,N_2917,N_2937);
or U3172 (N_3172,N_2991,N_2949);
or U3173 (N_3173,N_3017,N_2901);
and U3174 (N_3174,N_3000,N_2981);
nor U3175 (N_3175,N_3009,N_2888);
nor U3176 (N_3176,N_2996,N_3019);
xor U3177 (N_3177,N_2945,N_2908);
nand U3178 (N_3178,N_3020,N_2953);
and U3179 (N_3179,N_2940,N_2969);
and U3180 (N_3180,N_2908,N_2934);
nand U3181 (N_3181,N_2896,N_2894);
and U3182 (N_3182,N_2883,N_2966);
or U3183 (N_3183,N_2999,N_2962);
xor U3184 (N_3184,N_2989,N_3026);
nor U3185 (N_3185,N_2955,N_2954);
or U3186 (N_3186,N_3024,N_2914);
and U3187 (N_3187,N_2898,N_3008);
nor U3188 (N_3188,N_2928,N_3011);
nor U3189 (N_3189,N_2906,N_2960);
and U3190 (N_3190,N_2913,N_2894);
nor U3191 (N_3191,N_2993,N_2914);
xor U3192 (N_3192,N_3038,N_2986);
nand U3193 (N_3193,N_3038,N_2983);
nand U3194 (N_3194,N_2942,N_2957);
or U3195 (N_3195,N_2978,N_2924);
or U3196 (N_3196,N_2943,N_2938);
or U3197 (N_3197,N_2912,N_2961);
nand U3198 (N_3198,N_3024,N_2911);
nand U3199 (N_3199,N_2903,N_2958);
nand U3200 (N_3200,N_3043,N_3052);
nor U3201 (N_3201,N_3061,N_3192);
nand U3202 (N_3202,N_3097,N_3110);
and U3203 (N_3203,N_3142,N_3096);
or U3204 (N_3204,N_3104,N_3041);
and U3205 (N_3205,N_3076,N_3123);
and U3206 (N_3206,N_3174,N_3119);
nand U3207 (N_3207,N_3048,N_3117);
or U3208 (N_3208,N_3160,N_3045);
or U3209 (N_3209,N_3060,N_3063);
nor U3210 (N_3210,N_3196,N_3157);
or U3211 (N_3211,N_3101,N_3171);
nand U3212 (N_3212,N_3079,N_3078);
nand U3213 (N_3213,N_3083,N_3177);
or U3214 (N_3214,N_3172,N_3159);
or U3215 (N_3215,N_3158,N_3155);
or U3216 (N_3216,N_3120,N_3134);
or U3217 (N_3217,N_3153,N_3087);
nor U3218 (N_3218,N_3173,N_3146);
xnor U3219 (N_3219,N_3054,N_3126);
nand U3220 (N_3220,N_3132,N_3133);
nand U3221 (N_3221,N_3175,N_3191);
or U3222 (N_3222,N_3184,N_3189);
and U3223 (N_3223,N_3190,N_3149);
or U3224 (N_3224,N_3199,N_3185);
nor U3225 (N_3225,N_3151,N_3113);
or U3226 (N_3226,N_3072,N_3129);
nor U3227 (N_3227,N_3050,N_3165);
or U3228 (N_3228,N_3108,N_3154);
nor U3229 (N_3229,N_3086,N_3057);
xor U3230 (N_3230,N_3118,N_3062);
nand U3231 (N_3231,N_3059,N_3122);
nor U3232 (N_3232,N_3127,N_3064);
and U3233 (N_3233,N_3055,N_3049);
xnor U3234 (N_3234,N_3091,N_3112);
xor U3235 (N_3235,N_3109,N_3114);
and U3236 (N_3236,N_3156,N_3116);
and U3237 (N_3237,N_3102,N_3082);
nor U3238 (N_3238,N_3182,N_3095);
and U3239 (N_3239,N_3161,N_3084);
or U3240 (N_3240,N_3197,N_3071);
xor U3241 (N_3241,N_3181,N_3106);
nand U3242 (N_3242,N_3089,N_3067);
nand U3243 (N_3243,N_3140,N_3170);
or U3244 (N_3244,N_3058,N_3105);
nand U3245 (N_3245,N_3125,N_3046);
and U3246 (N_3246,N_3141,N_3176);
nor U3247 (N_3247,N_3093,N_3088);
and U3248 (N_3248,N_3128,N_3152);
xnor U3249 (N_3249,N_3103,N_3187);
nor U3250 (N_3250,N_3195,N_3186);
nand U3251 (N_3251,N_3066,N_3092);
and U3252 (N_3252,N_3070,N_3051);
nand U3253 (N_3253,N_3139,N_3150);
nand U3254 (N_3254,N_3065,N_3131);
nand U3255 (N_3255,N_3193,N_3056);
and U3256 (N_3256,N_3098,N_3100);
nand U3257 (N_3257,N_3162,N_3166);
and U3258 (N_3258,N_3111,N_3068);
nand U3259 (N_3259,N_3040,N_3042);
xnor U3260 (N_3260,N_3130,N_3144);
nand U3261 (N_3261,N_3164,N_3047);
xor U3262 (N_3262,N_3169,N_3147);
xor U3263 (N_3263,N_3138,N_3053);
xnor U3264 (N_3264,N_3163,N_3167);
and U3265 (N_3265,N_3194,N_3080);
nor U3266 (N_3266,N_3115,N_3044);
nor U3267 (N_3267,N_3121,N_3188);
or U3268 (N_3268,N_3085,N_3107);
nand U3269 (N_3269,N_3135,N_3178);
nor U3270 (N_3270,N_3077,N_3168);
or U3271 (N_3271,N_3137,N_3075);
nand U3272 (N_3272,N_3099,N_3124);
and U3273 (N_3273,N_3198,N_3074);
nand U3274 (N_3274,N_3073,N_3143);
nand U3275 (N_3275,N_3094,N_3069);
xnor U3276 (N_3276,N_3081,N_3183);
nand U3277 (N_3277,N_3180,N_3136);
xor U3278 (N_3278,N_3179,N_3148);
nand U3279 (N_3279,N_3145,N_3090);
xnor U3280 (N_3280,N_3051,N_3073);
and U3281 (N_3281,N_3198,N_3135);
or U3282 (N_3282,N_3132,N_3175);
nand U3283 (N_3283,N_3109,N_3096);
nor U3284 (N_3284,N_3139,N_3156);
or U3285 (N_3285,N_3159,N_3071);
nand U3286 (N_3286,N_3085,N_3139);
nor U3287 (N_3287,N_3098,N_3085);
xor U3288 (N_3288,N_3125,N_3103);
nor U3289 (N_3289,N_3076,N_3193);
nand U3290 (N_3290,N_3167,N_3110);
or U3291 (N_3291,N_3170,N_3076);
xor U3292 (N_3292,N_3082,N_3115);
and U3293 (N_3293,N_3071,N_3162);
and U3294 (N_3294,N_3096,N_3084);
and U3295 (N_3295,N_3144,N_3122);
or U3296 (N_3296,N_3101,N_3160);
nor U3297 (N_3297,N_3111,N_3122);
xnor U3298 (N_3298,N_3052,N_3151);
nand U3299 (N_3299,N_3123,N_3090);
nor U3300 (N_3300,N_3114,N_3187);
xnor U3301 (N_3301,N_3161,N_3052);
or U3302 (N_3302,N_3131,N_3080);
nand U3303 (N_3303,N_3160,N_3163);
xor U3304 (N_3304,N_3110,N_3076);
and U3305 (N_3305,N_3110,N_3127);
nand U3306 (N_3306,N_3190,N_3082);
nor U3307 (N_3307,N_3183,N_3089);
nand U3308 (N_3308,N_3133,N_3189);
or U3309 (N_3309,N_3135,N_3197);
nor U3310 (N_3310,N_3073,N_3125);
or U3311 (N_3311,N_3076,N_3109);
or U3312 (N_3312,N_3129,N_3112);
nand U3313 (N_3313,N_3046,N_3175);
nor U3314 (N_3314,N_3071,N_3170);
nor U3315 (N_3315,N_3184,N_3074);
and U3316 (N_3316,N_3078,N_3118);
and U3317 (N_3317,N_3047,N_3163);
xnor U3318 (N_3318,N_3196,N_3068);
xor U3319 (N_3319,N_3113,N_3115);
nand U3320 (N_3320,N_3193,N_3068);
nand U3321 (N_3321,N_3176,N_3152);
nor U3322 (N_3322,N_3115,N_3070);
or U3323 (N_3323,N_3048,N_3120);
or U3324 (N_3324,N_3050,N_3049);
or U3325 (N_3325,N_3097,N_3178);
xor U3326 (N_3326,N_3197,N_3091);
nand U3327 (N_3327,N_3058,N_3190);
xor U3328 (N_3328,N_3062,N_3088);
nand U3329 (N_3329,N_3184,N_3151);
and U3330 (N_3330,N_3177,N_3072);
nand U3331 (N_3331,N_3101,N_3107);
xor U3332 (N_3332,N_3055,N_3137);
or U3333 (N_3333,N_3097,N_3088);
nor U3334 (N_3334,N_3130,N_3167);
xnor U3335 (N_3335,N_3164,N_3144);
nand U3336 (N_3336,N_3069,N_3042);
and U3337 (N_3337,N_3119,N_3167);
xor U3338 (N_3338,N_3131,N_3195);
nand U3339 (N_3339,N_3112,N_3087);
or U3340 (N_3340,N_3166,N_3068);
nand U3341 (N_3341,N_3054,N_3063);
and U3342 (N_3342,N_3131,N_3115);
and U3343 (N_3343,N_3160,N_3147);
or U3344 (N_3344,N_3067,N_3149);
nor U3345 (N_3345,N_3144,N_3156);
xor U3346 (N_3346,N_3174,N_3086);
nor U3347 (N_3347,N_3186,N_3111);
xor U3348 (N_3348,N_3065,N_3104);
nand U3349 (N_3349,N_3098,N_3079);
xor U3350 (N_3350,N_3091,N_3071);
nor U3351 (N_3351,N_3168,N_3199);
nor U3352 (N_3352,N_3188,N_3080);
nand U3353 (N_3353,N_3178,N_3105);
nor U3354 (N_3354,N_3126,N_3128);
or U3355 (N_3355,N_3164,N_3181);
and U3356 (N_3356,N_3079,N_3096);
nand U3357 (N_3357,N_3077,N_3199);
and U3358 (N_3358,N_3128,N_3072);
xnor U3359 (N_3359,N_3047,N_3121);
xor U3360 (N_3360,N_3213,N_3249);
xnor U3361 (N_3361,N_3292,N_3286);
and U3362 (N_3362,N_3350,N_3354);
nand U3363 (N_3363,N_3311,N_3340);
nand U3364 (N_3364,N_3332,N_3288);
nor U3365 (N_3365,N_3345,N_3283);
or U3366 (N_3366,N_3342,N_3268);
nor U3367 (N_3367,N_3298,N_3287);
nor U3368 (N_3368,N_3300,N_3281);
xor U3369 (N_3369,N_3293,N_3338);
nor U3370 (N_3370,N_3359,N_3230);
or U3371 (N_3371,N_3206,N_3226);
or U3372 (N_3372,N_3308,N_3262);
xnor U3373 (N_3373,N_3318,N_3344);
or U3374 (N_3374,N_3294,N_3279);
and U3375 (N_3375,N_3284,N_3355);
xnor U3376 (N_3376,N_3260,N_3301);
nand U3377 (N_3377,N_3222,N_3227);
or U3378 (N_3378,N_3304,N_3231);
and U3379 (N_3379,N_3312,N_3278);
and U3380 (N_3380,N_3316,N_3285);
and U3381 (N_3381,N_3330,N_3204);
and U3382 (N_3382,N_3233,N_3313);
or U3383 (N_3383,N_3236,N_3215);
or U3384 (N_3384,N_3218,N_3232);
xor U3385 (N_3385,N_3248,N_3256);
nand U3386 (N_3386,N_3282,N_3225);
and U3387 (N_3387,N_3269,N_3310);
nand U3388 (N_3388,N_3349,N_3351);
nand U3389 (N_3389,N_3235,N_3265);
and U3390 (N_3390,N_3295,N_3352);
nand U3391 (N_3391,N_3250,N_3242);
xnor U3392 (N_3392,N_3289,N_3254);
and U3393 (N_3393,N_3302,N_3228);
or U3394 (N_3394,N_3319,N_3234);
or U3395 (N_3395,N_3217,N_3221);
and U3396 (N_3396,N_3210,N_3327);
xnor U3397 (N_3397,N_3263,N_3322);
xnor U3398 (N_3398,N_3246,N_3291);
and U3399 (N_3399,N_3346,N_3325);
nand U3400 (N_3400,N_3307,N_3264);
and U3401 (N_3401,N_3219,N_3290);
nand U3402 (N_3402,N_3328,N_3238);
xnor U3403 (N_3403,N_3214,N_3241);
nand U3404 (N_3404,N_3200,N_3207);
xor U3405 (N_3405,N_3257,N_3297);
nor U3406 (N_3406,N_3333,N_3239);
xnor U3407 (N_3407,N_3209,N_3326);
nor U3408 (N_3408,N_3317,N_3202);
xnor U3409 (N_3409,N_3303,N_3271);
or U3410 (N_3410,N_3348,N_3323);
nand U3411 (N_3411,N_3357,N_3347);
nand U3412 (N_3412,N_3272,N_3331);
and U3413 (N_3413,N_3277,N_3314);
xnor U3414 (N_3414,N_3220,N_3324);
nor U3415 (N_3415,N_3212,N_3353);
nor U3416 (N_3416,N_3261,N_3216);
nor U3417 (N_3417,N_3243,N_3358);
xor U3418 (N_3418,N_3229,N_3356);
and U3419 (N_3419,N_3334,N_3320);
or U3420 (N_3420,N_3253,N_3224);
nand U3421 (N_3421,N_3255,N_3240);
or U3422 (N_3422,N_3296,N_3237);
or U3423 (N_3423,N_3335,N_3341);
xor U3424 (N_3424,N_3339,N_3306);
nand U3425 (N_3425,N_3252,N_3321);
nor U3426 (N_3426,N_3267,N_3247);
or U3427 (N_3427,N_3274,N_3251);
nor U3428 (N_3428,N_3336,N_3223);
nor U3429 (N_3429,N_3343,N_3315);
or U3430 (N_3430,N_3299,N_3337);
nor U3431 (N_3431,N_3266,N_3245);
nor U3432 (N_3432,N_3208,N_3305);
nand U3433 (N_3433,N_3203,N_3201);
or U3434 (N_3434,N_3205,N_3259);
xnor U3435 (N_3435,N_3329,N_3280);
or U3436 (N_3436,N_3258,N_3273);
and U3437 (N_3437,N_3270,N_3309);
or U3438 (N_3438,N_3211,N_3276);
or U3439 (N_3439,N_3244,N_3275);
or U3440 (N_3440,N_3295,N_3337);
xnor U3441 (N_3441,N_3221,N_3259);
xor U3442 (N_3442,N_3203,N_3351);
nor U3443 (N_3443,N_3310,N_3257);
or U3444 (N_3444,N_3269,N_3205);
nor U3445 (N_3445,N_3213,N_3254);
nor U3446 (N_3446,N_3206,N_3208);
xor U3447 (N_3447,N_3228,N_3211);
nor U3448 (N_3448,N_3218,N_3228);
and U3449 (N_3449,N_3248,N_3207);
nor U3450 (N_3450,N_3240,N_3258);
or U3451 (N_3451,N_3329,N_3352);
nor U3452 (N_3452,N_3308,N_3312);
nand U3453 (N_3453,N_3304,N_3303);
nor U3454 (N_3454,N_3279,N_3301);
and U3455 (N_3455,N_3306,N_3242);
xor U3456 (N_3456,N_3208,N_3337);
nand U3457 (N_3457,N_3222,N_3280);
or U3458 (N_3458,N_3353,N_3307);
nor U3459 (N_3459,N_3282,N_3276);
nor U3460 (N_3460,N_3333,N_3226);
nand U3461 (N_3461,N_3214,N_3352);
and U3462 (N_3462,N_3305,N_3264);
or U3463 (N_3463,N_3216,N_3308);
xor U3464 (N_3464,N_3284,N_3237);
and U3465 (N_3465,N_3243,N_3204);
xor U3466 (N_3466,N_3314,N_3281);
xnor U3467 (N_3467,N_3205,N_3321);
or U3468 (N_3468,N_3236,N_3334);
or U3469 (N_3469,N_3349,N_3314);
nor U3470 (N_3470,N_3341,N_3356);
nor U3471 (N_3471,N_3243,N_3279);
and U3472 (N_3472,N_3299,N_3314);
xnor U3473 (N_3473,N_3334,N_3288);
or U3474 (N_3474,N_3268,N_3309);
or U3475 (N_3475,N_3268,N_3308);
xor U3476 (N_3476,N_3285,N_3208);
xnor U3477 (N_3477,N_3222,N_3310);
or U3478 (N_3478,N_3336,N_3272);
nand U3479 (N_3479,N_3204,N_3314);
nand U3480 (N_3480,N_3331,N_3313);
nand U3481 (N_3481,N_3214,N_3273);
xnor U3482 (N_3482,N_3261,N_3310);
and U3483 (N_3483,N_3208,N_3306);
nand U3484 (N_3484,N_3202,N_3357);
nor U3485 (N_3485,N_3306,N_3300);
xor U3486 (N_3486,N_3252,N_3307);
or U3487 (N_3487,N_3341,N_3217);
nand U3488 (N_3488,N_3252,N_3211);
or U3489 (N_3489,N_3243,N_3242);
or U3490 (N_3490,N_3312,N_3319);
and U3491 (N_3491,N_3287,N_3345);
nand U3492 (N_3492,N_3224,N_3330);
nor U3493 (N_3493,N_3348,N_3246);
xor U3494 (N_3494,N_3226,N_3302);
nor U3495 (N_3495,N_3252,N_3216);
and U3496 (N_3496,N_3326,N_3285);
nand U3497 (N_3497,N_3250,N_3328);
and U3498 (N_3498,N_3341,N_3236);
and U3499 (N_3499,N_3295,N_3297);
xor U3500 (N_3500,N_3277,N_3284);
nor U3501 (N_3501,N_3279,N_3219);
or U3502 (N_3502,N_3299,N_3315);
xnor U3503 (N_3503,N_3246,N_3269);
xor U3504 (N_3504,N_3277,N_3224);
or U3505 (N_3505,N_3337,N_3233);
nor U3506 (N_3506,N_3294,N_3230);
nand U3507 (N_3507,N_3283,N_3349);
xnor U3508 (N_3508,N_3312,N_3287);
or U3509 (N_3509,N_3247,N_3225);
or U3510 (N_3510,N_3343,N_3303);
nor U3511 (N_3511,N_3255,N_3335);
xor U3512 (N_3512,N_3302,N_3325);
nor U3513 (N_3513,N_3333,N_3262);
and U3514 (N_3514,N_3356,N_3351);
nor U3515 (N_3515,N_3234,N_3215);
nor U3516 (N_3516,N_3207,N_3294);
nor U3517 (N_3517,N_3203,N_3321);
nor U3518 (N_3518,N_3254,N_3226);
xnor U3519 (N_3519,N_3309,N_3328);
and U3520 (N_3520,N_3455,N_3436);
and U3521 (N_3521,N_3423,N_3481);
xor U3522 (N_3522,N_3442,N_3371);
and U3523 (N_3523,N_3502,N_3463);
xnor U3524 (N_3524,N_3495,N_3387);
nand U3525 (N_3525,N_3470,N_3381);
or U3526 (N_3526,N_3438,N_3370);
xnor U3527 (N_3527,N_3459,N_3376);
and U3528 (N_3528,N_3511,N_3474);
and U3529 (N_3529,N_3514,N_3403);
nor U3530 (N_3530,N_3417,N_3448);
and U3531 (N_3531,N_3487,N_3504);
and U3532 (N_3532,N_3503,N_3453);
xor U3533 (N_3533,N_3496,N_3444);
xnor U3534 (N_3534,N_3475,N_3374);
nor U3535 (N_3535,N_3405,N_3422);
or U3536 (N_3536,N_3426,N_3458);
xor U3537 (N_3537,N_3489,N_3429);
nor U3538 (N_3538,N_3362,N_3388);
nand U3539 (N_3539,N_3435,N_3369);
xnor U3540 (N_3540,N_3394,N_3437);
nor U3541 (N_3541,N_3404,N_3415);
nand U3542 (N_3542,N_3501,N_3378);
or U3543 (N_3543,N_3457,N_3377);
or U3544 (N_3544,N_3434,N_3412);
or U3545 (N_3545,N_3446,N_3391);
nand U3546 (N_3546,N_3418,N_3397);
nand U3547 (N_3547,N_3367,N_3409);
or U3548 (N_3548,N_3414,N_3461);
or U3549 (N_3549,N_3408,N_3373);
nor U3550 (N_3550,N_3462,N_3445);
xnor U3551 (N_3551,N_3395,N_3472);
and U3552 (N_3552,N_3439,N_3433);
xor U3553 (N_3553,N_3513,N_3384);
nand U3554 (N_3554,N_3383,N_3450);
or U3555 (N_3555,N_3431,N_3485);
nor U3556 (N_3556,N_3407,N_3482);
xnor U3557 (N_3557,N_3401,N_3477);
nor U3558 (N_3558,N_3424,N_3443);
xor U3559 (N_3559,N_3515,N_3427);
and U3560 (N_3560,N_3406,N_3508);
nand U3561 (N_3561,N_3466,N_3430);
xor U3562 (N_3562,N_3484,N_3416);
or U3563 (N_3563,N_3483,N_3432);
xnor U3564 (N_3564,N_3493,N_3402);
nor U3565 (N_3565,N_3399,N_3421);
nor U3566 (N_3566,N_3413,N_3440);
nand U3567 (N_3567,N_3447,N_3497);
nand U3568 (N_3568,N_3396,N_3449);
xor U3569 (N_3569,N_3400,N_3390);
or U3570 (N_3570,N_3425,N_3389);
or U3571 (N_3571,N_3468,N_3491);
xor U3572 (N_3572,N_3519,N_3366);
xnor U3573 (N_3573,N_3509,N_3360);
xor U3574 (N_3574,N_3494,N_3398);
nor U3575 (N_3575,N_3363,N_3368);
or U3576 (N_3576,N_3490,N_3452);
and U3577 (N_3577,N_3465,N_3505);
nor U3578 (N_3578,N_3361,N_3488);
or U3579 (N_3579,N_3392,N_3467);
xnor U3580 (N_3580,N_3441,N_3498);
nand U3581 (N_3581,N_3428,N_3456);
or U3582 (N_3582,N_3454,N_3419);
or U3583 (N_3583,N_3385,N_3365);
or U3584 (N_3584,N_3375,N_3451);
nor U3585 (N_3585,N_3460,N_3379);
xnor U3586 (N_3586,N_3486,N_3411);
nor U3587 (N_3587,N_3506,N_3471);
xnor U3588 (N_3588,N_3517,N_3476);
nand U3589 (N_3589,N_3499,N_3393);
nand U3590 (N_3590,N_3507,N_3410);
or U3591 (N_3591,N_3469,N_3512);
nand U3592 (N_3592,N_3492,N_3420);
and U3593 (N_3593,N_3480,N_3518);
or U3594 (N_3594,N_3380,N_3516);
nand U3595 (N_3595,N_3500,N_3386);
nor U3596 (N_3596,N_3510,N_3372);
xnor U3597 (N_3597,N_3478,N_3382);
or U3598 (N_3598,N_3479,N_3464);
xor U3599 (N_3599,N_3473,N_3364);
or U3600 (N_3600,N_3426,N_3397);
xnor U3601 (N_3601,N_3414,N_3402);
nor U3602 (N_3602,N_3510,N_3435);
xnor U3603 (N_3603,N_3379,N_3361);
xor U3604 (N_3604,N_3504,N_3485);
nor U3605 (N_3605,N_3492,N_3432);
or U3606 (N_3606,N_3422,N_3377);
nor U3607 (N_3607,N_3383,N_3441);
and U3608 (N_3608,N_3391,N_3457);
nor U3609 (N_3609,N_3423,N_3499);
xnor U3610 (N_3610,N_3373,N_3512);
xnor U3611 (N_3611,N_3401,N_3499);
or U3612 (N_3612,N_3423,N_3414);
nand U3613 (N_3613,N_3517,N_3388);
or U3614 (N_3614,N_3482,N_3388);
nor U3615 (N_3615,N_3486,N_3467);
or U3616 (N_3616,N_3503,N_3460);
or U3617 (N_3617,N_3411,N_3507);
nand U3618 (N_3618,N_3436,N_3424);
and U3619 (N_3619,N_3488,N_3391);
nand U3620 (N_3620,N_3502,N_3414);
nand U3621 (N_3621,N_3403,N_3485);
and U3622 (N_3622,N_3493,N_3386);
or U3623 (N_3623,N_3445,N_3513);
or U3624 (N_3624,N_3483,N_3485);
or U3625 (N_3625,N_3496,N_3367);
and U3626 (N_3626,N_3519,N_3449);
nand U3627 (N_3627,N_3508,N_3408);
xor U3628 (N_3628,N_3479,N_3383);
nor U3629 (N_3629,N_3367,N_3416);
or U3630 (N_3630,N_3417,N_3503);
or U3631 (N_3631,N_3408,N_3459);
xnor U3632 (N_3632,N_3448,N_3453);
and U3633 (N_3633,N_3361,N_3446);
and U3634 (N_3634,N_3408,N_3489);
xnor U3635 (N_3635,N_3457,N_3378);
nor U3636 (N_3636,N_3426,N_3450);
nand U3637 (N_3637,N_3454,N_3519);
nand U3638 (N_3638,N_3474,N_3398);
or U3639 (N_3639,N_3376,N_3372);
xor U3640 (N_3640,N_3381,N_3426);
xor U3641 (N_3641,N_3434,N_3448);
nor U3642 (N_3642,N_3473,N_3449);
nand U3643 (N_3643,N_3473,N_3474);
nor U3644 (N_3644,N_3501,N_3371);
nor U3645 (N_3645,N_3396,N_3382);
nor U3646 (N_3646,N_3446,N_3449);
and U3647 (N_3647,N_3426,N_3500);
and U3648 (N_3648,N_3474,N_3419);
nand U3649 (N_3649,N_3504,N_3496);
and U3650 (N_3650,N_3445,N_3498);
or U3651 (N_3651,N_3504,N_3450);
nand U3652 (N_3652,N_3510,N_3364);
and U3653 (N_3653,N_3384,N_3493);
or U3654 (N_3654,N_3430,N_3496);
and U3655 (N_3655,N_3362,N_3399);
or U3656 (N_3656,N_3480,N_3404);
and U3657 (N_3657,N_3477,N_3372);
or U3658 (N_3658,N_3506,N_3403);
and U3659 (N_3659,N_3390,N_3391);
nand U3660 (N_3660,N_3478,N_3481);
nor U3661 (N_3661,N_3463,N_3481);
and U3662 (N_3662,N_3481,N_3453);
and U3663 (N_3663,N_3459,N_3466);
nor U3664 (N_3664,N_3478,N_3370);
and U3665 (N_3665,N_3517,N_3453);
nor U3666 (N_3666,N_3442,N_3398);
nand U3667 (N_3667,N_3373,N_3479);
xnor U3668 (N_3668,N_3393,N_3514);
xor U3669 (N_3669,N_3394,N_3450);
and U3670 (N_3670,N_3440,N_3439);
nor U3671 (N_3671,N_3497,N_3378);
or U3672 (N_3672,N_3386,N_3495);
xor U3673 (N_3673,N_3447,N_3445);
xnor U3674 (N_3674,N_3406,N_3476);
xnor U3675 (N_3675,N_3490,N_3460);
or U3676 (N_3676,N_3389,N_3506);
nor U3677 (N_3677,N_3478,N_3472);
nand U3678 (N_3678,N_3375,N_3364);
and U3679 (N_3679,N_3506,N_3510);
xor U3680 (N_3680,N_3675,N_3564);
nor U3681 (N_3681,N_3619,N_3523);
nand U3682 (N_3682,N_3594,N_3540);
xor U3683 (N_3683,N_3581,N_3657);
and U3684 (N_3684,N_3679,N_3575);
xor U3685 (N_3685,N_3546,N_3624);
xor U3686 (N_3686,N_3595,N_3625);
nor U3687 (N_3687,N_3570,N_3664);
nand U3688 (N_3688,N_3620,N_3653);
xor U3689 (N_3689,N_3605,N_3636);
xor U3690 (N_3690,N_3678,N_3650);
nor U3691 (N_3691,N_3545,N_3643);
xnor U3692 (N_3692,N_3649,N_3577);
nor U3693 (N_3693,N_3626,N_3542);
and U3694 (N_3694,N_3580,N_3654);
nand U3695 (N_3695,N_3662,N_3558);
and U3696 (N_3696,N_3640,N_3633);
nor U3697 (N_3697,N_3567,N_3586);
or U3698 (N_3698,N_3529,N_3589);
nand U3699 (N_3699,N_3539,N_3606);
nor U3700 (N_3700,N_3565,N_3556);
and U3701 (N_3701,N_3617,N_3566);
or U3702 (N_3702,N_3599,N_3602);
nand U3703 (N_3703,N_3631,N_3646);
and U3704 (N_3704,N_3637,N_3593);
and U3705 (N_3705,N_3521,N_3655);
and U3706 (N_3706,N_3562,N_3669);
and U3707 (N_3707,N_3568,N_3559);
nor U3708 (N_3708,N_3590,N_3663);
nor U3709 (N_3709,N_3533,N_3557);
nand U3710 (N_3710,N_3607,N_3608);
nor U3711 (N_3711,N_3642,N_3547);
nand U3712 (N_3712,N_3674,N_3527);
or U3713 (N_3713,N_3660,N_3612);
or U3714 (N_3714,N_3644,N_3591);
and U3715 (N_3715,N_3658,N_3613);
and U3716 (N_3716,N_3628,N_3596);
nor U3717 (N_3717,N_3544,N_3538);
and U3718 (N_3718,N_3615,N_3603);
and U3719 (N_3719,N_3647,N_3651);
nand U3720 (N_3720,N_3569,N_3610);
or U3721 (N_3721,N_3629,N_3616);
xor U3722 (N_3722,N_3531,N_3584);
nand U3723 (N_3723,N_3548,N_3532);
xor U3724 (N_3724,N_3661,N_3676);
nand U3725 (N_3725,N_3588,N_3551);
and U3726 (N_3726,N_3522,N_3534);
nor U3727 (N_3727,N_3555,N_3578);
nand U3728 (N_3728,N_3666,N_3587);
nand U3729 (N_3729,N_3535,N_3528);
xor U3730 (N_3730,N_3592,N_3579);
and U3731 (N_3731,N_3671,N_3673);
and U3732 (N_3732,N_3561,N_3672);
or U3733 (N_3733,N_3665,N_3656);
xnor U3734 (N_3734,N_3601,N_3550);
nand U3735 (N_3735,N_3621,N_3585);
xor U3736 (N_3736,N_3667,N_3635);
nand U3737 (N_3737,N_3623,N_3597);
or U3738 (N_3738,N_3630,N_3614);
and U3739 (N_3739,N_3572,N_3520);
or U3740 (N_3740,N_3560,N_3530);
and U3741 (N_3741,N_3639,N_3598);
and U3742 (N_3742,N_3638,N_3554);
nor U3743 (N_3743,N_3573,N_3677);
and U3744 (N_3744,N_3536,N_3549);
and U3745 (N_3745,N_3552,N_3553);
nand U3746 (N_3746,N_3604,N_3537);
nand U3747 (N_3747,N_3543,N_3582);
nand U3748 (N_3748,N_3622,N_3600);
nor U3749 (N_3749,N_3611,N_3648);
or U3750 (N_3750,N_3525,N_3632);
xnor U3751 (N_3751,N_3609,N_3563);
and U3752 (N_3752,N_3645,N_3524);
and U3753 (N_3753,N_3641,N_3576);
and U3754 (N_3754,N_3652,N_3541);
xor U3755 (N_3755,N_3574,N_3526);
xor U3756 (N_3756,N_3668,N_3627);
nor U3757 (N_3757,N_3634,N_3583);
and U3758 (N_3758,N_3659,N_3571);
or U3759 (N_3759,N_3670,N_3618);
nand U3760 (N_3760,N_3618,N_3559);
xor U3761 (N_3761,N_3586,N_3588);
and U3762 (N_3762,N_3569,N_3625);
and U3763 (N_3763,N_3657,N_3533);
nand U3764 (N_3764,N_3575,N_3547);
xor U3765 (N_3765,N_3614,N_3580);
xor U3766 (N_3766,N_3622,N_3560);
nand U3767 (N_3767,N_3602,N_3630);
and U3768 (N_3768,N_3679,N_3658);
nand U3769 (N_3769,N_3626,N_3532);
nor U3770 (N_3770,N_3654,N_3590);
and U3771 (N_3771,N_3539,N_3668);
nor U3772 (N_3772,N_3662,N_3590);
nor U3773 (N_3773,N_3660,N_3653);
and U3774 (N_3774,N_3622,N_3571);
and U3775 (N_3775,N_3634,N_3616);
nand U3776 (N_3776,N_3525,N_3612);
or U3777 (N_3777,N_3619,N_3611);
and U3778 (N_3778,N_3673,N_3570);
xnor U3779 (N_3779,N_3641,N_3535);
or U3780 (N_3780,N_3553,N_3610);
nand U3781 (N_3781,N_3543,N_3583);
and U3782 (N_3782,N_3660,N_3645);
nor U3783 (N_3783,N_3588,N_3560);
xnor U3784 (N_3784,N_3642,N_3628);
nor U3785 (N_3785,N_3544,N_3628);
nor U3786 (N_3786,N_3531,N_3636);
nor U3787 (N_3787,N_3564,N_3530);
nor U3788 (N_3788,N_3677,N_3597);
or U3789 (N_3789,N_3522,N_3651);
or U3790 (N_3790,N_3558,N_3581);
and U3791 (N_3791,N_3535,N_3569);
xor U3792 (N_3792,N_3578,N_3547);
and U3793 (N_3793,N_3520,N_3629);
nor U3794 (N_3794,N_3626,N_3599);
and U3795 (N_3795,N_3631,N_3570);
nor U3796 (N_3796,N_3660,N_3627);
and U3797 (N_3797,N_3619,N_3666);
xor U3798 (N_3798,N_3626,N_3628);
and U3799 (N_3799,N_3648,N_3526);
and U3800 (N_3800,N_3647,N_3535);
and U3801 (N_3801,N_3619,N_3556);
nand U3802 (N_3802,N_3560,N_3584);
nand U3803 (N_3803,N_3673,N_3552);
nor U3804 (N_3804,N_3527,N_3660);
or U3805 (N_3805,N_3640,N_3671);
xor U3806 (N_3806,N_3592,N_3611);
nand U3807 (N_3807,N_3607,N_3632);
nand U3808 (N_3808,N_3654,N_3624);
nor U3809 (N_3809,N_3610,N_3616);
or U3810 (N_3810,N_3578,N_3605);
or U3811 (N_3811,N_3640,N_3622);
nor U3812 (N_3812,N_3538,N_3528);
nor U3813 (N_3813,N_3538,N_3644);
xnor U3814 (N_3814,N_3582,N_3625);
nor U3815 (N_3815,N_3525,N_3628);
nand U3816 (N_3816,N_3597,N_3653);
and U3817 (N_3817,N_3524,N_3571);
xor U3818 (N_3818,N_3547,N_3678);
xor U3819 (N_3819,N_3641,N_3555);
or U3820 (N_3820,N_3619,N_3524);
xnor U3821 (N_3821,N_3672,N_3589);
nor U3822 (N_3822,N_3653,N_3640);
or U3823 (N_3823,N_3676,N_3654);
or U3824 (N_3824,N_3601,N_3543);
nor U3825 (N_3825,N_3640,N_3523);
or U3826 (N_3826,N_3654,N_3599);
nor U3827 (N_3827,N_3585,N_3654);
and U3828 (N_3828,N_3617,N_3669);
or U3829 (N_3829,N_3549,N_3666);
xor U3830 (N_3830,N_3531,N_3567);
nor U3831 (N_3831,N_3630,N_3588);
and U3832 (N_3832,N_3626,N_3563);
nor U3833 (N_3833,N_3601,N_3647);
or U3834 (N_3834,N_3676,N_3652);
nor U3835 (N_3835,N_3613,N_3602);
and U3836 (N_3836,N_3562,N_3549);
nand U3837 (N_3837,N_3520,N_3583);
xnor U3838 (N_3838,N_3596,N_3574);
and U3839 (N_3839,N_3619,N_3522);
nand U3840 (N_3840,N_3711,N_3774);
and U3841 (N_3841,N_3708,N_3757);
or U3842 (N_3842,N_3832,N_3831);
nor U3843 (N_3843,N_3691,N_3771);
nand U3844 (N_3844,N_3786,N_3761);
or U3845 (N_3845,N_3740,N_3836);
nand U3846 (N_3846,N_3826,N_3764);
nor U3847 (N_3847,N_3723,N_3687);
xnor U3848 (N_3848,N_3809,N_3713);
nand U3849 (N_3849,N_3770,N_3794);
or U3850 (N_3850,N_3818,N_3769);
and U3851 (N_3851,N_3763,N_3698);
xnor U3852 (N_3852,N_3760,N_3800);
nand U3853 (N_3853,N_3738,N_3783);
and U3854 (N_3854,N_3690,N_3829);
nor U3855 (N_3855,N_3696,N_3807);
nor U3856 (N_3856,N_3727,N_3775);
nor U3857 (N_3857,N_3735,N_3767);
and U3858 (N_3858,N_3754,N_3728);
or U3859 (N_3859,N_3741,N_3835);
xnor U3860 (N_3860,N_3838,N_3787);
xnor U3861 (N_3861,N_3824,N_3801);
nor U3862 (N_3862,N_3748,N_3689);
and U3863 (N_3863,N_3755,N_3699);
nor U3864 (N_3864,N_3780,N_3681);
xor U3865 (N_3865,N_3744,N_3789);
or U3866 (N_3866,N_3795,N_3680);
nand U3867 (N_3867,N_3804,N_3765);
xnor U3868 (N_3868,N_3730,N_3700);
and U3869 (N_3869,N_3709,N_3703);
and U3870 (N_3870,N_3803,N_3697);
or U3871 (N_3871,N_3686,N_3822);
xor U3872 (N_3872,N_3837,N_3782);
nor U3873 (N_3873,N_3793,N_3833);
nand U3874 (N_3874,N_3682,N_3693);
nand U3875 (N_3875,N_3802,N_3811);
nand U3876 (N_3876,N_3720,N_3776);
and U3877 (N_3877,N_3726,N_3798);
and U3878 (N_3878,N_3733,N_3839);
nand U3879 (N_3879,N_3692,N_3821);
xnor U3880 (N_3880,N_3815,N_3704);
or U3881 (N_3881,N_3830,N_3784);
nor U3882 (N_3882,N_3751,N_3695);
nor U3883 (N_3883,N_3791,N_3788);
and U3884 (N_3884,N_3820,N_3823);
nand U3885 (N_3885,N_3745,N_3756);
and U3886 (N_3886,N_3799,N_3819);
nand U3887 (N_3887,N_3828,N_3773);
and U3888 (N_3888,N_3772,N_3739);
or U3889 (N_3889,N_3694,N_3718);
and U3890 (N_3890,N_3777,N_3810);
or U3891 (N_3891,N_3707,N_3759);
and U3892 (N_3892,N_3701,N_3805);
nor U3893 (N_3893,N_3806,N_3719);
and U3894 (N_3894,N_3685,N_3779);
xor U3895 (N_3895,N_3796,N_3825);
nand U3896 (N_3896,N_3729,N_3714);
nand U3897 (N_3897,N_3731,N_3734);
xnor U3898 (N_3898,N_3753,N_3827);
nor U3899 (N_3899,N_3749,N_3814);
xnor U3900 (N_3900,N_3752,N_3746);
nor U3901 (N_3901,N_3768,N_3797);
nor U3902 (N_3902,N_3724,N_3712);
xnor U3903 (N_3903,N_3684,N_3816);
nand U3904 (N_3904,N_3781,N_3736);
and U3905 (N_3905,N_3722,N_3747);
nand U3906 (N_3906,N_3715,N_3725);
or U3907 (N_3907,N_3683,N_3785);
nand U3908 (N_3908,N_3742,N_3710);
or U3909 (N_3909,N_3766,N_3702);
nand U3910 (N_3910,N_3750,N_3808);
nor U3911 (N_3911,N_3792,N_3737);
or U3912 (N_3912,N_3813,N_3717);
nand U3913 (N_3913,N_3721,N_3706);
nand U3914 (N_3914,N_3778,N_3743);
or U3915 (N_3915,N_3817,N_3705);
nor U3916 (N_3916,N_3758,N_3834);
or U3917 (N_3917,N_3688,N_3790);
xor U3918 (N_3918,N_3762,N_3732);
or U3919 (N_3919,N_3812,N_3716);
xnor U3920 (N_3920,N_3692,N_3783);
xnor U3921 (N_3921,N_3769,N_3723);
or U3922 (N_3922,N_3685,N_3765);
nand U3923 (N_3923,N_3707,N_3789);
nand U3924 (N_3924,N_3745,N_3686);
and U3925 (N_3925,N_3815,N_3763);
xnor U3926 (N_3926,N_3734,N_3803);
or U3927 (N_3927,N_3708,N_3832);
and U3928 (N_3928,N_3723,N_3690);
nand U3929 (N_3929,N_3742,N_3732);
nor U3930 (N_3930,N_3774,N_3700);
xnor U3931 (N_3931,N_3836,N_3693);
and U3932 (N_3932,N_3709,N_3826);
or U3933 (N_3933,N_3681,N_3802);
nand U3934 (N_3934,N_3751,N_3709);
nand U3935 (N_3935,N_3721,N_3825);
nor U3936 (N_3936,N_3785,N_3717);
or U3937 (N_3937,N_3791,N_3822);
or U3938 (N_3938,N_3680,N_3731);
nor U3939 (N_3939,N_3783,N_3739);
nor U3940 (N_3940,N_3714,N_3696);
nand U3941 (N_3941,N_3802,N_3694);
nor U3942 (N_3942,N_3680,N_3736);
xnor U3943 (N_3943,N_3751,N_3804);
or U3944 (N_3944,N_3711,N_3821);
nor U3945 (N_3945,N_3786,N_3693);
and U3946 (N_3946,N_3806,N_3749);
or U3947 (N_3947,N_3735,N_3800);
nor U3948 (N_3948,N_3701,N_3692);
xnor U3949 (N_3949,N_3736,N_3759);
and U3950 (N_3950,N_3756,N_3691);
xnor U3951 (N_3951,N_3733,N_3794);
or U3952 (N_3952,N_3681,N_3694);
and U3953 (N_3953,N_3729,N_3777);
and U3954 (N_3954,N_3831,N_3692);
xnor U3955 (N_3955,N_3717,N_3698);
xnor U3956 (N_3956,N_3680,N_3740);
nor U3957 (N_3957,N_3784,N_3734);
xnor U3958 (N_3958,N_3751,N_3682);
xnor U3959 (N_3959,N_3809,N_3712);
and U3960 (N_3960,N_3832,N_3836);
nand U3961 (N_3961,N_3721,N_3798);
or U3962 (N_3962,N_3824,N_3760);
nand U3963 (N_3963,N_3837,N_3747);
and U3964 (N_3964,N_3681,N_3820);
xor U3965 (N_3965,N_3744,N_3769);
and U3966 (N_3966,N_3760,N_3778);
xor U3967 (N_3967,N_3807,N_3727);
and U3968 (N_3968,N_3683,N_3688);
xnor U3969 (N_3969,N_3720,N_3764);
xnor U3970 (N_3970,N_3808,N_3773);
or U3971 (N_3971,N_3745,N_3753);
and U3972 (N_3972,N_3819,N_3691);
xnor U3973 (N_3973,N_3801,N_3683);
nor U3974 (N_3974,N_3818,N_3771);
and U3975 (N_3975,N_3725,N_3772);
nor U3976 (N_3976,N_3811,N_3800);
xnor U3977 (N_3977,N_3692,N_3787);
or U3978 (N_3978,N_3680,N_3755);
nor U3979 (N_3979,N_3690,N_3737);
xnor U3980 (N_3980,N_3825,N_3681);
nor U3981 (N_3981,N_3728,N_3740);
or U3982 (N_3982,N_3785,N_3839);
and U3983 (N_3983,N_3716,N_3720);
xnor U3984 (N_3984,N_3750,N_3759);
xor U3985 (N_3985,N_3698,N_3758);
xnor U3986 (N_3986,N_3725,N_3684);
xor U3987 (N_3987,N_3828,N_3732);
or U3988 (N_3988,N_3814,N_3761);
nor U3989 (N_3989,N_3696,N_3694);
nand U3990 (N_3990,N_3753,N_3824);
or U3991 (N_3991,N_3720,N_3781);
nand U3992 (N_3992,N_3685,N_3700);
nand U3993 (N_3993,N_3725,N_3827);
nand U3994 (N_3994,N_3688,N_3823);
nor U3995 (N_3995,N_3834,N_3744);
nor U3996 (N_3996,N_3768,N_3765);
nand U3997 (N_3997,N_3835,N_3709);
and U3998 (N_3998,N_3827,N_3712);
and U3999 (N_3999,N_3798,N_3746);
nand U4000 (N_4000,N_3896,N_3988);
nand U4001 (N_4001,N_3977,N_3877);
nor U4002 (N_4002,N_3918,N_3887);
xnor U4003 (N_4003,N_3933,N_3912);
nand U4004 (N_4004,N_3966,N_3844);
xnor U4005 (N_4005,N_3930,N_3850);
and U4006 (N_4006,N_3953,N_3889);
nor U4007 (N_4007,N_3904,N_3847);
xnor U4008 (N_4008,N_3888,N_3867);
nand U4009 (N_4009,N_3922,N_3995);
xor U4010 (N_4010,N_3948,N_3964);
xor U4011 (N_4011,N_3932,N_3911);
nor U4012 (N_4012,N_3996,N_3979);
or U4013 (N_4013,N_3982,N_3949);
nor U4014 (N_4014,N_3917,N_3848);
nand U4015 (N_4015,N_3860,N_3872);
nor U4016 (N_4016,N_3855,N_3876);
nand U4017 (N_4017,N_3992,N_3921);
or U4018 (N_4018,N_3919,N_3871);
nor U4019 (N_4019,N_3882,N_3986);
and U4020 (N_4020,N_3874,N_3853);
or U4021 (N_4021,N_3936,N_3895);
xor U4022 (N_4022,N_3925,N_3903);
nand U4023 (N_4023,N_3974,N_3934);
xor U4024 (N_4024,N_3957,N_3913);
and U4025 (N_4025,N_3849,N_3898);
xnor U4026 (N_4026,N_3868,N_3969);
or U4027 (N_4027,N_3989,N_3907);
xnor U4028 (N_4028,N_3971,N_3875);
xnor U4029 (N_4029,N_3946,N_3983);
nand U4030 (N_4030,N_3962,N_3928);
nand U4031 (N_4031,N_3883,N_3924);
and U4032 (N_4032,N_3916,N_3885);
nand U4033 (N_4033,N_3905,N_3959);
and U4034 (N_4034,N_3991,N_3968);
or U4035 (N_4035,N_3920,N_3937);
and U4036 (N_4036,N_3929,N_3842);
nor U4037 (N_4037,N_3902,N_3908);
nand U4038 (N_4038,N_3857,N_3861);
or U4039 (N_4039,N_3951,N_3945);
nor U4040 (N_4040,N_3944,N_3854);
nor U4041 (N_4041,N_3859,N_3985);
and U4042 (N_4042,N_3863,N_3958);
nor U4043 (N_4043,N_3938,N_3845);
and U4044 (N_4044,N_3955,N_3880);
and U4045 (N_4045,N_3981,N_3942);
xnor U4046 (N_4046,N_3906,N_3993);
nand U4047 (N_4047,N_3960,N_3998);
xnor U4048 (N_4048,N_3900,N_3956);
or U4049 (N_4049,N_3973,N_3997);
nor U4050 (N_4050,N_3897,N_3892);
xnor U4051 (N_4051,N_3950,N_3910);
nor U4052 (N_4052,N_3965,N_3947);
xor U4053 (N_4053,N_3878,N_3967);
or U4054 (N_4054,N_3846,N_3869);
nand U4055 (N_4055,N_3940,N_3994);
or U4056 (N_4056,N_3923,N_3961);
xnor U4057 (N_4057,N_3901,N_3864);
nor U4058 (N_4058,N_3963,N_3884);
and U4059 (N_4059,N_3939,N_3870);
nand U4060 (N_4060,N_3999,N_3935);
nand U4061 (N_4061,N_3915,N_3990);
or U4062 (N_4062,N_3865,N_3899);
nor U4063 (N_4063,N_3927,N_3941);
nor U4064 (N_4064,N_3926,N_3909);
or U4065 (N_4065,N_3978,N_3952);
and U4066 (N_4066,N_3841,N_3891);
or U4067 (N_4067,N_3943,N_3975);
xnor U4068 (N_4068,N_3879,N_3972);
and U4069 (N_4069,N_3881,N_3873);
or U4070 (N_4070,N_3931,N_3976);
xnor U4071 (N_4071,N_3894,N_3970);
and U4072 (N_4072,N_3890,N_3858);
or U4073 (N_4073,N_3856,N_3886);
xor U4074 (N_4074,N_3914,N_3893);
or U4075 (N_4075,N_3862,N_3840);
nor U4076 (N_4076,N_3866,N_3980);
nor U4077 (N_4077,N_3843,N_3987);
or U4078 (N_4078,N_3852,N_3851);
or U4079 (N_4079,N_3954,N_3984);
or U4080 (N_4080,N_3930,N_3871);
xnor U4081 (N_4081,N_3912,N_3882);
and U4082 (N_4082,N_3905,N_3910);
and U4083 (N_4083,N_3917,N_3942);
or U4084 (N_4084,N_3961,N_3908);
and U4085 (N_4085,N_3889,N_3909);
and U4086 (N_4086,N_3969,N_3991);
nand U4087 (N_4087,N_3958,N_3853);
and U4088 (N_4088,N_3904,N_3949);
xor U4089 (N_4089,N_3882,N_3884);
nand U4090 (N_4090,N_3975,N_3916);
nand U4091 (N_4091,N_3987,N_3933);
xnor U4092 (N_4092,N_3866,N_3908);
nand U4093 (N_4093,N_3862,N_3863);
xnor U4094 (N_4094,N_3865,N_3999);
and U4095 (N_4095,N_3952,N_3935);
xor U4096 (N_4096,N_3878,N_3851);
and U4097 (N_4097,N_3895,N_3868);
and U4098 (N_4098,N_3891,N_3956);
xnor U4099 (N_4099,N_3990,N_3966);
nor U4100 (N_4100,N_3905,N_3947);
nor U4101 (N_4101,N_3961,N_3856);
nand U4102 (N_4102,N_3995,N_3914);
xor U4103 (N_4103,N_3934,N_3956);
nor U4104 (N_4104,N_3961,N_3863);
or U4105 (N_4105,N_3982,N_3963);
and U4106 (N_4106,N_3995,N_3886);
nor U4107 (N_4107,N_3897,N_3997);
nand U4108 (N_4108,N_3975,N_3995);
nor U4109 (N_4109,N_3949,N_3957);
xnor U4110 (N_4110,N_3841,N_3897);
xor U4111 (N_4111,N_3957,N_3872);
or U4112 (N_4112,N_3977,N_3864);
nand U4113 (N_4113,N_3972,N_3980);
nor U4114 (N_4114,N_3989,N_3885);
and U4115 (N_4115,N_3870,N_3880);
xor U4116 (N_4116,N_3905,N_3869);
nor U4117 (N_4117,N_3850,N_3886);
nand U4118 (N_4118,N_3973,N_3896);
nand U4119 (N_4119,N_3986,N_3971);
and U4120 (N_4120,N_3940,N_3950);
nor U4121 (N_4121,N_3858,N_3924);
or U4122 (N_4122,N_3957,N_3934);
nor U4123 (N_4123,N_3894,N_3854);
and U4124 (N_4124,N_3939,N_3898);
nor U4125 (N_4125,N_3921,N_3880);
nor U4126 (N_4126,N_3860,N_3971);
nand U4127 (N_4127,N_3866,N_3871);
xor U4128 (N_4128,N_3901,N_3897);
nor U4129 (N_4129,N_3872,N_3876);
nor U4130 (N_4130,N_3956,N_3847);
or U4131 (N_4131,N_3911,N_3874);
nand U4132 (N_4132,N_3965,N_3935);
nand U4133 (N_4133,N_3952,N_3912);
nand U4134 (N_4134,N_3991,N_3984);
or U4135 (N_4135,N_3972,N_3923);
or U4136 (N_4136,N_3971,N_3987);
nand U4137 (N_4137,N_3976,N_3898);
nor U4138 (N_4138,N_3921,N_3966);
nor U4139 (N_4139,N_3936,N_3996);
nor U4140 (N_4140,N_3937,N_3957);
nor U4141 (N_4141,N_3893,N_3904);
and U4142 (N_4142,N_3974,N_3907);
nand U4143 (N_4143,N_3992,N_3842);
nor U4144 (N_4144,N_3965,N_3889);
or U4145 (N_4145,N_3858,N_3983);
nor U4146 (N_4146,N_3906,N_3941);
nor U4147 (N_4147,N_3851,N_3990);
xnor U4148 (N_4148,N_3999,N_3947);
nor U4149 (N_4149,N_3840,N_3866);
or U4150 (N_4150,N_3852,N_3953);
or U4151 (N_4151,N_3893,N_3901);
or U4152 (N_4152,N_3880,N_3845);
nor U4153 (N_4153,N_3993,N_3900);
or U4154 (N_4154,N_3850,N_3959);
and U4155 (N_4155,N_3907,N_3998);
xor U4156 (N_4156,N_3985,N_3934);
nand U4157 (N_4157,N_3926,N_3957);
nand U4158 (N_4158,N_3968,N_3863);
or U4159 (N_4159,N_3989,N_3960);
and U4160 (N_4160,N_4126,N_4146);
xor U4161 (N_4161,N_4054,N_4028);
nand U4162 (N_4162,N_4102,N_4062);
nor U4163 (N_4163,N_4159,N_4038);
nor U4164 (N_4164,N_4033,N_4053);
nand U4165 (N_4165,N_4088,N_4070);
nor U4166 (N_4166,N_4069,N_4066);
xor U4167 (N_4167,N_4117,N_4111);
xnor U4168 (N_4168,N_4078,N_4089);
and U4169 (N_4169,N_4036,N_4009);
xor U4170 (N_4170,N_4112,N_4121);
nand U4171 (N_4171,N_4051,N_4076);
or U4172 (N_4172,N_4125,N_4080);
xor U4173 (N_4173,N_4086,N_4094);
and U4174 (N_4174,N_4074,N_4105);
and U4175 (N_4175,N_4158,N_4100);
xnor U4176 (N_4176,N_4030,N_4075);
or U4177 (N_4177,N_4073,N_4021);
and U4178 (N_4178,N_4000,N_4002);
nor U4179 (N_4179,N_4046,N_4031);
nor U4180 (N_4180,N_4063,N_4150);
and U4181 (N_4181,N_4026,N_4151);
nand U4182 (N_4182,N_4097,N_4143);
and U4183 (N_4183,N_4119,N_4090);
nand U4184 (N_4184,N_4006,N_4098);
nor U4185 (N_4185,N_4017,N_4005);
nor U4186 (N_4186,N_4141,N_4060);
and U4187 (N_4187,N_4101,N_4012);
xnor U4188 (N_4188,N_4118,N_4145);
and U4189 (N_4189,N_4108,N_4014);
xor U4190 (N_4190,N_4148,N_4127);
nand U4191 (N_4191,N_4055,N_4039);
and U4192 (N_4192,N_4131,N_4123);
nor U4193 (N_4193,N_4103,N_4156);
xnor U4194 (N_4194,N_4140,N_4040);
nand U4195 (N_4195,N_4029,N_4122);
or U4196 (N_4196,N_4025,N_4099);
or U4197 (N_4197,N_4023,N_4041);
nor U4198 (N_4198,N_4109,N_4013);
nor U4199 (N_4199,N_4047,N_4139);
xor U4200 (N_4200,N_4059,N_4136);
nor U4201 (N_4201,N_4106,N_4057);
or U4202 (N_4202,N_4149,N_4032);
or U4203 (N_4203,N_4085,N_4113);
or U4204 (N_4204,N_4095,N_4129);
nand U4205 (N_4205,N_4011,N_4044);
or U4206 (N_4206,N_4056,N_4152);
xnor U4207 (N_4207,N_4071,N_4043);
nor U4208 (N_4208,N_4091,N_4142);
and U4209 (N_4209,N_4010,N_4133);
xor U4210 (N_4210,N_4003,N_4134);
xor U4211 (N_4211,N_4157,N_4132);
and U4212 (N_4212,N_4058,N_4022);
nand U4213 (N_4213,N_4016,N_4037);
xnor U4214 (N_4214,N_4093,N_4135);
and U4215 (N_4215,N_4104,N_4116);
or U4216 (N_4216,N_4137,N_4082);
xnor U4217 (N_4217,N_4042,N_4096);
xor U4218 (N_4218,N_4092,N_4128);
or U4219 (N_4219,N_4154,N_4001);
xnor U4220 (N_4220,N_4087,N_4045);
nand U4221 (N_4221,N_4144,N_4077);
and U4222 (N_4222,N_4083,N_4027);
nor U4223 (N_4223,N_4138,N_4120);
nor U4224 (N_4224,N_4007,N_4079);
nor U4225 (N_4225,N_4020,N_4110);
or U4226 (N_4226,N_4067,N_4049);
and U4227 (N_4227,N_4068,N_4153);
or U4228 (N_4228,N_4065,N_4124);
or U4229 (N_4229,N_4081,N_4015);
nor U4230 (N_4230,N_4072,N_4018);
xnor U4231 (N_4231,N_4052,N_4114);
and U4232 (N_4232,N_4035,N_4155);
xor U4233 (N_4233,N_4084,N_4034);
or U4234 (N_4234,N_4024,N_4019);
nand U4235 (N_4235,N_4147,N_4004);
nor U4236 (N_4236,N_4048,N_4064);
nand U4237 (N_4237,N_4130,N_4115);
and U4238 (N_4238,N_4107,N_4050);
nand U4239 (N_4239,N_4008,N_4061);
nor U4240 (N_4240,N_4075,N_4067);
xor U4241 (N_4241,N_4156,N_4125);
nor U4242 (N_4242,N_4046,N_4157);
or U4243 (N_4243,N_4077,N_4039);
nand U4244 (N_4244,N_4012,N_4072);
and U4245 (N_4245,N_4072,N_4124);
nor U4246 (N_4246,N_4040,N_4119);
xor U4247 (N_4247,N_4000,N_4128);
nor U4248 (N_4248,N_4048,N_4156);
nand U4249 (N_4249,N_4142,N_4011);
nor U4250 (N_4250,N_4142,N_4144);
nor U4251 (N_4251,N_4008,N_4151);
or U4252 (N_4252,N_4005,N_4045);
and U4253 (N_4253,N_4095,N_4058);
nor U4254 (N_4254,N_4058,N_4044);
nor U4255 (N_4255,N_4098,N_4129);
or U4256 (N_4256,N_4034,N_4093);
and U4257 (N_4257,N_4028,N_4016);
and U4258 (N_4258,N_4033,N_4067);
nor U4259 (N_4259,N_4112,N_4051);
nand U4260 (N_4260,N_4149,N_4104);
and U4261 (N_4261,N_4060,N_4015);
and U4262 (N_4262,N_4115,N_4009);
and U4263 (N_4263,N_4048,N_4046);
nor U4264 (N_4264,N_4140,N_4132);
and U4265 (N_4265,N_4015,N_4086);
nor U4266 (N_4266,N_4140,N_4130);
or U4267 (N_4267,N_4154,N_4018);
xnor U4268 (N_4268,N_4105,N_4055);
xor U4269 (N_4269,N_4101,N_4051);
nand U4270 (N_4270,N_4093,N_4008);
and U4271 (N_4271,N_4098,N_4108);
or U4272 (N_4272,N_4065,N_4096);
nand U4273 (N_4273,N_4036,N_4099);
or U4274 (N_4274,N_4141,N_4020);
xnor U4275 (N_4275,N_4109,N_4125);
nor U4276 (N_4276,N_4078,N_4021);
or U4277 (N_4277,N_4077,N_4007);
nor U4278 (N_4278,N_4156,N_4158);
nor U4279 (N_4279,N_4088,N_4116);
nand U4280 (N_4280,N_4136,N_4126);
and U4281 (N_4281,N_4138,N_4129);
or U4282 (N_4282,N_4040,N_4009);
nor U4283 (N_4283,N_4120,N_4113);
or U4284 (N_4284,N_4048,N_4044);
nor U4285 (N_4285,N_4058,N_4126);
and U4286 (N_4286,N_4022,N_4030);
xor U4287 (N_4287,N_4101,N_4048);
nand U4288 (N_4288,N_4154,N_4087);
nand U4289 (N_4289,N_4142,N_4054);
xor U4290 (N_4290,N_4108,N_4021);
or U4291 (N_4291,N_4078,N_4054);
nor U4292 (N_4292,N_4082,N_4117);
nor U4293 (N_4293,N_4102,N_4047);
nand U4294 (N_4294,N_4151,N_4043);
xnor U4295 (N_4295,N_4040,N_4011);
and U4296 (N_4296,N_4102,N_4011);
nor U4297 (N_4297,N_4023,N_4038);
xnor U4298 (N_4298,N_4042,N_4083);
and U4299 (N_4299,N_4087,N_4077);
xor U4300 (N_4300,N_4056,N_4011);
and U4301 (N_4301,N_4066,N_4049);
and U4302 (N_4302,N_4095,N_4025);
or U4303 (N_4303,N_4056,N_4014);
or U4304 (N_4304,N_4136,N_4047);
nor U4305 (N_4305,N_4004,N_4084);
nor U4306 (N_4306,N_4109,N_4048);
xnor U4307 (N_4307,N_4044,N_4131);
nor U4308 (N_4308,N_4020,N_4099);
and U4309 (N_4309,N_4023,N_4057);
nor U4310 (N_4310,N_4095,N_4081);
and U4311 (N_4311,N_4076,N_4132);
xor U4312 (N_4312,N_4081,N_4048);
or U4313 (N_4313,N_4108,N_4092);
nor U4314 (N_4314,N_4002,N_4134);
nand U4315 (N_4315,N_4042,N_4052);
and U4316 (N_4316,N_4137,N_4042);
and U4317 (N_4317,N_4085,N_4119);
and U4318 (N_4318,N_4056,N_4087);
nand U4319 (N_4319,N_4024,N_4092);
and U4320 (N_4320,N_4305,N_4190);
and U4321 (N_4321,N_4270,N_4298);
nand U4322 (N_4322,N_4224,N_4276);
nor U4323 (N_4323,N_4191,N_4275);
nor U4324 (N_4324,N_4223,N_4206);
nand U4325 (N_4325,N_4236,N_4204);
or U4326 (N_4326,N_4216,N_4296);
xor U4327 (N_4327,N_4240,N_4233);
xnor U4328 (N_4328,N_4168,N_4264);
nor U4329 (N_4329,N_4211,N_4217);
nor U4330 (N_4330,N_4239,N_4311);
xnor U4331 (N_4331,N_4172,N_4234);
nor U4332 (N_4332,N_4303,N_4319);
nand U4333 (N_4333,N_4251,N_4220);
or U4334 (N_4334,N_4222,N_4284);
and U4335 (N_4335,N_4258,N_4260);
nand U4336 (N_4336,N_4199,N_4177);
nand U4337 (N_4337,N_4281,N_4231);
or U4338 (N_4338,N_4252,N_4287);
and U4339 (N_4339,N_4318,N_4310);
xnor U4340 (N_4340,N_4205,N_4278);
nor U4341 (N_4341,N_4259,N_4263);
and U4342 (N_4342,N_4225,N_4174);
and U4343 (N_4343,N_4295,N_4246);
or U4344 (N_4344,N_4307,N_4219);
nor U4345 (N_4345,N_4294,N_4221);
and U4346 (N_4346,N_4286,N_4309);
nand U4347 (N_4347,N_4277,N_4288);
or U4348 (N_4348,N_4245,N_4198);
and U4349 (N_4349,N_4274,N_4185);
nor U4350 (N_4350,N_4243,N_4247);
nand U4351 (N_4351,N_4300,N_4186);
xnor U4352 (N_4352,N_4313,N_4304);
nor U4353 (N_4353,N_4256,N_4267);
and U4354 (N_4354,N_4180,N_4210);
and U4355 (N_4355,N_4279,N_4207);
xor U4356 (N_4356,N_4200,N_4209);
and U4357 (N_4357,N_4178,N_4215);
nand U4358 (N_4358,N_4194,N_4192);
and U4359 (N_4359,N_4189,N_4306);
or U4360 (N_4360,N_4299,N_4235);
xnor U4361 (N_4361,N_4292,N_4165);
and U4362 (N_4362,N_4293,N_4268);
nor U4363 (N_4363,N_4179,N_4280);
nand U4364 (N_4364,N_4261,N_4203);
and U4365 (N_4365,N_4208,N_4271);
nor U4366 (N_4366,N_4257,N_4266);
xnor U4367 (N_4367,N_4202,N_4181);
or U4368 (N_4368,N_4188,N_4171);
nor U4369 (N_4369,N_4315,N_4197);
nor U4370 (N_4370,N_4232,N_4170);
xor U4371 (N_4371,N_4226,N_4176);
or U4372 (N_4372,N_4282,N_4249);
nand U4373 (N_4373,N_4227,N_4255);
nor U4374 (N_4374,N_4193,N_4218);
and U4375 (N_4375,N_4160,N_4228);
or U4376 (N_4376,N_4254,N_4290);
nor U4377 (N_4377,N_4162,N_4312);
xor U4378 (N_4378,N_4166,N_4201);
nor U4379 (N_4379,N_4184,N_4161);
or U4380 (N_4380,N_4182,N_4229);
xor U4381 (N_4381,N_4164,N_4212);
nor U4382 (N_4382,N_4248,N_4237);
or U4383 (N_4383,N_4272,N_4283);
nor U4384 (N_4384,N_4173,N_4183);
nor U4385 (N_4385,N_4169,N_4291);
nor U4386 (N_4386,N_4187,N_4297);
or U4387 (N_4387,N_4262,N_4285);
or U4388 (N_4388,N_4301,N_4195);
nand U4389 (N_4389,N_4241,N_4289);
nor U4390 (N_4390,N_4317,N_4269);
nor U4391 (N_4391,N_4314,N_4302);
and U4392 (N_4392,N_4244,N_4316);
nand U4393 (N_4393,N_4230,N_4265);
or U4394 (N_4394,N_4175,N_4238);
xor U4395 (N_4395,N_4213,N_4163);
nor U4396 (N_4396,N_4273,N_4253);
or U4397 (N_4397,N_4242,N_4196);
or U4398 (N_4398,N_4308,N_4214);
nor U4399 (N_4399,N_4250,N_4167);
or U4400 (N_4400,N_4183,N_4278);
or U4401 (N_4401,N_4298,N_4165);
and U4402 (N_4402,N_4173,N_4160);
or U4403 (N_4403,N_4200,N_4216);
or U4404 (N_4404,N_4235,N_4274);
nor U4405 (N_4405,N_4210,N_4255);
and U4406 (N_4406,N_4296,N_4276);
xor U4407 (N_4407,N_4187,N_4276);
xor U4408 (N_4408,N_4244,N_4268);
or U4409 (N_4409,N_4200,N_4240);
and U4410 (N_4410,N_4161,N_4219);
nor U4411 (N_4411,N_4239,N_4232);
nand U4412 (N_4412,N_4306,N_4261);
or U4413 (N_4413,N_4235,N_4308);
or U4414 (N_4414,N_4203,N_4182);
xnor U4415 (N_4415,N_4168,N_4279);
xor U4416 (N_4416,N_4211,N_4224);
or U4417 (N_4417,N_4171,N_4222);
or U4418 (N_4418,N_4260,N_4247);
nor U4419 (N_4419,N_4231,N_4209);
nand U4420 (N_4420,N_4183,N_4210);
xor U4421 (N_4421,N_4187,N_4286);
and U4422 (N_4422,N_4222,N_4179);
or U4423 (N_4423,N_4304,N_4241);
nand U4424 (N_4424,N_4245,N_4257);
or U4425 (N_4425,N_4266,N_4296);
nand U4426 (N_4426,N_4173,N_4293);
nand U4427 (N_4427,N_4184,N_4251);
and U4428 (N_4428,N_4256,N_4191);
and U4429 (N_4429,N_4250,N_4202);
and U4430 (N_4430,N_4241,N_4265);
nor U4431 (N_4431,N_4310,N_4164);
nor U4432 (N_4432,N_4303,N_4236);
or U4433 (N_4433,N_4183,N_4191);
nor U4434 (N_4434,N_4251,N_4160);
nor U4435 (N_4435,N_4211,N_4245);
or U4436 (N_4436,N_4238,N_4176);
or U4437 (N_4437,N_4177,N_4217);
and U4438 (N_4438,N_4318,N_4202);
nor U4439 (N_4439,N_4310,N_4194);
nand U4440 (N_4440,N_4163,N_4237);
nor U4441 (N_4441,N_4293,N_4299);
or U4442 (N_4442,N_4168,N_4258);
xor U4443 (N_4443,N_4309,N_4208);
nand U4444 (N_4444,N_4247,N_4286);
nor U4445 (N_4445,N_4242,N_4280);
and U4446 (N_4446,N_4311,N_4184);
nor U4447 (N_4447,N_4241,N_4282);
and U4448 (N_4448,N_4282,N_4257);
or U4449 (N_4449,N_4277,N_4235);
or U4450 (N_4450,N_4164,N_4264);
and U4451 (N_4451,N_4223,N_4205);
nor U4452 (N_4452,N_4297,N_4192);
nand U4453 (N_4453,N_4168,N_4187);
nand U4454 (N_4454,N_4180,N_4231);
and U4455 (N_4455,N_4239,N_4252);
and U4456 (N_4456,N_4163,N_4233);
nor U4457 (N_4457,N_4264,N_4217);
xnor U4458 (N_4458,N_4191,N_4260);
nor U4459 (N_4459,N_4304,N_4264);
and U4460 (N_4460,N_4178,N_4291);
or U4461 (N_4461,N_4290,N_4287);
and U4462 (N_4462,N_4173,N_4166);
and U4463 (N_4463,N_4245,N_4190);
nor U4464 (N_4464,N_4168,N_4161);
and U4465 (N_4465,N_4187,N_4315);
or U4466 (N_4466,N_4285,N_4162);
nor U4467 (N_4467,N_4309,N_4198);
nor U4468 (N_4468,N_4288,N_4217);
or U4469 (N_4469,N_4285,N_4277);
and U4470 (N_4470,N_4251,N_4237);
xnor U4471 (N_4471,N_4230,N_4173);
or U4472 (N_4472,N_4295,N_4313);
xor U4473 (N_4473,N_4175,N_4205);
and U4474 (N_4474,N_4239,N_4318);
nand U4475 (N_4475,N_4167,N_4203);
and U4476 (N_4476,N_4209,N_4287);
nor U4477 (N_4477,N_4316,N_4296);
and U4478 (N_4478,N_4211,N_4277);
and U4479 (N_4479,N_4202,N_4258);
and U4480 (N_4480,N_4415,N_4356);
or U4481 (N_4481,N_4339,N_4325);
and U4482 (N_4482,N_4400,N_4338);
or U4483 (N_4483,N_4471,N_4467);
xnor U4484 (N_4484,N_4479,N_4378);
nor U4485 (N_4485,N_4324,N_4438);
nand U4486 (N_4486,N_4430,N_4348);
nand U4487 (N_4487,N_4459,N_4367);
xnor U4488 (N_4488,N_4421,N_4409);
nor U4489 (N_4489,N_4401,N_4387);
xor U4490 (N_4490,N_4350,N_4450);
and U4491 (N_4491,N_4455,N_4425);
nor U4492 (N_4492,N_4377,N_4392);
or U4493 (N_4493,N_4379,N_4423);
nor U4494 (N_4494,N_4451,N_4382);
nor U4495 (N_4495,N_4363,N_4362);
xnor U4496 (N_4496,N_4464,N_4352);
and U4497 (N_4497,N_4396,N_4447);
xor U4498 (N_4498,N_4446,N_4449);
xor U4499 (N_4499,N_4322,N_4354);
nand U4500 (N_4500,N_4341,N_4422);
nand U4501 (N_4501,N_4452,N_4351);
or U4502 (N_4502,N_4399,N_4327);
xor U4503 (N_4503,N_4374,N_4478);
nand U4504 (N_4504,N_4461,N_4357);
nand U4505 (N_4505,N_4458,N_4375);
xnor U4506 (N_4506,N_4381,N_4419);
and U4507 (N_4507,N_4465,N_4373);
nor U4508 (N_4508,N_4433,N_4372);
nand U4509 (N_4509,N_4466,N_4359);
and U4510 (N_4510,N_4389,N_4426);
xor U4511 (N_4511,N_4329,N_4427);
nor U4512 (N_4512,N_4408,N_4347);
and U4513 (N_4513,N_4411,N_4448);
and U4514 (N_4514,N_4476,N_4349);
nor U4515 (N_4515,N_4393,N_4380);
and U4516 (N_4516,N_4368,N_4388);
and U4517 (N_4517,N_4353,N_4462);
nand U4518 (N_4518,N_4385,N_4410);
nand U4519 (N_4519,N_4335,N_4343);
or U4520 (N_4520,N_4457,N_4355);
nand U4521 (N_4521,N_4337,N_4405);
and U4522 (N_4522,N_4397,N_4431);
nor U4523 (N_4523,N_4412,N_4414);
nand U4524 (N_4524,N_4436,N_4416);
or U4525 (N_4525,N_4386,N_4320);
nor U4526 (N_4526,N_4360,N_4332);
or U4527 (N_4527,N_4463,N_4366);
or U4528 (N_4528,N_4346,N_4358);
xor U4529 (N_4529,N_4326,N_4376);
nor U4530 (N_4530,N_4417,N_4453);
xor U4531 (N_4531,N_4334,N_4323);
xor U4532 (N_4532,N_4328,N_4435);
nand U4533 (N_4533,N_4444,N_4404);
xor U4534 (N_4534,N_4418,N_4406);
xor U4535 (N_4535,N_4434,N_4402);
or U4536 (N_4536,N_4333,N_4395);
or U4537 (N_4537,N_4331,N_4398);
nand U4538 (N_4538,N_4474,N_4340);
nor U4539 (N_4539,N_4330,N_4344);
or U4540 (N_4540,N_4336,N_4440);
xor U4541 (N_4541,N_4407,N_4445);
or U4542 (N_4542,N_4429,N_4477);
nand U4543 (N_4543,N_4443,N_4390);
xnor U4544 (N_4544,N_4420,N_4394);
nor U4545 (N_4545,N_4369,N_4460);
and U4546 (N_4546,N_4370,N_4441);
xor U4547 (N_4547,N_4413,N_4383);
and U4548 (N_4548,N_4454,N_4439);
or U4549 (N_4549,N_4365,N_4437);
xnor U4550 (N_4550,N_4456,N_4432);
nor U4551 (N_4551,N_4371,N_4342);
xor U4552 (N_4552,N_4472,N_4403);
nand U4553 (N_4553,N_4384,N_4475);
xnor U4554 (N_4554,N_4468,N_4364);
or U4555 (N_4555,N_4321,N_4469);
or U4556 (N_4556,N_4470,N_4442);
nor U4557 (N_4557,N_4361,N_4424);
nand U4558 (N_4558,N_4391,N_4428);
xor U4559 (N_4559,N_4473,N_4345);
or U4560 (N_4560,N_4425,N_4353);
and U4561 (N_4561,N_4442,N_4349);
nor U4562 (N_4562,N_4451,N_4363);
xnor U4563 (N_4563,N_4471,N_4387);
xor U4564 (N_4564,N_4430,N_4429);
nor U4565 (N_4565,N_4362,N_4475);
xor U4566 (N_4566,N_4392,N_4460);
or U4567 (N_4567,N_4371,N_4469);
and U4568 (N_4568,N_4340,N_4427);
nor U4569 (N_4569,N_4367,N_4476);
nand U4570 (N_4570,N_4474,N_4343);
nor U4571 (N_4571,N_4331,N_4396);
or U4572 (N_4572,N_4408,N_4320);
nand U4573 (N_4573,N_4447,N_4478);
or U4574 (N_4574,N_4455,N_4364);
or U4575 (N_4575,N_4337,N_4458);
and U4576 (N_4576,N_4369,N_4426);
nand U4577 (N_4577,N_4433,N_4437);
xnor U4578 (N_4578,N_4329,N_4392);
nor U4579 (N_4579,N_4411,N_4391);
xnor U4580 (N_4580,N_4357,N_4407);
nor U4581 (N_4581,N_4369,N_4410);
xor U4582 (N_4582,N_4325,N_4356);
xor U4583 (N_4583,N_4365,N_4436);
xnor U4584 (N_4584,N_4452,N_4397);
nand U4585 (N_4585,N_4393,N_4370);
and U4586 (N_4586,N_4406,N_4444);
and U4587 (N_4587,N_4416,N_4322);
nand U4588 (N_4588,N_4366,N_4372);
nor U4589 (N_4589,N_4331,N_4336);
xnor U4590 (N_4590,N_4430,N_4380);
and U4591 (N_4591,N_4455,N_4367);
or U4592 (N_4592,N_4443,N_4429);
nor U4593 (N_4593,N_4473,N_4446);
and U4594 (N_4594,N_4371,N_4403);
xnor U4595 (N_4595,N_4340,N_4459);
or U4596 (N_4596,N_4419,N_4464);
xnor U4597 (N_4597,N_4392,N_4361);
or U4598 (N_4598,N_4364,N_4325);
nand U4599 (N_4599,N_4439,N_4398);
nor U4600 (N_4600,N_4460,N_4449);
nand U4601 (N_4601,N_4367,N_4353);
and U4602 (N_4602,N_4418,N_4399);
or U4603 (N_4603,N_4374,N_4465);
and U4604 (N_4604,N_4462,N_4349);
xnor U4605 (N_4605,N_4454,N_4402);
nor U4606 (N_4606,N_4416,N_4333);
and U4607 (N_4607,N_4434,N_4381);
and U4608 (N_4608,N_4464,N_4417);
or U4609 (N_4609,N_4372,N_4376);
and U4610 (N_4610,N_4461,N_4409);
xnor U4611 (N_4611,N_4359,N_4344);
or U4612 (N_4612,N_4330,N_4462);
or U4613 (N_4613,N_4337,N_4377);
and U4614 (N_4614,N_4450,N_4476);
xnor U4615 (N_4615,N_4420,N_4417);
or U4616 (N_4616,N_4415,N_4419);
and U4617 (N_4617,N_4440,N_4477);
xnor U4618 (N_4618,N_4383,N_4467);
or U4619 (N_4619,N_4461,N_4399);
xor U4620 (N_4620,N_4453,N_4459);
nand U4621 (N_4621,N_4400,N_4367);
nor U4622 (N_4622,N_4444,N_4394);
nor U4623 (N_4623,N_4403,N_4451);
nand U4624 (N_4624,N_4326,N_4446);
nand U4625 (N_4625,N_4365,N_4414);
nor U4626 (N_4626,N_4378,N_4375);
nor U4627 (N_4627,N_4391,N_4405);
xnor U4628 (N_4628,N_4474,N_4338);
and U4629 (N_4629,N_4357,N_4365);
and U4630 (N_4630,N_4342,N_4367);
or U4631 (N_4631,N_4437,N_4438);
xor U4632 (N_4632,N_4353,N_4468);
or U4633 (N_4633,N_4407,N_4392);
or U4634 (N_4634,N_4389,N_4420);
xnor U4635 (N_4635,N_4335,N_4427);
and U4636 (N_4636,N_4363,N_4465);
or U4637 (N_4637,N_4435,N_4343);
nand U4638 (N_4638,N_4330,N_4352);
nand U4639 (N_4639,N_4441,N_4352);
or U4640 (N_4640,N_4635,N_4632);
nor U4641 (N_4641,N_4617,N_4506);
xor U4642 (N_4642,N_4624,N_4505);
and U4643 (N_4643,N_4529,N_4552);
nand U4644 (N_4644,N_4562,N_4571);
nor U4645 (N_4645,N_4502,N_4492);
nor U4646 (N_4646,N_4491,N_4511);
nor U4647 (N_4647,N_4582,N_4545);
xor U4648 (N_4648,N_4493,N_4533);
nor U4649 (N_4649,N_4621,N_4498);
nor U4650 (N_4650,N_4589,N_4625);
nor U4651 (N_4651,N_4541,N_4583);
nor U4652 (N_4652,N_4549,N_4577);
or U4653 (N_4653,N_4480,N_4628);
xor U4654 (N_4654,N_4598,N_4630);
xnor U4655 (N_4655,N_4581,N_4602);
nor U4656 (N_4656,N_4501,N_4608);
xnor U4657 (N_4657,N_4604,N_4567);
and U4658 (N_4658,N_4584,N_4613);
xnor U4659 (N_4659,N_4559,N_4597);
nand U4660 (N_4660,N_4586,N_4560);
nand U4661 (N_4661,N_4623,N_4573);
or U4662 (N_4662,N_4609,N_4481);
and U4663 (N_4663,N_4579,N_4580);
nor U4664 (N_4664,N_4515,N_4553);
xor U4665 (N_4665,N_4527,N_4513);
nand U4666 (N_4666,N_4569,N_4539);
xor U4667 (N_4667,N_4614,N_4575);
nand U4668 (N_4668,N_4530,N_4516);
nor U4669 (N_4669,N_4528,N_4565);
or U4670 (N_4670,N_4546,N_4547);
and U4671 (N_4671,N_4610,N_4524);
nor U4672 (N_4672,N_4537,N_4578);
and U4673 (N_4673,N_4607,N_4522);
nand U4674 (N_4674,N_4568,N_4518);
and U4675 (N_4675,N_4548,N_4519);
or U4676 (N_4676,N_4488,N_4482);
and U4677 (N_4677,N_4600,N_4639);
and U4678 (N_4678,N_4496,N_4558);
and U4679 (N_4679,N_4588,N_4532);
nor U4680 (N_4680,N_4561,N_4633);
nor U4681 (N_4681,N_4542,N_4521);
nand U4682 (N_4682,N_4556,N_4566);
or U4683 (N_4683,N_4626,N_4512);
and U4684 (N_4684,N_4611,N_4574);
nor U4685 (N_4685,N_4509,N_4544);
and U4686 (N_4686,N_4555,N_4629);
nor U4687 (N_4687,N_4536,N_4605);
and U4688 (N_4688,N_4563,N_4520);
nand U4689 (N_4689,N_4592,N_4531);
and U4690 (N_4690,N_4616,N_4483);
and U4691 (N_4691,N_4606,N_4622);
xor U4692 (N_4692,N_4534,N_4551);
or U4693 (N_4693,N_4636,N_4523);
nor U4694 (N_4694,N_4490,N_4538);
or U4695 (N_4695,N_4612,N_4572);
xor U4696 (N_4696,N_4485,N_4638);
and U4697 (N_4697,N_4484,N_4507);
or U4698 (N_4698,N_4601,N_4634);
or U4699 (N_4699,N_4593,N_4618);
xor U4700 (N_4700,N_4525,N_4596);
nand U4701 (N_4701,N_4543,N_4599);
xnor U4702 (N_4702,N_4486,N_4576);
and U4703 (N_4703,N_4500,N_4494);
nor U4704 (N_4704,N_4503,N_4517);
or U4705 (N_4705,N_4627,N_4510);
nand U4706 (N_4706,N_4497,N_4514);
nand U4707 (N_4707,N_4620,N_4564);
or U4708 (N_4708,N_4631,N_4508);
or U4709 (N_4709,N_4619,N_4637);
nand U4710 (N_4710,N_4557,N_4526);
nor U4711 (N_4711,N_4504,N_4570);
xnor U4712 (N_4712,N_4499,N_4535);
nand U4713 (N_4713,N_4489,N_4591);
nor U4714 (N_4714,N_4615,N_4540);
and U4715 (N_4715,N_4587,N_4550);
xor U4716 (N_4716,N_4603,N_4554);
xnor U4717 (N_4717,N_4595,N_4585);
or U4718 (N_4718,N_4594,N_4487);
nand U4719 (N_4719,N_4495,N_4590);
or U4720 (N_4720,N_4619,N_4570);
xnor U4721 (N_4721,N_4483,N_4575);
and U4722 (N_4722,N_4585,N_4604);
xnor U4723 (N_4723,N_4489,N_4561);
nor U4724 (N_4724,N_4502,N_4484);
nor U4725 (N_4725,N_4481,N_4589);
and U4726 (N_4726,N_4551,N_4526);
xor U4727 (N_4727,N_4588,N_4487);
nor U4728 (N_4728,N_4506,N_4627);
and U4729 (N_4729,N_4532,N_4639);
and U4730 (N_4730,N_4590,N_4535);
and U4731 (N_4731,N_4610,N_4584);
xnor U4732 (N_4732,N_4537,N_4483);
xor U4733 (N_4733,N_4592,N_4538);
and U4734 (N_4734,N_4509,N_4609);
nand U4735 (N_4735,N_4600,N_4543);
nor U4736 (N_4736,N_4560,N_4543);
and U4737 (N_4737,N_4528,N_4605);
nand U4738 (N_4738,N_4494,N_4502);
and U4739 (N_4739,N_4606,N_4488);
xnor U4740 (N_4740,N_4480,N_4561);
nand U4741 (N_4741,N_4543,N_4635);
or U4742 (N_4742,N_4621,N_4540);
xor U4743 (N_4743,N_4572,N_4535);
or U4744 (N_4744,N_4537,N_4507);
or U4745 (N_4745,N_4481,N_4627);
nand U4746 (N_4746,N_4618,N_4553);
xor U4747 (N_4747,N_4540,N_4536);
xnor U4748 (N_4748,N_4533,N_4515);
and U4749 (N_4749,N_4539,N_4584);
nand U4750 (N_4750,N_4499,N_4521);
nor U4751 (N_4751,N_4625,N_4638);
xnor U4752 (N_4752,N_4601,N_4576);
and U4753 (N_4753,N_4604,N_4580);
or U4754 (N_4754,N_4500,N_4635);
nand U4755 (N_4755,N_4503,N_4494);
or U4756 (N_4756,N_4491,N_4547);
nand U4757 (N_4757,N_4631,N_4578);
nand U4758 (N_4758,N_4508,N_4522);
and U4759 (N_4759,N_4516,N_4572);
xor U4760 (N_4760,N_4530,N_4535);
and U4761 (N_4761,N_4554,N_4587);
nand U4762 (N_4762,N_4638,N_4608);
xnor U4763 (N_4763,N_4519,N_4599);
nor U4764 (N_4764,N_4519,N_4514);
nor U4765 (N_4765,N_4544,N_4506);
nor U4766 (N_4766,N_4510,N_4529);
and U4767 (N_4767,N_4591,N_4560);
or U4768 (N_4768,N_4489,N_4617);
and U4769 (N_4769,N_4480,N_4502);
or U4770 (N_4770,N_4525,N_4610);
xor U4771 (N_4771,N_4626,N_4482);
or U4772 (N_4772,N_4483,N_4584);
and U4773 (N_4773,N_4572,N_4554);
and U4774 (N_4774,N_4611,N_4575);
or U4775 (N_4775,N_4561,N_4505);
xor U4776 (N_4776,N_4530,N_4576);
nor U4777 (N_4777,N_4548,N_4500);
nand U4778 (N_4778,N_4568,N_4612);
xor U4779 (N_4779,N_4561,N_4587);
and U4780 (N_4780,N_4538,N_4598);
or U4781 (N_4781,N_4566,N_4549);
or U4782 (N_4782,N_4486,N_4495);
xor U4783 (N_4783,N_4579,N_4511);
or U4784 (N_4784,N_4614,N_4583);
nor U4785 (N_4785,N_4591,N_4625);
nand U4786 (N_4786,N_4633,N_4615);
or U4787 (N_4787,N_4484,N_4543);
xnor U4788 (N_4788,N_4494,N_4486);
or U4789 (N_4789,N_4539,N_4576);
nor U4790 (N_4790,N_4599,N_4541);
or U4791 (N_4791,N_4626,N_4561);
xnor U4792 (N_4792,N_4582,N_4557);
nor U4793 (N_4793,N_4488,N_4559);
nor U4794 (N_4794,N_4637,N_4541);
or U4795 (N_4795,N_4636,N_4603);
nand U4796 (N_4796,N_4549,N_4618);
xnor U4797 (N_4797,N_4532,N_4555);
xor U4798 (N_4798,N_4590,N_4525);
and U4799 (N_4799,N_4515,N_4532);
nand U4800 (N_4800,N_4728,N_4748);
xnor U4801 (N_4801,N_4788,N_4755);
xor U4802 (N_4802,N_4768,N_4777);
nand U4803 (N_4803,N_4761,N_4749);
or U4804 (N_4804,N_4782,N_4776);
nand U4805 (N_4805,N_4715,N_4785);
and U4806 (N_4806,N_4690,N_4790);
nand U4807 (N_4807,N_4666,N_4744);
and U4808 (N_4808,N_4796,N_4721);
and U4809 (N_4809,N_4780,N_4798);
nor U4810 (N_4810,N_4651,N_4713);
and U4811 (N_4811,N_4732,N_4650);
and U4812 (N_4812,N_4704,N_4696);
xnor U4813 (N_4813,N_4694,N_4792);
nand U4814 (N_4814,N_4747,N_4655);
or U4815 (N_4815,N_4664,N_4712);
or U4816 (N_4816,N_4656,N_4675);
nand U4817 (N_4817,N_4671,N_4654);
and U4818 (N_4818,N_4731,N_4706);
and U4819 (N_4819,N_4778,N_4652);
or U4820 (N_4820,N_4701,N_4789);
and U4821 (N_4821,N_4719,N_4733);
or U4822 (N_4822,N_4767,N_4692);
xnor U4823 (N_4823,N_4759,N_4647);
and U4824 (N_4824,N_4663,N_4783);
or U4825 (N_4825,N_4668,N_4659);
xor U4826 (N_4826,N_4725,N_4724);
and U4827 (N_4827,N_4691,N_4660);
nor U4828 (N_4828,N_4645,N_4794);
and U4829 (N_4829,N_4752,N_4695);
nor U4830 (N_4830,N_4765,N_4770);
or U4831 (N_4831,N_4779,N_4750);
nor U4832 (N_4832,N_4722,N_4684);
nor U4833 (N_4833,N_4709,N_4677);
nand U4834 (N_4834,N_4689,N_4723);
and U4835 (N_4835,N_4760,N_4649);
or U4836 (N_4836,N_4742,N_4717);
nand U4837 (N_4837,N_4658,N_4730);
nor U4838 (N_4838,N_4795,N_4705);
or U4839 (N_4839,N_4754,N_4680);
nor U4840 (N_4840,N_4784,N_4769);
nand U4841 (N_4841,N_4710,N_4799);
xnor U4842 (N_4842,N_4640,N_4716);
and U4843 (N_4843,N_4676,N_4703);
nor U4844 (N_4844,N_4737,N_4787);
xor U4845 (N_4845,N_4682,N_4657);
nand U4846 (N_4846,N_4775,N_4688);
and U4847 (N_4847,N_4672,N_4758);
and U4848 (N_4848,N_4702,N_4653);
xnor U4849 (N_4849,N_4697,N_4674);
nor U4850 (N_4850,N_4735,N_4757);
and U4851 (N_4851,N_4736,N_4700);
xnor U4852 (N_4852,N_4686,N_4756);
nand U4853 (N_4853,N_4642,N_4727);
and U4854 (N_4854,N_4766,N_4739);
and U4855 (N_4855,N_4726,N_4648);
nand U4856 (N_4856,N_4687,N_4774);
or U4857 (N_4857,N_4745,N_4797);
nand U4858 (N_4858,N_4746,N_4667);
nand U4859 (N_4859,N_4771,N_4681);
xor U4860 (N_4860,N_4665,N_4643);
and U4861 (N_4861,N_4644,N_4707);
nand U4862 (N_4862,N_4678,N_4772);
and U4863 (N_4863,N_4669,N_4699);
nor U4864 (N_4864,N_4762,N_4734);
or U4865 (N_4865,N_4773,N_4793);
or U4866 (N_4866,N_4683,N_4670);
and U4867 (N_4867,N_4741,N_4679);
or U4868 (N_4868,N_4693,N_4763);
or U4869 (N_4869,N_4743,N_4791);
nor U4870 (N_4870,N_4661,N_4729);
and U4871 (N_4871,N_4740,N_4641);
xnor U4872 (N_4872,N_4714,N_4685);
and U4873 (N_4873,N_4718,N_4786);
xnor U4874 (N_4874,N_4781,N_4753);
or U4875 (N_4875,N_4673,N_4662);
and U4876 (N_4876,N_4711,N_4646);
and U4877 (N_4877,N_4720,N_4708);
nand U4878 (N_4878,N_4764,N_4751);
nor U4879 (N_4879,N_4698,N_4738);
nand U4880 (N_4880,N_4783,N_4748);
nor U4881 (N_4881,N_4796,N_4763);
nand U4882 (N_4882,N_4697,N_4760);
nand U4883 (N_4883,N_4771,N_4753);
nand U4884 (N_4884,N_4689,N_4799);
and U4885 (N_4885,N_4782,N_4760);
nor U4886 (N_4886,N_4662,N_4694);
and U4887 (N_4887,N_4771,N_4644);
nand U4888 (N_4888,N_4640,N_4715);
nor U4889 (N_4889,N_4644,N_4790);
nand U4890 (N_4890,N_4664,N_4671);
nand U4891 (N_4891,N_4734,N_4698);
or U4892 (N_4892,N_4663,N_4660);
and U4893 (N_4893,N_4764,N_4672);
and U4894 (N_4894,N_4686,N_4781);
and U4895 (N_4895,N_4671,N_4764);
nor U4896 (N_4896,N_4773,N_4652);
nand U4897 (N_4897,N_4734,N_4749);
and U4898 (N_4898,N_4684,N_4790);
xnor U4899 (N_4899,N_4719,N_4678);
nand U4900 (N_4900,N_4737,N_4771);
or U4901 (N_4901,N_4712,N_4786);
or U4902 (N_4902,N_4767,N_4699);
and U4903 (N_4903,N_4742,N_4713);
xnor U4904 (N_4904,N_4646,N_4654);
or U4905 (N_4905,N_4779,N_4710);
xor U4906 (N_4906,N_4736,N_4687);
nand U4907 (N_4907,N_4765,N_4691);
or U4908 (N_4908,N_4675,N_4689);
nor U4909 (N_4909,N_4776,N_4668);
nand U4910 (N_4910,N_4747,N_4741);
or U4911 (N_4911,N_4773,N_4686);
nand U4912 (N_4912,N_4714,N_4651);
xor U4913 (N_4913,N_4768,N_4645);
and U4914 (N_4914,N_4660,N_4680);
nand U4915 (N_4915,N_4743,N_4646);
xnor U4916 (N_4916,N_4772,N_4790);
nor U4917 (N_4917,N_4667,N_4754);
nand U4918 (N_4918,N_4763,N_4732);
nand U4919 (N_4919,N_4659,N_4683);
or U4920 (N_4920,N_4708,N_4650);
nand U4921 (N_4921,N_4661,N_4726);
or U4922 (N_4922,N_4755,N_4747);
or U4923 (N_4923,N_4710,N_4697);
nand U4924 (N_4924,N_4734,N_4788);
xnor U4925 (N_4925,N_4694,N_4655);
nand U4926 (N_4926,N_4727,N_4647);
nand U4927 (N_4927,N_4708,N_4766);
and U4928 (N_4928,N_4774,N_4700);
or U4929 (N_4929,N_4697,N_4745);
or U4930 (N_4930,N_4640,N_4790);
or U4931 (N_4931,N_4745,N_4783);
or U4932 (N_4932,N_4703,N_4656);
and U4933 (N_4933,N_4705,N_4749);
and U4934 (N_4934,N_4653,N_4736);
xor U4935 (N_4935,N_4736,N_4645);
xor U4936 (N_4936,N_4727,N_4798);
or U4937 (N_4937,N_4795,N_4699);
nor U4938 (N_4938,N_4681,N_4737);
and U4939 (N_4939,N_4716,N_4764);
nand U4940 (N_4940,N_4739,N_4758);
or U4941 (N_4941,N_4778,N_4796);
or U4942 (N_4942,N_4749,N_4756);
xor U4943 (N_4943,N_4699,N_4734);
nand U4944 (N_4944,N_4670,N_4779);
nand U4945 (N_4945,N_4752,N_4798);
and U4946 (N_4946,N_4663,N_4706);
or U4947 (N_4947,N_4762,N_4729);
and U4948 (N_4948,N_4739,N_4724);
or U4949 (N_4949,N_4772,N_4679);
nor U4950 (N_4950,N_4735,N_4669);
xnor U4951 (N_4951,N_4679,N_4743);
and U4952 (N_4952,N_4724,N_4694);
nor U4953 (N_4953,N_4640,N_4738);
nor U4954 (N_4954,N_4665,N_4789);
or U4955 (N_4955,N_4717,N_4722);
and U4956 (N_4956,N_4769,N_4744);
xnor U4957 (N_4957,N_4771,N_4662);
xnor U4958 (N_4958,N_4678,N_4657);
and U4959 (N_4959,N_4647,N_4730);
nand U4960 (N_4960,N_4806,N_4828);
xnor U4961 (N_4961,N_4921,N_4894);
or U4962 (N_4962,N_4863,N_4928);
and U4963 (N_4963,N_4835,N_4889);
and U4964 (N_4964,N_4900,N_4862);
and U4965 (N_4965,N_4896,N_4949);
or U4966 (N_4966,N_4925,N_4833);
xor U4967 (N_4967,N_4881,N_4824);
nand U4968 (N_4968,N_4887,N_4866);
or U4969 (N_4969,N_4830,N_4868);
or U4970 (N_4970,N_4829,N_4870);
xor U4971 (N_4971,N_4879,N_4840);
or U4972 (N_4972,N_4893,N_4916);
nor U4973 (N_4973,N_4853,N_4860);
nor U4974 (N_4974,N_4891,N_4836);
nand U4975 (N_4975,N_4924,N_4895);
nor U4976 (N_4976,N_4848,N_4857);
nand U4977 (N_4977,N_4858,N_4826);
nor U4978 (N_4978,N_4953,N_4904);
and U4979 (N_4979,N_4909,N_4855);
or U4980 (N_4980,N_4934,N_4849);
and U4981 (N_4981,N_4902,N_4841);
nand U4982 (N_4982,N_4832,N_4801);
or U4983 (N_4983,N_4851,N_4910);
nand U4984 (N_4984,N_4913,N_4956);
nor U4985 (N_4985,N_4877,N_4922);
and U4986 (N_4986,N_4936,N_4897);
nor U4987 (N_4987,N_4844,N_4814);
or U4988 (N_4988,N_4873,N_4861);
nand U4989 (N_4989,N_4867,N_4952);
xor U4990 (N_4990,N_4937,N_4957);
nand U4991 (N_4991,N_4959,N_4819);
nand U4992 (N_4992,N_4815,N_4812);
and U4993 (N_4993,N_4874,N_4808);
and U4994 (N_4994,N_4818,N_4883);
xor U4995 (N_4995,N_4923,N_4906);
nor U4996 (N_4996,N_4856,N_4859);
xor U4997 (N_4997,N_4898,N_4875);
xor U4998 (N_4998,N_4813,N_4825);
nor U4999 (N_4999,N_4847,N_4876);
xnor U5000 (N_5000,N_4912,N_4842);
or U5001 (N_5001,N_4948,N_4920);
xor U5002 (N_5002,N_4886,N_4890);
and U5003 (N_5003,N_4929,N_4919);
xnor U5004 (N_5004,N_4803,N_4831);
or U5005 (N_5005,N_4809,N_4943);
nand U5006 (N_5006,N_4892,N_4838);
nand U5007 (N_5007,N_4872,N_4880);
or U5008 (N_5008,N_4869,N_4946);
and U5009 (N_5009,N_4945,N_4944);
xnor U5010 (N_5010,N_4811,N_4914);
or U5011 (N_5011,N_4843,N_4822);
xnor U5012 (N_5012,N_4800,N_4820);
nand U5013 (N_5013,N_4882,N_4804);
xor U5014 (N_5014,N_4915,N_4938);
and U5015 (N_5015,N_4927,N_4888);
or U5016 (N_5016,N_4878,N_4823);
xor U5017 (N_5017,N_4954,N_4852);
nor U5018 (N_5018,N_4930,N_4865);
nand U5019 (N_5019,N_4940,N_4931);
nand U5020 (N_5020,N_4807,N_4810);
nor U5021 (N_5021,N_4850,N_4839);
nand U5022 (N_5022,N_4942,N_4926);
and U5023 (N_5023,N_4816,N_4941);
nor U5024 (N_5024,N_4854,N_4951);
nand U5025 (N_5025,N_4939,N_4834);
nand U5026 (N_5026,N_4908,N_4947);
and U5027 (N_5027,N_4845,N_4950);
and U5028 (N_5028,N_4905,N_4958);
xnor U5029 (N_5029,N_4846,N_4933);
xor U5030 (N_5030,N_4899,N_4802);
xnor U5031 (N_5031,N_4901,N_4955);
xor U5032 (N_5032,N_4821,N_4885);
nor U5033 (N_5033,N_4884,N_4817);
and U5034 (N_5034,N_4935,N_4907);
xor U5035 (N_5035,N_4917,N_4918);
or U5036 (N_5036,N_4805,N_4903);
and U5037 (N_5037,N_4864,N_4827);
and U5038 (N_5038,N_4932,N_4871);
nand U5039 (N_5039,N_4911,N_4837);
nand U5040 (N_5040,N_4869,N_4812);
xnor U5041 (N_5041,N_4801,N_4916);
xnor U5042 (N_5042,N_4814,N_4836);
and U5043 (N_5043,N_4810,N_4922);
and U5044 (N_5044,N_4865,N_4852);
nand U5045 (N_5045,N_4828,N_4879);
and U5046 (N_5046,N_4836,N_4908);
nand U5047 (N_5047,N_4877,N_4957);
and U5048 (N_5048,N_4820,N_4818);
and U5049 (N_5049,N_4871,N_4803);
xor U5050 (N_5050,N_4882,N_4903);
and U5051 (N_5051,N_4918,N_4955);
and U5052 (N_5052,N_4870,N_4814);
xor U5053 (N_5053,N_4827,N_4910);
nor U5054 (N_5054,N_4834,N_4835);
or U5055 (N_5055,N_4838,N_4876);
nand U5056 (N_5056,N_4846,N_4911);
and U5057 (N_5057,N_4817,N_4938);
xor U5058 (N_5058,N_4815,N_4801);
xor U5059 (N_5059,N_4953,N_4830);
or U5060 (N_5060,N_4898,N_4868);
nand U5061 (N_5061,N_4820,N_4846);
and U5062 (N_5062,N_4945,N_4894);
nor U5063 (N_5063,N_4871,N_4851);
nor U5064 (N_5064,N_4803,N_4855);
nor U5065 (N_5065,N_4834,N_4885);
and U5066 (N_5066,N_4947,N_4818);
or U5067 (N_5067,N_4831,N_4887);
and U5068 (N_5068,N_4822,N_4866);
and U5069 (N_5069,N_4943,N_4900);
xor U5070 (N_5070,N_4846,N_4829);
xnor U5071 (N_5071,N_4842,N_4836);
nor U5072 (N_5072,N_4849,N_4947);
or U5073 (N_5073,N_4867,N_4932);
nand U5074 (N_5074,N_4959,N_4931);
or U5075 (N_5075,N_4846,N_4900);
nand U5076 (N_5076,N_4873,N_4816);
nand U5077 (N_5077,N_4891,N_4811);
nand U5078 (N_5078,N_4940,N_4877);
or U5079 (N_5079,N_4894,N_4939);
and U5080 (N_5080,N_4906,N_4900);
or U5081 (N_5081,N_4802,N_4892);
xor U5082 (N_5082,N_4898,N_4944);
nor U5083 (N_5083,N_4867,N_4847);
xor U5084 (N_5084,N_4956,N_4882);
and U5085 (N_5085,N_4838,N_4817);
nand U5086 (N_5086,N_4828,N_4857);
and U5087 (N_5087,N_4932,N_4879);
or U5088 (N_5088,N_4877,N_4862);
nand U5089 (N_5089,N_4939,N_4875);
and U5090 (N_5090,N_4897,N_4911);
and U5091 (N_5091,N_4827,N_4853);
nor U5092 (N_5092,N_4945,N_4805);
or U5093 (N_5093,N_4886,N_4904);
or U5094 (N_5094,N_4943,N_4848);
nand U5095 (N_5095,N_4857,N_4805);
and U5096 (N_5096,N_4834,N_4826);
or U5097 (N_5097,N_4808,N_4800);
nor U5098 (N_5098,N_4815,N_4948);
nand U5099 (N_5099,N_4869,N_4867);
nor U5100 (N_5100,N_4933,N_4910);
nor U5101 (N_5101,N_4930,N_4830);
nand U5102 (N_5102,N_4860,N_4872);
nor U5103 (N_5103,N_4830,N_4858);
nand U5104 (N_5104,N_4803,N_4920);
and U5105 (N_5105,N_4824,N_4953);
nand U5106 (N_5106,N_4924,N_4856);
and U5107 (N_5107,N_4832,N_4887);
or U5108 (N_5108,N_4819,N_4800);
nor U5109 (N_5109,N_4806,N_4853);
xor U5110 (N_5110,N_4909,N_4926);
and U5111 (N_5111,N_4912,N_4920);
nor U5112 (N_5112,N_4910,N_4934);
xor U5113 (N_5113,N_4953,N_4835);
or U5114 (N_5114,N_4947,N_4837);
nand U5115 (N_5115,N_4822,N_4944);
xnor U5116 (N_5116,N_4911,N_4925);
xnor U5117 (N_5117,N_4873,N_4869);
nand U5118 (N_5118,N_4948,N_4808);
or U5119 (N_5119,N_4944,N_4916);
nor U5120 (N_5120,N_5010,N_5040);
and U5121 (N_5121,N_5029,N_5094);
nor U5122 (N_5122,N_4995,N_5116);
or U5123 (N_5123,N_5103,N_5100);
nor U5124 (N_5124,N_5046,N_5048);
nand U5125 (N_5125,N_5024,N_4965);
xor U5126 (N_5126,N_5030,N_5035);
xnor U5127 (N_5127,N_5004,N_5033);
and U5128 (N_5128,N_5070,N_4990);
or U5129 (N_5129,N_5003,N_4977);
xor U5130 (N_5130,N_5013,N_5002);
nand U5131 (N_5131,N_5025,N_4988);
nand U5132 (N_5132,N_5015,N_5084);
xnor U5133 (N_5133,N_4973,N_5011);
or U5134 (N_5134,N_5026,N_5108);
xor U5135 (N_5135,N_5064,N_4997);
nor U5136 (N_5136,N_5078,N_4981);
nor U5137 (N_5137,N_5032,N_4991);
and U5138 (N_5138,N_5049,N_5117);
and U5139 (N_5139,N_5088,N_4970);
or U5140 (N_5140,N_5069,N_5045);
xnor U5141 (N_5141,N_5068,N_5034);
or U5142 (N_5142,N_5067,N_5089);
and U5143 (N_5143,N_5060,N_5096);
or U5144 (N_5144,N_4975,N_5043);
nand U5145 (N_5145,N_5053,N_4974);
or U5146 (N_5146,N_5031,N_5039);
and U5147 (N_5147,N_4966,N_5090);
nand U5148 (N_5148,N_5109,N_5056);
nand U5149 (N_5149,N_5110,N_5000);
and U5150 (N_5150,N_5087,N_5072);
and U5151 (N_5151,N_4964,N_4982);
and U5152 (N_5152,N_5057,N_5106);
xor U5153 (N_5153,N_5023,N_4987);
or U5154 (N_5154,N_5085,N_4983);
and U5155 (N_5155,N_5073,N_5018);
or U5156 (N_5156,N_5092,N_5062);
nor U5157 (N_5157,N_5017,N_4968);
or U5158 (N_5158,N_4994,N_5079);
or U5159 (N_5159,N_5021,N_5065);
and U5160 (N_5160,N_5008,N_4989);
nand U5161 (N_5161,N_5077,N_4992);
or U5162 (N_5162,N_4993,N_4960);
or U5163 (N_5163,N_5050,N_5022);
or U5164 (N_5164,N_5055,N_4980);
or U5165 (N_5165,N_5047,N_5012);
and U5166 (N_5166,N_4984,N_5111);
or U5167 (N_5167,N_4979,N_5093);
nor U5168 (N_5168,N_5037,N_5083);
or U5169 (N_5169,N_4985,N_5063);
nor U5170 (N_5170,N_5098,N_5006);
and U5171 (N_5171,N_5014,N_4986);
nand U5172 (N_5172,N_4961,N_5105);
or U5173 (N_5173,N_5099,N_5066);
xnor U5174 (N_5174,N_5076,N_5054);
and U5175 (N_5175,N_5016,N_5028);
xnor U5176 (N_5176,N_5005,N_4996);
nand U5177 (N_5177,N_5086,N_5052);
nor U5178 (N_5178,N_5041,N_5020);
nand U5179 (N_5179,N_5081,N_5059);
nor U5180 (N_5180,N_5042,N_5009);
and U5181 (N_5181,N_4967,N_5118);
or U5182 (N_5182,N_5101,N_4978);
nand U5183 (N_5183,N_5095,N_5027);
nor U5184 (N_5184,N_5058,N_5082);
nand U5185 (N_5185,N_5007,N_5019);
or U5186 (N_5186,N_4972,N_5038);
nand U5187 (N_5187,N_5102,N_5051);
nand U5188 (N_5188,N_5001,N_4969);
and U5189 (N_5189,N_5113,N_5075);
xnor U5190 (N_5190,N_5119,N_5044);
and U5191 (N_5191,N_5104,N_4976);
nand U5192 (N_5192,N_5112,N_5080);
nor U5193 (N_5193,N_4962,N_4999);
nor U5194 (N_5194,N_4971,N_5074);
nand U5195 (N_5195,N_5097,N_5091);
nand U5196 (N_5196,N_5061,N_5107);
xnor U5197 (N_5197,N_5036,N_4998);
nand U5198 (N_5198,N_5071,N_4963);
or U5199 (N_5199,N_5114,N_5115);
xnor U5200 (N_5200,N_4978,N_5099);
and U5201 (N_5201,N_5099,N_4986);
xor U5202 (N_5202,N_5117,N_4970);
or U5203 (N_5203,N_5051,N_5081);
nor U5204 (N_5204,N_5015,N_5020);
xor U5205 (N_5205,N_5086,N_5009);
nand U5206 (N_5206,N_4965,N_4993);
xor U5207 (N_5207,N_5012,N_5069);
xnor U5208 (N_5208,N_5035,N_5073);
nor U5209 (N_5209,N_5051,N_5016);
nor U5210 (N_5210,N_5047,N_5070);
xor U5211 (N_5211,N_5050,N_4989);
and U5212 (N_5212,N_5069,N_4976);
and U5213 (N_5213,N_5007,N_5011);
nor U5214 (N_5214,N_5093,N_5055);
and U5215 (N_5215,N_5063,N_4968);
nand U5216 (N_5216,N_5091,N_5083);
xor U5217 (N_5217,N_5064,N_5023);
xnor U5218 (N_5218,N_5014,N_5057);
or U5219 (N_5219,N_4967,N_5105);
nor U5220 (N_5220,N_5045,N_5074);
and U5221 (N_5221,N_5080,N_5101);
and U5222 (N_5222,N_4990,N_5030);
and U5223 (N_5223,N_5103,N_4981);
nand U5224 (N_5224,N_5011,N_5066);
xnor U5225 (N_5225,N_5046,N_5105);
nor U5226 (N_5226,N_5033,N_5069);
nand U5227 (N_5227,N_4962,N_5110);
or U5228 (N_5228,N_4978,N_5089);
nor U5229 (N_5229,N_5050,N_4961);
xnor U5230 (N_5230,N_5084,N_4961);
nor U5231 (N_5231,N_4996,N_4960);
nor U5232 (N_5232,N_5089,N_4960);
nand U5233 (N_5233,N_4981,N_5009);
xnor U5234 (N_5234,N_4980,N_4975);
xnor U5235 (N_5235,N_5027,N_4972);
xor U5236 (N_5236,N_5089,N_5103);
nor U5237 (N_5237,N_5016,N_4987);
xor U5238 (N_5238,N_5099,N_4983);
and U5239 (N_5239,N_5000,N_5032);
nor U5240 (N_5240,N_5101,N_5056);
and U5241 (N_5241,N_4963,N_5089);
xor U5242 (N_5242,N_4985,N_4976);
nand U5243 (N_5243,N_5026,N_4993);
and U5244 (N_5244,N_4998,N_5074);
or U5245 (N_5245,N_5102,N_4970);
or U5246 (N_5246,N_5032,N_5065);
and U5247 (N_5247,N_5091,N_5052);
xnor U5248 (N_5248,N_5042,N_4999);
nand U5249 (N_5249,N_4972,N_4961);
or U5250 (N_5250,N_4982,N_5013);
nand U5251 (N_5251,N_4961,N_5040);
nand U5252 (N_5252,N_5067,N_5079);
and U5253 (N_5253,N_5068,N_5062);
and U5254 (N_5254,N_4988,N_5017);
nand U5255 (N_5255,N_5076,N_5098);
nor U5256 (N_5256,N_5071,N_5063);
and U5257 (N_5257,N_5088,N_5097);
or U5258 (N_5258,N_5048,N_4994);
nand U5259 (N_5259,N_5095,N_5039);
xor U5260 (N_5260,N_4986,N_5106);
nor U5261 (N_5261,N_4999,N_5114);
and U5262 (N_5262,N_5047,N_5094);
nor U5263 (N_5263,N_5103,N_5080);
and U5264 (N_5264,N_5037,N_5084);
nand U5265 (N_5265,N_5049,N_4978);
xnor U5266 (N_5266,N_4979,N_5115);
xor U5267 (N_5267,N_5057,N_4988);
xnor U5268 (N_5268,N_5052,N_5075);
nand U5269 (N_5269,N_5069,N_4995);
or U5270 (N_5270,N_5058,N_4994);
or U5271 (N_5271,N_4991,N_5009);
xor U5272 (N_5272,N_5109,N_5110);
and U5273 (N_5273,N_5012,N_4987);
nor U5274 (N_5274,N_5102,N_5041);
and U5275 (N_5275,N_5093,N_5005);
nand U5276 (N_5276,N_4998,N_5004);
and U5277 (N_5277,N_5102,N_5087);
xnor U5278 (N_5278,N_5078,N_5039);
xor U5279 (N_5279,N_5110,N_5074);
nor U5280 (N_5280,N_5213,N_5171);
nor U5281 (N_5281,N_5216,N_5223);
or U5282 (N_5282,N_5265,N_5148);
and U5283 (N_5283,N_5184,N_5207);
nor U5284 (N_5284,N_5256,N_5212);
and U5285 (N_5285,N_5166,N_5120);
and U5286 (N_5286,N_5152,N_5214);
and U5287 (N_5287,N_5160,N_5122);
nor U5288 (N_5288,N_5201,N_5240);
nor U5289 (N_5289,N_5276,N_5204);
nor U5290 (N_5290,N_5170,N_5225);
or U5291 (N_5291,N_5134,N_5217);
nor U5292 (N_5292,N_5180,N_5215);
nor U5293 (N_5293,N_5123,N_5261);
xor U5294 (N_5294,N_5250,N_5144);
nand U5295 (N_5295,N_5138,N_5202);
nand U5296 (N_5296,N_5177,N_5263);
nand U5297 (N_5297,N_5167,N_5242);
nand U5298 (N_5298,N_5262,N_5222);
xnor U5299 (N_5299,N_5219,N_5271);
nand U5300 (N_5300,N_5231,N_5136);
and U5301 (N_5301,N_5142,N_5158);
or U5302 (N_5302,N_5179,N_5221);
or U5303 (N_5303,N_5198,N_5127);
and U5304 (N_5304,N_5203,N_5189);
and U5305 (N_5305,N_5188,N_5165);
nand U5306 (N_5306,N_5176,N_5257);
or U5307 (N_5307,N_5270,N_5149);
xnor U5308 (N_5308,N_5157,N_5192);
or U5309 (N_5309,N_5133,N_5187);
nor U5310 (N_5310,N_5233,N_5185);
or U5311 (N_5311,N_5156,N_5267);
nor U5312 (N_5312,N_5235,N_5124);
and U5313 (N_5313,N_5255,N_5206);
and U5314 (N_5314,N_5178,N_5135);
or U5315 (N_5315,N_5154,N_5153);
nand U5316 (N_5316,N_5228,N_5232);
or U5317 (N_5317,N_5208,N_5163);
xnor U5318 (N_5318,N_5181,N_5162);
or U5319 (N_5319,N_5139,N_5269);
xnor U5320 (N_5320,N_5248,N_5194);
and U5321 (N_5321,N_5275,N_5183);
xnor U5322 (N_5322,N_5273,N_5258);
or U5323 (N_5323,N_5200,N_5268);
or U5324 (N_5324,N_5229,N_5264);
nor U5325 (N_5325,N_5132,N_5161);
or U5326 (N_5326,N_5141,N_5243);
or U5327 (N_5327,N_5126,N_5199);
or U5328 (N_5328,N_5173,N_5147);
or U5329 (N_5329,N_5237,N_5164);
nor U5330 (N_5330,N_5209,N_5211);
or U5331 (N_5331,N_5140,N_5196);
and U5332 (N_5332,N_5174,N_5131);
xor U5333 (N_5333,N_5279,N_5182);
nor U5334 (N_5334,N_5159,N_5266);
and U5335 (N_5335,N_5252,N_5128);
xor U5336 (N_5336,N_5121,N_5239);
nand U5337 (N_5337,N_5251,N_5253);
xnor U5338 (N_5338,N_5260,N_5278);
nor U5339 (N_5339,N_5227,N_5169);
xor U5340 (N_5340,N_5146,N_5245);
and U5341 (N_5341,N_5175,N_5218);
xnor U5342 (N_5342,N_5220,N_5168);
or U5343 (N_5343,N_5254,N_5259);
nor U5344 (N_5344,N_5155,N_5230);
and U5345 (N_5345,N_5238,N_5151);
nand U5346 (N_5346,N_5137,N_5125);
and U5347 (N_5347,N_5246,N_5150);
nand U5348 (N_5348,N_5186,N_5205);
or U5349 (N_5349,N_5130,N_5241);
nand U5350 (N_5350,N_5197,N_5234);
nor U5351 (N_5351,N_5224,N_5190);
nor U5352 (N_5352,N_5193,N_5247);
nand U5353 (N_5353,N_5145,N_5272);
xor U5354 (N_5354,N_5191,N_5277);
or U5355 (N_5355,N_5143,N_5226);
nand U5356 (N_5356,N_5274,N_5172);
nor U5357 (N_5357,N_5195,N_5129);
or U5358 (N_5358,N_5244,N_5236);
or U5359 (N_5359,N_5249,N_5210);
or U5360 (N_5360,N_5120,N_5257);
nor U5361 (N_5361,N_5226,N_5249);
nor U5362 (N_5362,N_5189,N_5198);
nor U5363 (N_5363,N_5279,N_5273);
xor U5364 (N_5364,N_5176,N_5234);
and U5365 (N_5365,N_5246,N_5198);
or U5366 (N_5366,N_5177,N_5198);
and U5367 (N_5367,N_5242,N_5178);
nor U5368 (N_5368,N_5218,N_5231);
or U5369 (N_5369,N_5234,N_5212);
or U5370 (N_5370,N_5209,N_5134);
nor U5371 (N_5371,N_5208,N_5148);
nand U5372 (N_5372,N_5219,N_5176);
and U5373 (N_5373,N_5191,N_5148);
nand U5374 (N_5374,N_5157,N_5166);
or U5375 (N_5375,N_5121,N_5184);
xnor U5376 (N_5376,N_5187,N_5145);
xnor U5377 (N_5377,N_5177,N_5276);
nor U5378 (N_5378,N_5213,N_5268);
nor U5379 (N_5379,N_5269,N_5151);
xnor U5380 (N_5380,N_5253,N_5227);
nand U5381 (N_5381,N_5212,N_5136);
or U5382 (N_5382,N_5149,N_5167);
or U5383 (N_5383,N_5129,N_5147);
nand U5384 (N_5384,N_5225,N_5202);
nor U5385 (N_5385,N_5121,N_5135);
nor U5386 (N_5386,N_5254,N_5245);
xnor U5387 (N_5387,N_5137,N_5254);
and U5388 (N_5388,N_5159,N_5185);
and U5389 (N_5389,N_5192,N_5254);
xnor U5390 (N_5390,N_5202,N_5226);
or U5391 (N_5391,N_5232,N_5261);
nor U5392 (N_5392,N_5206,N_5236);
and U5393 (N_5393,N_5266,N_5176);
nand U5394 (N_5394,N_5216,N_5212);
xnor U5395 (N_5395,N_5144,N_5162);
and U5396 (N_5396,N_5187,N_5224);
xor U5397 (N_5397,N_5158,N_5148);
or U5398 (N_5398,N_5180,N_5205);
and U5399 (N_5399,N_5123,N_5213);
or U5400 (N_5400,N_5262,N_5244);
nand U5401 (N_5401,N_5220,N_5232);
xor U5402 (N_5402,N_5134,N_5266);
or U5403 (N_5403,N_5172,N_5144);
and U5404 (N_5404,N_5220,N_5223);
or U5405 (N_5405,N_5209,N_5124);
nand U5406 (N_5406,N_5267,N_5223);
or U5407 (N_5407,N_5167,N_5146);
or U5408 (N_5408,N_5262,N_5153);
and U5409 (N_5409,N_5276,N_5231);
or U5410 (N_5410,N_5261,N_5180);
or U5411 (N_5411,N_5136,N_5121);
nor U5412 (N_5412,N_5138,N_5216);
or U5413 (N_5413,N_5182,N_5220);
nor U5414 (N_5414,N_5225,N_5244);
nor U5415 (N_5415,N_5265,N_5174);
nand U5416 (N_5416,N_5176,N_5208);
xnor U5417 (N_5417,N_5176,N_5144);
nor U5418 (N_5418,N_5240,N_5249);
nand U5419 (N_5419,N_5214,N_5188);
and U5420 (N_5420,N_5251,N_5237);
nor U5421 (N_5421,N_5192,N_5228);
nand U5422 (N_5422,N_5250,N_5201);
nor U5423 (N_5423,N_5198,N_5274);
nand U5424 (N_5424,N_5271,N_5152);
and U5425 (N_5425,N_5257,N_5265);
or U5426 (N_5426,N_5211,N_5259);
or U5427 (N_5427,N_5277,N_5124);
and U5428 (N_5428,N_5249,N_5167);
and U5429 (N_5429,N_5255,N_5225);
xor U5430 (N_5430,N_5222,N_5242);
nand U5431 (N_5431,N_5213,N_5223);
xor U5432 (N_5432,N_5160,N_5172);
or U5433 (N_5433,N_5234,N_5235);
nor U5434 (N_5434,N_5125,N_5258);
and U5435 (N_5435,N_5254,N_5216);
xnor U5436 (N_5436,N_5159,N_5256);
xnor U5437 (N_5437,N_5232,N_5176);
nor U5438 (N_5438,N_5238,N_5120);
or U5439 (N_5439,N_5271,N_5227);
xnor U5440 (N_5440,N_5377,N_5376);
nor U5441 (N_5441,N_5292,N_5352);
xnor U5442 (N_5442,N_5382,N_5336);
or U5443 (N_5443,N_5323,N_5430);
xor U5444 (N_5444,N_5318,N_5399);
or U5445 (N_5445,N_5406,N_5414);
and U5446 (N_5446,N_5415,N_5360);
and U5447 (N_5447,N_5299,N_5284);
nor U5448 (N_5448,N_5340,N_5293);
nor U5449 (N_5449,N_5387,N_5413);
or U5450 (N_5450,N_5422,N_5344);
and U5451 (N_5451,N_5427,N_5356);
xnor U5452 (N_5452,N_5313,N_5349);
or U5453 (N_5453,N_5398,N_5353);
and U5454 (N_5454,N_5416,N_5426);
xor U5455 (N_5455,N_5329,N_5290);
and U5456 (N_5456,N_5371,N_5358);
nand U5457 (N_5457,N_5332,N_5306);
nor U5458 (N_5458,N_5404,N_5312);
or U5459 (N_5459,N_5429,N_5319);
nand U5460 (N_5460,N_5378,N_5309);
nand U5461 (N_5461,N_5432,N_5367);
xor U5462 (N_5462,N_5295,N_5384);
nor U5463 (N_5463,N_5433,N_5420);
and U5464 (N_5464,N_5391,N_5408);
nor U5465 (N_5465,N_5390,N_5411);
xor U5466 (N_5466,N_5351,N_5369);
nand U5467 (N_5467,N_5335,N_5316);
or U5468 (N_5468,N_5389,N_5394);
and U5469 (N_5469,N_5421,N_5302);
nor U5470 (N_5470,N_5437,N_5350);
or U5471 (N_5471,N_5438,N_5326);
nor U5472 (N_5472,N_5305,N_5405);
nand U5473 (N_5473,N_5333,N_5343);
xor U5474 (N_5474,N_5310,N_5431);
nand U5475 (N_5475,N_5304,N_5373);
and U5476 (N_5476,N_5403,N_5379);
xor U5477 (N_5477,N_5417,N_5339);
or U5478 (N_5478,N_5386,N_5396);
and U5479 (N_5479,N_5428,N_5372);
nor U5480 (N_5480,N_5357,N_5285);
or U5481 (N_5481,N_5280,N_5400);
and U5482 (N_5482,N_5342,N_5423);
and U5483 (N_5483,N_5324,N_5364);
nor U5484 (N_5484,N_5392,N_5375);
or U5485 (N_5485,N_5380,N_5425);
or U5486 (N_5486,N_5412,N_5348);
nor U5487 (N_5487,N_5393,N_5436);
and U5488 (N_5488,N_5334,N_5419);
xor U5489 (N_5489,N_5322,N_5381);
and U5490 (N_5490,N_5315,N_5365);
xnor U5491 (N_5491,N_5402,N_5338);
and U5492 (N_5492,N_5317,N_5283);
nor U5493 (N_5493,N_5298,N_5355);
nor U5494 (N_5494,N_5409,N_5370);
xnor U5495 (N_5495,N_5300,N_5282);
nor U5496 (N_5496,N_5330,N_5347);
xor U5497 (N_5497,N_5363,N_5286);
and U5498 (N_5498,N_5401,N_5424);
or U5499 (N_5499,N_5374,N_5435);
or U5500 (N_5500,N_5327,N_5311);
xor U5501 (N_5501,N_5368,N_5434);
nor U5502 (N_5502,N_5354,N_5346);
or U5503 (N_5503,N_5395,N_5294);
or U5504 (N_5504,N_5341,N_5325);
and U5505 (N_5505,N_5320,N_5301);
and U5506 (N_5506,N_5418,N_5407);
or U5507 (N_5507,N_5287,N_5291);
or U5508 (N_5508,N_5388,N_5297);
or U5509 (N_5509,N_5359,N_5321);
or U5510 (N_5510,N_5288,N_5383);
or U5511 (N_5511,N_5289,N_5314);
nor U5512 (N_5512,N_5303,N_5331);
nor U5513 (N_5513,N_5366,N_5296);
nor U5514 (N_5514,N_5328,N_5361);
and U5515 (N_5515,N_5281,N_5385);
and U5516 (N_5516,N_5362,N_5410);
and U5517 (N_5517,N_5397,N_5439);
nand U5518 (N_5518,N_5337,N_5345);
xnor U5519 (N_5519,N_5308,N_5307);
xnor U5520 (N_5520,N_5338,N_5306);
or U5521 (N_5521,N_5367,N_5404);
or U5522 (N_5522,N_5406,N_5299);
or U5523 (N_5523,N_5378,N_5284);
nor U5524 (N_5524,N_5408,N_5291);
and U5525 (N_5525,N_5347,N_5432);
nor U5526 (N_5526,N_5394,N_5298);
and U5527 (N_5527,N_5392,N_5287);
nor U5528 (N_5528,N_5438,N_5299);
or U5529 (N_5529,N_5312,N_5336);
nor U5530 (N_5530,N_5286,N_5347);
nor U5531 (N_5531,N_5313,N_5423);
or U5532 (N_5532,N_5428,N_5405);
or U5533 (N_5533,N_5367,N_5386);
or U5534 (N_5534,N_5415,N_5431);
or U5535 (N_5535,N_5367,N_5379);
xnor U5536 (N_5536,N_5285,N_5409);
xor U5537 (N_5537,N_5412,N_5375);
or U5538 (N_5538,N_5435,N_5307);
or U5539 (N_5539,N_5404,N_5348);
and U5540 (N_5540,N_5399,N_5354);
nor U5541 (N_5541,N_5356,N_5380);
xnor U5542 (N_5542,N_5323,N_5366);
and U5543 (N_5543,N_5425,N_5423);
xor U5544 (N_5544,N_5422,N_5373);
nand U5545 (N_5545,N_5430,N_5324);
nor U5546 (N_5546,N_5369,N_5429);
xor U5547 (N_5547,N_5379,N_5292);
nor U5548 (N_5548,N_5419,N_5329);
xnor U5549 (N_5549,N_5340,N_5302);
xor U5550 (N_5550,N_5320,N_5421);
xor U5551 (N_5551,N_5419,N_5406);
and U5552 (N_5552,N_5280,N_5424);
xnor U5553 (N_5553,N_5434,N_5401);
nor U5554 (N_5554,N_5377,N_5429);
or U5555 (N_5555,N_5392,N_5377);
nor U5556 (N_5556,N_5303,N_5290);
xnor U5557 (N_5557,N_5409,N_5385);
xor U5558 (N_5558,N_5339,N_5371);
nor U5559 (N_5559,N_5401,N_5373);
nand U5560 (N_5560,N_5304,N_5380);
or U5561 (N_5561,N_5420,N_5439);
or U5562 (N_5562,N_5402,N_5336);
nor U5563 (N_5563,N_5329,N_5338);
nand U5564 (N_5564,N_5365,N_5359);
or U5565 (N_5565,N_5336,N_5302);
nor U5566 (N_5566,N_5367,N_5336);
or U5567 (N_5567,N_5403,N_5342);
and U5568 (N_5568,N_5320,N_5311);
nor U5569 (N_5569,N_5438,N_5346);
and U5570 (N_5570,N_5347,N_5285);
and U5571 (N_5571,N_5410,N_5409);
nand U5572 (N_5572,N_5413,N_5360);
nand U5573 (N_5573,N_5322,N_5401);
and U5574 (N_5574,N_5401,N_5349);
and U5575 (N_5575,N_5404,N_5298);
xnor U5576 (N_5576,N_5418,N_5322);
xnor U5577 (N_5577,N_5289,N_5368);
and U5578 (N_5578,N_5426,N_5381);
nor U5579 (N_5579,N_5312,N_5403);
xor U5580 (N_5580,N_5300,N_5429);
and U5581 (N_5581,N_5370,N_5431);
nand U5582 (N_5582,N_5370,N_5297);
nand U5583 (N_5583,N_5409,N_5420);
nand U5584 (N_5584,N_5414,N_5438);
nand U5585 (N_5585,N_5364,N_5280);
or U5586 (N_5586,N_5338,N_5419);
xor U5587 (N_5587,N_5349,N_5365);
xnor U5588 (N_5588,N_5319,N_5370);
nor U5589 (N_5589,N_5428,N_5363);
xor U5590 (N_5590,N_5408,N_5359);
nand U5591 (N_5591,N_5283,N_5382);
xor U5592 (N_5592,N_5422,N_5314);
xor U5593 (N_5593,N_5403,N_5294);
or U5594 (N_5594,N_5371,N_5380);
and U5595 (N_5595,N_5315,N_5371);
xnor U5596 (N_5596,N_5320,N_5309);
nor U5597 (N_5597,N_5375,N_5365);
and U5598 (N_5598,N_5352,N_5325);
xnor U5599 (N_5599,N_5352,N_5314);
nand U5600 (N_5600,N_5502,N_5598);
nor U5601 (N_5601,N_5520,N_5448);
xnor U5602 (N_5602,N_5559,N_5585);
nor U5603 (N_5603,N_5569,N_5519);
nand U5604 (N_5604,N_5492,N_5482);
and U5605 (N_5605,N_5484,N_5527);
nor U5606 (N_5606,N_5551,N_5549);
nand U5607 (N_5607,N_5566,N_5550);
xnor U5608 (N_5608,N_5503,N_5583);
and U5609 (N_5609,N_5496,N_5447);
nor U5610 (N_5610,N_5444,N_5465);
xor U5611 (N_5611,N_5534,N_5556);
or U5612 (N_5612,N_5574,N_5446);
and U5613 (N_5613,N_5543,N_5541);
and U5614 (N_5614,N_5572,N_5495);
nor U5615 (N_5615,N_5557,N_5537);
and U5616 (N_5616,N_5562,N_5590);
xor U5617 (N_5617,N_5469,N_5518);
xnor U5618 (N_5618,N_5595,N_5466);
or U5619 (N_5619,N_5599,N_5460);
nor U5620 (N_5620,N_5545,N_5530);
and U5621 (N_5621,N_5544,N_5538);
or U5622 (N_5622,N_5494,N_5515);
or U5623 (N_5623,N_5561,N_5467);
nand U5624 (N_5624,N_5504,N_5594);
xnor U5625 (N_5625,N_5580,N_5476);
nand U5626 (N_5626,N_5506,N_5523);
xnor U5627 (N_5627,N_5485,N_5558);
and U5628 (N_5628,N_5459,N_5463);
or U5629 (N_5629,N_5499,N_5450);
and U5630 (N_5630,N_5440,N_5455);
nor U5631 (N_5631,N_5555,N_5531);
nand U5632 (N_5632,N_5554,N_5470);
nand U5633 (N_5633,N_5449,N_5576);
xnor U5634 (N_5634,N_5490,N_5524);
xor U5635 (N_5635,N_5553,N_5483);
and U5636 (N_5636,N_5567,N_5577);
nand U5637 (N_5637,N_5517,N_5468);
and U5638 (N_5638,N_5587,N_5453);
and U5639 (N_5639,N_5479,N_5474);
and U5640 (N_5640,N_5575,N_5451);
nand U5641 (N_5641,N_5548,N_5510);
and U5642 (N_5642,N_5563,N_5570);
nor U5643 (N_5643,N_5597,N_5445);
or U5644 (N_5644,N_5475,N_5591);
and U5645 (N_5645,N_5441,N_5462);
nor U5646 (N_5646,N_5489,N_5452);
nor U5647 (N_5647,N_5526,N_5525);
or U5648 (N_5648,N_5500,N_5501);
or U5649 (N_5649,N_5579,N_5514);
and U5650 (N_5650,N_5592,N_5471);
nand U5651 (N_5651,N_5578,N_5454);
nand U5652 (N_5652,N_5593,N_5505);
and U5653 (N_5653,N_5513,N_5461);
nand U5654 (N_5654,N_5532,N_5443);
and U5655 (N_5655,N_5582,N_5472);
or U5656 (N_5656,N_5539,N_5509);
and U5657 (N_5657,N_5457,N_5552);
nor U5658 (N_5658,N_5491,N_5568);
and U5659 (N_5659,N_5464,N_5581);
or U5660 (N_5660,N_5564,N_5486);
and U5661 (N_5661,N_5511,N_5589);
or U5662 (N_5662,N_5507,N_5529);
nand U5663 (N_5663,N_5473,N_5481);
xor U5664 (N_5664,N_5498,N_5586);
or U5665 (N_5665,N_5560,N_5508);
nand U5666 (N_5666,N_5458,N_5477);
nor U5667 (N_5667,N_5540,N_5528);
xor U5668 (N_5668,N_5596,N_5521);
and U5669 (N_5669,N_5480,N_5536);
nor U5670 (N_5670,N_5456,N_5478);
xor U5671 (N_5671,N_5493,N_5512);
nand U5672 (N_5672,N_5497,N_5565);
or U5673 (N_5673,N_5584,N_5588);
and U5674 (N_5674,N_5535,N_5488);
xor U5675 (N_5675,N_5542,N_5522);
xnor U5676 (N_5676,N_5533,N_5571);
or U5677 (N_5677,N_5547,N_5546);
xor U5678 (N_5678,N_5442,N_5487);
or U5679 (N_5679,N_5573,N_5516);
or U5680 (N_5680,N_5599,N_5536);
nand U5681 (N_5681,N_5476,N_5523);
xor U5682 (N_5682,N_5572,N_5579);
or U5683 (N_5683,N_5520,N_5546);
nand U5684 (N_5684,N_5571,N_5540);
nand U5685 (N_5685,N_5566,N_5453);
nand U5686 (N_5686,N_5497,N_5577);
nor U5687 (N_5687,N_5502,N_5496);
nand U5688 (N_5688,N_5545,N_5544);
or U5689 (N_5689,N_5529,N_5564);
xnor U5690 (N_5690,N_5592,N_5554);
nor U5691 (N_5691,N_5505,N_5571);
nor U5692 (N_5692,N_5465,N_5560);
xnor U5693 (N_5693,N_5535,N_5514);
xnor U5694 (N_5694,N_5444,N_5592);
nand U5695 (N_5695,N_5549,N_5593);
xnor U5696 (N_5696,N_5527,N_5556);
and U5697 (N_5697,N_5514,N_5552);
nor U5698 (N_5698,N_5506,N_5590);
and U5699 (N_5699,N_5445,N_5543);
nand U5700 (N_5700,N_5515,N_5486);
nand U5701 (N_5701,N_5490,N_5554);
nand U5702 (N_5702,N_5481,N_5445);
or U5703 (N_5703,N_5495,N_5449);
nor U5704 (N_5704,N_5445,N_5498);
nand U5705 (N_5705,N_5447,N_5511);
or U5706 (N_5706,N_5464,N_5486);
nor U5707 (N_5707,N_5476,N_5518);
xor U5708 (N_5708,N_5508,N_5577);
nand U5709 (N_5709,N_5507,N_5586);
and U5710 (N_5710,N_5446,N_5505);
xnor U5711 (N_5711,N_5501,N_5555);
xor U5712 (N_5712,N_5447,N_5553);
nor U5713 (N_5713,N_5475,N_5469);
and U5714 (N_5714,N_5572,N_5570);
nand U5715 (N_5715,N_5560,N_5589);
or U5716 (N_5716,N_5465,N_5593);
and U5717 (N_5717,N_5512,N_5513);
and U5718 (N_5718,N_5577,N_5571);
or U5719 (N_5719,N_5470,N_5566);
nor U5720 (N_5720,N_5491,N_5482);
or U5721 (N_5721,N_5570,N_5448);
nand U5722 (N_5722,N_5589,N_5528);
nor U5723 (N_5723,N_5501,N_5489);
or U5724 (N_5724,N_5502,N_5508);
nor U5725 (N_5725,N_5487,N_5482);
xnor U5726 (N_5726,N_5459,N_5515);
and U5727 (N_5727,N_5534,N_5560);
nand U5728 (N_5728,N_5550,N_5560);
nand U5729 (N_5729,N_5531,N_5536);
and U5730 (N_5730,N_5547,N_5496);
xnor U5731 (N_5731,N_5467,N_5495);
xnor U5732 (N_5732,N_5517,N_5483);
nor U5733 (N_5733,N_5572,N_5466);
and U5734 (N_5734,N_5568,N_5511);
nand U5735 (N_5735,N_5450,N_5463);
or U5736 (N_5736,N_5463,N_5471);
nand U5737 (N_5737,N_5555,N_5445);
or U5738 (N_5738,N_5540,N_5585);
or U5739 (N_5739,N_5557,N_5594);
nand U5740 (N_5740,N_5598,N_5451);
xor U5741 (N_5741,N_5483,N_5464);
or U5742 (N_5742,N_5568,N_5579);
or U5743 (N_5743,N_5486,N_5552);
or U5744 (N_5744,N_5553,N_5498);
xor U5745 (N_5745,N_5516,N_5473);
and U5746 (N_5746,N_5442,N_5580);
and U5747 (N_5747,N_5575,N_5526);
xor U5748 (N_5748,N_5556,N_5586);
or U5749 (N_5749,N_5535,N_5532);
xnor U5750 (N_5750,N_5561,N_5440);
xnor U5751 (N_5751,N_5586,N_5598);
or U5752 (N_5752,N_5552,N_5574);
and U5753 (N_5753,N_5465,N_5509);
nor U5754 (N_5754,N_5458,N_5555);
nor U5755 (N_5755,N_5490,N_5566);
nand U5756 (N_5756,N_5589,N_5580);
xnor U5757 (N_5757,N_5463,N_5588);
xnor U5758 (N_5758,N_5586,N_5447);
nand U5759 (N_5759,N_5511,N_5506);
nand U5760 (N_5760,N_5656,N_5757);
or U5761 (N_5761,N_5715,N_5736);
or U5762 (N_5762,N_5627,N_5735);
nor U5763 (N_5763,N_5745,N_5658);
and U5764 (N_5764,N_5665,N_5640);
or U5765 (N_5765,N_5685,N_5604);
or U5766 (N_5766,N_5648,N_5631);
and U5767 (N_5767,N_5605,N_5706);
xnor U5768 (N_5768,N_5726,N_5678);
nand U5769 (N_5769,N_5663,N_5701);
nand U5770 (N_5770,N_5750,N_5689);
nand U5771 (N_5771,N_5661,N_5672);
and U5772 (N_5772,N_5638,N_5655);
nor U5773 (N_5773,N_5653,N_5606);
xor U5774 (N_5774,N_5700,N_5718);
nor U5775 (N_5775,N_5660,N_5751);
nand U5776 (N_5776,N_5617,N_5623);
nand U5777 (N_5777,N_5740,N_5633);
nand U5778 (N_5778,N_5729,N_5723);
or U5779 (N_5779,N_5666,N_5668);
or U5780 (N_5780,N_5727,N_5612);
and U5781 (N_5781,N_5744,N_5710);
nor U5782 (N_5782,N_5704,N_5622);
nor U5783 (N_5783,N_5650,N_5637);
xor U5784 (N_5784,N_5691,N_5688);
xor U5785 (N_5785,N_5636,N_5624);
or U5786 (N_5786,N_5614,N_5755);
xnor U5787 (N_5787,N_5670,N_5674);
or U5788 (N_5788,N_5708,N_5748);
or U5789 (N_5789,N_5680,N_5702);
nand U5790 (N_5790,N_5707,N_5692);
xnor U5791 (N_5791,N_5616,N_5669);
and U5792 (N_5792,N_5644,N_5676);
and U5793 (N_5793,N_5603,N_5758);
and U5794 (N_5794,N_5737,N_5721);
xor U5795 (N_5795,N_5709,N_5630);
and U5796 (N_5796,N_5643,N_5652);
xor U5797 (N_5797,N_5716,N_5693);
or U5798 (N_5798,N_5724,N_5645);
xnor U5799 (N_5799,N_5618,N_5635);
and U5800 (N_5800,N_5742,N_5690);
nand U5801 (N_5801,N_5732,N_5639);
or U5802 (N_5802,N_5681,N_5615);
nand U5803 (N_5803,N_5620,N_5684);
and U5804 (N_5804,N_5728,N_5659);
nor U5805 (N_5805,N_5698,N_5647);
and U5806 (N_5806,N_5642,N_5632);
or U5807 (N_5807,N_5646,N_5696);
nor U5808 (N_5808,N_5613,N_5601);
xor U5809 (N_5809,N_5720,N_5714);
xor U5810 (N_5810,N_5654,N_5675);
nand U5811 (N_5811,N_5753,N_5625);
xnor U5812 (N_5812,N_5686,N_5600);
and U5813 (N_5813,N_5621,N_5722);
nand U5814 (N_5814,N_5711,N_5743);
and U5815 (N_5815,N_5741,N_5739);
nor U5816 (N_5816,N_5756,N_5667);
xor U5817 (N_5817,N_5607,N_5759);
nor U5818 (N_5818,N_5602,N_5731);
and U5819 (N_5819,N_5611,N_5609);
and U5820 (N_5820,N_5629,N_5664);
xnor U5821 (N_5821,N_5717,N_5677);
or U5822 (N_5822,N_5628,N_5682);
nor U5823 (N_5823,N_5752,N_5705);
and U5824 (N_5824,N_5671,N_5754);
xor U5825 (N_5825,N_5730,N_5694);
and U5826 (N_5826,N_5713,N_5734);
nor U5827 (N_5827,N_5651,N_5687);
or U5828 (N_5828,N_5697,N_5733);
or U5829 (N_5829,N_5610,N_5738);
nor U5830 (N_5830,N_5608,N_5699);
and U5831 (N_5831,N_5746,N_5649);
xnor U5832 (N_5832,N_5747,N_5619);
xnor U5833 (N_5833,N_5695,N_5725);
nand U5834 (N_5834,N_5719,N_5712);
nor U5835 (N_5835,N_5673,N_5703);
xnor U5836 (N_5836,N_5683,N_5662);
xor U5837 (N_5837,N_5679,N_5641);
and U5838 (N_5838,N_5749,N_5626);
or U5839 (N_5839,N_5657,N_5634);
and U5840 (N_5840,N_5666,N_5721);
nand U5841 (N_5841,N_5688,N_5613);
xor U5842 (N_5842,N_5644,N_5754);
and U5843 (N_5843,N_5739,N_5628);
xor U5844 (N_5844,N_5661,N_5677);
or U5845 (N_5845,N_5628,N_5622);
and U5846 (N_5846,N_5654,N_5679);
and U5847 (N_5847,N_5746,N_5729);
nand U5848 (N_5848,N_5638,N_5729);
and U5849 (N_5849,N_5649,N_5715);
or U5850 (N_5850,N_5744,N_5749);
nand U5851 (N_5851,N_5702,N_5699);
nand U5852 (N_5852,N_5746,N_5739);
xnor U5853 (N_5853,N_5742,N_5665);
xnor U5854 (N_5854,N_5748,N_5703);
xnor U5855 (N_5855,N_5622,N_5735);
xnor U5856 (N_5856,N_5627,N_5729);
nand U5857 (N_5857,N_5661,N_5714);
nand U5858 (N_5858,N_5682,N_5617);
nor U5859 (N_5859,N_5685,N_5719);
nor U5860 (N_5860,N_5723,N_5674);
and U5861 (N_5861,N_5688,N_5643);
nand U5862 (N_5862,N_5753,N_5689);
or U5863 (N_5863,N_5623,N_5625);
nand U5864 (N_5864,N_5696,N_5729);
nor U5865 (N_5865,N_5638,N_5619);
nor U5866 (N_5866,N_5711,N_5650);
nor U5867 (N_5867,N_5650,N_5698);
nor U5868 (N_5868,N_5719,N_5737);
xnor U5869 (N_5869,N_5733,N_5683);
or U5870 (N_5870,N_5658,N_5673);
nand U5871 (N_5871,N_5685,N_5740);
nand U5872 (N_5872,N_5759,N_5747);
nor U5873 (N_5873,N_5753,N_5614);
xor U5874 (N_5874,N_5674,N_5672);
or U5875 (N_5875,N_5630,N_5631);
or U5876 (N_5876,N_5655,N_5688);
or U5877 (N_5877,N_5680,N_5618);
nor U5878 (N_5878,N_5678,N_5723);
xor U5879 (N_5879,N_5640,N_5635);
and U5880 (N_5880,N_5742,N_5679);
xnor U5881 (N_5881,N_5727,N_5749);
nand U5882 (N_5882,N_5670,N_5726);
xor U5883 (N_5883,N_5704,N_5669);
nor U5884 (N_5884,N_5720,N_5754);
nand U5885 (N_5885,N_5624,N_5661);
nand U5886 (N_5886,N_5614,N_5746);
nor U5887 (N_5887,N_5623,N_5658);
and U5888 (N_5888,N_5689,N_5608);
nand U5889 (N_5889,N_5689,N_5620);
and U5890 (N_5890,N_5722,N_5758);
nand U5891 (N_5891,N_5657,N_5610);
nor U5892 (N_5892,N_5727,N_5705);
and U5893 (N_5893,N_5744,N_5649);
or U5894 (N_5894,N_5748,N_5607);
xnor U5895 (N_5895,N_5635,N_5676);
or U5896 (N_5896,N_5703,N_5749);
or U5897 (N_5897,N_5688,N_5730);
and U5898 (N_5898,N_5631,N_5747);
or U5899 (N_5899,N_5694,N_5754);
or U5900 (N_5900,N_5666,N_5686);
or U5901 (N_5901,N_5665,N_5685);
or U5902 (N_5902,N_5617,N_5711);
and U5903 (N_5903,N_5670,N_5695);
and U5904 (N_5904,N_5664,N_5634);
or U5905 (N_5905,N_5711,N_5611);
nor U5906 (N_5906,N_5671,N_5642);
xor U5907 (N_5907,N_5724,N_5703);
or U5908 (N_5908,N_5635,N_5751);
xnor U5909 (N_5909,N_5695,N_5635);
nor U5910 (N_5910,N_5708,N_5610);
or U5911 (N_5911,N_5710,N_5685);
and U5912 (N_5912,N_5701,N_5620);
nor U5913 (N_5913,N_5723,N_5719);
nand U5914 (N_5914,N_5617,N_5665);
xor U5915 (N_5915,N_5619,N_5681);
nor U5916 (N_5916,N_5708,N_5613);
nand U5917 (N_5917,N_5661,N_5692);
nand U5918 (N_5918,N_5695,N_5619);
and U5919 (N_5919,N_5692,N_5664);
nand U5920 (N_5920,N_5879,N_5810);
xor U5921 (N_5921,N_5910,N_5793);
nand U5922 (N_5922,N_5892,N_5838);
and U5923 (N_5923,N_5916,N_5884);
xnor U5924 (N_5924,N_5893,N_5874);
nand U5925 (N_5925,N_5829,N_5780);
nor U5926 (N_5926,N_5881,N_5882);
xor U5927 (N_5927,N_5913,N_5886);
nor U5928 (N_5928,N_5836,N_5767);
xnor U5929 (N_5929,N_5773,N_5908);
nand U5930 (N_5930,N_5912,N_5860);
nand U5931 (N_5931,N_5903,N_5788);
and U5932 (N_5932,N_5777,N_5847);
or U5933 (N_5933,N_5854,N_5863);
nand U5934 (N_5934,N_5848,N_5868);
or U5935 (N_5935,N_5877,N_5831);
xnor U5936 (N_5936,N_5891,N_5785);
nor U5937 (N_5937,N_5878,N_5887);
and U5938 (N_5938,N_5872,N_5808);
nor U5939 (N_5939,N_5915,N_5858);
nand U5940 (N_5940,N_5842,N_5799);
and U5941 (N_5941,N_5862,N_5800);
nor U5942 (N_5942,N_5781,N_5770);
nand U5943 (N_5943,N_5864,N_5883);
and U5944 (N_5944,N_5827,N_5784);
xor U5945 (N_5945,N_5904,N_5821);
and U5946 (N_5946,N_5789,N_5859);
and U5947 (N_5947,N_5762,N_5824);
and U5948 (N_5948,N_5814,N_5772);
or U5949 (N_5949,N_5764,N_5801);
nor U5950 (N_5950,N_5811,N_5841);
and U5951 (N_5951,N_5797,N_5790);
nand U5952 (N_5952,N_5898,N_5825);
nand U5953 (N_5953,N_5798,N_5866);
xor U5954 (N_5954,N_5765,N_5917);
and U5955 (N_5955,N_5919,N_5771);
and U5956 (N_5956,N_5806,N_5876);
nand U5957 (N_5957,N_5865,N_5769);
and U5958 (N_5958,N_5817,N_5786);
nor U5959 (N_5959,N_5796,N_5783);
nand U5960 (N_5960,N_5766,N_5795);
and U5961 (N_5961,N_5867,N_5901);
nand U5962 (N_5962,N_5914,N_5844);
xor U5963 (N_5963,N_5816,N_5835);
nand U5964 (N_5964,N_5779,N_5778);
nor U5965 (N_5965,N_5822,N_5819);
and U5966 (N_5966,N_5846,N_5907);
xor U5967 (N_5967,N_5871,N_5776);
and U5968 (N_5968,N_5826,N_5902);
nand U5969 (N_5969,N_5852,N_5894);
or U5970 (N_5970,N_5760,N_5861);
or U5971 (N_5971,N_5813,N_5889);
nand U5972 (N_5972,N_5787,N_5794);
nand U5973 (N_5973,N_5807,N_5791);
or U5974 (N_5974,N_5820,N_5890);
and U5975 (N_5975,N_5763,N_5888);
nand U5976 (N_5976,N_5873,N_5849);
or U5977 (N_5977,N_5775,N_5856);
and U5978 (N_5978,N_5896,N_5815);
nor U5979 (N_5979,N_5875,N_5828);
xnor U5980 (N_5980,N_5774,N_5768);
nor U5981 (N_5981,N_5918,N_5900);
or U5982 (N_5982,N_5851,N_5833);
and U5983 (N_5983,N_5830,N_5895);
and U5984 (N_5984,N_5834,N_5761);
nor U5985 (N_5985,N_5869,N_5839);
and U5986 (N_5986,N_5899,N_5906);
nor U5987 (N_5987,N_5880,N_5805);
or U5988 (N_5988,N_5857,N_5853);
nor U5989 (N_5989,N_5905,N_5845);
and U5990 (N_5990,N_5809,N_5782);
xnor U5991 (N_5991,N_5802,N_5885);
or U5992 (N_5992,N_5897,N_5792);
or U5993 (N_5993,N_5909,N_5850);
nand U5994 (N_5994,N_5843,N_5804);
or U5995 (N_5995,N_5837,N_5812);
nor U5996 (N_5996,N_5803,N_5823);
nand U5997 (N_5997,N_5840,N_5855);
or U5998 (N_5998,N_5911,N_5870);
nor U5999 (N_5999,N_5818,N_5832);
nor U6000 (N_6000,N_5768,N_5804);
nor U6001 (N_6001,N_5801,N_5860);
nand U6002 (N_6002,N_5794,N_5824);
nand U6003 (N_6003,N_5803,N_5918);
or U6004 (N_6004,N_5818,N_5839);
and U6005 (N_6005,N_5879,N_5869);
and U6006 (N_6006,N_5769,N_5810);
or U6007 (N_6007,N_5777,N_5868);
xnor U6008 (N_6008,N_5907,N_5792);
nor U6009 (N_6009,N_5892,N_5894);
nor U6010 (N_6010,N_5863,N_5861);
nand U6011 (N_6011,N_5779,N_5918);
nor U6012 (N_6012,N_5910,N_5895);
and U6013 (N_6013,N_5835,N_5802);
nor U6014 (N_6014,N_5872,N_5864);
nand U6015 (N_6015,N_5889,N_5771);
xnor U6016 (N_6016,N_5812,N_5806);
xnor U6017 (N_6017,N_5802,N_5773);
nor U6018 (N_6018,N_5911,N_5851);
and U6019 (N_6019,N_5871,N_5804);
and U6020 (N_6020,N_5761,N_5774);
xnor U6021 (N_6021,N_5902,N_5885);
xor U6022 (N_6022,N_5805,N_5905);
nand U6023 (N_6023,N_5881,N_5769);
or U6024 (N_6024,N_5845,N_5794);
or U6025 (N_6025,N_5841,N_5889);
or U6026 (N_6026,N_5835,N_5807);
nor U6027 (N_6027,N_5801,N_5895);
xnor U6028 (N_6028,N_5907,N_5814);
or U6029 (N_6029,N_5840,N_5884);
nand U6030 (N_6030,N_5901,N_5887);
nand U6031 (N_6031,N_5774,N_5846);
nand U6032 (N_6032,N_5910,N_5787);
and U6033 (N_6033,N_5888,N_5825);
nand U6034 (N_6034,N_5916,N_5855);
nor U6035 (N_6035,N_5867,N_5834);
xor U6036 (N_6036,N_5764,N_5789);
xor U6037 (N_6037,N_5781,N_5810);
or U6038 (N_6038,N_5841,N_5885);
and U6039 (N_6039,N_5769,N_5875);
nor U6040 (N_6040,N_5830,N_5768);
or U6041 (N_6041,N_5785,N_5893);
or U6042 (N_6042,N_5766,N_5880);
nand U6043 (N_6043,N_5906,N_5771);
and U6044 (N_6044,N_5871,N_5766);
or U6045 (N_6045,N_5809,N_5781);
nor U6046 (N_6046,N_5837,N_5891);
or U6047 (N_6047,N_5785,N_5861);
nand U6048 (N_6048,N_5856,N_5763);
nand U6049 (N_6049,N_5902,N_5898);
or U6050 (N_6050,N_5799,N_5762);
xnor U6051 (N_6051,N_5774,N_5835);
nor U6052 (N_6052,N_5811,N_5866);
xnor U6053 (N_6053,N_5889,N_5897);
nor U6054 (N_6054,N_5783,N_5906);
or U6055 (N_6055,N_5911,N_5876);
or U6056 (N_6056,N_5859,N_5779);
nand U6057 (N_6057,N_5871,N_5792);
nand U6058 (N_6058,N_5807,N_5788);
or U6059 (N_6059,N_5909,N_5885);
and U6060 (N_6060,N_5804,N_5838);
and U6061 (N_6061,N_5879,N_5895);
nor U6062 (N_6062,N_5773,N_5845);
nand U6063 (N_6063,N_5775,N_5919);
nand U6064 (N_6064,N_5833,N_5856);
or U6065 (N_6065,N_5902,N_5899);
nor U6066 (N_6066,N_5909,N_5838);
xnor U6067 (N_6067,N_5877,N_5839);
or U6068 (N_6068,N_5849,N_5813);
nand U6069 (N_6069,N_5776,N_5884);
nand U6070 (N_6070,N_5911,N_5853);
or U6071 (N_6071,N_5789,N_5809);
or U6072 (N_6072,N_5766,N_5862);
xnor U6073 (N_6073,N_5897,N_5838);
nand U6074 (N_6074,N_5860,N_5889);
nand U6075 (N_6075,N_5883,N_5855);
xnor U6076 (N_6076,N_5857,N_5900);
or U6077 (N_6077,N_5862,N_5914);
nor U6078 (N_6078,N_5866,N_5768);
and U6079 (N_6079,N_5898,N_5840);
nand U6080 (N_6080,N_6066,N_5924);
nand U6081 (N_6081,N_6019,N_6047);
and U6082 (N_6082,N_5923,N_5955);
xnor U6083 (N_6083,N_6006,N_6029);
nand U6084 (N_6084,N_5952,N_6031);
or U6085 (N_6085,N_6008,N_6002);
nand U6086 (N_6086,N_5942,N_6035);
and U6087 (N_6087,N_5966,N_5983);
xnor U6088 (N_6088,N_5929,N_5953);
xnor U6089 (N_6089,N_5957,N_6076);
or U6090 (N_6090,N_5936,N_5943);
nor U6091 (N_6091,N_5945,N_6062);
or U6092 (N_6092,N_5980,N_5947);
xnor U6093 (N_6093,N_5928,N_5938);
nor U6094 (N_6094,N_5988,N_5963);
and U6095 (N_6095,N_6053,N_6042);
nand U6096 (N_6096,N_6070,N_6048);
xor U6097 (N_6097,N_6056,N_6072);
nor U6098 (N_6098,N_5939,N_6038);
or U6099 (N_6099,N_5971,N_5981);
nor U6100 (N_6100,N_6028,N_6030);
or U6101 (N_6101,N_6025,N_6049);
or U6102 (N_6102,N_5997,N_5930);
or U6103 (N_6103,N_5964,N_6014);
and U6104 (N_6104,N_6052,N_6010);
nor U6105 (N_6105,N_6011,N_5990);
and U6106 (N_6106,N_5979,N_5986);
and U6107 (N_6107,N_6020,N_6055);
xor U6108 (N_6108,N_5933,N_5992);
and U6109 (N_6109,N_5999,N_5973);
xnor U6110 (N_6110,N_5991,N_6051);
or U6111 (N_6111,N_6009,N_5941);
xnor U6112 (N_6112,N_6057,N_5984);
and U6113 (N_6113,N_6043,N_5968);
xnor U6114 (N_6114,N_6067,N_6024);
or U6115 (N_6115,N_6060,N_6039);
or U6116 (N_6116,N_6041,N_5934);
and U6117 (N_6117,N_6022,N_6075);
xnor U6118 (N_6118,N_6071,N_5921);
nand U6119 (N_6119,N_6078,N_5927);
xnor U6120 (N_6120,N_5969,N_5949);
and U6121 (N_6121,N_5967,N_5994);
nand U6122 (N_6122,N_6027,N_6018);
and U6123 (N_6123,N_5978,N_6044);
nand U6124 (N_6124,N_6058,N_6017);
and U6125 (N_6125,N_6037,N_5993);
or U6126 (N_6126,N_6004,N_5975);
xor U6127 (N_6127,N_5970,N_5935);
and U6128 (N_6128,N_6003,N_5972);
and U6129 (N_6129,N_5977,N_5922);
nor U6130 (N_6130,N_6033,N_6034);
or U6131 (N_6131,N_6073,N_5925);
nor U6132 (N_6132,N_6069,N_6061);
nand U6133 (N_6133,N_6005,N_5926);
or U6134 (N_6134,N_5962,N_6013);
or U6135 (N_6135,N_5958,N_6077);
nand U6136 (N_6136,N_6016,N_5931);
nor U6137 (N_6137,N_6045,N_5996);
and U6138 (N_6138,N_6000,N_5951);
nor U6139 (N_6139,N_5976,N_5954);
nor U6140 (N_6140,N_6026,N_5946);
or U6141 (N_6141,N_6001,N_5920);
nand U6142 (N_6142,N_5932,N_5960);
or U6143 (N_6143,N_5956,N_6063);
and U6144 (N_6144,N_5937,N_6015);
and U6145 (N_6145,N_6074,N_6007);
and U6146 (N_6146,N_5995,N_6012);
and U6147 (N_6147,N_6050,N_6036);
or U6148 (N_6148,N_5987,N_6064);
nand U6149 (N_6149,N_5998,N_5965);
nand U6150 (N_6150,N_6040,N_6068);
xnor U6151 (N_6151,N_5944,N_5985);
xnor U6152 (N_6152,N_5950,N_6021);
and U6153 (N_6153,N_5982,N_6054);
nor U6154 (N_6154,N_5974,N_6023);
and U6155 (N_6155,N_5948,N_5989);
xor U6156 (N_6156,N_6032,N_6046);
or U6157 (N_6157,N_6059,N_5959);
or U6158 (N_6158,N_5940,N_6065);
or U6159 (N_6159,N_6079,N_5961);
or U6160 (N_6160,N_6049,N_5987);
or U6161 (N_6161,N_5987,N_6030);
nor U6162 (N_6162,N_6036,N_5972);
xnor U6163 (N_6163,N_5935,N_6006);
xor U6164 (N_6164,N_5991,N_5934);
and U6165 (N_6165,N_5983,N_6059);
xnor U6166 (N_6166,N_6053,N_5936);
nor U6167 (N_6167,N_5960,N_6070);
or U6168 (N_6168,N_5956,N_5994);
nor U6169 (N_6169,N_5943,N_5970);
nor U6170 (N_6170,N_5955,N_6079);
and U6171 (N_6171,N_5940,N_6030);
nor U6172 (N_6172,N_5943,N_6052);
or U6173 (N_6173,N_5921,N_5997);
nor U6174 (N_6174,N_6071,N_5957);
or U6175 (N_6175,N_5959,N_5970);
nand U6176 (N_6176,N_6067,N_5948);
nand U6177 (N_6177,N_6043,N_6025);
xnor U6178 (N_6178,N_5962,N_6022);
nor U6179 (N_6179,N_5937,N_6016);
nor U6180 (N_6180,N_6045,N_5993);
nor U6181 (N_6181,N_6056,N_5996);
or U6182 (N_6182,N_6054,N_6047);
xnor U6183 (N_6183,N_6040,N_5990);
xor U6184 (N_6184,N_6073,N_5984);
and U6185 (N_6185,N_6060,N_6014);
nand U6186 (N_6186,N_5928,N_5952);
or U6187 (N_6187,N_5939,N_5941);
xnor U6188 (N_6188,N_5934,N_5964);
or U6189 (N_6189,N_5953,N_5967);
and U6190 (N_6190,N_6025,N_5956);
or U6191 (N_6191,N_6062,N_6032);
and U6192 (N_6192,N_5950,N_6079);
xor U6193 (N_6193,N_6033,N_5988);
nand U6194 (N_6194,N_5956,N_5958);
nand U6195 (N_6195,N_5922,N_5960);
xor U6196 (N_6196,N_5979,N_5981);
nand U6197 (N_6197,N_5958,N_6027);
nor U6198 (N_6198,N_6026,N_5967);
nand U6199 (N_6199,N_5954,N_6025);
or U6200 (N_6200,N_6000,N_6041);
or U6201 (N_6201,N_5926,N_5931);
or U6202 (N_6202,N_5930,N_6042);
and U6203 (N_6203,N_5990,N_6007);
xnor U6204 (N_6204,N_5947,N_5982);
and U6205 (N_6205,N_6028,N_6018);
nand U6206 (N_6206,N_6012,N_6009);
or U6207 (N_6207,N_6046,N_6076);
nand U6208 (N_6208,N_5974,N_6022);
nor U6209 (N_6209,N_6015,N_5947);
and U6210 (N_6210,N_6015,N_6067);
xor U6211 (N_6211,N_6046,N_5927);
or U6212 (N_6212,N_5972,N_5992);
nand U6213 (N_6213,N_5960,N_5936);
nor U6214 (N_6214,N_6075,N_5995);
nand U6215 (N_6215,N_5969,N_6026);
or U6216 (N_6216,N_6035,N_5933);
or U6217 (N_6217,N_5958,N_5959);
xnor U6218 (N_6218,N_6056,N_6079);
nand U6219 (N_6219,N_5982,N_6061);
or U6220 (N_6220,N_5923,N_6034);
and U6221 (N_6221,N_5979,N_6039);
or U6222 (N_6222,N_5954,N_5923);
nand U6223 (N_6223,N_6006,N_5923);
xnor U6224 (N_6224,N_5991,N_6022);
or U6225 (N_6225,N_6013,N_6065);
and U6226 (N_6226,N_5941,N_5994);
or U6227 (N_6227,N_6073,N_6033);
or U6228 (N_6228,N_5991,N_5949);
nand U6229 (N_6229,N_5921,N_5923);
xnor U6230 (N_6230,N_5937,N_6021);
xnor U6231 (N_6231,N_5940,N_6015);
nor U6232 (N_6232,N_6022,N_5944);
and U6233 (N_6233,N_6070,N_5930);
nand U6234 (N_6234,N_6073,N_6029);
nor U6235 (N_6235,N_6028,N_6017);
nor U6236 (N_6236,N_6078,N_5986);
nor U6237 (N_6237,N_6072,N_5934);
and U6238 (N_6238,N_5969,N_6005);
xnor U6239 (N_6239,N_6023,N_6014);
and U6240 (N_6240,N_6173,N_6146);
xnor U6241 (N_6241,N_6231,N_6147);
nand U6242 (N_6242,N_6167,N_6083);
nor U6243 (N_6243,N_6103,N_6131);
xnor U6244 (N_6244,N_6104,N_6117);
or U6245 (N_6245,N_6148,N_6157);
nand U6246 (N_6246,N_6215,N_6156);
or U6247 (N_6247,N_6208,N_6188);
xor U6248 (N_6248,N_6097,N_6094);
nand U6249 (N_6249,N_6153,N_6114);
nand U6250 (N_6250,N_6149,N_6119);
and U6251 (N_6251,N_6154,N_6120);
nor U6252 (N_6252,N_6162,N_6144);
or U6253 (N_6253,N_6199,N_6232);
or U6254 (N_6254,N_6093,N_6150);
or U6255 (N_6255,N_6102,N_6080);
and U6256 (N_6256,N_6181,N_6155);
nand U6257 (N_6257,N_6115,N_6234);
nand U6258 (N_6258,N_6122,N_6211);
and U6259 (N_6259,N_6163,N_6192);
nor U6260 (N_6260,N_6207,N_6107);
nand U6261 (N_6261,N_6229,N_6137);
nand U6262 (N_6262,N_6227,N_6233);
and U6263 (N_6263,N_6218,N_6121);
xnor U6264 (N_6264,N_6223,N_6179);
nand U6265 (N_6265,N_6186,N_6221);
and U6266 (N_6266,N_6089,N_6197);
or U6267 (N_6267,N_6101,N_6140);
xor U6268 (N_6268,N_6110,N_6217);
nand U6269 (N_6269,N_6184,N_6098);
and U6270 (N_6270,N_6081,N_6171);
xor U6271 (N_6271,N_6185,N_6202);
xnor U6272 (N_6272,N_6213,N_6168);
and U6273 (N_6273,N_6151,N_6203);
and U6274 (N_6274,N_6092,N_6205);
and U6275 (N_6275,N_6135,N_6105);
or U6276 (N_6276,N_6164,N_6193);
or U6277 (N_6277,N_6142,N_6145);
nand U6278 (N_6278,N_6198,N_6224);
nor U6279 (N_6279,N_6169,N_6176);
nand U6280 (N_6280,N_6165,N_6230);
xnor U6281 (N_6281,N_6143,N_6087);
nor U6282 (N_6282,N_6138,N_6136);
or U6283 (N_6283,N_6123,N_6200);
nand U6284 (N_6284,N_6161,N_6100);
and U6285 (N_6285,N_6096,N_6177);
xor U6286 (N_6286,N_6191,N_6216);
or U6287 (N_6287,N_6174,N_6084);
nand U6288 (N_6288,N_6095,N_6201);
nor U6289 (N_6289,N_6133,N_6139);
or U6290 (N_6290,N_6228,N_6159);
xor U6291 (N_6291,N_6111,N_6222);
xnor U6292 (N_6292,N_6112,N_6226);
or U6293 (N_6293,N_6116,N_6109);
and U6294 (N_6294,N_6196,N_6190);
or U6295 (N_6295,N_6210,N_6175);
nand U6296 (N_6296,N_6099,N_6158);
nor U6297 (N_6297,N_6219,N_6209);
and U6298 (N_6298,N_6206,N_6178);
or U6299 (N_6299,N_6127,N_6172);
nor U6300 (N_6300,N_6214,N_6130);
or U6301 (N_6301,N_6183,N_6189);
and U6302 (N_6302,N_6086,N_6195);
and U6303 (N_6303,N_6090,N_6091);
xor U6304 (N_6304,N_6082,N_6239);
or U6305 (N_6305,N_6182,N_6106);
or U6306 (N_6306,N_6141,N_6237);
nor U6307 (N_6307,N_6220,N_6236);
and U6308 (N_6308,N_6118,N_6204);
or U6309 (N_6309,N_6128,N_6160);
or U6310 (N_6310,N_6113,N_6124);
or U6311 (N_6311,N_6225,N_6152);
nor U6312 (N_6312,N_6108,N_6129);
or U6313 (N_6313,N_6194,N_6132);
and U6314 (N_6314,N_6170,N_6134);
xnor U6315 (N_6315,N_6180,N_6238);
and U6316 (N_6316,N_6235,N_6085);
nand U6317 (N_6317,N_6126,N_6187);
nand U6318 (N_6318,N_6088,N_6125);
or U6319 (N_6319,N_6212,N_6166);
and U6320 (N_6320,N_6210,N_6087);
nor U6321 (N_6321,N_6212,N_6184);
nor U6322 (N_6322,N_6194,N_6206);
and U6323 (N_6323,N_6158,N_6219);
or U6324 (N_6324,N_6164,N_6238);
or U6325 (N_6325,N_6223,N_6085);
or U6326 (N_6326,N_6145,N_6161);
xnor U6327 (N_6327,N_6196,N_6182);
and U6328 (N_6328,N_6177,N_6089);
and U6329 (N_6329,N_6151,N_6133);
nand U6330 (N_6330,N_6147,N_6168);
or U6331 (N_6331,N_6098,N_6121);
and U6332 (N_6332,N_6213,N_6199);
nand U6333 (N_6333,N_6090,N_6219);
and U6334 (N_6334,N_6084,N_6145);
nand U6335 (N_6335,N_6111,N_6141);
or U6336 (N_6336,N_6186,N_6207);
and U6337 (N_6337,N_6120,N_6094);
xnor U6338 (N_6338,N_6220,N_6225);
nand U6339 (N_6339,N_6152,N_6132);
xnor U6340 (N_6340,N_6115,N_6226);
and U6341 (N_6341,N_6228,N_6132);
xor U6342 (N_6342,N_6110,N_6129);
nand U6343 (N_6343,N_6085,N_6204);
nor U6344 (N_6344,N_6236,N_6179);
nand U6345 (N_6345,N_6090,N_6108);
nor U6346 (N_6346,N_6184,N_6233);
xnor U6347 (N_6347,N_6102,N_6151);
or U6348 (N_6348,N_6184,N_6140);
and U6349 (N_6349,N_6136,N_6153);
nor U6350 (N_6350,N_6107,N_6104);
and U6351 (N_6351,N_6153,N_6137);
xor U6352 (N_6352,N_6157,N_6084);
and U6353 (N_6353,N_6158,N_6177);
or U6354 (N_6354,N_6129,N_6210);
or U6355 (N_6355,N_6105,N_6232);
xnor U6356 (N_6356,N_6141,N_6177);
nor U6357 (N_6357,N_6182,N_6129);
or U6358 (N_6358,N_6235,N_6093);
nor U6359 (N_6359,N_6227,N_6088);
or U6360 (N_6360,N_6204,N_6125);
or U6361 (N_6361,N_6161,N_6217);
xor U6362 (N_6362,N_6114,N_6161);
or U6363 (N_6363,N_6128,N_6091);
nand U6364 (N_6364,N_6172,N_6151);
nand U6365 (N_6365,N_6137,N_6145);
nor U6366 (N_6366,N_6164,N_6231);
nand U6367 (N_6367,N_6126,N_6165);
nor U6368 (N_6368,N_6105,N_6141);
or U6369 (N_6369,N_6149,N_6235);
xnor U6370 (N_6370,N_6200,N_6102);
and U6371 (N_6371,N_6167,N_6130);
nor U6372 (N_6372,N_6105,N_6228);
and U6373 (N_6373,N_6175,N_6144);
nand U6374 (N_6374,N_6166,N_6099);
or U6375 (N_6375,N_6214,N_6116);
nand U6376 (N_6376,N_6207,N_6139);
and U6377 (N_6377,N_6207,N_6130);
xor U6378 (N_6378,N_6153,N_6161);
nand U6379 (N_6379,N_6113,N_6204);
xnor U6380 (N_6380,N_6121,N_6180);
nor U6381 (N_6381,N_6199,N_6118);
nor U6382 (N_6382,N_6160,N_6223);
xnor U6383 (N_6383,N_6081,N_6130);
or U6384 (N_6384,N_6231,N_6168);
and U6385 (N_6385,N_6231,N_6221);
xnor U6386 (N_6386,N_6191,N_6169);
nand U6387 (N_6387,N_6201,N_6122);
nand U6388 (N_6388,N_6183,N_6169);
nor U6389 (N_6389,N_6211,N_6112);
or U6390 (N_6390,N_6142,N_6233);
nand U6391 (N_6391,N_6107,N_6226);
or U6392 (N_6392,N_6176,N_6214);
and U6393 (N_6393,N_6160,N_6191);
nor U6394 (N_6394,N_6236,N_6225);
nor U6395 (N_6395,N_6178,N_6101);
xnor U6396 (N_6396,N_6180,N_6084);
and U6397 (N_6397,N_6139,N_6089);
or U6398 (N_6398,N_6090,N_6237);
nand U6399 (N_6399,N_6162,N_6138);
nand U6400 (N_6400,N_6266,N_6253);
xnor U6401 (N_6401,N_6378,N_6366);
nand U6402 (N_6402,N_6276,N_6341);
and U6403 (N_6403,N_6326,N_6286);
nor U6404 (N_6404,N_6395,N_6296);
nand U6405 (N_6405,N_6290,N_6312);
nor U6406 (N_6406,N_6375,N_6351);
or U6407 (N_6407,N_6371,N_6343);
xor U6408 (N_6408,N_6386,N_6263);
nor U6409 (N_6409,N_6323,N_6272);
nand U6410 (N_6410,N_6259,N_6324);
and U6411 (N_6411,N_6338,N_6251);
or U6412 (N_6412,N_6269,N_6317);
and U6413 (N_6413,N_6254,N_6244);
xnor U6414 (N_6414,N_6289,N_6340);
and U6415 (N_6415,N_6275,N_6325);
nand U6416 (N_6416,N_6242,N_6358);
or U6417 (N_6417,N_6398,N_6241);
or U6418 (N_6418,N_6359,N_6288);
nand U6419 (N_6419,N_6397,N_6299);
nor U6420 (N_6420,N_6303,N_6334);
nor U6421 (N_6421,N_6311,N_6295);
nor U6422 (N_6422,N_6256,N_6240);
and U6423 (N_6423,N_6328,N_6387);
or U6424 (N_6424,N_6377,N_6383);
and U6425 (N_6425,N_6390,N_6292);
or U6426 (N_6426,N_6318,N_6307);
or U6427 (N_6427,N_6319,N_6285);
nand U6428 (N_6428,N_6339,N_6279);
xnor U6429 (N_6429,N_6368,N_6283);
and U6430 (N_6430,N_6332,N_6360);
and U6431 (N_6431,N_6249,N_6393);
or U6432 (N_6432,N_6373,N_6287);
xnor U6433 (N_6433,N_6273,N_6258);
nor U6434 (N_6434,N_6374,N_6322);
and U6435 (N_6435,N_6362,N_6297);
nand U6436 (N_6436,N_6267,N_6284);
and U6437 (N_6437,N_6293,N_6392);
nor U6438 (N_6438,N_6309,N_6274);
nor U6439 (N_6439,N_6335,N_6260);
or U6440 (N_6440,N_6252,N_6321);
and U6441 (N_6441,N_6261,N_6278);
or U6442 (N_6442,N_6384,N_6347);
and U6443 (N_6443,N_6300,N_6294);
nand U6444 (N_6444,N_6389,N_6245);
or U6445 (N_6445,N_6350,N_6320);
and U6446 (N_6446,N_6361,N_6337);
nor U6447 (N_6447,N_6342,N_6280);
or U6448 (N_6448,N_6376,N_6363);
or U6449 (N_6449,N_6354,N_6316);
xor U6450 (N_6450,N_6255,N_6301);
and U6451 (N_6451,N_6344,N_6348);
xor U6452 (N_6452,N_6247,N_6372);
nor U6453 (N_6453,N_6381,N_6304);
xor U6454 (N_6454,N_6385,N_6305);
xor U6455 (N_6455,N_6357,N_6308);
or U6456 (N_6456,N_6356,N_6302);
nor U6457 (N_6457,N_6310,N_6346);
nor U6458 (N_6458,N_6329,N_6379);
or U6459 (N_6459,N_6291,N_6355);
or U6460 (N_6460,N_6248,N_6396);
nand U6461 (N_6461,N_6353,N_6349);
nor U6462 (N_6462,N_6330,N_6282);
nor U6463 (N_6463,N_6365,N_6243);
xnor U6464 (N_6464,N_6281,N_6250);
nor U6465 (N_6465,N_6382,N_6314);
or U6466 (N_6466,N_6333,N_6264);
nand U6467 (N_6467,N_6277,N_6298);
and U6468 (N_6468,N_6370,N_6399);
and U6469 (N_6469,N_6367,N_6306);
or U6470 (N_6470,N_6369,N_6327);
xnor U6471 (N_6471,N_6265,N_6364);
or U6472 (N_6472,N_6271,N_6336);
nor U6473 (N_6473,N_6391,N_6262);
xnor U6474 (N_6474,N_6315,N_6345);
or U6475 (N_6475,N_6352,N_6313);
or U6476 (N_6476,N_6331,N_6257);
or U6477 (N_6477,N_6246,N_6270);
nor U6478 (N_6478,N_6394,N_6380);
xor U6479 (N_6479,N_6388,N_6268);
nand U6480 (N_6480,N_6397,N_6373);
nor U6481 (N_6481,N_6318,N_6383);
and U6482 (N_6482,N_6324,N_6353);
and U6483 (N_6483,N_6381,N_6240);
nand U6484 (N_6484,N_6320,N_6246);
or U6485 (N_6485,N_6277,N_6301);
nor U6486 (N_6486,N_6266,N_6261);
nand U6487 (N_6487,N_6376,N_6282);
xnor U6488 (N_6488,N_6307,N_6337);
nand U6489 (N_6489,N_6285,N_6298);
or U6490 (N_6490,N_6292,N_6287);
or U6491 (N_6491,N_6397,N_6319);
xnor U6492 (N_6492,N_6323,N_6358);
nand U6493 (N_6493,N_6381,N_6311);
nand U6494 (N_6494,N_6245,N_6267);
or U6495 (N_6495,N_6339,N_6385);
xor U6496 (N_6496,N_6289,N_6353);
nand U6497 (N_6497,N_6395,N_6369);
nand U6498 (N_6498,N_6380,N_6363);
or U6499 (N_6499,N_6388,N_6345);
nand U6500 (N_6500,N_6369,N_6246);
nor U6501 (N_6501,N_6334,N_6392);
and U6502 (N_6502,N_6259,N_6350);
or U6503 (N_6503,N_6372,N_6305);
nor U6504 (N_6504,N_6305,N_6327);
and U6505 (N_6505,N_6368,N_6343);
xor U6506 (N_6506,N_6281,N_6345);
and U6507 (N_6507,N_6264,N_6374);
and U6508 (N_6508,N_6310,N_6268);
xor U6509 (N_6509,N_6388,N_6306);
or U6510 (N_6510,N_6362,N_6266);
or U6511 (N_6511,N_6259,N_6268);
or U6512 (N_6512,N_6356,N_6308);
xor U6513 (N_6513,N_6281,N_6363);
and U6514 (N_6514,N_6294,N_6281);
or U6515 (N_6515,N_6281,N_6370);
nor U6516 (N_6516,N_6252,N_6390);
xnor U6517 (N_6517,N_6273,N_6352);
or U6518 (N_6518,N_6262,N_6389);
xnor U6519 (N_6519,N_6337,N_6359);
nor U6520 (N_6520,N_6347,N_6304);
and U6521 (N_6521,N_6354,N_6329);
xnor U6522 (N_6522,N_6305,N_6259);
xnor U6523 (N_6523,N_6277,N_6348);
nor U6524 (N_6524,N_6314,N_6321);
xor U6525 (N_6525,N_6399,N_6298);
xnor U6526 (N_6526,N_6307,N_6354);
and U6527 (N_6527,N_6361,N_6312);
nor U6528 (N_6528,N_6331,N_6333);
xnor U6529 (N_6529,N_6319,N_6274);
or U6530 (N_6530,N_6327,N_6357);
xor U6531 (N_6531,N_6349,N_6384);
nand U6532 (N_6532,N_6332,N_6342);
and U6533 (N_6533,N_6270,N_6396);
nor U6534 (N_6534,N_6378,N_6342);
and U6535 (N_6535,N_6294,N_6359);
xor U6536 (N_6536,N_6246,N_6301);
and U6537 (N_6537,N_6346,N_6301);
and U6538 (N_6538,N_6265,N_6247);
or U6539 (N_6539,N_6272,N_6253);
xnor U6540 (N_6540,N_6355,N_6313);
nor U6541 (N_6541,N_6358,N_6252);
or U6542 (N_6542,N_6275,N_6362);
xnor U6543 (N_6543,N_6363,N_6247);
xor U6544 (N_6544,N_6294,N_6385);
or U6545 (N_6545,N_6311,N_6360);
or U6546 (N_6546,N_6330,N_6384);
nand U6547 (N_6547,N_6331,N_6386);
and U6548 (N_6548,N_6331,N_6264);
and U6549 (N_6549,N_6241,N_6246);
nand U6550 (N_6550,N_6349,N_6373);
and U6551 (N_6551,N_6322,N_6288);
nand U6552 (N_6552,N_6285,N_6277);
nand U6553 (N_6553,N_6309,N_6314);
nor U6554 (N_6554,N_6384,N_6355);
and U6555 (N_6555,N_6399,N_6344);
and U6556 (N_6556,N_6245,N_6345);
xnor U6557 (N_6557,N_6366,N_6386);
xor U6558 (N_6558,N_6368,N_6326);
xor U6559 (N_6559,N_6287,N_6248);
nor U6560 (N_6560,N_6481,N_6400);
or U6561 (N_6561,N_6541,N_6410);
and U6562 (N_6562,N_6407,N_6488);
and U6563 (N_6563,N_6540,N_6491);
nand U6564 (N_6564,N_6433,N_6442);
or U6565 (N_6565,N_6431,N_6483);
xor U6566 (N_6566,N_6469,N_6518);
nand U6567 (N_6567,N_6409,N_6444);
xnor U6568 (N_6568,N_6496,N_6454);
and U6569 (N_6569,N_6545,N_6430);
nor U6570 (N_6570,N_6429,N_6477);
and U6571 (N_6571,N_6402,N_6445);
or U6572 (N_6572,N_6417,N_6459);
xnor U6573 (N_6573,N_6494,N_6464);
nor U6574 (N_6574,N_6493,N_6449);
xnor U6575 (N_6575,N_6471,N_6549);
or U6576 (N_6576,N_6447,N_6425);
xnor U6577 (N_6577,N_6415,N_6466);
and U6578 (N_6578,N_6453,N_6420);
nand U6579 (N_6579,N_6538,N_6486);
or U6580 (N_6580,N_6474,N_6476);
xnor U6581 (N_6581,N_6551,N_6547);
nor U6582 (N_6582,N_6537,N_6472);
nor U6583 (N_6583,N_6475,N_6534);
nand U6584 (N_6584,N_6467,N_6519);
and U6585 (N_6585,N_6441,N_6437);
or U6586 (N_6586,N_6531,N_6497);
xor U6587 (N_6587,N_6416,N_6499);
or U6588 (N_6588,N_6542,N_6461);
or U6589 (N_6589,N_6487,N_6527);
or U6590 (N_6590,N_6452,N_6543);
nand U6591 (N_6591,N_6455,N_6530);
or U6592 (N_6592,N_6546,N_6553);
nor U6593 (N_6593,N_6432,N_6470);
or U6594 (N_6594,N_6423,N_6501);
xor U6595 (N_6595,N_6460,N_6536);
and U6596 (N_6596,N_6507,N_6502);
nor U6597 (N_6597,N_6510,N_6480);
nand U6598 (N_6598,N_6490,N_6424);
and U6599 (N_6599,N_6558,N_6411);
xnor U6600 (N_6600,N_6427,N_6500);
nor U6601 (N_6601,N_6406,N_6413);
or U6602 (N_6602,N_6448,N_6495);
and U6603 (N_6603,N_6463,N_6539);
and U6604 (N_6604,N_6462,N_6446);
nor U6605 (N_6605,N_6485,N_6506);
xnor U6606 (N_6606,N_6405,N_6555);
or U6607 (N_6607,N_6465,N_6440);
and U6608 (N_6608,N_6532,N_6522);
nor U6609 (N_6609,N_6509,N_6514);
nand U6610 (N_6610,N_6548,N_6443);
nand U6611 (N_6611,N_6505,N_6438);
xnor U6612 (N_6612,N_6529,N_6528);
or U6613 (N_6613,N_6404,N_6556);
nand U6614 (N_6614,N_6523,N_6414);
nor U6615 (N_6615,N_6428,N_6412);
and U6616 (N_6616,N_6439,N_6408);
or U6617 (N_6617,N_6451,N_6456);
or U6618 (N_6618,N_6554,N_6434);
and U6619 (N_6619,N_6473,N_6482);
nor U6620 (N_6620,N_6478,N_6489);
or U6621 (N_6621,N_6418,N_6401);
nor U6622 (N_6622,N_6484,N_6511);
nand U6623 (N_6623,N_6513,N_6544);
nand U6624 (N_6624,N_6422,N_6535);
and U6625 (N_6625,N_6517,N_6498);
nand U6626 (N_6626,N_6403,N_6479);
xnor U6627 (N_6627,N_6457,N_6468);
nor U6628 (N_6628,N_6435,N_6524);
nand U6629 (N_6629,N_6508,N_6557);
nand U6630 (N_6630,N_6516,N_6559);
nand U6631 (N_6631,N_6552,N_6521);
xnor U6632 (N_6632,N_6550,N_6421);
nor U6633 (N_6633,N_6492,N_6520);
xnor U6634 (N_6634,N_6526,N_6436);
nand U6635 (N_6635,N_6512,N_6533);
and U6636 (N_6636,N_6525,N_6450);
nand U6637 (N_6637,N_6458,N_6515);
or U6638 (N_6638,N_6503,N_6504);
and U6639 (N_6639,N_6426,N_6419);
nor U6640 (N_6640,N_6541,N_6519);
or U6641 (N_6641,N_6489,N_6525);
xor U6642 (N_6642,N_6500,N_6465);
or U6643 (N_6643,N_6487,N_6517);
nor U6644 (N_6644,N_6523,N_6547);
or U6645 (N_6645,N_6426,N_6470);
or U6646 (N_6646,N_6478,N_6445);
nor U6647 (N_6647,N_6433,N_6460);
xnor U6648 (N_6648,N_6541,N_6432);
or U6649 (N_6649,N_6516,N_6415);
nor U6650 (N_6650,N_6552,N_6491);
xnor U6651 (N_6651,N_6484,N_6426);
nor U6652 (N_6652,N_6544,N_6459);
and U6653 (N_6653,N_6490,N_6507);
nor U6654 (N_6654,N_6443,N_6435);
xnor U6655 (N_6655,N_6500,N_6482);
xor U6656 (N_6656,N_6539,N_6411);
nand U6657 (N_6657,N_6476,N_6504);
and U6658 (N_6658,N_6418,N_6520);
xnor U6659 (N_6659,N_6516,N_6434);
xnor U6660 (N_6660,N_6488,N_6422);
and U6661 (N_6661,N_6483,N_6409);
nand U6662 (N_6662,N_6470,N_6524);
and U6663 (N_6663,N_6438,N_6500);
nand U6664 (N_6664,N_6419,N_6535);
and U6665 (N_6665,N_6418,N_6541);
or U6666 (N_6666,N_6527,N_6471);
nand U6667 (N_6667,N_6472,N_6556);
xnor U6668 (N_6668,N_6534,N_6424);
nor U6669 (N_6669,N_6408,N_6419);
nand U6670 (N_6670,N_6460,N_6469);
nor U6671 (N_6671,N_6499,N_6526);
xor U6672 (N_6672,N_6501,N_6528);
or U6673 (N_6673,N_6414,N_6489);
and U6674 (N_6674,N_6490,N_6543);
xor U6675 (N_6675,N_6519,N_6546);
xor U6676 (N_6676,N_6513,N_6430);
nor U6677 (N_6677,N_6514,N_6452);
xnor U6678 (N_6678,N_6461,N_6550);
or U6679 (N_6679,N_6486,N_6508);
xnor U6680 (N_6680,N_6558,N_6424);
xor U6681 (N_6681,N_6499,N_6506);
nor U6682 (N_6682,N_6401,N_6406);
nand U6683 (N_6683,N_6416,N_6427);
nor U6684 (N_6684,N_6479,N_6497);
nand U6685 (N_6685,N_6491,N_6498);
nor U6686 (N_6686,N_6402,N_6554);
or U6687 (N_6687,N_6487,N_6416);
nor U6688 (N_6688,N_6436,N_6449);
xor U6689 (N_6689,N_6445,N_6483);
or U6690 (N_6690,N_6482,N_6550);
and U6691 (N_6691,N_6522,N_6487);
nor U6692 (N_6692,N_6466,N_6520);
xor U6693 (N_6693,N_6495,N_6423);
xor U6694 (N_6694,N_6438,N_6471);
or U6695 (N_6695,N_6450,N_6541);
and U6696 (N_6696,N_6509,N_6452);
nor U6697 (N_6697,N_6474,N_6440);
and U6698 (N_6698,N_6532,N_6407);
nand U6699 (N_6699,N_6484,N_6523);
nor U6700 (N_6700,N_6521,N_6453);
and U6701 (N_6701,N_6447,N_6503);
nor U6702 (N_6702,N_6406,N_6519);
and U6703 (N_6703,N_6437,N_6444);
nand U6704 (N_6704,N_6503,N_6414);
or U6705 (N_6705,N_6464,N_6416);
nand U6706 (N_6706,N_6553,N_6535);
xor U6707 (N_6707,N_6480,N_6513);
nor U6708 (N_6708,N_6543,N_6507);
and U6709 (N_6709,N_6529,N_6520);
nor U6710 (N_6710,N_6552,N_6498);
xor U6711 (N_6711,N_6533,N_6402);
xnor U6712 (N_6712,N_6465,N_6445);
xnor U6713 (N_6713,N_6545,N_6412);
nor U6714 (N_6714,N_6525,N_6559);
and U6715 (N_6715,N_6505,N_6495);
nand U6716 (N_6716,N_6551,N_6485);
and U6717 (N_6717,N_6407,N_6471);
nor U6718 (N_6718,N_6477,N_6491);
or U6719 (N_6719,N_6526,N_6401);
or U6720 (N_6720,N_6674,N_6569);
nand U6721 (N_6721,N_6570,N_6612);
or U6722 (N_6722,N_6639,N_6624);
xnor U6723 (N_6723,N_6646,N_6704);
nand U6724 (N_6724,N_6626,N_6564);
and U6725 (N_6725,N_6606,N_6631);
nor U6726 (N_6726,N_6677,N_6621);
or U6727 (N_6727,N_6701,N_6579);
xor U6728 (N_6728,N_6574,N_6689);
xnor U6729 (N_6729,N_6685,N_6708);
xor U6730 (N_6730,N_6647,N_6585);
and U6731 (N_6731,N_6660,N_6661);
nor U6732 (N_6732,N_6607,N_6697);
or U6733 (N_6733,N_6693,N_6627);
nand U6734 (N_6734,N_6658,N_6637);
xnor U6735 (N_6735,N_6649,N_6571);
xor U6736 (N_6736,N_6586,N_6614);
nand U6737 (N_6737,N_6640,N_6625);
xnor U6738 (N_6738,N_6590,N_6623);
xor U6739 (N_6739,N_6609,N_6713);
and U6740 (N_6740,N_6691,N_6589);
nand U6741 (N_6741,N_6615,N_6657);
xnor U6742 (N_6742,N_6694,N_6618);
nor U6743 (N_6743,N_6619,N_6703);
nor U6744 (N_6744,N_6715,N_6671);
and U6745 (N_6745,N_6659,N_6710);
or U6746 (N_6746,N_6702,N_6645);
nor U6747 (N_6747,N_6666,N_6563);
and U6748 (N_6748,N_6641,N_6642);
nor U6749 (N_6749,N_6672,N_6599);
nor U6750 (N_6750,N_6651,N_6673);
xor U6751 (N_6751,N_6578,N_6565);
and U6752 (N_6752,N_6678,N_6718);
and U6753 (N_6753,N_6605,N_6633);
or U6754 (N_6754,N_6650,N_6603);
nor U6755 (N_6755,N_6705,N_6665);
xor U6756 (N_6756,N_6617,N_6695);
xnor U6757 (N_6757,N_6616,N_6652);
or U6758 (N_6758,N_6596,N_6613);
and U6759 (N_6759,N_6577,N_6682);
nand U6760 (N_6760,N_6676,N_6573);
nand U6761 (N_6761,N_6561,N_6698);
xor U6762 (N_6762,N_6632,N_6668);
nor U6763 (N_6763,N_6654,N_6560);
nand U6764 (N_6764,N_6719,N_6629);
nor U6765 (N_6765,N_6593,N_6669);
and U6766 (N_6766,N_6610,N_6663);
nor U6767 (N_6767,N_6587,N_6601);
xnor U6768 (N_6768,N_6670,N_6716);
and U6769 (N_6769,N_6622,N_6602);
and U6770 (N_6770,N_6594,N_6636);
xnor U6771 (N_6771,N_6584,N_6608);
xor U6772 (N_6772,N_6644,N_6684);
xnor U6773 (N_6773,N_6583,N_6580);
nand U6774 (N_6774,N_6591,N_6683);
nand U6775 (N_6775,N_6575,N_6709);
xnor U6776 (N_6776,N_6634,N_6581);
xor U6777 (N_6777,N_6597,N_6686);
xor U6778 (N_6778,N_6706,N_6648);
or U6779 (N_6779,N_6717,N_6568);
nand U6780 (N_6780,N_6696,N_6604);
nor U6781 (N_6781,N_6667,N_6679);
nor U6782 (N_6782,N_6681,N_6572);
xor U6783 (N_6783,N_6712,N_6638);
nor U6784 (N_6784,N_6598,N_6664);
or U6785 (N_6785,N_6595,N_6711);
nand U6786 (N_6786,N_6714,N_6620);
xnor U6787 (N_6787,N_6576,N_6567);
and U6788 (N_6788,N_6643,N_6566);
or U6789 (N_6789,N_6582,N_6588);
nand U6790 (N_6790,N_6600,N_6680);
xnor U6791 (N_6791,N_6611,N_6656);
and U6792 (N_6792,N_6630,N_6692);
xnor U6793 (N_6793,N_6653,N_6662);
or U6794 (N_6794,N_6699,N_6707);
and U6795 (N_6795,N_6700,N_6687);
or U6796 (N_6796,N_6690,N_6562);
nor U6797 (N_6797,N_6655,N_6688);
nand U6798 (N_6798,N_6675,N_6635);
nand U6799 (N_6799,N_6592,N_6628);
nand U6800 (N_6800,N_6718,N_6669);
nor U6801 (N_6801,N_6715,N_6584);
and U6802 (N_6802,N_6595,N_6596);
nor U6803 (N_6803,N_6595,N_6577);
or U6804 (N_6804,N_6699,N_6602);
nand U6805 (N_6805,N_6659,N_6704);
nand U6806 (N_6806,N_6601,N_6600);
nor U6807 (N_6807,N_6655,N_6568);
nor U6808 (N_6808,N_6675,N_6595);
nor U6809 (N_6809,N_6563,N_6593);
xor U6810 (N_6810,N_6676,N_6639);
or U6811 (N_6811,N_6637,N_6677);
nor U6812 (N_6812,N_6612,N_6637);
and U6813 (N_6813,N_6699,N_6588);
nand U6814 (N_6814,N_6654,N_6588);
nand U6815 (N_6815,N_6663,N_6674);
and U6816 (N_6816,N_6670,N_6659);
nand U6817 (N_6817,N_6654,N_6661);
nand U6818 (N_6818,N_6703,N_6661);
nor U6819 (N_6819,N_6582,N_6673);
nand U6820 (N_6820,N_6675,N_6651);
xor U6821 (N_6821,N_6597,N_6571);
nor U6822 (N_6822,N_6641,N_6673);
or U6823 (N_6823,N_6572,N_6689);
nand U6824 (N_6824,N_6573,N_6708);
and U6825 (N_6825,N_6680,N_6716);
and U6826 (N_6826,N_6684,N_6629);
and U6827 (N_6827,N_6708,N_6613);
xor U6828 (N_6828,N_6637,N_6568);
xnor U6829 (N_6829,N_6693,N_6610);
or U6830 (N_6830,N_6626,N_6603);
or U6831 (N_6831,N_6654,N_6677);
nand U6832 (N_6832,N_6644,N_6710);
nor U6833 (N_6833,N_6714,N_6709);
xnor U6834 (N_6834,N_6621,N_6627);
xnor U6835 (N_6835,N_6663,N_6642);
nor U6836 (N_6836,N_6634,N_6599);
xnor U6837 (N_6837,N_6563,N_6704);
xnor U6838 (N_6838,N_6712,N_6632);
and U6839 (N_6839,N_6598,N_6623);
xnor U6840 (N_6840,N_6574,N_6567);
or U6841 (N_6841,N_6569,N_6620);
and U6842 (N_6842,N_6595,N_6705);
xnor U6843 (N_6843,N_6577,N_6658);
nor U6844 (N_6844,N_6587,N_6701);
nor U6845 (N_6845,N_6577,N_6704);
nand U6846 (N_6846,N_6628,N_6627);
xor U6847 (N_6847,N_6653,N_6679);
xnor U6848 (N_6848,N_6639,N_6567);
and U6849 (N_6849,N_6656,N_6566);
or U6850 (N_6850,N_6702,N_6695);
nand U6851 (N_6851,N_6623,N_6624);
nor U6852 (N_6852,N_6683,N_6663);
and U6853 (N_6853,N_6716,N_6584);
nand U6854 (N_6854,N_6560,N_6617);
or U6855 (N_6855,N_6660,N_6716);
nand U6856 (N_6856,N_6678,N_6569);
and U6857 (N_6857,N_6714,N_6689);
or U6858 (N_6858,N_6593,N_6684);
xor U6859 (N_6859,N_6566,N_6649);
xor U6860 (N_6860,N_6675,N_6604);
and U6861 (N_6861,N_6713,N_6665);
or U6862 (N_6862,N_6693,N_6563);
xor U6863 (N_6863,N_6632,N_6646);
nor U6864 (N_6864,N_6667,N_6713);
xor U6865 (N_6865,N_6638,N_6656);
xor U6866 (N_6866,N_6711,N_6563);
or U6867 (N_6867,N_6676,N_6652);
xor U6868 (N_6868,N_6563,N_6605);
nand U6869 (N_6869,N_6662,N_6596);
nand U6870 (N_6870,N_6566,N_6642);
xnor U6871 (N_6871,N_6715,N_6678);
nand U6872 (N_6872,N_6713,N_6607);
or U6873 (N_6873,N_6713,N_6642);
and U6874 (N_6874,N_6572,N_6675);
nor U6875 (N_6875,N_6613,N_6597);
and U6876 (N_6876,N_6566,N_6694);
or U6877 (N_6877,N_6573,N_6579);
xor U6878 (N_6878,N_6630,N_6585);
xnor U6879 (N_6879,N_6694,N_6593);
nor U6880 (N_6880,N_6741,N_6852);
and U6881 (N_6881,N_6871,N_6726);
nand U6882 (N_6882,N_6805,N_6721);
nor U6883 (N_6883,N_6762,N_6730);
nor U6884 (N_6884,N_6820,N_6786);
nor U6885 (N_6885,N_6767,N_6723);
and U6886 (N_6886,N_6750,N_6831);
nand U6887 (N_6887,N_6783,N_6749);
nand U6888 (N_6888,N_6864,N_6804);
nor U6889 (N_6889,N_6785,N_6821);
and U6890 (N_6890,N_6791,N_6859);
nor U6891 (N_6891,N_6722,N_6838);
and U6892 (N_6892,N_6769,N_6737);
nand U6893 (N_6893,N_6728,N_6744);
nor U6894 (N_6894,N_6873,N_6828);
nand U6895 (N_6895,N_6846,N_6729);
nor U6896 (N_6896,N_6827,N_6819);
or U6897 (N_6897,N_6810,N_6853);
nand U6898 (N_6898,N_6866,N_6860);
nand U6899 (N_6899,N_6836,N_6862);
nor U6900 (N_6900,N_6840,N_6752);
and U6901 (N_6901,N_6832,N_6724);
or U6902 (N_6902,N_6841,N_6878);
xnor U6903 (N_6903,N_6758,N_6787);
and U6904 (N_6904,N_6754,N_6867);
nor U6905 (N_6905,N_6796,N_6770);
and U6906 (N_6906,N_6748,N_6835);
nor U6907 (N_6907,N_6826,N_6868);
nor U6908 (N_6908,N_6809,N_6822);
nand U6909 (N_6909,N_6772,N_6742);
nor U6910 (N_6910,N_6800,N_6794);
nand U6911 (N_6911,N_6837,N_6830);
nand U6912 (N_6912,N_6773,N_6825);
or U6913 (N_6913,N_6782,N_6760);
xor U6914 (N_6914,N_6848,N_6815);
and U6915 (N_6915,N_6874,N_6823);
and U6916 (N_6916,N_6855,N_6842);
xor U6917 (N_6917,N_6824,N_6793);
nand U6918 (N_6918,N_6776,N_6829);
nand U6919 (N_6919,N_6764,N_6774);
nor U6920 (N_6920,N_6807,N_6735);
and U6921 (N_6921,N_6869,N_6799);
or U6922 (N_6922,N_6775,N_6759);
nor U6923 (N_6923,N_6813,N_6751);
or U6924 (N_6924,N_6757,N_6734);
nand U6925 (N_6925,N_6756,N_6797);
nand U6926 (N_6926,N_6738,N_6814);
nand U6927 (N_6927,N_6863,N_6747);
nand U6928 (N_6928,N_6788,N_6798);
and U6929 (N_6929,N_6789,N_6865);
xnor U6930 (N_6930,N_6745,N_6850);
nand U6931 (N_6931,N_6795,N_6849);
nand U6932 (N_6932,N_6872,N_6736);
and U6933 (N_6933,N_6780,N_6765);
or U6934 (N_6934,N_6802,N_6879);
nand U6935 (N_6935,N_6870,N_6854);
xnor U6936 (N_6936,N_6740,N_6818);
xnor U6937 (N_6937,N_6803,N_6851);
nand U6938 (N_6938,N_6743,N_6781);
xnor U6939 (N_6939,N_6801,N_6766);
and U6940 (N_6940,N_6861,N_6843);
nor U6941 (N_6941,N_6845,N_6817);
nand U6942 (N_6942,N_6856,N_6720);
and U6943 (N_6943,N_6763,N_6790);
nand U6944 (N_6944,N_6732,N_6844);
nor U6945 (N_6945,N_6746,N_6847);
xor U6946 (N_6946,N_6727,N_6857);
nor U6947 (N_6947,N_6877,N_6733);
nand U6948 (N_6948,N_6753,N_6778);
xnor U6949 (N_6949,N_6739,N_6811);
or U6950 (N_6950,N_6833,N_6816);
and U6951 (N_6951,N_6839,N_6725);
or U6952 (N_6952,N_6731,N_6768);
nor U6953 (N_6953,N_6858,N_6784);
and U6954 (N_6954,N_6834,N_6808);
and U6955 (N_6955,N_6876,N_6806);
and U6956 (N_6956,N_6771,N_6779);
nand U6957 (N_6957,N_6761,N_6875);
xnor U6958 (N_6958,N_6812,N_6755);
nand U6959 (N_6959,N_6777,N_6792);
and U6960 (N_6960,N_6819,N_6768);
nand U6961 (N_6961,N_6817,N_6871);
nor U6962 (N_6962,N_6864,N_6786);
or U6963 (N_6963,N_6867,N_6873);
nor U6964 (N_6964,N_6878,N_6741);
xnor U6965 (N_6965,N_6812,N_6774);
or U6966 (N_6966,N_6757,N_6731);
nand U6967 (N_6967,N_6748,N_6824);
or U6968 (N_6968,N_6740,N_6744);
nand U6969 (N_6969,N_6726,N_6851);
nor U6970 (N_6970,N_6839,N_6784);
nor U6971 (N_6971,N_6839,N_6832);
nand U6972 (N_6972,N_6783,N_6756);
or U6973 (N_6973,N_6879,N_6862);
and U6974 (N_6974,N_6842,N_6749);
or U6975 (N_6975,N_6878,N_6781);
and U6976 (N_6976,N_6856,N_6742);
xor U6977 (N_6977,N_6744,N_6794);
nand U6978 (N_6978,N_6863,N_6846);
xnor U6979 (N_6979,N_6845,N_6848);
nand U6980 (N_6980,N_6747,N_6828);
and U6981 (N_6981,N_6859,N_6738);
and U6982 (N_6982,N_6759,N_6870);
and U6983 (N_6983,N_6879,N_6741);
or U6984 (N_6984,N_6771,N_6833);
or U6985 (N_6985,N_6740,N_6783);
nand U6986 (N_6986,N_6745,N_6766);
or U6987 (N_6987,N_6828,N_6762);
and U6988 (N_6988,N_6794,N_6831);
nand U6989 (N_6989,N_6745,N_6767);
and U6990 (N_6990,N_6825,N_6772);
and U6991 (N_6991,N_6786,N_6874);
or U6992 (N_6992,N_6820,N_6768);
nand U6993 (N_6993,N_6840,N_6848);
nand U6994 (N_6994,N_6800,N_6729);
and U6995 (N_6995,N_6868,N_6854);
or U6996 (N_6996,N_6727,N_6856);
nor U6997 (N_6997,N_6823,N_6783);
nand U6998 (N_6998,N_6856,N_6793);
nor U6999 (N_6999,N_6789,N_6786);
or U7000 (N_7000,N_6793,N_6744);
nand U7001 (N_7001,N_6827,N_6795);
or U7002 (N_7002,N_6757,N_6761);
xnor U7003 (N_7003,N_6828,N_6844);
xor U7004 (N_7004,N_6803,N_6724);
and U7005 (N_7005,N_6732,N_6819);
nand U7006 (N_7006,N_6809,N_6839);
xor U7007 (N_7007,N_6845,N_6761);
nor U7008 (N_7008,N_6792,N_6766);
nor U7009 (N_7009,N_6738,N_6733);
xnor U7010 (N_7010,N_6733,N_6765);
and U7011 (N_7011,N_6818,N_6776);
xnor U7012 (N_7012,N_6788,N_6866);
or U7013 (N_7013,N_6772,N_6820);
and U7014 (N_7014,N_6866,N_6808);
or U7015 (N_7015,N_6763,N_6815);
and U7016 (N_7016,N_6756,N_6827);
nor U7017 (N_7017,N_6738,N_6721);
and U7018 (N_7018,N_6772,N_6843);
nor U7019 (N_7019,N_6841,N_6787);
nor U7020 (N_7020,N_6878,N_6758);
nand U7021 (N_7021,N_6841,N_6791);
or U7022 (N_7022,N_6788,N_6848);
or U7023 (N_7023,N_6820,N_6868);
and U7024 (N_7024,N_6792,N_6850);
nand U7025 (N_7025,N_6733,N_6865);
xor U7026 (N_7026,N_6858,N_6852);
nand U7027 (N_7027,N_6751,N_6761);
and U7028 (N_7028,N_6816,N_6743);
nor U7029 (N_7029,N_6788,N_6757);
or U7030 (N_7030,N_6755,N_6801);
xnor U7031 (N_7031,N_6844,N_6728);
or U7032 (N_7032,N_6757,N_6841);
nor U7033 (N_7033,N_6759,N_6840);
nand U7034 (N_7034,N_6784,N_6807);
xnor U7035 (N_7035,N_6847,N_6842);
xor U7036 (N_7036,N_6841,N_6785);
and U7037 (N_7037,N_6856,N_6758);
nor U7038 (N_7038,N_6779,N_6861);
or U7039 (N_7039,N_6873,N_6831);
nor U7040 (N_7040,N_6888,N_7021);
nor U7041 (N_7041,N_6914,N_6881);
or U7042 (N_7042,N_6981,N_7005);
and U7043 (N_7043,N_7019,N_7039);
or U7044 (N_7044,N_6901,N_6934);
and U7045 (N_7045,N_6972,N_6916);
or U7046 (N_7046,N_6909,N_6929);
and U7047 (N_7047,N_6883,N_7026);
or U7048 (N_7048,N_7036,N_6890);
or U7049 (N_7049,N_6894,N_6985);
xnor U7050 (N_7050,N_7006,N_6925);
xnor U7051 (N_7051,N_6963,N_6922);
nand U7052 (N_7052,N_6898,N_6994);
nor U7053 (N_7053,N_6954,N_7017);
and U7054 (N_7054,N_7010,N_6998);
nand U7055 (N_7055,N_7007,N_6880);
or U7056 (N_7056,N_6990,N_6900);
nand U7057 (N_7057,N_6882,N_7034);
or U7058 (N_7058,N_6932,N_7008);
nand U7059 (N_7059,N_6906,N_7033);
and U7060 (N_7060,N_6889,N_7009);
or U7061 (N_7061,N_6957,N_7022);
nor U7062 (N_7062,N_7004,N_6975);
and U7063 (N_7063,N_6965,N_6886);
and U7064 (N_7064,N_6945,N_6895);
and U7065 (N_7065,N_6977,N_6943);
nor U7066 (N_7066,N_7027,N_6885);
or U7067 (N_7067,N_6938,N_6988);
xor U7068 (N_7068,N_6921,N_7016);
xor U7069 (N_7069,N_6920,N_6941);
or U7070 (N_7070,N_7030,N_6903);
and U7071 (N_7071,N_6911,N_6986);
nand U7072 (N_7072,N_6951,N_7031);
xor U7073 (N_7073,N_7020,N_6924);
nand U7074 (N_7074,N_7001,N_6939);
and U7075 (N_7075,N_7014,N_6960);
and U7076 (N_7076,N_7000,N_6896);
xnor U7077 (N_7077,N_6899,N_6973);
xor U7078 (N_7078,N_7018,N_6980);
xnor U7079 (N_7079,N_6908,N_6967);
nand U7080 (N_7080,N_6917,N_6907);
xnor U7081 (N_7081,N_6935,N_6969);
xor U7082 (N_7082,N_7037,N_6955);
or U7083 (N_7083,N_6961,N_7013);
nor U7084 (N_7084,N_7035,N_6946);
and U7085 (N_7085,N_7032,N_6942);
and U7086 (N_7086,N_6966,N_6905);
nand U7087 (N_7087,N_6971,N_6897);
or U7088 (N_7088,N_6997,N_6956);
nand U7089 (N_7089,N_7025,N_6978);
or U7090 (N_7090,N_6964,N_6962);
and U7091 (N_7091,N_6991,N_6919);
nor U7092 (N_7092,N_6902,N_6995);
nand U7093 (N_7093,N_6910,N_6958);
nand U7094 (N_7094,N_6970,N_7023);
nor U7095 (N_7095,N_6928,N_6944);
and U7096 (N_7096,N_6947,N_6940);
and U7097 (N_7097,N_6989,N_7012);
nor U7098 (N_7098,N_6993,N_6933);
nand U7099 (N_7099,N_6923,N_6893);
and U7100 (N_7100,N_6959,N_6982);
nor U7101 (N_7101,N_6983,N_6968);
nand U7102 (N_7102,N_6992,N_6953);
nand U7103 (N_7103,N_6948,N_6984);
nand U7104 (N_7104,N_6987,N_7011);
nor U7105 (N_7105,N_6927,N_7028);
nor U7106 (N_7106,N_6926,N_6976);
nor U7107 (N_7107,N_6915,N_6913);
nand U7108 (N_7108,N_6979,N_7038);
or U7109 (N_7109,N_6952,N_6949);
nor U7110 (N_7110,N_6918,N_6974);
xnor U7111 (N_7111,N_6937,N_6887);
xor U7112 (N_7112,N_7029,N_6936);
nand U7113 (N_7113,N_6904,N_6931);
nor U7114 (N_7114,N_6930,N_6999);
and U7115 (N_7115,N_7015,N_6891);
nand U7116 (N_7116,N_7024,N_6892);
and U7117 (N_7117,N_7003,N_6884);
xnor U7118 (N_7118,N_6950,N_6912);
nor U7119 (N_7119,N_7002,N_6996);
xor U7120 (N_7120,N_6915,N_6957);
nor U7121 (N_7121,N_6928,N_6880);
xor U7122 (N_7122,N_6951,N_7014);
nor U7123 (N_7123,N_6983,N_6932);
nor U7124 (N_7124,N_6886,N_6882);
nor U7125 (N_7125,N_6942,N_6954);
or U7126 (N_7126,N_6967,N_7009);
and U7127 (N_7127,N_6921,N_6996);
nand U7128 (N_7128,N_6892,N_6897);
and U7129 (N_7129,N_6992,N_6963);
nor U7130 (N_7130,N_6925,N_6957);
nor U7131 (N_7131,N_6918,N_6941);
and U7132 (N_7132,N_7023,N_6984);
xor U7133 (N_7133,N_6948,N_6991);
or U7134 (N_7134,N_6912,N_6960);
and U7135 (N_7135,N_7016,N_7007);
nor U7136 (N_7136,N_6919,N_6958);
nor U7137 (N_7137,N_6907,N_6981);
nand U7138 (N_7138,N_6893,N_7025);
or U7139 (N_7139,N_6886,N_7002);
nand U7140 (N_7140,N_6922,N_6957);
xor U7141 (N_7141,N_6994,N_6894);
and U7142 (N_7142,N_7004,N_6908);
xor U7143 (N_7143,N_6887,N_6938);
and U7144 (N_7144,N_6915,N_6912);
xor U7145 (N_7145,N_7017,N_6905);
xnor U7146 (N_7146,N_6907,N_6993);
nor U7147 (N_7147,N_7014,N_7013);
xor U7148 (N_7148,N_6928,N_6916);
or U7149 (N_7149,N_7024,N_6957);
or U7150 (N_7150,N_6945,N_6880);
and U7151 (N_7151,N_6985,N_6926);
xnor U7152 (N_7152,N_6900,N_6886);
nand U7153 (N_7153,N_6999,N_7001);
nor U7154 (N_7154,N_6955,N_6943);
and U7155 (N_7155,N_6941,N_6978);
nor U7156 (N_7156,N_6921,N_6920);
or U7157 (N_7157,N_6946,N_7004);
and U7158 (N_7158,N_7025,N_6973);
nor U7159 (N_7159,N_6956,N_6911);
or U7160 (N_7160,N_6991,N_6909);
nor U7161 (N_7161,N_6904,N_6956);
xor U7162 (N_7162,N_7035,N_6931);
nand U7163 (N_7163,N_6934,N_7036);
xnor U7164 (N_7164,N_6992,N_6918);
and U7165 (N_7165,N_6882,N_6923);
and U7166 (N_7166,N_6986,N_6997);
xor U7167 (N_7167,N_6952,N_6889);
and U7168 (N_7168,N_6924,N_6983);
xnor U7169 (N_7169,N_6984,N_6953);
nand U7170 (N_7170,N_6942,N_6974);
and U7171 (N_7171,N_7025,N_6913);
and U7172 (N_7172,N_6949,N_6888);
xor U7173 (N_7173,N_6920,N_6950);
and U7174 (N_7174,N_6914,N_7026);
nand U7175 (N_7175,N_6904,N_6883);
or U7176 (N_7176,N_7026,N_6889);
or U7177 (N_7177,N_7024,N_7006);
or U7178 (N_7178,N_6884,N_7014);
nand U7179 (N_7179,N_7030,N_6900);
and U7180 (N_7180,N_6901,N_7031);
or U7181 (N_7181,N_7010,N_6995);
or U7182 (N_7182,N_6955,N_6887);
xnor U7183 (N_7183,N_6937,N_6896);
or U7184 (N_7184,N_7019,N_6953);
xor U7185 (N_7185,N_7004,N_6965);
nand U7186 (N_7186,N_7036,N_6988);
xor U7187 (N_7187,N_6995,N_6997);
xnor U7188 (N_7188,N_6951,N_7028);
nand U7189 (N_7189,N_7021,N_6954);
and U7190 (N_7190,N_6954,N_6919);
nand U7191 (N_7191,N_6950,N_6943);
nand U7192 (N_7192,N_7033,N_7001);
xnor U7193 (N_7193,N_6947,N_6970);
nand U7194 (N_7194,N_7030,N_7017);
xnor U7195 (N_7195,N_6996,N_6941);
and U7196 (N_7196,N_6958,N_6943);
and U7197 (N_7197,N_6946,N_6891);
and U7198 (N_7198,N_7011,N_6989);
or U7199 (N_7199,N_6961,N_6919);
nor U7200 (N_7200,N_7040,N_7152);
xnor U7201 (N_7201,N_7184,N_7057);
or U7202 (N_7202,N_7168,N_7051);
or U7203 (N_7203,N_7139,N_7050);
xor U7204 (N_7204,N_7156,N_7115);
xnor U7205 (N_7205,N_7189,N_7082);
or U7206 (N_7206,N_7077,N_7113);
nand U7207 (N_7207,N_7159,N_7148);
nor U7208 (N_7208,N_7197,N_7195);
or U7209 (N_7209,N_7106,N_7178);
nand U7210 (N_7210,N_7171,N_7186);
xnor U7211 (N_7211,N_7138,N_7103);
nand U7212 (N_7212,N_7073,N_7068);
or U7213 (N_7213,N_7058,N_7101);
nand U7214 (N_7214,N_7070,N_7155);
nor U7215 (N_7215,N_7078,N_7137);
nand U7216 (N_7216,N_7169,N_7066);
nand U7217 (N_7217,N_7194,N_7170);
and U7218 (N_7218,N_7188,N_7191);
or U7219 (N_7219,N_7094,N_7192);
nor U7220 (N_7220,N_7112,N_7124);
nor U7221 (N_7221,N_7198,N_7085);
nand U7222 (N_7222,N_7072,N_7143);
xnor U7223 (N_7223,N_7172,N_7132);
nand U7224 (N_7224,N_7097,N_7162);
nand U7225 (N_7225,N_7177,N_7117);
and U7226 (N_7226,N_7063,N_7096);
nor U7227 (N_7227,N_7111,N_7089);
nor U7228 (N_7228,N_7108,N_7056);
nor U7229 (N_7229,N_7190,N_7181);
nor U7230 (N_7230,N_7100,N_7146);
nor U7231 (N_7231,N_7087,N_7067);
or U7232 (N_7232,N_7157,N_7174);
and U7233 (N_7233,N_7061,N_7081);
nor U7234 (N_7234,N_7153,N_7105);
and U7235 (N_7235,N_7166,N_7116);
xor U7236 (N_7236,N_7052,N_7158);
and U7237 (N_7237,N_7144,N_7154);
and U7238 (N_7238,N_7193,N_7048);
or U7239 (N_7239,N_7131,N_7180);
nor U7240 (N_7240,N_7187,N_7109);
xor U7241 (N_7241,N_7069,N_7150);
nand U7242 (N_7242,N_7053,N_7183);
nand U7243 (N_7243,N_7175,N_7062);
or U7244 (N_7244,N_7182,N_7092);
or U7245 (N_7245,N_7133,N_7128);
and U7246 (N_7246,N_7054,N_7104);
nor U7247 (N_7247,N_7071,N_7075);
xnor U7248 (N_7248,N_7130,N_7149);
xnor U7249 (N_7249,N_7119,N_7080);
nor U7250 (N_7250,N_7114,N_7126);
xor U7251 (N_7251,N_7084,N_7042);
nor U7252 (N_7252,N_7163,N_7147);
nor U7253 (N_7253,N_7043,N_7076);
or U7254 (N_7254,N_7074,N_7091);
nor U7255 (N_7255,N_7098,N_7121);
nand U7256 (N_7256,N_7167,N_7118);
nor U7257 (N_7257,N_7123,N_7045);
or U7258 (N_7258,N_7041,N_7161);
nor U7259 (N_7259,N_7095,N_7060);
nor U7260 (N_7260,N_7099,N_7151);
or U7261 (N_7261,N_7064,N_7083);
nand U7262 (N_7262,N_7164,N_7088);
xor U7263 (N_7263,N_7044,N_7140);
xnor U7264 (N_7264,N_7093,N_7135);
xnor U7265 (N_7265,N_7125,N_7110);
xor U7266 (N_7266,N_7055,N_7122);
nor U7267 (N_7267,N_7185,N_7086);
nor U7268 (N_7268,N_7176,N_7160);
and U7269 (N_7269,N_7127,N_7142);
or U7270 (N_7270,N_7173,N_7141);
xnor U7271 (N_7271,N_7059,N_7047);
nand U7272 (N_7272,N_7079,N_7129);
or U7273 (N_7273,N_7165,N_7049);
or U7274 (N_7274,N_7090,N_7179);
or U7275 (N_7275,N_7145,N_7046);
nand U7276 (N_7276,N_7196,N_7199);
or U7277 (N_7277,N_7134,N_7102);
or U7278 (N_7278,N_7120,N_7107);
xnor U7279 (N_7279,N_7136,N_7065);
and U7280 (N_7280,N_7048,N_7160);
and U7281 (N_7281,N_7069,N_7167);
xnor U7282 (N_7282,N_7181,N_7095);
and U7283 (N_7283,N_7172,N_7080);
nand U7284 (N_7284,N_7103,N_7063);
and U7285 (N_7285,N_7125,N_7092);
nor U7286 (N_7286,N_7166,N_7184);
nor U7287 (N_7287,N_7107,N_7068);
and U7288 (N_7288,N_7052,N_7058);
nor U7289 (N_7289,N_7068,N_7183);
nand U7290 (N_7290,N_7159,N_7170);
and U7291 (N_7291,N_7176,N_7173);
or U7292 (N_7292,N_7068,N_7086);
nand U7293 (N_7293,N_7168,N_7049);
nand U7294 (N_7294,N_7096,N_7083);
xor U7295 (N_7295,N_7072,N_7123);
and U7296 (N_7296,N_7096,N_7052);
nand U7297 (N_7297,N_7133,N_7172);
or U7298 (N_7298,N_7045,N_7057);
or U7299 (N_7299,N_7185,N_7063);
and U7300 (N_7300,N_7163,N_7167);
or U7301 (N_7301,N_7133,N_7109);
xor U7302 (N_7302,N_7160,N_7151);
nand U7303 (N_7303,N_7183,N_7189);
xor U7304 (N_7304,N_7100,N_7095);
and U7305 (N_7305,N_7129,N_7176);
xnor U7306 (N_7306,N_7179,N_7081);
nor U7307 (N_7307,N_7083,N_7153);
xor U7308 (N_7308,N_7159,N_7179);
or U7309 (N_7309,N_7112,N_7145);
xnor U7310 (N_7310,N_7183,N_7165);
or U7311 (N_7311,N_7103,N_7155);
or U7312 (N_7312,N_7104,N_7150);
and U7313 (N_7313,N_7162,N_7193);
nand U7314 (N_7314,N_7190,N_7054);
nor U7315 (N_7315,N_7071,N_7147);
xnor U7316 (N_7316,N_7064,N_7130);
and U7317 (N_7317,N_7042,N_7182);
and U7318 (N_7318,N_7122,N_7101);
and U7319 (N_7319,N_7193,N_7158);
and U7320 (N_7320,N_7159,N_7095);
nand U7321 (N_7321,N_7117,N_7096);
or U7322 (N_7322,N_7079,N_7062);
nand U7323 (N_7323,N_7166,N_7056);
and U7324 (N_7324,N_7167,N_7060);
and U7325 (N_7325,N_7088,N_7156);
nand U7326 (N_7326,N_7089,N_7119);
and U7327 (N_7327,N_7194,N_7044);
or U7328 (N_7328,N_7139,N_7190);
or U7329 (N_7329,N_7054,N_7118);
and U7330 (N_7330,N_7198,N_7110);
and U7331 (N_7331,N_7072,N_7191);
and U7332 (N_7332,N_7170,N_7180);
and U7333 (N_7333,N_7135,N_7140);
or U7334 (N_7334,N_7062,N_7168);
nor U7335 (N_7335,N_7052,N_7177);
nand U7336 (N_7336,N_7166,N_7103);
xnor U7337 (N_7337,N_7071,N_7041);
xnor U7338 (N_7338,N_7150,N_7116);
nor U7339 (N_7339,N_7183,N_7057);
or U7340 (N_7340,N_7055,N_7079);
and U7341 (N_7341,N_7158,N_7135);
nand U7342 (N_7342,N_7112,N_7134);
nand U7343 (N_7343,N_7080,N_7152);
xor U7344 (N_7344,N_7167,N_7096);
and U7345 (N_7345,N_7107,N_7117);
xnor U7346 (N_7346,N_7135,N_7091);
nand U7347 (N_7347,N_7190,N_7056);
nor U7348 (N_7348,N_7096,N_7049);
and U7349 (N_7349,N_7138,N_7149);
xnor U7350 (N_7350,N_7190,N_7183);
xor U7351 (N_7351,N_7049,N_7149);
nand U7352 (N_7352,N_7062,N_7098);
or U7353 (N_7353,N_7118,N_7077);
and U7354 (N_7354,N_7172,N_7058);
nand U7355 (N_7355,N_7178,N_7184);
nor U7356 (N_7356,N_7129,N_7077);
nand U7357 (N_7357,N_7178,N_7077);
xnor U7358 (N_7358,N_7139,N_7086);
nor U7359 (N_7359,N_7044,N_7119);
or U7360 (N_7360,N_7356,N_7255);
nand U7361 (N_7361,N_7222,N_7353);
and U7362 (N_7362,N_7221,N_7233);
or U7363 (N_7363,N_7244,N_7266);
and U7364 (N_7364,N_7336,N_7333);
or U7365 (N_7365,N_7298,N_7245);
nand U7366 (N_7366,N_7279,N_7291);
and U7367 (N_7367,N_7345,N_7276);
or U7368 (N_7368,N_7312,N_7268);
and U7369 (N_7369,N_7235,N_7231);
nor U7370 (N_7370,N_7350,N_7224);
or U7371 (N_7371,N_7307,N_7343);
nor U7372 (N_7372,N_7277,N_7220);
xor U7373 (N_7373,N_7346,N_7202);
nand U7374 (N_7374,N_7234,N_7314);
xnor U7375 (N_7375,N_7294,N_7267);
or U7376 (N_7376,N_7299,N_7216);
xor U7377 (N_7377,N_7309,N_7223);
nand U7378 (N_7378,N_7273,N_7200);
and U7379 (N_7379,N_7238,N_7306);
nand U7380 (N_7380,N_7254,N_7349);
and U7381 (N_7381,N_7342,N_7215);
xor U7382 (N_7382,N_7229,N_7219);
and U7383 (N_7383,N_7331,N_7293);
nor U7384 (N_7384,N_7351,N_7317);
xnor U7385 (N_7385,N_7263,N_7227);
xnor U7386 (N_7386,N_7288,N_7329);
xnor U7387 (N_7387,N_7287,N_7205);
and U7388 (N_7388,N_7211,N_7246);
xnor U7389 (N_7389,N_7302,N_7348);
and U7390 (N_7390,N_7247,N_7250);
nand U7391 (N_7391,N_7338,N_7323);
or U7392 (N_7392,N_7284,N_7282);
or U7393 (N_7393,N_7334,N_7337);
xnor U7394 (N_7394,N_7322,N_7259);
nand U7395 (N_7395,N_7249,N_7251);
xor U7396 (N_7396,N_7217,N_7204);
nand U7397 (N_7397,N_7261,N_7327);
and U7398 (N_7398,N_7218,N_7341);
nand U7399 (N_7399,N_7260,N_7280);
or U7400 (N_7400,N_7258,N_7308);
nand U7401 (N_7401,N_7236,N_7328);
and U7402 (N_7402,N_7257,N_7325);
nand U7403 (N_7403,N_7335,N_7315);
xnor U7404 (N_7404,N_7228,N_7283);
or U7405 (N_7405,N_7241,N_7270);
nor U7406 (N_7406,N_7275,N_7303);
nor U7407 (N_7407,N_7262,N_7237);
nand U7408 (N_7408,N_7340,N_7278);
xor U7409 (N_7409,N_7347,N_7212);
nor U7410 (N_7410,N_7296,N_7264);
or U7411 (N_7411,N_7300,N_7344);
or U7412 (N_7412,N_7256,N_7316);
or U7413 (N_7413,N_7326,N_7214);
nor U7414 (N_7414,N_7239,N_7285);
and U7415 (N_7415,N_7355,N_7324);
nand U7416 (N_7416,N_7269,N_7208);
nor U7417 (N_7417,N_7359,N_7292);
nand U7418 (N_7418,N_7265,N_7318);
and U7419 (N_7419,N_7332,N_7248);
and U7420 (N_7420,N_7330,N_7274);
or U7421 (N_7421,N_7242,N_7310);
nand U7422 (N_7422,N_7321,N_7295);
nor U7423 (N_7423,N_7313,N_7207);
and U7424 (N_7424,N_7290,N_7281);
or U7425 (N_7425,N_7304,N_7253);
xnor U7426 (N_7426,N_7209,N_7301);
or U7427 (N_7427,N_7203,N_7210);
nor U7428 (N_7428,N_7225,N_7354);
and U7429 (N_7429,N_7230,N_7358);
and U7430 (N_7430,N_7297,N_7201);
nor U7431 (N_7431,N_7289,N_7232);
and U7432 (N_7432,N_7243,N_7213);
or U7433 (N_7433,N_7286,N_7240);
nand U7434 (N_7434,N_7305,N_7311);
nand U7435 (N_7435,N_7226,N_7357);
xor U7436 (N_7436,N_7252,N_7206);
xor U7437 (N_7437,N_7271,N_7352);
and U7438 (N_7438,N_7320,N_7339);
and U7439 (N_7439,N_7319,N_7272);
or U7440 (N_7440,N_7230,N_7305);
nor U7441 (N_7441,N_7249,N_7283);
nand U7442 (N_7442,N_7297,N_7286);
xnor U7443 (N_7443,N_7280,N_7276);
xor U7444 (N_7444,N_7201,N_7335);
nor U7445 (N_7445,N_7227,N_7232);
xor U7446 (N_7446,N_7262,N_7250);
and U7447 (N_7447,N_7330,N_7283);
xor U7448 (N_7448,N_7323,N_7274);
nor U7449 (N_7449,N_7226,N_7205);
nand U7450 (N_7450,N_7225,N_7262);
nand U7451 (N_7451,N_7295,N_7234);
or U7452 (N_7452,N_7346,N_7200);
nand U7453 (N_7453,N_7206,N_7319);
or U7454 (N_7454,N_7295,N_7267);
nand U7455 (N_7455,N_7307,N_7207);
xnor U7456 (N_7456,N_7245,N_7286);
or U7457 (N_7457,N_7226,N_7208);
nand U7458 (N_7458,N_7311,N_7231);
nor U7459 (N_7459,N_7256,N_7317);
xor U7460 (N_7460,N_7316,N_7236);
xor U7461 (N_7461,N_7324,N_7330);
or U7462 (N_7462,N_7202,N_7277);
and U7463 (N_7463,N_7240,N_7304);
nand U7464 (N_7464,N_7263,N_7276);
nand U7465 (N_7465,N_7264,N_7302);
xor U7466 (N_7466,N_7294,N_7291);
nand U7467 (N_7467,N_7285,N_7225);
and U7468 (N_7468,N_7256,N_7204);
xor U7469 (N_7469,N_7278,N_7322);
xor U7470 (N_7470,N_7321,N_7252);
xor U7471 (N_7471,N_7267,N_7276);
or U7472 (N_7472,N_7349,N_7253);
or U7473 (N_7473,N_7334,N_7209);
xor U7474 (N_7474,N_7257,N_7223);
nand U7475 (N_7475,N_7331,N_7253);
nand U7476 (N_7476,N_7237,N_7318);
xnor U7477 (N_7477,N_7316,N_7289);
and U7478 (N_7478,N_7232,N_7359);
nor U7479 (N_7479,N_7306,N_7334);
nor U7480 (N_7480,N_7235,N_7218);
and U7481 (N_7481,N_7323,N_7355);
or U7482 (N_7482,N_7359,N_7343);
nand U7483 (N_7483,N_7224,N_7296);
nor U7484 (N_7484,N_7300,N_7248);
or U7485 (N_7485,N_7281,N_7354);
and U7486 (N_7486,N_7326,N_7262);
xnor U7487 (N_7487,N_7217,N_7201);
nor U7488 (N_7488,N_7208,N_7222);
nor U7489 (N_7489,N_7265,N_7229);
or U7490 (N_7490,N_7211,N_7339);
or U7491 (N_7491,N_7312,N_7324);
or U7492 (N_7492,N_7240,N_7337);
nor U7493 (N_7493,N_7310,N_7229);
and U7494 (N_7494,N_7297,N_7240);
xnor U7495 (N_7495,N_7305,N_7303);
nand U7496 (N_7496,N_7359,N_7289);
or U7497 (N_7497,N_7239,N_7301);
xor U7498 (N_7498,N_7261,N_7242);
nand U7499 (N_7499,N_7279,N_7265);
xnor U7500 (N_7500,N_7318,N_7321);
or U7501 (N_7501,N_7211,N_7203);
nor U7502 (N_7502,N_7359,N_7287);
nand U7503 (N_7503,N_7245,N_7237);
or U7504 (N_7504,N_7267,N_7343);
or U7505 (N_7505,N_7323,N_7347);
xor U7506 (N_7506,N_7278,N_7262);
nand U7507 (N_7507,N_7267,N_7217);
nor U7508 (N_7508,N_7226,N_7209);
nor U7509 (N_7509,N_7301,N_7272);
nor U7510 (N_7510,N_7270,N_7231);
xor U7511 (N_7511,N_7267,N_7229);
or U7512 (N_7512,N_7281,N_7231);
nor U7513 (N_7513,N_7200,N_7332);
xnor U7514 (N_7514,N_7328,N_7264);
and U7515 (N_7515,N_7234,N_7239);
nor U7516 (N_7516,N_7317,N_7328);
xor U7517 (N_7517,N_7316,N_7330);
nand U7518 (N_7518,N_7337,N_7287);
xnor U7519 (N_7519,N_7249,N_7301);
or U7520 (N_7520,N_7389,N_7412);
xor U7521 (N_7521,N_7395,N_7436);
xor U7522 (N_7522,N_7509,N_7388);
nand U7523 (N_7523,N_7478,N_7433);
and U7524 (N_7524,N_7380,N_7425);
and U7525 (N_7525,N_7367,N_7508);
xor U7526 (N_7526,N_7443,N_7365);
xnor U7527 (N_7527,N_7427,N_7360);
or U7528 (N_7528,N_7470,N_7453);
xnor U7529 (N_7529,N_7454,N_7485);
nand U7530 (N_7530,N_7421,N_7446);
or U7531 (N_7531,N_7500,N_7384);
or U7532 (N_7532,N_7396,N_7397);
nand U7533 (N_7533,N_7456,N_7448);
nand U7534 (N_7534,N_7410,N_7383);
xnor U7535 (N_7535,N_7392,N_7512);
nor U7536 (N_7536,N_7375,N_7484);
nor U7537 (N_7537,N_7420,N_7471);
nor U7538 (N_7538,N_7435,N_7428);
or U7539 (N_7539,N_7422,N_7404);
or U7540 (N_7540,N_7407,N_7477);
or U7541 (N_7541,N_7489,N_7403);
nand U7542 (N_7542,N_7400,N_7447);
nand U7543 (N_7543,N_7487,N_7439);
or U7544 (N_7544,N_7501,N_7363);
and U7545 (N_7545,N_7473,N_7513);
and U7546 (N_7546,N_7494,N_7515);
nor U7547 (N_7547,N_7480,N_7475);
and U7548 (N_7548,N_7462,N_7458);
and U7549 (N_7549,N_7492,N_7419);
and U7550 (N_7550,N_7370,N_7503);
nand U7551 (N_7551,N_7393,N_7430);
nor U7552 (N_7552,N_7382,N_7387);
and U7553 (N_7553,N_7364,N_7399);
xnor U7554 (N_7554,N_7426,N_7416);
xnor U7555 (N_7555,N_7413,N_7423);
nor U7556 (N_7556,N_7381,N_7459);
nand U7557 (N_7557,N_7402,N_7451);
nand U7558 (N_7558,N_7479,N_7468);
and U7559 (N_7559,N_7372,N_7408);
nand U7560 (N_7560,N_7371,N_7409);
xnor U7561 (N_7561,N_7418,N_7432);
and U7562 (N_7562,N_7502,N_7376);
xor U7563 (N_7563,N_7449,N_7398);
or U7564 (N_7564,N_7505,N_7514);
xor U7565 (N_7565,N_7411,N_7431);
xor U7566 (N_7566,N_7424,N_7401);
xnor U7567 (N_7567,N_7390,N_7438);
nand U7568 (N_7568,N_7474,N_7497);
xnor U7569 (N_7569,N_7499,N_7429);
xnor U7570 (N_7570,N_7414,N_7440);
nor U7571 (N_7571,N_7482,N_7444);
nor U7572 (N_7572,N_7461,N_7361);
xnor U7573 (N_7573,N_7434,N_7394);
xor U7574 (N_7574,N_7483,N_7507);
nand U7575 (N_7575,N_7460,N_7374);
and U7576 (N_7576,N_7493,N_7465);
or U7577 (N_7577,N_7441,N_7377);
xnor U7578 (N_7578,N_7516,N_7415);
and U7579 (N_7579,N_7467,N_7486);
nand U7580 (N_7580,N_7504,N_7442);
and U7581 (N_7581,N_7455,N_7373);
nand U7582 (N_7582,N_7405,N_7391);
or U7583 (N_7583,N_7406,N_7457);
and U7584 (N_7584,N_7506,N_7437);
nand U7585 (N_7585,N_7495,N_7379);
or U7586 (N_7586,N_7481,N_7510);
and U7587 (N_7587,N_7452,N_7496);
or U7588 (N_7588,N_7366,N_7386);
nor U7589 (N_7589,N_7472,N_7469);
nor U7590 (N_7590,N_7385,N_7519);
nor U7591 (N_7591,N_7498,N_7476);
and U7592 (N_7592,N_7488,N_7378);
or U7593 (N_7593,N_7417,N_7369);
nor U7594 (N_7594,N_7466,N_7362);
and U7595 (N_7595,N_7450,N_7517);
or U7596 (N_7596,N_7368,N_7511);
nand U7597 (N_7597,N_7445,N_7491);
or U7598 (N_7598,N_7490,N_7464);
and U7599 (N_7599,N_7463,N_7518);
or U7600 (N_7600,N_7393,N_7426);
or U7601 (N_7601,N_7426,N_7386);
nand U7602 (N_7602,N_7473,N_7471);
and U7603 (N_7603,N_7429,N_7386);
nand U7604 (N_7604,N_7395,N_7519);
xor U7605 (N_7605,N_7491,N_7449);
nand U7606 (N_7606,N_7464,N_7497);
nand U7607 (N_7607,N_7380,N_7455);
nand U7608 (N_7608,N_7420,N_7430);
nand U7609 (N_7609,N_7407,N_7452);
and U7610 (N_7610,N_7361,N_7372);
xnor U7611 (N_7611,N_7486,N_7390);
nor U7612 (N_7612,N_7477,N_7400);
nor U7613 (N_7613,N_7377,N_7402);
and U7614 (N_7614,N_7438,N_7458);
nor U7615 (N_7615,N_7467,N_7435);
nor U7616 (N_7616,N_7517,N_7369);
and U7617 (N_7617,N_7363,N_7389);
or U7618 (N_7618,N_7503,N_7470);
and U7619 (N_7619,N_7393,N_7479);
xor U7620 (N_7620,N_7413,N_7396);
xnor U7621 (N_7621,N_7487,N_7382);
xnor U7622 (N_7622,N_7402,N_7403);
nor U7623 (N_7623,N_7509,N_7478);
nand U7624 (N_7624,N_7466,N_7380);
nor U7625 (N_7625,N_7482,N_7426);
nand U7626 (N_7626,N_7485,N_7401);
nor U7627 (N_7627,N_7442,N_7398);
or U7628 (N_7628,N_7482,N_7468);
nor U7629 (N_7629,N_7476,N_7387);
or U7630 (N_7630,N_7402,N_7391);
nand U7631 (N_7631,N_7464,N_7491);
nor U7632 (N_7632,N_7374,N_7372);
xnor U7633 (N_7633,N_7450,N_7393);
or U7634 (N_7634,N_7416,N_7398);
or U7635 (N_7635,N_7398,N_7381);
xnor U7636 (N_7636,N_7420,N_7443);
nor U7637 (N_7637,N_7384,N_7422);
and U7638 (N_7638,N_7392,N_7453);
xor U7639 (N_7639,N_7396,N_7372);
and U7640 (N_7640,N_7473,N_7511);
and U7641 (N_7641,N_7483,N_7445);
nor U7642 (N_7642,N_7467,N_7501);
or U7643 (N_7643,N_7364,N_7480);
or U7644 (N_7644,N_7363,N_7513);
nor U7645 (N_7645,N_7403,N_7442);
nand U7646 (N_7646,N_7453,N_7505);
and U7647 (N_7647,N_7407,N_7476);
and U7648 (N_7648,N_7433,N_7364);
nor U7649 (N_7649,N_7383,N_7449);
nor U7650 (N_7650,N_7377,N_7373);
or U7651 (N_7651,N_7406,N_7391);
and U7652 (N_7652,N_7481,N_7373);
and U7653 (N_7653,N_7407,N_7421);
and U7654 (N_7654,N_7494,N_7498);
nor U7655 (N_7655,N_7429,N_7445);
xnor U7656 (N_7656,N_7445,N_7424);
nor U7657 (N_7657,N_7368,N_7378);
nand U7658 (N_7658,N_7492,N_7390);
and U7659 (N_7659,N_7457,N_7461);
xor U7660 (N_7660,N_7410,N_7445);
and U7661 (N_7661,N_7447,N_7508);
and U7662 (N_7662,N_7475,N_7516);
xnor U7663 (N_7663,N_7473,N_7470);
nand U7664 (N_7664,N_7396,N_7471);
nor U7665 (N_7665,N_7518,N_7433);
and U7666 (N_7666,N_7493,N_7425);
and U7667 (N_7667,N_7397,N_7364);
nand U7668 (N_7668,N_7364,N_7379);
and U7669 (N_7669,N_7424,N_7463);
and U7670 (N_7670,N_7429,N_7403);
and U7671 (N_7671,N_7485,N_7451);
nand U7672 (N_7672,N_7495,N_7387);
nand U7673 (N_7673,N_7368,N_7468);
nand U7674 (N_7674,N_7446,N_7465);
nor U7675 (N_7675,N_7441,N_7470);
or U7676 (N_7676,N_7420,N_7489);
xnor U7677 (N_7677,N_7442,N_7469);
nor U7678 (N_7678,N_7431,N_7438);
and U7679 (N_7679,N_7443,N_7360);
xor U7680 (N_7680,N_7600,N_7586);
and U7681 (N_7681,N_7593,N_7671);
nor U7682 (N_7682,N_7634,N_7532);
or U7683 (N_7683,N_7540,N_7596);
and U7684 (N_7684,N_7618,N_7584);
nor U7685 (N_7685,N_7614,N_7580);
or U7686 (N_7686,N_7533,N_7642);
xnor U7687 (N_7687,N_7590,N_7635);
and U7688 (N_7688,N_7660,N_7655);
and U7689 (N_7689,N_7672,N_7613);
nor U7690 (N_7690,N_7581,N_7645);
and U7691 (N_7691,N_7551,N_7530);
nand U7692 (N_7692,N_7619,N_7542);
or U7693 (N_7693,N_7572,N_7569);
xnor U7694 (N_7694,N_7534,N_7641);
nor U7695 (N_7695,N_7675,N_7562);
and U7696 (N_7696,N_7624,N_7563);
and U7697 (N_7697,N_7541,N_7663);
xor U7698 (N_7698,N_7667,N_7571);
or U7699 (N_7699,N_7610,N_7656);
nand U7700 (N_7700,N_7545,N_7529);
nor U7701 (N_7701,N_7676,N_7623);
or U7702 (N_7702,N_7615,N_7579);
or U7703 (N_7703,N_7668,N_7520);
and U7704 (N_7704,N_7664,N_7604);
xor U7705 (N_7705,N_7621,N_7670);
nand U7706 (N_7706,N_7538,N_7564);
nand U7707 (N_7707,N_7555,N_7574);
nor U7708 (N_7708,N_7612,N_7666);
and U7709 (N_7709,N_7561,N_7547);
xnor U7710 (N_7710,N_7558,N_7679);
nor U7711 (N_7711,N_7611,N_7657);
and U7712 (N_7712,N_7554,N_7594);
nor U7713 (N_7713,N_7662,N_7626);
or U7714 (N_7714,N_7616,N_7552);
and U7715 (N_7715,N_7560,N_7539);
nor U7716 (N_7716,N_7633,N_7628);
nand U7717 (N_7717,N_7591,N_7627);
and U7718 (N_7718,N_7567,N_7557);
nor U7719 (N_7719,N_7531,N_7526);
nor U7720 (N_7720,N_7559,N_7592);
xor U7721 (N_7721,N_7622,N_7654);
nand U7722 (N_7722,N_7661,N_7602);
and U7723 (N_7723,N_7608,N_7648);
and U7724 (N_7724,N_7605,N_7639);
or U7725 (N_7725,N_7638,N_7588);
and U7726 (N_7726,N_7548,N_7636);
xnor U7727 (N_7727,N_7550,N_7603);
nand U7728 (N_7728,N_7543,N_7523);
nor U7729 (N_7729,N_7637,N_7598);
or U7730 (N_7730,N_7631,N_7524);
xnor U7731 (N_7731,N_7599,N_7646);
xor U7732 (N_7732,N_7528,N_7544);
and U7733 (N_7733,N_7620,N_7658);
xor U7734 (N_7734,N_7647,N_7607);
or U7735 (N_7735,N_7632,N_7578);
and U7736 (N_7736,N_7625,N_7650);
nand U7737 (N_7737,N_7653,N_7665);
and U7738 (N_7738,N_7643,N_7577);
and U7739 (N_7739,N_7573,N_7549);
nor U7740 (N_7740,N_7630,N_7649);
nand U7741 (N_7741,N_7570,N_7587);
or U7742 (N_7742,N_7575,N_7673);
xor U7743 (N_7743,N_7566,N_7651);
or U7744 (N_7744,N_7585,N_7522);
nor U7745 (N_7745,N_7659,N_7576);
nor U7746 (N_7746,N_7644,N_7674);
nor U7747 (N_7747,N_7582,N_7553);
nor U7748 (N_7748,N_7536,N_7617);
or U7749 (N_7749,N_7527,N_7565);
and U7750 (N_7750,N_7546,N_7537);
and U7751 (N_7751,N_7609,N_7669);
xnor U7752 (N_7752,N_7595,N_7525);
or U7753 (N_7753,N_7601,N_7521);
nor U7754 (N_7754,N_7606,N_7677);
nor U7755 (N_7755,N_7589,N_7629);
nor U7756 (N_7756,N_7568,N_7583);
xor U7757 (N_7757,N_7535,N_7678);
and U7758 (N_7758,N_7597,N_7556);
and U7759 (N_7759,N_7652,N_7640);
or U7760 (N_7760,N_7661,N_7662);
nor U7761 (N_7761,N_7663,N_7553);
xor U7762 (N_7762,N_7628,N_7569);
nand U7763 (N_7763,N_7607,N_7638);
xnor U7764 (N_7764,N_7557,N_7627);
and U7765 (N_7765,N_7656,N_7595);
or U7766 (N_7766,N_7585,N_7587);
nor U7767 (N_7767,N_7672,N_7615);
nand U7768 (N_7768,N_7589,N_7543);
nand U7769 (N_7769,N_7524,N_7627);
or U7770 (N_7770,N_7618,N_7586);
or U7771 (N_7771,N_7546,N_7523);
nor U7772 (N_7772,N_7522,N_7576);
nand U7773 (N_7773,N_7552,N_7664);
xnor U7774 (N_7774,N_7591,N_7618);
xor U7775 (N_7775,N_7677,N_7648);
or U7776 (N_7776,N_7639,N_7541);
and U7777 (N_7777,N_7639,N_7524);
and U7778 (N_7778,N_7649,N_7563);
or U7779 (N_7779,N_7547,N_7564);
xor U7780 (N_7780,N_7595,N_7631);
and U7781 (N_7781,N_7545,N_7602);
xnor U7782 (N_7782,N_7650,N_7581);
or U7783 (N_7783,N_7544,N_7561);
nand U7784 (N_7784,N_7642,N_7605);
nor U7785 (N_7785,N_7666,N_7542);
nor U7786 (N_7786,N_7596,N_7603);
and U7787 (N_7787,N_7656,N_7630);
nand U7788 (N_7788,N_7672,N_7609);
xnor U7789 (N_7789,N_7602,N_7568);
nand U7790 (N_7790,N_7538,N_7600);
xnor U7791 (N_7791,N_7655,N_7574);
nand U7792 (N_7792,N_7660,N_7565);
and U7793 (N_7793,N_7545,N_7596);
nor U7794 (N_7794,N_7548,N_7589);
xnor U7795 (N_7795,N_7656,N_7632);
and U7796 (N_7796,N_7529,N_7597);
and U7797 (N_7797,N_7602,N_7594);
and U7798 (N_7798,N_7598,N_7678);
nor U7799 (N_7799,N_7581,N_7635);
and U7800 (N_7800,N_7632,N_7582);
nand U7801 (N_7801,N_7616,N_7639);
or U7802 (N_7802,N_7558,N_7672);
xnor U7803 (N_7803,N_7641,N_7586);
nand U7804 (N_7804,N_7641,N_7632);
and U7805 (N_7805,N_7652,N_7613);
or U7806 (N_7806,N_7572,N_7646);
or U7807 (N_7807,N_7611,N_7636);
and U7808 (N_7808,N_7576,N_7580);
and U7809 (N_7809,N_7557,N_7552);
xnor U7810 (N_7810,N_7544,N_7594);
nor U7811 (N_7811,N_7555,N_7583);
nand U7812 (N_7812,N_7666,N_7569);
xnor U7813 (N_7813,N_7559,N_7670);
and U7814 (N_7814,N_7630,N_7629);
and U7815 (N_7815,N_7603,N_7673);
nand U7816 (N_7816,N_7630,N_7581);
and U7817 (N_7817,N_7663,N_7542);
nor U7818 (N_7818,N_7592,N_7652);
nand U7819 (N_7819,N_7601,N_7675);
or U7820 (N_7820,N_7615,N_7618);
or U7821 (N_7821,N_7536,N_7633);
nor U7822 (N_7822,N_7567,N_7610);
nand U7823 (N_7823,N_7529,N_7535);
and U7824 (N_7824,N_7583,N_7547);
nand U7825 (N_7825,N_7612,N_7527);
nand U7826 (N_7826,N_7583,N_7587);
and U7827 (N_7827,N_7642,N_7568);
or U7828 (N_7828,N_7671,N_7565);
nor U7829 (N_7829,N_7526,N_7580);
nor U7830 (N_7830,N_7591,N_7675);
nor U7831 (N_7831,N_7664,N_7527);
and U7832 (N_7832,N_7583,N_7664);
nand U7833 (N_7833,N_7633,N_7602);
or U7834 (N_7834,N_7618,N_7585);
and U7835 (N_7835,N_7678,N_7577);
nand U7836 (N_7836,N_7662,N_7609);
nand U7837 (N_7837,N_7542,N_7559);
and U7838 (N_7838,N_7577,N_7535);
or U7839 (N_7839,N_7614,N_7597);
nand U7840 (N_7840,N_7796,N_7832);
or U7841 (N_7841,N_7730,N_7792);
xnor U7842 (N_7842,N_7761,N_7815);
and U7843 (N_7843,N_7797,N_7738);
xor U7844 (N_7844,N_7803,N_7691);
and U7845 (N_7845,N_7734,N_7784);
xor U7846 (N_7846,N_7723,N_7735);
nor U7847 (N_7847,N_7726,N_7813);
nor U7848 (N_7848,N_7682,N_7766);
or U7849 (N_7849,N_7810,N_7789);
xnor U7850 (N_7850,N_7748,N_7839);
xnor U7851 (N_7851,N_7764,N_7768);
and U7852 (N_7852,N_7747,N_7785);
or U7853 (N_7853,N_7685,N_7760);
nand U7854 (N_7854,N_7774,N_7772);
nor U7855 (N_7855,N_7838,N_7762);
or U7856 (N_7856,N_7802,N_7782);
or U7857 (N_7857,N_7756,N_7758);
and U7858 (N_7858,N_7688,N_7806);
nand U7859 (N_7859,N_7777,N_7709);
or U7860 (N_7860,N_7821,N_7720);
or U7861 (N_7861,N_7719,N_7713);
xnor U7862 (N_7862,N_7716,N_7739);
or U7863 (N_7863,N_7827,N_7835);
xnor U7864 (N_7864,N_7805,N_7696);
nand U7865 (N_7865,N_7717,N_7740);
nor U7866 (N_7866,N_7697,N_7795);
nor U7867 (N_7867,N_7771,N_7819);
xor U7868 (N_7868,N_7725,N_7822);
and U7869 (N_7869,N_7800,N_7718);
nor U7870 (N_7870,N_7829,N_7715);
xnor U7871 (N_7871,N_7729,N_7763);
and U7872 (N_7872,N_7834,N_7828);
nor U7873 (N_7873,N_7831,N_7698);
or U7874 (N_7874,N_7707,N_7799);
nand U7875 (N_7875,N_7769,N_7750);
or U7876 (N_7876,N_7686,N_7701);
or U7877 (N_7877,N_7692,N_7775);
nand U7878 (N_7878,N_7733,N_7779);
or U7879 (N_7879,N_7804,N_7703);
nand U7880 (N_7880,N_7817,N_7783);
or U7881 (N_7881,N_7780,N_7753);
xor U7882 (N_7882,N_7830,N_7773);
or U7883 (N_7883,N_7745,N_7714);
xor U7884 (N_7884,N_7711,N_7743);
nand U7885 (N_7885,N_7825,N_7757);
xor U7886 (N_7886,N_7798,N_7728);
nor U7887 (N_7887,N_7808,N_7749);
nand U7888 (N_7888,N_7681,N_7801);
nor U7889 (N_7889,N_7684,N_7793);
xnor U7890 (N_7890,N_7765,N_7820);
or U7891 (N_7891,N_7823,N_7695);
nor U7892 (N_7892,N_7741,N_7818);
or U7893 (N_7893,N_7754,N_7755);
nand U7894 (N_7894,N_7816,N_7732);
and U7895 (N_7895,N_7787,N_7699);
nor U7896 (N_7896,N_7778,N_7693);
xnor U7897 (N_7897,N_7708,N_7700);
nand U7898 (N_7898,N_7812,N_7710);
or U7899 (N_7899,N_7833,N_7702);
xnor U7900 (N_7900,N_7724,N_7683);
nand U7901 (N_7901,N_7786,N_7704);
nand U7902 (N_7902,N_7788,N_7731);
xor U7903 (N_7903,N_7790,N_7837);
nor U7904 (N_7904,N_7687,N_7744);
nor U7905 (N_7905,N_7737,N_7705);
or U7906 (N_7906,N_7722,N_7824);
or U7907 (N_7907,N_7807,N_7742);
nor U7908 (N_7908,N_7809,N_7712);
nand U7909 (N_7909,N_7770,N_7781);
xnor U7910 (N_7910,N_7694,N_7791);
nor U7911 (N_7911,N_7814,N_7836);
and U7912 (N_7912,N_7752,N_7736);
nor U7913 (N_7913,N_7794,N_7680);
nand U7914 (N_7914,N_7826,N_7721);
xor U7915 (N_7915,N_7767,N_7689);
xnor U7916 (N_7916,N_7727,N_7706);
nand U7917 (N_7917,N_7746,N_7751);
or U7918 (N_7918,N_7759,N_7690);
or U7919 (N_7919,N_7811,N_7776);
xnor U7920 (N_7920,N_7705,N_7787);
and U7921 (N_7921,N_7771,N_7770);
xor U7922 (N_7922,N_7830,N_7796);
and U7923 (N_7923,N_7746,N_7814);
or U7924 (N_7924,N_7817,N_7699);
nand U7925 (N_7925,N_7816,N_7742);
xor U7926 (N_7926,N_7791,N_7745);
or U7927 (N_7927,N_7695,N_7803);
nor U7928 (N_7928,N_7775,N_7689);
nor U7929 (N_7929,N_7728,N_7770);
xor U7930 (N_7930,N_7693,N_7838);
nand U7931 (N_7931,N_7712,N_7810);
nor U7932 (N_7932,N_7754,N_7685);
and U7933 (N_7933,N_7737,N_7709);
nand U7934 (N_7934,N_7801,N_7827);
xor U7935 (N_7935,N_7741,N_7776);
or U7936 (N_7936,N_7776,N_7683);
nor U7937 (N_7937,N_7711,N_7724);
nand U7938 (N_7938,N_7701,N_7721);
xnor U7939 (N_7939,N_7837,N_7762);
and U7940 (N_7940,N_7767,N_7810);
and U7941 (N_7941,N_7822,N_7837);
xor U7942 (N_7942,N_7707,N_7829);
or U7943 (N_7943,N_7772,N_7700);
and U7944 (N_7944,N_7729,N_7826);
xor U7945 (N_7945,N_7831,N_7814);
nand U7946 (N_7946,N_7763,N_7828);
and U7947 (N_7947,N_7741,N_7822);
and U7948 (N_7948,N_7781,N_7833);
or U7949 (N_7949,N_7709,N_7747);
nor U7950 (N_7950,N_7782,N_7821);
or U7951 (N_7951,N_7778,N_7762);
nand U7952 (N_7952,N_7781,N_7828);
xnor U7953 (N_7953,N_7813,N_7717);
xnor U7954 (N_7954,N_7792,N_7688);
xor U7955 (N_7955,N_7692,N_7810);
and U7956 (N_7956,N_7806,N_7732);
nand U7957 (N_7957,N_7744,N_7681);
and U7958 (N_7958,N_7684,N_7755);
or U7959 (N_7959,N_7706,N_7745);
nand U7960 (N_7960,N_7701,N_7773);
and U7961 (N_7961,N_7814,N_7749);
xor U7962 (N_7962,N_7789,N_7773);
and U7963 (N_7963,N_7778,N_7793);
or U7964 (N_7964,N_7786,N_7727);
nand U7965 (N_7965,N_7748,N_7781);
xnor U7966 (N_7966,N_7803,N_7704);
and U7967 (N_7967,N_7703,N_7751);
nor U7968 (N_7968,N_7820,N_7782);
or U7969 (N_7969,N_7697,N_7823);
nand U7970 (N_7970,N_7795,N_7782);
nand U7971 (N_7971,N_7801,N_7803);
nor U7972 (N_7972,N_7826,N_7776);
and U7973 (N_7973,N_7820,N_7812);
or U7974 (N_7974,N_7721,N_7811);
and U7975 (N_7975,N_7832,N_7830);
nor U7976 (N_7976,N_7711,N_7740);
nand U7977 (N_7977,N_7713,N_7689);
nand U7978 (N_7978,N_7736,N_7813);
nand U7979 (N_7979,N_7780,N_7688);
xnor U7980 (N_7980,N_7811,N_7681);
or U7981 (N_7981,N_7684,N_7762);
xor U7982 (N_7982,N_7739,N_7740);
nor U7983 (N_7983,N_7718,N_7814);
nand U7984 (N_7984,N_7702,N_7726);
nor U7985 (N_7985,N_7751,N_7802);
and U7986 (N_7986,N_7750,N_7779);
nor U7987 (N_7987,N_7835,N_7686);
or U7988 (N_7988,N_7804,N_7811);
nor U7989 (N_7989,N_7700,N_7691);
nand U7990 (N_7990,N_7818,N_7762);
nor U7991 (N_7991,N_7708,N_7764);
nand U7992 (N_7992,N_7834,N_7722);
xor U7993 (N_7993,N_7753,N_7771);
nand U7994 (N_7994,N_7799,N_7791);
or U7995 (N_7995,N_7813,N_7801);
nand U7996 (N_7996,N_7785,N_7816);
and U7997 (N_7997,N_7773,N_7750);
and U7998 (N_7998,N_7684,N_7716);
and U7999 (N_7999,N_7821,N_7775);
or U8000 (N_8000,N_7937,N_7992);
xnor U8001 (N_8001,N_7935,N_7892);
xor U8002 (N_8002,N_7952,N_7915);
nor U8003 (N_8003,N_7862,N_7972);
and U8004 (N_8004,N_7923,N_7857);
nor U8005 (N_8005,N_7850,N_7906);
nand U8006 (N_8006,N_7842,N_7844);
xnor U8007 (N_8007,N_7948,N_7887);
nor U8008 (N_8008,N_7910,N_7969);
nand U8009 (N_8009,N_7851,N_7918);
nand U8010 (N_8010,N_7947,N_7954);
and U8011 (N_8011,N_7977,N_7990);
and U8012 (N_8012,N_7919,N_7939);
and U8013 (N_8013,N_7934,N_7973);
nand U8014 (N_8014,N_7994,N_7998);
and U8015 (N_8015,N_7908,N_7840);
nand U8016 (N_8016,N_7894,N_7925);
nand U8017 (N_8017,N_7896,N_7905);
and U8018 (N_8018,N_7921,N_7980);
or U8019 (N_8019,N_7997,N_7899);
or U8020 (N_8020,N_7922,N_7875);
nor U8021 (N_8021,N_7983,N_7995);
nand U8022 (N_8022,N_7962,N_7932);
and U8023 (N_8023,N_7984,N_7903);
and U8024 (N_8024,N_7871,N_7889);
and U8025 (N_8025,N_7938,N_7946);
nor U8026 (N_8026,N_7907,N_7898);
xnor U8027 (N_8027,N_7970,N_7913);
xor U8028 (N_8028,N_7988,N_7869);
nand U8029 (N_8029,N_7927,N_7863);
xor U8030 (N_8030,N_7859,N_7979);
nand U8031 (N_8031,N_7885,N_7858);
xnor U8032 (N_8032,N_7928,N_7936);
and U8033 (N_8033,N_7971,N_7901);
xor U8034 (N_8034,N_7843,N_7877);
or U8035 (N_8035,N_7909,N_7880);
xnor U8036 (N_8036,N_7968,N_7849);
xor U8037 (N_8037,N_7895,N_7974);
xnor U8038 (N_8038,N_7860,N_7867);
or U8039 (N_8039,N_7848,N_7949);
xnor U8040 (N_8040,N_7855,N_7941);
nand U8041 (N_8041,N_7961,N_7940);
nor U8042 (N_8042,N_7965,N_7986);
and U8043 (N_8043,N_7917,N_7847);
or U8044 (N_8044,N_7856,N_7882);
xor U8045 (N_8045,N_7841,N_7886);
nor U8046 (N_8046,N_7866,N_7993);
and U8047 (N_8047,N_7964,N_7879);
nand U8048 (N_8048,N_7924,N_7951);
nand U8049 (N_8049,N_7874,N_7981);
xor U8050 (N_8050,N_7991,N_7904);
xnor U8051 (N_8051,N_7897,N_7891);
nand U8052 (N_8052,N_7865,N_7942);
nor U8053 (N_8053,N_7955,N_7890);
or U8054 (N_8054,N_7999,N_7873);
nor U8055 (N_8055,N_7945,N_7933);
xnor U8056 (N_8056,N_7912,N_7846);
nor U8057 (N_8057,N_7956,N_7916);
and U8058 (N_8058,N_7868,N_7845);
and U8059 (N_8059,N_7920,N_7931);
nand U8060 (N_8060,N_7958,N_7930);
xor U8061 (N_8061,N_7987,N_7989);
nand U8062 (N_8062,N_7854,N_7985);
nor U8063 (N_8063,N_7976,N_7953);
nor U8064 (N_8064,N_7950,N_7878);
xor U8065 (N_8065,N_7963,N_7914);
and U8066 (N_8066,N_7876,N_7883);
nor U8067 (N_8067,N_7929,N_7870);
nand U8068 (N_8068,N_7943,N_7966);
nor U8069 (N_8069,N_7893,N_7902);
and U8070 (N_8070,N_7881,N_7982);
nor U8071 (N_8071,N_7911,N_7861);
nand U8072 (N_8072,N_7960,N_7852);
xor U8073 (N_8073,N_7884,N_7957);
nand U8074 (N_8074,N_7959,N_7853);
and U8075 (N_8075,N_7996,N_7975);
xor U8076 (N_8076,N_7872,N_7864);
nand U8077 (N_8077,N_7900,N_7978);
nand U8078 (N_8078,N_7944,N_7926);
nand U8079 (N_8079,N_7888,N_7967);
and U8080 (N_8080,N_7996,N_7974);
nor U8081 (N_8081,N_7937,N_7954);
nand U8082 (N_8082,N_7971,N_7934);
nor U8083 (N_8083,N_7857,N_7968);
or U8084 (N_8084,N_7944,N_7923);
xnor U8085 (N_8085,N_7873,N_7872);
or U8086 (N_8086,N_7890,N_7850);
nor U8087 (N_8087,N_7912,N_7868);
and U8088 (N_8088,N_7902,N_7969);
and U8089 (N_8089,N_7911,N_7893);
xnor U8090 (N_8090,N_7875,N_7970);
nand U8091 (N_8091,N_7863,N_7958);
nor U8092 (N_8092,N_7991,N_7984);
nor U8093 (N_8093,N_7875,N_7937);
and U8094 (N_8094,N_7863,N_7911);
nand U8095 (N_8095,N_7893,N_7845);
xor U8096 (N_8096,N_7916,N_7962);
nor U8097 (N_8097,N_7958,N_7931);
nor U8098 (N_8098,N_7843,N_7853);
xor U8099 (N_8099,N_7982,N_7971);
nor U8100 (N_8100,N_7882,N_7991);
xor U8101 (N_8101,N_7975,N_7903);
nand U8102 (N_8102,N_7890,N_7880);
nand U8103 (N_8103,N_7941,N_7876);
nor U8104 (N_8104,N_7978,N_7992);
nand U8105 (N_8105,N_7846,N_7882);
xor U8106 (N_8106,N_7927,N_7841);
xnor U8107 (N_8107,N_7976,N_7914);
xnor U8108 (N_8108,N_7866,N_7913);
nor U8109 (N_8109,N_7846,N_7995);
and U8110 (N_8110,N_7857,N_7879);
and U8111 (N_8111,N_7844,N_7870);
and U8112 (N_8112,N_7856,N_7983);
xnor U8113 (N_8113,N_7938,N_7994);
xor U8114 (N_8114,N_7923,N_7945);
nand U8115 (N_8115,N_7982,N_7901);
nand U8116 (N_8116,N_7953,N_7892);
or U8117 (N_8117,N_7897,N_7980);
or U8118 (N_8118,N_7921,N_7895);
xor U8119 (N_8119,N_7862,N_7948);
nand U8120 (N_8120,N_7940,N_7908);
xnor U8121 (N_8121,N_7947,N_7940);
or U8122 (N_8122,N_7938,N_7940);
or U8123 (N_8123,N_7983,N_7852);
or U8124 (N_8124,N_7931,N_7905);
nor U8125 (N_8125,N_7939,N_7981);
and U8126 (N_8126,N_7945,N_7983);
nand U8127 (N_8127,N_7901,N_7920);
or U8128 (N_8128,N_7905,N_7904);
or U8129 (N_8129,N_7913,N_7863);
and U8130 (N_8130,N_7999,N_7985);
nor U8131 (N_8131,N_7919,N_7950);
or U8132 (N_8132,N_7891,N_7920);
xnor U8133 (N_8133,N_7885,N_7882);
or U8134 (N_8134,N_7887,N_7982);
nor U8135 (N_8135,N_7868,N_7891);
or U8136 (N_8136,N_7844,N_7881);
or U8137 (N_8137,N_7876,N_7990);
nor U8138 (N_8138,N_7943,N_7981);
or U8139 (N_8139,N_7875,N_7903);
nor U8140 (N_8140,N_7994,N_7881);
nor U8141 (N_8141,N_7857,N_7892);
nor U8142 (N_8142,N_7939,N_7922);
nand U8143 (N_8143,N_7985,N_7852);
xnor U8144 (N_8144,N_7849,N_7916);
xor U8145 (N_8145,N_7893,N_7883);
nor U8146 (N_8146,N_7982,N_7965);
and U8147 (N_8147,N_7878,N_7874);
nor U8148 (N_8148,N_7894,N_7948);
nor U8149 (N_8149,N_7948,N_7891);
and U8150 (N_8150,N_7840,N_7990);
and U8151 (N_8151,N_7960,N_7988);
nand U8152 (N_8152,N_7920,N_7847);
nand U8153 (N_8153,N_7875,N_7847);
nor U8154 (N_8154,N_7940,N_7914);
nand U8155 (N_8155,N_7926,N_7970);
and U8156 (N_8156,N_7946,N_7980);
and U8157 (N_8157,N_7924,N_7853);
nor U8158 (N_8158,N_7989,N_7853);
nand U8159 (N_8159,N_7882,N_7927);
nor U8160 (N_8160,N_8159,N_8155);
and U8161 (N_8161,N_8142,N_8073);
xor U8162 (N_8162,N_8001,N_8042);
nand U8163 (N_8163,N_8030,N_8057);
and U8164 (N_8164,N_8126,N_8134);
or U8165 (N_8165,N_8033,N_8091);
nand U8166 (N_8166,N_8068,N_8148);
nor U8167 (N_8167,N_8083,N_8045);
or U8168 (N_8168,N_8016,N_8021);
nor U8169 (N_8169,N_8075,N_8052);
nor U8170 (N_8170,N_8081,N_8055);
nand U8171 (N_8171,N_8003,N_8028);
and U8172 (N_8172,N_8061,N_8103);
and U8173 (N_8173,N_8124,N_8090);
nor U8174 (N_8174,N_8004,N_8144);
nor U8175 (N_8175,N_8022,N_8077);
xnor U8176 (N_8176,N_8146,N_8060);
and U8177 (N_8177,N_8015,N_8065);
and U8178 (N_8178,N_8141,N_8130);
nor U8179 (N_8179,N_8106,N_8132);
and U8180 (N_8180,N_8070,N_8105);
and U8181 (N_8181,N_8100,N_8131);
or U8182 (N_8182,N_8121,N_8064);
nand U8183 (N_8183,N_8069,N_8128);
nor U8184 (N_8184,N_8035,N_8102);
nor U8185 (N_8185,N_8108,N_8002);
xnor U8186 (N_8186,N_8074,N_8029);
nor U8187 (N_8187,N_8044,N_8113);
nand U8188 (N_8188,N_8118,N_8063);
xnor U8189 (N_8189,N_8154,N_8094);
nand U8190 (N_8190,N_8085,N_8007);
nor U8191 (N_8191,N_8151,N_8125);
and U8192 (N_8192,N_8025,N_8017);
nor U8193 (N_8193,N_8082,N_8153);
nor U8194 (N_8194,N_8088,N_8080);
nand U8195 (N_8195,N_8006,N_8135);
nor U8196 (N_8196,N_8157,N_8032);
and U8197 (N_8197,N_8127,N_8104);
and U8198 (N_8198,N_8110,N_8048);
nand U8199 (N_8199,N_8031,N_8005);
nand U8200 (N_8200,N_8027,N_8036);
nor U8201 (N_8201,N_8079,N_8111);
and U8202 (N_8202,N_8037,N_8140);
and U8203 (N_8203,N_8117,N_8020);
and U8204 (N_8204,N_8152,N_8051);
and U8205 (N_8205,N_8112,N_8043);
xnor U8206 (N_8206,N_8013,N_8034);
xor U8207 (N_8207,N_8000,N_8122);
nor U8208 (N_8208,N_8024,N_8138);
and U8209 (N_8209,N_8040,N_8053);
or U8210 (N_8210,N_8115,N_8119);
or U8211 (N_8211,N_8041,N_8129);
xnor U8212 (N_8212,N_8095,N_8067);
nand U8213 (N_8213,N_8156,N_8008);
xnor U8214 (N_8214,N_8066,N_8023);
nand U8215 (N_8215,N_8076,N_8133);
xnor U8216 (N_8216,N_8058,N_8026);
nand U8217 (N_8217,N_8123,N_8039);
nor U8218 (N_8218,N_8158,N_8084);
and U8219 (N_8219,N_8145,N_8096);
nor U8220 (N_8220,N_8147,N_8009);
or U8221 (N_8221,N_8093,N_8014);
xor U8222 (N_8222,N_8056,N_8010);
and U8223 (N_8223,N_8011,N_8078);
or U8224 (N_8224,N_8054,N_8116);
or U8225 (N_8225,N_8062,N_8149);
or U8226 (N_8226,N_8089,N_8114);
and U8227 (N_8227,N_8047,N_8143);
or U8228 (N_8228,N_8046,N_8120);
nor U8229 (N_8229,N_8019,N_8101);
xnor U8230 (N_8230,N_8099,N_8050);
and U8231 (N_8231,N_8087,N_8071);
and U8232 (N_8232,N_8038,N_8107);
xnor U8233 (N_8233,N_8098,N_8072);
nand U8234 (N_8234,N_8139,N_8086);
or U8235 (N_8235,N_8136,N_8137);
or U8236 (N_8236,N_8150,N_8109);
and U8237 (N_8237,N_8049,N_8092);
nand U8238 (N_8238,N_8059,N_8097);
nand U8239 (N_8239,N_8012,N_8018);
and U8240 (N_8240,N_8089,N_8060);
or U8241 (N_8241,N_8002,N_8158);
xnor U8242 (N_8242,N_8115,N_8151);
xor U8243 (N_8243,N_8048,N_8021);
or U8244 (N_8244,N_8141,N_8074);
xnor U8245 (N_8245,N_8144,N_8032);
xnor U8246 (N_8246,N_8127,N_8031);
nand U8247 (N_8247,N_8090,N_8057);
and U8248 (N_8248,N_8151,N_8077);
nor U8249 (N_8249,N_8000,N_8107);
nand U8250 (N_8250,N_8108,N_8049);
xor U8251 (N_8251,N_8103,N_8073);
xnor U8252 (N_8252,N_8107,N_8008);
or U8253 (N_8253,N_8158,N_8096);
nor U8254 (N_8254,N_8155,N_8006);
nor U8255 (N_8255,N_8099,N_8083);
xnor U8256 (N_8256,N_8112,N_8073);
and U8257 (N_8257,N_8009,N_8077);
nand U8258 (N_8258,N_8052,N_8030);
and U8259 (N_8259,N_8124,N_8019);
or U8260 (N_8260,N_8113,N_8132);
nor U8261 (N_8261,N_8150,N_8086);
nor U8262 (N_8262,N_8097,N_8076);
or U8263 (N_8263,N_8063,N_8070);
xnor U8264 (N_8264,N_8117,N_8069);
nor U8265 (N_8265,N_8076,N_8042);
nand U8266 (N_8266,N_8121,N_8050);
nor U8267 (N_8267,N_8070,N_8143);
xor U8268 (N_8268,N_8126,N_8004);
and U8269 (N_8269,N_8098,N_8058);
and U8270 (N_8270,N_8114,N_8049);
xnor U8271 (N_8271,N_8017,N_8073);
nor U8272 (N_8272,N_8095,N_8091);
xor U8273 (N_8273,N_8034,N_8030);
and U8274 (N_8274,N_8035,N_8150);
nor U8275 (N_8275,N_8152,N_8070);
nand U8276 (N_8276,N_8094,N_8078);
or U8277 (N_8277,N_8077,N_8143);
xnor U8278 (N_8278,N_8084,N_8098);
and U8279 (N_8279,N_8129,N_8073);
xor U8280 (N_8280,N_8005,N_8130);
xor U8281 (N_8281,N_8095,N_8002);
or U8282 (N_8282,N_8105,N_8093);
or U8283 (N_8283,N_8071,N_8028);
xnor U8284 (N_8284,N_8080,N_8131);
xnor U8285 (N_8285,N_8030,N_8056);
nor U8286 (N_8286,N_8000,N_8011);
nor U8287 (N_8287,N_8032,N_8059);
or U8288 (N_8288,N_8034,N_8027);
nor U8289 (N_8289,N_8070,N_8038);
xnor U8290 (N_8290,N_8031,N_8146);
or U8291 (N_8291,N_8060,N_8156);
and U8292 (N_8292,N_8064,N_8098);
and U8293 (N_8293,N_8137,N_8119);
or U8294 (N_8294,N_8023,N_8018);
nor U8295 (N_8295,N_8030,N_8107);
and U8296 (N_8296,N_8150,N_8139);
xnor U8297 (N_8297,N_8086,N_8061);
or U8298 (N_8298,N_8122,N_8022);
nor U8299 (N_8299,N_8059,N_8093);
nor U8300 (N_8300,N_8008,N_8002);
nor U8301 (N_8301,N_8067,N_8147);
xor U8302 (N_8302,N_8015,N_8132);
xor U8303 (N_8303,N_8019,N_8153);
xnor U8304 (N_8304,N_8019,N_8063);
nand U8305 (N_8305,N_8056,N_8018);
and U8306 (N_8306,N_8125,N_8147);
xnor U8307 (N_8307,N_8107,N_8058);
nand U8308 (N_8308,N_8118,N_8100);
nor U8309 (N_8309,N_8051,N_8083);
nand U8310 (N_8310,N_8007,N_8104);
xor U8311 (N_8311,N_8055,N_8105);
and U8312 (N_8312,N_8101,N_8138);
and U8313 (N_8313,N_8015,N_8045);
xnor U8314 (N_8314,N_8158,N_8115);
or U8315 (N_8315,N_8056,N_8142);
nand U8316 (N_8316,N_8085,N_8141);
nand U8317 (N_8317,N_8138,N_8058);
nand U8318 (N_8318,N_8125,N_8116);
and U8319 (N_8319,N_8088,N_8016);
or U8320 (N_8320,N_8249,N_8280);
nor U8321 (N_8321,N_8300,N_8243);
xor U8322 (N_8322,N_8203,N_8213);
or U8323 (N_8323,N_8186,N_8306);
nor U8324 (N_8324,N_8301,N_8171);
xor U8325 (N_8325,N_8211,N_8319);
xnor U8326 (N_8326,N_8170,N_8183);
and U8327 (N_8327,N_8262,N_8252);
nand U8328 (N_8328,N_8205,N_8289);
nor U8329 (N_8329,N_8304,N_8308);
and U8330 (N_8330,N_8225,N_8310);
or U8331 (N_8331,N_8281,N_8266);
and U8332 (N_8332,N_8233,N_8163);
xnor U8333 (N_8333,N_8272,N_8264);
nand U8334 (N_8334,N_8317,N_8167);
and U8335 (N_8335,N_8294,N_8284);
nand U8336 (N_8336,N_8241,N_8296);
xnor U8337 (N_8337,N_8188,N_8277);
nor U8338 (N_8338,N_8192,N_8212);
and U8339 (N_8339,N_8221,N_8292);
and U8340 (N_8340,N_8283,N_8290);
nand U8341 (N_8341,N_8191,N_8298);
and U8342 (N_8342,N_8295,N_8314);
or U8343 (N_8343,N_8215,N_8311);
nand U8344 (N_8344,N_8232,N_8162);
and U8345 (N_8345,N_8302,N_8216);
and U8346 (N_8346,N_8226,N_8263);
or U8347 (N_8347,N_8208,N_8313);
and U8348 (N_8348,N_8161,N_8316);
or U8349 (N_8349,N_8229,N_8201);
and U8350 (N_8350,N_8223,N_8199);
and U8351 (N_8351,N_8297,N_8180);
and U8352 (N_8352,N_8242,N_8190);
and U8353 (N_8353,N_8187,N_8270);
or U8354 (N_8354,N_8210,N_8178);
and U8355 (N_8355,N_8165,N_8278);
nand U8356 (N_8356,N_8244,N_8204);
xnor U8357 (N_8357,N_8315,N_8287);
xnor U8358 (N_8358,N_8237,N_8197);
or U8359 (N_8359,N_8307,N_8275);
or U8360 (N_8360,N_8220,N_8247);
or U8361 (N_8361,N_8254,N_8267);
and U8362 (N_8362,N_8184,N_8164);
nor U8363 (N_8363,N_8166,N_8279);
or U8364 (N_8364,N_8257,N_8193);
nor U8365 (N_8365,N_8258,N_8318);
nand U8366 (N_8366,N_8282,N_8269);
or U8367 (N_8367,N_8248,N_8206);
nor U8368 (N_8368,N_8238,N_8288);
or U8369 (N_8369,N_8219,N_8268);
nand U8370 (N_8370,N_8202,N_8218);
nor U8371 (N_8371,N_8274,N_8239);
and U8372 (N_8372,N_8169,N_8265);
or U8373 (N_8373,N_8261,N_8312);
nand U8374 (N_8374,N_8224,N_8256);
nand U8375 (N_8375,N_8293,N_8240);
nand U8376 (N_8376,N_8236,N_8179);
xor U8377 (N_8377,N_8160,N_8271);
xnor U8378 (N_8378,N_8255,N_8217);
nand U8379 (N_8379,N_8273,N_8299);
or U8380 (N_8380,N_8194,N_8228);
nand U8381 (N_8381,N_8230,N_8207);
or U8382 (N_8382,N_8181,N_8276);
nor U8383 (N_8383,N_8231,N_8222);
nor U8384 (N_8384,N_8291,N_8198);
nand U8385 (N_8385,N_8173,N_8259);
nand U8386 (N_8386,N_8235,N_8214);
nor U8387 (N_8387,N_8246,N_8227);
and U8388 (N_8388,N_8260,N_8245);
nand U8389 (N_8389,N_8234,N_8200);
nand U8390 (N_8390,N_8209,N_8305);
nand U8391 (N_8391,N_8195,N_8303);
nand U8392 (N_8392,N_8174,N_8172);
nand U8393 (N_8393,N_8196,N_8251);
or U8394 (N_8394,N_8168,N_8182);
or U8395 (N_8395,N_8175,N_8185);
nor U8396 (N_8396,N_8176,N_8250);
nor U8397 (N_8397,N_8285,N_8253);
and U8398 (N_8398,N_8177,N_8189);
nand U8399 (N_8399,N_8309,N_8286);
or U8400 (N_8400,N_8205,N_8197);
or U8401 (N_8401,N_8301,N_8250);
and U8402 (N_8402,N_8262,N_8161);
or U8403 (N_8403,N_8181,N_8310);
xnor U8404 (N_8404,N_8199,N_8192);
and U8405 (N_8405,N_8235,N_8299);
nor U8406 (N_8406,N_8258,N_8170);
xor U8407 (N_8407,N_8263,N_8292);
and U8408 (N_8408,N_8293,N_8161);
xnor U8409 (N_8409,N_8283,N_8284);
or U8410 (N_8410,N_8209,N_8197);
nor U8411 (N_8411,N_8271,N_8222);
and U8412 (N_8412,N_8228,N_8258);
nor U8413 (N_8413,N_8172,N_8304);
nand U8414 (N_8414,N_8249,N_8205);
xnor U8415 (N_8415,N_8166,N_8163);
nor U8416 (N_8416,N_8274,N_8308);
xor U8417 (N_8417,N_8287,N_8198);
nor U8418 (N_8418,N_8177,N_8289);
nor U8419 (N_8419,N_8195,N_8251);
xor U8420 (N_8420,N_8236,N_8282);
or U8421 (N_8421,N_8286,N_8211);
nand U8422 (N_8422,N_8233,N_8300);
and U8423 (N_8423,N_8282,N_8212);
nand U8424 (N_8424,N_8265,N_8160);
or U8425 (N_8425,N_8170,N_8285);
or U8426 (N_8426,N_8238,N_8279);
nand U8427 (N_8427,N_8287,N_8241);
nand U8428 (N_8428,N_8167,N_8299);
or U8429 (N_8429,N_8292,N_8171);
xnor U8430 (N_8430,N_8308,N_8215);
nor U8431 (N_8431,N_8197,N_8183);
and U8432 (N_8432,N_8302,N_8212);
or U8433 (N_8433,N_8238,N_8318);
xnor U8434 (N_8434,N_8278,N_8292);
xnor U8435 (N_8435,N_8273,N_8185);
xnor U8436 (N_8436,N_8219,N_8261);
xor U8437 (N_8437,N_8219,N_8246);
nand U8438 (N_8438,N_8299,N_8227);
or U8439 (N_8439,N_8198,N_8269);
nand U8440 (N_8440,N_8169,N_8196);
nor U8441 (N_8441,N_8229,N_8276);
nor U8442 (N_8442,N_8244,N_8199);
nor U8443 (N_8443,N_8260,N_8276);
and U8444 (N_8444,N_8187,N_8181);
and U8445 (N_8445,N_8246,N_8280);
and U8446 (N_8446,N_8307,N_8258);
or U8447 (N_8447,N_8246,N_8266);
xnor U8448 (N_8448,N_8231,N_8256);
xnor U8449 (N_8449,N_8304,N_8272);
xnor U8450 (N_8450,N_8170,N_8202);
and U8451 (N_8451,N_8267,N_8217);
xnor U8452 (N_8452,N_8317,N_8283);
and U8453 (N_8453,N_8316,N_8319);
nor U8454 (N_8454,N_8272,N_8166);
nand U8455 (N_8455,N_8252,N_8175);
and U8456 (N_8456,N_8221,N_8297);
or U8457 (N_8457,N_8234,N_8163);
and U8458 (N_8458,N_8162,N_8265);
xor U8459 (N_8459,N_8267,N_8265);
xor U8460 (N_8460,N_8304,N_8277);
or U8461 (N_8461,N_8267,N_8226);
nor U8462 (N_8462,N_8319,N_8296);
nor U8463 (N_8463,N_8279,N_8219);
nor U8464 (N_8464,N_8314,N_8265);
and U8465 (N_8465,N_8311,N_8181);
nor U8466 (N_8466,N_8293,N_8209);
xnor U8467 (N_8467,N_8230,N_8168);
nand U8468 (N_8468,N_8236,N_8233);
nand U8469 (N_8469,N_8245,N_8287);
or U8470 (N_8470,N_8163,N_8214);
nor U8471 (N_8471,N_8258,N_8234);
or U8472 (N_8472,N_8221,N_8271);
xnor U8473 (N_8473,N_8218,N_8279);
xor U8474 (N_8474,N_8282,N_8246);
or U8475 (N_8475,N_8167,N_8267);
and U8476 (N_8476,N_8267,N_8263);
nor U8477 (N_8477,N_8179,N_8173);
and U8478 (N_8478,N_8274,N_8279);
and U8479 (N_8479,N_8160,N_8168);
and U8480 (N_8480,N_8394,N_8400);
nor U8481 (N_8481,N_8425,N_8439);
and U8482 (N_8482,N_8387,N_8350);
xnor U8483 (N_8483,N_8346,N_8376);
or U8484 (N_8484,N_8321,N_8384);
nand U8485 (N_8485,N_8379,N_8443);
nor U8486 (N_8486,N_8385,N_8388);
and U8487 (N_8487,N_8419,N_8408);
nor U8488 (N_8488,N_8479,N_8327);
xnor U8489 (N_8489,N_8468,N_8364);
nand U8490 (N_8490,N_8344,N_8389);
or U8491 (N_8491,N_8465,N_8462);
and U8492 (N_8492,N_8454,N_8447);
or U8493 (N_8493,N_8471,N_8457);
and U8494 (N_8494,N_8459,N_8435);
and U8495 (N_8495,N_8338,N_8352);
nand U8496 (N_8496,N_8402,N_8444);
nand U8497 (N_8497,N_8428,N_8417);
nand U8498 (N_8498,N_8329,N_8372);
or U8499 (N_8499,N_8446,N_8368);
and U8500 (N_8500,N_8455,N_8354);
nor U8501 (N_8501,N_8328,N_8467);
and U8502 (N_8502,N_8440,N_8353);
and U8503 (N_8503,N_8431,N_8423);
and U8504 (N_8504,N_8334,N_8342);
and U8505 (N_8505,N_8436,N_8332);
and U8506 (N_8506,N_8351,N_8476);
and U8507 (N_8507,N_8361,N_8386);
nor U8508 (N_8508,N_8367,N_8362);
xnor U8509 (N_8509,N_8463,N_8399);
xor U8510 (N_8510,N_8424,N_8373);
nor U8511 (N_8511,N_8477,N_8437);
nand U8512 (N_8512,N_8324,N_8356);
and U8513 (N_8513,N_8348,N_8438);
nor U8514 (N_8514,N_8358,N_8366);
and U8515 (N_8515,N_8369,N_8375);
xnor U8516 (N_8516,N_8448,N_8320);
nor U8517 (N_8517,N_8331,N_8359);
or U8518 (N_8518,N_8405,N_8434);
xor U8519 (N_8519,N_8360,N_8411);
xor U8520 (N_8520,N_8326,N_8426);
nor U8521 (N_8521,N_8456,N_8371);
nand U8522 (N_8522,N_8422,N_8430);
xnor U8523 (N_8523,N_8470,N_8343);
nand U8524 (N_8524,N_8377,N_8441);
and U8525 (N_8525,N_8410,N_8378);
and U8526 (N_8526,N_8381,N_8432);
xor U8527 (N_8527,N_8337,N_8412);
nor U8528 (N_8528,N_8429,N_8451);
xnor U8529 (N_8529,N_8392,N_8458);
or U8530 (N_8530,N_8433,N_8404);
and U8531 (N_8531,N_8453,N_8395);
and U8532 (N_8532,N_8415,N_8445);
and U8533 (N_8533,N_8357,N_8478);
or U8534 (N_8534,N_8427,N_8396);
nor U8535 (N_8535,N_8420,N_8421);
xnor U8536 (N_8536,N_8341,N_8473);
nand U8537 (N_8537,N_8401,N_8374);
nand U8538 (N_8538,N_8413,N_8336);
and U8539 (N_8539,N_8347,N_8335);
xor U8540 (N_8540,N_8355,N_8442);
nand U8541 (N_8541,N_8475,N_8325);
and U8542 (N_8542,N_8363,N_8330);
and U8543 (N_8543,N_8365,N_8414);
nand U8544 (N_8544,N_8323,N_8382);
or U8545 (N_8545,N_8345,N_8460);
nand U8546 (N_8546,N_8406,N_8391);
or U8547 (N_8547,N_8403,N_8416);
and U8548 (N_8548,N_8452,N_8464);
nand U8549 (N_8549,N_8461,N_8333);
and U8550 (N_8550,N_8469,N_8398);
and U8551 (N_8551,N_8340,N_8450);
nand U8552 (N_8552,N_8466,N_8390);
and U8553 (N_8553,N_8472,N_8397);
nand U8554 (N_8554,N_8418,N_8383);
or U8555 (N_8555,N_8393,N_8349);
xor U8556 (N_8556,N_8370,N_8449);
or U8557 (N_8557,N_8407,N_8339);
or U8558 (N_8558,N_8380,N_8409);
or U8559 (N_8559,N_8322,N_8474);
nor U8560 (N_8560,N_8406,N_8390);
nor U8561 (N_8561,N_8321,N_8471);
nand U8562 (N_8562,N_8377,N_8416);
and U8563 (N_8563,N_8467,N_8320);
or U8564 (N_8564,N_8415,N_8348);
xnor U8565 (N_8565,N_8428,N_8462);
xnor U8566 (N_8566,N_8356,N_8355);
and U8567 (N_8567,N_8335,N_8474);
or U8568 (N_8568,N_8453,N_8371);
and U8569 (N_8569,N_8421,N_8372);
nand U8570 (N_8570,N_8424,N_8387);
xor U8571 (N_8571,N_8387,N_8383);
and U8572 (N_8572,N_8443,N_8469);
nand U8573 (N_8573,N_8421,N_8395);
nor U8574 (N_8574,N_8459,N_8331);
nand U8575 (N_8575,N_8461,N_8420);
nor U8576 (N_8576,N_8380,N_8395);
and U8577 (N_8577,N_8403,N_8339);
or U8578 (N_8578,N_8471,N_8371);
or U8579 (N_8579,N_8424,N_8426);
or U8580 (N_8580,N_8415,N_8357);
xnor U8581 (N_8581,N_8373,N_8358);
nor U8582 (N_8582,N_8449,N_8407);
or U8583 (N_8583,N_8389,N_8477);
and U8584 (N_8584,N_8471,N_8377);
nor U8585 (N_8585,N_8336,N_8427);
xnor U8586 (N_8586,N_8433,N_8432);
or U8587 (N_8587,N_8439,N_8456);
xnor U8588 (N_8588,N_8341,N_8452);
nand U8589 (N_8589,N_8450,N_8421);
xor U8590 (N_8590,N_8383,N_8347);
and U8591 (N_8591,N_8339,N_8357);
xnor U8592 (N_8592,N_8380,N_8433);
xnor U8593 (N_8593,N_8415,N_8429);
or U8594 (N_8594,N_8368,N_8377);
xnor U8595 (N_8595,N_8381,N_8410);
nor U8596 (N_8596,N_8331,N_8411);
xnor U8597 (N_8597,N_8470,N_8466);
nor U8598 (N_8598,N_8320,N_8392);
or U8599 (N_8599,N_8461,N_8459);
nor U8600 (N_8600,N_8396,N_8463);
nand U8601 (N_8601,N_8473,N_8453);
and U8602 (N_8602,N_8449,N_8458);
nor U8603 (N_8603,N_8442,N_8426);
nor U8604 (N_8604,N_8402,N_8424);
nor U8605 (N_8605,N_8344,N_8420);
and U8606 (N_8606,N_8324,N_8405);
xor U8607 (N_8607,N_8419,N_8328);
xor U8608 (N_8608,N_8348,N_8367);
or U8609 (N_8609,N_8436,N_8456);
xor U8610 (N_8610,N_8325,N_8470);
nand U8611 (N_8611,N_8392,N_8466);
or U8612 (N_8612,N_8478,N_8383);
or U8613 (N_8613,N_8409,N_8476);
xnor U8614 (N_8614,N_8433,N_8394);
xor U8615 (N_8615,N_8330,N_8443);
xnor U8616 (N_8616,N_8417,N_8355);
or U8617 (N_8617,N_8429,N_8355);
or U8618 (N_8618,N_8393,N_8445);
or U8619 (N_8619,N_8402,N_8327);
nand U8620 (N_8620,N_8359,N_8358);
nor U8621 (N_8621,N_8379,N_8411);
nand U8622 (N_8622,N_8456,N_8471);
xnor U8623 (N_8623,N_8391,N_8460);
nor U8624 (N_8624,N_8417,N_8410);
or U8625 (N_8625,N_8444,N_8416);
and U8626 (N_8626,N_8409,N_8474);
xor U8627 (N_8627,N_8412,N_8396);
xor U8628 (N_8628,N_8346,N_8389);
nand U8629 (N_8629,N_8414,N_8442);
and U8630 (N_8630,N_8383,N_8379);
or U8631 (N_8631,N_8434,N_8359);
nor U8632 (N_8632,N_8411,N_8441);
nand U8633 (N_8633,N_8372,N_8436);
xor U8634 (N_8634,N_8451,N_8397);
and U8635 (N_8635,N_8358,N_8458);
nor U8636 (N_8636,N_8473,N_8329);
or U8637 (N_8637,N_8352,N_8365);
xnor U8638 (N_8638,N_8449,N_8403);
nand U8639 (N_8639,N_8424,N_8386);
nand U8640 (N_8640,N_8490,N_8524);
nand U8641 (N_8641,N_8493,N_8558);
or U8642 (N_8642,N_8545,N_8523);
and U8643 (N_8643,N_8481,N_8583);
xor U8644 (N_8644,N_8561,N_8483);
nor U8645 (N_8645,N_8639,N_8637);
nor U8646 (N_8646,N_8613,N_8500);
xnor U8647 (N_8647,N_8597,N_8636);
nand U8648 (N_8648,N_8496,N_8528);
and U8649 (N_8649,N_8628,N_8592);
and U8650 (N_8650,N_8608,N_8516);
or U8651 (N_8651,N_8556,N_8601);
or U8652 (N_8652,N_8522,N_8638);
nor U8653 (N_8653,N_8527,N_8499);
xnor U8654 (N_8654,N_8492,N_8559);
nand U8655 (N_8655,N_8508,N_8562);
or U8656 (N_8656,N_8624,N_8615);
and U8657 (N_8657,N_8485,N_8541);
or U8658 (N_8658,N_8495,N_8482);
or U8659 (N_8659,N_8521,N_8599);
and U8660 (N_8660,N_8629,N_8633);
or U8661 (N_8661,N_8498,N_8544);
xor U8662 (N_8662,N_8486,N_8570);
and U8663 (N_8663,N_8563,N_8487);
xor U8664 (N_8664,N_8512,N_8536);
nor U8665 (N_8665,N_8614,N_8553);
or U8666 (N_8666,N_8564,N_8548);
nand U8667 (N_8667,N_8491,N_8611);
and U8668 (N_8668,N_8589,N_8598);
and U8669 (N_8669,N_8502,N_8554);
nand U8670 (N_8670,N_8625,N_8538);
or U8671 (N_8671,N_8576,N_8568);
or U8672 (N_8672,N_8619,N_8566);
or U8673 (N_8673,N_8616,N_8543);
and U8674 (N_8674,N_8579,N_8525);
nor U8675 (N_8675,N_8519,N_8551);
xor U8676 (N_8676,N_8622,N_8480);
nand U8677 (N_8677,N_8489,N_8635);
nand U8678 (N_8678,N_8582,N_8552);
or U8679 (N_8679,N_8631,N_8586);
or U8680 (N_8680,N_8600,N_8526);
xor U8681 (N_8681,N_8603,N_8511);
and U8682 (N_8682,N_8606,N_8501);
or U8683 (N_8683,N_8510,N_8595);
or U8684 (N_8684,N_8604,N_8497);
nand U8685 (N_8685,N_8540,N_8605);
nor U8686 (N_8686,N_8509,N_8575);
nor U8687 (N_8687,N_8537,N_8535);
or U8688 (N_8688,N_8587,N_8594);
nor U8689 (N_8689,N_8618,N_8577);
xnor U8690 (N_8690,N_8602,N_8571);
nand U8691 (N_8691,N_8488,N_8621);
and U8692 (N_8692,N_8533,N_8534);
and U8693 (N_8693,N_8531,N_8529);
nand U8694 (N_8694,N_8627,N_8507);
nand U8695 (N_8695,N_8574,N_8550);
nand U8696 (N_8696,N_8549,N_8610);
and U8697 (N_8697,N_8634,N_8612);
nand U8698 (N_8698,N_8494,N_8626);
or U8699 (N_8699,N_8565,N_8530);
nor U8700 (N_8700,N_8557,N_8584);
and U8701 (N_8701,N_8484,N_8532);
nor U8702 (N_8702,N_8542,N_8555);
xnor U8703 (N_8703,N_8588,N_8567);
xnor U8704 (N_8704,N_8572,N_8560);
nand U8705 (N_8705,N_8569,N_8505);
nor U8706 (N_8706,N_8609,N_8539);
xor U8707 (N_8707,N_8506,N_8620);
nand U8708 (N_8708,N_8518,N_8617);
and U8709 (N_8709,N_8630,N_8578);
and U8710 (N_8710,N_8632,N_8514);
xor U8711 (N_8711,N_8596,N_8580);
or U8712 (N_8712,N_8573,N_8623);
nand U8713 (N_8713,N_8590,N_8591);
nor U8714 (N_8714,N_8547,N_8503);
or U8715 (N_8715,N_8504,N_8593);
and U8716 (N_8716,N_8607,N_8517);
or U8717 (N_8717,N_8581,N_8520);
and U8718 (N_8718,N_8546,N_8515);
nand U8719 (N_8719,N_8513,N_8585);
nor U8720 (N_8720,N_8494,N_8632);
nor U8721 (N_8721,N_8526,N_8521);
or U8722 (N_8722,N_8614,N_8604);
xor U8723 (N_8723,N_8542,N_8617);
xnor U8724 (N_8724,N_8563,N_8603);
and U8725 (N_8725,N_8558,N_8526);
xor U8726 (N_8726,N_8493,N_8561);
and U8727 (N_8727,N_8628,N_8521);
nor U8728 (N_8728,N_8565,N_8639);
nand U8729 (N_8729,N_8595,N_8509);
or U8730 (N_8730,N_8515,N_8582);
nand U8731 (N_8731,N_8521,N_8601);
and U8732 (N_8732,N_8618,N_8599);
nor U8733 (N_8733,N_8613,N_8502);
and U8734 (N_8734,N_8595,N_8620);
or U8735 (N_8735,N_8563,N_8541);
and U8736 (N_8736,N_8559,N_8574);
nand U8737 (N_8737,N_8505,N_8581);
and U8738 (N_8738,N_8491,N_8542);
xor U8739 (N_8739,N_8490,N_8599);
nor U8740 (N_8740,N_8612,N_8557);
xnor U8741 (N_8741,N_8540,N_8579);
nor U8742 (N_8742,N_8532,N_8564);
xnor U8743 (N_8743,N_8613,N_8633);
or U8744 (N_8744,N_8510,N_8636);
xor U8745 (N_8745,N_8497,N_8616);
or U8746 (N_8746,N_8489,N_8537);
and U8747 (N_8747,N_8505,N_8551);
and U8748 (N_8748,N_8575,N_8622);
nor U8749 (N_8749,N_8544,N_8540);
and U8750 (N_8750,N_8614,N_8505);
and U8751 (N_8751,N_8511,N_8536);
nand U8752 (N_8752,N_8528,N_8555);
nand U8753 (N_8753,N_8514,N_8630);
nand U8754 (N_8754,N_8490,N_8580);
nor U8755 (N_8755,N_8638,N_8622);
and U8756 (N_8756,N_8534,N_8545);
and U8757 (N_8757,N_8498,N_8493);
xnor U8758 (N_8758,N_8547,N_8568);
xor U8759 (N_8759,N_8621,N_8611);
xnor U8760 (N_8760,N_8482,N_8484);
nand U8761 (N_8761,N_8521,N_8520);
nand U8762 (N_8762,N_8489,N_8534);
and U8763 (N_8763,N_8579,N_8527);
or U8764 (N_8764,N_8534,N_8630);
and U8765 (N_8765,N_8568,N_8637);
xor U8766 (N_8766,N_8531,N_8559);
nand U8767 (N_8767,N_8497,N_8617);
or U8768 (N_8768,N_8549,N_8560);
or U8769 (N_8769,N_8613,N_8554);
nand U8770 (N_8770,N_8578,N_8510);
nor U8771 (N_8771,N_8568,N_8626);
or U8772 (N_8772,N_8534,N_8562);
nor U8773 (N_8773,N_8492,N_8575);
nor U8774 (N_8774,N_8529,N_8525);
or U8775 (N_8775,N_8580,N_8633);
xnor U8776 (N_8776,N_8505,N_8539);
nand U8777 (N_8777,N_8500,N_8612);
nor U8778 (N_8778,N_8499,N_8513);
and U8779 (N_8779,N_8586,N_8497);
nor U8780 (N_8780,N_8578,N_8581);
xnor U8781 (N_8781,N_8536,N_8555);
xnor U8782 (N_8782,N_8636,N_8634);
and U8783 (N_8783,N_8511,N_8548);
and U8784 (N_8784,N_8543,N_8577);
xor U8785 (N_8785,N_8604,N_8483);
nor U8786 (N_8786,N_8520,N_8544);
nor U8787 (N_8787,N_8532,N_8552);
nand U8788 (N_8788,N_8543,N_8613);
nand U8789 (N_8789,N_8575,N_8533);
or U8790 (N_8790,N_8585,N_8613);
xor U8791 (N_8791,N_8572,N_8566);
or U8792 (N_8792,N_8607,N_8488);
or U8793 (N_8793,N_8548,N_8600);
nand U8794 (N_8794,N_8599,N_8586);
nand U8795 (N_8795,N_8601,N_8505);
and U8796 (N_8796,N_8539,N_8503);
xor U8797 (N_8797,N_8585,N_8637);
and U8798 (N_8798,N_8620,N_8621);
or U8799 (N_8799,N_8633,N_8575);
nand U8800 (N_8800,N_8666,N_8690);
and U8801 (N_8801,N_8799,N_8794);
nand U8802 (N_8802,N_8750,N_8655);
nor U8803 (N_8803,N_8729,N_8650);
nor U8804 (N_8804,N_8778,N_8702);
nand U8805 (N_8805,N_8685,N_8663);
or U8806 (N_8806,N_8755,N_8733);
and U8807 (N_8807,N_8765,N_8659);
nand U8808 (N_8808,N_8726,N_8725);
or U8809 (N_8809,N_8641,N_8746);
nand U8810 (N_8810,N_8691,N_8642);
xor U8811 (N_8811,N_8752,N_8644);
or U8812 (N_8812,N_8703,N_8751);
xor U8813 (N_8813,N_8737,N_8734);
nor U8814 (N_8814,N_8764,N_8773);
or U8815 (N_8815,N_8745,N_8679);
xor U8816 (N_8816,N_8645,N_8687);
or U8817 (N_8817,N_8721,N_8742);
nor U8818 (N_8818,N_8724,N_8732);
and U8819 (N_8819,N_8762,N_8664);
or U8820 (N_8820,N_8793,N_8789);
xor U8821 (N_8821,N_8672,N_8766);
xor U8822 (N_8822,N_8795,N_8707);
nand U8823 (N_8823,N_8722,N_8782);
nand U8824 (N_8824,N_8647,N_8718);
xnor U8825 (N_8825,N_8786,N_8728);
nand U8826 (N_8826,N_8753,N_8798);
nor U8827 (N_8827,N_8720,N_8667);
or U8828 (N_8828,N_8681,N_8715);
nor U8829 (N_8829,N_8797,N_8706);
xor U8830 (N_8830,N_8709,N_8704);
xnor U8831 (N_8831,N_8754,N_8684);
nand U8832 (N_8832,N_8714,N_8759);
nand U8833 (N_8833,N_8670,N_8796);
xnor U8834 (N_8834,N_8669,N_8723);
nand U8835 (N_8835,N_8708,N_8770);
nor U8836 (N_8836,N_8719,N_8701);
nor U8837 (N_8837,N_8693,N_8717);
or U8838 (N_8838,N_8710,N_8674);
nand U8839 (N_8839,N_8777,N_8740);
xor U8840 (N_8840,N_8682,N_8785);
or U8841 (N_8841,N_8712,N_8774);
and U8842 (N_8842,N_8767,N_8643);
and U8843 (N_8843,N_8692,N_8738);
and U8844 (N_8844,N_8716,N_8668);
nand U8845 (N_8845,N_8665,N_8695);
xor U8846 (N_8846,N_8735,N_8649);
and U8847 (N_8847,N_8739,N_8658);
nor U8848 (N_8848,N_8673,N_8705);
and U8849 (N_8849,N_8779,N_8736);
xor U8850 (N_8850,N_8758,N_8652);
nor U8851 (N_8851,N_8713,N_8662);
or U8852 (N_8852,N_8677,N_8743);
nor U8853 (N_8853,N_8688,N_8780);
nor U8854 (N_8854,N_8730,N_8760);
xnor U8855 (N_8855,N_8711,N_8657);
nand U8856 (N_8856,N_8781,N_8792);
and U8857 (N_8857,N_8646,N_8787);
or U8858 (N_8858,N_8661,N_8727);
xnor U8859 (N_8859,N_8776,N_8775);
nor U8860 (N_8860,N_8790,N_8694);
xor U8861 (N_8861,N_8741,N_8788);
and U8862 (N_8862,N_8783,N_8768);
xnor U8863 (N_8863,N_8771,N_8772);
nor U8864 (N_8864,N_8748,N_8749);
xor U8865 (N_8865,N_8697,N_8660);
xor U8866 (N_8866,N_8680,N_8653);
nor U8867 (N_8867,N_8784,N_8744);
xor U8868 (N_8868,N_8675,N_8696);
or U8869 (N_8869,N_8683,N_8640);
nor U8870 (N_8870,N_8756,N_8747);
nor U8871 (N_8871,N_8671,N_8689);
or U8872 (N_8872,N_8698,N_8699);
nand U8873 (N_8873,N_8648,N_8654);
nand U8874 (N_8874,N_8678,N_8651);
and U8875 (N_8875,N_8731,N_8676);
xor U8876 (N_8876,N_8791,N_8763);
and U8877 (N_8877,N_8686,N_8757);
xor U8878 (N_8878,N_8769,N_8761);
nor U8879 (N_8879,N_8656,N_8700);
nand U8880 (N_8880,N_8718,N_8657);
nand U8881 (N_8881,N_8684,N_8656);
nand U8882 (N_8882,N_8720,N_8672);
and U8883 (N_8883,N_8794,N_8742);
nand U8884 (N_8884,N_8795,N_8725);
nor U8885 (N_8885,N_8746,N_8678);
or U8886 (N_8886,N_8697,N_8757);
nor U8887 (N_8887,N_8794,N_8687);
nand U8888 (N_8888,N_8799,N_8700);
xor U8889 (N_8889,N_8748,N_8678);
xor U8890 (N_8890,N_8735,N_8710);
nor U8891 (N_8891,N_8671,N_8707);
nand U8892 (N_8892,N_8744,N_8699);
and U8893 (N_8893,N_8662,N_8765);
nand U8894 (N_8894,N_8717,N_8649);
or U8895 (N_8895,N_8652,N_8788);
nor U8896 (N_8896,N_8777,N_8714);
or U8897 (N_8897,N_8674,N_8797);
and U8898 (N_8898,N_8724,N_8713);
nor U8899 (N_8899,N_8761,N_8753);
or U8900 (N_8900,N_8795,N_8655);
nor U8901 (N_8901,N_8656,N_8773);
nand U8902 (N_8902,N_8783,N_8724);
and U8903 (N_8903,N_8716,N_8747);
nand U8904 (N_8904,N_8742,N_8774);
and U8905 (N_8905,N_8772,N_8761);
and U8906 (N_8906,N_8683,N_8651);
and U8907 (N_8907,N_8682,N_8717);
nor U8908 (N_8908,N_8783,N_8757);
xor U8909 (N_8909,N_8711,N_8755);
nor U8910 (N_8910,N_8653,N_8757);
and U8911 (N_8911,N_8752,N_8779);
nand U8912 (N_8912,N_8674,N_8681);
nor U8913 (N_8913,N_8760,N_8710);
or U8914 (N_8914,N_8746,N_8668);
or U8915 (N_8915,N_8674,N_8787);
nand U8916 (N_8916,N_8653,N_8656);
or U8917 (N_8917,N_8744,N_8766);
xnor U8918 (N_8918,N_8723,N_8733);
nand U8919 (N_8919,N_8692,N_8749);
and U8920 (N_8920,N_8728,N_8708);
or U8921 (N_8921,N_8664,N_8773);
nand U8922 (N_8922,N_8779,N_8721);
nand U8923 (N_8923,N_8753,N_8787);
xnor U8924 (N_8924,N_8666,N_8655);
xnor U8925 (N_8925,N_8659,N_8673);
or U8926 (N_8926,N_8661,N_8776);
and U8927 (N_8927,N_8732,N_8664);
nor U8928 (N_8928,N_8799,N_8726);
nor U8929 (N_8929,N_8657,N_8790);
xnor U8930 (N_8930,N_8716,N_8674);
and U8931 (N_8931,N_8712,N_8794);
or U8932 (N_8932,N_8662,N_8677);
nand U8933 (N_8933,N_8664,N_8716);
xnor U8934 (N_8934,N_8648,N_8773);
or U8935 (N_8935,N_8785,N_8653);
and U8936 (N_8936,N_8690,N_8765);
nor U8937 (N_8937,N_8687,N_8731);
xor U8938 (N_8938,N_8651,N_8797);
and U8939 (N_8939,N_8738,N_8776);
xnor U8940 (N_8940,N_8770,N_8677);
xnor U8941 (N_8941,N_8696,N_8678);
xor U8942 (N_8942,N_8685,N_8742);
xnor U8943 (N_8943,N_8768,N_8698);
or U8944 (N_8944,N_8714,N_8778);
and U8945 (N_8945,N_8703,N_8784);
nand U8946 (N_8946,N_8659,N_8786);
nand U8947 (N_8947,N_8743,N_8796);
nand U8948 (N_8948,N_8769,N_8671);
and U8949 (N_8949,N_8645,N_8640);
and U8950 (N_8950,N_8704,N_8726);
or U8951 (N_8951,N_8710,N_8794);
nand U8952 (N_8952,N_8644,N_8688);
nand U8953 (N_8953,N_8649,N_8795);
or U8954 (N_8954,N_8749,N_8720);
or U8955 (N_8955,N_8707,N_8730);
xnor U8956 (N_8956,N_8654,N_8653);
nand U8957 (N_8957,N_8680,N_8641);
xor U8958 (N_8958,N_8705,N_8749);
nor U8959 (N_8959,N_8676,N_8732);
nand U8960 (N_8960,N_8945,N_8893);
nand U8961 (N_8961,N_8901,N_8902);
nand U8962 (N_8962,N_8944,N_8856);
or U8963 (N_8963,N_8952,N_8843);
xor U8964 (N_8964,N_8879,N_8864);
xor U8965 (N_8965,N_8836,N_8829);
or U8966 (N_8966,N_8827,N_8896);
and U8967 (N_8967,N_8905,N_8957);
or U8968 (N_8968,N_8809,N_8823);
nor U8969 (N_8969,N_8848,N_8806);
or U8970 (N_8970,N_8814,N_8835);
nor U8971 (N_8971,N_8953,N_8895);
and U8972 (N_8972,N_8904,N_8873);
nor U8973 (N_8973,N_8840,N_8807);
and U8974 (N_8974,N_8886,N_8825);
xor U8975 (N_8975,N_8851,N_8940);
nand U8976 (N_8976,N_8892,N_8899);
or U8977 (N_8977,N_8815,N_8818);
nor U8978 (N_8978,N_8833,N_8946);
and U8979 (N_8979,N_8919,N_8861);
nor U8980 (N_8980,N_8900,N_8894);
or U8981 (N_8981,N_8800,N_8849);
nor U8982 (N_8982,N_8918,N_8841);
or U8983 (N_8983,N_8819,N_8883);
nor U8984 (N_8984,N_8926,N_8948);
and U8985 (N_8985,N_8871,N_8824);
nor U8986 (N_8986,N_8921,N_8950);
nor U8987 (N_8987,N_8903,N_8942);
nor U8988 (N_8988,N_8949,N_8958);
nand U8989 (N_8989,N_8947,N_8860);
nand U8990 (N_8990,N_8934,N_8804);
or U8991 (N_8991,N_8844,N_8898);
xnor U8992 (N_8992,N_8917,N_8935);
xnor U8993 (N_8993,N_8854,N_8859);
nor U8994 (N_8994,N_8914,N_8846);
xnor U8995 (N_8995,N_8887,N_8909);
nor U8996 (N_8996,N_8868,N_8915);
and U8997 (N_8997,N_8813,N_8925);
nand U8998 (N_8998,N_8938,N_8885);
nor U8999 (N_8999,N_8862,N_8884);
nor U9000 (N_9000,N_8869,N_8801);
nor U9001 (N_9001,N_8954,N_8872);
nand U9002 (N_9002,N_8897,N_8805);
nand U9003 (N_9003,N_8816,N_8910);
or U9004 (N_9004,N_8877,N_8932);
nor U9005 (N_9005,N_8880,N_8924);
nand U9006 (N_9006,N_8955,N_8951);
and U9007 (N_9007,N_8878,N_8817);
nand U9008 (N_9008,N_8930,N_8890);
and U9009 (N_9009,N_8831,N_8839);
nand U9010 (N_9010,N_8876,N_8881);
xnor U9011 (N_9011,N_8838,N_8907);
xnor U9012 (N_9012,N_8845,N_8870);
xnor U9013 (N_9013,N_8874,N_8888);
xor U9014 (N_9014,N_8852,N_8933);
or U9015 (N_9015,N_8891,N_8937);
xor U9016 (N_9016,N_8906,N_8853);
xor U9017 (N_9017,N_8837,N_8865);
or U9018 (N_9018,N_8889,N_8922);
nor U9019 (N_9019,N_8834,N_8857);
or U9020 (N_9020,N_8811,N_8850);
or U9021 (N_9021,N_8821,N_8863);
xnor U9022 (N_9022,N_8858,N_8866);
nand U9023 (N_9023,N_8908,N_8802);
and U9024 (N_9024,N_8943,N_8936);
and U9025 (N_9025,N_8927,N_8847);
nand U9026 (N_9026,N_8822,N_8830);
or U9027 (N_9027,N_8803,N_8928);
nand U9028 (N_9028,N_8959,N_8911);
nand U9029 (N_9029,N_8913,N_8832);
or U9030 (N_9030,N_8956,N_8810);
or U9031 (N_9031,N_8941,N_8939);
xor U9032 (N_9032,N_8867,N_8855);
or U9033 (N_9033,N_8912,N_8828);
nor U9034 (N_9034,N_8808,N_8875);
nand U9035 (N_9035,N_8923,N_8929);
nor U9036 (N_9036,N_8842,N_8920);
nor U9037 (N_9037,N_8820,N_8931);
or U9038 (N_9038,N_8812,N_8916);
nand U9039 (N_9039,N_8882,N_8826);
xor U9040 (N_9040,N_8852,N_8880);
xnor U9041 (N_9041,N_8876,N_8884);
nand U9042 (N_9042,N_8863,N_8824);
xor U9043 (N_9043,N_8908,N_8866);
or U9044 (N_9044,N_8908,N_8905);
xor U9045 (N_9045,N_8849,N_8951);
xor U9046 (N_9046,N_8897,N_8943);
xor U9047 (N_9047,N_8815,N_8916);
nor U9048 (N_9048,N_8911,N_8827);
nand U9049 (N_9049,N_8946,N_8838);
nand U9050 (N_9050,N_8883,N_8848);
nand U9051 (N_9051,N_8868,N_8860);
nor U9052 (N_9052,N_8882,N_8949);
nand U9053 (N_9053,N_8922,N_8924);
nor U9054 (N_9054,N_8850,N_8896);
nor U9055 (N_9055,N_8926,N_8952);
xor U9056 (N_9056,N_8924,N_8948);
nand U9057 (N_9057,N_8869,N_8842);
xnor U9058 (N_9058,N_8814,N_8820);
or U9059 (N_9059,N_8956,N_8831);
and U9060 (N_9060,N_8907,N_8949);
nand U9061 (N_9061,N_8906,N_8857);
nand U9062 (N_9062,N_8926,N_8903);
nor U9063 (N_9063,N_8938,N_8810);
or U9064 (N_9064,N_8854,N_8956);
nor U9065 (N_9065,N_8905,N_8818);
or U9066 (N_9066,N_8817,N_8937);
or U9067 (N_9067,N_8953,N_8802);
nand U9068 (N_9068,N_8888,N_8924);
or U9069 (N_9069,N_8910,N_8810);
nand U9070 (N_9070,N_8928,N_8946);
nor U9071 (N_9071,N_8921,N_8863);
or U9072 (N_9072,N_8882,N_8843);
nor U9073 (N_9073,N_8815,N_8927);
xnor U9074 (N_9074,N_8857,N_8952);
and U9075 (N_9075,N_8905,N_8895);
xnor U9076 (N_9076,N_8838,N_8908);
xnor U9077 (N_9077,N_8951,N_8807);
nand U9078 (N_9078,N_8938,N_8927);
nand U9079 (N_9079,N_8844,N_8902);
or U9080 (N_9080,N_8827,N_8837);
xor U9081 (N_9081,N_8887,N_8916);
xnor U9082 (N_9082,N_8933,N_8825);
nor U9083 (N_9083,N_8845,N_8932);
and U9084 (N_9084,N_8931,N_8898);
nor U9085 (N_9085,N_8821,N_8940);
or U9086 (N_9086,N_8841,N_8864);
or U9087 (N_9087,N_8807,N_8855);
xor U9088 (N_9088,N_8866,N_8854);
xor U9089 (N_9089,N_8933,N_8881);
or U9090 (N_9090,N_8912,N_8825);
or U9091 (N_9091,N_8917,N_8899);
nor U9092 (N_9092,N_8852,N_8957);
xor U9093 (N_9093,N_8866,N_8824);
nor U9094 (N_9094,N_8881,N_8934);
nand U9095 (N_9095,N_8940,N_8910);
or U9096 (N_9096,N_8848,N_8946);
nand U9097 (N_9097,N_8886,N_8826);
nand U9098 (N_9098,N_8851,N_8952);
or U9099 (N_9099,N_8924,N_8891);
xnor U9100 (N_9100,N_8939,N_8935);
nor U9101 (N_9101,N_8883,N_8887);
or U9102 (N_9102,N_8845,N_8888);
nand U9103 (N_9103,N_8945,N_8834);
nand U9104 (N_9104,N_8859,N_8947);
and U9105 (N_9105,N_8884,N_8892);
xor U9106 (N_9106,N_8956,N_8851);
nor U9107 (N_9107,N_8860,N_8894);
nand U9108 (N_9108,N_8829,N_8850);
nand U9109 (N_9109,N_8937,N_8922);
or U9110 (N_9110,N_8913,N_8825);
nor U9111 (N_9111,N_8818,N_8810);
and U9112 (N_9112,N_8895,N_8930);
xnor U9113 (N_9113,N_8800,N_8912);
nor U9114 (N_9114,N_8928,N_8955);
or U9115 (N_9115,N_8887,N_8934);
nor U9116 (N_9116,N_8863,N_8849);
and U9117 (N_9117,N_8950,N_8810);
and U9118 (N_9118,N_8952,N_8822);
and U9119 (N_9119,N_8938,N_8895);
or U9120 (N_9120,N_9051,N_8965);
xor U9121 (N_9121,N_8967,N_9062);
or U9122 (N_9122,N_9021,N_9115);
nand U9123 (N_9123,N_9011,N_8987);
and U9124 (N_9124,N_8976,N_9081);
and U9125 (N_9125,N_9056,N_8964);
xor U9126 (N_9126,N_9028,N_9007);
nand U9127 (N_9127,N_9009,N_8990);
and U9128 (N_9128,N_9111,N_9096);
xnor U9129 (N_9129,N_9116,N_9080);
nor U9130 (N_9130,N_9084,N_9068);
nand U9131 (N_9131,N_8985,N_8984);
nor U9132 (N_9132,N_8973,N_9103);
xor U9133 (N_9133,N_9057,N_9061);
nand U9134 (N_9134,N_9088,N_9101);
or U9135 (N_9135,N_9064,N_9041);
nand U9136 (N_9136,N_9082,N_9054);
or U9137 (N_9137,N_9053,N_9038);
nand U9138 (N_9138,N_9107,N_9099);
or U9139 (N_9139,N_9024,N_9070);
or U9140 (N_9140,N_8995,N_9117);
nand U9141 (N_9141,N_9002,N_9067);
xor U9142 (N_9142,N_9044,N_9016);
and U9143 (N_9143,N_9055,N_9093);
nand U9144 (N_9144,N_9045,N_9098);
nand U9145 (N_9145,N_9005,N_9076);
and U9146 (N_9146,N_8988,N_9105);
nor U9147 (N_9147,N_9008,N_9106);
and U9148 (N_9148,N_9110,N_9029);
nand U9149 (N_9149,N_9074,N_9050);
nor U9150 (N_9150,N_9071,N_9059);
or U9151 (N_9151,N_9060,N_9034);
nor U9152 (N_9152,N_8991,N_9047);
xor U9153 (N_9153,N_9040,N_8997);
nand U9154 (N_9154,N_9087,N_9036);
or U9155 (N_9155,N_9023,N_9119);
or U9156 (N_9156,N_9118,N_9026);
xnor U9157 (N_9157,N_9043,N_9025);
and U9158 (N_9158,N_8996,N_9073);
and U9159 (N_9159,N_9058,N_8977);
nor U9160 (N_9160,N_8978,N_9018);
or U9161 (N_9161,N_9046,N_9048);
and U9162 (N_9162,N_8981,N_9001);
or U9163 (N_9163,N_9027,N_9108);
nand U9164 (N_9164,N_9042,N_9004);
xnor U9165 (N_9165,N_9019,N_9014);
xor U9166 (N_9166,N_9097,N_9109);
nor U9167 (N_9167,N_8966,N_9006);
xnor U9168 (N_9168,N_9072,N_9033);
or U9169 (N_9169,N_9013,N_8986);
nand U9170 (N_9170,N_8975,N_9075);
and U9171 (N_9171,N_8971,N_8998);
nor U9172 (N_9172,N_9078,N_8972);
xor U9173 (N_9173,N_9015,N_9083);
nand U9174 (N_9174,N_8983,N_8993);
nand U9175 (N_9175,N_8979,N_9079);
or U9176 (N_9176,N_8994,N_9095);
xor U9177 (N_9177,N_8989,N_9037);
xor U9178 (N_9178,N_9065,N_9000);
xnor U9179 (N_9179,N_9030,N_8960);
or U9180 (N_9180,N_9114,N_9035);
and U9181 (N_9181,N_8969,N_9003);
xor U9182 (N_9182,N_9089,N_9049);
nand U9183 (N_9183,N_8970,N_9094);
or U9184 (N_9184,N_8992,N_9010);
or U9185 (N_9185,N_9100,N_8968);
nor U9186 (N_9186,N_8982,N_8999);
nor U9187 (N_9187,N_8962,N_9032);
or U9188 (N_9188,N_9092,N_9077);
nor U9189 (N_9189,N_9113,N_9104);
xnor U9190 (N_9190,N_8963,N_9017);
nor U9191 (N_9191,N_9012,N_9085);
nand U9192 (N_9192,N_9086,N_9091);
or U9193 (N_9193,N_8961,N_9063);
nor U9194 (N_9194,N_9069,N_9066);
xor U9195 (N_9195,N_9031,N_9022);
xnor U9196 (N_9196,N_9020,N_8974);
or U9197 (N_9197,N_9052,N_8980);
xnor U9198 (N_9198,N_9090,N_9102);
nand U9199 (N_9199,N_9112,N_9039);
xnor U9200 (N_9200,N_9057,N_9085);
and U9201 (N_9201,N_9053,N_9115);
xnor U9202 (N_9202,N_9106,N_9024);
nand U9203 (N_9203,N_9045,N_8999);
or U9204 (N_9204,N_9093,N_9001);
xnor U9205 (N_9205,N_9043,N_9000);
and U9206 (N_9206,N_9064,N_9006);
nor U9207 (N_9207,N_9106,N_9090);
and U9208 (N_9208,N_9084,N_9087);
and U9209 (N_9209,N_8993,N_9016);
xor U9210 (N_9210,N_9001,N_9056);
and U9211 (N_9211,N_9093,N_9048);
or U9212 (N_9212,N_9070,N_8965);
nor U9213 (N_9213,N_9072,N_9107);
xnor U9214 (N_9214,N_9028,N_9080);
nor U9215 (N_9215,N_8996,N_9087);
and U9216 (N_9216,N_8985,N_8993);
nor U9217 (N_9217,N_9093,N_9019);
or U9218 (N_9218,N_9019,N_9106);
nor U9219 (N_9219,N_8978,N_9008);
and U9220 (N_9220,N_8972,N_9024);
or U9221 (N_9221,N_9078,N_9049);
and U9222 (N_9222,N_9075,N_9002);
nand U9223 (N_9223,N_8980,N_9015);
xor U9224 (N_9224,N_9036,N_9001);
nor U9225 (N_9225,N_9041,N_9073);
or U9226 (N_9226,N_9084,N_9054);
nor U9227 (N_9227,N_9115,N_9069);
or U9228 (N_9228,N_9057,N_8968);
nor U9229 (N_9229,N_9068,N_9036);
nand U9230 (N_9230,N_9104,N_9027);
and U9231 (N_9231,N_9099,N_9045);
nand U9232 (N_9232,N_8970,N_9095);
xor U9233 (N_9233,N_9034,N_8978);
or U9234 (N_9234,N_9087,N_8992);
xnor U9235 (N_9235,N_9000,N_8998);
nand U9236 (N_9236,N_9007,N_8987);
and U9237 (N_9237,N_9015,N_9106);
or U9238 (N_9238,N_9034,N_8965);
nand U9239 (N_9239,N_9010,N_9099);
nor U9240 (N_9240,N_9011,N_9031);
or U9241 (N_9241,N_8990,N_9015);
and U9242 (N_9242,N_8978,N_9028);
nor U9243 (N_9243,N_9014,N_8973);
nand U9244 (N_9244,N_8984,N_8966);
or U9245 (N_9245,N_9118,N_8989);
nand U9246 (N_9246,N_8984,N_9040);
or U9247 (N_9247,N_9084,N_9106);
xnor U9248 (N_9248,N_9073,N_8984);
nand U9249 (N_9249,N_9088,N_9059);
and U9250 (N_9250,N_9034,N_9016);
or U9251 (N_9251,N_8998,N_9074);
or U9252 (N_9252,N_9032,N_9062);
nor U9253 (N_9253,N_9043,N_8995);
nand U9254 (N_9254,N_9001,N_9029);
nor U9255 (N_9255,N_9017,N_9111);
nand U9256 (N_9256,N_9051,N_9011);
or U9257 (N_9257,N_9034,N_9041);
nor U9258 (N_9258,N_9060,N_8971);
nor U9259 (N_9259,N_8976,N_9089);
or U9260 (N_9260,N_8973,N_9004);
xor U9261 (N_9261,N_9083,N_9040);
or U9262 (N_9262,N_9090,N_8981);
and U9263 (N_9263,N_9061,N_8994);
xnor U9264 (N_9264,N_9079,N_9100);
and U9265 (N_9265,N_9118,N_9002);
nor U9266 (N_9266,N_8991,N_8975);
nand U9267 (N_9267,N_9046,N_8994);
xnor U9268 (N_9268,N_8966,N_9010);
nand U9269 (N_9269,N_9037,N_9099);
or U9270 (N_9270,N_9073,N_8998);
nor U9271 (N_9271,N_9084,N_8965);
xnor U9272 (N_9272,N_9082,N_9044);
and U9273 (N_9273,N_8984,N_9033);
xnor U9274 (N_9274,N_9098,N_8983);
nor U9275 (N_9275,N_9061,N_9074);
or U9276 (N_9276,N_9088,N_9040);
and U9277 (N_9277,N_8981,N_9039);
or U9278 (N_9278,N_8973,N_9032);
and U9279 (N_9279,N_8978,N_8981);
xor U9280 (N_9280,N_9128,N_9239);
or U9281 (N_9281,N_9224,N_9244);
xor U9282 (N_9282,N_9220,N_9175);
nand U9283 (N_9283,N_9135,N_9237);
xnor U9284 (N_9284,N_9173,N_9161);
or U9285 (N_9285,N_9156,N_9136);
xor U9286 (N_9286,N_9236,N_9124);
nand U9287 (N_9287,N_9160,N_9186);
or U9288 (N_9288,N_9273,N_9142);
xnor U9289 (N_9289,N_9200,N_9232);
nand U9290 (N_9290,N_9197,N_9246);
xor U9291 (N_9291,N_9223,N_9176);
nor U9292 (N_9292,N_9169,N_9209);
nand U9293 (N_9293,N_9155,N_9205);
xnor U9294 (N_9294,N_9201,N_9153);
xnor U9295 (N_9295,N_9148,N_9178);
xnor U9296 (N_9296,N_9274,N_9183);
nor U9297 (N_9297,N_9171,N_9269);
nor U9298 (N_9298,N_9132,N_9133);
and U9299 (N_9299,N_9249,N_9179);
nand U9300 (N_9300,N_9177,N_9241);
nand U9301 (N_9301,N_9272,N_9130);
nor U9302 (N_9302,N_9131,N_9255);
xor U9303 (N_9303,N_9193,N_9222);
or U9304 (N_9304,N_9143,N_9234);
xnor U9305 (N_9305,N_9191,N_9260);
nand U9306 (N_9306,N_9259,N_9151);
and U9307 (N_9307,N_9154,N_9158);
nor U9308 (N_9308,N_9270,N_9267);
and U9309 (N_9309,N_9219,N_9262);
xnor U9310 (N_9310,N_9229,N_9121);
and U9311 (N_9311,N_9170,N_9276);
and U9312 (N_9312,N_9181,N_9214);
nand U9313 (N_9313,N_9189,N_9264);
xor U9314 (N_9314,N_9275,N_9163);
nor U9315 (N_9315,N_9231,N_9206);
xnor U9316 (N_9316,N_9167,N_9164);
nand U9317 (N_9317,N_9226,N_9213);
xor U9318 (N_9318,N_9159,N_9196);
xnor U9319 (N_9319,N_9221,N_9138);
nand U9320 (N_9320,N_9217,N_9247);
and U9321 (N_9321,N_9194,N_9125);
or U9322 (N_9322,N_9278,N_9207);
nor U9323 (N_9323,N_9187,N_9180);
or U9324 (N_9324,N_9251,N_9218);
nand U9325 (N_9325,N_9225,N_9242);
nor U9326 (N_9326,N_9185,N_9238);
nor U9327 (N_9327,N_9266,N_9126);
xnor U9328 (N_9328,N_9122,N_9174);
and U9329 (N_9329,N_9145,N_9139);
xor U9330 (N_9330,N_9199,N_9172);
xor U9331 (N_9331,N_9263,N_9257);
nor U9332 (N_9332,N_9190,N_9215);
or U9333 (N_9333,N_9252,N_9265);
or U9334 (N_9334,N_9123,N_9157);
and U9335 (N_9335,N_9208,N_9134);
or U9336 (N_9336,N_9230,N_9258);
and U9337 (N_9337,N_9198,N_9243);
and U9338 (N_9338,N_9168,N_9150);
xor U9339 (N_9339,N_9245,N_9250);
nor U9340 (N_9340,N_9152,N_9235);
or U9341 (N_9341,N_9228,N_9147);
xnor U9342 (N_9342,N_9204,N_9253);
nor U9343 (N_9343,N_9144,N_9127);
nor U9344 (N_9344,N_9129,N_9146);
or U9345 (N_9345,N_9202,N_9233);
nand U9346 (N_9346,N_9254,N_9184);
and U9347 (N_9347,N_9268,N_9166);
nor U9348 (N_9348,N_9149,N_9256);
and U9349 (N_9349,N_9195,N_9240);
or U9350 (N_9350,N_9137,N_9216);
nor U9351 (N_9351,N_9279,N_9261);
nor U9352 (N_9352,N_9182,N_9248);
xor U9353 (N_9353,N_9162,N_9192);
nor U9354 (N_9354,N_9277,N_9203);
xnor U9355 (N_9355,N_9120,N_9211);
or U9356 (N_9356,N_9140,N_9188);
nand U9357 (N_9357,N_9227,N_9210);
xor U9358 (N_9358,N_9165,N_9141);
and U9359 (N_9359,N_9212,N_9271);
nor U9360 (N_9360,N_9274,N_9165);
nor U9361 (N_9361,N_9155,N_9127);
nand U9362 (N_9362,N_9186,N_9155);
nor U9363 (N_9363,N_9271,N_9196);
nand U9364 (N_9364,N_9204,N_9230);
or U9365 (N_9365,N_9213,N_9270);
or U9366 (N_9366,N_9262,N_9129);
xor U9367 (N_9367,N_9220,N_9180);
xnor U9368 (N_9368,N_9265,N_9145);
nor U9369 (N_9369,N_9276,N_9144);
and U9370 (N_9370,N_9198,N_9180);
nor U9371 (N_9371,N_9272,N_9251);
nor U9372 (N_9372,N_9238,N_9258);
xor U9373 (N_9373,N_9232,N_9228);
nand U9374 (N_9374,N_9212,N_9141);
or U9375 (N_9375,N_9244,N_9147);
or U9376 (N_9376,N_9147,N_9205);
or U9377 (N_9377,N_9222,N_9173);
xnor U9378 (N_9378,N_9154,N_9239);
nor U9379 (N_9379,N_9193,N_9250);
nand U9380 (N_9380,N_9215,N_9209);
nand U9381 (N_9381,N_9199,N_9179);
nor U9382 (N_9382,N_9170,N_9178);
xor U9383 (N_9383,N_9251,N_9179);
or U9384 (N_9384,N_9172,N_9177);
and U9385 (N_9385,N_9246,N_9182);
nor U9386 (N_9386,N_9145,N_9212);
xnor U9387 (N_9387,N_9275,N_9164);
xnor U9388 (N_9388,N_9138,N_9268);
and U9389 (N_9389,N_9144,N_9254);
xor U9390 (N_9390,N_9197,N_9251);
nor U9391 (N_9391,N_9150,N_9218);
or U9392 (N_9392,N_9131,N_9269);
or U9393 (N_9393,N_9132,N_9194);
nor U9394 (N_9394,N_9246,N_9230);
or U9395 (N_9395,N_9276,N_9273);
and U9396 (N_9396,N_9248,N_9235);
and U9397 (N_9397,N_9268,N_9159);
nand U9398 (N_9398,N_9279,N_9230);
nand U9399 (N_9399,N_9188,N_9154);
nand U9400 (N_9400,N_9244,N_9148);
nor U9401 (N_9401,N_9139,N_9236);
nand U9402 (N_9402,N_9193,N_9195);
nand U9403 (N_9403,N_9270,N_9156);
or U9404 (N_9404,N_9210,N_9258);
or U9405 (N_9405,N_9254,N_9229);
xnor U9406 (N_9406,N_9257,N_9275);
and U9407 (N_9407,N_9218,N_9236);
or U9408 (N_9408,N_9274,N_9204);
nor U9409 (N_9409,N_9230,N_9133);
xor U9410 (N_9410,N_9234,N_9176);
nand U9411 (N_9411,N_9271,N_9257);
nand U9412 (N_9412,N_9227,N_9142);
nor U9413 (N_9413,N_9130,N_9128);
or U9414 (N_9414,N_9171,N_9239);
nor U9415 (N_9415,N_9167,N_9129);
and U9416 (N_9416,N_9230,N_9209);
or U9417 (N_9417,N_9206,N_9249);
or U9418 (N_9418,N_9146,N_9192);
nor U9419 (N_9419,N_9218,N_9239);
xor U9420 (N_9420,N_9267,N_9207);
nand U9421 (N_9421,N_9147,N_9178);
nor U9422 (N_9422,N_9196,N_9164);
and U9423 (N_9423,N_9134,N_9254);
nand U9424 (N_9424,N_9278,N_9155);
and U9425 (N_9425,N_9130,N_9129);
xor U9426 (N_9426,N_9153,N_9200);
and U9427 (N_9427,N_9265,N_9183);
and U9428 (N_9428,N_9240,N_9256);
xnor U9429 (N_9429,N_9134,N_9182);
nand U9430 (N_9430,N_9216,N_9274);
nand U9431 (N_9431,N_9269,N_9125);
nand U9432 (N_9432,N_9132,N_9200);
xor U9433 (N_9433,N_9169,N_9249);
and U9434 (N_9434,N_9208,N_9279);
xor U9435 (N_9435,N_9215,N_9275);
and U9436 (N_9436,N_9242,N_9134);
nand U9437 (N_9437,N_9279,N_9180);
xor U9438 (N_9438,N_9236,N_9132);
or U9439 (N_9439,N_9261,N_9267);
xnor U9440 (N_9440,N_9364,N_9313);
or U9441 (N_9441,N_9355,N_9308);
nand U9442 (N_9442,N_9370,N_9283);
and U9443 (N_9443,N_9390,N_9292);
or U9444 (N_9444,N_9327,N_9360);
nor U9445 (N_9445,N_9321,N_9282);
nand U9446 (N_9446,N_9286,N_9324);
xor U9447 (N_9447,N_9307,N_9394);
xnor U9448 (N_9448,N_9330,N_9369);
or U9449 (N_9449,N_9317,N_9302);
or U9450 (N_9450,N_9410,N_9335);
nor U9451 (N_9451,N_9357,N_9391);
and U9452 (N_9452,N_9366,N_9363);
and U9453 (N_9453,N_9295,N_9289);
nand U9454 (N_9454,N_9425,N_9306);
nand U9455 (N_9455,N_9381,N_9359);
nor U9456 (N_9456,N_9436,N_9427);
nand U9457 (N_9457,N_9431,N_9429);
or U9458 (N_9458,N_9392,N_9416);
or U9459 (N_9459,N_9382,N_9304);
nand U9460 (N_9460,N_9393,N_9400);
or U9461 (N_9461,N_9349,N_9426);
xor U9462 (N_9462,N_9379,N_9389);
nor U9463 (N_9463,N_9388,N_9341);
nand U9464 (N_9464,N_9417,N_9344);
or U9465 (N_9465,N_9418,N_9409);
nor U9466 (N_9466,N_9316,N_9420);
xnor U9467 (N_9467,N_9377,N_9315);
nor U9468 (N_9468,N_9354,N_9339);
or U9469 (N_9469,N_9385,N_9280);
xor U9470 (N_9470,N_9299,N_9296);
xor U9471 (N_9471,N_9380,N_9326);
xor U9472 (N_9472,N_9323,N_9343);
xor U9473 (N_9473,N_9411,N_9438);
nor U9474 (N_9474,N_9348,N_9293);
nand U9475 (N_9475,N_9414,N_9333);
and U9476 (N_9476,N_9421,N_9432);
nand U9477 (N_9477,N_9309,N_9372);
nor U9478 (N_9478,N_9297,N_9350);
nand U9479 (N_9479,N_9331,N_9430);
nor U9480 (N_9480,N_9378,N_9374);
nor U9481 (N_9481,N_9395,N_9287);
xor U9482 (N_9482,N_9361,N_9373);
and U9483 (N_9483,N_9401,N_9294);
nand U9484 (N_9484,N_9435,N_9328);
or U9485 (N_9485,N_9310,N_9383);
and U9486 (N_9486,N_9371,N_9437);
nand U9487 (N_9487,N_9403,N_9358);
nor U9488 (N_9488,N_9386,N_9329);
nand U9489 (N_9489,N_9281,N_9291);
and U9490 (N_9490,N_9413,N_9424);
nor U9491 (N_9491,N_9314,N_9322);
nand U9492 (N_9492,N_9334,N_9347);
nor U9493 (N_9493,N_9408,N_9303);
xnor U9494 (N_9494,N_9422,N_9415);
nor U9495 (N_9495,N_9301,N_9311);
nor U9496 (N_9496,N_9407,N_9397);
and U9497 (N_9497,N_9338,N_9362);
and U9498 (N_9498,N_9434,N_9412);
xor U9499 (N_9499,N_9340,N_9305);
xor U9500 (N_9500,N_9433,N_9337);
nand U9501 (N_9501,N_9368,N_9290);
nand U9502 (N_9502,N_9365,N_9351);
nor U9503 (N_9503,N_9399,N_9439);
and U9504 (N_9504,N_9345,N_9353);
or U9505 (N_9505,N_9428,N_9356);
nand U9506 (N_9506,N_9325,N_9300);
nor U9507 (N_9507,N_9398,N_9375);
and U9508 (N_9508,N_9318,N_9402);
or U9509 (N_9509,N_9406,N_9367);
nor U9510 (N_9510,N_9312,N_9342);
or U9511 (N_9511,N_9288,N_9319);
nand U9512 (N_9512,N_9404,N_9396);
nand U9513 (N_9513,N_9423,N_9332);
xnor U9514 (N_9514,N_9387,N_9320);
or U9515 (N_9515,N_9346,N_9352);
xor U9516 (N_9516,N_9284,N_9405);
xnor U9517 (N_9517,N_9285,N_9376);
nor U9518 (N_9518,N_9384,N_9336);
xnor U9519 (N_9519,N_9298,N_9419);
nand U9520 (N_9520,N_9326,N_9387);
nor U9521 (N_9521,N_9410,N_9397);
and U9522 (N_9522,N_9356,N_9283);
xnor U9523 (N_9523,N_9409,N_9348);
xnor U9524 (N_9524,N_9323,N_9432);
or U9525 (N_9525,N_9397,N_9331);
nand U9526 (N_9526,N_9296,N_9335);
and U9527 (N_9527,N_9318,N_9290);
nor U9528 (N_9528,N_9328,N_9389);
nand U9529 (N_9529,N_9289,N_9378);
or U9530 (N_9530,N_9323,N_9326);
nand U9531 (N_9531,N_9345,N_9323);
xor U9532 (N_9532,N_9422,N_9402);
or U9533 (N_9533,N_9407,N_9289);
xor U9534 (N_9534,N_9413,N_9428);
and U9535 (N_9535,N_9383,N_9403);
nand U9536 (N_9536,N_9370,N_9308);
and U9537 (N_9537,N_9362,N_9378);
nor U9538 (N_9538,N_9367,N_9297);
or U9539 (N_9539,N_9415,N_9404);
xnor U9540 (N_9540,N_9402,N_9352);
and U9541 (N_9541,N_9325,N_9399);
nor U9542 (N_9542,N_9423,N_9393);
nand U9543 (N_9543,N_9400,N_9298);
and U9544 (N_9544,N_9352,N_9421);
or U9545 (N_9545,N_9285,N_9322);
nand U9546 (N_9546,N_9386,N_9391);
xor U9547 (N_9547,N_9425,N_9285);
xor U9548 (N_9548,N_9289,N_9300);
and U9549 (N_9549,N_9438,N_9345);
or U9550 (N_9550,N_9342,N_9432);
and U9551 (N_9551,N_9404,N_9365);
or U9552 (N_9552,N_9432,N_9327);
and U9553 (N_9553,N_9365,N_9325);
nand U9554 (N_9554,N_9306,N_9391);
and U9555 (N_9555,N_9428,N_9340);
and U9556 (N_9556,N_9374,N_9389);
and U9557 (N_9557,N_9374,N_9345);
nand U9558 (N_9558,N_9367,N_9293);
or U9559 (N_9559,N_9320,N_9339);
or U9560 (N_9560,N_9435,N_9358);
nand U9561 (N_9561,N_9352,N_9432);
or U9562 (N_9562,N_9346,N_9330);
nor U9563 (N_9563,N_9416,N_9353);
nand U9564 (N_9564,N_9302,N_9427);
xnor U9565 (N_9565,N_9400,N_9408);
and U9566 (N_9566,N_9351,N_9383);
or U9567 (N_9567,N_9330,N_9391);
nand U9568 (N_9568,N_9430,N_9434);
nor U9569 (N_9569,N_9329,N_9395);
xnor U9570 (N_9570,N_9429,N_9332);
nor U9571 (N_9571,N_9348,N_9299);
and U9572 (N_9572,N_9411,N_9439);
and U9573 (N_9573,N_9383,N_9311);
or U9574 (N_9574,N_9420,N_9317);
or U9575 (N_9575,N_9331,N_9389);
and U9576 (N_9576,N_9412,N_9321);
or U9577 (N_9577,N_9376,N_9349);
nand U9578 (N_9578,N_9336,N_9389);
xnor U9579 (N_9579,N_9409,N_9337);
nor U9580 (N_9580,N_9315,N_9286);
xnor U9581 (N_9581,N_9327,N_9323);
nand U9582 (N_9582,N_9415,N_9331);
nand U9583 (N_9583,N_9399,N_9305);
nand U9584 (N_9584,N_9373,N_9309);
xnor U9585 (N_9585,N_9432,N_9398);
nor U9586 (N_9586,N_9365,N_9362);
nor U9587 (N_9587,N_9353,N_9319);
nand U9588 (N_9588,N_9360,N_9330);
and U9589 (N_9589,N_9420,N_9296);
or U9590 (N_9590,N_9329,N_9302);
or U9591 (N_9591,N_9392,N_9302);
or U9592 (N_9592,N_9395,N_9294);
or U9593 (N_9593,N_9383,N_9357);
nor U9594 (N_9594,N_9426,N_9358);
nor U9595 (N_9595,N_9403,N_9368);
or U9596 (N_9596,N_9323,N_9324);
xor U9597 (N_9597,N_9376,N_9357);
and U9598 (N_9598,N_9432,N_9329);
nand U9599 (N_9599,N_9421,N_9396);
and U9600 (N_9600,N_9570,N_9598);
xor U9601 (N_9601,N_9504,N_9554);
nand U9602 (N_9602,N_9488,N_9569);
and U9603 (N_9603,N_9454,N_9555);
nor U9604 (N_9604,N_9580,N_9517);
nand U9605 (N_9605,N_9553,N_9465);
and U9606 (N_9606,N_9571,N_9591);
or U9607 (N_9607,N_9584,N_9448);
xor U9608 (N_9608,N_9452,N_9573);
nand U9609 (N_9609,N_9519,N_9544);
or U9610 (N_9610,N_9466,N_9581);
xnor U9611 (N_9611,N_9560,N_9552);
nor U9612 (N_9612,N_9493,N_9518);
or U9613 (N_9613,N_9523,N_9509);
nor U9614 (N_9614,N_9542,N_9576);
nor U9615 (N_9615,N_9478,N_9530);
or U9616 (N_9616,N_9533,N_9582);
nor U9617 (N_9617,N_9513,N_9541);
or U9618 (N_9618,N_9521,N_9492);
nor U9619 (N_9619,N_9597,N_9549);
nor U9620 (N_9620,N_9461,N_9443);
and U9621 (N_9621,N_9477,N_9540);
or U9622 (N_9622,N_9498,N_9506);
and U9623 (N_9623,N_9494,N_9497);
xnor U9624 (N_9624,N_9588,N_9495);
xnor U9625 (N_9625,N_9470,N_9459);
nand U9626 (N_9626,N_9496,N_9473);
nand U9627 (N_9627,N_9535,N_9468);
nand U9628 (N_9628,N_9464,N_9550);
xnor U9629 (N_9629,N_9455,N_9579);
nor U9630 (N_9630,N_9556,N_9456);
and U9631 (N_9631,N_9536,N_9528);
xnor U9632 (N_9632,N_9480,N_9472);
and U9633 (N_9633,N_9514,N_9537);
nor U9634 (N_9634,N_9475,N_9564);
nor U9635 (N_9635,N_9534,N_9460);
nand U9636 (N_9636,N_9462,N_9515);
nor U9637 (N_9637,N_9561,N_9444);
nand U9638 (N_9638,N_9594,N_9503);
and U9639 (N_9639,N_9551,N_9527);
and U9640 (N_9640,N_9538,N_9512);
nor U9641 (N_9641,N_9463,N_9562);
xnor U9642 (N_9642,N_9568,N_9440);
and U9643 (N_9643,N_9489,N_9511);
or U9644 (N_9644,N_9445,N_9547);
nand U9645 (N_9645,N_9575,N_9479);
nand U9646 (N_9646,N_9502,N_9557);
or U9647 (N_9647,N_9545,N_9508);
nor U9648 (N_9648,N_9548,N_9599);
and U9649 (N_9649,N_9520,N_9563);
xor U9650 (N_9650,N_9500,N_9543);
xor U9651 (N_9651,N_9487,N_9590);
nand U9652 (N_9652,N_9469,N_9450);
nor U9653 (N_9653,N_9578,N_9446);
xnor U9654 (N_9654,N_9572,N_9451);
and U9655 (N_9655,N_9583,N_9586);
nand U9656 (N_9656,N_9484,N_9565);
or U9657 (N_9657,N_9467,N_9458);
or U9658 (N_9658,N_9505,N_9510);
and U9659 (N_9659,N_9566,N_9592);
and U9660 (N_9660,N_9526,N_9593);
and U9661 (N_9661,N_9474,N_9524);
or U9662 (N_9662,N_9589,N_9574);
xnor U9663 (N_9663,N_9499,N_9587);
or U9664 (N_9664,N_9471,N_9485);
xnor U9665 (N_9665,N_9539,N_9559);
nand U9666 (N_9666,N_9585,N_9447);
nand U9667 (N_9667,N_9516,N_9577);
and U9668 (N_9668,N_9501,N_9529);
nor U9669 (N_9669,N_9507,N_9546);
nand U9670 (N_9670,N_9532,N_9457);
nor U9671 (N_9671,N_9596,N_9531);
xor U9672 (N_9672,N_9442,N_9449);
xnor U9673 (N_9673,N_9486,N_9522);
nor U9674 (N_9674,N_9595,N_9490);
or U9675 (N_9675,N_9482,N_9567);
and U9676 (N_9676,N_9525,N_9491);
or U9677 (N_9677,N_9558,N_9441);
and U9678 (N_9678,N_9476,N_9453);
xor U9679 (N_9679,N_9483,N_9481);
or U9680 (N_9680,N_9584,N_9576);
or U9681 (N_9681,N_9538,N_9442);
nand U9682 (N_9682,N_9583,N_9568);
or U9683 (N_9683,N_9568,N_9555);
nor U9684 (N_9684,N_9536,N_9493);
or U9685 (N_9685,N_9542,N_9564);
nand U9686 (N_9686,N_9541,N_9510);
nand U9687 (N_9687,N_9599,N_9482);
or U9688 (N_9688,N_9571,N_9491);
nand U9689 (N_9689,N_9528,N_9589);
and U9690 (N_9690,N_9526,N_9578);
xnor U9691 (N_9691,N_9582,N_9443);
or U9692 (N_9692,N_9575,N_9588);
xnor U9693 (N_9693,N_9499,N_9456);
nor U9694 (N_9694,N_9570,N_9589);
xnor U9695 (N_9695,N_9524,N_9527);
nor U9696 (N_9696,N_9444,N_9538);
xnor U9697 (N_9697,N_9586,N_9463);
nand U9698 (N_9698,N_9464,N_9513);
nor U9699 (N_9699,N_9473,N_9519);
or U9700 (N_9700,N_9446,N_9496);
or U9701 (N_9701,N_9490,N_9516);
nor U9702 (N_9702,N_9550,N_9596);
nand U9703 (N_9703,N_9545,N_9449);
or U9704 (N_9704,N_9551,N_9528);
nor U9705 (N_9705,N_9495,N_9486);
nand U9706 (N_9706,N_9599,N_9504);
nor U9707 (N_9707,N_9561,N_9531);
nor U9708 (N_9708,N_9454,N_9598);
or U9709 (N_9709,N_9579,N_9504);
nor U9710 (N_9710,N_9514,N_9586);
nor U9711 (N_9711,N_9513,N_9458);
nor U9712 (N_9712,N_9448,N_9541);
nand U9713 (N_9713,N_9490,N_9504);
nor U9714 (N_9714,N_9590,N_9486);
xor U9715 (N_9715,N_9550,N_9546);
xnor U9716 (N_9716,N_9443,N_9485);
or U9717 (N_9717,N_9513,N_9533);
nor U9718 (N_9718,N_9559,N_9549);
nand U9719 (N_9719,N_9529,N_9496);
xnor U9720 (N_9720,N_9460,N_9524);
and U9721 (N_9721,N_9566,N_9595);
nand U9722 (N_9722,N_9515,N_9595);
nand U9723 (N_9723,N_9500,N_9480);
or U9724 (N_9724,N_9484,N_9513);
nor U9725 (N_9725,N_9575,N_9516);
or U9726 (N_9726,N_9589,N_9559);
and U9727 (N_9727,N_9527,N_9479);
xnor U9728 (N_9728,N_9555,N_9584);
or U9729 (N_9729,N_9556,N_9565);
and U9730 (N_9730,N_9482,N_9529);
nor U9731 (N_9731,N_9589,N_9592);
and U9732 (N_9732,N_9512,N_9511);
and U9733 (N_9733,N_9540,N_9449);
or U9734 (N_9734,N_9496,N_9542);
nand U9735 (N_9735,N_9468,N_9444);
nor U9736 (N_9736,N_9488,N_9545);
xnor U9737 (N_9737,N_9452,N_9539);
and U9738 (N_9738,N_9572,N_9499);
nand U9739 (N_9739,N_9575,N_9538);
nand U9740 (N_9740,N_9521,N_9501);
and U9741 (N_9741,N_9465,N_9495);
nor U9742 (N_9742,N_9587,N_9511);
nand U9743 (N_9743,N_9498,N_9560);
and U9744 (N_9744,N_9489,N_9545);
nor U9745 (N_9745,N_9558,N_9502);
or U9746 (N_9746,N_9470,N_9495);
nand U9747 (N_9747,N_9559,N_9493);
or U9748 (N_9748,N_9517,N_9462);
nand U9749 (N_9749,N_9490,N_9522);
xor U9750 (N_9750,N_9442,N_9458);
or U9751 (N_9751,N_9464,N_9484);
or U9752 (N_9752,N_9566,N_9511);
xor U9753 (N_9753,N_9552,N_9466);
nor U9754 (N_9754,N_9536,N_9519);
and U9755 (N_9755,N_9515,N_9513);
nor U9756 (N_9756,N_9595,N_9513);
nor U9757 (N_9757,N_9556,N_9448);
or U9758 (N_9758,N_9472,N_9505);
xor U9759 (N_9759,N_9513,N_9507);
nor U9760 (N_9760,N_9752,N_9699);
xor U9761 (N_9761,N_9663,N_9736);
and U9762 (N_9762,N_9708,N_9653);
or U9763 (N_9763,N_9735,N_9737);
and U9764 (N_9764,N_9624,N_9739);
nor U9765 (N_9765,N_9647,N_9727);
and U9766 (N_9766,N_9731,N_9628);
xnor U9767 (N_9767,N_9668,N_9648);
xnor U9768 (N_9768,N_9703,N_9645);
nand U9769 (N_9769,N_9720,N_9675);
and U9770 (N_9770,N_9695,N_9664);
or U9771 (N_9771,N_9758,N_9693);
and U9772 (N_9772,N_9747,N_9607);
and U9773 (N_9773,N_9618,N_9714);
nor U9774 (N_9774,N_9610,N_9751);
and U9775 (N_9775,N_9682,N_9712);
or U9776 (N_9776,N_9632,N_9723);
and U9777 (N_9777,N_9603,N_9621);
xnor U9778 (N_9778,N_9608,N_9696);
or U9779 (N_9779,N_9717,N_9754);
xnor U9780 (N_9780,N_9684,N_9685);
and U9781 (N_9781,N_9634,N_9745);
nor U9782 (N_9782,N_9622,N_9721);
or U9783 (N_9783,N_9635,N_9719);
xor U9784 (N_9784,N_9750,N_9672);
nor U9785 (N_9785,N_9626,N_9669);
or U9786 (N_9786,N_9673,N_9753);
or U9787 (N_9787,N_9604,N_9704);
nor U9788 (N_9788,N_9630,N_9679);
and U9789 (N_9789,N_9744,N_9600);
nor U9790 (N_9790,N_9688,N_9724);
xnor U9791 (N_9791,N_9658,N_9759);
or U9792 (N_9792,N_9722,N_9683);
or U9793 (N_9793,N_9706,N_9749);
xor U9794 (N_9794,N_9649,N_9659);
xor U9795 (N_9795,N_9715,N_9641);
nand U9796 (N_9796,N_9646,N_9740);
and U9797 (N_9797,N_9652,N_9707);
nand U9798 (N_9798,N_9726,N_9619);
xor U9799 (N_9799,N_9611,N_9665);
and U9800 (N_9800,N_9625,N_9667);
nor U9801 (N_9801,N_9666,N_9657);
or U9802 (N_9802,N_9651,N_9656);
xor U9803 (N_9803,N_9748,N_9705);
nand U9804 (N_9804,N_9644,N_9654);
or U9805 (N_9805,N_9709,N_9690);
nor U9806 (N_9806,N_9616,N_9633);
nand U9807 (N_9807,N_9756,N_9738);
nor U9808 (N_9808,N_9741,N_9734);
xor U9809 (N_9809,N_9711,N_9623);
nor U9810 (N_9810,N_9755,N_9661);
xnor U9811 (N_9811,N_9609,N_9643);
or U9812 (N_9812,N_9700,N_9746);
and U9813 (N_9813,N_9601,N_9743);
xnor U9814 (N_9814,N_9691,N_9697);
nand U9815 (N_9815,N_9725,N_9733);
xnor U9816 (N_9816,N_9698,N_9655);
nand U9817 (N_9817,N_9680,N_9710);
nor U9818 (N_9818,N_9677,N_9606);
and U9819 (N_9819,N_9612,N_9671);
xor U9820 (N_9820,N_9686,N_9742);
or U9821 (N_9821,N_9615,N_9678);
xor U9822 (N_9822,N_9613,N_9631);
xor U9823 (N_9823,N_9617,N_9729);
nand U9824 (N_9824,N_9681,N_9662);
or U9825 (N_9825,N_9676,N_9718);
or U9826 (N_9826,N_9605,N_9602);
and U9827 (N_9827,N_9716,N_9687);
nor U9828 (N_9828,N_9637,N_9692);
or U9829 (N_9829,N_9701,N_9638);
or U9830 (N_9830,N_9694,N_9757);
xnor U9831 (N_9831,N_9627,N_9713);
and U9832 (N_9832,N_9642,N_9689);
nor U9833 (N_9833,N_9614,N_9730);
nand U9834 (N_9834,N_9636,N_9702);
nand U9835 (N_9835,N_9660,N_9670);
or U9836 (N_9836,N_9650,N_9674);
or U9837 (N_9837,N_9629,N_9728);
nor U9838 (N_9838,N_9640,N_9732);
xor U9839 (N_9839,N_9620,N_9639);
nand U9840 (N_9840,N_9724,N_9610);
nor U9841 (N_9841,N_9650,N_9676);
nor U9842 (N_9842,N_9678,N_9700);
or U9843 (N_9843,N_9703,N_9668);
xnor U9844 (N_9844,N_9756,N_9603);
nand U9845 (N_9845,N_9608,N_9743);
nor U9846 (N_9846,N_9696,N_9609);
nand U9847 (N_9847,N_9679,N_9746);
nor U9848 (N_9848,N_9752,N_9719);
nand U9849 (N_9849,N_9752,N_9685);
nand U9850 (N_9850,N_9630,N_9651);
or U9851 (N_9851,N_9712,N_9618);
xnor U9852 (N_9852,N_9664,N_9708);
and U9853 (N_9853,N_9621,N_9692);
xor U9854 (N_9854,N_9635,N_9631);
and U9855 (N_9855,N_9687,N_9679);
and U9856 (N_9856,N_9652,N_9682);
nor U9857 (N_9857,N_9688,N_9655);
nand U9858 (N_9858,N_9705,N_9609);
or U9859 (N_9859,N_9671,N_9753);
nand U9860 (N_9860,N_9691,N_9616);
xnor U9861 (N_9861,N_9620,N_9699);
or U9862 (N_9862,N_9622,N_9713);
or U9863 (N_9863,N_9654,N_9683);
or U9864 (N_9864,N_9700,N_9653);
nand U9865 (N_9865,N_9679,N_9753);
or U9866 (N_9866,N_9654,N_9616);
nand U9867 (N_9867,N_9756,N_9651);
and U9868 (N_9868,N_9642,N_9670);
or U9869 (N_9869,N_9688,N_9646);
or U9870 (N_9870,N_9655,N_9676);
xnor U9871 (N_9871,N_9679,N_9635);
nand U9872 (N_9872,N_9665,N_9670);
or U9873 (N_9873,N_9671,N_9627);
nor U9874 (N_9874,N_9739,N_9614);
and U9875 (N_9875,N_9656,N_9731);
and U9876 (N_9876,N_9658,N_9612);
or U9877 (N_9877,N_9605,N_9724);
or U9878 (N_9878,N_9648,N_9667);
or U9879 (N_9879,N_9709,N_9732);
or U9880 (N_9880,N_9672,N_9654);
nand U9881 (N_9881,N_9673,N_9642);
nand U9882 (N_9882,N_9676,N_9661);
or U9883 (N_9883,N_9711,N_9652);
nor U9884 (N_9884,N_9707,N_9656);
xor U9885 (N_9885,N_9668,N_9614);
or U9886 (N_9886,N_9701,N_9743);
xor U9887 (N_9887,N_9617,N_9736);
nor U9888 (N_9888,N_9654,N_9755);
nor U9889 (N_9889,N_9690,N_9746);
or U9890 (N_9890,N_9602,N_9628);
nor U9891 (N_9891,N_9615,N_9608);
xnor U9892 (N_9892,N_9720,N_9695);
or U9893 (N_9893,N_9621,N_9634);
xor U9894 (N_9894,N_9701,N_9738);
nor U9895 (N_9895,N_9693,N_9612);
or U9896 (N_9896,N_9609,N_9662);
and U9897 (N_9897,N_9635,N_9684);
and U9898 (N_9898,N_9657,N_9686);
or U9899 (N_9899,N_9677,N_9716);
and U9900 (N_9900,N_9724,N_9614);
or U9901 (N_9901,N_9690,N_9609);
or U9902 (N_9902,N_9629,N_9643);
nor U9903 (N_9903,N_9733,N_9682);
xor U9904 (N_9904,N_9677,N_9647);
and U9905 (N_9905,N_9685,N_9739);
or U9906 (N_9906,N_9728,N_9751);
nor U9907 (N_9907,N_9615,N_9612);
nor U9908 (N_9908,N_9728,N_9680);
nand U9909 (N_9909,N_9656,N_9637);
xor U9910 (N_9910,N_9749,N_9614);
and U9911 (N_9911,N_9644,N_9631);
and U9912 (N_9912,N_9720,N_9640);
nor U9913 (N_9913,N_9742,N_9639);
nor U9914 (N_9914,N_9716,N_9668);
or U9915 (N_9915,N_9733,N_9643);
or U9916 (N_9916,N_9604,N_9728);
xnor U9917 (N_9917,N_9686,N_9606);
nor U9918 (N_9918,N_9678,N_9725);
or U9919 (N_9919,N_9645,N_9634);
nand U9920 (N_9920,N_9873,N_9888);
xor U9921 (N_9921,N_9781,N_9902);
xnor U9922 (N_9922,N_9765,N_9911);
nor U9923 (N_9923,N_9866,N_9838);
xor U9924 (N_9924,N_9876,N_9784);
and U9925 (N_9925,N_9889,N_9763);
nor U9926 (N_9926,N_9825,N_9832);
or U9927 (N_9927,N_9835,N_9792);
and U9928 (N_9928,N_9857,N_9865);
or U9929 (N_9929,N_9874,N_9836);
and U9930 (N_9930,N_9848,N_9789);
nor U9931 (N_9931,N_9912,N_9846);
nor U9932 (N_9932,N_9913,N_9831);
nand U9933 (N_9933,N_9783,N_9870);
xor U9934 (N_9934,N_9790,N_9868);
nand U9935 (N_9935,N_9890,N_9778);
xor U9936 (N_9936,N_9905,N_9794);
or U9937 (N_9937,N_9806,N_9909);
and U9938 (N_9938,N_9906,N_9884);
and U9939 (N_9939,N_9849,N_9775);
nand U9940 (N_9940,N_9845,N_9771);
and U9941 (N_9941,N_9894,N_9880);
or U9942 (N_9942,N_9760,N_9847);
nand U9943 (N_9943,N_9841,N_9893);
nor U9944 (N_9944,N_9915,N_9795);
nand U9945 (N_9945,N_9780,N_9769);
xor U9946 (N_9946,N_9916,N_9816);
xor U9947 (N_9947,N_9834,N_9858);
nor U9948 (N_9948,N_9774,N_9814);
nor U9949 (N_9949,N_9811,N_9854);
xor U9950 (N_9950,N_9833,N_9918);
nor U9951 (N_9951,N_9859,N_9910);
nor U9952 (N_9952,N_9869,N_9785);
nand U9953 (N_9953,N_9813,N_9875);
xor U9954 (N_9954,N_9844,N_9850);
and U9955 (N_9955,N_9819,N_9864);
and U9956 (N_9956,N_9881,N_9878);
or U9957 (N_9957,N_9882,N_9860);
xor U9958 (N_9958,N_9914,N_9762);
nand U9959 (N_9959,N_9862,N_9787);
nand U9960 (N_9960,N_9853,N_9899);
nor U9961 (N_9961,N_9786,N_9823);
nand U9962 (N_9962,N_9827,N_9871);
xor U9963 (N_9963,N_9805,N_9828);
nor U9964 (N_9964,N_9830,N_9826);
or U9965 (N_9965,N_9804,N_9779);
or U9966 (N_9966,N_9896,N_9761);
nor U9967 (N_9967,N_9852,N_9837);
and U9968 (N_9968,N_9788,N_9821);
nand U9969 (N_9969,N_9901,N_9883);
and U9970 (N_9970,N_9798,N_9812);
nor U9971 (N_9971,N_9840,N_9815);
nand U9972 (N_9972,N_9917,N_9839);
nor U9973 (N_9973,N_9809,N_9892);
nand U9974 (N_9974,N_9908,N_9810);
and U9975 (N_9975,N_9898,N_9800);
nand U9976 (N_9976,N_9768,N_9886);
or U9977 (N_9977,N_9863,N_9773);
nand U9978 (N_9978,N_9818,N_9801);
or U9979 (N_9979,N_9776,N_9900);
or U9980 (N_9980,N_9766,N_9843);
nor U9981 (N_9981,N_9887,N_9777);
xor U9982 (N_9982,N_9904,N_9807);
nor U9983 (N_9983,N_9764,N_9802);
and U9984 (N_9984,N_9856,N_9772);
and U9985 (N_9985,N_9797,N_9803);
or U9986 (N_9986,N_9879,N_9907);
nor U9987 (N_9987,N_9919,N_9770);
and U9988 (N_9988,N_9796,N_9822);
xor U9989 (N_9989,N_9897,N_9820);
xnor U9990 (N_9990,N_9895,N_9842);
nor U9991 (N_9991,N_9817,N_9855);
nand U9992 (N_9992,N_9791,N_9799);
or U9993 (N_9993,N_9885,N_9782);
nand U9994 (N_9994,N_9793,N_9872);
and U9995 (N_9995,N_9808,N_9829);
and U9996 (N_9996,N_9867,N_9824);
and U9997 (N_9997,N_9767,N_9903);
xor U9998 (N_9998,N_9891,N_9877);
xor U9999 (N_9999,N_9851,N_9861);
and U10000 (N_10000,N_9770,N_9870);
or U10001 (N_10001,N_9805,N_9822);
and U10002 (N_10002,N_9828,N_9813);
and U10003 (N_10003,N_9837,N_9870);
and U10004 (N_10004,N_9901,N_9897);
and U10005 (N_10005,N_9777,N_9907);
nor U10006 (N_10006,N_9872,N_9791);
and U10007 (N_10007,N_9906,N_9843);
xnor U10008 (N_10008,N_9900,N_9772);
nand U10009 (N_10009,N_9837,N_9838);
and U10010 (N_10010,N_9833,N_9825);
nor U10011 (N_10011,N_9865,N_9813);
xor U10012 (N_10012,N_9853,N_9791);
nor U10013 (N_10013,N_9772,N_9847);
nand U10014 (N_10014,N_9875,N_9855);
xnor U10015 (N_10015,N_9915,N_9881);
and U10016 (N_10016,N_9906,N_9832);
nand U10017 (N_10017,N_9788,N_9839);
nor U10018 (N_10018,N_9781,N_9855);
or U10019 (N_10019,N_9909,N_9850);
nand U10020 (N_10020,N_9838,N_9909);
and U10021 (N_10021,N_9881,N_9887);
nor U10022 (N_10022,N_9873,N_9806);
xnor U10023 (N_10023,N_9789,N_9884);
xnor U10024 (N_10024,N_9844,N_9841);
nand U10025 (N_10025,N_9837,N_9909);
xnor U10026 (N_10026,N_9901,N_9884);
xor U10027 (N_10027,N_9805,N_9776);
nand U10028 (N_10028,N_9873,N_9908);
xor U10029 (N_10029,N_9788,N_9792);
nand U10030 (N_10030,N_9871,N_9838);
nor U10031 (N_10031,N_9817,N_9878);
xor U10032 (N_10032,N_9841,N_9826);
and U10033 (N_10033,N_9915,N_9818);
nor U10034 (N_10034,N_9842,N_9846);
nand U10035 (N_10035,N_9788,N_9812);
nand U10036 (N_10036,N_9810,N_9769);
xnor U10037 (N_10037,N_9853,N_9862);
or U10038 (N_10038,N_9915,N_9883);
and U10039 (N_10039,N_9840,N_9810);
nor U10040 (N_10040,N_9824,N_9901);
nor U10041 (N_10041,N_9790,N_9910);
nor U10042 (N_10042,N_9845,N_9860);
and U10043 (N_10043,N_9763,N_9907);
nand U10044 (N_10044,N_9777,N_9779);
xor U10045 (N_10045,N_9886,N_9840);
xnor U10046 (N_10046,N_9762,N_9887);
nand U10047 (N_10047,N_9760,N_9826);
xor U10048 (N_10048,N_9772,N_9812);
or U10049 (N_10049,N_9862,N_9912);
nor U10050 (N_10050,N_9908,N_9814);
nor U10051 (N_10051,N_9880,N_9829);
nand U10052 (N_10052,N_9821,N_9893);
or U10053 (N_10053,N_9772,N_9859);
or U10054 (N_10054,N_9817,N_9904);
and U10055 (N_10055,N_9912,N_9906);
or U10056 (N_10056,N_9780,N_9809);
and U10057 (N_10057,N_9919,N_9820);
or U10058 (N_10058,N_9868,N_9847);
nand U10059 (N_10059,N_9836,N_9802);
nor U10060 (N_10060,N_9843,N_9789);
nand U10061 (N_10061,N_9875,N_9826);
and U10062 (N_10062,N_9840,N_9820);
and U10063 (N_10063,N_9806,N_9849);
xnor U10064 (N_10064,N_9839,N_9915);
nand U10065 (N_10065,N_9828,N_9902);
nand U10066 (N_10066,N_9837,N_9896);
xor U10067 (N_10067,N_9793,N_9760);
nor U10068 (N_10068,N_9812,N_9776);
xnor U10069 (N_10069,N_9902,N_9865);
xnor U10070 (N_10070,N_9777,N_9867);
xnor U10071 (N_10071,N_9884,N_9856);
nand U10072 (N_10072,N_9872,N_9902);
and U10073 (N_10073,N_9895,N_9811);
nand U10074 (N_10074,N_9844,N_9775);
and U10075 (N_10075,N_9871,N_9842);
nor U10076 (N_10076,N_9902,N_9859);
xnor U10077 (N_10077,N_9890,N_9769);
or U10078 (N_10078,N_9904,N_9760);
nand U10079 (N_10079,N_9912,N_9899);
and U10080 (N_10080,N_10052,N_10004);
or U10081 (N_10081,N_9995,N_10067);
and U10082 (N_10082,N_10061,N_9974);
or U10083 (N_10083,N_10054,N_10068);
and U10084 (N_10084,N_10000,N_9931);
and U10085 (N_10085,N_10040,N_9994);
nor U10086 (N_10086,N_10045,N_10005);
and U10087 (N_10087,N_9958,N_9956);
and U10088 (N_10088,N_10053,N_9941);
xnor U10089 (N_10089,N_10066,N_10014);
and U10090 (N_10090,N_10036,N_10006);
or U10091 (N_10091,N_10035,N_9942);
nor U10092 (N_10092,N_9935,N_10022);
xor U10093 (N_10093,N_9945,N_10059);
or U10094 (N_10094,N_9993,N_10037);
or U10095 (N_10095,N_9949,N_10019);
or U10096 (N_10096,N_9999,N_9985);
nand U10097 (N_10097,N_9982,N_9988);
nand U10098 (N_10098,N_9973,N_9966);
and U10099 (N_10099,N_10016,N_10033);
xnor U10100 (N_10100,N_10008,N_10015);
and U10101 (N_10101,N_9965,N_10058);
nand U10102 (N_10102,N_10055,N_9959);
or U10103 (N_10103,N_10027,N_10047);
nand U10104 (N_10104,N_9975,N_10034);
nor U10105 (N_10105,N_9921,N_10060);
xnor U10106 (N_10106,N_9926,N_10042);
nand U10107 (N_10107,N_9950,N_10023);
nor U10108 (N_10108,N_10077,N_9951);
and U10109 (N_10109,N_10043,N_10071);
xnor U10110 (N_10110,N_9987,N_10039);
xnor U10111 (N_10111,N_9940,N_10076);
nor U10112 (N_10112,N_9944,N_9990);
nor U10113 (N_10113,N_10046,N_10018);
or U10114 (N_10114,N_9943,N_9963);
nand U10115 (N_10115,N_9969,N_10007);
or U10116 (N_10116,N_10057,N_9954);
xnor U10117 (N_10117,N_9947,N_9962);
and U10118 (N_10118,N_9928,N_10002);
xor U10119 (N_10119,N_9961,N_10011);
nand U10120 (N_10120,N_9983,N_9968);
nor U10121 (N_10121,N_10024,N_9992);
xor U10122 (N_10122,N_9934,N_10074);
or U10123 (N_10123,N_10017,N_9979);
and U10124 (N_10124,N_10041,N_10070);
nor U10125 (N_10125,N_10032,N_10078);
nand U10126 (N_10126,N_9989,N_9977);
nand U10127 (N_10127,N_9924,N_10013);
xor U10128 (N_10128,N_10003,N_10056);
and U10129 (N_10129,N_10064,N_9957);
nand U10130 (N_10130,N_10029,N_9922);
and U10131 (N_10131,N_10051,N_9981);
and U10132 (N_10132,N_10079,N_9964);
nand U10133 (N_10133,N_9976,N_9998);
xnor U10134 (N_10134,N_10069,N_9923);
xnor U10135 (N_10135,N_9920,N_10020);
and U10136 (N_10136,N_9978,N_9996);
xnor U10137 (N_10137,N_9927,N_9991);
xnor U10138 (N_10138,N_9955,N_9932);
or U10139 (N_10139,N_10001,N_10073);
xor U10140 (N_10140,N_9952,N_10026);
nor U10141 (N_10141,N_10048,N_10031);
or U10142 (N_10142,N_9971,N_9997);
or U10143 (N_10143,N_9936,N_9948);
and U10144 (N_10144,N_10028,N_9967);
nor U10145 (N_10145,N_10012,N_9933);
or U10146 (N_10146,N_10025,N_10062);
and U10147 (N_10147,N_10050,N_10038);
or U10148 (N_10148,N_9937,N_10049);
or U10149 (N_10149,N_9925,N_9986);
nor U10150 (N_10150,N_10021,N_9929);
nand U10151 (N_10151,N_9938,N_9953);
nand U10152 (N_10152,N_10065,N_9984);
nor U10153 (N_10153,N_9970,N_10010);
and U10154 (N_10154,N_9980,N_10030);
xor U10155 (N_10155,N_10009,N_9930);
xnor U10156 (N_10156,N_10063,N_9939);
nand U10157 (N_10157,N_10075,N_10044);
xnor U10158 (N_10158,N_9972,N_9946);
or U10159 (N_10159,N_10072,N_9960);
nand U10160 (N_10160,N_9962,N_9971);
xnor U10161 (N_10161,N_9948,N_9966);
xor U10162 (N_10162,N_10056,N_10057);
nand U10163 (N_10163,N_9998,N_10053);
nand U10164 (N_10164,N_10072,N_9947);
nand U10165 (N_10165,N_9997,N_9941);
xor U10166 (N_10166,N_10078,N_9958);
nor U10167 (N_10167,N_9998,N_10035);
nand U10168 (N_10168,N_10003,N_9972);
nand U10169 (N_10169,N_10008,N_9954);
and U10170 (N_10170,N_10056,N_9941);
and U10171 (N_10171,N_10004,N_10074);
nand U10172 (N_10172,N_10042,N_10057);
nor U10173 (N_10173,N_9982,N_10065);
xnor U10174 (N_10174,N_10078,N_9936);
nand U10175 (N_10175,N_9978,N_10021);
nand U10176 (N_10176,N_9952,N_10032);
and U10177 (N_10177,N_10011,N_10007);
xor U10178 (N_10178,N_9938,N_9990);
and U10179 (N_10179,N_10032,N_9959);
xnor U10180 (N_10180,N_9941,N_9964);
xnor U10181 (N_10181,N_10025,N_9994);
and U10182 (N_10182,N_10035,N_9970);
nand U10183 (N_10183,N_9982,N_10031);
or U10184 (N_10184,N_9939,N_10013);
xor U10185 (N_10185,N_10077,N_10079);
xnor U10186 (N_10186,N_9997,N_10024);
or U10187 (N_10187,N_9972,N_10078);
and U10188 (N_10188,N_9976,N_9980);
and U10189 (N_10189,N_10045,N_10010);
nor U10190 (N_10190,N_9950,N_10073);
or U10191 (N_10191,N_9927,N_9952);
xnor U10192 (N_10192,N_9942,N_10028);
and U10193 (N_10193,N_10068,N_10062);
and U10194 (N_10194,N_10016,N_10013);
or U10195 (N_10195,N_9961,N_10073);
nor U10196 (N_10196,N_10012,N_10070);
xor U10197 (N_10197,N_9957,N_9993);
and U10198 (N_10198,N_9925,N_10042);
or U10199 (N_10199,N_9934,N_9926);
nor U10200 (N_10200,N_9932,N_9969);
nand U10201 (N_10201,N_10023,N_10072);
nand U10202 (N_10202,N_9999,N_10056);
nor U10203 (N_10203,N_10058,N_10041);
nand U10204 (N_10204,N_9968,N_9972);
nand U10205 (N_10205,N_9990,N_9921);
and U10206 (N_10206,N_9963,N_10062);
nand U10207 (N_10207,N_10010,N_10013);
or U10208 (N_10208,N_10061,N_9952);
xor U10209 (N_10209,N_9941,N_10015);
nor U10210 (N_10210,N_10010,N_10079);
nand U10211 (N_10211,N_10013,N_9971);
or U10212 (N_10212,N_9959,N_9999);
nor U10213 (N_10213,N_10009,N_9959);
nor U10214 (N_10214,N_10076,N_9975);
and U10215 (N_10215,N_9943,N_9983);
nand U10216 (N_10216,N_9992,N_10036);
or U10217 (N_10217,N_10004,N_10028);
or U10218 (N_10218,N_9926,N_9924);
and U10219 (N_10219,N_9948,N_9967);
and U10220 (N_10220,N_9996,N_9979);
and U10221 (N_10221,N_9988,N_10020);
and U10222 (N_10222,N_9995,N_9954);
or U10223 (N_10223,N_9973,N_10052);
nand U10224 (N_10224,N_10025,N_9969);
nand U10225 (N_10225,N_9941,N_10058);
xor U10226 (N_10226,N_10066,N_9974);
nand U10227 (N_10227,N_9953,N_10001);
nor U10228 (N_10228,N_10008,N_10038);
or U10229 (N_10229,N_10020,N_9986);
nor U10230 (N_10230,N_10001,N_10008);
and U10231 (N_10231,N_10043,N_10068);
or U10232 (N_10232,N_9987,N_9920);
nor U10233 (N_10233,N_10075,N_9993);
or U10234 (N_10234,N_10045,N_10003);
nand U10235 (N_10235,N_9952,N_10017);
nor U10236 (N_10236,N_9920,N_9947);
nand U10237 (N_10237,N_10078,N_10076);
or U10238 (N_10238,N_9920,N_10016);
or U10239 (N_10239,N_9929,N_10011);
xor U10240 (N_10240,N_10114,N_10175);
nand U10241 (N_10241,N_10229,N_10107);
or U10242 (N_10242,N_10196,N_10156);
or U10243 (N_10243,N_10168,N_10176);
and U10244 (N_10244,N_10150,N_10223);
nand U10245 (N_10245,N_10096,N_10113);
nand U10246 (N_10246,N_10082,N_10202);
nor U10247 (N_10247,N_10190,N_10139);
nand U10248 (N_10248,N_10101,N_10085);
nand U10249 (N_10249,N_10219,N_10203);
and U10250 (N_10250,N_10171,N_10206);
or U10251 (N_10251,N_10126,N_10216);
nor U10252 (N_10252,N_10160,N_10142);
xor U10253 (N_10253,N_10111,N_10132);
xor U10254 (N_10254,N_10125,N_10090);
xnor U10255 (N_10255,N_10129,N_10182);
nand U10256 (N_10256,N_10163,N_10173);
nor U10257 (N_10257,N_10106,N_10094);
and U10258 (N_10258,N_10121,N_10097);
or U10259 (N_10259,N_10110,N_10108);
nand U10260 (N_10260,N_10158,N_10170);
and U10261 (N_10261,N_10169,N_10239);
and U10262 (N_10262,N_10215,N_10145);
xor U10263 (N_10263,N_10135,N_10212);
nand U10264 (N_10264,N_10102,N_10207);
or U10265 (N_10265,N_10232,N_10086);
nor U10266 (N_10266,N_10172,N_10091);
nor U10267 (N_10267,N_10220,N_10116);
nand U10268 (N_10268,N_10187,N_10205);
or U10269 (N_10269,N_10217,N_10133);
nand U10270 (N_10270,N_10164,N_10230);
nand U10271 (N_10271,N_10128,N_10138);
xnor U10272 (N_10272,N_10087,N_10181);
xor U10273 (N_10273,N_10123,N_10161);
xor U10274 (N_10274,N_10191,N_10180);
nand U10275 (N_10275,N_10198,N_10152);
xor U10276 (N_10276,N_10165,N_10208);
xnor U10277 (N_10277,N_10186,N_10100);
nand U10278 (N_10278,N_10146,N_10231);
and U10279 (N_10279,N_10224,N_10083);
or U10280 (N_10280,N_10183,N_10235);
xor U10281 (N_10281,N_10127,N_10140);
or U10282 (N_10282,N_10131,N_10117);
and U10283 (N_10283,N_10234,N_10195);
nand U10284 (N_10284,N_10098,N_10227);
nor U10285 (N_10285,N_10159,N_10174);
and U10286 (N_10286,N_10179,N_10192);
nor U10287 (N_10287,N_10103,N_10136);
nand U10288 (N_10288,N_10194,N_10120);
and U10289 (N_10289,N_10222,N_10201);
and U10290 (N_10290,N_10193,N_10148);
and U10291 (N_10291,N_10084,N_10233);
and U10292 (N_10292,N_10112,N_10099);
nand U10293 (N_10293,N_10167,N_10213);
xor U10294 (N_10294,N_10185,N_10119);
nand U10295 (N_10295,N_10162,N_10221);
or U10296 (N_10296,N_10144,N_10109);
xor U10297 (N_10297,N_10093,N_10088);
xor U10298 (N_10298,N_10189,N_10130);
and U10299 (N_10299,N_10095,N_10238);
nand U10300 (N_10300,N_10092,N_10143);
and U10301 (N_10301,N_10134,N_10105);
nand U10302 (N_10302,N_10155,N_10226);
xnor U10303 (N_10303,N_10154,N_10153);
nor U10304 (N_10304,N_10177,N_10214);
nor U10305 (N_10305,N_10157,N_10200);
or U10306 (N_10306,N_10184,N_10237);
or U10307 (N_10307,N_10218,N_10204);
or U10308 (N_10308,N_10080,N_10149);
or U10309 (N_10309,N_10228,N_10225);
and U10310 (N_10310,N_10137,N_10104);
xnor U10311 (N_10311,N_10188,N_10122);
or U10312 (N_10312,N_10147,N_10209);
nor U10313 (N_10313,N_10089,N_10178);
or U10314 (N_10314,N_10210,N_10197);
nor U10315 (N_10315,N_10124,N_10211);
or U10316 (N_10316,N_10141,N_10236);
nand U10317 (N_10317,N_10151,N_10081);
xor U10318 (N_10318,N_10166,N_10199);
nand U10319 (N_10319,N_10118,N_10115);
nor U10320 (N_10320,N_10129,N_10179);
nand U10321 (N_10321,N_10188,N_10133);
or U10322 (N_10322,N_10083,N_10173);
nor U10323 (N_10323,N_10221,N_10136);
nor U10324 (N_10324,N_10224,N_10191);
or U10325 (N_10325,N_10205,N_10122);
xnor U10326 (N_10326,N_10229,N_10219);
xnor U10327 (N_10327,N_10147,N_10237);
nand U10328 (N_10328,N_10235,N_10093);
xor U10329 (N_10329,N_10172,N_10109);
nand U10330 (N_10330,N_10147,N_10150);
and U10331 (N_10331,N_10194,N_10207);
nand U10332 (N_10332,N_10083,N_10129);
nor U10333 (N_10333,N_10136,N_10106);
nor U10334 (N_10334,N_10213,N_10087);
xnor U10335 (N_10335,N_10213,N_10154);
or U10336 (N_10336,N_10203,N_10118);
nor U10337 (N_10337,N_10202,N_10195);
or U10338 (N_10338,N_10215,N_10119);
nand U10339 (N_10339,N_10225,N_10172);
nor U10340 (N_10340,N_10086,N_10172);
and U10341 (N_10341,N_10102,N_10205);
and U10342 (N_10342,N_10180,N_10212);
or U10343 (N_10343,N_10158,N_10235);
xnor U10344 (N_10344,N_10170,N_10234);
nor U10345 (N_10345,N_10210,N_10090);
nand U10346 (N_10346,N_10147,N_10127);
xnor U10347 (N_10347,N_10174,N_10111);
xnor U10348 (N_10348,N_10093,N_10128);
or U10349 (N_10349,N_10133,N_10239);
xnor U10350 (N_10350,N_10122,N_10080);
nand U10351 (N_10351,N_10118,N_10108);
xnor U10352 (N_10352,N_10172,N_10099);
nand U10353 (N_10353,N_10238,N_10179);
or U10354 (N_10354,N_10119,N_10083);
and U10355 (N_10355,N_10192,N_10096);
and U10356 (N_10356,N_10170,N_10106);
xor U10357 (N_10357,N_10105,N_10153);
nand U10358 (N_10358,N_10148,N_10171);
or U10359 (N_10359,N_10142,N_10201);
and U10360 (N_10360,N_10114,N_10220);
xnor U10361 (N_10361,N_10162,N_10236);
or U10362 (N_10362,N_10175,N_10117);
xnor U10363 (N_10363,N_10189,N_10175);
nand U10364 (N_10364,N_10227,N_10161);
or U10365 (N_10365,N_10146,N_10223);
and U10366 (N_10366,N_10147,N_10119);
nand U10367 (N_10367,N_10137,N_10156);
nand U10368 (N_10368,N_10132,N_10237);
xnor U10369 (N_10369,N_10100,N_10162);
or U10370 (N_10370,N_10091,N_10227);
and U10371 (N_10371,N_10082,N_10081);
nor U10372 (N_10372,N_10161,N_10174);
nand U10373 (N_10373,N_10089,N_10191);
and U10374 (N_10374,N_10222,N_10115);
or U10375 (N_10375,N_10134,N_10081);
nand U10376 (N_10376,N_10131,N_10120);
or U10377 (N_10377,N_10112,N_10101);
nor U10378 (N_10378,N_10234,N_10106);
or U10379 (N_10379,N_10222,N_10153);
or U10380 (N_10380,N_10218,N_10109);
xnor U10381 (N_10381,N_10193,N_10081);
nand U10382 (N_10382,N_10151,N_10239);
nand U10383 (N_10383,N_10236,N_10173);
and U10384 (N_10384,N_10125,N_10212);
nand U10385 (N_10385,N_10091,N_10235);
or U10386 (N_10386,N_10084,N_10177);
xor U10387 (N_10387,N_10137,N_10158);
nor U10388 (N_10388,N_10230,N_10235);
nand U10389 (N_10389,N_10080,N_10168);
nor U10390 (N_10390,N_10126,N_10158);
xor U10391 (N_10391,N_10119,N_10224);
nand U10392 (N_10392,N_10141,N_10158);
nand U10393 (N_10393,N_10088,N_10185);
nor U10394 (N_10394,N_10089,N_10083);
xor U10395 (N_10395,N_10211,N_10123);
nand U10396 (N_10396,N_10224,N_10147);
and U10397 (N_10397,N_10088,N_10203);
and U10398 (N_10398,N_10163,N_10126);
xnor U10399 (N_10399,N_10116,N_10189);
and U10400 (N_10400,N_10346,N_10297);
xor U10401 (N_10401,N_10271,N_10397);
or U10402 (N_10402,N_10329,N_10347);
and U10403 (N_10403,N_10258,N_10368);
or U10404 (N_10404,N_10316,N_10356);
or U10405 (N_10405,N_10375,N_10332);
and U10406 (N_10406,N_10282,N_10250);
nand U10407 (N_10407,N_10277,N_10374);
xor U10408 (N_10408,N_10262,N_10280);
and U10409 (N_10409,N_10377,N_10362);
or U10410 (N_10410,N_10321,N_10295);
nand U10411 (N_10411,N_10313,N_10359);
xor U10412 (N_10412,N_10357,N_10275);
and U10413 (N_10413,N_10340,N_10394);
xnor U10414 (N_10414,N_10281,N_10351);
nand U10415 (N_10415,N_10353,N_10274);
nor U10416 (N_10416,N_10283,N_10391);
nand U10417 (N_10417,N_10370,N_10293);
nor U10418 (N_10418,N_10330,N_10276);
xnor U10419 (N_10419,N_10335,N_10298);
and U10420 (N_10420,N_10327,N_10311);
nand U10421 (N_10421,N_10251,N_10382);
and U10422 (N_10422,N_10317,N_10367);
or U10423 (N_10423,N_10256,N_10264);
xor U10424 (N_10424,N_10318,N_10396);
nor U10425 (N_10425,N_10319,N_10325);
and U10426 (N_10426,N_10369,N_10333);
and U10427 (N_10427,N_10380,N_10389);
nor U10428 (N_10428,N_10244,N_10289);
nand U10429 (N_10429,N_10399,N_10290);
xor U10430 (N_10430,N_10272,N_10286);
xnor U10431 (N_10431,N_10247,N_10383);
nor U10432 (N_10432,N_10331,N_10296);
nor U10433 (N_10433,N_10301,N_10269);
and U10434 (N_10434,N_10305,N_10336);
and U10435 (N_10435,N_10285,N_10348);
xor U10436 (N_10436,N_10373,N_10334);
nor U10437 (N_10437,N_10254,N_10393);
or U10438 (N_10438,N_10288,N_10379);
nor U10439 (N_10439,N_10342,N_10339);
xnor U10440 (N_10440,N_10243,N_10246);
nand U10441 (N_10441,N_10384,N_10259);
nand U10442 (N_10442,N_10261,N_10260);
nand U10443 (N_10443,N_10381,N_10345);
or U10444 (N_10444,N_10303,N_10365);
xnor U10445 (N_10445,N_10278,N_10364);
and U10446 (N_10446,N_10372,N_10360);
nor U10447 (N_10447,N_10291,N_10248);
and U10448 (N_10448,N_10371,N_10268);
nand U10449 (N_10449,N_10299,N_10320);
nor U10450 (N_10450,N_10265,N_10287);
or U10451 (N_10451,N_10245,N_10349);
and U10452 (N_10452,N_10249,N_10302);
xnor U10453 (N_10453,N_10252,N_10322);
or U10454 (N_10454,N_10257,N_10354);
or U10455 (N_10455,N_10338,N_10324);
and U10456 (N_10456,N_10241,N_10314);
or U10457 (N_10457,N_10310,N_10385);
xnor U10458 (N_10458,N_10294,N_10366);
and U10459 (N_10459,N_10387,N_10284);
xnor U10460 (N_10460,N_10266,N_10323);
and U10461 (N_10461,N_10392,N_10304);
or U10462 (N_10462,N_10263,N_10328);
or U10463 (N_10463,N_10388,N_10270);
and U10464 (N_10464,N_10361,N_10378);
xnor U10465 (N_10465,N_10343,N_10341);
or U10466 (N_10466,N_10255,N_10352);
and U10467 (N_10467,N_10386,N_10337);
nor U10468 (N_10468,N_10309,N_10308);
and U10469 (N_10469,N_10315,N_10306);
xnor U10470 (N_10470,N_10376,N_10395);
nor U10471 (N_10471,N_10292,N_10355);
nor U10472 (N_10472,N_10350,N_10326);
or U10473 (N_10473,N_10267,N_10240);
nand U10474 (N_10474,N_10273,N_10390);
and U10475 (N_10475,N_10279,N_10300);
nand U10476 (N_10476,N_10358,N_10307);
or U10477 (N_10477,N_10242,N_10363);
or U10478 (N_10478,N_10312,N_10344);
or U10479 (N_10479,N_10253,N_10398);
xnor U10480 (N_10480,N_10295,N_10277);
nor U10481 (N_10481,N_10367,N_10307);
or U10482 (N_10482,N_10260,N_10240);
or U10483 (N_10483,N_10330,N_10381);
and U10484 (N_10484,N_10324,N_10254);
nand U10485 (N_10485,N_10248,N_10254);
nor U10486 (N_10486,N_10323,N_10256);
nor U10487 (N_10487,N_10359,N_10327);
nor U10488 (N_10488,N_10360,N_10383);
xnor U10489 (N_10489,N_10346,N_10342);
or U10490 (N_10490,N_10315,N_10293);
nand U10491 (N_10491,N_10288,N_10310);
xnor U10492 (N_10492,N_10298,N_10381);
xnor U10493 (N_10493,N_10278,N_10267);
nand U10494 (N_10494,N_10295,N_10269);
nor U10495 (N_10495,N_10292,N_10273);
nor U10496 (N_10496,N_10278,N_10380);
and U10497 (N_10497,N_10361,N_10240);
or U10498 (N_10498,N_10313,N_10342);
or U10499 (N_10499,N_10264,N_10310);
and U10500 (N_10500,N_10291,N_10345);
xnor U10501 (N_10501,N_10248,N_10326);
nor U10502 (N_10502,N_10383,N_10384);
xnor U10503 (N_10503,N_10345,N_10273);
xor U10504 (N_10504,N_10313,N_10257);
nand U10505 (N_10505,N_10288,N_10344);
or U10506 (N_10506,N_10259,N_10306);
nor U10507 (N_10507,N_10380,N_10255);
and U10508 (N_10508,N_10271,N_10247);
and U10509 (N_10509,N_10375,N_10248);
and U10510 (N_10510,N_10294,N_10271);
or U10511 (N_10511,N_10312,N_10242);
or U10512 (N_10512,N_10281,N_10271);
nor U10513 (N_10513,N_10319,N_10290);
nor U10514 (N_10514,N_10329,N_10266);
or U10515 (N_10515,N_10392,N_10288);
nand U10516 (N_10516,N_10306,N_10333);
nand U10517 (N_10517,N_10257,N_10314);
nor U10518 (N_10518,N_10336,N_10301);
xnor U10519 (N_10519,N_10358,N_10394);
nand U10520 (N_10520,N_10395,N_10389);
nor U10521 (N_10521,N_10262,N_10265);
xor U10522 (N_10522,N_10385,N_10324);
xnor U10523 (N_10523,N_10305,N_10369);
nand U10524 (N_10524,N_10348,N_10329);
nor U10525 (N_10525,N_10280,N_10379);
and U10526 (N_10526,N_10384,N_10241);
nor U10527 (N_10527,N_10249,N_10309);
and U10528 (N_10528,N_10296,N_10245);
nand U10529 (N_10529,N_10252,N_10350);
nand U10530 (N_10530,N_10260,N_10274);
nor U10531 (N_10531,N_10331,N_10266);
xnor U10532 (N_10532,N_10272,N_10378);
xnor U10533 (N_10533,N_10248,N_10388);
xor U10534 (N_10534,N_10306,N_10349);
and U10535 (N_10535,N_10375,N_10349);
nand U10536 (N_10536,N_10271,N_10343);
nor U10537 (N_10537,N_10241,N_10332);
xnor U10538 (N_10538,N_10247,N_10292);
xnor U10539 (N_10539,N_10332,N_10250);
nand U10540 (N_10540,N_10353,N_10344);
or U10541 (N_10541,N_10367,N_10247);
xnor U10542 (N_10542,N_10298,N_10325);
nor U10543 (N_10543,N_10383,N_10394);
nand U10544 (N_10544,N_10312,N_10396);
xnor U10545 (N_10545,N_10252,N_10396);
xor U10546 (N_10546,N_10288,N_10342);
nand U10547 (N_10547,N_10388,N_10292);
nand U10548 (N_10548,N_10334,N_10357);
and U10549 (N_10549,N_10373,N_10379);
and U10550 (N_10550,N_10374,N_10278);
and U10551 (N_10551,N_10309,N_10334);
xor U10552 (N_10552,N_10325,N_10288);
or U10553 (N_10553,N_10262,N_10333);
nand U10554 (N_10554,N_10373,N_10283);
nand U10555 (N_10555,N_10302,N_10248);
nor U10556 (N_10556,N_10300,N_10398);
nor U10557 (N_10557,N_10381,N_10354);
nor U10558 (N_10558,N_10334,N_10312);
xnor U10559 (N_10559,N_10393,N_10316);
nand U10560 (N_10560,N_10526,N_10530);
xnor U10561 (N_10561,N_10401,N_10549);
xor U10562 (N_10562,N_10551,N_10519);
xor U10563 (N_10563,N_10436,N_10463);
and U10564 (N_10564,N_10419,N_10439);
xor U10565 (N_10565,N_10480,N_10426);
xnor U10566 (N_10566,N_10534,N_10459);
and U10567 (N_10567,N_10457,N_10450);
nand U10568 (N_10568,N_10402,N_10531);
xor U10569 (N_10569,N_10427,N_10453);
xor U10570 (N_10570,N_10500,N_10489);
nand U10571 (N_10571,N_10403,N_10458);
or U10572 (N_10572,N_10490,N_10416);
xnor U10573 (N_10573,N_10466,N_10470);
and U10574 (N_10574,N_10412,N_10456);
or U10575 (N_10575,N_10522,N_10468);
xor U10576 (N_10576,N_10516,N_10409);
nand U10577 (N_10577,N_10484,N_10407);
nor U10578 (N_10578,N_10438,N_10481);
nand U10579 (N_10579,N_10405,N_10454);
nand U10580 (N_10580,N_10503,N_10512);
nor U10581 (N_10581,N_10511,N_10462);
nor U10582 (N_10582,N_10492,N_10498);
nand U10583 (N_10583,N_10537,N_10477);
xnor U10584 (N_10584,N_10533,N_10421);
or U10585 (N_10585,N_10449,N_10528);
and U10586 (N_10586,N_10487,N_10485);
or U10587 (N_10587,N_10418,N_10495);
or U10588 (N_10588,N_10432,N_10555);
and U10589 (N_10589,N_10536,N_10502);
and U10590 (N_10590,N_10504,N_10451);
nand U10591 (N_10591,N_10482,N_10417);
nand U10592 (N_10592,N_10505,N_10429);
xor U10593 (N_10593,N_10483,N_10400);
nor U10594 (N_10594,N_10446,N_10521);
or U10595 (N_10595,N_10541,N_10506);
or U10596 (N_10596,N_10424,N_10434);
or U10597 (N_10597,N_10471,N_10491);
and U10598 (N_10598,N_10479,N_10431);
and U10599 (N_10599,N_10444,N_10497);
or U10600 (N_10600,N_10540,N_10513);
and U10601 (N_10601,N_10488,N_10452);
or U10602 (N_10602,N_10556,N_10435);
xnor U10603 (N_10603,N_10411,N_10441);
nand U10604 (N_10604,N_10535,N_10496);
nor U10605 (N_10605,N_10554,N_10428);
and U10606 (N_10606,N_10553,N_10425);
nand U10607 (N_10607,N_10547,N_10532);
nor U10608 (N_10608,N_10406,N_10447);
nand U10609 (N_10609,N_10475,N_10465);
nor U10610 (N_10610,N_10461,N_10442);
and U10611 (N_10611,N_10408,N_10548);
or U10612 (N_10612,N_10493,N_10507);
and U10613 (N_10613,N_10515,N_10415);
nand U10614 (N_10614,N_10520,N_10552);
and U10615 (N_10615,N_10542,N_10430);
nor U10616 (N_10616,N_10543,N_10440);
or U10617 (N_10617,N_10464,N_10437);
nand U10618 (N_10618,N_10539,N_10523);
or U10619 (N_10619,N_10509,N_10460);
nand U10620 (N_10620,N_10524,N_10474);
and U10621 (N_10621,N_10544,N_10510);
nor U10622 (N_10622,N_10545,N_10469);
nor U10623 (N_10623,N_10525,N_10448);
or U10624 (N_10624,N_10455,N_10494);
nand U10625 (N_10625,N_10558,N_10546);
or U10626 (N_10626,N_10527,N_10445);
nand U10627 (N_10627,N_10433,N_10473);
nor U10628 (N_10628,N_10413,N_10467);
nand U10629 (N_10629,N_10443,N_10559);
and U10630 (N_10630,N_10557,N_10404);
nor U10631 (N_10631,N_10410,N_10508);
and U10632 (N_10632,N_10472,N_10422);
xnor U10633 (N_10633,N_10420,N_10529);
or U10634 (N_10634,N_10550,N_10499);
xnor U10635 (N_10635,N_10517,N_10423);
and U10636 (N_10636,N_10476,N_10478);
and U10637 (N_10637,N_10518,N_10538);
xor U10638 (N_10638,N_10414,N_10501);
or U10639 (N_10639,N_10514,N_10486);
nand U10640 (N_10640,N_10445,N_10468);
xnor U10641 (N_10641,N_10414,N_10483);
nand U10642 (N_10642,N_10404,N_10521);
xor U10643 (N_10643,N_10511,N_10473);
nand U10644 (N_10644,N_10409,N_10534);
nand U10645 (N_10645,N_10484,N_10552);
xnor U10646 (N_10646,N_10436,N_10482);
xnor U10647 (N_10647,N_10441,N_10481);
xnor U10648 (N_10648,N_10518,N_10491);
and U10649 (N_10649,N_10411,N_10498);
or U10650 (N_10650,N_10446,N_10557);
or U10651 (N_10651,N_10512,N_10520);
or U10652 (N_10652,N_10501,N_10467);
xnor U10653 (N_10653,N_10516,N_10527);
nor U10654 (N_10654,N_10512,N_10404);
nor U10655 (N_10655,N_10525,N_10551);
or U10656 (N_10656,N_10535,N_10482);
and U10657 (N_10657,N_10544,N_10416);
nand U10658 (N_10658,N_10425,N_10461);
nor U10659 (N_10659,N_10461,N_10524);
or U10660 (N_10660,N_10516,N_10422);
and U10661 (N_10661,N_10507,N_10557);
and U10662 (N_10662,N_10533,N_10501);
nand U10663 (N_10663,N_10524,N_10498);
xor U10664 (N_10664,N_10439,N_10487);
and U10665 (N_10665,N_10428,N_10414);
nand U10666 (N_10666,N_10402,N_10510);
or U10667 (N_10667,N_10519,N_10494);
xor U10668 (N_10668,N_10490,N_10558);
nand U10669 (N_10669,N_10544,N_10554);
or U10670 (N_10670,N_10526,N_10483);
nor U10671 (N_10671,N_10539,N_10434);
xor U10672 (N_10672,N_10413,N_10469);
nor U10673 (N_10673,N_10495,N_10534);
nor U10674 (N_10674,N_10405,N_10538);
and U10675 (N_10675,N_10491,N_10489);
xor U10676 (N_10676,N_10550,N_10474);
nand U10677 (N_10677,N_10474,N_10467);
nor U10678 (N_10678,N_10545,N_10548);
nor U10679 (N_10679,N_10548,N_10529);
or U10680 (N_10680,N_10425,N_10435);
nor U10681 (N_10681,N_10547,N_10557);
xor U10682 (N_10682,N_10432,N_10431);
nor U10683 (N_10683,N_10516,N_10460);
nand U10684 (N_10684,N_10409,N_10507);
nor U10685 (N_10685,N_10542,N_10432);
nor U10686 (N_10686,N_10477,N_10446);
nand U10687 (N_10687,N_10527,N_10513);
nand U10688 (N_10688,N_10453,N_10500);
xor U10689 (N_10689,N_10487,N_10496);
xnor U10690 (N_10690,N_10461,N_10459);
and U10691 (N_10691,N_10542,N_10466);
nor U10692 (N_10692,N_10438,N_10440);
nand U10693 (N_10693,N_10404,N_10425);
nor U10694 (N_10694,N_10472,N_10530);
nand U10695 (N_10695,N_10472,N_10412);
xor U10696 (N_10696,N_10517,N_10421);
nand U10697 (N_10697,N_10421,N_10434);
nand U10698 (N_10698,N_10544,N_10530);
nor U10699 (N_10699,N_10473,N_10519);
or U10700 (N_10700,N_10475,N_10481);
and U10701 (N_10701,N_10512,N_10484);
nor U10702 (N_10702,N_10423,N_10525);
nand U10703 (N_10703,N_10417,N_10434);
nor U10704 (N_10704,N_10545,N_10462);
xor U10705 (N_10705,N_10460,N_10407);
or U10706 (N_10706,N_10535,N_10532);
xnor U10707 (N_10707,N_10508,N_10481);
nand U10708 (N_10708,N_10449,N_10508);
and U10709 (N_10709,N_10542,N_10406);
nor U10710 (N_10710,N_10438,N_10420);
xnor U10711 (N_10711,N_10529,N_10500);
xnor U10712 (N_10712,N_10517,N_10451);
and U10713 (N_10713,N_10520,N_10557);
xor U10714 (N_10714,N_10514,N_10489);
nor U10715 (N_10715,N_10502,N_10472);
xor U10716 (N_10716,N_10516,N_10552);
nand U10717 (N_10717,N_10487,N_10435);
and U10718 (N_10718,N_10553,N_10559);
nand U10719 (N_10719,N_10534,N_10546);
xor U10720 (N_10720,N_10694,N_10641);
nor U10721 (N_10721,N_10696,N_10701);
and U10722 (N_10722,N_10585,N_10590);
and U10723 (N_10723,N_10693,N_10597);
xnor U10724 (N_10724,N_10710,N_10661);
nor U10725 (N_10725,N_10651,N_10708);
nand U10726 (N_10726,N_10596,N_10578);
and U10727 (N_10727,N_10591,N_10668);
xor U10728 (N_10728,N_10581,N_10574);
and U10729 (N_10729,N_10647,N_10659);
nor U10730 (N_10730,N_10677,N_10588);
nand U10731 (N_10731,N_10582,N_10717);
xor U10732 (N_10732,N_10594,N_10570);
xor U10733 (N_10733,N_10687,N_10667);
xnor U10734 (N_10734,N_10627,N_10719);
xor U10735 (N_10735,N_10691,N_10617);
nand U10736 (N_10736,N_10601,N_10619);
nand U10737 (N_10737,N_10600,N_10637);
or U10738 (N_10738,N_10663,N_10676);
xor U10739 (N_10739,N_10613,N_10683);
xnor U10740 (N_10740,N_10656,N_10699);
or U10741 (N_10741,N_10589,N_10603);
or U10742 (N_10742,N_10624,N_10629);
and U10743 (N_10743,N_10623,N_10568);
and U10744 (N_10744,N_10564,N_10658);
nand U10745 (N_10745,N_10572,N_10673);
or U10746 (N_10746,N_10604,N_10631);
nand U10747 (N_10747,N_10702,N_10657);
nor U10748 (N_10748,N_10680,N_10621);
and U10749 (N_10749,N_10586,N_10669);
or U10750 (N_10750,N_10714,N_10697);
xor U10751 (N_10751,N_10618,N_10615);
or U10752 (N_10752,N_10638,N_10614);
nor U10753 (N_10753,N_10703,N_10654);
nand U10754 (N_10754,N_10571,N_10704);
and U10755 (N_10755,N_10579,N_10635);
nand U10756 (N_10756,N_10715,N_10711);
and U10757 (N_10757,N_10632,N_10587);
nand U10758 (N_10758,N_10655,N_10607);
xor U10759 (N_10759,N_10608,N_10695);
or U10760 (N_10760,N_10679,N_10672);
xnor U10761 (N_10761,N_10573,N_10674);
nand U10762 (N_10762,N_10630,N_10653);
xor U10763 (N_10763,N_10716,N_10639);
xnor U10764 (N_10764,N_10584,N_10593);
and U10765 (N_10765,N_10684,N_10665);
nand U10766 (N_10766,N_10648,N_10622);
nor U10767 (N_10767,N_10628,N_10569);
nor U10768 (N_10768,N_10625,N_10636);
nand U10769 (N_10769,N_10712,N_10566);
nand U10770 (N_10770,N_10698,N_10670);
nand U10771 (N_10771,N_10664,N_10678);
and U10772 (N_10772,N_10685,N_10562);
nor U10773 (N_10773,N_10666,N_10690);
and U10774 (N_10774,N_10583,N_10643);
nand U10775 (N_10775,N_10646,N_10686);
nand U10776 (N_10776,N_10709,N_10692);
and U10777 (N_10777,N_10706,N_10689);
xor U10778 (N_10778,N_10700,N_10605);
nand U10779 (N_10779,N_10660,N_10563);
nor U10780 (N_10780,N_10645,N_10705);
xnor U10781 (N_10781,N_10565,N_10681);
nor U10782 (N_10782,N_10671,N_10575);
or U10783 (N_10783,N_10713,N_10598);
nor U10784 (N_10784,N_10649,N_10577);
or U10785 (N_10785,N_10662,N_10718);
nor U10786 (N_10786,N_10688,N_10560);
nor U10787 (N_10787,N_10561,N_10634);
and U10788 (N_10788,N_10602,N_10707);
xnor U10789 (N_10789,N_10611,N_10606);
nor U10790 (N_10790,N_10626,N_10652);
xor U10791 (N_10791,N_10620,N_10633);
xor U10792 (N_10792,N_10650,N_10616);
and U10793 (N_10793,N_10644,N_10612);
nor U10794 (N_10794,N_10567,N_10610);
nor U10795 (N_10795,N_10682,N_10592);
xnor U10796 (N_10796,N_10609,N_10640);
or U10797 (N_10797,N_10580,N_10576);
nor U10798 (N_10798,N_10642,N_10595);
nand U10799 (N_10799,N_10675,N_10599);
nor U10800 (N_10800,N_10632,N_10629);
and U10801 (N_10801,N_10632,N_10652);
nor U10802 (N_10802,N_10680,N_10595);
xor U10803 (N_10803,N_10717,N_10646);
nand U10804 (N_10804,N_10578,N_10709);
xor U10805 (N_10805,N_10711,N_10709);
or U10806 (N_10806,N_10636,N_10705);
nor U10807 (N_10807,N_10614,N_10658);
nor U10808 (N_10808,N_10623,N_10630);
nand U10809 (N_10809,N_10583,N_10609);
and U10810 (N_10810,N_10691,N_10578);
or U10811 (N_10811,N_10625,N_10560);
or U10812 (N_10812,N_10624,N_10602);
and U10813 (N_10813,N_10598,N_10603);
nor U10814 (N_10814,N_10653,N_10595);
xor U10815 (N_10815,N_10563,N_10678);
xnor U10816 (N_10816,N_10617,N_10668);
nor U10817 (N_10817,N_10627,N_10705);
or U10818 (N_10818,N_10630,N_10626);
xor U10819 (N_10819,N_10632,N_10581);
nand U10820 (N_10820,N_10631,N_10705);
or U10821 (N_10821,N_10614,N_10664);
nor U10822 (N_10822,N_10630,N_10599);
xnor U10823 (N_10823,N_10660,N_10662);
nor U10824 (N_10824,N_10624,N_10636);
nand U10825 (N_10825,N_10622,N_10667);
nor U10826 (N_10826,N_10655,N_10597);
or U10827 (N_10827,N_10630,N_10714);
and U10828 (N_10828,N_10656,N_10703);
nand U10829 (N_10829,N_10579,N_10700);
or U10830 (N_10830,N_10638,N_10606);
xnor U10831 (N_10831,N_10688,N_10676);
or U10832 (N_10832,N_10717,N_10714);
nand U10833 (N_10833,N_10601,N_10633);
xnor U10834 (N_10834,N_10650,N_10702);
or U10835 (N_10835,N_10571,N_10607);
or U10836 (N_10836,N_10605,N_10633);
nand U10837 (N_10837,N_10684,N_10676);
nor U10838 (N_10838,N_10703,N_10696);
xor U10839 (N_10839,N_10579,N_10641);
nand U10840 (N_10840,N_10682,N_10607);
nor U10841 (N_10841,N_10626,N_10710);
and U10842 (N_10842,N_10574,N_10705);
or U10843 (N_10843,N_10606,N_10645);
and U10844 (N_10844,N_10667,N_10628);
nand U10845 (N_10845,N_10604,N_10574);
and U10846 (N_10846,N_10696,N_10564);
or U10847 (N_10847,N_10686,N_10666);
xor U10848 (N_10848,N_10597,N_10564);
or U10849 (N_10849,N_10614,N_10657);
and U10850 (N_10850,N_10666,N_10590);
nor U10851 (N_10851,N_10711,N_10601);
xor U10852 (N_10852,N_10658,N_10655);
nor U10853 (N_10853,N_10665,N_10669);
and U10854 (N_10854,N_10688,N_10651);
xor U10855 (N_10855,N_10663,N_10683);
nor U10856 (N_10856,N_10711,N_10658);
nor U10857 (N_10857,N_10662,N_10639);
nand U10858 (N_10858,N_10640,N_10620);
nand U10859 (N_10859,N_10695,N_10586);
nor U10860 (N_10860,N_10571,N_10635);
nor U10861 (N_10861,N_10567,N_10624);
and U10862 (N_10862,N_10694,N_10670);
nor U10863 (N_10863,N_10634,N_10685);
or U10864 (N_10864,N_10610,N_10599);
xnor U10865 (N_10865,N_10660,N_10644);
or U10866 (N_10866,N_10615,N_10560);
and U10867 (N_10867,N_10712,N_10618);
xnor U10868 (N_10868,N_10677,N_10626);
or U10869 (N_10869,N_10663,N_10695);
or U10870 (N_10870,N_10612,N_10631);
nor U10871 (N_10871,N_10613,N_10658);
and U10872 (N_10872,N_10598,N_10687);
nand U10873 (N_10873,N_10658,N_10610);
and U10874 (N_10874,N_10703,N_10637);
and U10875 (N_10875,N_10582,N_10632);
xnor U10876 (N_10876,N_10615,N_10661);
xor U10877 (N_10877,N_10632,N_10670);
and U10878 (N_10878,N_10684,N_10564);
nand U10879 (N_10879,N_10614,N_10684);
nand U10880 (N_10880,N_10831,N_10769);
nand U10881 (N_10881,N_10746,N_10740);
and U10882 (N_10882,N_10739,N_10817);
or U10883 (N_10883,N_10851,N_10869);
xor U10884 (N_10884,N_10840,N_10835);
xnor U10885 (N_10885,N_10824,N_10809);
and U10886 (N_10886,N_10850,N_10820);
or U10887 (N_10887,N_10808,N_10759);
or U10888 (N_10888,N_10781,N_10826);
or U10889 (N_10889,N_10842,N_10816);
or U10890 (N_10890,N_10731,N_10878);
or U10891 (N_10891,N_10829,N_10868);
nand U10892 (N_10892,N_10786,N_10763);
or U10893 (N_10893,N_10794,N_10762);
nand U10894 (N_10894,N_10742,N_10775);
nor U10895 (N_10895,N_10795,N_10862);
nor U10896 (N_10896,N_10784,N_10844);
and U10897 (N_10897,N_10877,N_10753);
nand U10898 (N_10898,N_10803,N_10825);
nor U10899 (N_10899,N_10870,N_10756);
or U10900 (N_10900,N_10791,N_10744);
xor U10901 (N_10901,N_10777,N_10773);
and U10902 (N_10902,N_10818,N_10755);
nor U10903 (N_10903,N_10819,N_10738);
and U10904 (N_10904,N_10858,N_10843);
xnor U10905 (N_10905,N_10792,N_10864);
xnor U10906 (N_10906,N_10758,N_10785);
or U10907 (N_10907,N_10853,N_10872);
and U10908 (N_10908,N_10730,N_10866);
and U10909 (N_10909,N_10836,N_10724);
or U10910 (N_10910,N_10726,N_10747);
xnor U10911 (N_10911,N_10827,N_10774);
xor U10912 (N_10912,N_10722,N_10749);
and U10913 (N_10913,N_10736,N_10783);
nand U10914 (N_10914,N_10790,N_10799);
nand U10915 (N_10915,N_10779,N_10751);
or U10916 (N_10916,N_10754,N_10834);
xor U10917 (N_10917,N_10838,N_10855);
and U10918 (N_10918,N_10806,N_10802);
xor U10919 (N_10919,N_10796,N_10801);
xor U10920 (N_10920,N_10778,N_10768);
nand U10921 (N_10921,N_10760,N_10772);
nor U10922 (N_10922,N_10788,N_10805);
nor U10923 (N_10923,N_10734,N_10797);
and U10924 (N_10924,N_10752,N_10847);
nand U10925 (N_10925,N_10861,N_10743);
nor U10926 (N_10926,N_10839,N_10776);
nand U10927 (N_10927,N_10745,N_10807);
nor U10928 (N_10928,N_10871,N_10757);
or U10929 (N_10929,N_10782,N_10863);
nor U10930 (N_10930,N_10879,N_10764);
or U10931 (N_10931,N_10767,N_10787);
nor U10932 (N_10932,N_10798,N_10728);
and U10933 (N_10933,N_10735,N_10780);
xor U10934 (N_10934,N_10837,N_10852);
and U10935 (N_10935,N_10748,N_10765);
nor U10936 (N_10936,N_10854,N_10857);
and U10937 (N_10937,N_10800,N_10789);
nand U10938 (N_10938,N_10741,N_10811);
xnor U10939 (N_10939,N_10732,N_10812);
nor U10940 (N_10940,N_10873,N_10733);
xor U10941 (N_10941,N_10848,N_10721);
nor U10942 (N_10942,N_10729,N_10867);
or U10943 (N_10943,N_10723,N_10828);
xnor U10944 (N_10944,N_10833,N_10813);
nand U10945 (N_10945,N_10727,N_10750);
nor U10946 (N_10946,N_10849,N_10804);
and U10947 (N_10947,N_10770,N_10771);
and U10948 (N_10948,N_10793,N_10720);
xor U10949 (N_10949,N_10856,N_10822);
nand U10950 (N_10950,N_10814,N_10815);
nand U10951 (N_10951,N_10766,N_10821);
nand U10952 (N_10952,N_10761,N_10841);
and U10953 (N_10953,N_10875,N_10845);
nor U10954 (N_10954,N_10737,N_10832);
and U10955 (N_10955,N_10865,N_10823);
nor U10956 (N_10956,N_10874,N_10846);
nor U10957 (N_10957,N_10859,N_10876);
or U10958 (N_10958,N_10810,N_10860);
nand U10959 (N_10959,N_10830,N_10725);
xor U10960 (N_10960,N_10741,N_10821);
nor U10961 (N_10961,N_10728,N_10736);
or U10962 (N_10962,N_10870,N_10729);
nand U10963 (N_10963,N_10851,N_10875);
or U10964 (N_10964,N_10846,N_10841);
nand U10965 (N_10965,N_10844,N_10815);
and U10966 (N_10966,N_10726,N_10771);
nor U10967 (N_10967,N_10830,N_10842);
and U10968 (N_10968,N_10792,N_10723);
and U10969 (N_10969,N_10871,N_10729);
nor U10970 (N_10970,N_10759,N_10805);
nor U10971 (N_10971,N_10804,N_10756);
and U10972 (N_10972,N_10764,N_10790);
xor U10973 (N_10973,N_10865,N_10778);
or U10974 (N_10974,N_10738,N_10787);
or U10975 (N_10975,N_10773,N_10741);
nand U10976 (N_10976,N_10797,N_10795);
and U10977 (N_10977,N_10778,N_10743);
nand U10978 (N_10978,N_10787,N_10797);
nor U10979 (N_10979,N_10730,N_10759);
xnor U10980 (N_10980,N_10750,N_10759);
nor U10981 (N_10981,N_10849,N_10801);
xnor U10982 (N_10982,N_10847,N_10742);
nor U10983 (N_10983,N_10819,N_10727);
or U10984 (N_10984,N_10793,N_10732);
nand U10985 (N_10985,N_10808,N_10833);
nor U10986 (N_10986,N_10755,N_10780);
or U10987 (N_10987,N_10800,N_10790);
nor U10988 (N_10988,N_10814,N_10737);
nor U10989 (N_10989,N_10808,N_10814);
nor U10990 (N_10990,N_10725,N_10847);
xor U10991 (N_10991,N_10778,N_10815);
or U10992 (N_10992,N_10724,N_10730);
and U10993 (N_10993,N_10744,N_10853);
or U10994 (N_10994,N_10765,N_10786);
nor U10995 (N_10995,N_10797,N_10785);
nor U10996 (N_10996,N_10775,N_10862);
and U10997 (N_10997,N_10766,N_10772);
nor U10998 (N_10998,N_10875,N_10865);
nand U10999 (N_10999,N_10758,N_10781);
or U11000 (N_11000,N_10746,N_10745);
nor U11001 (N_11001,N_10854,N_10796);
or U11002 (N_11002,N_10752,N_10857);
nor U11003 (N_11003,N_10800,N_10756);
and U11004 (N_11004,N_10729,N_10810);
and U11005 (N_11005,N_10742,N_10752);
nor U11006 (N_11006,N_10765,N_10733);
nand U11007 (N_11007,N_10810,N_10766);
or U11008 (N_11008,N_10846,N_10809);
nor U11009 (N_11009,N_10750,N_10801);
and U11010 (N_11010,N_10804,N_10867);
nor U11011 (N_11011,N_10855,N_10756);
nor U11012 (N_11012,N_10812,N_10761);
and U11013 (N_11013,N_10761,N_10827);
nor U11014 (N_11014,N_10831,N_10877);
xor U11015 (N_11015,N_10860,N_10766);
or U11016 (N_11016,N_10801,N_10832);
xor U11017 (N_11017,N_10754,N_10819);
and U11018 (N_11018,N_10790,N_10798);
xnor U11019 (N_11019,N_10849,N_10760);
nand U11020 (N_11020,N_10876,N_10872);
and U11021 (N_11021,N_10795,N_10812);
xor U11022 (N_11022,N_10721,N_10852);
or U11023 (N_11023,N_10776,N_10742);
nand U11024 (N_11024,N_10761,N_10752);
nand U11025 (N_11025,N_10821,N_10772);
nand U11026 (N_11026,N_10858,N_10815);
nand U11027 (N_11027,N_10768,N_10862);
nor U11028 (N_11028,N_10843,N_10789);
and U11029 (N_11029,N_10818,N_10793);
and U11030 (N_11030,N_10738,N_10800);
or U11031 (N_11031,N_10836,N_10849);
and U11032 (N_11032,N_10744,N_10873);
xor U11033 (N_11033,N_10841,N_10850);
xor U11034 (N_11034,N_10726,N_10828);
nand U11035 (N_11035,N_10775,N_10832);
or U11036 (N_11036,N_10740,N_10823);
or U11037 (N_11037,N_10862,N_10820);
nand U11038 (N_11038,N_10777,N_10814);
xor U11039 (N_11039,N_10772,N_10807);
xnor U11040 (N_11040,N_11013,N_10921);
xnor U11041 (N_11041,N_10947,N_11023);
nand U11042 (N_11042,N_10881,N_10903);
nor U11043 (N_11043,N_11016,N_11039);
nor U11044 (N_11044,N_11031,N_10968);
nand U11045 (N_11045,N_10949,N_10977);
nand U11046 (N_11046,N_10988,N_10953);
and U11047 (N_11047,N_10914,N_10969);
nand U11048 (N_11048,N_11011,N_10961);
nand U11049 (N_11049,N_10962,N_11022);
nor U11050 (N_11050,N_10916,N_10910);
or U11051 (N_11051,N_11019,N_10993);
xnor U11052 (N_11052,N_10981,N_10918);
nor U11053 (N_11053,N_10941,N_10913);
or U11054 (N_11054,N_10912,N_10898);
xor U11055 (N_11055,N_10985,N_10885);
or U11056 (N_11056,N_10952,N_10960);
and U11057 (N_11057,N_10928,N_10989);
nand U11058 (N_11058,N_10930,N_10958);
nand U11059 (N_11059,N_10964,N_11004);
nor U11060 (N_11060,N_11018,N_10896);
nand U11061 (N_11061,N_11028,N_10939);
and U11062 (N_11062,N_10927,N_10976);
nand U11063 (N_11063,N_10967,N_10932);
nor U11064 (N_11064,N_10999,N_11014);
or U11065 (N_11065,N_10938,N_10984);
xnor U11066 (N_11066,N_10917,N_10929);
and U11067 (N_11067,N_10966,N_11002);
xor U11068 (N_11068,N_10986,N_10888);
nand U11069 (N_11069,N_10899,N_10924);
nand U11070 (N_11070,N_10959,N_10973);
xnor U11071 (N_11071,N_10950,N_10894);
nand U11072 (N_11072,N_10905,N_10978);
and U11073 (N_11073,N_10884,N_10880);
xor U11074 (N_11074,N_10995,N_10900);
xnor U11075 (N_11075,N_10925,N_10911);
xor U11076 (N_11076,N_10886,N_10987);
and U11077 (N_11077,N_10994,N_10890);
nand U11078 (N_11078,N_10972,N_10943);
and U11079 (N_11079,N_10992,N_10934);
or U11080 (N_11080,N_10957,N_11035);
nor U11081 (N_11081,N_10895,N_10990);
and U11082 (N_11082,N_11020,N_11029);
or U11083 (N_11083,N_10909,N_10982);
nand U11084 (N_11084,N_11000,N_11037);
or U11085 (N_11085,N_11012,N_11005);
nand U11086 (N_11086,N_11021,N_10904);
or U11087 (N_11087,N_10974,N_10954);
or U11088 (N_11088,N_10979,N_10906);
nor U11089 (N_11089,N_10883,N_10956);
nand U11090 (N_11090,N_10935,N_10902);
nand U11091 (N_11091,N_10889,N_10948);
nand U11092 (N_11092,N_10998,N_10975);
or U11093 (N_11093,N_10887,N_10971);
or U11094 (N_11094,N_11010,N_10965);
or U11095 (N_11095,N_11015,N_10919);
or U11096 (N_11096,N_10945,N_11026);
nor U11097 (N_11097,N_11027,N_11030);
or U11098 (N_11098,N_10996,N_11017);
or U11099 (N_11099,N_10897,N_10908);
and U11100 (N_11100,N_10951,N_10907);
or U11101 (N_11101,N_10920,N_10931);
and U11102 (N_11102,N_10901,N_11006);
xnor U11103 (N_11103,N_11024,N_11032);
nand U11104 (N_11104,N_11036,N_10922);
and U11105 (N_11105,N_11034,N_11008);
or U11106 (N_11106,N_10980,N_10926);
xor U11107 (N_11107,N_10915,N_11038);
xnor U11108 (N_11108,N_10937,N_10892);
nand U11109 (N_11109,N_11033,N_10940);
nand U11110 (N_11110,N_10997,N_10944);
and U11111 (N_11111,N_10923,N_10933);
xor U11112 (N_11112,N_10893,N_11007);
nor U11113 (N_11113,N_11009,N_10946);
or U11114 (N_11114,N_10942,N_10970);
nand U11115 (N_11115,N_10963,N_11001);
nand U11116 (N_11116,N_10891,N_11003);
or U11117 (N_11117,N_10936,N_10991);
xnor U11118 (N_11118,N_10882,N_10983);
xnor U11119 (N_11119,N_11025,N_10955);
xnor U11120 (N_11120,N_10964,N_11016);
nand U11121 (N_11121,N_10895,N_10899);
nand U11122 (N_11122,N_10974,N_10880);
nand U11123 (N_11123,N_10972,N_11035);
and U11124 (N_11124,N_11003,N_10954);
nand U11125 (N_11125,N_10960,N_10896);
nand U11126 (N_11126,N_10928,N_11035);
or U11127 (N_11127,N_10990,N_10884);
nand U11128 (N_11128,N_11030,N_10932);
and U11129 (N_11129,N_10924,N_10946);
xnor U11130 (N_11130,N_10934,N_10932);
nand U11131 (N_11131,N_10893,N_11033);
xnor U11132 (N_11132,N_10975,N_10899);
nand U11133 (N_11133,N_10982,N_10915);
nand U11134 (N_11134,N_10916,N_10983);
nor U11135 (N_11135,N_10964,N_10948);
xnor U11136 (N_11136,N_10940,N_11027);
nor U11137 (N_11137,N_10995,N_11023);
nand U11138 (N_11138,N_10952,N_10913);
and U11139 (N_11139,N_10967,N_11007);
nand U11140 (N_11140,N_11011,N_10901);
nand U11141 (N_11141,N_10903,N_10990);
nand U11142 (N_11142,N_11015,N_11001);
and U11143 (N_11143,N_10954,N_10978);
or U11144 (N_11144,N_10942,N_10941);
or U11145 (N_11145,N_11007,N_11022);
and U11146 (N_11146,N_11001,N_10971);
and U11147 (N_11147,N_10987,N_11016);
or U11148 (N_11148,N_11009,N_10933);
xor U11149 (N_11149,N_11009,N_10966);
xnor U11150 (N_11150,N_11006,N_10884);
nor U11151 (N_11151,N_10895,N_10967);
nand U11152 (N_11152,N_10963,N_10976);
xnor U11153 (N_11153,N_10929,N_10984);
nor U11154 (N_11154,N_11015,N_10961);
xnor U11155 (N_11155,N_10923,N_10912);
nor U11156 (N_11156,N_10974,N_10931);
nand U11157 (N_11157,N_10955,N_10978);
nand U11158 (N_11158,N_10896,N_10918);
or U11159 (N_11159,N_11009,N_10923);
nor U11160 (N_11160,N_11022,N_10882);
nor U11161 (N_11161,N_10914,N_10897);
or U11162 (N_11162,N_10891,N_10924);
xor U11163 (N_11163,N_10947,N_10904);
xor U11164 (N_11164,N_10915,N_10992);
nand U11165 (N_11165,N_11020,N_10919);
xnor U11166 (N_11166,N_10939,N_10906);
or U11167 (N_11167,N_11037,N_10979);
xnor U11168 (N_11168,N_10905,N_10958);
or U11169 (N_11169,N_10948,N_10931);
and U11170 (N_11170,N_10934,N_10904);
and U11171 (N_11171,N_10956,N_10885);
nand U11172 (N_11172,N_10921,N_10886);
or U11173 (N_11173,N_10980,N_10975);
xnor U11174 (N_11174,N_10896,N_11014);
or U11175 (N_11175,N_10959,N_11033);
and U11176 (N_11176,N_10941,N_10890);
nor U11177 (N_11177,N_10883,N_10962);
nand U11178 (N_11178,N_10926,N_10957);
and U11179 (N_11179,N_10929,N_10989);
and U11180 (N_11180,N_11025,N_10941);
nor U11181 (N_11181,N_10921,N_10992);
xor U11182 (N_11182,N_10945,N_11036);
and U11183 (N_11183,N_10943,N_10888);
nor U11184 (N_11184,N_11018,N_11004);
nand U11185 (N_11185,N_10926,N_10901);
nand U11186 (N_11186,N_10909,N_10912);
nand U11187 (N_11187,N_10999,N_10948);
and U11188 (N_11188,N_10939,N_10937);
and U11189 (N_11189,N_10958,N_10922);
xor U11190 (N_11190,N_10895,N_11034);
nor U11191 (N_11191,N_10950,N_10956);
or U11192 (N_11192,N_10988,N_10918);
nor U11193 (N_11193,N_11011,N_10997);
xor U11194 (N_11194,N_10969,N_10910);
nor U11195 (N_11195,N_10880,N_10955);
xor U11196 (N_11196,N_11004,N_10905);
or U11197 (N_11197,N_11032,N_10996);
nor U11198 (N_11198,N_10983,N_10953);
xnor U11199 (N_11199,N_10946,N_10983);
and U11200 (N_11200,N_11064,N_11164);
nor U11201 (N_11201,N_11079,N_11161);
nand U11202 (N_11202,N_11199,N_11067);
or U11203 (N_11203,N_11175,N_11101);
nand U11204 (N_11204,N_11179,N_11166);
and U11205 (N_11205,N_11147,N_11050);
nand U11206 (N_11206,N_11138,N_11132);
xor U11207 (N_11207,N_11140,N_11070);
and U11208 (N_11208,N_11053,N_11169);
nand U11209 (N_11209,N_11194,N_11061);
and U11210 (N_11210,N_11190,N_11085);
nand U11211 (N_11211,N_11165,N_11174);
or U11212 (N_11212,N_11154,N_11089);
nor U11213 (N_11213,N_11171,N_11082);
and U11214 (N_11214,N_11058,N_11040);
nand U11215 (N_11215,N_11100,N_11110);
nor U11216 (N_11216,N_11097,N_11080);
and U11217 (N_11217,N_11156,N_11133);
nor U11218 (N_11218,N_11098,N_11111);
or U11219 (N_11219,N_11184,N_11178);
nand U11220 (N_11220,N_11074,N_11120);
xor U11221 (N_11221,N_11108,N_11115);
nor U11222 (N_11222,N_11045,N_11162);
xnor U11223 (N_11223,N_11196,N_11087);
or U11224 (N_11224,N_11103,N_11060);
xnor U11225 (N_11225,N_11136,N_11055);
xor U11226 (N_11226,N_11130,N_11091);
nand U11227 (N_11227,N_11168,N_11192);
nor U11228 (N_11228,N_11076,N_11094);
and U11229 (N_11229,N_11057,N_11145);
xnor U11230 (N_11230,N_11170,N_11127);
and U11231 (N_11231,N_11056,N_11105);
nor U11232 (N_11232,N_11177,N_11143);
nor U11233 (N_11233,N_11137,N_11153);
xor U11234 (N_11234,N_11066,N_11112);
or U11235 (N_11235,N_11123,N_11046);
xnor U11236 (N_11236,N_11104,N_11180);
and U11237 (N_11237,N_11191,N_11187);
xnor U11238 (N_11238,N_11099,N_11129);
nand U11239 (N_11239,N_11186,N_11193);
and U11240 (N_11240,N_11047,N_11197);
and U11241 (N_11241,N_11107,N_11146);
and U11242 (N_11242,N_11135,N_11072);
xor U11243 (N_11243,N_11078,N_11041);
nor U11244 (N_11244,N_11086,N_11158);
and U11245 (N_11245,N_11155,N_11151);
xor U11246 (N_11246,N_11126,N_11185);
nor U11247 (N_11247,N_11048,N_11149);
nor U11248 (N_11248,N_11157,N_11084);
or U11249 (N_11249,N_11139,N_11198);
or U11250 (N_11250,N_11077,N_11106);
xor U11251 (N_11251,N_11063,N_11065);
and U11252 (N_11252,N_11043,N_11068);
nor U11253 (N_11253,N_11118,N_11042);
nor U11254 (N_11254,N_11071,N_11081);
xnor U11255 (N_11255,N_11114,N_11172);
nand U11256 (N_11256,N_11054,N_11141);
xor U11257 (N_11257,N_11173,N_11128);
and U11258 (N_11258,N_11052,N_11090);
xnor U11259 (N_11259,N_11044,N_11119);
and U11260 (N_11260,N_11117,N_11116);
nor U11261 (N_11261,N_11113,N_11142);
nor U11262 (N_11262,N_11183,N_11181);
nor U11263 (N_11263,N_11095,N_11102);
nand U11264 (N_11264,N_11167,N_11131);
and U11265 (N_11265,N_11134,N_11069);
and U11266 (N_11266,N_11122,N_11195);
nand U11267 (N_11267,N_11189,N_11083);
nand U11268 (N_11268,N_11096,N_11093);
nor U11269 (N_11269,N_11188,N_11125);
xnor U11270 (N_11270,N_11051,N_11152);
nor U11271 (N_11271,N_11176,N_11124);
xor U11272 (N_11272,N_11150,N_11163);
xor U11273 (N_11273,N_11109,N_11059);
nor U11274 (N_11274,N_11088,N_11121);
and U11275 (N_11275,N_11144,N_11148);
nand U11276 (N_11276,N_11092,N_11182);
xnor U11277 (N_11277,N_11062,N_11160);
nand U11278 (N_11278,N_11049,N_11073);
or U11279 (N_11279,N_11075,N_11159);
or U11280 (N_11280,N_11103,N_11142);
nor U11281 (N_11281,N_11089,N_11104);
or U11282 (N_11282,N_11163,N_11133);
and U11283 (N_11283,N_11186,N_11057);
xor U11284 (N_11284,N_11042,N_11056);
nor U11285 (N_11285,N_11041,N_11188);
nor U11286 (N_11286,N_11070,N_11164);
and U11287 (N_11287,N_11160,N_11058);
xor U11288 (N_11288,N_11070,N_11089);
or U11289 (N_11289,N_11043,N_11186);
xor U11290 (N_11290,N_11180,N_11097);
and U11291 (N_11291,N_11125,N_11077);
nor U11292 (N_11292,N_11097,N_11188);
and U11293 (N_11293,N_11082,N_11180);
xor U11294 (N_11294,N_11048,N_11136);
nor U11295 (N_11295,N_11107,N_11171);
and U11296 (N_11296,N_11144,N_11081);
nor U11297 (N_11297,N_11101,N_11076);
xor U11298 (N_11298,N_11063,N_11126);
or U11299 (N_11299,N_11079,N_11065);
xor U11300 (N_11300,N_11134,N_11189);
xnor U11301 (N_11301,N_11160,N_11073);
and U11302 (N_11302,N_11048,N_11123);
nor U11303 (N_11303,N_11077,N_11101);
nor U11304 (N_11304,N_11145,N_11062);
nor U11305 (N_11305,N_11176,N_11106);
nand U11306 (N_11306,N_11166,N_11191);
xnor U11307 (N_11307,N_11161,N_11046);
xor U11308 (N_11308,N_11129,N_11071);
nor U11309 (N_11309,N_11105,N_11137);
nand U11310 (N_11310,N_11171,N_11096);
xor U11311 (N_11311,N_11136,N_11190);
xor U11312 (N_11312,N_11121,N_11110);
or U11313 (N_11313,N_11069,N_11087);
xor U11314 (N_11314,N_11059,N_11195);
nand U11315 (N_11315,N_11187,N_11049);
nor U11316 (N_11316,N_11074,N_11058);
nand U11317 (N_11317,N_11171,N_11066);
or U11318 (N_11318,N_11182,N_11086);
nor U11319 (N_11319,N_11074,N_11185);
and U11320 (N_11320,N_11138,N_11141);
nand U11321 (N_11321,N_11119,N_11176);
nand U11322 (N_11322,N_11164,N_11040);
nor U11323 (N_11323,N_11113,N_11085);
xnor U11324 (N_11324,N_11154,N_11140);
and U11325 (N_11325,N_11072,N_11042);
or U11326 (N_11326,N_11049,N_11196);
xnor U11327 (N_11327,N_11098,N_11049);
nor U11328 (N_11328,N_11172,N_11048);
nor U11329 (N_11329,N_11111,N_11179);
nand U11330 (N_11330,N_11124,N_11192);
and U11331 (N_11331,N_11053,N_11121);
nand U11332 (N_11332,N_11199,N_11143);
xnor U11333 (N_11333,N_11042,N_11070);
xnor U11334 (N_11334,N_11074,N_11194);
nor U11335 (N_11335,N_11081,N_11065);
and U11336 (N_11336,N_11153,N_11188);
and U11337 (N_11337,N_11116,N_11181);
nor U11338 (N_11338,N_11095,N_11120);
and U11339 (N_11339,N_11121,N_11066);
nand U11340 (N_11340,N_11196,N_11127);
or U11341 (N_11341,N_11191,N_11174);
nand U11342 (N_11342,N_11176,N_11088);
or U11343 (N_11343,N_11058,N_11059);
or U11344 (N_11344,N_11170,N_11064);
xor U11345 (N_11345,N_11188,N_11096);
nand U11346 (N_11346,N_11053,N_11071);
nor U11347 (N_11347,N_11087,N_11188);
or U11348 (N_11348,N_11070,N_11186);
or U11349 (N_11349,N_11166,N_11137);
or U11350 (N_11350,N_11083,N_11165);
and U11351 (N_11351,N_11186,N_11140);
and U11352 (N_11352,N_11171,N_11167);
or U11353 (N_11353,N_11106,N_11067);
or U11354 (N_11354,N_11110,N_11127);
xor U11355 (N_11355,N_11152,N_11141);
xnor U11356 (N_11356,N_11115,N_11068);
or U11357 (N_11357,N_11176,N_11065);
xnor U11358 (N_11358,N_11126,N_11045);
xnor U11359 (N_11359,N_11124,N_11043);
nor U11360 (N_11360,N_11222,N_11308);
nor U11361 (N_11361,N_11228,N_11253);
and U11362 (N_11362,N_11355,N_11224);
nor U11363 (N_11363,N_11242,N_11268);
nand U11364 (N_11364,N_11205,N_11338);
nand U11365 (N_11365,N_11225,N_11325);
nor U11366 (N_11366,N_11203,N_11288);
nor U11367 (N_11367,N_11356,N_11216);
xor U11368 (N_11368,N_11285,N_11235);
nor U11369 (N_11369,N_11358,N_11316);
nand U11370 (N_11370,N_11299,N_11321);
and U11371 (N_11371,N_11256,N_11324);
xor U11372 (N_11372,N_11234,N_11238);
or U11373 (N_11373,N_11221,N_11293);
xnor U11374 (N_11374,N_11319,N_11204);
or U11375 (N_11375,N_11352,N_11271);
and U11376 (N_11376,N_11229,N_11315);
or U11377 (N_11377,N_11211,N_11275);
nor U11378 (N_11378,N_11359,N_11334);
xnor U11379 (N_11379,N_11241,N_11236);
or U11380 (N_11380,N_11313,N_11220);
and U11381 (N_11381,N_11263,N_11303);
nor U11382 (N_11382,N_11245,N_11255);
xor U11383 (N_11383,N_11342,N_11344);
xor U11384 (N_11384,N_11298,N_11232);
nor U11385 (N_11385,N_11200,N_11257);
nand U11386 (N_11386,N_11294,N_11348);
nand U11387 (N_11387,N_11331,N_11300);
xor U11388 (N_11388,N_11329,N_11231);
nand U11389 (N_11389,N_11286,N_11304);
nand U11390 (N_11390,N_11320,N_11297);
xor U11391 (N_11391,N_11357,N_11354);
or U11392 (N_11392,N_11290,N_11261);
or U11393 (N_11393,N_11206,N_11323);
nand U11394 (N_11394,N_11289,N_11322);
nand U11395 (N_11395,N_11353,N_11283);
nand U11396 (N_11396,N_11247,N_11274);
nor U11397 (N_11397,N_11328,N_11291);
and U11398 (N_11398,N_11260,N_11239);
nand U11399 (N_11399,N_11351,N_11250);
xnor U11400 (N_11400,N_11267,N_11207);
and U11401 (N_11401,N_11270,N_11292);
nand U11402 (N_11402,N_11233,N_11332);
nor U11403 (N_11403,N_11347,N_11223);
nor U11404 (N_11404,N_11210,N_11341);
nor U11405 (N_11405,N_11310,N_11251);
nand U11406 (N_11406,N_11244,N_11213);
or U11407 (N_11407,N_11301,N_11230);
or U11408 (N_11408,N_11284,N_11227);
and U11409 (N_11409,N_11214,N_11278);
and U11410 (N_11410,N_11266,N_11287);
xnor U11411 (N_11411,N_11340,N_11208);
nor U11412 (N_11412,N_11350,N_11277);
nand U11413 (N_11413,N_11279,N_11307);
nand U11414 (N_11414,N_11309,N_11265);
xor U11415 (N_11415,N_11248,N_11312);
and U11416 (N_11416,N_11217,N_11249);
xnor U11417 (N_11417,N_11243,N_11259);
nand U11418 (N_11418,N_11314,N_11306);
or U11419 (N_11419,N_11252,N_11311);
or U11420 (N_11420,N_11218,N_11345);
or U11421 (N_11421,N_11246,N_11343);
nor U11422 (N_11422,N_11269,N_11282);
nand U11423 (N_11423,N_11226,N_11272);
or U11424 (N_11424,N_11317,N_11336);
nand U11425 (N_11425,N_11280,N_11296);
xnor U11426 (N_11426,N_11281,N_11215);
nor U11427 (N_11427,N_11209,N_11330);
or U11428 (N_11428,N_11349,N_11318);
and U11429 (N_11429,N_11276,N_11258);
nor U11430 (N_11430,N_11202,N_11302);
xnor U11431 (N_11431,N_11254,N_11262);
nand U11432 (N_11432,N_11264,N_11305);
or U11433 (N_11433,N_11273,N_11212);
or U11434 (N_11434,N_11240,N_11335);
and U11435 (N_11435,N_11327,N_11295);
xnor U11436 (N_11436,N_11201,N_11339);
nor U11437 (N_11437,N_11237,N_11219);
or U11438 (N_11438,N_11326,N_11346);
nor U11439 (N_11439,N_11333,N_11337);
nor U11440 (N_11440,N_11265,N_11291);
nand U11441 (N_11441,N_11310,N_11357);
nand U11442 (N_11442,N_11343,N_11332);
xor U11443 (N_11443,N_11321,N_11320);
xor U11444 (N_11444,N_11272,N_11336);
nand U11445 (N_11445,N_11257,N_11273);
nor U11446 (N_11446,N_11219,N_11297);
and U11447 (N_11447,N_11296,N_11335);
and U11448 (N_11448,N_11245,N_11208);
xnor U11449 (N_11449,N_11218,N_11295);
or U11450 (N_11450,N_11283,N_11241);
or U11451 (N_11451,N_11298,N_11336);
and U11452 (N_11452,N_11223,N_11275);
and U11453 (N_11453,N_11245,N_11321);
or U11454 (N_11454,N_11219,N_11319);
nor U11455 (N_11455,N_11303,N_11316);
or U11456 (N_11456,N_11212,N_11293);
xnor U11457 (N_11457,N_11352,N_11228);
nor U11458 (N_11458,N_11350,N_11222);
xnor U11459 (N_11459,N_11354,N_11342);
and U11460 (N_11460,N_11267,N_11321);
xnor U11461 (N_11461,N_11338,N_11216);
xor U11462 (N_11462,N_11323,N_11297);
and U11463 (N_11463,N_11211,N_11215);
nor U11464 (N_11464,N_11345,N_11328);
and U11465 (N_11465,N_11357,N_11341);
xnor U11466 (N_11466,N_11354,N_11233);
or U11467 (N_11467,N_11321,N_11282);
or U11468 (N_11468,N_11215,N_11261);
nor U11469 (N_11469,N_11218,N_11259);
xor U11470 (N_11470,N_11243,N_11298);
nand U11471 (N_11471,N_11316,N_11326);
xor U11472 (N_11472,N_11336,N_11294);
or U11473 (N_11473,N_11355,N_11335);
xor U11474 (N_11474,N_11207,N_11223);
xnor U11475 (N_11475,N_11358,N_11229);
or U11476 (N_11476,N_11303,N_11302);
and U11477 (N_11477,N_11355,N_11232);
xor U11478 (N_11478,N_11291,N_11257);
xnor U11479 (N_11479,N_11347,N_11272);
and U11480 (N_11480,N_11269,N_11349);
nand U11481 (N_11481,N_11217,N_11301);
nor U11482 (N_11482,N_11240,N_11331);
or U11483 (N_11483,N_11247,N_11267);
xor U11484 (N_11484,N_11327,N_11279);
xnor U11485 (N_11485,N_11269,N_11292);
nand U11486 (N_11486,N_11339,N_11318);
nor U11487 (N_11487,N_11304,N_11231);
nand U11488 (N_11488,N_11249,N_11237);
nor U11489 (N_11489,N_11320,N_11275);
or U11490 (N_11490,N_11200,N_11353);
xnor U11491 (N_11491,N_11220,N_11296);
and U11492 (N_11492,N_11321,N_11244);
xor U11493 (N_11493,N_11259,N_11354);
and U11494 (N_11494,N_11339,N_11329);
xor U11495 (N_11495,N_11311,N_11216);
or U11496 (N_11496,N_11249,N_11244);
nor U11497 (N_11497,N_11285,N_11240);
nand U11498 (N_11498,N_11246,N_11287);
nand U11499 (N_11499,N_11244,N_11340);
or U11500 (N_11500,N_11242,N_11308);
and U11501 (N_11501,N_11205,N_11309);
nor U11502 (N_11502,N_11214,N_11291);
or U11503 (N_11503,N_11233,N_11316);
nor U11504 (N_11504,N_11230,N_11333);
nor U11505 (N_11505,N_11264,N_11263);
nand U11506 (N_11506,N_11222,N_11264);
nor U11507 (N_11507,N_11214,N_11213);
or U11508 (N_11508,N_11299,N_11272);
or U11509 (N_11509,N_11338,N_11325);
nand U11510 (N_11510,N_11314,N_11335);
nor U11511 (N_11511,N_11298,N_11270);
and U11512 (N_11512,N_11345,N_11298);
xnor U11513 (N_11513,N_11244,N_11317);
nand U11514 (N_11514,N_11269,N_11237);
or U11515 (N_11515,N_11232,N_11312);
nand U11516 (N_11516,N_11343,N_11216);
or U11517 (N_11517,N_11228,N_11279);
xnor U11518 (N_11518,N_11271,N_11316);
or U11519 (N_11519,N_11207,N_11203);
or U11520 (N_11520,N_11388,N_11447);
nor U11521 (N_11521,N_11370,N_11365);
or U11522 (N_11522,N_11476,N_11462);
xnor U11523 (N_11523,N_11366,N_11402);
and U11524 (N_11524,N_11409,N_11401);
xnor U11525 (N_11525,N_11493,N_11516);
or U11526 (N_11526,N_11491,N_11427);
xor U11527 (N_11527,N_11441,N_11423);
nor U11528 (N_11528,N_11430,N_11501);
or U11529 (N_11529,N_11385,N_11383);
nor U11530 (N_11530,N_11478,N_11456);
or U11531 (N_11531,N_11407,N_11368);
nand U11532 (N_11532,N_11420,N_11472);
xnor U11533 (N_11533,N_11468,N_11475);
xor U11534 (N_11534,N_11486,N_11463);
nor U11535 (N_11535,N_11375,N_11504);
and U11536 (N_11536,N_11473,N_11469);
xnor U11537 (N_11537,N_11363,N_11386);
nand U11538 (N_11538,N_11442,N_11377);
or U11539 (N_11539,N_11513,N_11519);
and U11540 (N_11540,N_11380,N_11371);
nor U11541 (N_11541,N_11431,N_11412);
nor U11542 (N_11542,N_11507,N_11429);
nand U11543 (N_11543,N_11360,N_11499);
nor U11544 (N_11544,N_11416,N_11408);
or U11545 (N_11545,N_11506,N_11502);
nor U11546 (N_11546,N_11367,N_11426);
xnor U11547 (N_11547,N_11428,N_11433);
and U11548 (N_11548,N_11500,N_11418);
or U11549 (N_11549,N_11411,N_11439);
or U11550 (N_11550,N_11517,N_11452);
and U11551 (N_11551,N_11440,N_11448);
xor U11552 (N_11552,N_11490,N_11424);
and U11553 (N_11553,N_11419,N_11396);
nand U11554 (N_11554,N_11470,N_11384);
and U11555 (N_11555,N_11459,N_11458);
nor U11556 (N_11556,N_11497,N_11378);
and U11557 (N_11557,N_11436,N_11509);
and U11558 (N_11558,N_11464,N_11446);
xnor U11559 (N_11559,N_11484,N_11466);
or U11560 (N_11560,N_11389,N_11455);
or U11561 (N_11561,N_11505,N_11451);
or U11562 (N_11562,N_11437,N_11421);
and U11563 (N_11563,N_11480,N_11364);
and U11564 (N_11564,N_11373,N_11415);
and U11565 (N_11565,N_11449,N_11392);
xnor U11566 (N_11566,N_11438,N_11381);
xor U11567 (N_11567,N_11514,N_11410);
xor U11568 (N_11568,N_11362,N_11376);
or U11569 (N_11569,N_11465,N_11432);
or U11570 (N_11570,N_11403,N_11454);
xnor U11571 (N_11571,N_11481,N_11417);
or U11572 (N_11572,N_11372,N_11510);
nor U11573 (N_11573,N_11453,N_11379);
nand U11574 (N_11574,N_11474,N_11445);
nor U11575 (N_11575,N_11414,N_11483);
nand U11576 (N_11576,N_11404,N_11361);
and U11577 (N_11577,N_11390,N_11515);
nor U11578 (N_11578,N_11406,N_11498);
xor U11579 (N_11579,N_11425,N_11479);
xnor U11580 (N_11580,N_11508,N_11518);
or U11581 (N_11581,N_11387,N_11492);
nor U11582 (N_11582,N_11434,N_11487);
xor U11583 (N_11583,N_11369,N_11495);
nand U11584 (N_11584,N_11489,N_11435);
nand U11585 (N_11585,N_11391,N_11471);
and U11586 (N_11586,N_11482,N_11413);
xnor U11587 (N_11587,N_11485,N_11477);
and U11588 (N_11588,N_11503,N_11394);
and U11589 (N_11589,N_11450,N_11405);
or U11590 (N_11590,N_11397,N_11512);
xnor U11591 (N_11591,N_11443,N_11488);
and U11592 (N_11592,N_11422,N_11467);
nor U11593 (N_11593,N_11393,N_11511);
nand U11594 (N_11594,N_11460,N_11382);
nand U11595 (N_11595,N_11395,N_11461);
and U11596 (N_11596,N_11398,N_11399);
nand U11597 (N_11597,N_11444,N_11374);
nor U11598 (N_11598,N_11457,N_11496);
nand U11599 (N_11599,N_11400,N_11494);
nor U11600 (N_11600,N_11435,N_11451);
and U11601 (N_11601,N_11420,N_11436);
nand U11602 (N_11602,N_11426,N_11509);
nand U11603 (N_11603,N_11374,N_11362);
nor U11604 (N_11604,N_11389,N_11500);
xnor U11605 (N_11605,N_11374,N_11454);
nor U11606 (N_11606,N_11367,N_11483);
and U11607 (N_11607,N_11508,N_11388);
nand U11608 (N_11608,N_11484,N_11467);
and U11609 (N_11609,N_11406,N_11510);
nor U11610 (N_11610,N_11373,N_11449);
or U11611 (N_11611,N_11372,N_11366);
nand U11612 (N_11612,N_11509,N_11469);
or U11613 (N_11613,N_11393,N_11481);
nor U11614 (N_11614,N_11390,N_11379);
xnor U11615 (N_11615,N_11455,N_11414);
nor U11616 (N_11616,N_11389,N_11452);
xnor U11617 (N_11617,N_11373,N_11471);
and U11618 (N_11618,N_11456,N_11411);
or U11619 (N_11619,N_11495,N_11399);
nand U11620 (N_11620,N_11506,N_11481);
and U11621 (N_11621,N_11497,N_11436);
and U11622 (N_11622,N_11374,N_11503);
or U11623 (N_11623,N_11451,N_11464);
xor U11624 (N_11624,N_11419,N_11401);
and U11625 (N_11625,N_11434,N_11443);
nor U11626 (N_11626,N_11408,N_11383);
nand U11627 (N_11627,N_11390,N_11360);
nor U11628 (N_11628,N_11408,N_11460);
and U11629 (N_11629,N_11375,N_11512);
xnor U11630 (N_11630,N_11446,N_11430);
nor U11631 (N_11631,N_11401,N_11453);
nor U11632 (N_11632,N_11512,N_11362);
xnor U11633 (N_11633,N_11403,N_11367);
nand U11634 (N_11634,N_11485,N_11518);
xor U11635 (N_11635,N_11394,N_11418);
xor U11636 (N_11636,N_11424,N_11476);
xor U11637 (N_11637,N_11440,N_11361);
nand U11638 (N_11638,N_11508,N_11450);
xnor U11639 (N_11639,N_11510,N_11363);
and U11640 (N_11640,N_11482,N_11372);
or U11641 (N_11641,N_11432,N_11499);
xor U11642 (N_11642,N_11502,N_11430);
nand U11643 (N_11643,N_11439,N_11451);
xnor U11644 (N_11644,N_11430,N_11450);
nand U11645 (N_11645,N_11464,N_11483);
or U11646 (N_11646,N_11378,N_11494);
xor U11647 (N_11647,N_11398,N_11518);
nor U11648 (N_11648,N_11463,N_11427);
nand U11649 (N_11649,N_11373,N_11495);
nand U11650 (N_11650,N_11467,N_11510);
nand U11651 (N_11651,N_11386,N_11371);
nand U11652 (N_11652,N_11517,N_11433);
or U11653 (N_11653,N_11415,N_11480);
nor U11654 (N_11654,N_11430,N_11485);
and U11655 (N_11655,N_11420,N_11409);
nor U11656 (N_11656,N_11458,N_11497);
xor U11657 (N_11657,N_11461,N_11517);
nand U11658 (N_11658,N_11484,N_11380);
nor U11659 (N_11659,N_11452,N_11459);
nor U11660 (N_11660,N_11375,N_11455);
and U11661 (N_11661,N_11506,N_11465);
xnor U11662 (N_11662,N_11500,N_11468);
or U11663 (N_11663,N_11419,N_11365);
nand U11664 (N_11664,N_11406,N_11400);
or U11665 (N_11665,N_11375,N_11377);
xor U11666 (N_11666,N_11406,N_11392);
or U11667 (N_11667,N_11360,N_11370);
nor U11668 (N_11668,N_11508,N_11436);
xnor U11669 (N_11669,N_11478,N_11491);
or U11670 (N_11670,N_11519,N_11518);
or U11671 (N_11671,N_11410,N_11512);
xnor U11672 (N_11672,N_11382,N_11458);
nor U11673 (N_11673,N_11364,N_11406);
or U11674 (N_11674,N_11373,N_11394);
nand U11675 (N_11675,N_11420,N_11393);
xnor U11676 (N_11676,N_11503,N_11502);
nand U11677 (N_11677,N_11443,N_11517);
nand U11678 (N_11678,N_11374,N_11414);
and U11679 (N_11679,N_11429,N_11366);
and U11680 (N_11680,N_11548,N_11541);
or U11681 (N_11681,N_11653,N_11660);
and U11682 (N_11682,N_11639,N_11624);
xnor U11683 (N_11683,N_11600,N_11599);
and U11684 (N_11684,N_11606,N_11674);
nand U11685 (N_11685,N_11554,N_11588);
or U11686 (N_11686,N_11623,N_11612);
or U11687 (N_11687,N_11520,N_11627);
and U11688 (N_11688,N_11549,N_11531);
and U11689 (N_11689,N_11592,N_11577);
nand U11690 (N_11690,N_11540,N_11539);
nor U11691 (N_11691,N_11630,N_11525);
xnor U11692 (N_11692,N_11656,N_11560);
xor U11693 (N_11693,N_11602,N_11594);
and U11694 (N_11694,N_11526,N_11565);
nand U11695 (N_11695,N_11557,N_11537);
xnor U11696 (N_11696,N_11619,N_11590);
and U11697 (N_11697,N_11665,N_11614);
and U11698 (N_11698,N_11637,N_11533);
or U11699 (N_11699,N_11673,N_11626);
and U11700 (N_11700,N_11532,N_11561);
xnor U11701 (N_11701,N_11555,N_11635);
or U11702 (N_11702,N_11567,N_11649);
nor U11703 (N_11703,N_11579,N_11569);
nand U11704 (N_11704,N_11542,N_11631);
xor U11705 (N_11705,N_11593,N_11644);
nor U11706 (N_11706,N_11607,N_11667);
and U11707 (N_11707,N_11574,N_11583);
nand U11708 (N_11708,N_11617,N_11530);
and U11709 (N_11709,N_11563,N_11662);
nand U11710 (N_11710,N_11605,N_11632);
nand U11711 (N_11711,N_11647,N_11650);
xor U11712 (N_11712,N_11634,N_11556);
and U11713 (N_11713,N_11578,N_11595);
nor U11714 (N_11714,N_11638,N_11678);
xnor U11715 (N_11715,N_11589,N_11559);
and U11716 (N_11716,N_11604,N_11669);
and U11717 (N_11717,N_11545,N_11566);
xor U11718 (N_11718,N_11581,N_11544);
nand U11719 (N_11719,N_11571,N_11645);
nand U11720 (N_11720,N_11622,N_11524);
xor U11721 (N_11721,N_11663,N_11664);
and U11722 (N_11722,N_11679,N_11633);
nand U11723 (N_11723,N_11528,N_11616);
or U11724 (N_11724,N_11553,N_11584);
nand U11725 (N_11725,N_11675,N_11640);
and U11726 (N_11726,N_11642,N_11575);
nor U11727 (N_11727,N_11534,N_11618);
and U11728 (N_11728,N_11547,N_11576);
nor U11729 (N_11729,N_11676,N_11641);
or U11730 (N_11730,N_11543,N_11671);
or U11731 (N_11731,N_11587,N_11643);
xor U11732 (N_11732,N_11573,N_11562);
xor U11733 (N_11733,N_11611,N_11629);
nor U11734 (N_11734,N_11636,N_11648);
or U11735 (N_11735,N_11628,N_11523);
nor U11736 (N_11736,N_11677,N_11522);
xnor U11737 (N_11737,N_11657,N_11598);
or U11738 (N_11738,N_11597,N_11596);
nor U11739 (N_11739,N_11527,N_11655);
and U11740 (N_11740,N_11558,N_11568);
nor U11741 (N_11741,N_11625,N_11654);
nand U11742 (N_11742,N_11550,N_11538);
or U11743 (N_11743,N_11582,N_11646);
and U11744 (N_11744,N_11651,N_11570);
xnor U11745 (N_11745,N_11536,N_11615);
nand U11746 (N_11746,N_11603,N_11610);
xor U11747 (N_11747,N_11552,N_11586);
nor U11748 (N_11748,N_11564,N_11585);
nor U11749 (N_11749,N_11580,N_11652);
and U11750 (N_11750,N_11620,N_11551);
xor U11751 (N_11751,N_11546,N_11672);
xor U11752 (N_11752,N_11608,N_11613);
nand U11753 (N_11753,N_11661,N_11659);
xor U11754 (N_11754,N_11521,N_11572);
nor U11755 (N_11755,N_11670,N_11666);
nand U11756 (N_11756,N_11529,N_11621);
or U11757 (N_11757,N_11601,N_11609);
xor U11758 (N_11758,N_11668,N_11535);
and U11759 (N_11759,N_11658,N_11591);
nand U11760 (N_11760,N_11630,N_11663);
or U11761 (N_11761,N_11543,N_11523);
and U11762 (N_11762,N_11521,N_11573);
or U11763 (N_11763,N_11669,N_11670);
and U11764 (N_11764,N_11593,N_11522);
or U11765 (N_11765,N_11530,N_11621);
or U11766 (N_11766,N_11617,N_11607);
and U11767 (N_11767,N_11575,N_11653);
or U11768 (N_11768,N_11679,N_11628);
xnor U11769 (N_11769,N_11618,N_11569);
nand U11770 (N_11770,N_11521,N_11587);
nor U11771 (N_11771,N_11529,N_11617);
nor U11772 (N_11772,N_11537,N_11646);
nand U11773 (N_11773,N_11606,N_11615);
xor U11774 (N_11774,N_11617,N_11545);
and U11775 (N_11775,N_11587,N_11639);
nor U11776 (N_11776,N_11663,N_11679);
nand U11777 (N_11777,N_11545,N_11669);
and U11778 (N_11778,N_11581,N_11535);
and U11779 (N_11779,N_11575,N_11544);
nand U11780 (N_11780,N_11600,N_11549);
xnor U11781 (N_11781,N_11566,N_11547);
nand U11782 (N_11782,N_11522,N_11595);
nor U11783 (N_11783,N_11602,N_11656);
nand U11784 (N_11784,N_11666,N_11587);
or U11785 (N_11785,N_11533,N_11662);
or U11786 (N_11786,N_11557,N_11564);
and U11787 (N_11787,N_11660,N_11566);
and U11788 (N_11788,N_11564,N_11595);
nand U11789 (N_11789,N_11650,N_11593);
or U11790 (N_11790,N_11676,N_11617);
or U11791 (N_11791,N_11532,N_11574);
nor U11792 (N_11792,N_11541,N_11560);
xor U11793 (N_11793,N_11582,N_11533);
nor U11794 (N_11794,N_11541,N_11671);
or U11795 (N_11795,N_11619,N_11585);
and U11796 (N_11796,N_11565,N_11563);
or U11797 (N_11797,N_11609,N_11524);
nand U11798 (N_11798,N_11660,N_11632);
and U11799 (N_11799,N_11579,N_11575);
and U11800 (N_11800,N_11527,N_11638);
xnor U11801 (N_11801,N_11638,N_11561);
nor U11802 (N_11802,N_11610,N_11599);
or U11803 (N_11803,N_11601,N_11665);
nor U11804 (N_11804,N_11643,N_11575);
or U11805 (N_11805,N_11658,N_11594);
and U11806 (N_11806,N_11622,N_11664);
and U11807 (N_11807,N_11674,N_11603);
nor U11808 (N_11808,N_11530,N_11610);
xnor U11809 (N_11809,N_11579,N_11649);
nand U11810 (N_11810,N_11520,N_11668);
xor U11811 (N_11811,N_11628,N_11549);
and U11812 (N_11812,N_11622,N_11653);
and U11813 (N_11813,N_11638,N_11547);
nor U11814 (N_11814,N_11544,N_11550);
xor U11815 (N_11815,N_11560,N_11628);
and U11816 (N_11816,N_11611,N_11526);
or U11817 (N_11817,N_11621,N_11574);
nor U11818 (N_11818,N_11619,N_11520);
and U11819 (N_11819,N_11629,N_11564);
xor U11820 (N_11820,N_11678,N_11600);
and U11821 (N_11821,N_11604,N_11529);
xor U11822 (N_11822,N_11660,N_11673);
nand U11823 (N_11823,N_11576,N_11562);
and U11824 (N_11824,N_11638,N_11670);
nor U11825 (N_11825,N_11672,N_11676);
or U11826 (N_11826,N_11559,N_11526);
and U11827 (N_11827,N_11649,N_11597);
nor U11828 (N_11828,N_11653,N_11630);
nand U11829 (N_11829,N_11559,N_11597);
or U11830 (N_11830,N_11627,N_11565);
nor U11831 (N_11831,N_11629,N_11671);
or U11832 (N_11832,N_11617,N_11652);
and U11833 (N_11833,N_11578,N_11541);
xnor U11834 (N_11834,N_11540,N_11572);
or U11835 (N_11835,N_11578,N_11587);
and U11836 (N_11836,N_11632,N_11671);
nand U11837 (N_11837,N_11591,N_11530);
nand U11838 (N_11838,N_11567,N_11573);
nor U11839 (N_11839,N_11611,N_11542);
or U11840 (N_11840,N_11728,N_11784);
or U11841 (N_11841,N_11839,N_11816);
xor U11842 (N_11842,N_11808,N_11782);
or U11843 (N_11843,N_11701,N_11739);
nor U11844 (N_11844,N_11780,N_11813);
and U11845 (N_11845,N_11700,N_11748);
xor U11846 (N_11846,N_11747,N_11705);
and U11847 (N_11847,N_11802,N_11697);
and U11848 (N_11848,N_11837,N_11758);
nand U11849 (N_11849,N_11717,N_11795);
or U11850 (N_11850,N_11726,N_11734);
or U11851 (N_11851,N_11722,N_11754);
or U11852 (N_11852,N_11715,N_11681);
or U11853 (N_11853,N_11742,N_11755);
or U11854 (N_11854,N_11823,N_11828);
xnor U11855 (N_11855,N_11835,N_11720);
nor U11856 (N_11856,N_11829,N_11767);
nor U11857 (N_11857,N_11769,N_11692);
and U11858 (N_11858,N_11749,N_11800);
nor U11859 (N_11859,N_11759,N_11727);
or U11860 (N_11860,N_11792,N_11736);
and U11861 (N_11861,N_11833,N_11811);
xnor U11862 (N_11862,N_11830,N_11744);
or U11863 (N_11863,N_11689,N_11826);
or U11864 (N_11864,N_11824,N_11738);
xor U11865 (N_11865,N_11791,N_11695);
and U11866 (N_11866,N_11714,N_11818);
and U11867 (N_11867,N_11756,N_11690);
nand U11868 (N_11868,N_11694,N_11702);
nor U11869 (N_11869,N_11757,N_11729);
and U11870 (N_11870,N_11821,N_11741);
or U11871 (N_11871,N_11730,N_11682);
nor U11872 (N_11872,N_11737,N_11834);
and U11873 (N_11873,N_11781,N_11685);
nand U11874 (N_11874,N_11760,N_11819);
and U11875 (N_11875,N_11735,N_11723);
and U11876 (N_11876,N_11787,N_11790);
nor U11877 (N_11877,N_11761,N_11680);
xnor U11878 (N_11878,N_11832,N_11794);
nand U11879 (N_11879,N_11820,N_11838);
nand U11880 (N_11880,N_11712,N_11778);
nand U11881 (N_11881,N_11716,N_11807);
or U11882 (N_11882,N_11711,N_11733);
nand U11883 (N_11883,N_11703,N_11724);
or U11884 (N_11884,N_11793,N_11709);
and U11885 (N_11885,N_11698,N_11772);
xnor U11886 (N_11886,N_11810,N_11718);
xnor U11887 (N_11887,N_11693,N_11688);
xor U11888 (N_11888,N_11777,N_11801);
and U11889 (N_11889,N_11708,N_11684);
nand U11890 (N_11890,N_11836,N_11768);
and U11891 (N_11891,N_11732,N_11827);
nand U11892 (N_11892,N_11797,N_11746);
nor U11893 (N_11893,N_11773,N_11799);
nand U11894 (N_11894,N_11707,N_11770);
or U11895 (N_11895,N_11783,N_11805);
and U11896 (N_11896,N_11696,N_11779);
and U11897 (N_11897,N_11763,N_11753);
nor U11898 (N_11898,N_11774,N_11804);
xnor U11899 (N_11899,N_11691,N_11752);
nand U11900 (N_11900,N_11817,N_11785);
nor U11901 (N_11901,N_11798,N_11683);
or U11902 (N_11902,N_11721,N_11825);
xor U11903 (N_11903,N_11751,N_11765);
and U11904 (N_11904,N_11740,N_11812);
nor U11905 (N_11905,N_11766,N_11786);
nand U11906 (N_11906,N_11719,N_11762);
and U11907 (N_11907,N_11789,N_11725);
or U11908 (N_11908,N_11788,N_11699);
and U11909 (N_11909,N_11806,N_11776);
nand U11910 (N_11910,N_11775,N_11814);
and U11911 (N_11911,N_11743,N_11796);
and U11912 (N_11912,N_11731,N_11809);
or U11913 (N_11913,N_11771,N_11686);
or U11914 (N_11914,N_11706,N_11713);
xor U11915 (N_11915,N_11704,N_11710);
nand U11916 (N_11916,N_11750,N_11764);
xor U11917 (N_11917,N_11745,N_11815);
nor U11918 (N_11918,N_11822,N_11803);
nand U11919 (N_11919,N_11831,N_11687);
or U11920 (N_11920,N_11744,N_11805);
nand U11921 (N_11921,N_11733,N_11695);
xor U11922 (N_11922,N_11754,N_11788);
nor U11923 (N_11923,N_11759,N_11705);
xor U11924 (N_11924,N_11696,N_11747);
xnor U11925 (N_11925,N_11710,N_11753);
or U11926 (N_11926,N_11780,N_11808);
nand U11927 (N_11927,N_11738,N_11756);
nor U11928 (N_11928,N_11712,N_11764);
xor U11929 (N_11929,N_11778,N_11707);
xor U11930 (N_11930,N_11710,N_11751);
nor U11931 (N_11931,N_11714,N_11771);
xnor U11932 (N_11932,N_11756,N_11732);
and U11933 (N_11933,N_11777,N_11705);
nand U11934 (N_11934,N_11706,N_11805);
xnor U11935 (N_11935,N_11814,N_11835);
nand U11936 (N_11936,N_11710,N_11722);
nor U11937 (N_11937,N_11790,N_11680);
xnor U11938 (N_11938,N_11778,N_11736);
nand U11939 (N_11939,N_11785,N_11839);
xor U11940 (N_11940,N_11680,N_11737);
or U11941 (N_11941,N_11758,N_11757);
nor U11942 (N_11942,N_11692,N_11827);
xor U11943 (N_11943,N_11683,N_11782);
xor U11944 (N_11944,N_11803,N_11808);
or U11945 (N_11945,N_11799,N_11833);
xnor U11946 (N_11946,N_11766,N_11742);
or U11947 (N_11947,N_11686,N_11813);
nand U11948 (N_11948,N_11787,N_11767);
or U11949 (N_11949,N_11733,N_11792);
and U11950 (N_11950,N_11739,N_11709);
or U11951 (N_11951,N_11759,N_11684);
nor U11952 (N_11952,N_11776,N_11756);
nor U11953 (N_11953,N_11776,N_11814);
or U11954 (N_11954,N_11734,N_11787);
or U11955 (N_11955,N_11681,N_11794);
nand U11956 (N_11956,N_11826,N_11806);
or U11957 (N_11957,N_11733,N_11707);
nand U11958 (N_11958,N_11723,N_11769);
nand U11959 (N_11959,N_11813,N_11764);
xor U11960 (N_11960,N_11779,N_11717);
nand U11961 (N_11961,N_11814,N_11737);
xnor U11962 (N_11962,N_11681,N_11780);
nand U11963 (N_11963,N_11709,N_11719);
and U11964 (N_11964,N_11706,N_11703);
and U11965 (N_11965,N_11747,N_11836);
xor U11966 (N_11966,N_11778,N_11749);
nor U11967 (N_11967,N_11811,N_11710);
and U11968 (N_11968,N_11731,N_11838);
or U11969 (N_11969,N_11705,N_11707);
or U11970 (N_11970,N_11717,N_11740);
xnor U11971 (N_11971,N_11789,N_11697);
or U11972 (N_11972,N_11683,N_11719);
nor U11973 (N_11973,N_11688,N_11822);
xnor U11974 (N_11974,N_11737,N_11733);
nor U11975 (N_11975,N_11695,N_11779);
nand U11976 (N_11976,N_11774,N_11806);
xnor U11977 (N_11977,N_11776,N_11749);
and U11978 (N_11978,N_11720,N_11738);
nor U11979 (N_11979,N_11787,N_11707);
nand U11980 (N_11980,N_11705,N_11735);
xor U11981 (N_11981,N_11753,N_11831);
nor U11982 (N_11982,N_11726,N_11753);
nand U11983 (N_11983,N_11833,N_11705);
xnor U11984 (N_11984,N_11716,N_11818);
xor U11985 (N_11985,N_11786,N_11698);
nor U11986 (N_11986,N_11713,N_11725);
nor U11987 (N_11987,N_11778,N_11696);
or U11988 (N_11988,N_11796,N_11834);
and U11989 (N_11989,N_11740,N_11795);
nand U11990 (N_11990,N_11755,N_11723);
nand U11991 (N_11991,N_11823,N_11818);
or U11992 (N_11992,N_11837,N_11790);
nand U11993 (N_11993,N_11808,N_11771);
and U11994 (N_11994,N_11683,N_11794);
nor U11995 (N_11995,N_11708,N_11808);
or U11996 (N_11996,N_11819,N_11769);
xor U11997 (N_11997,N_11700,N_11801);
or U11998 (N_11998,N_11819,N_11810);
nor U11999 (N_11999,N_11789,N_11831);
nand U12000 (N_12000,N_11946,N_11901);
and U12001 (N_12001,N_11850,N_11870);
nand U12002 (N_12002,N_11886,N_11900);
nor U12003 (N_12003,N_11883,N_11882);
nand U12004 (N_12004,N_11998,N_11920);
xor U12005 (N_12005,N_11919,N_11983);
and U12006 (N_12006,N_11871,N_11855);
nand U12007 (N_12007,N_11967,N_11931);
or U12008 (N_12008,N_11916,N_11986);
xor U12009 (N_12009,N_11896,N_11852);
nor U12010 (N_12010,N_11941,N_11868);
and U12011 (N_12011,N_11964,N_11980);
nand U12012 (N_12012,N_11911,N_11914);
and U12013 (N_12013,N_11957,N_11926);
or U12014 (N_12014,N_11993,N_11866);
nand U12015 (N_12015,N_11972,N_11862);
nor U12016 (N_12016,N_11930,N_11895);
nand U12017 (N_12017,N_11969,N_11987);
and U12018 (N_12018,N_11859,N_11943);
or U12019 (N_12019,N_11977,N_11939);
nor U12020 (N_12020,N_11922,N_11966);
nor U12021 (N_12021,N_11953,N_11898);
or U12022 (N_12022,N_11867,N_11924);
xor U12023 (N_12023,N_11959,N_11945);
and U12024 (N_12024,N_11944,N_11912);
or U12025 (N_12025,N_11846,N_11872);
or U12026 (N_12026,N_11981,N_11928);
nand U12027 (N_12027,N_11929,N_11947);
nor U12028 (N_12028,N_11950,N_11910);
nor U12029 (N_12029,N_11840,N_11904);
nor U12030 (N_12030,N_11856,N_11954);
and U12031 (N_12031,N_11978,N_11940);
nor U12032 (N_12032,N_11933,N_11937);
and U12033 (N_12033,N_11845,N_11877);
nand U12034 (N_12034,N_11970,N_11995);
xor U12035 (N_12035,N_11951,N_11932);
nor U12036 (N_12036,N_11874,N_11844);
nand U12037 (N_12037,N_11881,N_11992);
xnor U12038 (N_12038,N_11878,N_11893);
or U12039 (N_12039,N_11905,N_11842);
xnor U12040 (N_12040,N_11892,N_11849);
and U12041 (N_12041,N_11889,N_11885);
nor U12042 (N_12042,N_11869,N_11903);
nor U12043 (N_12043,N_11962,N_11949);
nor U12044 (N_12044,N_11884,N_11975);
or U12045 (N_12045,N_11973,N_11974);
or U12046 (N_12046,N_11935,N_11984);
and U12047 (N_12047,N_11907,N_11958);
and U12048 (N_12048,N_11841,N_11913);
or U12049 (N_12049,N_11880,N_11915);
nand U12050 (N_12050,N_11997,N_11938);
nor U12051 (N_12051,N_11876,N_11971);
nand U12052 (N_12052,N_11858,N_11988);
or U12053 (N_12053,N_11965,N_11989);
nor U12054 (N_12054,N_11906,N_11865);
and U12055 (N_12055,N_11860,N_11891);
and U12056 (N_12056,N_11909,N_11934);
nand U12057 (N_12057,N_11985,N_11990);
nand U12058 (N_12058,N_11897,N_11890);
nand U12059 (N_12059,N_11899,N_11925);
nor U12060 (N_12060,N_11908,N_11848);
and U12061 (N_12061,N_11887,N_11982);
or U12062 (N_12062,N_11923,N_11936);
or U12063 (N_12063,N_11927,N_11918);
and U12064 (N_12064,N_11948,N_11994);
or U12065 (N_12065,N_11879,N_11902);
nand U12066 (N_12066,N_11955,N_11979);
xnor U12067 (N_12067,N_11999,N_11873);
or U12068 (N_12068,N_11863,N_11853);
nand U12069 (N_12069,N_11917,N_11847);
nor U12070 (N_12070,N_11843,N_11960);
nand U12071 (N_12071,N_11942,N_11963);
xor U12072 (N_12072,N_11991,N_11952);
nand U12073 (N_12073,N_11888,N_11996);
or U12074 (N_12074,N_11961,N_11921);
nand U12075 (N_12075,N_11956,N_11851);
or U12076 (N_12076,N_11857,N_11875);
or U12077 (N_12077,N_11976,N_11968);
and U12078 (N_12078,N_11894,N_11864);
xnor U12079 (N_12079,N_11861,N_11854);
nor U12080 (N_12080,N_11957,N_11925);
xnor U12081 (N_12081,N_11978,N_11918);
and U12082 (N_12082,N_11902,N_11875);
xor U12083 (N_12083,N_11868,N_11942);
nor U12084 (N_12084,N_11985,N_11886);
nand U12085 (N_12085,N_11907,N_11991);
xnor U12086 (N_12086,N_11991,N_11938);
nor U12087 (N_12087,N_11867,N_11922);
or U12088 (N_12088,N_11992,N_11970);
nor U12089 (N_12089,N_11951,N_11848);
or U12090 (N_12090,N_11987,N_11928);
and U12091 (N_12091,N_11951,N_11918);
and U12092 (N_12092,N_11870,N_11921);
nand U12093 (N_12093,N_11857,N_11960);
and U12094 (N_12094,N_11965,N_11937);
nand U12095 (N_12095,N_11977,N_11980);
nand U12096 (N_12096,N_11934,N_11860);
xor U12097 (N_12097,N_11867,N_11927);
and U12098 (N_12098,N_11881,N_11896);
nand U12099 (N_12099,N_11975,N_11924);
xnor U12100 (N_12100,N_11902,N_11852);
and U12101 (N_12101,N_11841,N_11843);
xnor U12102 (N_12102,N_11847,N_11926);
nor U12103 (N_12103,N_11886,N_11874);
nor U12104 (N_12104,N_11947,N_11907);
nor U12105 (N_12105,N_11997,N_11889);
and U12106 (N_12106,N_11882,N_11923);
xor U12107 (N_12107,N_11886,N_11868);
nor U12108 (N_12108,N_11936,N_11863);
or U12109 (N_12109,N_11855,N_11863);
and U12110 (N_12110,N_11913,N_11860);
and U12111 (N_12111,N_11852,N_11913);
nand U12112 (N_12112,N_11985,N_11898);
and U12113 (N_12113,N_11942,N_11966);
and U12114 (N_12114,N_11941,N_11968);
nor U12115 (N_12115,N_11978,N_11993);
xor U12116 (N_12116,N_11864,N_11970);
and U12117 (N_12117,N_11927,N_11963);
nor U12118 (N_12118,N_11890,N_11996);
or U12119 (N_12119,N_11881,N_11967);
and U12120 (N_12120,N_11888,N_11990);
and U12121 (N_12121,N_11940,N_11880);
nor U12122 (N_12122,N_11853,N_11848);
xor U12123 (N_12123,N_11973,N_11915);
nor U12124 (N_12124,N_11881,N_11856);
xnor U12125 (N_12125,N_11869,N_11902);
nand U12126 (N_12126,N_11955,N_11959);
or U12127 (N_12127,N_11846,N_11858);
and U12128 (N_12128,N_11938,N_11846);
nand U12129 (N_12129,N_11986,N_11950);
nor U12130 (N_12130,N_11862,N_11997);
nor U12131 (N_12131,N_11931,N_11937);
and U12132 (N_12132,N_11998,N_11907);
nand U12133 (N_12133,N_11866,N_11922);
nor U12134 (N_12134,N_11856,N_11974);
or U12135 (N_12135,N_11967,N_11968);
and U12136 (N_12136,N_11884,N_11942);
xor U12137 (N_12137,N_11902,N_11905);
or U12138 (N_12138,N_11920,N_11968);
and U12139 (N_12139,N_11873,N_11983);
and U12140 (N_12140,N_11950,N_11972);
and U12141 (N_12141,N_11922,N_11992);
and U12142 (N_12142,N_11878,N_11902);
and U12143 (N_12143,N_11892,N_11961);
xor U12144 (N_12144,N_11858,N_11951);
nand U12145 (N_12145,N_11952,N_11949);
and U12146 (N_12146,N_11904,N_11923);
and U12147 (N_12147,N_11861,N_11944);
nand U12148 (N_12148,N_11920,N_11996);
nand U12149 (N_12149,N_11876,N_11877);
nand U12150 (N_12150,N_11854,N_11870);
nor U12151 (N_12151,N_11982,N_11877);
nand U12152 (N_12152,N_11958,N_11884);
or U12153 (N_12153,N_11854,N_11868);
xnor U12154 (N_12154,N_11986,N_11943);
or U12155 (N_12155,N_11979,N_11950);
nor U12156 (N_12156,N_11873,N_11937);
xnor U12157 (N_12157,N_11944,N_11960);
or U12158 (N_12158,N_11857,N_11850);
nand U12159 (N_12159,N_11913,N_11909);
nand U12160 (N_12160,N_12044,N_12061);
and U12161 (N_12161,N_12056,N_12013);
nand U12162 (N_12162,N_12120,N_12027);
nand U12163 (N_12163,N_12019,N_12079);
xnor U12164 (N_12164,N_12149,N_12025);
xor U12165 (N_12165,N_12121,N_12026);
or U12166 (N_12166,N_12111,N_12141);
xnor U12167 (N_12167,N_12138,N_12012);
nor U12168 (N_12168,N_12050,N_12046);
xor U12169 (N_12169,N_12131,N_12024);
and U12170 (N_12170,N_12128,N_12101);
nand U12171 (N_12171,N_12070,N_12067);
nor U12172 (N_12172,N_12072,N_12097);
xor U12173 (N_12173,N_12100,N_12035);
xnor U12174 (N_12174,N_12135,N_12126);
and U12175 (N_12175,N_12114,N_12124);
xnor U12176 (N_12176,N_12154,N_12155);
or U12177 (N_12177,N_12021,N_12116);
nand U12178 (N_12178,N_12125,N_12087);
and U12179 (N_12179,N_12069,N_12038);
and U12180 (N_12180,N_12017,N_12142);
or U12181 (N_12181,N_12104,N_12055);
nand U12182 (N_12182,N_12099,N_12049);
or U12183 (N_12183,N_12148,N_12058);
xor U12184 (N_12184,N_12053,N_12068);
nor U12185 (N_12185,N_12051,N_12036);
xnor U12186 (N_12186,N_12113,N_12134);
or U12187 (N_12187,N_12045,N_12062);
nand U12188 (N_12188,N_12086,N_12090);
nand U12189 (N_12189,N_12136,N_12005);
and U12190 (N_12190,N_12004,N_12084);
nand U12191 (N_12191,N_12127,N_12066);
and U12192 (N_12192,N_12144,N_12006);
or U12193 (N_12193,N_12075,N_12054);
or U12194 (N_12194,N_12000,N_12112);
or U12195 (N_12195,N_12096,N_12089);
nor U12196 (N_12196,N_12071,N_12040);
xnor U12197 (N_12197,N_12147,N_12028);
and U12198 (N_12198,N_12042,N_12106);
xor U12199 (N_12199,N_12007,N_12143);
xor U12200 (N_12200,N_12139,N_12151);
nand U12201 (N_12201,N_12020,N_12029);
or U12202 (N_12202,N_12091,N_12016);
nor U12203 (N_12203,N_12060,N_12105);
or U12204 (N_12204,N_12015,N_12085);
xnor U12205 (N_12205,N_12157,N_12150);
or U12206 (N_12206,N_12047,N_12103);
xor U12207 (N_12207,N_12001,N_12115);
or U12208 (N_12208,N_12153,N_12109);
nor U12209 (N_12209,N_12145,N_12059);
or U12210 (N_12210,N_12158,N_12098);
or U12211 (N_12211,N_12014,N_12063);
xnor U12212 (N_12212,N_12009,N_12011);
xor U12213 (N_12213,N_12088,N_12159);
nor U12214 (N_12214,N_12092,N_12082);
nor U12215 (N_12215,N_12152,N_12041);
or U12216 (N_12216,N_12140,N_12094);
nor U12217 (N_12217,N_12093,N_12107);
xnor U12218 (N_12218,N_12123,N_12102);
nor U12219 (N_12219,N_12119,N_12129);
nor U12220 (N_12220,N_12078,N_12037);
xor U12221 (N_12221,N_12034,N_12132);
and U12222 (N_12222,N_12108,N_12039);
xnor U12223 (N_12223,N_12110,N_12023);
xnor U12224 (N_12224,N_12018,N_12076);
xnor U12225 (N_12225,N_12057,N_12032);
nor U12226 (N_12226,N_12065,N_12008);
or U12227 (N_12227,N_12080,N_12010);
or U12228 (N_12228,N_12048,N_12002);
or U12229 (N_12229,N_12130,N_12064);
and U12230 (N_12230,N_12081,N_12003);
xnor U12231 (N_12231,N_12146,N_12022);
nand U12232 (N_12232,N_12095,N_12030);
or U12233 (N_12233,N_12122,N_12074);
nand U12234 (N_12234,N_12073,N_12137);
nand U12235 (N_12235,N_12133,N_12117);
nor U12236 (N_12236,N_12083,N_12052);
nand U12237 (N_12237,N_12118,N_12156);
nand U12238 (N_12238,N_12033,N_12077);
xor U12239 (N_12239,N_12031,N_12043);
and U12240 (N_12240,N_12093,N_12008);
or U12241 (N_12241,N_12119,N_12046);
xnor U12242 (N_12242,N_12095,N_12101);
or U12243 (N_12243,N_12134,N_12056);
nor U12244 (N_12244,N_12063,N_12143);
nand U12245 (N_12245,N_12034,N_12062);
or U12246 (N_12246,N_12009,N_12031);
nor U12247 (N_12247,N_12016,N_12063);
xor U12248 (N_12248,N_12058,N_12064);
and U12249 (N_12249,N_12080,N_12051);
nor U12250 (N_12250,N_12015,N_12125);
or U12251 (N_12251,N_12102,N_12047);
nor U12252 (N_12252,N_12078,N_12027);
nor U12253 (N_12253,N_12158,N_12060);
xor U12254 (N_12254,N_12134,N_12137);
and U12255 (N_12255,N_12014,N_12042);
and U12256 (N_12256,N_12048,N_12028);
xnor U12257 (N_12257,N_12094,N_12042);
and U12258 (N_12258,N_12105,N_12010);
nand U12259 (N_12259,N_12085,N_12077);
nor U12260 (N_12260,N_12031,N_12013);
or U12261 (N_12261,N_12009,N_12020);
xor U12262 (N_12262,N_12145,N_12015);
xor U12263 (N_12263,N_12052,N_12103);
and U12264 (N_12264,N_12088,N_12019);
and U12265 (N_12265,N_12148,N_12082);
nand U12266 (N_12266,N_12099,N_12056);
xor U12267 (N_12267,N_12096,N_12125);
or U12268 (N_12268,N_12153,N_12151);
xor U12269 (N_12269,N_12096,N_12009);
xnor U12270 (N_12270,N_12029,N_12048);
or U12271 (N_12271,N_12098,N_12063);
or U12272 (N_12272,N_12009,N_12024);
xnor U12273 (N_12273,N_12086,N_12069);
nor U12274 (N_12274,N_12008,N_12021);
or U12275 (N_12275,N_12014,N_12152);
or U12276 (N_12276,N_12140,N_12120);
and U12277 (N_12277,N_12058,N_12051);
xnor U12278 (N_12278,N_12022,N_12125);
or U12279 (N_12279,N_12155,N_12121);
nand U12280 (N_12280,N_12143,N_12138);
and U12281 (N_12281,N_12090,N_12080);
xor U12282 (N_12282,N_12050,N_12036);
and U12283 (N_12283,N_12066,N_12018);
and U12284 (N_12284,N_12150,N_12025);
nand U12285 (N_12285,N_12114,N_12039);
nand U12286 (N_12286,N_12060,N_12143);
xor U12287 (N_12287,N_12049,N_12130);
or U12288 (N_12288,N_12047,N_12039);
or U12289 (N_12289,N_12089,N_12112);
and U12290 (N_12290,N_12116,N_12070);
nand U12291 (N_12291,N_12049,N_12034);
nand U12292 (N_12292,N_12061,N_12040);
or U12293 (N_12293,N_12066,N_12022);
xnor U12294 (N_12294,N_12069,N_12091);
nor U12295 (N_12295,N_12035,N_12132);
and U12296 (N_12296,N_12138,N_12127);
nor U12297 (N_12297,N_12097,N_12155);
and U12298 (N_12298,N_12098,N_12050);
nor U12299 (N_12299,N_12024,N_12120);
and U12300 (N_12300,N_12120,N_12148);
and U12301 (N_12301,N_12083,N_12078);
nand U12302 (N_12302,N_12061,N_12020);
xnor U12303 (N_12303,N_12067,N_12017);
or U12304 (N_12304,N_12085,N_12133);
and U12305 (N_12305,N_12096,N_12133);
or U12306 (N_12306,N_12134,N_12154);
nor U12307 (N_12307,N_12125,N_12138);
or U12308 (N_12308,N_12093,N_12142);
xor U12309 (N_12309,N_12065,N_12073);
or U12310 (N_12310,N_12148,N_12025);
or U12311 (N_12311,N_12094,N_12078);
and U12312 (N_12312,N_12031,N_12075);
or U12313 (N_12313,N_12120,N_12022);
xor U12314 (N_12314,N_12093,N_12154);
nor U12315 (N_12315,N_12065,N_12157);
or U12316 (N_12316,N_12106,N_12035);
nor U12317 (N_12317,N_12149,N_12114);
nor U12318 (N_12318,N_12024,N_12026);
nand U12319 (N_12319,N_12011,N_12100);
and U12320 (N_12320,N_12276,N_12234);
and U12321 (N_12321,N_12212,N_12224);
nand U12322 (N_12322,N_12178,N_12239);
and U12323 (N_12323,N_12227,N_12269);
and U12324 (N_12324,N_12197,N_12259);
nor U12325 (N_12325,N_12255,N_12194);
nand U12326 (N_12326,N_12284,N_12294);
and U12327 (N_12327,N_12289,N_12281);
or U12328 (N_12328,N_12202,N_12165);
or U12329 (N_12329,N_12189,N_12176);
and U12330 (N_12330,N_12287,N_12179);
xor U12331 (N_12331,N_12272,N_12282);
and U12332 (N_12332,N_12306,N_12251);
and U12333 (N_12333,N_12244,N_12240);
or U12334 (N_12334,N_12160,N_12229);
nand U12335 (N_12335,N_12270,N_12310);
nor U12336 (N_12336,N_12233,N_12290);
and U12337 (N_12337,N_12182,N_12291);
and U12338 (N_12338,N_12312,N_12236);
nor U12339 (N_12339,N_12273,N_12308);
nor U12340 (N_12340,N_12218,N_12200);
nor U12341 (N_12341,N_12245,N_12219);
nand U12342 (N_12342,N_12199,N_12238);
nor U12343 (N_12343,N_12297,N_12210);
or U12344 (N_12344,N_12173,N_12167);
and U12345 (N_12345,N_12267,N_12293);
and U12346 (N_12346,N_12230,N_12303);
and U12347 (N_12347,N_12296,N_12193);
and U12348 (N_12348,N_12161,N_12265);
nor U12349 (N_12349,N_12249,N_12274);
and U12350 (N_12350,N_12248,N_12184);
xor U12351 (N_12351,N_12307,N_12260);
nor U12352 (N_12352,N_12225,N_12231);
xor U12353 (N_12353,N_12278,N_12207);
or U12354 (N_12354,N_12174,N_12163);
and U12355 (N_12355,N_12209,N_12188);
nor U12356 (N_12356,N_12316,N_12313);
and U12357 (N_12357,N_12166,N_12170);
and U12358 (N_12358,N_12301,N_12319);
or U12359 (N_12359,N_12263,N_12286);
nand U12360 (N_12360,N_12264,N_12277);
xnor U12361 (N_12361,N_12315,N_12211);
nand U12362 (N_12362,N_12217,N_12271);
or U12363 (N_12363,N_12314,N_12206);
and U12364 (N_12364,N_12298,N_12256);
or U12365 (N_12365,N_12223,N_12214);
and U12366 (N_12366,N_12253,N_12257);
xnor U12367 (N_12367,N_12288,N_12164);
nand U12368 (N_12368,N_12262,N_12232);
nor U12369 (N_12369,N_12201,N_12246);
or U12370 (N_12370,N_12190,N_12228);
xnor U12371 (N_12371,N_12241,N_12203);
nand U12372 (N_12372,N_12292,N_12183);
nand U12373 (N_12373,N_12185,N_12213);
nor U12374 (N_12374,N_12235,N_12279);
or U12375 (N_12375,N_12243,N_12247);
nand U12376 (N_12376,N_12226,N_12300);
nor U12377 (N_12377,N_12280,N_12252);
xor U12378 (N_12378,N_12258,N_12198);
or U12379 (N_12379,N_12285,N_12266);
or U12380 (N_12380,N_12309,N_12221);
or U12381 (N_12381,N_12242,N_12204);
xor U12382 (N_12382,N_12250,N_12254);
and U12383 (N_12383,N_12175,N_12196);
xor U12384 (N_12384,N_12311,N_12317);
xnor U12385 (N_12385,N_12318,N_12283);
or U12386 (N_12386,N_12171,N_12177);
nor U12387 (N_12387,N_12208,N_12172);
nand U12388 (N_12388,N_12295,N_12220);
or U12389 (N_12389,N_12299,N_12215);
xnor U12390 (N_12390,N_12216,N_12169);
xor U12391 (N_12391,N_12237,N_12192);
nor U12392 (N_12392,N_12275,N_12305);
or U12393 (N_12393,N_12261,N_12168);
and U12394 (N_12394,N_12186,N_12304);
xor U12395 (N_12395,N_12222,N_12187);
and U12396 (N_12396,N_12181,N_12195);
xnor U12397 (N_12397,N_12191,N_12162);
or U12398 (N_12398,N_12268,N_12205);
and U12399 (N_12399,N_12180,N_12302);
nand U12400 (N_12400,N_12300,N_12173);
and U12401 (N_12401,N_12243,N_12266);
nor U12402 (N_12402,N_12293,N_12160);
and U12403 (N_12403,N_12260,N_12245);
xor U12404 (N_12404,N_12162,N_12223);
or U12405 (N_12405,N_12291,N_12309);
or U12406 (N_12406,N_12178,N_12202);
and U12407 (N_12407,N_12305,N_12171);
or U12408 (N_12408,N_12299,N_12250);
and U12409 (N_12409,N_12242,N_12231);
nor U12410 (N_12410,N_12169,N_12284);
nand U12411 (N_12411,N_12169,N_12192);
nand U12412 (N_12412,N_12315,N_12171);
nand U12413 (N_12413,N_12293,N_12244);
nand U12414 (N_12414,N_12211,N_12277);
or U12415 (N_12415,N_12245,N_12243);
xnor U12416 (N_12416,N_12265,N_12189);
nor U12417 (N_12417,N_12191,N_12238);
nand U12418 (N_12418,N_12212,N_12319);
or U12419 (N_12419,N_12285,N_12298);
nor U12420 (N_12420,N_12171,N_12201);
nor U12421 (N_12421,N_12270,N_12251);
or U12422 (N_12422,N_12198,N_12292);
nand U12423 (N_12423,N_12180,N_12279);
nand U12424 (N_12424,N_12195,N_12228);
nand U12425 (N_12425,N_12193,N_12167);
or U12426 (N_12426,N_12280,N_12315);
and U12427 (N_12427,N_12308,N_12245);
and U12428 (N_12428,N_12292,N_12250);
nor U12429 (N_12429,N_12162,N_12302);
xnor U12430 (N_12430,N_12239,N_12303);
nand U12431 (N_12431,N_12211,N_12160);
and U12432 (N_12432,N_12297,N_12221);
and U12433 (N_12433,N_12188,N_12261);
nor U12434 (N_12434,N_12236,N_12270);
nand U12435 (N_12435,N_12275,N_12272);
xnor U12436 (N_12436,N_12218,N_12237);
nor U12437 (N_12437,N_12191,N_12273);
and U12438 (N_12438,N_12225,N_12261);
nor U12439 (N_12439,N_12253,N_12277);
xor U12440 (N_12440,N_12237,N_12291);
nand U12441 (N_12441,N_12252,N_12262);
nor U12442 (N_12442,N_12248,N_12284);
nand U12443 (N_12443,N_12297,N_12176);
or U12444 (N_12444,N_12215,N_12270);
xor U12445 (N_12445,N_12268,N_12254);
or U12446 (N_12446,N_12289,N_12309);
nand U12447 (N_12447,N_12226,N_12192);
or U12448 (N_12448,N_12299,N_12303);
and U12449 (N_12449,N_12238,N_12313);
xnor U12450 (N_12450,N_12162,N_12206);
and U12451 (N_12451,N_12277,N_12199);
or U12452 (N_12452,N_12211,N_12305);
and U12453 (N_12453,N_12237,N_12210);
xor U12454 (N_12454,N_12205,N_12262);
nand U12455 (N_12455,N_12276,N_12310);
nor U12456 (N_12456,N_12186,N_12169);
and U12457 (N_12457,N_12247,N_12279);
nand U12458 (N_12458,N_12243,N_12251);
and U12459 (N_12459,N_12193,N_12318);
nand U12460 (N_12460,N_12260,N_12199);
xor U12461 (N_12461,N_12215,N_12242);
xor U12462 (N_12462,N_12279,N_12217);
and U12463 (N_12463,N_12214,N_12316);
or U12464 (N_12464,N_12167,N_12273);
xor U12465 (N_12465,N_12209,N_12220);
xor U12466 (N_12466,N_12187,N_12167);
nand U12467 (N_12467,N_12229,N_12219);
nor U12468 (N_12468,N_12297,N_12231);
or U12469 (N_12469,N_12242,N_12246);
or U12470 (N_12470,N_12262,N_12222);
nor U12471 (N_12471,N_12223,N_12308);
and U12472 (N_12472,N_12255,N_12246);
and U12473 (N_12473,N_12213,N_12280);
nor U12474 (N_12474,N_12264,N_12299);
xor U12475 (N_12475,N_12284,N_12230);
nand U12476 (N_12476,N_12166,N_12192);
or U12477 (N_12477,N_12208,N_12293);
nand U12478 (N_12478,N_12173,N_12172);
xor U12479 (N_12479,N_12216,N_12218);
or U12480 (N_12480,N_12425,N_12476);
nor U12481 (N_12481,N_12329,N_12355);
nand U12482 (N_12482,N_12451,N_12336);
nand U12483 (N_12483,N_12434,N_12373);
or U12484 (N_12484,N_12472,N_12369);
xnor U12485 (N_12485,N_12403,N_12432);
or U12486 (N_12486,N_12465,N_12335);
nor U12487 (N_12487,N_12469,N_12364);
nand U12488 (N_12488,N_12352,N_12439);
and U12489 (N_12489,N_12368,N_12407);
xor U12490 (N_12490,N_12383,N_12421);
or U12491 (N_12491,N_12413,N_12365);
nand U12492 (N_12492,N_12477,N_12463);
or U12493 (N_12493,N_12417,N_12321);
or U12494 (N_12494,N_12479,N_12399);
nand U12495 (N_12495,N_12328,N_12366);
or U12496 (N_12496,N_12447,N_12395);
nor U12497 (N_12497,N_12408,N_12378);
or U12498 (N_12498,N_12393,N_12411);
nand U12499 (N_12499,N_12384,N_12330);
nand U12500 (N_12500,N_12431,N_12449);
nor U12501 (N_12501,N_12429,N_12380);
xnor U12502 (N_12502,N_12385,N_12337);
nor U12503 (N_12503,N_12388,N_12333);
xor U12504 (N_12504,N_12339,N_12433);
nor U12505 (N_12505,N_12442,N_12426);
xor U12506 (N_12506,N_12381,N_12400);
nand U12507 (N_12507,N_12418,N_12345);
nor U12508 (N_12508,N_12467,N_12386);
and U12509 (N_12509,N_12455,N_12445);
and U12510 (N_12510,N_12359,N_12406);
xor U12511 (N_12511,N_12446,N_12327);
nor U12512 (N_12512,N_12402,N_12342);
and U12513 (N_12513,N_12340,N_12448);
or U12514 (N_12514,N_12322,N_12438);
nand U12515 (N_12515,N_12414,N_12356);
nor U12516 (N_12516,N_12363,N_12350);
or U12517 (N_12517,N_12344,N_12443);
and U12518 (N_12518,N_12361,N_12351);
nor U12519 (N_12519,N_12412,N_12367);
nand U12520 (N_12520,N_12453,N_12473);
nand U12521 (N_12521,N_12474,N_12401);
xor U12522 (N_12522,N_12362,N_12358);
or U12523 (N_12523,N_12320,N_12441);
nand U12524 (N_12524,N_12440,N_12404);
or U12525 (N_12525,N_12471,N_12454);
nor U12526 (N_12526,N_12452,N_12338);
nor U12527 (N_12527,N_12326,N_12391);
nor U12528 (N_12528,N_12357,N_12475);
and U12529 (N_12529,N_12375,N_12379);
nand U12530 (N_12530,N_12405,N_12334);
nand U12531 (N_12531,N_12466,N_12347);
xnor U12532 (N_12532,N_12464,N_12450);
nand U12533 (N_12533,N_12456,N_12470);
nand U12534 (N_12534,N_12422,N_12360);
nand U12535 (N_12535,N_12461,N_12371);
and U12536 (N_12536,N_12435,N_12420);
nor U12537 (N_12537,N_12382,N_12398);
nor U12538 (N_12538,N_12346,N_12419);
xnor U12539 (N_12539,N_12372,N_12437);
or U12540 (N_12540,N_12377,N_12458);
xnor U12541 (N_12541,N_12331,N_12468);
or U12542 (N_12542,N_12462,N_12416);
and U12543 (N_12543,N_12374,N_12397);
and U12544 (N_12544,N_12376,N_12459);
or U12545 (N_12545,N_12430,N_12424);
or U12546 (N_12546,N_12428,N_12332);
and U12547 (N_12547,N_12478,N_12325);
or U12548 (N_12548,N_12349,N_12324);
nor U12549 (N_12549,N_12354,N_12410);
nand U12550 (N_12550,N_12436,N_12387);
nand U12551 (N_12551,N_12394,N_12343);
nor U12552 (N_12552,N_12423,N_12457);
nor U12553 (N_12553,N_12415,N_12341);
xor U12554 (N_12554,N_12389,N_12392);
nand U12555 (N_12555,N_12396,N_12370);
and U12556 (N_12556,N_12353,N_12409);
or U12557 (N_12557,N_12427,N_12390);
or U12558 (N_12558,N_12460,N_12348);
or U12559 (N_12559,N_12323,N_12444);
nand U12560 (N_12560,N_12394,N_12348);
nand U12561 (N_12561,N_12370,N_12429);
nand U12562 (N_12562,N_12397,N_12393);
or U12563 (N_12563,N_12431,N_12400);
or U12564 (N_12564,N_12321,N_12335);
nand U12565 (N_12565,N_12320,N_12361);
nand U12566 (N_12566,N_12423,N_12439);
nor U12567 (N_12567,N_12457,N_12363);
and U12568 (N_12568,N_12460,N_12370);
or U12569 (N_12569,N_12452,N_12477);
or U12570 (N_12570,N_12379,N_12361);
xnor U12571 (N_12571,N_12404,N_12452);
nor U12572 (N_12572,N_12437,N_12457);
and U12573 (N_12573,N_12420,N_12389);
or U12574 (N_12574,N_12362,N_12332);
nand U12575 (N_12575,N_12350,N_12345);
xor U12576 (N_12576,N_12346,N_12437);
and U12577 (N_12577,N_12331,N_12403);
or U12578 (N_12578,N_12443,N_12390);
nor U12579 (N_12579,N_12458,N_12463);
nand U12580 (N_12580,N_12476,N_12397);
and U12581 (N_12581,N_12400,N_12468);
nand U12582 (N_12582,N_12402,N_12433);
nand U12583 (N_12583,N_12323,N_12414);
xor U12584 (N_12584,N_12417,N_12353);
xnor U12585 (N_12585,N_12450,N_12368);
and U12586 (N_12586,N_12420,N_12371);
xor U12587 (N_12587,N_12431,N_12394);
and U12588 (N_12588,N_12382,N_12407);
nor U12589 (N_12589,N_12430,N_12359);
or U12590 (N_12590,N_12411,N_12374);
nand U12591 (N_12591,N_12426,N_12455);
and U12592 (N_12592,N_12375,N_12479);
nor U12593 (N_12593,N_12433,N_12342);
xnor U12594 (N_12594,N_12354,N_12452);
nor U12595 (N_12595,N_12427,N_12396);
nand U12596 (N_12596,N_12439,N_12479);
nor U12597 (N_12597,N_12466,N_12326);
nor U12598 (N_12598,N_12339,N_12441);
and U12599 (N_12599,N_12436,N_12372);
or U12600 (N_12600,N_12479,N_12400);
nor U12601 (N_12601,N_12475,N_12438);
and U12602 (N_12602,N_12344,N_12404);
and U12603 (N_12603,N_12456,N_12371);
nor U12604 (N_12604,N_12478,N_12352);
xor U12605 (N_12605,N_12474,N_12435);
or U12606 (N_12606,N_12434,N_12439);
xor U12607 (N_12607,N_12423,N_12452);
nor U12608 (N_12608,N_12455,N_12339);
xnor U12609 (N_12609,N_12392,N_12327);
nand U12610 (N_12610,N_12474,N_12470);
xnor U12611 (N_12611,N_12377,N_12331);
or U12612 (N_12612,N_12474,N_12392);
nand U12613 (N_12613,N_12371,N_12388);
and U12614 (N_12614,N_12377,N_12479);
and U12615 (N_12615,N_12468,N_12329);
or U12616 (N_12616,N_12433,N_12338);
nand U12617 (N_12617,N_12457,N_12335);
nand U12618 (N_12618,N_12361,N_12420);
nand U12619 (N_12619,N_12417,N_12385);
and U12620 (N_12620,N_12407,N_12347);
xor U12621 (N_12621,N_12383,N_12428);
xnor U12622 (N_12622,N_12407,N_12367);
nor U12623 (N_12623,N_12368,N_12399);
or U12624 (N_12624,N_12378,N_12465);
nor U12625 (N_12625,N_12392,N_12337);
nor U12626 (N_12626,N_12371,N_12475);
nand U12627 (N_12627,N_12455,N_12367);
and U12628 (N_12628,N_12399,N_12433);
or U12629 (N_12629,N_12473,N_12427);
and U12630 (N_12630,N_12346,N_12368);
and U12631 (N_12631,N_12466,N_12415);
or U12632 (N_12632,N_12323,N_12325);
or U12633 (N_12633,N_12453,N_12332);
xor U12634 (N_12634,N_12373,N_12339);
xnor U12635 (N_12635,N_12393,N_12401);
xnor U12636 (N_12636,N_12328,N_12451);
or U12637 (N_12637,N_12467,N_12325);
and U12638 (N_12638,N_12356,N_12469);
xnor U12639 (N_12639,N_12446,N_12469);
or U12640 (N_12640,N_12541,N_12580);
or U12641 (N_12641,N_12516,N_12510);
nand U12642 (N_12642,N_12635,N_12576);
or U12643 (N_12643,N_12524,N_12486);
nor U12644 (N_12644,N_12592,N_12564);
and U12645 (N_12645,N_12559,N_12613);
nor U12646 (N_12646,N_12591,N_12594);
nor U12647 (N_12647,N_12543,N_12551);
nand U12648 (N_12648,N_12507,N_12546);
nor U12649 (N_12649,N_12518,N_12511);
nand U12650 (N_12650,N_12604,N_12491);
or U12651 (N_12651,N_12545,N_12586);
or U12652 (N_12652,N_12553,N_12584);
or U12653 (N_12653,N_12505,N_12636);
nor U12654 (N_12654,N_12497,N_12630);
or U12655 (N_12655,N_12590,N_12597);
xnor U12656 (N_12656,N_12612,N_12611);
nor U12657 (N_12657,N_12484,N_12629);
nand U12658 (N_12658,N_12632,N_12607);
xor U12659 (N_12659,N_12614,N_12521);
nor U12660 (N_12660,N_12523,N_12485);
or U12661 (N_12661,N_12582,N_12618);
nand U12662 (N_12662,N_12492,N_12487);
and U12663 (N_12663,N_12627,N_12498);
and U12664 (N_12664,N_12619,N_12534);
nor U12665 (N_12665,N_12493,N_12624);
nand U12666 (N_12666,N_12481,N_12608);
and U12667 (N_12667,N_12529,N_12573);
nand U12668 (N_12668,N_12517,N_12552);
xor U12669 (N_12669,N_12620,N_12480);
or U12670 (N_12670,N_12557,N_12500);
nand U12671 (N_12671,N_12528,N_12525);
and U12672 (N_12672,N_12571,N_12526);
xnor U12673 (N_12673,N_12483,N_12502);
nand U12674 (N_12674,N_12555,N_12578);
and U12675 (N_12675,N_12572,N_12574);
nand U12676 (N_12676,N_12522,N_12570);
xor U12677 (N_12677,N_12621,N_12494);
and U12678 (N_12678,N_12554,N_12588);
xor U12679 (N_12679,N_12565,N_12605);
or U12680 (N_12680,N_12514,N_12616);
nor U12681 (N_12681,N_12567,N_12577);
and U12682 (N_12682,N_12598,N_12581);
xnor U12683 (N_12683,N_12499,N_12560);
nor U12684 (N_12684,N_12515,N_12527);
nand U12685 (N_12685,N_12530,N_12503);
and U12686 (N_12686,N_12532,N_12562);
nor U12687 (N_12687,N_12628,N_12549);
or U12688 (N_12688,N_12561,N_12482);
xnor U12689 (N_12689,N_12533,N_12513);
nor U12690 (N_12690,N_12639,N_12575);
nor U12691 (N_12691,N_12539,N_12634);
xnor U12692 (N_12692,N_12495,N_12535);
nand U12693 (N_12693,N_12531,N_12537);
xor U12694 (N_12694,N_12508,N_12544);
nor U12695 (N_12695,N_12593,N_12589);
nand U12696 (N_12696,N_12490,N_12601);
xor U12697 (N_12697,N_12509,N_12548);
or U12698 (N_12698,N_12568,N_12536);
nand U12699 (N_12699,N_12501,N_12606);
or U12700 (N_12700,N_12542,N_12596);
nand U12701 (N_12701,N_12512,N_12504);
and U12702 (N_12702,N_12610,N_12626);
nor U12703 (N_12703,N_12585,N_12550);
or U12704 (N_12704,N_12625,N_12637);
or U12705 (N_12705,N_12633,N_12563);
and U12706 (N_12706,N_12547,N_12595);
nor U12707 (N_12707,N_12623,N_12558);
nor U12708 (N_12708,N_12602,N_12519);
nor U12709 (N_12709,N_12622,N_12540);
nand U12710 (N_12710,N_12600,N_12599);
nand U12711 (N_12711,N_12489,N_12566);
nor U12712 (N_12712,N_12609,N_12506);
nor U12713 (N_12713,N_12520,N_12631);
nand U12714 (N_12714,N_12617,N_12556);
or U12715 (N_12715,N_12587,N_12488);
nor U12716 (N_12716,N_12615,N_12579);
or U12717 (N_12717,N_12638,N_12538);
or U12718 (N_12718,N_12569,N_12496);
xnor U12719 (N_12719,N_12583,N_12603);
nand U12720 (N_12720,N_12591,N_12551);
nor U12721 (N_12721,N_12617,N_12638);
and U12722 (N_12722,N_12539,N_12491);
nor U12723 (N_12723,N_12487,N_12514);
xnor U12724 (N_12724,N_12500,N_12620);
nand U12725 (N_12725,N_12483,N_12579);
nand U12726 (N_12726,N_12556,N_12613);
nor U12727 (N_12727,N_12567,N_12540);
nand U12728 (N_12728,N_12604,N_12513);
or U12729 (N_12729,N_12620,N_12577);
nor U12730 (N_12730,N_12626,N_12611);
xor U12731 (N_12731,N_12572,N_12488);
nand U12732 (N_12732,N_12529,N_12575);
nor U12733 (N_12733,N_12500,N_12516);
nor U12734 (N_12734,N_12595,N_12492);
and U12735 (N_12735,N_12490,N_12547);
and U12736 (N_12736,N_12566,N_12545);
nor U12737 (N_12737,N_12584,N_12493);
and U12738 (N_12738,N_12523,N_12551);
xnor U12739 (N_12739,N_12554,N_12547);
nor U12740 (N_12740,N_12548,N_12573);
and U12741 (N_12741,N_12613,N_12596);
and U12742 (N_12742,N_12543,N_12531);
nor U12743 (N_12743,N_12632,N_12577);
and U12744 (N_12744,N_12527,N_12510);
and U12745 (N_12745,N_12587,N_12578);
xor U12746 (N_12746,N_12630,N_12487);
nor U12747 (N_12747,N_12513,N_12639);
nand U12748 (N_12748,N_12512,N_12574);
nand U12749 (N_12749,N_12491,N_12543);
and U12750 (N_12750,N_12562,N_12601);
and U12751 (N_12751,N_12569,N_12517);
and U12752 (N_12752,N_12604,N_12628);
nand U12753 (N_12753,N_12560,N_12543);
nor U12754 (N_12754,N_12495,N_12620);
or U12755 (N_12755,N_12484,N_12623);
nor U12756 (N_12756,N_12621,N_12543);
and U12757 (N_12757,N_12638,N_12561);
xnor U12758 (N_12758,N_12610,N_12488);
xnor U12759 (N_12759,N_12483,N_12613);
nor U12760 (N_12760,N_12577,N_12627);
or U12761 (N_12761,N_12601,N_12581);
nand U12762 (N_12762,N_12514,N_12527);
xor U12763 (N_12763,N_12523,N_12597);
or U12764 (N_12764,N_12507,N_12630);
nand U12765 (N_12765,N_12532,N_12506);
xor U12766 (N_12766,N_12603,N_12508);
and U12767 (N_12767,N_12579,N_12503);
xor U12768 (N_12768,N_12487,N_12631);
nand U12769 (N_12769,N_12529,N_12604);
or U12770 (N_12770,N_12587,N_12627);
and U12771 (N_12771,N_12480,N_12509);
nand U12772 (N_12772,N_12594,N_12629);
and U12773 (N_12773,N_12587,N_12579);
xnor U12774 (N_12774,N_12513,N_12500);
or U12775 (N_12775,N_12512,N_12578);
nor U12776 (N_12776,N_12588,N_12522);
nor U12777 (N_12777,N_12599,N_12597);
and U12778 (N_12778,N_12499,N_12502);
xnor U12779 (N_12779,N_12609,N_12497);
nor U12780 (N_12780,N_12560,N_12545);
nand U12781 (N_12781,N_12606,N_12521);
and U12782 (N_12782,N_12530,N_12586);
and U12783 (N_12783,N_12591,N_12637);
or U12784 (N_12784,N_12527,N_12632);
or U12785 (N_12785,N_12630,N_12565);
xor U12786 (N_12786,N_12507,N_12555);
nand U12787 (N_12787,N_12500,N_12496);
nand U12788 (N_12788,N_12612,N_12563);
nor U12789 (N_12789,N_12484,N_12599);
nor U12790 (N_12790,N_12616,N_12500);
and U12791 (N_12791,N_12511,N_12606);
and U12792 (N_12792,N_12620,N_12576);
nand U12793 (N_12793,N_12587,N_12534);
or U12794 (N_12794,N_12592,N_12588);
or U12795 (N_12795,N_12565,N_12608);
xnor U12796 (N_12796,N_12578,N_12506);
xnor U12797 (N_12797,N_12607,N_12637);
xor U12798 (N_12798,N_12637,N_12506);
and U12799 (N_12799,N_12502,N_12527);
nand U12800 (N_12800,N_12760,N_12658);
nand U12801 (N_12801,N_12780,N_12688);
or U12802 (N_12802,N_12732,N_12773);
nand U12803 (N_12803,N_12678,N_12708);
nor U12804 (N_12804,N_12738,N_12718);
nor U12805 (N_12805,N_12721,N_12735);
nand U12806 (N_12806,N_12770,N_12743);
xnor U12807 (N_12807,N_12713,N_12795);
nand U12808 (N_12808,N_12691,N_12750);
nor U12809 (N_12809,N_12788,N_12765);
xnor U12810 (N_12810,N_12663,N_12677);
xnor U12811 (N_12811,N_12669,N_12702);
nand U12812 (N_12812,N_12674,N_12671);
nand U12813 (N_12813,N_12796,N_12726);
nor U12814 (N_12814,N_12690,N_12720);
and U12815 (N_12815,N_12781,N_12797);
or U12816 (N_12816,N_12661,N_12745);
xor U12817 (N_12817,N_12689,N_12642);
and U12818 (N_12818,N_12789,N_12649);
nand U12819 (N_12819,N_12653,N_12685);
and U12820 (N_12820,N_12764,N_12662);
xnor U12821 (N_12821,N_12752,N_12709);
nor U12822 (N_12822,N_12654,N_12751);
and U12823 (N_12823,N_12763,N_12737);
and U12824 (N_12824,N_12683,N_12739);
nand U12825 (N_12825,N_12723,N_12651);
or U12826 (N_12826,N_12777,N_12759);
and U12827 (N_12827,N_12657,N_12755);
nand U12828 (N_12828,N_12798,N_12650);
nand U12829 (N_12829,N_12736,N_12730);
nor U12830 (N_12830,N_12676,N_12693);
nor U12831 (N_12831,N_12766,N_12733);
nor U12832 (N_12832,N_12655,N_12784);
nor U12833 (N_12833,N_12734,N_12761);
and U12834 (N_12834,N_12758,N_12717);
nor U12835 (N_12835,N_12722,N_12779);
nor U12836 (N_12836,N_12668,N_12775);
and U12837 (N_12837,N_12731,N_12748);
nor U12838 (N_12838,N_12692,N_12786);
nand U12839 (N_12839,N_12799,N_12645);
or U12840 (N_12840,N_12778,N_12785);
and U12841 (N_12841,N_12646,N_12664);
or U12842 (N_12842,N_12647,N_12719);
and U12843 (N_12843,N_12741,N_12707);
xnor U12844 (N_12844,N_12697,N_12768);
nand U12845 (N_12845,N_12793,N_12675);
xnor U12846 (N_12846,N_12652,N_12641);
nor U12847 (N_12847,N_12791,N_12700);
nor U12848 (N_12848,N_12772,N_12782);
nor U12849 (N_12849,N_12747,N_12680);
xnor U12850 (N_12850,N_12712,N_12746);
xor U12851 (N_12851,N_12753,N_12716);
xnor U12852 (N_12852,N_12749,N_12684);
and U12853 (N_12853,N_12757,N_12769);
nor U12854 (N_12854,N_12698,N_12776);
or U12855 (N_12855,N_12783,N_12771);
nand U12856 (N_12856,N_12670,N_12665);
nor U12857 (N_12857,N_12724,N_12727);
or U12858 (N_12858,N_12767,N_12715);
xor U12859 (N_12859,N_12660,N_12648);
or U12860 (N_12860,N_12666,N_12706);
xnor U12861 (N_12861,N_12711,N_12744);
and U12862 (N_12862,N_12729,N_12754);
xnor U12863 (N_12863,N_12679,N_12714);
xnor U12864 (N_12864,N_12695,N_12725);
nor U12865 (N_12865,N_12686,N_12643);
and U12866 (N_12866,N_12728,N_12703);
or U12867 (N_12867,N_12710,N_12681);
and U12868 (N_12868,N_12696,N_12687);
nand U12869 (N_12869,N_12792,N_12701);
xnor U12870 (N_12870,N_12667,N_12699);
nor U12871 (N_12871,N_12704,N_12740);
xor U12872 (N_12872,N_12640,N_12694);
nand U12873 (N_12873,N_12705,N_12756);
nand U12874 (N_12874,N_12790,N_12742);
xnor U12875 (N_12875,N_12794,N_12673);
nor U12876 (N_12876,N_12774,N_12672);
or U12877 (N_12877,N_12656,N_12644);
and U12878 (N_12878,N_12762,N_12659);
xor U12879 (N_12879,N_12787,N_12682);
nor U12880 (N_12880,N_12727,N_12650);
nand U12881 (N_12881,N_12739,N_12798);
nand U12882 (N_12882,N_12732,N_12710);
nand U12883 (N_12883,N_12795,N_12686);
or U12884 (N_12884,N_12766,N_12735);
and U12885 (N_12885,N_12798,N_12791);
nand U12886 (N_12886,N_12670,N_12698);
xor U12887 (N_12887,N_12773,N_12673);
nor U12888 (N_12888,N_12723,N_12702);
or U12889 (N_12889,N_12751,N_12655);
and U12890 (N_12890,N_12778,N_12743);
nand U12891 (N_12891,N_12741,N_12646);
or U12892 (N_12892,N_12689,N_12766);
or U12893 (N_12893,N_12797,N_12790);
nand U12894 (N_12894,N_12702,N_12653);
or U12895 (N_12895,N_12705,N_12733);
xnor U12896 (N_12896,N_12773,N_12677);
nor U12897 (N_12897,N_12662,N_12714);
nand U12898 (N_12898,N_12658,N_12762);
nand U12899 (N_12899,N_12753,N_12659);
nand U12900 (N_12900,N_12685,N_12672);
or U12901 (N_12901,N_12698,N_12743);
and U12902 (N_12902,N_12685,N_12676);
xnor U12903 (N_12903,N_12776,N_12694);
and U12904 (N_12904,N_12791,N_12783);
and U12905 (N_12905,N_12781,N_12758);
xor U12906 (N_12906,N_12697,N_12710);
nor U12907 (N_12907,N_12775,N_12779);
or U12908 (N_12908,N_12672,N_12735);
nand U12909 (N_12909,N_12656,N_12797);
nand U12910 (N_12910,N_12749,N_12687);
xnor U12911 (N_12911,N_12727,N_12715);
or U12912 (N_12912,N_12714,N_12784);
and U12913 (N_12913,N_12666,N_12652);
nor U12914 (N_12914,N_12737,N_12777);
nor U12915 (N_12915,N_12667,N_12646);
xnor U12916 (N_12916,N_12744,N_12678);
or U12917 (N_12917,N_12761,N_12737);
xnor U12918 (N_12918,N_12673,N_12700);
nand U12919 (N_12919,N_12650,N_12660);
and U12920 (N_12920,N_12732,N_12746);
nand U12921 (N_12921,N_12734,N_12746);
nor U12922 (N_12922,N_12776,N_12702);
nor U12923 (N_12923,N_12743,N_12709);
nand U12924 (N_12924,N_12693,N_12787);
and U12925 (N_12925,N_12644,N_12661);
nor U12926 (N_12926,N_12682,N_12647);
nand U12927 (N_12927,N_12749,N_12663);
and U12928 (N_12928,N_12733,N_12699);
nor U12929 (N_12929,N_12677,N_12754);
or U12930 (N_12930,N_12706,N_12663);
nand U12931 (N_12931,N_12656,N_12673);
and U12932 (N_12932,N_12708,N_12674);
and U12933 (N_12933,N_12784,N_12664);
nor U12934 (N_12934,N_12675,N_12662);
and U12935 (N_12935,N_12731,N_12644);
nand U12936 (N_12936,N_12713,N_12751);
or U12937 (N_12937,N_12739,N_12680);
or U12938 (N_12938,N_12715,N_12743);
and U12939 (N_12939,N_12684,N_12678);
and U12940 (N_12940,N_12743,N_12741);
or U12941 (N_12941,N_12749,N_12747);
and U12942 (N_12942,N_12649,N_12640);
xnor U12943 (N_12943,N_12665,N_12767);
or U12944 (N_12944,N_12651,N_12748);
nand U12945 (N_12945,N_12694,N_12795);
xor U12946 (N_12946,N_12675,N_12709);
xnor U12947 (N_12947,N_12662,N_12713);
nand U12948 (N_12948,N_12743,N_12654);
xnor U12949 (N_12949,N_12717,N_12697);
and U12950 (N_12950,N_12751,N_12729);
nand U12951 (N_12951,N_12707,N_12701);
xnor U12952 (N_12952,N_12648,N_12777);
nor U12953 (N_12953,N_12777,N_12792);
nor U12954 (N_12954,N_12761,N_12683);
xnor U12955 (N_12955,N_12727,N_12771);
nor U12956 (N_12956,N_12669,N_12730);
nor U12957 (N_12957,N_12710,N_12667);
xnor U12958 (N_12958,N_12782,N_12760);
xnor U12959 (N_12959,N_12773,N_12665);
nand U12960 (N_12960,N_12822,N_12917);
nor U12961 (N_12961,N_12861,N_12930);
and U12962 (N_12962,N_12921,N_12910);
and U12963 (N_12963,N_12811,N_12838);
or U12964 (N_12964,N_12867,N_12834);
nand U12965 (N_12965,N_12853,N_12871);
nor U12966 (N_12966,N_12892,N_12901);
xnor U12967 (N_12967,N_12886,N_12957);
nor U12968 (N_12968,N_12854,N_12889);
or U12969 (N_12969,N_12809,N_12878);
or U12970 (N_12970,N_12817,N_12888);
nand U12971 (N_12971,N_12880,N_12879);
or U12972 (N_12972,N_12856,N_12939);
or U12973 (N_12973,N_12909,N_12897);
nand U12974 (N_12974,N_12925,N_12833);
and U12975 (N_12975,N_12802,N_12873);
or U12976 (N_12976,N_12842,N_12936);
and U12977 (N_12977,N_12902,N_12916);
nand U12978 (N_12978,N_12810,N_12850);
xnor U12979 (N_12979,N_12948,N_12928);
nand U12980 (N_12980,N_12815,N_12814);
and U12981 (N_12981,N_12941,N_12821);
nor U12982 (N_12982,N_12929,N_12841);
xnor U12983 (N_12983,N_12887,N_12950);
xor U12984 (N_12984,N_12832,N_12931);
nand U12985 (N_12985,N_12919,N_12884);
nand U12986 (N_12986,N_12857,N_12839);
nand U12987 (N_12987,N_12947,N_12940);
nor U12988 (N_12988,N_12818,N_12900);
xnor U12989 (N_12989,N_12835,N_12837);
xor U12990 (N_12990,N_12846,N_12903);
nor U12991 (N_12991,N_12932,N_12843);
nand U12992 (N_12992,N_12905,N_12907);
xnor U12993 (N_12993,N_12866,N_12920);
nand U12994 (N_12994,N_12825,N_12926);
xnor U12995 (N_12995,N_12849,N_12869);
or U12996 (N_12996,N_12954,N_12912);
nand U12997 (N_12997,N_12938,N_12836);
and U12998 (N_12998,N_12826,N_12956);
or U12999 (N_12999,N_12895,N_12915);
nor U13000 (N_13000,N_12911,N_12891);
or U13001 (N_13001,N_12949,N_12830);
nor U13002 (N_13002,N_12800,N_12819);
or U13003 (N_13003,N_12934,N_12844);
nor U13004 (N_13004,N_12813,N_12862);
and U13005 (N_13005,N_12823,N_12807);
and U13006 (N_13006,N_12847,N_12935);
and U13007 (N_13007,N_12933,N_12872);
nor U13008 (N_13008,N_12904,N_12881);
nor U13009 (N_13009,N_12896,N_12943);
xnor U13010 (N_13010,N_12852,N_12876);
or U13011 (N_13011,N_12840,N_12918);
xor U13012 (N_13012,N_12870,N_12945);
or U13013 (N_13013,N_12828,N_12927);
nor U13014 (N_13014,N_12820,N_12894);
and U13015 (N_13015,N_12882,N_12829);
xor U13016 (N_13016,N_12874,N_12959);
xnor U13017 (N_13017,N_12922,N_12805);
nor U13018 (N_13018,N_12906,N_12937);
nor U13019 (N_13019,N_12944,N_12958);
and U13020 (N_13020,N_12893,N_12923);
nor U13021 (N_13021,N_12899,N_12868);
or U13022 (N_13022,N_12848,N_12855);
or U13023 (N_13023,N_12953,N_12942);
xor U13024 (N_13024,N_12890,N_12875);
nand U13025 (N_13025,N_12951,N_12824);
or U13026 (N_13026,N_12803,N_12806);
xnor U13027 (N_13027,N_12812,N_12908);
nand U13028 (N_13028,N_12883,N_12865);
nor U13029 (N_13029,N_12827,N_12801);
nand U13030 (N_13030,N_12898,N_12831);
xor U13031 (N_13031,N_12808,N_12816);
and U13032 (N_13032,N_12860,N_12877);
and U13033 (N_13033,N_12859,N_12914);
or U13034 (N_13034,N_12952,N_12913);
and U13035 (N_13035,N_12863,N_12851);
nand U13036 (N_13036,N_12858,N_12946);
xnor U13037 (N_13037,N_12864,N_12885);
nand U13038 (N_13038,N_12845,N_12804);
nor U13039 (N_13039,N_12955,N_12924);
and U13040 (N_13040,N_12812,N_12913);
nor U13041 (N_13041,N_12802,N_12894);
nand U13042 (N_13042,N_12936,N_12917);
nor U13043 (N_13043,N_12803,N_12813);
or U13044 (N_13044,N_12910,N_12893);
nor U13045 (N_13045,N_12812,N_12887);
and U13046 (N_13046,N_12823,N_12922);
nor U13047 (N_13047,N_12912,N_12834);
nor U13048 (N_13048,N_12955,N_12933);
xor U13049 (N_13049,N_12870,N_12839);
nand U13050 (N_13050,N_12836,N_12897);
nand U13051 (N_13051,N_12814,N_12892);
nand U13052 (N_13052,N_12909,N_12837);
nand U13053 (N_13053,N_12900,N_12833);
nand U13054 (N_13054,N_12863,N_12957);
nor U13055 (N_13055,N_12813,N_12891);
xnor U13056 (N_13056,N_12880,N_12864);
nand U13057 (N_13057,N_12819,N_12806);
and U13058 (N_13058,N_12899,N_12870);
and U13059 (N_13059,N_12959,N_12830);
nand U13060 (N_13060,N_12841,N_12938);
nand U13061 (N_13061,N_12861,N_12950);
nand U13062 (N_13062,N_12885,N_12887);
or U13063 (N_13063,N_12923,N_12860);
or U13064 (N_13064,N_12806,N_12952);
or U13065 (N_13065,N_12910,N_12800);
nor U13066 (N_13066,N_12921,N_12804);
xor U13067 (N_13067,N_12944,N_12842);
xor U13068 (N_13068,N_12915,N_12812);
and U13069 (N_13069,N_12802,N_12845);
nor U13070 (N_13070,N_12816,N_12862);
nor U13071 (N_13071,N_12958,N_12887);
or U13072 (N_13072,N_12936,N_12825);
nand U13073 (N_13073,N_12811,N_12920);
nand U13074 (N_13074,N_12953,N_12845);
nand U13075 (N_13075,N_12890,N_12880);
xor U13076 (N_13076,N_12829,N_12921);
nor U13077 (N_13077,N_12927,N_12958);
and U13078 (N_13078,N_12820,N_12889);
xor U13079 (N_13079,N_12833,N_12935);
or U13080 (N_13080,N_12801,N_12865);
nor U13081 (N_13081,N_12804,N_12927);
nor U13082 (N_13082,N_12833,N_12920);
nor U13083 (N_13083,N_12808,N_12952);
or U13084 (N_13084,N_12902,N_12914);
nand U13085 (N_13085,N_12869,N_12879);
and U13086 (N_13086,N_12828,N_12918);
nand U13087 (N_13087,N_12930,N_12928);
nor U13088 (N_13088,N_12941,N_12936);
and U13089 (N_13089,N_12898,N_12927);
xor U13090 (N_13090,N_12835,N_12917);
or U13091 (N_13091,N_12863,N_12890);
and U13092 (N_13092,N_12952,N_12908);
or U13093 (N_13093,N_12890,N_12874);
xor U13094 (N_13094,N_12836,N_12803);
nand U13095 (N_13095,N_12849,N_12910);
or U13096 (N_13096,N_12881,N_12889);
xnor U13097 (N_13097,N_12800,N_12909);
xnor U13098 (N_13098,N_12943,N_12893);
or U13099 (N_13099,N_12912,N_12940);
and U13100 (N_13100,N_12807,N_12863);
nand U13101 (N_13101,N_12865,N_12930);
and U13102 (N_13102,N_12831,N_12874);
xor U13103 (N_13103,N_12830,N_12915);
nor U13104 (N_13104,N_12940,N_12883);
xor U13105 (N_13105,N_12914,N_12872);
nor U13106 (N_13106,N_12894,N_12816);
and U13107 (N_13107,N_12875,N_12923);
nor U13108 (N_13108,N_12890,N_12817);
xnor U13109 (N_13109,N_12815,N_12881);
and U13110 (N_13110,N_12807,N_12835);
and U13111 (N_13111,N_12815,N_12884);
and U13112 (N_13112,N_12948,N_12934);
nor U13113 (N_13113,N_12935,N_12884);
or U13114 (N_13114,N_12808,N_12955);
nor U13115 (N_13115,N_12811,N_12959);
and U13116 (N_13116,N_12943,N_12852);
nand U13117 (N_13117,N_12885,N_12936);
nor U13118 (N_13118,N_12837,N_12914);
or U13119 (N_13119,N_12806,N_12863);
xor U13120 (N_13120,N_13046,N_13095);
nand U13121 (N_13121,N_13018,N_12976);
xor U13122 (N_13122,N_12991,N_13073);
nand U13123 (N_13123,N_13034,N_13003);
and U13124 (N_13124,N_12981,N_13047);
or U13125 (N_13125,N_13067,N_13044);
or U13126 (N_13126,N_13086,N_13068);
nand U13127 (N_13127,N_13010,N_13059);
and U13128 (N_13128,N_13006,N_13062);
xor U13129 (N_13129,N_13114,N_13085);
xnor U13130 (N_13130,N_13050,N_13075);
nor U13131 (N_13131,N_12990,N_13007);
xor U13132 (N_13132,N_13101,N_12963);
xnor U13133 (N_13133,N_13109,N_13032);
or U13134 (N_13134,N_12965,N_12970);
nor U13135 (N_13135,N_13113,N_12972);
xor U13136 (N_13136,N_13098,N_13087);
nor U13137 (N_13137,N_13004,N_13096);
xor U13138 (N_13138,N_13091,N_13024);
and U13139 (N_13139,N_12984,N_12993);
or U13140 (N_13140,N_13060,N_12998);
nor U13141 (N_13141,N_13014,N_12961);
or U13142 (N_13142,N_13036,N_12978);
xor U13143 (N_13143,N_13053,N_13015);
nor U13144 (N_13144,N_13037,N_13012);
or U13145 (N_13145,N_12996,N_13117);
and U13146 (N_13146,N_13052,N_13066);
xor U13147 (N_13147,N_13074,N_12980);
nand U13148 (N_13148,N_13033,N_13042);
and U13149 (N_13149,N_13035,N_12986);
and U13150 (N_13150,N_13116,N_13056);
nor U13151 (N_13151,N_13069,N_12977);
nor U13152 (N_13152,N_13118,N_13030);
nand U13153 (N_13153,N_12988,N_13076);
nand U13154 (N_13154,N_12995,N_13013);
xor U13155 (N_13155,N_13102,N_13111);
xor U13156 (N_13156,N_13031,N_12973);
xnor U13157 (N_13157,N_13061,N_13028);
xor U13158 (N_13158,N_12968,N_13005);
and U13159 (N_13159,N_12989,N_13019);
xor U13160 (N_13160,N_13112,N_13088);
nand U13161 (N_13161,N_13039,N_13078);
xor U13162 (N_13162,N_13104,N_13089);
or U13163 (N_13163,N_13016,N_13064);
or U13164 (N_13164,N_13025,N_12966);
or U13165 (N_13165,N_13038,N_13029);
nor U13166 (N_13166,N_13081,N_12997);
nor U13167 (N_13167,N_13103,N_12994);
nor U13168 (N_13168,N_13110,N_13009);
xor U13169 (N_13169,N_13023,N_13020);
nor U13170 (N_13170,N_13000,N_13093);
or U13171 (N_13171,N_13079,N_13107);
and U13172 (N_13172,N_13065,N_13027);
xnor U13173 (N_13173,N_13084,N_13045);
and U13174 (N_13174,N_12982,N_13071);
nand U13175 (N_13175,N_12974,N_13063);
and U13176 (N_13176,N_13090,N_13051);
or U13177 (N_13177,N_12960,N_13058);
nand U13178 (N_13178,N_12969,N_13100);
xnor U13179 (N_13179,N_13070,N_13119);
and U13180 (N_13180,N_13108,N_13055);
nand U13181 (N_13181,N_13097,N_13080);
nor U13182 (N_13182,N_12985,N_13077);
and U13183 (N_13183,N_13040,N_12999);
nor U13184 (N_13184,N_13082,N_12992);
and U13185 (N_13185,N_12967,N_12979);
or U13186 (N_13186,N_13092,N_12987);
or U13187 (N_13187,N_13083,N_12964);
xnor U13188 (N_13188,N_13002,N_13026);
nand U13189 (N_13189,N_13021,N_13106);
xnor U13190 (N_13190,N_12962,N_13001);
and U13191 (N_13191,N_13057,N_12983);
nand U13192 (N_13192,N_13072,N_13008);
or U13193 (N_13193,N_13054,N_13017);
xor U13194 (N_13194,N_13011,N_13099);
nor U13195 (N_13195,N_13094,N_12975);
and U13196 (N_13196,N_13105,N_13115);
xor U13197 (N_13197,N_13048,N_13041);
nand U13198 (N_13198,N_13043,N_12971);
nor U13199 (N_13199,N_13049,N_13022);
nor U13200 (N_13200,N_13092,N_13082);
or U13201 (N_13201,N_13098,N_12966);
and U13202 (N_13202,N_12996,N_12998);
nor U13203 (N_13203,N_13066,N_13023);
nor U13204 (N_13204,N_13069,N_12974);
xnor U13205 (N_13205,N_12961,N_13087);
xor U13206 (N_13206,N_13035,N_12965);
and U13207 (N_13207,N_13038,N_13103);
nand U13208 (N_13208,N_13003,N_12990);
nand U13209 (N_13209,N_13062,N_12960);
nand U13210 (N_13210,N_13026,N_13063);
nor U13211 (N_13211,N_12964,N_12980);
and U13212 (N_13212,N_13022,N_13083);
or U13213 (N_13213,N_13119,N_13015);
xor U13214 (N_13214,N_12960,N_12986);
or U13215 (N_13215,N_13051,N_13076);
and U13216 (N_13216,N_13076,N_13013);
nand U13217 (N_13217,N_13068,N_13091);
or U13218 (N_13218,N_13027,N_13014);
and U13219 (N_13219,N_13042,N_13044);
or U13220 (N_13220,N_13101,N_13010);
or U13221 (N_13221,N_12980,N_12987);
and U13222 (N_13222,N_13031,N_13057);
and U13223 (N_13223,N_13021,N_12963);
nand U13224 (N_13224,N_12970,N_13028);
xnor U13225 (N_13225,N_13063,N_13083);
nor U13226 (N_13226,N_13096,N_12979);
xnor U13227 (N_13227,N_12977,N_13054);
nor U13228 (N_13228,N_13090,N_12979);
xnor U13229 (N_13229,N_12974,N_13016);
or U13230 (N_13230,N_13096,N_13072);
and U13231 (N_13231,N_13062,N_13033);
and U13232 (N_13232,N_13027,N_12978);
nor U13233 (N_13233,N_13108,N_12964);
nand U13234 (N_13234,N_13026,N_13024);
nor U13235 (N_13235,N_13106,N_13016);
nor U13236 (N_13236,N_13084,N_13005);
and U13237 (N_13237,N_13075,N_12984);
xor U13238 (N_13238,N_13028,N_13014);
or U13239 (N_13239,N_13057,N_13056);
xnor U13240 (N_13240,N_13089,N_13096);
and U13241 (N_13241,N_13025,N_13105);
or U13242 (N_13242,N_13011,N_13001);
nand U13243 (N_13243,N_13059,N_13005);
nand U13244 (N_13244,N_12981,N_13076);
or U13245 (N_13245,N_12963,N_13074);
xor U13246 (N_13246,N_13085,N_13099);
or U13247 (N_13247,N_13030,N_13087);
or U13248 (N_13248,N_12965,N_13056);
xor U13249 (N_13249,N_13004,N_12995);
or U13250 (N_13250,N_13112,N_13003);
and U13251 (N_13251,N_13109,N_13063);
or U13252 (N_13252,N_12997,N_13098);
and U13253 (N_13253,N_13096,N_12990);
xor U13254 (N_13254,N_12971,N_12973);
nand U13255 (N_13255,N_12986,N_13045);
or U13256 (N_13256,N_12963,N_13038);
nor U13257 (N_13257,N_13064,N_13066);
or U13258 (N_13258,N_13060,N_13115);
xor U13259 (N_13259,N_12987,N_12979);
or U13260 (N_13260,N_13015,N_12966);
xnor U13261 (N_13261,N_13076,N_13049);
or U13262 (N_13262,N_12980,N_12995);
nor U13263 (N_13263,N_13029,N_13045);
nand U13264 (N_13264,N_13058,N_13114);
or U13265 (N_13265,N_13106,N_13076);
and U13266 (N_13266,N_12974,N_13059);
xnor U13267 (N_13267,N_13054,N_13092);
nor U13268 (N_13268,N_13002,N_12964);
nand U13269 (N_13269,N_13108,N_13084);
xor U13270 (N_13270,N_13111,N_12999);
nand U13271 (N_13271,N_13027,N_13115);
or U13272 (N_13272,N_12979,N_13012);
or U13273 (N_13273,N_12988,N_13000);
nor U13274 (N_13274,N_13048,N_12988);
xnor U13275 (N_13275,N_13005,N_13047);
and U13276 (N_13276,N_13117,N_13045);
or U13277 (N_13277,N_12983,N_12977);
and U13278 (N_13278,N_13061,N_13029);
and U13279 (N_13279,N_13089,N_13037);
and U13280 (N_13280,N_13121,N_13223);
and U13281 (N_13281,N_13210,N_13276);
xor U13282 (N_13282,N_13145,N_13158);
or U13283 (N_13283,N_13209,N_13155);
or U13284 (N_13284,N_13207,N_13161);
nor U13285 (N_13285,N_13228,N_13186);
or U13286 (N_13286,N_13180,N_13165);
and U13287 (N_13287,N_13179,N_13205);
or U13288 (N_13288,N_13224,N_13142);
xnor U13289 (N_13289,N_13256,N_13174);
or U13290 (N_13290,N_13215,N_13201);
or U13291 (N_13291,N_13129,N_13160);
and U13292 (N_13292,N_13131,N_13130);
nand U13293 (N_13293,N_13154,N_13173);
nor U13294 (N_13294,N_13254,N_13136);
nand U13295 (N_13295,N_13237,N_13194);
xor U13296 (N_13296,N_13144,N_13192);
or U13297 (N_13297,N_13200,N_13225);
nor U13298 (N_13298,N_13133,N_13253);
nor U13299 (N_13299,N_13208,N_13218);
nand U13300 (N_13300,N_13272,N_13206);
xor U13301 (N_13301,N_13170,N_13277);
and U13302 (N_13302,N_13127,N_13204);
or U13303 (N_13303,N_13120,N_13214);
or U13304 (N_13304,N_13163,N_13222);
and U13305 (N_13305,N_13134,N_13159);
nand U13306 (N_13306,N_13252,N_13126);
nor U13307 (N_13307,N_13211,N_13122);
xnor U13308 (N_13308,N_13216,N_13274);
nand U13309 (N_13309,N_13229,N_13140);
or U13310 (N_13310,N_13259,N_13148);
nor U13311 (N_13311,N_13188,N_13124);
nor U13312 (N_13312,N_13150,N_13169);
nand U13313 (N_13313,N_13230,N_13191);
nor U13314 (N_13314,N_13238,N_13199);
or U13315 (N_13315,N_13213,N_13242);
and U13316 (N_13316,N_13239,N_13171);
nand U13317 (N_13317,N_13132,N_13181);
or U13318 (N_13318,N_13197,N_13263);
xnor U13319 (N_13319,N_13249,N_13203);
and U13320 (N_13320,N_13260,N_13231);
xor U13321 (N_13321,N_13187,N_13258);
and U13322 (N_13322,N_13196,N_13273);
or U13323 (N_13323,N_13212,N_13241);
and U13324 (N_13324,N_13139,N_13264);
or U13325 (N_13325,N_13275,N_13235);
xor U13326 (N_13326,N_13141,N_13164);
and U13327 (N_13327,N_13146,N_13219);
or U13328 (N_13328,N_13202,N_13243);
and U13329 (N_13329,N_13162,N_13236);
nor U13330 (N_13330,N_13267,N_13250);
nand U13331 (N_13331,N_13177,N_13189);
and U13332 (N_13332,N_13227,N_13278);
or U13333 (N_13333,N_13269,N_13153);
xor U13334 (N_13334,N_13157,N_13247);
nor U13335 (N_13335,N_13175,N_13152);
xor U13336 (N_13336,N_13125,N_13156);
nor U13337 (N_13337,N_13251,N_13268);
xor U13338 (N_13338,N_13172,N_13220);
nor U13339 (N_13339,N_13232,N_13176);
xnor U13340 (N_13340,N_13183,N_13245);
nor U13341 (N_13341,N_13255,N_13217);
or U13342 (N_13342,N_13266,N_13149);
xnor U13343 (N_13343,N_13248,N_13198);
nand U13344 (N_13344,N_13143,N_13167);
nand U13345 (N_13345,N_13184,N_13240);
nor U13346 (N_13346,N_13123,N_13166);
and U13347 (N_13347,N_13182,N_13195);
nor U13348 (N_13348,N_13135,N_13185);
and U13349 (N_13349,N_13168,N_13233);
xor U13350 (N_13350,N_13257,N_13244);
nand U13351 (N_13351,N_13178,N_13234);
nor U13352 (N_13352,N_13190,N_13138);
nor U13353 (N_13353,N_13128,N_13279);
xnor U13354 (N_13354,N_13147,N_13265);
nand U13355 (N_13355,N_13137,N_13221);
nand U13356 (N_13356,N_13246,N_13226);
nor U13357 (N_13357,N_13261,N_13193);
xor U13358 (N_13358,N_13151,N_13270);
nand U13359 (N_13359,N_13262,N_13271);
or U13360 (N_13360,N_13157,N_13208);
or U13361 (N_13361,N_13246,N_13134);
and U13362 (N_13362,N_13255,N_13272);
nor U13363 (N_13363,N_13225,N_13244);
nor U13364 (N_13364,N_13238,N_13208);
xor U13365 (N_13365,N_13142,N_13212);
and U13366 (N_13366,N_13175,N_13214);
nand U13367 (N_13367,N_13248,N_13214);
or U13368 (N_13368,N_13145,N_13134);
and U13369 (N_13369,N_13158,N_13165);
nor U13370 (N_13370,N_13159,N_13245);
nand U13371 (N_13371,N_13179,N_13211);
xor U13372 (N_13372,N_13228,N_13145);
or U13373 (N_13373,N_13239,N_13210);
xor U13374 (N_13374,N_13172,N_13129);
nand U13375 (N_13375,N_13244,N_13240);
xnor U13376 (N_13376,N_13219,N_13247);
and U13377 (N_13377,N_13135,N_13246);
or U13378 (N_13378,N_13271,N_13274);
or U13379 (N_13379,N_13131,N_13198);
or U13380 (N_13380,N_13231,N_13128);
nand U13381 (N_13381,N_13124,N_13274);
nor U13382 (N_13382,N_13175,N_13157);
and U13383 (N_13383,N_13160,N_13174);
nand U13384 (N_13384,N_13255,N_13150);
nand U13385 (N_13385,N_13253,N_13155);
or U13386 (N_13386,N_13220,N_13240);
and U13387 (N_13387,N_13141,N_13216);
nor U13388 (N_13388,N_13234,N_13196);
nor U13389 (N_13389,N_13271,N_13165);
nor U13390 (N_13390,N_13126,N_13216);
nand U13391 (N_13391,N_13244,N_13139);
nand U13392 (N_13392,N_13156,N_13248);
and U13393 (N_13393,N_13200,N_13253);
or U13394 (N_13394,N_13183,N_13133);
nand U13395 (N_13395,N_13132,N_13164);
or U13396 (N_13396,N_13134,N_13176);
and U13397 (N_13397,N_13231,N_13127);
and U13398 (N_13398,N_13193,N_13129);
or U13399 (N_13399,N_13137,N_13266);
nor U13400 (N_13400,N_13235,N_13174);
nor U13401 (N_13401,N_13256,N_13226);
xor U13402 (N_13402,N_13206,N_13212);
nand U13403 (N_13403,N_13123,N_13275);
nor U13404 (N_13404,N_13249,N_13149);
or U13405 (N_13405,N_13170,N_13155);
xnor U13406 (N_13406,N_13222,N_13191);
nor U13407 (N_13407,N_13259,N_13220);
nand U13408 (N_13408,N_13263,N_13159);
xor U13409 (N_13409,N_13172,N_13224);
xor U13410 (N_13410,N_13175,N_13256);
and U13411 (N_13411,N_13162,N_13124);
or U13412 (N_13412,N_13199,N_13259);
nand U13413 (N_13413,N_13263,N_13133);
nand U13414 (N_13414,N_13164,N_13199);
and U13415 (N_13415,N_13121,N_13131);
and U13416 (N_13416,N_13198,N_13138);
xor U13417 (N_13417,N_13245,N_13223);
and U13418 (N_13418,N_13232,N_13278);
xor U13419 (N_13419,N_13275,N_13208);
and U13420 (N_13420,N_13170,N_13211);
nor U13421 (N_13421,N_13212,N_13214);
xor U13422 (N_13422,N_13239,N_13156);
and U13423 (N_13423,N_13259,N_13226);
and U13424 (N_13424,N_13245,N_13132);
or U13425 (N_13425,N_13173,N_13225);
or U13426 (N_13426,N_13181,N_13215);
nand U13427 (N_13427,N_13195,N_13128);
and U13428 (N_13428,N_13268,N_13257);
nand U13429 (N_13429,N_13216,N_13266);
nand U13430 (N_13430,N_13188,N_13240);
nand U13431 (N_13431,N_13131,N_13185);
xnor U13432 (N_13432,N_13254,N_13264);
or U13433 (N_13433,N_13266,N_13136);
xor U13434 (N_13434,N_13179,N_13180);
and U13435 (N_13435,N_13226,N_13278);
xor U13436 (N_13436,N_13187,N_13141);
nor U13437 (N_13437,N_13160,N_13148);
or U13438 (N_13438,N_13199,N_13223);
and U13439 (N_13439,N_13256,N_13263);
and U13440 (N_13440,N_13365,N_13391);
nor U13441 (N_13441,N_13410,N_13420);
nor U13442 (N_13442,N_13293,N_13401);
and U13443 (N_13443,N_13340,N_13439);
or U13444 (N_13444,N_13411,N_13322);
and U13445 (N_13445,N_13357,N_13429);
nand U13446 (N_13446,N_13435,N_13368);
or U13447 (N_13447,N_13416,N_13379);
or U13448 (N_13448,N_13402,N_13407);
nor U13449 (N_13449,N_13290,N_13362);
nor U13450 (N_13450,N_13284,N_13383);
and U13451 (N_13451,N_13343,N_13282);
and U13452 (N_13452,N_13331,N_13397);
nand U13453 (N_13453,N_13395,N_13325);
or U13454 (N_13454,N_13388,N_13366);
and U13455 (N_13455,N_13393,N_13375);
nor U13456 (N_13456,N_13417,N_13430);
or U13457 (N_13457,N_13334,N_13385);
xor U13458 (N_13458,N_13319,N_13310);
xnor U13459 (N_13459,N_13311,N_13419);
and U13460 (N_13460,N_13315,N_13291);
nand U13461 (N_13461,N_13317,N_13288);
and U13462 (N_13462,N_13403,N_13376);
or U13463 (N_13463,N_13352,N_13333);
nand U13464 (N_13464,N_13386,N_13399);
nand U13465 (N_13465,N_13421,N_13327);
xnor U13466 (N_13466,N_13348,N_13381);
xor U13467 (N_13467,N_13301,N_13287);
or U13468 (N_13468,N_13286,N_13387);
nor U13469 (N_13469,N_13423,N_13305);
xnor U13470 (N_13470,N_13338,N_13324);
nor U13471 (N_13471,N_13413,N_13280);
nand U13472 (N_13472,N_13398,N_13296);
nand U13473 (N_13473,N_13426,N_13408);
and U13474 (N_13474,N_13371,N_13400);
nor U13475 (N_13475,N_13339,N_13297);
and U13476 (N_13476,N_13374,N_13309);
xnor U13477 (N_13477,N_13285,N_13303);
nand U13478 (N_13478,N_13369,N_13330);
and U13479 (N_13479,N_13412,N_13431);
and U13480 (N_13480,N_13292,N_13304);
nand U13481 (N_13481,N_13358,N_13359);
nor U13482 (N_13482,N_13406,N_13328);
and U13483 (N_13483,N_13382,N_13326);
and U13484 (N_13484,N_13436,N_13313);
nand U13485 (N_13485,N_13363,N_13329);
nor U13486 (N_13486,N_13380,N_13370);
or U13487 (N_13487,N_13294,N_13356);
or U13488 (N_13488,N_13298,N_13372);
nand U13489 (N_13489,N_13427,N_13378);
nor U13490 (N_13490,N_13355,N_13384);
and U13491 (N_13491,N_13323,N_13433);
or U13492 (N_13492,N_13390,N_13422);
nand U13493 (N_13493,N_13396,N_13364);
nor U13494 (N_13494,N_13418,N_13346);
and U13495 (N_13495,N_13360,N_13361);
nand U13496 (N_13496,N_13354,N_13351);
nand U13497 (N_13497,N_13409,N_13321);
xnor U13498 (N_13498,N_13350,N_13367);
nor U13499 (N_13499,N_13335,N_13300);
nor U13500 (N_13500,N_13405,N_13373);
and U13501 (N_13501,N_13302,N_13306);
and U13502 (N_13502,N_13295,N_13342);
nand U13503 (N_13503,N_13299,N_13404);
nand U13504 (N_13504,N_13320,N_13377);
nand U13505 (N_13505,N_13308,N_13314);
nand U13506 (N_13506,N_13347,N_13414);
nand U13507 (N_13507,N_13289,N_13345);
xnor U13508 (N_13508,N_13316,N_13392);
nand U13509 (N_13509,N_13281,N_13389);
and U13510 (N_13510,N_13341,N_13336);
xnor U13511 (N_13511,N_13428,N_13434);
and U13512 (N_13512,N_13332,N_13424);
and U13513 (N_13513,N_13353,N_13349);
or U13514 (N_13514,N_13337,N_13344);
nor U13515 (N_13515,N_13425,N_13437);
and U13516 (N_13516,N_13394,N_13318);
nor U13517 (N_13517,N_13312,N_13415);
xor U13518 (N_13518,N_13283,N_13432);
or U13519 (N_13519,N_13307,N_13438);
and U13520 (N_13520,N_13284,N_13398);
nand U13521 (N_13521,N_13356,N_13317);
nand U13522 (N_13522,N_13287,N_13396);
nand U13523 (N_13523,N_13363,N_13281);
xnor U13524 (N_13524,N_13385,N_13432);
or U13525 (N_13525,N_13333,N_13424);
or U13526 (N_13526,N_13361,N_13437);
and U13527 (N_13527,N_13303,N_13427);
nor U13528 (N_13528,N_13379,N_13281);
xor U13529 (N_13529,N_13345,N_13288);
nand U13530 (N_13530,N_13343,N_13383);
and U13531 (N_13531,N_13411,N_13396);
or U13532 (N_13532,N_13295,N_13414);
xnor U13533 (N_13533,N_13338,N_13359);
nand U13534 (N_13534,N_13351,N_13355);
nor U13535 (N_13535,N_13422,N_13378);
nand U13536 (N_13536,N_13368,N_13321);
and U13537 (N_13537,N_13285,N_13305);
or U13538 (N_13538,N_13396,N_13302);
and U13539 (N_13539,N_13315,N_13399);
and U13540 (N_13540,N_13310,N_13436);
and U13541 (N_13541,N_13369,N_13421);
xor U13542 (N_13542,N_13282,N_13422);
or U13543 (N_13543,N_13336,N_13340);
and U13544 (N_13544,N_13362,N_13364);
or U13545 (N_13545,N_13406,N_13388);
or U13546 (N_13546,N_13405,N_13314);
xor U13547 (N_13547,N_13363,N_13318);
nand U13548 (N_13548,N_13334,N_13322);
or U13549 (N_13549,N_13336,N_13370);
and U13550 (N_13550,N_13347,N_13384);
and U13551 (N_13551,N_13321,N_13394);
xor U13552 (N_13552,N_13345,N_13410);
and U13553 (N_13553,N_13321,N_13305);
nand U13554 (N_13554,N_13385,N_13402);
nand U13555 (N_13555,N_13351,N_13432);
xor U13556 (N_13556,N_13382,N_13380);
or U13557 (N_13557,N_13346,N_13305);
or U13558 (N_13558,N_13350,N_13291);
nand U13559 (N_13559,N_13282,N_13394);
or U13560 (N_13560,N_13350,N_13380);
xnor U13561 (N_13561,N_13324,N_13287);
nand U13562 (N_13562,N_13325,N_13405);
nor U13563 (N_13563,N_13332,N_13439);
nand U13564 (N_13564,N_13371,N_13327);
and U13565 (N_13565,N_13349,N_13439);
nand U13566 (N_13566,N_13400,N_13366);
and U13567 (N_13567,N_13337,N_13295);
xnor U13568 (N_13568,N_13424,N_13410);
nor U13569 (N_13569,N_13436,N_13425);
nor U13570 (N_13570,N_13379,N_13301);
and U13571 (N_13571,N_13353,N_13427);
and U13572 (N_13572,N_13393,N_13407);
nor U13573 (N_13573,N_13375,N_13340);
nor U13574 (N_13574,N_13324,N_13284);
xnor U13575 (N_13575,N_13362,N_13296);
xor U13576 (N_13576,N_13297,N_13289);
and U13577 (N_13577,N_13366,N_13281);
nand U13578 (N_13578,N_13295,N_13363);
and U13579 (N_13579,N_13349,N_13356);
nor U13580 (N_13580,N_13354,N_13429);
nor U13581 (N_13581,N_13331,N_13282);
and U13582 (N_13582,N_13295,N_13298);
xnor U13583 (N_13583,N_13371,N_13372);
or U13584 (N_13584,N_13288,N_13389);
xnor U13585 (N_13585,N_13353,N_13388);
and U13586 (N_13586,N_13398,N_13374);
nand U13587 (N_13587,N_13430,N_13312);
and U13588 (N_13588,N_13396,N_13408);
nand U13589 (N_13589,N_13369,N_13408);
or U13590 (N_13590,N_13409,N_13354);
xnor U13591 (N_13591,N_13331,N_13309);
and U13592 (N_13592,N_13333,N_13378);
nor U13593 (N_13593,N_13430,N_13393);
xor U13594 (N_13594,N_13433,N_13421);
nand U13595 (N_13595,N_13388,N_13354);
or U13596 (N_13596,N_13306,N_13341);
xnor U13597 (N_13597,N_13408,N_13435);
nor U13598 (N_13598,N_13351,N_13287);
nand U13599 (N_13599,N_13378,N_13375);
nand U13600 (N_13600,N_13591,N_13444);
xor U13601 (N_13601,N_13536,N_13473);
and U13602 (N_13602,N_13488,N_13442);
nor U13603 (N_13603,N_13570,N_13564);
and U13604 (N_13604,N_13453,N_13579);
xor U13605 (N_13605,N_13554,N_13469);
xor U13606 (N_13606,N_13563,N_13542);
xnor U13607 (N_13607,N_13466,N_13578);
xnor U13608 (N_13608,N_13511,N_13477);
nand U13609 (N_13609,N_13472,N_13474);
nor U13610 (N_13610,N_13491,N_13452);
and U13611 (N_13611,N_13520,N_13582);
xnor U13612 (N_13612,N_13565,N_13569);
nand U13613 (N_13613,N_13489,N_13562);
nor U13614 (N_13614,N_13513,N_13599);
and U13615 (N_13615,N_13467,N_13567);
nand U13616 (N_13616,N_13538,N_13456);
or U13617 (N_13617,N_13528,N_13535);
xor U13618 (N_13618,N_13503,N_13481);
or U13619 (N_13619,N_13449,N_13470);
and U13620 (N_13620,N_13446,N_13580);
or U13621 (N_13621,N_13471,N_13496);
nand U13622 (N_13622,N_13465,N_13508);
or U13623 (N_13623,N_13586,N_13549);
and U13624 (N_13624,N_13484,N_13498);
xnor U13625 (N_13625,N_13559,N_13464);
or U13626 (N_13626,N_13590,N_13478);
xor U13627 (N_13627,N_13475,N_13462);
nor U13628 (N_13628,N_13593,N_13501);
and U13629 (N_13629,N_13552,N_13486);
xor U13630 (N_13630,N_13455,N_13541);
or U13631 (N_13631,N_13537,N_13583);
or U13632 (N_13632,N_13525,N_13499);
nor U13633 (N_13633,N_13566,N_13548);
or U13634 (N_13634,N_13440,N_13550);
or U13635 (N_13635,N_13598,N_13544);
or U13636 (N_13636,N_13460,N_13507);
or U13637 (N_13637,N_13457,N_13519);
or U13638 (N_13638,N_13494,N_13575);
and U13639 (N_13639,N_13558,N_13527);
and U13640 (N_13640,N_13506,N_13584);
xnor U13641 (N_13641,N_13533,N_13451);
nand U13642 (N_13642,N_13581,N_13551);
nand U13643 (N_13643,N_13585,N_13447);
nand U13644 (N_13644,N_13445,N_13458);
nor U13645 (N_13645,N_13577,N_13556);
nor U13646 (N_13646,N_13509,N_13592);
or U13647 (N_13647,N_13512,N_13596);
xor U13648 (N_13648,N_13573,N_13574);
xnor U13649 (N_13649,N_13479,N_13500);
xor U13650 (N_13650,N_13505,N_13504);
nor U13651 (N_13651,N_13545,N_13463);
and U13652 (N_13652,N_13497,N_13557);
nor U13653 (N_13653,N_13561,N_13532);
or U13654 (N_13654,N_13441,N_13546);
or U13655 (N_13655,N_13526,N_13510);
and U13656 (N_13656,N_13568,N_13576);
xor U13657 (N_13657,N_13553,N_13597);
xnor U13658 (N_13658,N_13461,N_13515);
nor U13659 (N_13659,N_13529,N_13490);
nand U13660 (N_13660,N_13595,N_13572);
nor U13661 (N_13661,N_13514,N_13560);
and U13662 (N_13662,N_13443,N_13516);
nor U13663 (N_13663,N_13485,N_13459);
nand U13664 (N_13664,N_13492,N_13571);
and U13665 (N_13665,N_13448,N_13540);
xnor U13666 (N_13666,N_13493,N_13534);
xnor U13667 (N_13667,N_13487,N_13450);
nor U13668 (N_13668,N_13480,N_13518);
and U13669 (N_13669,N_13547,N_13539);
nor U13670 (N_13670,N_13476,N_13454);
xor U13671 (N_13671,N_13531,N_13523);
and U13672 (N_13672,N_13482,N_13530);
nor U13673 (N_13673,N_13502,N_13468);
nor U13674 (N_13674,N_13589,N_13524);
nand U13675 (N_13675,N_13555,N_13587);
and U13676 (N_13676,N_13588,N_13522);
nor U13677 (N_13677,N_13594,N_13543);
and U13678 (N_13678,N_13517,N_13521);
xnor U13679 (N_13679,N_13483,N_13495);
xor U13680 (N_13680,N_13550,N_13589);
nand U13681 (N_13681,N_13445,N_13460);
xnor U13682 (N_13682,N_13574,N_13509);
xor U13683 (N_13683,N_13531,N_13504);
or U13684 (N_13684,N_13476,N_13452);
xnor U13685 (N_13685,N_13523,N_13524);
xor U13686 (N_13686,N_13447,N_13462);
or U13687 (N_13687,N_13450,N_13475);
nor U13688 (N_13688,N_13505,N_13540);
nand U13689 (N_13689,N_13577,N_13505);
or U13690 (N_13690,N_13507,N_13443);
nand U13691 (N_13691,N_13454,N_13593);
nor U13692 (N_13692,N_13599,N_13489);
nand U13693 (N_13693,N_13512,N_13440);
nor U13694 (N_13694,N_13505,N_13499);
or U13695 (N_13695,N_13497,N_13468);
or U13696 (N_13696,N_13537,N_13476);
nand U13697 (N_13697,N_13574,N_13450);
xor U13698 (N_13698,N_13578,N_13465);
nand U13699 (N_13699,N_13583,N_13516);
xor U13700 (N_13700,N_13457,N_13507);
nor U13701 (N_13701,N_13565,N_13595);
xor U13702 (N_13702,N_13541,N_13566);
xor U13703 (N_13703,N_13486,N_13549);
nor U13704 (N_13704,N_13514,N_13534);
or U13705 (N_13705,N_13555,N_13441);
nor U13706 (N_13706,N_13453,N_13469);
or U13707 (N_13707,N_13546,N_13589);
nor U13708 (N_13708,N_13566,N_13554);
nor U13709 (N_13709,N_13548,N_13442);
nor U13710 (N_13710,N_13473,N_13592);
nand U13711 (N_13711,N_13528,N_13518);
nand U13712 (N_13712,N_13475,N_13529);
or U13713 (N_13713,N_13477,N_13478);
xor U13714 (N_13714,N_13566,N_13466);
nand U13715 (N_13715,N_13504,N_13577);
or U13716 (N_13716,N_13504,N_13472);
or U13717 (N_13717,N_13563,N_13532);
xor U13718 (N_13718,N_13540,N_13453);
and U13719 (N_13719,N_13560,N_13599);
nand U13720 (N_13720,N_13458,N_13547);
or U13721 (N_13721,N_13575,N_13561);
or U13722 (N_13722,N_13468,N_13536);
xor U13723 (N_13723,N_13555,N_13497);
or U13724 (N_13724,N_13456,N_13448);
nand U13725 (N_13725,N_13480,N_13543);
xor U13726 (N_13726,N_13572,N_13454);
xnor U13727 (N_13727,N_13569,N_13519);
nand U13728 (N_13728,N_13582,N_13590);
nand U13729 (N_13729,N_13517,N_13559);
nand U13730 (N_13730,N_13511,N_13459);
xnor U13731 (N_13731,N_13571,N_13442);
and U13732 (N_13732,N_13477,N_13569);
or U13733 (N_13733,N_13443,N_13448);
nor U13734 (N_13734,N_13506,N_13541);
nor U13735 (N_13735,N_13544,N_13572);
nor U13736 (N_13736,N_13446,N_13584);
nor U13737 (N_13737,N_13544,N_13499);
or U13738 (N_13738,N_13440,N_13474);
xor U13739 (N_13739,N_13452,N_13551);
nand U13740 (N_13740,N_13556,N_13583);
or U13741 (N_13741,N_13577,N_13561);
or U13742 (N_13742,N_13478,N_13597);
or U13743 (N_13743,N_13506,N_13543);
nor U13744 (N_13744,N_13569,N_13512);
xnor U13745 (N_13745,N_13572,N_13589);
nor U13746 (N_13746,N_13564,N_13576);
xnor U13747 (N_13747,N_13535,N_13597);
and U13748 (N_13748,N_13573,N_13542);
nor U13749 (N_13749,N_13475,N_13528);
nand U13750 (N_13750,N_13537,N_13509);
and U13751 (N_13751,N_13571,N_13472);
and U13752 (N_13752,N_13515,N_13468);
xor U13753 (N_13753,N_13599,N_13444);
nand U13754 (N_13754,N_13526,N_13493);
or U13755 (N_13755,N_13550,N_13444);
xnor U13756 (N_13756,N_13572,N_13450);
xor U13757 (N_13757,N_13539,N_13477);
or U13758 (N_13758,N_13456,N_13530);
xor U13759 (N_13759,N_13523,N_13528);
nor U13760 (N_13760,N_13604,N_13732);
nand U13761 (N_13761,N_13651,N_13756);
and U13762 (N_13762,N_13610,N_13718);
and U13763 (N_13763,N_13676,N_13662);
nor U13764 (N_13764,N_13634,N_13744);
nor U13765 (N_13765,N_13609,N_13614);
and U13766 (N_13766,N_13658,N_13612);
xnor U13767 (N_13767,N_13638,N_13708);
and U13768 (N_13768,N_13671,N_13600);
and U13769 (N_13769,N_13643,N_13706);
xnor U13770 (N_13770,N_13606,N_13738);
xnor U13771 (N_13771,N_13703,N_13728);
xnor U13772 (N_13772,N_13664,N_13680);
nor U13773 (N_13773,N_13733,N_13675);
and U13774 (N_13774,N_13617,N_13754);
xnor U13775 (N_13775,N_13700,N_13655);
nor U13776 (N_13776,N_13698,N_13699);
nand U13777 (N_13777,N_13684,N_13729);
nand U13778 (N_13778,N_13626,N_13711);
nand U13779 (N_13779,N_13715,N_13727);
or U13780 (N_13780,N_13619,N_13724);
nand U13781 (N_13781,N_13613,N_13618);
nand U13782 (N_13782,N_13678,N_13747);
and U13783 (N_13783,N_13639,N_13605);
nand U13784 (N_13784,N_13697,N_13755);
nand U13785 (N_13785,N_13702,N_13622);
xor U13786 (N_13786,N_13681,N_13674);
or U13787 (N_13787,N_13739,N_13752);
xor U13788 (N_13788,N_13685,N_13652);
or U13789 (N_13789,N_13661,N_13737);
xor U13790 (N_13790,N_13633,N_13736);
and U13791 (N_13791,N_13644,N_13672);
xor U13792 (N_13792,N_13602,N_13656);
xor U13793 (N_13793,N_13628,N_13745);
or U13794 (N_13794,N_13657,N_13713);
and U13795 (N_13795,N_13712,N_13731);
nor U13796 (N_13796,N_13630,N_13743);
or U13797 (N_13797,N_13694,N_13714);
nand U13798 (N_13798,N_13689,N_13627);
or U13799 (N_13799,N_13757,N_13642);
nand U13800 (N_13800,N_13691,N_13753);
and U13801 (N_13801,N_13635,N_13704);
or U13802 (N_13802,N_13723,N_13663);
nor U13803 (N_13803,N_13607,N_13659);
xor U13804 (N_13804,N_13624,N_13632);
and U13805 (N_13805,N_13645,N_13603);
and U13806 (N_13806,N_13648,N_13726);
xor U13807 (N_13807,N_13749,N_13696);
nor U13808 (N_13808,N_13621,N_13647);
nor U13809 (N_13809,N_13722,N_13620);
nand U13810 (N_13810,N_13758,N_13751);
nand U13811 (N_13811,N_13683,N_13730);
xor U13812 (N_13812,N_13750,N_13705);
or U13813 (N_13813,N_13616,N_13660);
or U13814 (N_13814,N_13721,N_13650);
xnor U13815 (N_13815,N_13695,N_13710);
nor U13816 (N_13816,N_13742,N_13673);
xnor U13817 (N_13817,N_13666,N_13759);
nand U13818 (N_13818,N_13631,N_13690);
nand U13819 (N_13819,N_13625,N_13623);
nand U13820 (N_13820,N_13629,N_13669);
xor U13821 (N_13821,N_13682,N_13693);
and U13822 (N_13822,N_13679,N_13641);
xor U13823 (N_13823,N_13665,N_13717);
and U13824 (N_13824,N_13611,N_13740);
nor U13825 (N_13825,N_13654,N_13701);
or U13826 (N_13826,N_13637,N_13677);
or U13827 (N_13827,N_13601,N_13707);
xor U13828 (N_13828,N_13608,N_13716);
xnor U13829 (N_13829,N_13649,N_13615);
or U13830 (N_13830,N_13646,N_13709);
or U13831 (N_13831,N_13686,N_13668);
nor U13832 (N_13832,N_13687,N_13667);
and U13833 (N_13833,N_13720,N_13692);
or U13834 (N_13834,N_13719,N_13653);
or U13835 (N_13835,N_13725,N_13746);
nand U13836 (N_13836,N_13748,N_13636);
or U13837 (N_13837,N_13688,N_13640);
and U13838 (N_13838,N_13741,N_13734);
nor U13839 (N_13839,N_13670,N_13735);
xor U13840 (N_13840,N_13725,N_13636);
nor U13841 (N_13841,N_13615,N_13678);
and U13842 (N_13842,N_13635,N_13636);
and U13843 (N_13843,N_13671,N_13707);
or U13844 (N_13844,N_13622,N_13698);
nand U13845 (N_13845,N_13750,N_13717);
nand U13846 (N_13846,N_13744,N_13713);
nor U13847 (N_13847,N_13607,N_13707);
xnor U13848 (N_13848,N_13621,N_13755);
nor U13849 (N_13849,N_13678,N_13602);
or U13850 (N_13850,N_13745,N_13710);
xor U13851 (N_13851,N_13730,N_13627);
or U13852 (N_13852,N_13745,N_13643);
and U13853 (N_13853,N_13642,N_13737);
xor U13854 (N_13854,N_13675,N_13604);
nor U13855 (N_13855,N_13748,N_13626);
xor U13856 (N_13856,N_13662,N_13759);
nor U13857 (N_13857,N_13672,N_13745);
nand U13858 (N_13858,N_13628,N_13721);
or U13859 (N_13859,N_13619,N_13710);
and U13860 (N_13860,N_13711,N_13751);
and U13861 (N_13861,N_13613,N_13647);
xor U13862 (N_13862,N_13727,N_13676);
xor U13863 (N_13863,N_13684,N_13601);
and U13864 (N_13864,N_13692,N_13602);
nand U13865 (N_13865,N_13627,N_13645);
and U13866 (N_13866,N_13684,N_13665);
or U13867 (N_13867,N_13647,N_13663);
and U13868 (N_13868,N_13655,N_13674);
nand U13869 (N_13869,N_13636,N_13730);
xnor U13870 (N_13870,N_13742,N_13648);
xor U13871 (N_13871,N_13715,N_13742);
or U13872 (N_13872,N_13609,N_13717);
nor U13873 (N_13873,N_13643,N_13679);
xnor U13874 (N_13874,N_13643,N_13735);
xor U13875 (N_13875,N_13736,N_13708);
xnor U13876 (N_13876,N_13663,N_13642);
nand U13877 (N_13877,N_13601,N_13664);
nand U13878 (N_13878,N_13720,N_13638);
or U13879 (N_13879,N_13623,N_13636);
or U13880 (N_13880,N_13731,N_13715);
and U13881 (N_13881,N_13732,N_13721);
nor U13882 (N_13882,N_13612,N_13642);
nor U13883 (N_13883,N_13668,N_13607);
or U13884 (N_13884,N_13626,N_13684);
and U13885 (N_13885,N_13751,N_13671);
xnor U13886 (N_13886,N_13709,N_13713);
and U13887 (N_13887,N_13601,N_13663);
and U13888 (N_13888,N_13618,N_13687);
nand U13889 (N_13889,N_13608,N_13695);
nor U13890 (N_13890,N_13676,N_13665);
xnor U13891 (N_13891,N_13734,N_13717);
nor U13892 (N_13892,N_13645,N_13722);
nor U13893 (N_13893,N_13756,N_13663);
or U13894 (N_13894,N_13621,N_13633);
or U13895 (N_13895,N_13643,N_13611);
or U13896 (N_13896,N_13719,N_13740);
or U13897 (N_13897,N_13724,N_13695);
xnor U13898 (N_13898,N_13692,N_13678);
nor U13899 (N_13899,N_13750,N_13604);
and U13900 (N_13900,N_13628,N_13619);
and U13901 (N_13901,N_13692,N_13675);
and U13902 (N_13902,N_13715,N_13636);
nor U13903 (N_13903,N_13634,N_13641);
nand U13904 (N_13904,N_13701,N_13699);
nand U13905 (N_13905,N_13647,N_13682);
xnor U13906 (N_13906,N_13604,N_13727);
or U13907 (N_13907,N_13715,N_13707);
and U13908 (N_13908,N_13729,N_13744);
nand U13909 (N_13909,N_13726,N_13604);
or U13910 (N_13910,N_13724,N_13729);
nor U13911 (N_13911,N_13630,N_13624);
nand U13912 (N_13912,N_13636,N_13681);
nand U13913 (N_13913,N_13666,N_13643);
nor U13914 (N_13914,N_13736,N_13614);
or U13915 (N_13915,N_13640,N_13734);
xor U13916 (N_13916,N_13696,N_13661);
xor U13917 (N_13917,N_13708,N_13651);
nand U13918 (N_13918,N_13734,N_13664);
or U13919 (N_13919,N_13616,N_13676);
nor U13920 (N_13920,N_13796,N_13874);
and U13921 (N_13921,N_13830,N_13808);
or U13922 (N_13922,N_13803,N_13783);
and U13923 (N_13923,N_13843,N_13817);
or U13924 (N_13924,N_13907,N_13814);
and U13925 (N_13925,N_13906,N_13799);
and U13926 (N_13926,N_13816,N_13894);
nor U13927 (N_13927,N_13898,N_13837);
nand U13928 (N_13928,N_13798,N_13910);
nor U13929 (N_13929,N_13809,N_13868);
or U13930 (N_13930,N_13805,N_13865);
or U13931 (N_13931,N_13899,N_13876);
nor U13932 (N_13932,N_13835,N_13883);
and U13933 (N_13933,N_13797,N_13795);
nand U13934 (N_13934,N_13813,N_13790);
nor U13935 (N_13935,N_13834,N_13774);
nand U13936 (N_13936,N_13818,N_13806);
nor U13937 (N_13937,N_13789,N_13776);
and U13938 (N_13938,N_13903,N_13765);
nor U13939 (N_13939,N_13823,N_13915);
and U13940 (N_13940,N_13885,N_13872);
or U13941 (N_13941,N_13879,N_13788);
nand U13942 (N_13942,N_13794,N_13918);
and U13943 (N_13943,N_13833,N_13841);
xor U13944 (N_13944,N_13802,N_13780);
xor U13945 (N_13945,N_13896,N_13862);
nor U13946 (N_13946,N_13858,N_13863);
or U13947 (N_13947,N_13856,N_13845);
nand U13948 (N_13948,N_13861,N_13839);
xor U13949 (N_13949,N_13836,N_13786);
nand U13950 (N_13950,N_13764,N_13912);
xnor U13951 (N_13951,N_13873,N_13913);
or U13952 (N_13952,N_13888,N_13866);
nor U13953 (N_13953,N_13769,N_13775);
and U13954 (N_13954,N_13807,N_13778);
xnor U13955 (N_13955,N_13821,N_13804);
nor U13956 (N_13956,N_13893,N_13880);
xor U13957 (N_13957,N_13772,N_13771);
and U13958 (N_13958,N_13777,N_13911);
and U13959 (N_13959,N_13792,N_13857);
xor U13960 (N_13960,N_13800,N_13890);
and U13961 (N_13961,N_13815,N_13827);
or U13962 (N_13962,N_13869,N_13826);
nor U13963 (N_13963,N_13779,N_13919);
nand U13964 (N_13964,N_13832,N_13828);
and U13965 (N_13965,N_13822,N_13842);
nor U13966 (N_13966,N_13891,N_13824);
and U13967 (N_13967,N_13870,N_13909);
xor U13968 (N_13968,N_13787,N_13895);
and U13969 (N_13969,N_13852,N_13760);
xor U13970 (N_13970,N_13851,N_13914);
nor U13971 (N_13971,N_13811,N_13901);
nand U13972 (N_13972,N_13782,N_13902);
and U13973 (N_13973,N_13785,N_13768);
nand U13974 (N_13974,N_13877,N_13829);
nor U13975 (N_13975,N_13849,N_13761);
nand U13976 (N_13976,N_13905,N_13773);
and U13977 (N_13977,N_13860,N_13875);
nand U13978 (N_13978,N_13867,N_13825);
nor U13979 (N_13979,N_13853,N_13770);
or U13980 (N_13980,N_13882,N_13801);
nor U13981 (N_13981,N_13886,N_13900);
nor U13982 (N_13982,N_13762,N_13844);
nor U13983 (N_13983,N_13855,N_13848);
nor U13984 (N_13984,N_13917,N_13850);
nand U13985 (N_13985,N_13840,N_13791);
xor U13986 (N_13986,N_13810,N_13793);
nand U13987 (N_13987,N_13812,N_13897);
and U13988 (N_13988,N_13784,N_13887);
xor U13989 (N_13989,N_13916,N_13781);
xnor U13990 (N_13990,N_13766,N_13819);
and U13991 (N_13991,N_13838,N_13831);
nor U13992 (N_13992,N_13864,N_13847);
xnor U13993 (N_13993,N_13892,N_13763);
nand U13994 (N_13994,N_13889,N_13878);
xnor U13995 (N_13995,N_13767,N_13820);
and U13996 (N_13996,N_13846,N_13854);
nor U13997 (N_13997,N_13908,N_13884);
nand U13998 (N_13998,N_13871,N_13904);
nor U13999 (N_13999,N_13859,N_13881);
or U14000 (N_14000,N_13784,N_13893);
nor U14001 (N_14001,N_13871,N_13783);
or U14002 (N_14002,N_13767,N_13881);
or U14003 (N_14003,N_13831,N_13913);
and U14004 (N_14004,N_13895,N_13789);
nand U14005 (N_14005,N_13844,N_13876);
nand U14006 (N_14006,N_13889,N_13879);
nor U14007 (N_14007,N_13846,N_13806);
xor U14008 (N_14008,N_13819,N_13832);
xnor U14009 (N_14009,N_13894,N_13917);
or U14010 (N_14010,N_13794,N_13789);
or U14011 (N_14011,N_13916,N_13812);
and U14012 (N_14012,N_13910,N_13773);
and U14013 (N_14013,N_13904,N_13807);
xnor U14014 (N_14014,N_13856,N_13841);
and U14015 (N_14015,N_13813,N_13895);
nand U14016 (N_14016,N_13809,N_13779);
and U14017 (N_14017,N_13868,N_13762);
nor U14018 (N_14018,N_13878,N_13909);
xnor U14019 (N_14019,N_13835,N_13914);
or U14020 (N_14020,N_13875,N_13815);
nand U14021 (N_14021,N_13808,N_13780);
nor U14022 (N_14022,N_13855,N_13846);
and U14023 (N_14023,N_13803,N_13822);
and U14024 (N_14024,N_13855,N_13830);
and U14025 (N_14025,N_13808,N_13876);
xor U14026 (N_14026,N_13774,N_13825);
or U14027 (N_14027,N_13823,N_13818);
xnor U14028 (N_14028,N_13824,N_13837);
nor U14029 (N_14029,N_13829,N_13801);
and U14030 (N_14030,N_13793,N_13819);
xor U14031 (N_14031,N_13918,N_13804);
and U14032 (N_14032,N_13856,N_13804);
or U14033 (N_14033,N_13903,N_13863);
or U14034 (N_14034,N_13826,N_13854);
nand U14035 (N_14035,N_13895,N_13833);
nand U14036 (N_14036,N_13779,N_13781);
and U14037 (N_14037,N_13775,N_13911);
or U14038 (N_14038,N_13856,N_13824);
or U14039 (N_14039,N_13904,N_13856);
nor U14040 (N_14040,N_13801,N_13854);
or U14041 (N_14041,N_13817,N_13916);
and U14042 (N_14042,N_13797,N_13844);
nand U14043 (N_14043,N_13770,N_13799);
nor U14044 (N_14044,N_13763,N_13884);
or U14045 (N_14045,N_13878,N_13886);
nand U14046 (N_14046,N_13888,N_13881);
nor U14047 (N_14047,N_13834,N_13879);
or U14048 (N_14048,N_13854,N_13794);
nor U14049 (N_14049,N_13766,N_13769);
xor U14050 (N_14050,N_13866,N_13787);
xor U14051 (N_14051,N_13915,N_13880);
xnor U14052 (N_14052,N_13818,N_13773);
and U14053 (N_14053,N_13815,N_13772);
and U14054 (N_14054,N_13836,N_13816);
nor U14055 (N_14055,N_13903,N_13891);
xnor U14056 (N_14056,N_13912,N_13872);
and U14057 (N_14057,N_13897,N_13825);
xor U14058 (N_14058,N_13814,N_13875);
nor U14059 (N_14059,N_13887,N_13763);
and U14060 (N_14060,N_13896,N_13849);
xor U14061 (N_14061,N_13805,N_13889);
nor U14062 (N_14062,N_13855,N_13887);
nand U14063 (N_14063,N_13850,N_13794);
nor U14064 (N_14064,N_13914,N_13783);
or U14065 (N_14065,N_13829,N_13788);
xnor U14066 (N_14066,N_13788,N_13855);
and U14067 (N_14067,N_13866,N_13835);
nor U14068 (N_14068,N_13809,N_13776);
xnor U14069 (N_14069,N_13764,N_13813);
xnor U14070 (N_14070,N_13789,N_13874);
and U14071 (N_14071,N_13852,N_13918);
xnor U14072 (N_14072,N_13915,N_13919);
xnor U14073 (N_14073,N_13773,N_13807);
xnor U14074 (N_14074,N_13854,N_13825);
nand U14075 (N_14075,N_13858,N_13884);
or U14076 (N_14076,N_13848,N_13865);
nand U14077 (N_14077,N_13888,N_13839);
nand U14078 (N_14078,N_13840,N_13762);
or U14079 (N_14079,N_13899,N_13789);
or U14080 (N_14080,N_13936,N_13941);
and U14081 (N_14081,N_13921,N_13980);
or U14082 (N_14082,N_13973,N_14039);
and U14083 (N_14083,N_14015,N_14017);
and U14084 (N_14084,N_14011,N_13954);
nor U14085 (N_14085,N_14068,N_14013);
and U14086 (N_14086,N_14022,N_13990);
and U14087 (N_14087,N_14063,N_13987);
and U14088 (N_14088,N_14060,N_13984);
or U14089 (N_14089,N_13953,N_14061);
nand U14090 (N_14090,N_13946,N_13983);
nor U14091 (N_14091,N_13940,N_13935);
and U14092 (N_14092,N_13971,N_14024);
nor U14093 (N_14093,N_14001,N_14009);
and U14094 (N_14094,N_13957,N_13930);
nor U14095 (N_14095,N_13950,N_13989);
or U14096 (N_14096,N_13993,N_13988);
xnor U14097 (N_14097,N_14002,N_14040);
and U14098 (N_14098,N_14019,N_13982);
or U14099 (N_14099,N_13962,N_13924);
nand U14100 (N_14100,N_14048,N_14042);
nor U14101 (N_14101,N_13927,N_14043);
xnor U14102 (N_14102,N_14076,N_13942);
or U14103 (N_14103,N_14047,N_14062);
xnor U14104 (N_14104,N_14012,N_13981);
and U14105 (N_14105,N_14044,N_13949);
xnor U14106 (N_14106,N_13938,N_14000);
nor U14107 (N_14107,N_13934,N_14008);
nand U14108 (N_14108,N_14053,N_14038);
xor U14109 (N_14109,N_13986,N_14051);
nor U14110 (N_14110,N_13968,N_13997);
nand U14111 (N_14111,N_14057,N_13948);
and U14112 (N_14112,N_14072,N_14026);
nand U14113 (N_14113,N_14078,N_13977);
xnor U14114 (N_14114,N_13965,N_13976);
xor U14115 (N_14115,N_13939,N_14052);
or U14116 (N_14116,N_14059,N_14049);
nor U14117 (N_14117,N_14066,N_13994);
nor U14118 (N_14118,N_14004,N_14014);
or U14119 (N_14119,N_14027,N_13932);
or U14120 (N_14120,N_13944,N_14041);
nor U14121 (N_14121,N_13960,N_14030);
nor U14122 (N_14122,N_13923,N_13956);
nor U14123 (N_14123,N_14020,N_13951);
xnor U14124 (N_14124,N_14079,N_14077);
xor U14125 (N_14125,N_14065,N_13998);
or U14126 (N_14126,N_13967,N_14034);
nor U14127 (N_14127,N_14029,N_13952);
and U14128 (N_14128,N_13985,N_14070);
nand U14129 (N_14129,N_13996,N_13963);
xor U14130 (N_14130,N_13943,N_13975);
nand U14131 (N_14131,N_13964,N_13929);
and U14132 (N_14132,N_13920,N_14007);
and U14133 (N_14133,N_14016,N_13955);
and U14134 (N_14134,N_14074,N_13922);
nor U14135 (N_14135,N_13995,N_14046);
xor U14136 (N_14136,N_13945,N_14037);
xor U14137 (N_14137,N_13928,N_13961);
or U14138 (N_14138,N_14032,N_13979);
nor U14139 (N_14139,N_14036,N_14033);
and U14140 (N_14140,N_14050,N_13974);
and U14141 (N_14141,N_13978,N_14003);
xor U14142 (N_14142,N_14069,N_14010);
or U14143 (N_14143,N_13933,N_14055);
or U14144 (N_14144,N_13991,N_13969);
xor U14145 (N_14145,N_13937,N_14075);
and U14146 (N_14146,N_13931,N_14021);
nor U14147 (N_14147,N_13966,N_14067);
or U14148 (N_14148,N_13926,N_13999);
or U14149 (N_14149,N_14056,N_14005);
nand U14150 (N_14150,N_14031,N_14071);
or U14151 (N_14151,N_14006,N_14035);
or U14152 (N_14152,N_14064,N_13970);
nor U14153 (N_14153,N_13992,N_13972);
nor U14154 (N_14154,N_14054,N_13958);
xor U14155 (N_14155,N_14058,N_13925);
xor U14156 (N_14156,N_13959,N_14023);
nand U14157 (N_14157,N_13947,N_14028);
nor U14158 (N_14158,N_14045,N_14073);
nand U14159 (N_14159,N_14018,N_14025);
and U14160 (N_14160,N_13953,N_13952);
and U14161 (N_14161,N_13963,N_13995);
nand U14162 (N_14162,N_13973,N_13971);
nand U14163 (N_14163,N_14006,N_13983);
nor U14164 (N_14164,N_14002,N_13979);
and U14165 (N_14165,N_13946,N_14020);
and U14166 (N_14166,N_14060,N_14074);
nor U14167 (N_14167,N_13998,N_14016);
nor U14168 (N_14168,N_14005,N_13962);
nor U14169 (N_14169,N_13965,N_14006);
nand U14170 (N_14170,N_14077,N_13985);
xor U14171 (N_14171,N_14070,N_14077);
nand U14172 (N_14172,N_13933,N_14003);
nor U14173 (N_14173,N_13924,N_14066);
or U14174 (N_14174,N_13983,N_14040);
nand U14175 (N_14175,N_13990,N_13927);
or U14176 (N_14176,N_14009,N_13987);
nand U14177 (N_14177,N_13955,N_13927);
or U14178 (N_14178,N_13941,N_14038);
and U14179 (N_14179,N_13934,N_14055);
nand U14180 (N_14180,N_13931,N_13947);
and U14181 (N_14181,N_13989,N_14050);
nand U14182 (N_14182,N_14066,N_14021);
nor U14183 (N_14183,N_14065,N_14048);
nand U14184 (N_14184,N_14044,N_13920);
and U14185 (N_14185,N_14041,N_14069);
or U14186 (N_14186,N_13969,N_13936);
xor U14187 (N_14187,N_13940,N_14012);
nor U14188 (N_14188,N_13930,N_14023);
nor U14189 (N_14189,N_13935,N_14044);
nor U14190 (N_14190,N_14078,N_14033);
xor U14191 (N_14191,N_14022,N_13966);
xor U14192 (N_14192,N_13927,N_13926);
nand U14193 (N_14193,N_14018,N_13991);
and U14194 (N_14194,N_14074,N_14028);
or U14195 (N_14195,N_14040,N_14005);
and U14196 (N_14196,N_14010,N_13941);
xor U14197 (N_14197,N_14032,N_13956);
and U14198 (N_14198,N_13985,N_14012);
or U14199 (N_14199,N_13976,N_13927);
and U14200 (N_14200,N_13955,N_14076);
nor U14201 (N_14201,N_14078,N_14058);
and U14202 (N_14202,N_13988,N_13976);
xnor U14203 (N_14203,N_13987,N_14019);
nor U14204 (N_14204,N_13978,N_13950);
or U14205 (N_14205,N_13942,N_14022);
xor U14206 (N_14206,N_14018,N_14044);
nand U14207 (N_14207,N_13977,N_14041);
and U14208 (N_14208,N_13930,N_14027);
nor U14209 (N_14209,N_13922,N_14038);
nand U14210 (N_14210,N_13944,N_13963);
nand U14211 (N_14211,N_14022,N_13976);
nor U14212 (N_14212,N_14021,N_13944);
nor U14213 (N_14213,N_14059,N_13991);
or U14214 (N_14214,N_14008,N_13978);
nor U14215 (N_14215,N_13959,N_13983);
and U14216 (N_14216,N_13925,N_14031);
or U14217 (N_14217,N_14057,N_13989);
nand U14218 (N_14218,N_14028,N_14043);
nor U14219 (N_14219,N_14051,N_14067);
nor U14220 (N_14220,N_13925,N_14019);
and U14221 (N_14221,N_14060,N_14039);
nor U14222 (N_14222,N_13957,N_14034);
and U14223 (N_14223,N_14062,N_13934);
nor U14224 (N_14224,N_13986,N_13960);
nand U14225 (N_14225,N_13962,N_13922);
nor U14226 (N_14226,N_14054,N_14005);
nor U14227 (N_14227,N_14047,N_13936);
xnor U14228 (N_14228,N_13987,N_13968);
xnor U14229 (N_14229,N_13934,N_13951);
and U14230 (N_14230,N_13941,N_14050);
or U14231 (N_14231,N_13955,N_13991);
or U14232 (N_14232,N_14047,N_13998);
and U14233 (N_14233,N_14003,N_14030);
nor U14234 (N_14234,N_13939,N_14070);
nand U14235 (N_14235,N_14063,N_13928);
and U14236 (N_14236,N_13995,N_13941);
nor U14237 (N_14237,N_13976,N_13971);
nor U14238 (N_14238,N_13965,N_13931);
or U14239 (N_14239,N_14062,N_13931);
nand U14240 (N_14240,N_14189,N_14233);
or U14241 (N_14241,N_14174,N_14099);
nor U14242 (N_14242,N_14183,N_14091);
and U14243 (N_14243,N_14104,N_14190);
nand U14244 (N_14244,N_14197,N_14156);
and U14245 (N_14245,N_14141,N_14132);
and U14246 (N_14246,N_14228,N_14222);
nor U14247 (N_14247,N_14084,N_14115);
or U14248 (N_14248,N_14165,N_14148);
or U14249 (N_14249,N_14163,N_14143);
and U14250 (N_14250,N_14216,N_14234);
or U14251 (N_14251,N_14198,N_14162);
nor U14252 (N_14252,N_14114,N_14166);
nor U14253 (N_14253,N_14127,N_14160);
nand U14254 (N_14254,N_14221,N_14144);
xor U14255 (N_14255,N_14173,N_14086);
nand U14256 (N_14256,N_14106,N_14113);
nor U14257 (N_14257,N_14210,N_14085);
and U14258 (N_14258,N_14168,N_14218);
nand U14259 (N_14259,N_14219,N_14192);
or U14260 (N_14260,N_14139,N_14147);
nor U14261 (N_14261,N_14149,N_14172);
and U14262 (N_14262,N_14153,N_14231);
and U14263 (N_14263,N_14184,N_14154);
nor U14264 (N_14264,N_14109,N_14229);
xor U14265 (N_14265,N_14169,N_14208);
nor U14266 (N_14266,N_14111,N_14237);
and U14267 (N_14267,N_14136,N_14080);
nor U14268 (N_14268,N_14176,N_14236);
and U14269 (N_14269,N_14205,N_14097);
or U14270 (N_14270,N_14187,N_14146);
and U14271 (N_14271,N_14100,N_14158);
nand U14272 (N_14272,N_14204,N_14171);
nor U14273 (N_14273,N_14098,N_14137);
or U14274 (N_14274,N_14094,N_14194);
nand U14275 (N_14275,N_14182,N_14203);
nand U14276 (N_14276,N_14207,N_14105);
xnor U14277 (N_14277,N_14090,N_14223);
nor U14278 (N_14278,N_14170,N_14101);
nand U14279 (N_14279,N_14112,N_14226);
or U14280 (N_14280,N_14134,N_14202);
xnor U14281 (N_14281,N_14186,N_14230);
and U14282 (N_14282,N_14110,N_14220);
nor U14283 (N_14283,N_14177,N_14239);
xnor U14284 (N_14284,N_14130,N_14188);
and U14285 (N_14285,N_14140,N_14103);
nand U14286 (N_14286,N_14157,N_14082);
nor U14287 (N_14287,N_14108,N_14209);
nor U14288 (N_14288,N_14119,N_14121);
nor U14289 (N_14289,N_14235,N_14199);
nand U14290 (N_14290,N_14178,N_14096);
xor U14291 (N_14291,N_14215,N_14095);
nor U14292 (N_14292,N_14227,N_14179);
nor U14293 (N_14293,N_14087,N_14180);
and U14294 (N_14294,N_14124,N_14145);
or U14295 (N_14295,N_14088,N_14195);
or U14296 (N_14296,N_14107,N_14122);
nor U14297 (N_14297,N_14150,N_14081);
nand U14298 (N_14298,N_14181,N_14126);
nand U14299 (N_14299,N_14120,N_14211);
xor U14300 (N_14300,N_14093,N_14092);
and U14301 (N_14301,N_14155,N_14138);
nand U14302 (N_14302,N_14175,N_14131);
or U14303 (N_14303,N_14217,N_14117);
xor U14304 (N_14304,N_14152,N_14238);
nor U14305 (N_14305,N_14212,N_14118);
and U14306 (N_14306,N_14129,N_14123);
nand U14307 (N_14307,N_14224,N_14185);
nand U14308 (N_14308,N_14201,N_14232);
or U14309 (N_14309,N_14225,N_14193);
or U14310 (N_14310,N_14083,N_14125);
or U14311 (N_14311,N_14159,N_14128);
and U14312 (N_14312,N_14213,N_14200);
xnor U14313 (N_14313,N_14161,N_14214);
or U14314 (N_14314,N_14135,N_14133);
and U14315 (N_14315,N_14191,N_14164);
and U14316 (N_14316,N_14102,N_14196);
and U14317 (N_14317,N_14151,N_14206);
nand U14318 (N_14318,N_14116,N_14167);
nor U14319 (N_14319,N_14142,N_14089);
nor U14320 (N_14320,N_14100,N_14188);
xor U14321 (N_14321,N_14215,N_14102);
nor U14322 (N_14322,N_14147,N_14106);
and U14323 (N_14323,N_14214,N_14150);
xor U14324 (N_14324,N_14084,N_14208);
nor U14325 (N_14325,N_14120,N_14126);
or U14326 (N_14326,N_14185,N_14196);
or U14327 (N_14327,N_14098,N_14154);
xnor U14328 (N_14328,N_14147,N_14173);
or U14329 (N_14329,N_14207,N_14166);
nor U14330 (N_14330,N_14083,N_14178);
nand U14331 (N_14331,N_14182,N_14167);
or U14332 (N_14332,N_14123,N_14084);
or U14333 (N_14333,N_14125,N_14197);
nand U14334 (N_14334,N_14232,N_14218);
nor U14335 (N_14335,N_14216,N_14090);
xnor U14336 (N_14336,N_14120,N_14124);
nand U14337 (N_14337,N_14121,N_14087);
nand U14338 (N_14338,N_14149,N_14238);
nor U14339 (N_14339,N_14098,N_14122);
nand U14340 (N_14340,N_14136,N_14227);
or U14341 (N_14341,N_14142,N_14104);
nor U14342 (N_14342,N_14080,N_14154);
xor U14343 (N_14343,N_14226,N_14113);
xor U14344 (N_14344,N_14092,N_14187);
nor U14345 (N_14345,N_14223,N_14091);
and U14346 (N_14346,N_14209,N_14237);
xor U14347 (N_14347,N_14082,N_14130);
nor U14348 (N_14348,N_14165,N_14163);
nor U14349 (N_14349,N_14080,N_14100);
nor U14350 (N_14350,N_14181,N_14188);
or U14351 (N_14351,N_14156,N_14142);
xnor U14352 (N_14352,N_14200,N_14099);
nand U14353 (N_14353,N_14172,N_14083);
nor U14354 (N_14354,N_14083,N_14085);
and U14355 (N_14355,N_14107,N_14227);
nand U14356 (N_14356,N_14123,N_14232);
or U14357 (N_14357,N_14111,N_14188);
nand U14358 (N_14358,N_14091,N_14190);
nor U14359 (N_14359,N_14095,N_14236);
or U14360 (N_14360,N_14093,N_14095);
xnor U14361 (N_14361,N_14235,N_14239);
xor U14362 (N_14362,N_14158,N_14099);
or U14363 (N_14363,N_14093,N_14200);
nor U14364 (N_14364,N_14118,N_14122);
nand U14365 (N_14365,N_14132,N_14205);
and U14366 (N_14366,N_14211,N_14196);
and U14367 (N_14367,N_14116,N_14153);
nand U14368 (N_14368,N_14196,N_14224);
xor U14369 (N_14369,N_14152,N_14196);
and U14370 (N_14370,N_14126,N_14116);
or U14371 (N_14371,N_14095,N_14117);
nand U14372 (N_14372,N_14215,N_14178);
nand U14373 (N_14373,N_14129,N_14219);
or U14374 (N_14374,N_14152,N_14111);
nor U14375 (N_14375,N_14106,N_14132);
nand U14376 (N_14376,N_14219,N_14149);
nand U14377 (N_14377,N_14161,N_14206);
nor U14378 (N_14378,N_14188,N_14204);
xnor U14379 (N_14379,N_14129,N_14160);
or U14380 (N_14380,N_14085,N_14185);
nand U14381 (N_14381,N_14125,N_14220);
xnor U14382 (N_14382,N_14118,N_14098);
nor U14383 (N_14383,N_14147,N_14103);
or U14384 (N_14384,N_14154,N_14086);
or U14385 (N_14385,N_14237,N_14134);
and U14386 (N_14386,N_14238,N_14236);
xor U14387 (N_14387,N_14178,N_14126);
and U14388 (N_14388,N_14086,N_14182);
xor U14389 (N_14389,N_14119,N_14113);
and U14390 (N_14390,N_14143,N_14174);
xor U14391 (N_14391,N_14210,N_14238);
and U14392 (N_14392,N_14106,N_14188);
or U14393 (N_14393,N_14087,N_14135);
nor U14394 (N_14394,N_14088,N_14108);
nor U14395 (N_14395,N_14153,N_14201);
nand U14396 (N_14396,N_14095,N_14218);
xor U14397 (N_14397,N_14099,N_14084);
and U14398 (N_14398,N_14217,N_14179);
or U14399 (N_14399,N_14108,N_14167);
nor U14400 (N_14400,N_14287,N_14262);
nand U14401 (N_14401,N_14334,N_14371);
nand U14402 (N_14402,N_14390,N_14320);
xnor U14403 (N_14403,N_14345,N_14283);
nand U14404 (N_14404,N_14360,N_14289);
xor U14405 (N_14405,N_14372,N_14336);
xnor U14406 (N_14406,N_14240,N_14356);
or U14407 (N_14407,N_14359,N_14308);
xnor U14408 (N_14408,N_14374,N_14248);
and U14409 (N_14409,N_14329,N_14286);
and U14410 (N_14410,N_14242,N_14255);
or U14411 (N_14411,N_14305,N_14285);
nor U14412 (N_14412,N_14250,N_14302);
xnor U14413 (N_14413,N_14266,N_14244);
nand U14414 (N_14414,N_14362,N_14269);
or U14415 (N_14415,N_14337,N_14272);
xnor U14416 (N_14416,N_14256,N_14297);
or U14417 (N_14417,N_14369,N_14274);
or U14418 (N_14418,N_14324,N_14261);
or U14419 (N_14419,N_14316,N_14260);
or U14420 (N_14420,N_14361,N_14399);
nor U14421 (N_14421,N_14314,N_14275);
nand U14422 (N_14422,N_14384,N_14385);
nor U14423 (N_14423,N_14296,N_14396);
xnor U14424 (N_14424,N_14273,N_14392);
nand U14425 (N_14425,N_14352,N_14382);
and U14426 (N_14426,N_14357,N_14249);
nor U14427 (N_14427,N_14282,N_14304);
or U14428 (N_14428,N_14292,N_14254);
nand U14429 (N_14429,N_14364,N_14279);
or U14430 (N_14430,N_14263,N_14317);
or U14431 (N_14431,N_14348,N_14258);
or U14432 (N_14432,N_14349,N_14398);
or U14433 (N_14433,N_14322,N_14340);
nor U14434 (N_14434,N_14265,N_14284);
and U14435 (N_14435,N_14315,N_14353);
or U14436 (N_14436,N_14303,N_14389);
or U14437 (N_14437,N_14344,N_14381);
and U14438 (N_14438,N_14391,N_14277);
and U14439 (N_14439,N_14300,N_14341);
xor U14440 (N_14440,N_14290,N_14380);
and U14441 (N_14441,N_14325,N_14376);
nor U14442 (N_14442,N_14306,N_14368);
xnor U14443 (N_14443,N_14331,N_14355);
nor U14444 (N_14444,N_14333,N_14332);
or U14445 (N_14445,N_14245,N_14267);
nor U14446 (N_14446,N_14373,N_14252);
xnor U14447 (N_14447,N_14387,N_14295);
and U14448 (N_14448,N_14335,N_14377);
nor U14449 (N_14449,N_14367,N_14299);
nor U14450 (N_14450,N_14365,N_14358);
xor U14451 (N_14451,N_14343,N_14318);
nand U14452 (N_14452,N_14241,N_14394);
or U14453 (N_14453,N_14350,N_14346);
or U14454 (N_14454,N_14339,N_14281);
or U14455 (N_14455,N_14375,N_14298);
or U14456 (N_14456,N_14301,N_14319);
and U14457 (N_14457,N_14351,N_14395);
xnor U14458 (N_14458,N_14251,N_14247);
or U14459 (N_14459,N_14328,N_14383);
and U14460 (N_14460,N_14309,N_14312);
nand U14461 (N_14461,N_14313,N_14276);
or U14462 (N_14462,N_14271,N_14278);
xor U14463 (N_14463,N_14253,N_14347);
xnor U14464 (N_14464,N_14246,N_14379);
xnor U14465 (N_14465,N_14291,N_14293);
and U14466 (N_14466,N_14363,N_14259);
or U14467 (N_14467,N_14397,N_14280);
nand U14468 (N_14468,N_14294,N_14388);
nand U14469 (N_14469,N_14342,N_14327);
or U14470 (N_14470,N_14310,N_14378);
nand U14471 (N_14471,N_14257,N_14338);
and U14472 (N_14472,N_14326,N_14330);
nor U14473 (N_14473,N_14264,N_14288);
or U14474 (N_14474,N_14243,N_14323);
nand U14475 (N_14475,N_14268,N_14321);
nand U14476 (N_14476,N_14370,N_14366);
nor U14477 (N_14477,N_14311,N_14270);
nand U14478 (N_14478,N_14354,N_14386);
nor U14479 (N_14479,N_14307,N_14393);
nand U14480 (N_14480,N_14297,N_14320);
nor U14481 (N_14481,N_14331,N_14361);
nand U14482 (N_14482,N_14344,N_14364);
and U14483 (N_14483,N_14254,N_14288);
xnor U14484 (N_14484,N_14304,N_14336);
nand U14485 (N_14485,N_14360,N_14313);
and U14486 (N_14486,N_14267,N_14290);
xor U14487 (N_14487,N_14256,N_14351);
nor U14488 (N_14488,N_14378,N_14260);
and U14489 (N_14489,N_14241,N_14387);
or U14490 (N_14490,N_14398,N_14356);
xor U14491 (N_14491,N_14385,N_14382);
xor U14492 (N_14492,N_14319,N_14242);
nor U14493 (N_14493,N_14287,N_14350);
nor U14494 (N_14494,N_14275,N_14298);
xor U14495 (N_14495,N_14377,N_14378);
and U14496 (N_14496,N_14249,N_14308);
xnor U14497 (N_14497,N_14310,N_14384);
nor U14498 (N_14498,N_14340,N_14331);
and U14499 (N_14499,N_14382,N_14383);
xor U14500 (N_14500,N_14266,N_14284);
xnor U14501 (N_14501,N_14302,N_14295);
nor U14502 (N_14502,N_14330,N_14343);
or U14503 (N_14503,N_14286,N_14347);
nand U14504 (N_14504,N_14323,N_14242);
nand U14505 (N_14505,N_14358,N_14357);
nor U14506 (N_14506,N_14257,N_14254);
xor U14507 (N_14507,N_14314,N_14343);
nor U14508 (N_14508,N_14362,N_14242);
nand U14509 (N_14509,N_14384,N_14319);
nor U14510 (N_14510,N_14372,N_14374);
xor U14511 (N_14511,N_14254,N_14323);
and U14512 (N_14512,N_14378,N_14255);
xor U14513 (N_14513,N_14305,N_14369);
xnor U14514 (N_14514,N_14266,N_14339);
nor U14515 (N_14515,N_14356,N_14254);
or U14516 (N_14516,N_14377,N_14309);
and U14517 (N_14517,N_14384,N_14336);
nand U14518 (N_14518,N_14276,N_14261);
nand U14519 (N_14519,N_14270,N_14370);
or U14520 (N_14520,N_14259,N_14285);
and U14521 (N_14521,N_14327,N_14282);
nand U14522 (N_14522,N_14315,N_14288);
xor U14523 (N_14523,N_14356,N_14332);
and U14524 (N_14524,N_14305,N_14299);
nand U14525 (N_14525,N_14370,N_14360);
nor U14526 (N_14526,N_14276,N_14323);
nor U14527 (N_14527,N_14381,N_14370);
nor U14528 (N_14528,N_14293,N_14246);
or U14529 (N_14529,N_14266,N_14328);
xnor U14530 (N_14530,N_14263,N_14262);
or U14531 (N_14531,N_14250,N_14387);
and U14532 (N_14532,N_14305,N_14399);
nand U14533 (N_14533,N_14267,N_14373);
or U14534 (N_14534,N_14388,N_14348);
or U14535 (N_14535,N_14240,N_14317);
and U14536 (N_14536,N_14354,N_14361);
or U14537 (N_14537,N_14269,N_14343);
or U14538 (N_14538,N_14246,N_14388);
xnor U14539 (N_14539,N_14289,N_14246);
nand U14540 (N_14540,N_14317,N_14298);
and U14541 (N_14541,N_14317,N_14384);
nand U14542 (N_14542,N_14243,N_14318);
nand U14543 (N_14543,N_14264,N_14276);
nand U14544 (N_14544,N_14392,N_14285);
nor U14545 (N_14545,N_14274,N_14293);
and U14546 (N_14546,N_14365,N_14337);
or U14547 (N_14547,N_14251,N_14397);
or U14548 (N_14548,N_14348,N_14362);
and U14549 (N_14549,N_14278,N_14360);
and U14550 (N_14550,N_14374,N_14366);
or U14551 (N_14551,N_14340,N_14299);
xor U14552 (N_14552,N_14345,N_14390);
and U14553 (N_14553,N_14251,N_14282);
nand U14554 (N_14554,N_14328,N_14376);
and U14555 (N_14555,N_14313,N_14309);
xnor U14556 (N_14556,N_14301,N_14268);
and U14557 (N_14557,N_14295,N_14285);
xor U14558 (N_14558,N_14330,N_14280);
or U14559 (N_14559,N_14256,N_14330);
xnor U14560 (N_14560,N_14549,N_14425);
nor U14561 (N_14561,N_14551,N_14438);
or U14562 (N_14562,N_14442,N_14518);
xnor U14563 (N_14563,N_14417,N_14456);
and U14564 (N_14564,N_14444,N_14403);
nand U14565 (N_14565,N_14486,N_14452);
nand U14566 (N_14566,N_14407,N_14517);
nor U14567 (N_14567,N_14419,N_14440);
or U14568 (N_14568,N_14516,N_14520);
nor U14569 (N_14569,N_14457,N_14544);
and U14570 (N_14570,N_14441,N_14465);
and U14571 (N_14571,N_14446,N_14526);
and U14572 (N_14572,N_14484,N_14489);
nor U14573 (N_14573,N_14476,N_14409);
nand U14574 (N_14574,N_14541,N_14470);
and U14575 (N_14575,N_14502,N_14401);
nor U14576 (N_14576,N_14427,N_14449);
xnor U14577 (N_14577,N_14492,N_14477);
nor U14578 (N_14578,N_14528,N_14506);
xnor U14579 (N_14579,N_14488,N_14525);
xnor U14580 (N_14580,N_14557,N_14429);
xnor U14581 (N_14581,N_14538,N_14478);
xnor U14582 (N_14582,N_14514,N_14521);
nand U14583 (N_14583,N_14519,N_14494);
nor U14584 (N_14584,N_14454,N_14443);
nand U14585 (N_14585,N_14460,N_14482);
xor U14586 (N_14586,N_14415,N_14522);
xor U14587 (N_14587,N_14402,N_14408);
nand U14588 (N_14588,N_14547,N_14431);
and U14589 (N_14589,N_14527,N_14423);
xnor U14590 (N_14590,N_14469,N_14416);
and U14591 (N_14591,N_14430,N_14453);
xnor U14592 (N_14592,N_14515,N_14435);
and U14593 (N_14593,N_14536,N_14533);
or U14594 (N_14594,N_14451,N_14507);
nand U14595 (N_14595,N_14436,N_14499);
nand U14596 (N_14596,N_14545,N_14542);
nand U14597 (N_14597,N_14432,N_14475);
nor U14598 (N_14598,N_14439,N_14474);
or U14599 (N_14599,N_14433,N_14422);
and U14600 (N_14600,N_14553,N_14413);
or U14601 (N_14601,N_14418,N_14464);
nand U14602 (N_14602,N_14498,N_14467);
nor U14603 (N_14603,N_14480,N_14400);
xnor U14604 (N_14604,N_14412,N_14420);
and U14605 (N_14605,N_14459,N_14428);
xor U14606 (N_14606,N_14463,N_14495);
xor U14607 (N_14607,N_14405,N_14468);
xnor U14608 (N_14608,N_14461,N_14410);
and U14609 (N_14609,N_14532,N_14458);
xor U14610 (N_14610,N_14471,N_14462);
xnor U14611 (N_14611,N_14546,N_14529);
or U14612 (N_14612,N_14426,N_14424);
or U14613 (N_14613,N_14421,N_14513);
nor U14614 (N_14614,N_14448,N_14503);
and U14615 (N_14615,N_14555,N_14404);
nand U14616 (N_14616,N_14496,N_14523);
xnor U14617 (N_14617,N_14455,N_14485);
nand U14618 (N_14618,N_14487,N_14483);
and U14619 (N_14619,N_14437,N_14493);
nor U14620 (N_14620,N_14450,N_14497);
or U14621 (N_14621,N_14543,N_14411);
or U14622 (N_14622,N_14406,N_14479);
xnor U14623 (N_14623,N_14509,N_14559);
nand U14624 (N_14624,N_14505,N_14491);
nand U14625 (N_14625,N_14414,N_14445);
nand U14626 (N_14626,N_14512,N_14552);
or U14627 (N_14627,N_14501,N_14472);
or U14628 (N_14628,N_14558,N_14540);
nor U14629 (N_14629,N_14511,N_14473);
and U14630 (N_14630,N_14539,N_14504);
xor U14631 (N_14631,N_14508,N_14534);
nor U14632 (N_14632,N_14531,N_14535);
and U14633 (N_14633,N_14530,N_14490);
nand U14634 (N_14634,N_14510,N_14447);
xnor U14635 (N_14635,N_14556,N_14500);
xor U14636 (N_14636,N_14537,N_14481);
nor U14637 (N_14637,N_14524,N_14466);
or U14638 (N_14638,N_14548,N_14554);
nor U14639 (N_14639,N_14434,N_14550);
and U14640 (N_14640,N_14502,N_14416);
nor U14641 (N_14641,N_14547,N_14528);
xnor U14642 (N_14642,N_14438,N_14417);
nand U14643 (N_14643,N_14488,N_14451);
xor U14644 (N_14644,N_14420,N_14470);
nand U14645 (N_14645,N_14514,N_14558);
xor U14646 (N_14646,N_14485,N_14499);
and U14647 (N_14647,N_14451,N_14498);
or U14648 (N_14648,N_14448,N_14466);
nand U14649 (N_14649,N_14476,N_14426);
or U14650 (N_14650,N_14464,N_14446);
nand U14651 (N_14651,N_14453,N_14409);
nand U14652 (N_14652,N_14436,N_14554);
and U14653 (N_14653,N_14425,N_14513);
xnor U14654 (N_14654,N_14492,N_14431);
and U14655 (N_14655,N_14511,N_14460);
xor U14656 (N_14656,N_14530,N_14554);
xnor U14657 (N_14657,N_14537,N_14475);
or U14658 (N_14658,N_14555,N_14544);
and U14659 (N_14659,N_14500,N_14442);
or U14660 (N_14660,N_14441,N_14501);
nor U14661 (N_14661,N_14471,N_14520);
nand U14662 (N_14662,N_14477,N_14502);
and U14663 (N_14663,N_14480,N_14440);
nand U14664 (N_14664,N_14455,N_14427);
or U14665 (N_14665,N_14509,N_14542);
or U14666 (N_14666,N_14538,N_14463);
and U14667 (N_14667,N_14489,N_14470);
nand U14668 (N_14668,N_14421,N_14523);
nand U14669 (N_14669,N_14494,N_14410);
nor U14670 (N_14670,N_14490,N_14517);
nor U14671 (N_14671,N_14403,N_14433);
nor U14672 (N_14672,N_14538,N_14551);
xor U14673 (N_14673,N_14541,N_14439);
xnor U14674 (N_14674,N_14422,N_14450);
and U14675 (N_14675,N_14424,N_14421);
nor U14676 (N_14676,N_14447,N_14457);
xor U14677 (N_14677,N_14476,N_14440);
and U14678 (N_14678,N_14518,N_14492);
nand U14679 (N_14679,N_14485,N_14461);
nand U14680 (N_14680,N_14402,N_14445);
nand U14681 (N_14681,N_14439,N_14494);
nand U14682 (N_14682,N_14492,N_14455);
nor U14683 (N_14683,N_14515,N_14411);
nor U14684 (N_14684,N_14478,N_14523);
or U14685 (N_14685,N_14525,N_14519);
xor U14686 (N_14686,N_14431,N_14548);
xor U14687 (N_14687,N_14527,N_14468);
xnor U14688 (N_14688,N_14413,N_14500);
or U14689 (N_14689,N_14459,N_14468);
nor U14690 (N_14690,N_14520,N_14436);
or U14691 (N_14691,N_14445,N_14476);
and U14692 (N_14692,N_14485,N_14536);
xnor U14693 (N_14693,N_14423,N_14406);
nor U14694 (N_14694,N_14478,N_14404);
nand U14695 (N_14695,N_14420,N_14478);
nor U14696 (N_14696,N_14439,N_14476);
xor U14697 (N_14697,N_14456,N_14403);
nor U14698 (N_14698,N_14488,N_14539);
nand U14699 (N_14699,N_14470,N_14428);
xor U14700 (N_14700,N_14538,N_14542);
nand U14701 (N_14701,N_14426,N_14468);
xnor U14702 (N_14702,N_14442,N_14479);
and U14703 (N_14703,N_14439,N_14502);
nand U14704 (N_14704,N_14464,N_14438);
or U14705 (N_14705,N_14529,N_14522);
nor U14706 (N_14706,N_14537,N_14469);
nor U14707 (N_14707,N_14508,N_14530);
and U14708 (N_14708,N_14468,N_14522);
xor U14709 (N_14709,N_14487,N_14456);
or U14710 (N_14710,N_14503,N_14415);
and U14711 (N_14711,N_14546,N_14552);
or U14712 (N_14712,N_14447,N_14482);
nand U14713 (N_14713,N_14498,N_14495);
xnor U14714 (N_14714,N_14426,N_14445);
nand U14715 (N_14715,N_14431,N_14458);
or U14716 (N_14716,N_14538,N_14493);
xnor U14717 (N_14717,N_14473,N_14435);
or U14718 (N_14718,N_14472,N_14502);
or U14719 (N_14719,N_14432,N_14406);
and U14720 (N_14720,N_14656,N_14606);
xnor U14721 (N_14721,N_14664,N_14709);
nand U14722 (N_14722,N_14580,N_14704);
xnor U14723 (N_14723,N_14625,N_14711);
xor U14724 (N_14724,N_14669,N_14659);
and U14725 (N_14725,N_14702,N_14650);
nor U14726 (N_14726,N_14629,N_14567);
nor U14727 (N_14727,N_14717,N_14647);
or U14728 (N_14728,N_14633,N_14662);
nor U14729 (N_14729,N_14707,N_14646);
nand U14730 (N_14730,N_14602,N_14619);
nand U14731 (N_14731,N_14611,N_14620);
or U14732 (N_14732,N_14665,N_14645);
nand U14733 (N_14733,N_14661,N_14560);
nand U14734 (N_14734,N_14701,N_14700);
nor U14735 (N_14735,N_14583,N_14618);
or U14736 (N_14736,N_14719,N_14687);
nor U14737 (N_14737,N_14688,N_14651);
nand U14738 (N_14738,N_14671,N_14684);
xor U14739 (N_14739,N_14696,N_14718);
nor U14740 (N_14740,N_14654,N_14571);
nand U14741 (N_14741,N_14603,N_14642);
xnor U14742 (N_14742,N_14639,N_14674);
xor U14743 (N_14743,N_14621,N_14623);
or U14744 (N_14744,N_14565,N_14607);
nor U14745 (N_14745,N_14569,N_14652);
xnor U14746 (N_14746,N_14628,N_14648);
and U14747 (N_14747,N_14694,N_14568);
nor U14748 (N_14748,N_14585,N_14708);
nor U14749 (N_14749,N_14562,N_14676);
nor U14750 (N_14750,N_14597,N_14706);
xnor U14751 (N_14751,N_14653,N_14561);
or U14752 (N_14752,N_14598,N_14643);
and U14753 (N_14753,N_14614,N_14681);
or U14754 (N_14754,N_14644,N_14692);
xor U14755 (N_14755,N_14663,N_14635);
nand U14756 (N_14756,N_14634,N_14587);
nor U14757 (N_14757,N_14579,N_14622);
nand U14758 (N_14758,N_14589,N_14596);
nand U14759 (N_14759,N_14592,N_14686);
or U14760 (N_14760,N_14605,N_14705);
nand U14761 (N_14761,N_14672,N_14612);
nand U14762 (N_14762,N_14689,N_14682);
or U14763 (N_14763,N_14574,N_14595);
or U14764 (N_14764,N_14575,N_14624);
or U14765 (N_14765,N_14712,N_14673);
and U14766 (N_14766,N_14649,N_14677);
xor U14767 (N_14767,N_14660,N_14637);
or U14768 (N_14768,N_14714,N_14599);
or U14769 (N_14769,N_14578,N_14703);
or U14770 (N_14770,N_14563,N_14668);
and U14771 (N_14771,N_14590,N_14617);
and U14772 (N_14772,N_14570,N_14608);
and U14773 (N_14773,N_14693,N_14594);
or U14774 (N_14774,N_14678,N_14610);
xor U14775 (N_14775,N_14670,N_14615);
nand U14776 (N_14776,N_14609,N_14591);
and U14777 (N_14777,N_14604,N_14600);
nor U14778 (N_14778,N_14641,N_14683);
or U14779 (N_14779,N_14666,N_14582);
nor U14780 (N_14780,N_14593,N_14627);
nor U14781 (N_14781,N_14630,N_14698);
xnor U14782 (N_14782,N_14667,N_14586);
nand U14783 (N_14783,N_14638,N_14697);
nand U14784 (N_14784,N_14588,N_14690);
xor U14785 (N_14785,N_14616,N_14613);
nand U14786 (N_14786,N_14658,N_14685);
or U14787 (N_14787,N_14566,N_14601);
nand U14788 (N_14788,N_14713,N_14657);
nor U14789 (N_14789,N_14710,N_14564);
xnor U14790 (N_14790,N_14573,N_14584);
xnor U14791 (N_14791,N_14680,N_14679);
or U14792 (N_14792,N_14715,N_14581);
nand U14793 (N_14793,N_14695,N_14631);
and U14794 (N_14794,N_14636,N_14572);
nand U14795 (N_14795,N_14675,N_14640);
nand U14796 (N_14796,N_14577,N_14632);
xor U14797 (N_14797,N_14576,N_14699);
nand U14798 (N_14798,N_14716,N_14655);
xnor U14799 (N_14799,N_14691,N_14626);
nor U14800 (N_14800,N_14677,N_14568);
nand U14801 (N_14801,N_14695,N_14692);
and U14802 (N_14802,N_14655,N_14610);
or U14803 (N_14803,N_14709,N_14602);
or U14804 (N_14804,N_14704,N_14671);
and U14805 (N_14805,N_14563,N_14689);
nand U14806 (N_14806,N_14619,N_14687);
nor U14807 (N_14807,N_14580,N_14614);
or U14808 (N_14808,N_14667,N_14719);
xor U14809 (N_14809,N_14620,N_14605);
and U14810 (N_14810,N_14645,N_14716);
nand U14811 (N_14811,N_14634,N_14615);
and U14812 (N_14812,N_14631,N_14711);
and U14813 (N_14813,N_14658,N_14719);
nand U14814 (N_14814,N_14652,N_14562);
nand U14815 (N_14815,N_14684,N_14643);
or U14816 (N_14816,N_14718,N_14573);
xor U14817 (N_14817,N_14583,N_14669);
and U14818 (N_14818,N_14581,N_14614);
or U14819 (N_14819,N_14619,N_14568);
or U14820 (N_14820,N_14616,N_14599);
or U14821 (N_14821,N_14643,N_14596);
and U14822 (N_14822,N_14591,N_14637);
xor U14823 (N_14823,N_14719,N_14608);
and U14824 (N_14824,N_14707,N_14617);
xor U14825 (N_14825,N_14594,N_14679);
nor U14826 (N_14826,N_14708,N_14699);
xnor U14827 (N_14827,N_14691,N_14635);
nor U14828 (N_14828,N_14583,N_14610);
xor U14829 (N_14829,N_14583,N_14691);
or U14830 (N_14830,N_14703,N_14637);
nand U14831 (N_14831,N_14656,N_14642);
nand U14832 (N_14832,N_14698,N_14667);
nor U14833 (N_14833,N_14648,N_14571);
nor U14834 (N_14834,N_14680,N_14689);
and U14835 (N_14835,N_14580,N_14687);
nor U14836 (N_14836,N_14648,N_14625);
nand U14837 (N_14837,N_14644,N_14623);
nor U14838 (N_14838,N_14597,N_14642);
nand U14839 (N_14839,N_14617,N_14603);
and U14840 (N_14840,N_14612,N_14679);
and U14841 (N_14841,N_14567,N_14668);
xnor U14842 (N_14842,N_14618,N_14600);
nand U14843 (N_14843,N_14666,N_14580);
or U14844 (N_14844,N_14627,N_14687);
or U14845 (N_14845,N_14668,N_14639);
xor U14846 (N_14846,N_14637,N_14600);
and U14847 (N_14847,N_14708,N_14709);
or U14848 (N_14848,N_14632,N_14709);
nand U14849 (N_14849,N_14719,N_14612);
xnor U14850 (N_14850,N_14567,N_14701);
or U14851 (N_14851,N_14587,N_14622);
xnor U14852 (N_14852,N_14612,N_14630);
nand U14853 (N_14853,N_14630,N_14689);
and U14854 (N_14854,N_14699,N_14679);
nand U14855 (N_14855,N_14663,N_14674);
nand U14856 (N_14856,N_14711,N_14600);
and U14857 (N_14857,N_14579,N_14585);
and U14858 (N_14858,N_14700,N_14594);
and U14859 (N_14859,N_14683,N_14598);
and U14860 (N_14860,N_14669,N_14644);
or U14861 (N_14861,N_14613,N_14579);
xor U14862 (N_14862,N_14568,N_14668);
nand U14863 (N_14863,N_14602,N_14566);
and U14864 (N_14864,N_14630,N_14683);
or U14865 (N_14865,N_14660,N_14650);
xor U14866 (N_14866,N_14696,N_14707);
or U14867 (N_14867,N_14564,N_14615);
nand U14868 (N_14868,N_14684,N_14621);
nor U14869 (N_14869,N_14691,N_14699);
nor U14870 (N_14870,N_14702,N_14610);
and U14871 (N_14871,N_14580,N_14699);
or U14872 (N_14872,N_14635,N_14563);
xnor U14873 (N_14873,N_14601,N_14625);
nor U14874 (N_14874,N_14717,N_14634);
xnor U14875 (N_14875,N_14704,N_14686);
and U14876 (N_14876,N_14706,N_14670);
and U14877 (N_14877,N_14628,N_14680);
or U14878 (N_14878,N_14598,N_14603);
nand U14879 (N_14879,N_14594,N_14563);
or U14880 (N_14880,N_14822,N_14730);
or U14881 (N_14881,N_14834,N_14868);
xnor U14882 (N_14882,N_14839,N_14803);
nand U14883 (N_14883,N_14739,N_14720);
xor U14884 (N_14884,N_14737,N_14798);
or U14885 (N_14885,N_14732,N_14761);
and U14886 (N_14886,N_14742,N_14815);
or U14887 (N_14887,N_14725,N_14807);
xnor U14888 (N_14888,N_14800,N_14846);
or U14889 (N_14889,N_14847,N_14759);
nor U14890 (N_14890,N_14872,N_14829);
and U14891 (N_14891,N_14844,N_14769);
nor U14892 (N_14892,N_14767,N_14802);
or U14893 (N_14893,N_14825,N_14875);
nor U14894 (N_14894,N_14797,N_14758);
xnor U14895 (N_14895,N_14853,N_14826);
nand U14896 (N_14896,N_14782,N_14836);
nor U14897 (N_14897,N_14820,N_14848);
xor U14898 (N_14898,N_14787,N_14781);
or U14899 (N_14899,N_14760,N_14775);
nor U14900 (N_14900,N_14762,N_14858);
or U14901 (N_14901,N_14879,N_14786);
nand U14902 (N_14902,N_14840,N_14727);
nand U14903 (N_14903,N_14813,N_14850);
nand U14904 (N_14904,N_14799,N_14766);
or U14905 (N_14905,N_14771,N_14866);
nand U14906 (N_14906,N_14827,N_14744);
and U14907 (N_14907,N_14804,N_14790);
nor U14908 (N_14908,N_14791,N_14755);
nand U14909 (N_14909,N_14877,N_14726);
nor U14910 (N_14910,N_14805,N_14831);
xnor U14911 (N_14911,N_14864,N_14854);
xor U14912 (N_14912,N_14749,N_14862);
nor U14913 (N_14913,N_14723,N_14842);
or U14914 (N_14914,N_14818,N_14838);
nor U14915 (N_14915,N_14777,N_14747);
xor U14916 (N_14916,N_14832,N_14876);
nand U14917 (N_14917,N_14772,N_14874);
nand U14918 (N_14918,N_14764,N_14855);
and U14919 (N_14919,N_14751,N_14823);
nand U14920 (N_14920,N_14752,N_14871);
and U14921 (N_14921,N_14808,N_14809);
nand U14922 (N_14922,N_14765,N_14841);
and U14923 (N_14923,N_14738,N_14722);
nand U14924 (N_14924,N_14878,N_14794);
xor U14925 (N_14925,N_14795,N_14830);
xnor U14926 (N_14926,N_14734,N_14821);
nor U14927 (N_14927,N_14770,N_14861);
and U14928 (N_14928,N_14754,N_14783);
xor U14929 (N_14929,N_14835,N_14793);
and U14930 (N_14930,N_14860,N_14837);
xnor U14931 (N_14931,N_14816,N_14763);
or U14932 (N_14932,N_14768,N_14857);
or U14933 (N_14933,N_14810,N_14788);
xnor U14934 (N_14934,N_14779,N_14869);
or U14935 (N_14935,N_14785,N_14870);
nand U14936 (N_14936,N_14814,N_14819);
xnor U14937 (N_14937,N_14741,N_14773);
nor U14938 (N_14938,N_14867,N_14743);
and U14939 (N_14939,N_14729,N_14774);
xor U14940 (N_14940,N_14828,N_14824);
or U14941 (N_14941,N_14851,N_14792);
and U14942 (N_14942,N_14740,N_14856);
nor U14943 (N_14943,N_14849,N_14756);
or U14944 (N_14944,N_14757,N_14731);
nand U14945 (N_14945,N_14811,N_14778);
nor U14946 (N_14946,N_14859,N_14806);
nand U14947 (N_14947,N_14745,N_14753);
nor U14948 (N_14948,N_14736,N_14746);
xor U14949 (N_14949,N_14817,N_14843);
xor U14950 (N_14950,N_14845,N_14863);
and U14951 (N_14951,N_14776,N_14796);
or U14952 (N_14952,N_14724,N_14750);
nor U14953 (N_14953,N_14852,N_14784);
nor U14954 (N_14954,N_14812,N_14865);
nand U14955 (N_14955,N_14780,N_14748);
or U14956 (N_14956,N_14735,N_14833);
nand U14957 (N_14957,N_14721,N_14789);
or U14958 (N_14958,N_14733,N_14728);
xor U14959 (N_14959,N_14801,N_14873);
or U14960 (N_14960,N_14760,N_14801);
and U14961 (N_14961,N_14735,N_14878);
xor U14962 (N_14962,N_14800,N_14777);
and U14963 (N_14963,N_14808,N_14749);
or U14964 (N_14964,N_14850,N_14828);
and U14965 (N_14965,N_14770,N_14812);
nor U14966 (N_14966,N_14747,N_14845);
and U14967 (N_14967,N_14860,N_14818);
nor U14968 (N_14968,N_14720,N_14813);
nor U14969 (N_14969,N_14861,N_14866);
and U14970 (N_14970,N_14739,N_14829);
or U14971 (N_14971,N_14722,N_14870);
or U14972 (N_14972,N_14872,N_14726);
and U14973 (N_14973,N_14842,N_14853);
and U14974 (N_14974,N_14850,N_14735);
and U14975 (N_14975,N_14729,N_14843);
and U14976 (N_14976,N_14766,N_14878);
nand U14977 (N_14977,N_14758,N_14848);
xor U14978 (N_14978,N_14758,N_14863);
and U14979 (N_14979,N_14873,N_14856);
nand U14980 (N_14980,N_14835,N_14724);
and U14981 (N_14981,N_14771,N_14733);
nand U14982 (N_14982,N_14722,N_14795);
nand U14983 (N_14983,N_14790,N_14834);
nand U14984 (N_14984,N_14750,N_14842);
or U14985 (N_14985,N_14812,N_14814);
or U14986 (N_14986,N_14818,N_14830);
and U14987 (N_14987,N_14747,N_14757);
nand U14988 (N_14988,N_14750,N_14862);
nand U14989 (N_14989,N_14823,N_14721);
or U14990 (N_14990,N_14793,N_14742);
or U14991 (N_14991,N_14829,N_14854);
nand U14992 (N_14992,N_14741,N_14751);
nand U14993 (N_14993,N_14800,N_14841);
nor U14994 (N_14994,N_14806,N_14798);
and U14995 (N_14995,N_14796,N_14800);
nand U14996 (N_14996,N_14809,N_14820);
xor U14997 (N_14997,N_14734,N_14769);
xor U14998 (N_14998,N_14726,N_14788);
or U14999 (N_14999,N_14859,N_14838);
or U15000 (N_15000,N_14835,N_14772);
nand U15001 (N_15001,N_14811,N_14828);
nor U15002 (N_15002,N_14807,N_14820);
nand U15003 (N_15003,N_14852,N_14761);
or U15004 (N_15004,N_14784,N_14847);
nor U15005 (N_15005,N_14793,N_14722);
xor U15006 (N_15006,N_14839,N_14810);
and U15007 (N_15007,N_14852,N_14811);
or U15008 (N_15008,N_14863,N_14735);
nand U15009 (N_15009,N_14849,N_14856);
nor U15010 (N_15010,N_14808,N_14870);
nor U15011 (N_15011,N_14759,N_14762);
nand U15012 (N_15012,N_14796,N_14734);
and U15013 (N_15013,N_14851,N_14774);
xnor U15014 (N_15014,N_14811,N_14834);
xor U15015 (N_15015,N_14770,N_14856);
xnor U15016 (N_15016,N_14870,N_14806);
xor U15017 (N_15017,N_14759,N_14734);
xnor U15018 (N_15018,N_14738,N_14844);
or U15019 (N_15019,N_14773,N_14864);
nand U15020 (N_15020,N_14724,N_14766);
nor U15021 (N_15021,N_14818,N_14753);
nand U15022 (N_15022,N_14721,N_14775);
nand U15023 (N_15023,N_14867,N_14795);
xor U15024 (N_15024,N_14737,N_14770);
xor U15025 (N_15025,N_14830,N_14846);
nor U15026 (N_15026,N_14851,N_14823);
and U15027 (N_15027,N_14829,N_14823);
nor U15028 (N_15028,N_14821,N_14847);
nor U15029 (N_15029,N_14822,N_14732);
nor U15030 (N_15030,N_14862,N_14855);
and U15031 (N_15031,N_14817,N_14782);
nor U15032 (N_15032,N_14847,N_14774);
nor U15033 (N_15033,N_14847,N_14787);
and U15034 (N_15034,N_14759,N_14763);
and U15035 (N_15035,N_14860,N_14805);
nand U15036 (N_15036,N_14830,N_14822);
nand U15037 (N_15037,N_14807,N_14784);
or U15038 (N_15038,N_14809,N_14798);
nand U15039 (N_15039,N_14805,N_14788);
xnor U15040 (N_15040,N_14991,N_14894);
xor U15041 (N_15041,N_14929,N_14911);
nor U15042 (N_15042,N_14950,N_15007);
nor U15043 (N_15043,N_15008,N_14931);
xor U15044 (N_15044,N_14985,N_15032);
nand U15045 (N_15045,N_14917,N_14883);
or U15046 (N_15046,N_14912,N_14885);
xnor U15047 (N_15047,N_14969,N_14952);
nand U15048 (N_15048,N_15006,N_15029);
nand U15049 (N_15049,N_15017,N_14891);
and U15050 (N_15050,N_14986,N_15019);
and U15051 (N_15051,N_14893,N_14998);
xor U15052 (N_15052,N_14930,N_14909);
xor U15053 (N_15053,N_14993,N_14996);
and U15054 (N_15054,N_14890,N_14895);
nand U15055 (N_15055,N_15035,N_14916);
xnor U15056 (N_15056,N_14980,N_14901);
nand U15057 (N_15057,N_14960,N_14948);
xor U15058 (N_15058,N_14937,N_14935);
xor U15059 (N_15059,N_15026,N_14896);
nand U15060 (N_15060,N_14926,N_14997);
xnor U15061 (N_15061,N_15001,N_14943);
nor U15062 (N_15062,N_14978,N_14964);
nor U15063 (N_15063,N_14915,N_14961);
xnor U15064 (N_15064,N_14983,N_15030);
or U15065 (N_15065,N_14965,N_14975);
or U15066 (N_15066,N_15004,N_14908);
or U15067 (N_15067,N_14966,N_14941);
and U15068 (N_15068,N_14962,N_15028);
nand U15069 (N_15069,N_15011,N_14899);
nand U15070 (N_15070,N_15039,N_14987);
nor U15071 (N_15071,N_15027,N_14944);
or U15072 (N_15072,N_14914,N_14971);
and U15073 (N_15073,N_14992,N_14927);
nor U15074 (N_15074,N_15033,N_15037);
or U15075 (N_15075,N_15013,N_14936);
or U15076 (N_15076,N_14967,N_14902);
nand U15077 (N_15077,N_14880,N_15021);
nor U15078 (N_15078,N_14898,N_14981);
xnor U15079 (N_15079,N_14897,N_14953);
or U15080 (N_15080,N_14979,N_14954);
and U15081 (N_15081,N_14945,N_14949);
or U15082 (N_15082,N_14918,N_15016);
and U15083 (N_15083,N_14900,N_14892);
nor U15084 (N_15084,N_14984,N_14976);
nor U15085 (N_15085,N_14888,N_14990);
or U15086 (N_15086,N_15024,N_14963);
nand U15087 (N_15087,N_15000,N_14940);
or U15088 (N_15088,N_15038,N_14939);
nor U15089 (N_15089,N_14958,N_14995);
or U15090 (N_15090,N_14913,N_14955);
nor U15091 (N_15091,N_14928,N_15018);
or U15092 (N_15092,N_14972,N_14881);
xor U15093 (N_15093,N_14977,N_14942);
nand U15094 (N_15094,N_15014,N_14994);
nor U15095 (N_15095,N_15036,N_15023);
and U15096 (N_15096,N_14933,N_15009);
nand U15097 (N_15097,N_15015,N_15031);
or U15098 (N_15098,N_15012,N_14886);
or U15099 (N_15099,N_15003,N_14921);
xor U15100 (N_15100,N_14910,N_15022);
nor U15101 (N_15101,N_14947,N_15005);
nor U15102 (N_15102,N_15020,N_14925);
or U15103 (N_15103,N_15025,N_14934);
nor U15104 (N_15104,N_14932,N_14924);
nand U15105 (N_15105,N_14904,N_14905);
xor U15106 (N_15106,N_14919,N_14906);
nor U15107 (N_15107,N_14988,N_14922);
xnor U15108 (N_15108,N_14887,N_14968);
or U15109 (N_15109,N_14957,N_14956);
xor U15110 (N_15110,N_14974,N_14920);
xor U15111 (N_15111,N_15002,N_14999);
nor U15112 (N_15112,N_15010,N_14959);
xnor U15113 (N_15113,N_14982,N_14938);
or U15114 (N_15114,N_14923,N_14946);
or U15115 (N_15115,N_14970,N_14907);
nor U15116 (N_15116,N_15034,N_14903);
and U15117 (N_15117,N_14882,N_14951);
xnor U15118 (N_15118,N_14884,N_14889);
or U15119 (N_15119,N_14989,N_14973);
nand U15120 (N_15120,N_14905,N_14968);
or U15121 (N_15121,N_14989,N_14899);
nor U15122 (N_15122,N_15033,N_14913);
or U15123 (N_15123,N_15016,N_15023);
nand U15124 (N_15124,N_14891,N_14912);
and U15125 (N_15125,N_15033,N_15011);
nor U15126 (N_15126,N_14933,N_15032);
nor U15127 (N_15127,N_14968,N_14977);
nor U15128 (N_15128,N_14915,N_15009);
or U15129 (N_15129,N_14895,N_14989);
or U15130 (N_15130,N_15011,N_14892);
and U15131 (N_15131,N_14940,N_14923);
and U15132 (N_15132,N_14988,N_15037);
xor U15133 (N_15133,N_14940,N_14930);
xnor U15134 (N_15134,N_14980,N_14893);
nor U15135 (N_15135,N_14927,N_14983);
and U15136 (N_15136,N_14907,N_15033);
or U15137 (N_15137,N_14996,N_14963);
nor U15138 (N_15138,N_15003,N_14982);
xor U15139 (N_15139,N_14984,N_14951);
nor U15140 (N_15140,N_14967,N_14974);
xor U15141 (N_15141,N_15011,N_15022);
nand U15142 (N_15142,N_14915,N_14980);
or U15143 (N_15143,N_14914,N_14935);
nand U15144 (N_15144,N_14966,N_14919);
and U15145 (N_15145,N_14998,N_14971);
and U15146 (N_15146,N_15026,N_14965);
or U15147 (N_15147,N_14964,N_14923);
or U15148 (N_15148,N_14998,N_14912);
or U15149 (N_15149,N_15006,N_14945);
xnor U15150 (N_15150,N_15005,N_14992);
and U15151 (N_15151,N_14907,N_14931);
xor U15152 (N_15152,N_14910,N_14925);
nand U15153 (N_15153,N_15031,N_14944);
or U15154 (N_15154,N_14895,N_15004);
nand U15155 (N_15155,N_15034,N_15019);
and U15156 (N_15156,N_14929,N_14902);
or U15157 (N_15157,N_14966,N_15006);
xor U15158 (N_15158,N_14988,N_14934);
xor U15159 (N_15159,N_14903,N_15033);
nand U15160 (N_15160,N_14902,N_15006);
and U15161 (N_15161,N_15033,N_14885);
xnor U15162 (N_15162,N_15001,N_14987);
nor U15163 (N_15163,N_14888,N_15012);
xnor U15164 (N_15164,N_14967,N_14887);
xor U15165 (N_15165,N_15024,N_14967);
or U15166 (N_15166,N_14908,N_14961);
and U15167 (N_15167,N_14976,N_14905);
xor U15168 (N_15168,N_14888,N_15025);
xor U15169 (N_15169,N_14886,N_15009);
or U15170 (N_15170,N_14884,N_15036);
nor U15171 (N_15171,N_14907,N_14973);
or U15172 (N_15172,N_15011,N_14984);
and U15173 (N_15173,N_14937,N_14925);
xor U15174 (N_15174,N_14889,N_15037);
or U15175 (N_15175,N_14975,N_14962);
or U15176 (N_15176,N_15038,N_14970);
xor U15177 (N_15177,N_14925,N_14915);
nor U15178 (N_15178,N_14996,N_14887);
nor U15179 (N_15179,N_14892,N_14971);
nand U15180 (N_15180,N_14961,N_14970);
nand U15181 (N_15181,N_14947,N_14938);
nor U15182 (N_15182,N_14946,N_14935);
and U15183 (N_15183,N_14931,N_14896);
and U15184 (N_15184,N_15001,N_14917);
xor U15185 (N_15185,N_14941,N_14937);
xnor U15186 (N_15186,N_14880,N_14997);
xnor U15187 (N_15187,N_15012,N_15007);
and U15188 (N_15188,N_14881,N_14982);
and U15189 (N_15189,N_14943,N_15028);
or U15190 (N_15190,N_14888,N_15018);
or U15191 (N_15191,N_15008,N_14989);
or U15192 (N_15192,N_15019,N_14898);
or U15193 (N_15193,N_14983,N_15018);
nand U15194 (N_15194,N_14921,N_14915);
or U15195 (N_15195,N_14882,N_15015);
or U15196 (N_15196,N_15016,N_15033);
and U15197 (N_15197,N_15004,N_14960);
xnor U15198 (N_15198,N_14980,N_14939);
nand U15199 (N_15199,N_14896,N_14951);
nor U15200 (N_15200,N_15105,N_15075);
and U15201 (N_15201,N_15117,N_15166);
nand U15202 (N_15202,N_15090,N_15148);
and U15203 (N_15203,N_15132,N_15174);
nand U15204 (N_15204,N_15058,N_15144);
nand U15205 (N_15205,N_15164,N_15165);
and U15206 (N_15206,N_15103,N_15096);
xor U15207 (N_15207,N_15068,N_15178);
nor U15208 (N_15208,N_15053,N_15170);
nor U15209 (N_15209,N_15089,N_15094);
nand U15210 (N_15210,N_15176,N_15142);
and U15211 (N_15211,N_15040,N_15121);
nand U15212 (N_15212,N_15085,N_15106);
nor U15213 (N_15213,N_15061,N_15043);
xor U15214 (N_15214,N_15155,N_15059);
nor U15215 (N_15215,N_15168,N_15189);
nor U15216 (N_15216,N_15050,N_15151);
or U15217 (N_15217,N_15112,N_15084);
and U15218 (N_15218,N_15041,N_15196);
xnor U15219 (N_15219,N_15129,N_15153);
nand U15220 (N_15220,N_15047,N_15093);
nand U15221 (N_15221,N_15192,N_15123);
nor U15222 (N_15222,N_15104,N_15197);
nor U15223 (N_15223,N_15167,N_15137);
and U15224 (N_15224,N_15115,N_15131);
xnor U15225 (N_15225,N_15118,N_15126);
or U15226 (N_15226,N_15172,N_15180);
nand U15227 (N_15227,N_15150,N_15071);
nand U15228 (N_15228,N_15177,N_15149);
nand U15229 (N_15229,N_15091,N_15154);
nand U15230 (N_15230,N_15152,N_15077);
or U15231 (N_15231,N_15046,N_15179);
and U15232 (N_15232,N_15169,N_15067);
or U15233 (N_15233,N_15147,N_15175);
nor U15234 (N_15234,N_15109,N_15082);
xnor U15235 (N_15235,N_15156,N_15124);
and U15236 (N_15236,N_15160,N_15199);
or U15237 (N_15237,N_15119,N_15145);
nand U15238 (N_15238,N_15055,N_15183);
xor U15239 (N_15239,N_15069,N_15057);
and U15240 (N_15240,N_15136,N_15140);
and U15241 (N_15241,N_15107,N_15101);
xor U15242 (N_15242,N_15079,N_15161);
and U15243 (N_15243,N_15044,N_15120);
or U15244 (N_15244,N_15081,N_15100);
and U15245 (N_15245,N_15135,N_15193);
or U15246 (N_15246,N_15056,N_15128);
and U15247 (N_15247,N_15143,N_15116);
nor U15248 (N_15248,N_15064,N_15083);
xor U15249 (N_15249,N_15073,N_15098);
and U15250 (N_15250,N_15163,N_15045);
nor U15251 (N_15251,N_15042,N_15185);
or U15252 (N_15252,N_15191,N_15078);
and U15253 (N_15253,N_15051,N_15099);
nand U15254 (N_15254,N_15111,N_15188);
nor U15255 (N_15255,N_15122,N_15066);
xnor U15256 (N_15256,N_15072,N_15171);
and U15257 (N_15257,N_15141,N_15097);
xnor U15258 (N_15258,N_15074,N_15062);
or U15259 (N_15259,N_15070,N_15146);
or U15260 (N_15260,N_15125,N_15048);
or U15261 (N_15261,N_15173,N_15186);
nor U15262 (N_15262,N_15133,N_15054);
nand U15263 (N_15263,N_15108,N_15114);
nor U15264 (N_15264,N_15065,N_15158);
nor U15265 (N_15265,N_15157,N_15110);
or U15266 (N_15266,N_15187,N_15162);
or U15267 (N_15267,N_15086,N_15060);
xnor U15268 (N_15268,N_15127,N_15134);
nand U15269 (N_15269,N_15194,N_15088);
nand U15270 (N_15270,N_15195,N_15095);
nor U15271 (N_15271,N_15102,N_15159);
xor U15272 (N_15272,N_15139,N_15092);
nor U15273 (N_15273,N_15190,N_15049);
nand U15274 (N_15274,N_15181,N_15184);
or U15275 (N_15275,N_15063,N_15087);
nor U15276 (N_15276,N_15080,N_15113);
or U15277 (N_15277,N_15182,N_15130);
xor U15278 (N_15278,N_15198,N_15076);
xnor U15279 (N_15279,N_15138,N_15052);
or U15280 (N_15280,N_15072,N_15063);
nand U15281 (N_15281,N_15093,N_15107);
nor U15282 (N_15282,N_15122,N_15186);
nand U15283 (N_15283,N_15128,N_15043);
nand U15284 (N_15284,N_15182,N_15195);
nand U15285 (N_15285,N_15184,N_15048);
or U15286 (N_15286,N_15175,N_15090);
xnor U15287 (N_15287,N_15091,N_15113);
xor U15288 (N_15288,N_15064,N_15197);
or U15289 (N_15289,N_15088,N_15179);
or U15290 (N_15290,N_15197,N_15056);
xnor U15291 (N_15291,N_15143,N_15154);
and U15292 (N_15292,N_15114,N_15132);
xnor U15293 (N_15293,N_15055,N_15046);
and U15294 (N_15294,N_15089,N_15139);
and U15295 (N_15295,N_15148,N_15143);
xor U15296 (N_15296,N_15190,N_15125);
nor U15297 (N_15297,N_15175,N_15103);
nor U15298 (N_15298,N_15118,N_15150);
xor U15299 (N_15299,N_15082,N_15089);
nor U15300 (N_15300,N_15061,N_15153);
or U15301 (N_15301,N_15116,N_15144);
or U15302 (N_15302,N_15085,N_15168);
or U15303 (N_15303,N_15126,N_15158);
nand U15304 (N_15304,N_15044,N_15127);
nand U15305 (N_15305,N_15081,N_15062);
or U15306 (N_15306,N_15146,N_15077);
and U15307 (N_15307,N_15131,N_15175);
xnor U15308 (N_15308,N_15171,N_15107);
nand U15309 (N_15309,N_15132,N_15044);
nand U15310 (N_15310,N_15142,N_15185);
xor U15311 (N_15311,N_15073,N_15086);
xnor U15312 (N_15312,N_15104,N_15043);
or U15313 (N_15313,N_15191,N_15168);
nor U15314 (N_15314,N_15116,N_15147);
xor U15315 (N_15315,N_15165,N_15075);
or U15316 (N_15316,N_15081,N_15192);
or U15317 (N_15317,N_15041,N_15073);
or U15318 (N_15318,N_15075,N_15100);
and U15319 (N_15319,N_15118,N_15155);
or U15320 (N_15320,N_15145,N_15199);
and U15321 (N_15321,N_15047,N_15112);
or U15322 (N_15322,N_15063,N_15190);
nand U15323 (N_15323,N_15085,N_15100);
nand U15324 (N_15324,N_15157,N_15107);
or U15325 (N_15325,N_15097,N_15148);
xnor U15326 (N_15326,N_15132,N_15081);
nor U15327 (N_15327,N_15076,N_15064);
or U15328 (N_15328,N_15118,N_15152);
nor U15329 (N_15329,N_15193,N_15164);
xnor U15330 (N_15330,N_15067,N_15093);
nor U15331 (N_15331,N_15140,N_15069);
xnor U15332 (N_15332,N_15119,N_15154);
or U15333 (N_15333,N_15165,N_15179);
nand U15334 (N_15334,N_15161,N_15154);
or U15335 (N_15335,N_15071,N_15180);
nand U15336 (N_15336,N_15183,N_15124);
or U15337 (N_15337,N_15080,N_15063);
nor U15338 (N_15338,N_15129,N_15052);
nor U15339 (N_15339,N_15045,N_15048);
xnor U15340 (N_15340,N_15151,N_15074);
or U15341 (N_15341,N_15110,N_15145);
nor U15342 (N_15342,N_15066,N_15052);
or U15343 (N_15343,N_15104,N_15064);
or U15344 (N_15344,N_15099,N_15152);
or U15345 (N_15345,N_15158,N_15181);
and U15346 (N_15346,N_15105,N_15137);
xnor U15347 (N_15347,N_15100,N_15186);
nor U15348 (N_15348,N_15165,N_15070);
and U15349 (N_15349,N_15176,N_15188);
xor U15350 (N_15350,N_15177,N_15196);
nor U15351 (N_15351,N_15135,N_15148);
nor U15352 (N_15352,N_15059,N_15041);
nand U15353 (N_15353,N_15075,N_15166);
nand U15354 (N_15354,N_15083,N_15162);
nor U15355 (N_15355,N_15059,N_15114);
nand U15356 (N_15356,N_15096,N_15157);
nand U15357 (N_15357,N_15180,N_15198);
or U15358 (N_15358,N_15146,N_15195);
nand U15359 (N_15359,N_15063,N_15156);
and U15360 (N_15360,N_15325,N_15259);
nand U15361 (N_15361,N_15237,N_15229);
xnor U15362 (N_15362,N_15293,N_15222);
nor U15363 (N_15363,N_15249,N_15320);
or U15364 (N_15364,N_15315,N_15269);
and U15365 (N_15365,N_15221,N_15228);
or U15366 (N_15366,N_15236,N_15232);
nand U15367 (N_15367,N_15209,N_15213);
nand U15368 (N_15368,N_15234,N_15220);
or U15369 (N_15369,N_15336,N_15214);
xor U15370 (N_15370,N_15289,N_15309);
nand U15371 (N_15371,N_15287,N_15201);
or U15372 (N_15372,N_15271,N_15273);
and U15373 (N_15373,N_15233,N_15266);
nand U15374 (N_15374,N_15255,N_15218);
xor U15375 (N_15375,N_15301,N_15351);
nor U15376 (N_15376,N_15247,N_15323);
nand U15377 (N_15377,N_15313,N_15311);
and U15378 (N_15378,N_15205,N_15217);
and U15379 (N_15379,N_15272,N_15203);
and U15380 (N_15380,N_15330,N_15308);
and U15381 (N_15381,N_15256,N_15244);
or U15382 (N_15382,N_15341,N_15202);
and U15383 (N_15383,N_15302,N_15200);
and U15384 (N_15384,N_15265,N_15274);
and U15385 (N_15385,N_15243,N_15204);
and U15386 (N_15386,N_15300,N_15291);
nand U15387 (N_15387,N_15253,N_15270);
xnor U15388 (N_15388,N_15230,N_15354);
nand U15389 (N_15389,N_15344,N_15292);
nor U15390 (N_15390,N_15339,N_15208);
and U15391 (N_15391,N_15285,N_15355);
or U15392 (N_15392,N_15248,N_15215);
nand U15393 (N_15393,N_15261,N_15326);
xor U15394 (N_15394,N_15210,N_15304);
nor U15395 (N_15395,N_15334,N_15267);
nand U15396 (N_15396,N_15345,N_15312);
and U15397 (N_15397,N_15216,N_15257);
or U15398 (N_15398,N_15246,N_15239);
xor U15399 (N_15399,N_15278,N_15240);
nor U15400 (N_15400,N_15321,N_15329);
nand U15401 (N_15401,N_15348,N_15262);
xnor U15402 (N_15402,N_15280,N_15242);
nand U15403 (N_15403,N_15324,N_15296);
or U15404 (N_15404,N_15207,N_15338);
nand U15405 (N_15405,N_15317,N_15241);
and U15406 (N_15406,N_15305,N_15277);
and U15407 (N_15407,N_15254,N_15314);
xor U15408 (N_15408,N_15286,N_15328);
nand U15409 (N_15409,N_15316,N_15288);
and U15410 (N_15410,N_15297,N_15342);
or U15411 (N_15411,N_15251,N_15306);
and U15412 (N_15412,N_15276,N_15332);
xor U15413 (N_15413,N_15211,N_15282);
nor U15414 (N_15414,N_15357,N_15319);
or U15415 (N_15415,N_15263,N_15327);
and U15416 (N_15416,N_15250,N_15260);
nand U15417 (N_15417,N_15235,N_15223);
nand U15418 (N_15418,N_15331,N_15227);
nand U15419 (N_15419,N_15347,N_15343);
nor U15420 (N_15420,N_15281,N_15352);
nor U15421 (N_15421,N_15358,N_15283);
xor U15422 (N_15422,N_15219,N_15346);
xor U15423 (N_15423,N_15303,N_15206);
nor U15424 (N_15424,N_15295,N_15298);
and U15425 (N_15425,N_15353,N_15275);
xor U15426 (N_15426,N_15225,N_15284);
nor U15427 (N_15427,N_15279,N_15337);
and U15428 (N_15428,N_15294,N_15224);
or U15429 (N_15429,N_15340,N_15350);
nor U15430 (N_15430,N_15252,N_15356);
nor U15431 (N_15431,N_15290,N_15310);
xnor U15432 (N_15432,N_15318,N_15231);
nor U15433 (N_15433,N_15238,N_15268);
nor U15434 (N_15434,N_15264,N_15245);
or U15435 (N_15435,N_15307,N_15258);
xnor U15436 (N_15436,N_15299,N_15333);
and U15437 (N_15437,N_15349,N_15212);
nand U15438 (N_15438,N_15226,N_15359);
nor U15439 (N_15439,N_15335,N_15322);
nand U15440 (N_15440,N_15238,N_15241);
or U15441 (N_15441,N_15219,N_15270);
nand U15442 (N_15442,N_15334,N_15307);
nor U15443 (N_15443,N_15204,N_15344);
xnor U15444 (N_15444,N_15327,N_15249);
nor U15445 (N_15445,N_15214,N_15306);
nand U15446 (N_15446,N_15352,N_15253);
or U15447 (N_15447,N_15234,N_15296);
and U15448 (N_15448,N_15262,N_15247);
and U15449 (N_15449,N_15324,N_15220);
nor U15450 (N_15450,N_15206,N_15248);
nand U15451 (N_15451,N_15349,N_15233);
and U15452 (N_15452,N_15277,N_15339);
or U15453 (N_15453,N_15211,N_15243);
xor U15454 (N_15454,N_15261,N_15257);
or U15455 (N_15455,N_15321,N_15264);
or U15456 (N_15456,N_15314,N_15234);
and U15457 (N_15457,N_15222,N_15257);
nor U15458 (N_15458,N_15332,N_15311);
nand U15459 (N_15459,N_15269,N_15332);
nor U15460 (N_15460,N_15334,N_15306);
nand U15461 (N_15461,N_15264,N_15200);
nand U15462 (N_15462,N_15260,N_15219);
xor U15463 (N_15463,N_15296,N_15337);
or U15464 (N_15464,N_15289,N_15222);
nand U15465 (N_15465,N_15316,N_15208);
nand U15466 (N_15466,N_15240,N_15353);
nand U15467 (N_15467,N_15316,N_15346);
nand U15468 (N_15468,N_15280,N_15327);
nor U15469 (N_15469,N_15251,N_15272);
nand U15470 (N_15470,N_15234,N_15233);
nand U15471 (N_15471,N_15273,N_15267);
or U15472 (N_15472,N_15204,N_15265);
and U15473 (N_15473,N_15308,N_15206);
nor U15474 (N_15474,N_15349,N_15273);
and U15475 (N_15475,N_15327,N_15242);
xor U15476 (N_15476,N_15293,N_15289);
and U15477 (N_15477,N_15240,N_15299);
nor U15478 (N_15478,N_15213,N_15217);
nand U15479 (N_15479,N_15207,N_15322);
and U15480 (N_15480,N_15245,N_15356);
nor U15481 (N_15481,N_15216,N_15303);
and U15482 (N_15482,N_15287,N_15226);
xor U15483 (N_15483,N_15254,N_15309);
xnor U15484 (N_15484,N_15267,N_15250);
nand U15485 (N_15485,N_15225,N_15234);
or U15486 (N_15486,N_15295,N_15320);
nand U15487 (N_15487,N_15338,N_15211);
nor U15488 (N_15488,N_15346,N_15294);
or U15489 (N_15489,N_15289,N_15242);
or U15490 (N_15490,N_15292,N_15351);
xor U15491 (N_15491,N_15209,N_15246);
nand U15492 (N_15492,N_15313,N_15316);
xnor U15493 (N_15493,N_15350,N_15330);
xor U15494 (N_15494,N_15263,N_15344);
xnor U15495 (N_15495,N_15348,N_15359);
nand U15496 (N_15496,N_15232,N_15290);
or U15497 (N_15497,N_15268,N_15212);
xor U15498 (N_15498,N_15257,N_15345);
and U15499 (N_15499,N_15238,N_15209);
xnor U15500 (N_15500,N_15324,N_15314);
nor U15501 (N_15501,N_15326,N_15288);
or U15502 (N_15502,N_15299,N_15311);
and U15503 (N_15503,N_15296,N_15352);
and U15504 (N_15504,N_15203,N_15283);
nor U15505 (N_15505,N_15223,N_15222);
or U15506 (N_15506,N_15329,N_15252);
nor U15507 (N_15507,N_15200,N_15323);
nand U15508 (N_15508,N_15353,N_15209);
xnor U15509 (N_15509,N_15336,N_15219);
xor U15510 (N_15510,N_15336,N_15273);
nor U15511 (N_15511,N_15222,N_15292);
nand U15512 (N_15512,N_15240,N_15220);
nor U15513 (N_15513,N_15331,N_15297);
nand U15514 (N_15514,N_15305,N_15230);
and U15515 (N_15515,N_15284,N_15233);
and U15516 (N_15516,N_15284,N_15290);
nor U15517 (N_15517,N_15206,N_15230);
and U15518 (N_15518,N_15270,N_15328);
and U15519 (N_15519,N_15331,N_15288);
and U15520 (N_15520,N_15391,N_15443);
nor U15521 (N_15521,N_15505,N_15510);
or U15522 (N_15522,N_15401,N_15430);
and U15523 (N_15523,N_15461,N_15479);
and U15524 (N_15524,N_15440,N_15385);
and U15525 (N_15525,N_15498,N_15394);
and U15526 (N_15526,N_15400,N_15519);
xnor U15527 (N_15527,N_15449,N_15492);
or U15528 (N_15528,N_15513,N_15414);
and U15529 (N_15529,N_15480,N_15428);
and U15530 (N_15530,N_15433,N_15368);
or U15531 (N_15531,N_15422,N_15420);
and U15532 (N_15532,N_15495,N_15389);
xnor U15533 (N_15533,N_15388,N_15484);
nor U15534 (N_15534,N_15506,N_15518);
and U15535 (N_15535,N_15502,N_15407);
or U15536 (N_15536,N_15489,N_15413);
xnor U15537 (N_15537,N_15517,N_15462);
or U15538 (N_15538,N_15367,N_15460);
and U15539 (N_15539,N_15438,N_15486);
nor U15540 (N_15540,N_15364,N_15437);
xnor U15541 (N_15541,N_15474,N_15471);
nor U15542 (N_15542,N_15415,N_15403);
nor U15543 (N_15543,N_15468,N_15393);
xnor U15544 (N_15544,N_15514,N_15507);
xnor U15545 (N_15545,N_15416,N_15465);
nor U15546 (N_15546,N_15483,N_15496);
or U15547 (N_15547,N_15423,N_15365);
nand U15548 (N_15548,N_15378,N_15409);
nand U15549 (N_15549,N_15490,N_15379);
xor U15550 (N_15550,N_15504,N_15412);
xnor U15551 (N_15551,N_15424,N_15361);
xor U15552 (N_15552,N_15360,N_15397);
and U15553 (N_15553,N_15398,N_15493);
nand U15554 (N_15554,N_15408,N_15478);
nand U15555 (N_15555,N_15451,N_15464);
nand U15556 (N_15556,N_15473,N_15395);
and U15557 (N_15557,N_15452,N_15445);
nor U15558 (N_15558,N_15441,N_15421);
nand U15559 (N_15559,N_15472,N_15491);
nand U15560 (N_15560,N_15463,N_15444);
nor U15561 (N_15561,N_15466,N_15384);
nand U15562 (N_15562,N_15455,N_15417);
nand U15563 (N_15563,N_15362,N_15481);
and U15564 (N_15564,N_15431,N_15516);
and U15565 (N_15565,N_15371,N_15439);
or U15566 (N_15566,N_15501,N_15456);
or U15567 (N_15567,N_15442,N_15488);
and U15568 (N_15568,N_15381,N_15467);
nor U15569 (N_15569,N_15429,N_15508);
or U15570 (N_15570,N_15503,N_15447);
nand U15571 (N_15571,N_15425,N_15454);
or U15572 (N_15572,N_15386,N_15448);
or U15573 (N_15573,N_15427,N_15457);
and U15574 (N_15574,N_15375,N_15459);
nor U15575 (N_15575,N_15511,N_15377);
nand U15576 (N_15576,N_15476,N_15515);
and U15577 (N_15577,N_15434,N_15366);
nor U15578 (N_15578,N_15494,N_15392);
and U15579 (N_15579,N_15399,N_15453);
xnor U15580 (N_15580,N_15369,N_15419);
xor U15581 (N_15581,N_15475,N_15432);
and U15582 (N_15582,N_15482,N_15387);
and U15583 (N_15583,N_15382,N_15512);
and U15584 (N_15584,N_15450,N_15370);
nand U15585 (N_15585,N_15373,N_15372);
and U15586 (N_15586,N_15405,N_15497);
nor U15587 (N_15587,N_15470,N_15390);
xor U15588 (N_15588,N_15499,N_15500);
or U15589 (N_15589,N_15404,N_15487);
nand U15590 (N_15590,N_15509,N_15418);
nand U15591 (N_15591,N_15396,N_15383);
and U15592 (N_15592,N_15426,N_15485);
nor U15593 (N_15593,N_15435,N_15469);
nand U15594 (N_15594,N_15406,N_15410);
nor U15595 (N_15595,N_15436,N_15446);
nand U15596 (N_15596,N_15363,N_15402);
nor U15597 (N_15597,N_15458,N_15411);
nor U15598 (N_15598,N_15477,N_15376);
nor U15599 (N_15599,N_15374,N_15380);
xnor U15600 (N_15600,N_15397,N_15457);
xnor U15601 (N_15601,N_15408,N_15449);
nand U15602 (N_15602,N_15429,N_15473);
nand U15603 (N_15603,N_15511,N_15498);
nor U15604 (N_15604,N_15378,N_15463);
xnor U15605 (N_15605,N_15444,N_15494);
nor U15606 (N_15606,N_15405,N_15421);
or U15607 (N_15607,N_15433,N_15482);
nor U15608 (N_15608,N_15386,N_15434);
nor U15609 (N_15609,N_15460,N_15399);
and U15610 (N_15610,N_15463,N_15383);
nor U15611 (N_15611,N_15487,N_15466);
nand U15612 (N_15612,N_15383,N_15447);
nor U15613 (N_15613,N_15365,N_15491);
nor U15614 (N_15614,N_15478,N_15409);
and U15615 (N_15615,N_15436,N_15371);
and U15616 (N_15616,N_15430,N_15428);
nand U15617 (N_15617,N_15513,N_15500);
nor U15618 (N_15618,N_15492,N_15460);
nand U15619 (N_15619,N_15440,N_15518);
or U15620 (N_15620,N_15361,N_15510);
and U15621 (N_15621,N_15376,N_15431);
xnor U15622 (N_15622,N_15360,N_15441);
or U15623 (N_15623,N_15506,N_15437);
or U15624 (N_15624,N_15480,N_15450);
xnor U15625 (N_15625,N_15475,N_15372);
nand U15626 (N_15626,N_15487,N_15403);
nor U15627 (N_15627,N_15367,N_15432);
xnor U15628 (N_15628,N_15454,N_15371);
nor U15629 (N_15629,N_15451,N_15448);
nor U15630 (N_15630,N_15476,N_15462);
nand U15631 (N_15631,N_15378,N_15466);
nand U15632 (N_15632,N_15497,N_15392);
xor U15633 (N_15633,N_15372,N_15411);
nand U15634 (N_15634,N_15477,N_15469);
or U15635 (N_15635,N_15457,N_15461);
xor U15636 (N_15636,N_15431,N_15502);
and U15637 (N_15637,N_15488,N_15435);
or U15638 (N_15638,N_15432,N_15409);
and U15639 (N_15639,N_15481,N_15510);
xor U15640 (N_15640,N_15454,N_15512);
nand U15641 (N_15641,N_15390,N_15448);
xnor U15642 (N_15642,N_15510,N_15471);
and U15643 (N_15643,N_15403,N_15511);
or U15644 (N_15644,N_15432,N_15407);
nor U15645 (N_15645,N_15375,N_15367);
xnor U15646 (N_15646,N_15377,N_15435);
xor U15647 (N_15647,N_15496,N_15392);
or U15648 (N_15648,N_15444,N_15466);
and U15649 (N_15649,N_15459,N_15367);
xor U15650 (N_15650,N_15417,N_15423);
xor U15651 (N_15651,N_15367,N_15456);
and U15652 (N_15652,N_15481,N_15370);
nor U15653 (N_15653,N_15463,N_15492);
or U15654 (N_15654,N_15480,N_15444);
nor U15655 (N_15655,N_15416,N_15436);
nor U15656 (N_15656,N_15408,N_15391);
nand U15657 (N_15657,N_15505,N_15386);
nand U15658 (N_15658,N_15413,N_15479);
nand U15659 (N_15659,N_15492,N_15455);
or U15660 (N_15660,N_15456,N_15450);
or U15661 (N_15661,N_15442,N_15380);
and U15662 (N_15662,N_15379,N_15415);
or U15663 (N_15663,N_15480,N_15461);
and U15664 (N_15664,N_15411,N_15361);
nand U15665 (N_15665,N_15410,N_15460);
nand U15666 (N_15666,N_15407,N_15394);
xor U15667 (N_15667,N_15504,N_15413);
and U15668 (N_15668,N_15503,N_15392);
nand U15669 (N_15669,N_15516,N_15491);
or U15670 (N_15670,N_15374,N_15412);
nor U15671 (N_15671,N_15362,N_15499);
nor U15672 (N_15672,N_15454,N_15517);
or U15673 (N_15673,N_15420,N_15405);
and U15674 (N_15674,N_15498,N_15409);
nor U15675 (N_15675,N_15410,N_15372);
nand U15676 (N_15676,N_15468,N_15450);
nand U15677 (N_15677,N_15452,N_15466);
nand U15678 (N_15678,N_15401,N_15416);
or U15679 (N_15679,N_15413,N_15465);
xor U15680 (N_15680,N_15568,N_15637);
or U15681 (N_15681,N_15592,N_15638);
nor U15682 (N_15682,N_15547,N_15653);
and U15683 (N_15683,N_15650,N_15675);
nand U15684 (N_15684,N_15591,N_15600);
nand U15685 (N_15685,N_15548,N_15564);
and U15686 (N_15686,N_15627,N_15562);
xnor U15687 (N_15687,N_15558,N_15586);
nand U15688 (N_15688,N_15556,N_15538);
nand U15689 (N_15689,N_15559,N_15595);
nor U15690 (N_15690,N_15671,N_15601);
or U15691 (N_15691,N_15529,N_15636);
or U15692 (N_15692,N_15525,N_15677);
nand U15693 (N_15693,N_15664,N_15521);
or U15694 (N_15694,N_15649,N_15641);
and U15695 (N_15695,N_15615,N_15554);
xnor U15696 (N_15696,N_15632,N_15647);
nor U15697 (N_15697,N_15646,N_15625);
xor U15698 (N_15698,N_15581,N_15678);
nor U15699 (N_15699,N_15672,N_15658);
and U15700 (N_15700,N_15634,N_15616);
or U15701 (N_15701,N_15531,N_15557);
xnor U15702 (N_15702,N_15530,N_15617);
and U15703 (N_15703,N_15673,N_15566);
xnor U15704 (N_15704,N_15631,N_15609);
nor U15705 (N_15705,N_15534,N_15665);
xor U15706 (N_15706,N_15611,N_15535);
and U15707 (N_15707,N_15654,N_15546);
xor U15708 (N_15708,N_15555,N_15603);
and U15709 (N_15709,N_15666,N_15662);
nor U15710 (N_15710,N_15583,N_15552);
or U15711 (N_15711,N_15594,N_15542);
xor U15712 (N_15712,N_15561,N_15602);
xor U15713 (N_15713,N_15565,N_15608);
nor U15714 (N_15714,N_15522,N_15620);
nor U15715 (N_15715,N_15560,N_15667);
and U15716 (N_15716,N_15536,N_15628);
and U15717 (N_15717,N_15520,N_15657);
and U15718 (N_15718,N_15596,N_15585);
or U15719 (N_15719,N_15579,N_15626);
and U15720 (N_15720,N_15670,N_15610);
or U15721 (N_15721,N_15533,N_15569);
or U15722 (N_15722,N_15618,N_15551);
nor U15723 (N_15723,N_15580,N_15635);
nor U15724 (N_15724,N_15643,N_15639);
or U15725 (N_15725,N_15540,N_15624);
xor U15726 (N_15726,N_15669,N_15607);
nor U15727 (N_15727,N_15528,N_15659);
and U15728 (N_15728,N_15572,N_15571);
nand U15729 (N_15729,N_15623,N_15679);
xnor U15730 (N_15730,N_15612,N_15606);
nand U15731 (N_15731,N_15676,N_15630);
nor U15732 (N_15732,N_15660,N_15577);
nand U15733 (N_15733,N_15590,N_15597);
xnor U15734 (N_15734,N_15613,N_15668);
nor U15735 (N_15735,N_15549,N_15661);
or U15736 (N_15736,N_15574,N_15582);
xnor U15737 (N_15737,N_15567,N_15656);
nor U15738 (N_15738,N_15633,N_15578);
nand U15739 (N_15739,N_15598,N_15674);
nor U15740 (N_15740,N_15593,N_15663);
nor U15741 (N_15741,N_15537,N_15651);
and U15742 (N_15742,N_15648,N_15645);
and U15743 (N_15743,N_15655,N_15573);
and U15744 (N_15744,N_15599,N_15652);
or U15745 (N_15745,N_15532,N_15589);
or U15746 (N_15746,N_15553,N_15604);
nand U15747 (N_15747,N_15621,N_15570);
nand U15748 (N_15748,N_15543,N_15622);
nand U15749 (N_15749,N_15575,N_15539);
and U15750 (N_15750,N_15576,N_15550);
and U15751 (N_15751,N_15587,N_15527);
or U15752 (N_15752,N_15545,N_15563);
nor U15753 (N_15753,N_15544,N_15644);
nand U15754 (N_15754,N_15629,N_15614);
nor U15755 (N_15755,N_15584,N_15642);
nor U15756 (N_15756,N_15524,N_15605);
and U15757 (N_15757,N_15523,N_15640);
and U15758 (N_15758,N_15588,N_15526);
xnor U15759 (N_15759,N_15619,N_15541);
nor U15760 (N_15760,N_15629,N_15571);
or U15761 (N_15761,N_15547,N_15563);
nand U15762 (N_15762,N_15636,N_15655);
nor U15763 (N_15763,N_15609,N_15544);
nor U15764 (N_15764,N_15538,N_15564);
or U15765 (N_15765,N_15633,N_15660);
and U15766 (N_15766,N_15647,N_15671);
nand U15767 (N_15767,N_15628,N_15648);
or U15768 (N_15768,N_15549,N_15538);
xnor U15769 (N_15769,N_15603,N_15620);
or U15770 (N_15770,N_15523,N_15602);
nand U15771 (N_15771,N_15570,N_15591);
nand U15772 (N_15772,N_15667,N_15678);
xnor U15773 (N_15773,N_15562,N_15640);
and U15774 (N_15774,N_15606,N_15651);
nand U15775 (N_15775,N_15572,N_15596);
or U15776 (N_15776,N_15653,N_15646);
nor U15777 (N_15777,N_15597,N_15643);
nand U15778 (N_15778,N_15620,N_15553);
nand U15779 (N_15779,N_15638,N_15544);
or U15780 (N_15780,N_15536,N_15592);
and U15781 (N_15781,N_15643,N_15650);
or U15782 (N_15782,N_15605,N_15673);
or U15783 (N_15783,N_15554,N_15625);
or U15784 (N_15784,N_15623,N_15633);
nand U15785 (N_15785,N_15542,N_15615);
nand U15786 (N_15786,N_15604,N_15600);
nand U15787 (N_15787,N_15533,N_15678);
or U15788 (N_15788,N_15540,N_15543);
and U15789 (N_15789,N_15658,N_15557);
nand U15790 (N_15790,N_15536,N_15650);
xor U15791 (N_15791,N_15536,N_15560);
xnor U15792 (N_15792,N_15599,N_15586);
or U15793 (N_15793,N_15673,N_15638);
and U15794 (N_15794,N_15578,N_15532);
and U15795 (N_15795,N_15630,N_15627);
nor U15796 (N_15796,N_15577,N_15641);
xor U15797 (N_15797,N_15541,N_15567);
nor U15798 (N_15798,N_15672,N_15650);
nor U15799 (N_15799,N_15529,N_15564);
xor U15800 (N_15800,N_15622,N_15539);
nand U15801 (N_15801,N_15626,N_15521);
nor U15802 (N_15802,N_15679,N_15529);
and U15803 (N_15803,N_15617,N_15531);
xnor U15804 (N_15804,N_15632,N_15658);
or U15805 (N_15805,N_15658,N_15588);
xor U15806 (N_15806,N_15550,N_15522);
and U15807 (N_15807,N_15661,N_15527);
and U15808 (N_15808,N_15569,N_15539);
xnor U15809 (N_15809,N_15574,N_15601);
and U15810 (N_15810,N_15528,N_15547);
and U15811 (N_15811,N_15525,N_15657);
nor U15812 (N_15812,N_15660,N_15647);
and U15813 (N_15813,N_15609,N_15632);
nand U15814 (N_15814,N_15639,N_15540);
or U15815 (N_15815,N_15538,N_15590);
nand U15816 (N_15816,N_15676,N_15679);
or U15817 (N_15817,N_15578,N_15637);
nand U15818 (N_15818,N_15664,N_15555);
and U15819 (N_15819,N_15577,N_15575);
nand U15820 (N_15820,N_15615,N_15523);
and U15821 (N_15821,N_15593,N_15666);
or U15822 (N_15822,N_15672,N_15619);
nand U15823 (N_15823,N_15649,N_15597);
and U15824 (N_15824,N_15546,N_15676);
or U15825 (N_15825,N_15624,N_15543);
nand U15826 (N_15826,N_15600,N_15635);
nand U15827 (N_15827,N_15613,N_15528);
nand U15828 (N_15828,N_15558,N_15566);
nand U15829 (N_15829,N_15522,N_15648);
or U15830 (N_15830,N_15657,N_15565);
or U15831 (N_15831,N_15610,N_15656);
nand U15832 (N_15832,N_15675,N_15649);
nor U15833 (N_15833,N_15589,N_15614);
and U15834 (N_15834,N_15625,N_15679);
or U15835 (N_15835,N_15624,N_15568);
nor U15836 (N_15836,N_15523,N_15639);
and U15837 (N_15837,N_15653,N_15634);
xor U15838 (N_15838,N_15612,N_15546);
xor U15839 (N_15839,N_15650,N_15544);
nor U15840 (N_15840,N_15814,N_15802);
and U15841 (N_15841,N_15738,N_15789);
nand U15842 (N_15842,N_15779,N_15772);
nor U15843 (N_15843,N_15766,N_15699);
or U15844 (N_15844,N_15823,N_15806);
or U15845 (N_15845,N_15793,N_15709);
and U15846 (N_15846,N_15711,N_15834);
nor U15847 (N_15847,N_15783,N_15830);
nand U15848 (N_15848,N_15797,N_15721);
xor U15849 (N_15849,N_15715,N_15786);
or U15850 (N_15850,N_15712,N_15728);
nor U15851 (N_15851,N_15730,N_15799);
nor U15852 (N_15852,N_15832,N_15700);
or U15853 (N_15853,N_15810,N_15753);
or U15854 (N_15854,N_15778,N_15803);
xnor U15855 (N_15855,N_15685,N_15795);
xnor U15856 (N_15856,N_15749,N_15773);
and U15857 (N_15857,N_15831,N_15705);
or U15858 (N_15858,N_15737,N_15724);
nand U15859 (N_15859,N_15694,N_15757);
nor U15860 (N_15860,N_15718,N_15734);
nor U15861 (N_15861,N_15782,N_15771);
or U15862 (N_15862,N_15827,N_15731);
nand U15863 (N_15863,N_15798,N_15726);
or U15864 (N_15864,N_15774,N_15760);
xnor U15865 (N_15865,N_15689,N_15791);
nor U15866 (N_15866,N_15833,N_15720);
or U15867 (N_15867,N_15743,N_15698);
xor U15868 (N_15868,N_15765,N_15707);
nor U15869 (N_15869,N_15691,N_15836);
nand U15870 (N_15870,N_15751,N_15796);
and U15871 (N_15871,N_15829,N_15756);
or U15872 (N_15872,N_15838,N_15727);
or U15873 (N_15873,N_15736,N_15742);
nand U15874 (N_15874,N_15701,N_15818);
nor U15875 (N_15875,N_15807,N_15761);
or U15876 (N_15876,N_15781,N_15811);
xor U15877 (N_15877,N_15746,N_15735);
nor U15878 (N_15878,N_15695,N_15792);
nand U15879 (N_15879,N_15682,N_15717);
xor U15880 (N_15880,N_15755,N_15828);
xor U15881 (N_15881,N_15775,N_15770);
xnor U15882 (N_15882,N_15710,N_15713);
or U15883 (N_15883,N_15748,N_15784);
xnor U15884 (N_15884,N_15835,N_15733);
nand U15885 (N_15885,N_15801,N_15839);
and U15886 (N_15886,N_15697,N_15816);
xnor U15887 (N_15887,N_15692,N_15822);
nor U15888 (N_15888,N_15714,N_15812);
or U15889 (N_15889,N_15719,N_15725);
nor U15890 (N_15890,N_15794,N_15716);
or U15891 (N_15891,N_15815,N_15729);
nor U15892 (N_15892,N_15688,N_15684);
xor U15893 (N_15893,N_15758,N_15776);
xnor U15894 (N_15894,N_15777,N_15747);
xor U15895 (N_15895,N_15706,N_15752);
or U15896 (N_15896,N_15762,N_15763);
xor U15897 (N_15897,N_15808,N_15800);
xnor U15898 (N_15898,N_15817,N_15693);
nor U15899 (N_15899,N_15681,N_15764);
xnor U15900 (N_15900,N_15740,N_15813);
nor U15901 (N_15901,N_15820,N_15739);
xor U15902 (N_15902,N_15741,N_15722);
nor U15903 (N_15903,N_15754,N_15750);
nand U15904 (N_15904,N_15826,N_15805);
nor U15905 (N_15905,N_15702,N_15690);
nand U15906 (N_15906,N_15819,N_15825);
or U15907 (N_15907,N_15686,N_15759);
xor U15908 (N_15908,N_15824,N_15821);
and U15909 (N_15909,N_15790,N_15696);
nand U15910 (N_15910,N_15780,N_15744);
nand U15911 (N_15911,N_15745,N_15723);
xnor U15912 (N_15912,N_15804,N_15703);
nor U15913 (N_15913,N_15768,N_15683);
and U15914 (N_15914,N_15809,N_15732);
nand U15915 (N_15915,N_15787,N_15680);
and U15916 (N_15916,N_15708,N_15785);
xnor U15917 (N_15917,N_15837,N_15767);
or U15918 (N_15918,N_15704,N_15687);
or U15919 (N_15919,N_15788,N_15769);
nor U15920 (N_15920,N_15725,N_15816);
nor U15921 (N_15921,N_15699,N_15771);
and U15922 (N_15922,N_15774,N_15700);
nand U15923 (N_15923,N_15775,N_15801);
xor U15924 (N_15924,N_15774,N_15703);
xnor U15925 (N_15925,N_15711,N_15719);
or U15926 (N_15926,N_15729,N_15810);
nand U15927 (N_15927,N_15756,N_15834);
nand U15928 (N_15928,N_15818,N_15697);
and U15929 (N_15929,N_15838,N_15807);
xnor U15930 (N_15930,N_15710,N_15791);
xor U15931 (N_15931,N_15835,N_15739);
or U15932 (N_15932,N_15688,N_15769);
nor U15933 (N_15933,N_15823,N_15695);
or U15934 (N_15934,N_15770,N_15802);
nor U15935 (N_15935,N_15802,N_15750);
and U15936 (N_15936,N_15708,N_15690);
nand U15937 (N_15937,N_15809,N_15688);
nand U15938 (N_15938,N_15819,N_15757);
and U15939 (N_15939,N_15790,N_15814);
nand U15940 (N_15940,N_15735,N_15774);
nor U15941 (N_15941,N_15795,N_15796);
or U15942 (N_15942,N_15823,N_15756);
xor U15943 (N_15943,N_15751,N_15710);
nand U15944 (N_15944,N_15835,N_15806);
nor U15945 (N_15945,N_15835,N_15758);
or U15946 (N_15946,N_15703,N_15705);
nand U15947 (N_15947,N_15704,N_15709);
nand U15948 (N_15948,N_15839,N_15787);
xor U15949 (N_15949,N_15725,N_15731);
xnor U15950 (N_15950,N_15766,N_15728);
or U15951 (N_15951,N_15695,N_15736);
xnor U15952 (N_15952,N_15776,N_15739);
nand U15953 (N_15953,N_15812,N_15764);
xor U15954 (N_15954,N_15837,N_15763);
xor U15955 (N_15955,N_15778,N_15787);
or U15956 (N_15956,N_15829,N_15695);
or U15957 (N_15957,N_15726,N_15835);
or U15958 (N_15958,N_15725,N_15805);
and U15959 (N_15959,N_15750,N_15726);
xnor U15960 (N_15960,N_15802,N_15731);
and U15961 (N_15961,N_15752,N_15741);
xor U15962 (N_15962,N_15776,N_15734);
nor U15963 (N_15963,N_15743,N_15702);
xor U15964 (N_15964,N_15714,N_15776);
and U15965 (N_15965,N_15796,N_15776);
or U15966 (N_15966,N_15735,N_15821);
nand U15967 (N_15967,N_15758,N_15741);
nand U15968 (N_15968,N_15823,N_15814);
and U15969 (N_15969,N_15704,N_15828);
nand U15970 (N_15970,N_15808,N_15707);
or U15971 (N_15971,N_15837,N_15717);
or U15972 (N_15972,N_15768,N_15770);
and U15973 (N_15973,N_15685,N_15725);
or U15974 (N_15974,N_15729,N_15771);
and U15975 (N_15975,N_15822,N_15740);
and U15976 (N_15976,N_15696,N_15700);
nand U15977 (N_15977,N_15824,N_15796);
and U15978 (N_15978,N_15772,N_15690);
xor U15979 (N_15979,N_15774,N_15719);
xor U15980 (N_15980,N_15744,N_15693);
nor U15981 (N_15981,N_15765,N_15809);
xor U15982 (N_15982,N_15742,N_15703);
nor U15983 (N_15983,N_15680,N_15684);
nand U15984 (N_15984,N_15799,N_15768);
nor U15985 (N_15985,N_15752,N_15759);
nand U15986 (N_15986,N_15825,N_15831);
nand U15987 (N_15987,N_15759,N_15703);
or U15988 (N_15988,N_15781,N_15805);
and U15989 (N_15989,N_15804,N_15685);
xnor U15990 (N_15990,N_15800,N_15743);
and U15991 (N_15991,N_15817,N_15722);
xnor U15992 (N_15992,N_15737,N_15772);
nor U15993 (N_15993,N_15710,N_15769);
and U15994 (N_15994,N_15699,N_15749);
xor U15995 (N_15995,N_15819,N_15740);
nand U15996 (N_15996,N_15703,N_15693);
and U15997 (N_15997,N_15727,N_15772);
or U15998 (N_15998,N_15838,N_15724);
nand U15999 (N_15999,N_15744,N_15807);
or U16000 (N_16000,N_15948,N_15886);
and U16001 (N_16001,N_15979,N_15920);
xor U16002 (N_16002,N_15849,N_15859);
nand U16003 (N_16003,N_15980,N_15997);
nand U16004 (N_16004,N_15852,N_15900);
xnor U16005 (N_16005,N_15922,N_15888);
nand U16006 (N_16006,N_15950,N_15840);
nand U16007 (N_16007,N_15915,N_15893);
nand U16008 (N_16008,N_15941,N_15882);
and U16009 (N_16009,N_15887,N_15988);
nor U16010 (N_16010,N_15848,N_15961);
nand U16011 (N_16011,N_15914,N_15912);
or U16012 (N_16012,N_15935,N_15949);
nor U16013 (N_16013,N_15927,N_15861);
or U16014 (N_16014,N_15963,N_15860);
nand U16015 (N_16015,N_15937,N_15916);
or U16016 (N_16016,N_15946,N_15999);
or U16017 (N_16017,N_15991,N_15984);
and U16018 (N_16018,N_15952,N_15890);
nand U16019 (N_16019,N_15868,N_15934);
nor U16020 (N_16020,N_15926,N_15845);
nand U16021 (N_16021,N_15958,N_15876);
or U16022 (N_16022,N_15933,N_15929);
or U16023 (N_16023,N_15925,N_15974);
nor U16024 (N_16024,N_15919,N_15936);
nor U16025 (N_16025,N_15978,N_15905);
xor U16026 (N_16026,N_15921,N_15879);
and U16027 (N_16027,N_15871,N_15875);
and U16028 (N_16028,N_15990,N_15904);
nor U16029 (N_16029,N_15866,N_15970);
nand U16030 (N_16030,N_15851,N_15960);
nand U16031 (N_16031,N_15940,N_15867);
nand U16032 (N_16032,N_15923,N_15917);
xnor U16033 (N_16033,N_15853,N_15865);
or U16034 (N_16034,N_15944,N_15982);
nor U16035 (N_16035,N_15878,N_15895);
nor U16036 (N_16036,N_15842,N_15956);
nand U16037 (N_16037,N_15966,N_15889);
or U16038 (N_16038,N_15996,N_15939);
or U16039 (N_16039,N_15942,N_15924);
xor U16040 (N_16040,N_15930,N_15907);
or U16041 (N_16041,N_15987,N_15881);
and U16042 (N_16042,N_15869,N_15953);
and U16043 (N_16043,N_15903,N_15971);
and U16044 (N_16044,N_15894,N_15901);
or U16045 (N_16045,N_15891,N_15843);
xor U16046 (N_16046,N_15918,N_15972);
or U16047 (N_16047,N_15884,N_15947);
nand U16048 (N_16048,N_15962,N_15870);
or U16049 (N_16049,N_15985,N_15994);
xor U16050 (N_16050,N_15973,N_15898);
nand U16051 (N_16051,N_15976,N_15945);
xnor U16052 (N_16052,N_15844,N_15964);
nand U16053 (N_16053,N_15969,N_15856);
or U16054 (N_16054,N_15847,N_15897);
xnor U16055 (N_16055,N_15986,N_15855);
nand U16056 (N_16056,N_15880,N_15975);
nand U16057 (N_16057,N_15858,N_15885);
and U16058 (N_16058,N_15932,N_15899);
nor U16059 (N_16059,N_15998,N_15931);
nor U16060 (N_16060,N_15872,N_15951);
xor U16061 (N_16061,N_15902,N_15977);
nor U16062 (N_16062,N_15995,N_15943);
nor U16063 (N_16063,N_15989,N_15873);
nand U16064 (N_16064,N_15911,N_15959);
xnor U16065 (N_16065,N_15908,N_15909);
nand U16066 (N_16066,N_15864,N_15993);
xor U16067 (N_16067,N_15910,N_15846);
nor U16068 (N_16068,N_15906,N_15874);
nor U16069 (N_16069,N_15954,N_15892);
nand U16070 (N_16070,N_15841,N_15862);
nand U16071 (N_16071,N_15863,N_15968);
nand U16072 (N_16072,N_15965,N_15857);
and U16073 (N_16073,N_15850,N_15938);
or U16074 (N_16074,N_15877,N_15928);
xor U16075 (N_16075,N_15992,N_15983);
nand U16076 (N_16076,N_15883,N_15913);
or U16077 (N_16077,N_15955,N_15957);
nor U16078 (N_16078,N_15896,N_15967);
or U16079 (N_16079,N_15854,N_15981);
or U16080 (N_16080,N_15999,N_15957);
or U16081 (N_16081,N_15851,N_15933);
and U16082 (N_16082,N_15942,N_15990);
or U16083 (N_16083,N_15850,N_15981);
nor U16084 (N_16084,N_15905,N_15880);
and U16085 (N_16085,N_15847,N_15872);
nor U16086 (N_16086,N_15987,N_15902);
and U16087 (N_16087,N_15868,N_15972);
xnor U16088 (N_16088,N_15989,N_15866);
nand U16089 (N_16089,N_15974,N_15845);
nor U16090 (N_16090,N_15873,N_15892);
or U16091 (N_16091,N_15863,N_15937);
nand U16092 (N_16092,N_15960,N_15958);
or U16093 (N_16093,N_15958,N_15920);
or U16094 (N_16094,N_15858,N_15915);
and U16095 (N_16095,N_15934,N_15987);
and U16096 (N_16096,N_15904,N_15968);
nor U16097 (N_16097,N_15975,N_15970);
xor U16098 (N_16098,N_15994,N_15940);
and U16099 (N_16099,N_15994,N_15878);
and U16100 (N_16100,N_15971,N_15927);
nor U16101 (N_16101,N_15887,N_15871);
or U16102 (N_16102,N_15909,N_15943);
xnor U16103 (N_16103,N_15989,N_15980);
nor U16104 (N_16104,N_15958,N_15903);
nor U16105 (N_16105,N_15986,N_15900);
nand U16106 (N_16106,N_15976,N_15845);
xnor U16107 (N_16107,N_15895,N_15997);
xor U16108 (N_16108,N_15934,N_15899);
or U16109 (N_16109,N_15899,N_15952);
xor U16110 (N_16110,N_15849,N_15880);
or U16111 (N_16111,N_15991,N_15845);
nand U16112 (N_16112,N_15981,N_15911);
nand U16113 (N_16113,N_15959,N_15972);
xnor U16114 (N_16114,N_15881,N_15947);
nand U16115 (N_16115,N_15859,N_15860);
or U16116 (N_16116,N_15988,N_15900);
or U16117 (N_16117,N_15942,N_15861);
xnor U16118 (N_16118,N_15879,N_15967);
nand U16119 (N_16119,N_15938,N_15870);
or U16120 (N_16120,N_15958,N_15934);
xor U16121 (N_16121,N_15906,N_15963);
and U16122 (N_16122,N_15934,N_15882);
nand U16123 (N_16123,N_15845,N_15932);
nand U16124 (N_16124,N_15877,N_15853);
xor U16125 (N_16125,N_15899,N_15931);
nor U16126 (N_16126,N_15848,N_15940);
or U16127 (N_16127,N_15887,N_15851);
xor U16128 (N_16128,N_15928,N_15958);
xnor U16129 (N_16129,N_15929,N_15891);
and U16130 (N_16130,N_15958,N_15862);
xor U16131 (N_16131,N_15913,N_15870);
nor U16132 (N_16132,N_15963,N_15883);
nor U16133 (N_16133,N_15906,N_15960);
or U16134 (N_16134,N_15965,N_15874);
nand U16135 (N_16135,N_15909,N_15885);
or U16136 (N_16136,N_15861,N_15900);
and U16137 (N_16137,N_15967,N_15981);
or U16138 (N_16138,N_15860,N_15875);
xnor U16139 (N_16139,N_15987,N_15959);
and U16140 (N_16140,N_15849,N_15932);
and U16141 (N_16141,N_15975,N_15867);
nand U16142 (N_16142,N_15841,N_15992);
or U16143 (N_16143,N_15945,N_15885);
xor U16144 (N_16144,N_15870,N_15950);
xnor U16145 (N_16145,N_15860,N_15858);
xnor U16146 (N_16146,N_15898,N_15995);
or U16147 (N_16147,N_15960,N_15971);
xor U16148 (N_16148,N_15847,N_15876);
xor U16149 (N_16149,N_15981,N_15977);
or U16150 (N_16150,N_15985,N_15995);
nor U16151 (N_16151,N_15887,N_15890);
xnor U16152 (N_16152,N_15933,N_15924);
nor U16153 (N_16153,N_15931,N_15921);
nand U16154 (N_16154,N_15852,N_15948);
or U16155 (N_16155,N_15907,N_15846);
nor U16156 (N_16156,N_15972,N_15883);
or U16157 (N_16157,N_15969,N_15865);
nor U16158 (N_16158,N_15853,N_15850);
nand U16159 (N_16159,N_15866,N_15896);
or U16160 (N_16160,N_16008,N_16030);
nor U16161 (N_16161,N_16119,N_16031);
nor U16162 (N_16162,N_16064,N_16141);
nor U16163 (N_16163,N_16101,N_16013);
and U16164 (N_16164,N_16085,N_16086);
or U16165 (N_16165,N_16061,N_16106);
xor U16166 (N_16166,N_16103,N_16107);
nand U16167 (N_16167,N_16140,N_16063);
and U16168 (N_16168,N_16018,N_16081);
nand U16169 (N_16169,N_16058,N_16075);
nor U16170 (N_16170,N_16056,N_16045);
and U16171 (N_16171,N_16098,N_16012);
xnor U16172 (N_16172,N_16040,N_16122);
or U16173 (N_16173,N_16132,N_16087);
nor U16174 (N_16174,N_16108,N_16145);
xnor U16175 (N_16175,N_16026,N_16003);
nand U16176 (N_16176,N_16129,N_16046);
nor U16177 (N_16177,N_16148,N_16102);
or U16178 (N_16178,N_16002,N_16143);
or U16179 (N_16179,N_16051,N_16017);
nand U16180 (N_16180,N_16094,N_16009);
and U16181 (N_16181,N_16109,N_16110);
xor U16182 (N_16182,N_16076,N_16077);
nand U16183 (N_16183,N_16149,N_16156);
or U16184 (N_16184,N_16000,N_16069);
or U16185 (N_16185,N_16136,N_16139);
nand U16186 (N_16186,N_16055,N_16020);
nand U16187 (N_16187,N_16037,N_16135);
and U16188 (N_16188,N_16151,N_16089);
nand U16189 (N_16189,N_16041,N_16070);
xnor U16190 (N_16190,N_16091,N_16146);
nand U16191 (N_16191,N_16095,N_16042);
or U16192 (N_16192,N_16019,N_16127);
and U16193 (N_16193,N_16130,N_16027);
xnor U16194 (N_16194,N_16074,N_16072);
and U16195 (N_16195,N_16142,N_16112);
nor U16196 (N_16196,N_16053,N_16153);
nor U16197 (N_16197,N_16100,N_16134);
xnor U16198 (N_16198,N_16044,N_16120);
nor U16199 (N_16199,N_16138,N_16029);
and U16200 (N_16200,N_16039,N_16060);
xor U16201 (N_16201,N_16016,N_16154);
nor U16202 (N_16202,N_16006,N_16096);
xor U16203 (N_16203,N_16005,N_16057);
xnor U16204 (N_16204,N_16117,N_16032);
xnor U16205 (N_16205,N_16073,N_16092);
xnor U16206 (N_16206,N_16021,N_16099);
xor U16207 (N_16207,N_16155,N_16048);
nor U16208 (N_16208,N_16043,N_16025);
xor U16209 (N_16209,N_16083,N_16080);
or U16210 (N_16210,N_16001,N_16144);
xor U16211 (N_16211,N_16050,N_16115);
xnor U16212 (N_16212,N_16126,N_16078);
and U16213 (N_16213,N_16066,N_16022);
nor U16214 (N_16214,N_16097,N_16125);
and U16215 (N_16215,N_16123,N_16024);
xnor U16216 (N_16216,N_16111,N_16152);
xnor U16217 (N_16217,N_16038,N_16105);
and U16218 (N_16218,N_16068,N_16010);
and U16219 (N_16219,N_16067,N_16007);
and U16220 (N_16220,N_16015,N_16071);
nor U16221 (N_16221,N_16150,N_16082);
nand U16222 (N_16222,N_16054,N_16034);
nor U16223 (N_16223,N_16124,N_16118);
nand U16224 (N_16224,N_16157,N_16079);
nand U16225 (N_16225,N_16158,N_16052);
nand U16226 (N_16226,N_16033,N_16088);
xor U16227 (N_16227,N_16059,N_16113);
nand U16228 (N_16228,N_16131,N_16159);
and U16229 (N_16229,N_16028,N_16147);
and U16230 (N_16230,N_16011,N_16023);
nor U16231 (N_16231,N_16014,N_16114);
xnor U16232 (N_16232,N_16116,N_16084);
nand U16233 (N_16233,N_16049,N_16121);
nor U16234 (N_16234,N_16104,N_16047);
xnor U16235 (N_16235,N_16065,N_16137);
nand U16236 (N_16236,N_16093,N_16062);
nor U16237 (N_16237,N_16004,N_16036);
and U16238 (N_16238,N_16090,N_16035);
nor U16239 (N_16239,N_16133,N_16128);
nand U16240 (N_16240,N_16101,N_16131);
nor U16241 (N_16241,N_16148,N_16018);
or U16242 (N_16242,N_16130,N_16137);
xnor U16243 (N_16243,N_16156,N_16039);
nand U16244 (N_16244,N_16152,N_16090);
or U16245 (N_16245,N_16128,N_16054);
nand U16246 (N_16246,N_16156,N_16074);
nor U16247 (N_16247,N_16071,N_16126);
nand U16248 (N_16248,N_16054,N_16139);
xnor U16249 (N_16249,N_16146,N_16157);
or U16250 (N_16250,N_16107,N_16017);
nor U16251 (N_16251,N_16154,N_16030);
and U16252 (N_16252,N_16121,N_16019);
nand U16253 (N_16253,N_16078,N_16132);
xor U16254 (N_16254,N_16056,N_16098);
or U16255 (N_16255,N_16025,N_16054);
nor U16256 (N_16256,N_16007,N_16147);
or U16257 (N_16257,N_16124,N_16094);
nand U16258 (N_16258,N_16043,N_16124);
and U16259 (N_16259,N_16026,N_16053);
nor U16260 (N_16260,N_16065,N_16000);
or U16261 (N_16261,N_16020,N_16070);
nand U16262 (N_16262,N_16032,N_16111);
nor U16263 (N_16263,N_16028,N_16145);
nand U16264 (N_16264,N_16054,N_16001);
xor U16265 (N_16265,N_16006,N_16043);
and U16266 (N_16266,N_16138,N_16068);
or U16267 (N_16267,N_16156,N_16000);
nand U16268 (N_16268,N_16147,N_16015);
xor U16269 (N_16269,N_16119,N_16049);
and U16270 (N_16270,N_16070,N_16076);
xnor U16271 (N_16271,N_16050,N_16141);
nand U16272 (N_16272,N_16125,N_16098);
nand U16273 (N_16273,N_16010,N_16136);
and U16274 (N_16274,N_16012,N_16006);
xor U16275 (N_16275,N_16070,N_16134);
and U16276 (N_16276,N_16049,N_16036);
and U16277 (N_16277,N_16090,N_16080);
and U16278 (N_16278,N_16056,N_16127);
nor U16279 (N_16279,N_16010,N_16073);
nor U16280 (N_16280,N_16048,N_16036);
xor U16281 (N_16281,N_16012,N_16099);
or U16282 (N_16282,N_16139,N_16057);
or U16283 (N_16283,N_16027,N_16017);
nand U16284 (N_16284,N_16076,N_16008);
and U16285 (N_16285,N_16128,N_16138);
nand U16286 (N_16286,N_16021,N_16015);
and U16287 (N_16287,N_16049,N_16108);
nor U16288 (N_16288,N_16003,N_16130);
xor U16289 (N_16289,N_16005,N_16043);
or U16290 (N_16290,N_16156,N_16092);
nor U16291 (N_16291,N_16133,N_16009);
nor U16292 (N_16292,N_16137,N_16091);
and U16293 (N_16293,N_16154,N_16117);
nor U16294 (N_16294,N_16145,N_16102);
and U16295 (N_16295,N_16094,N_16119);
xnor U16296 (N_16296,N_16054,N_16121);
and U16297 (N_16297,N_16066,N_16159);
nor U16298 (N_16298,N_16144,N_16029);
nor U16299 (N_16299,N_16060,N_16077);
and U16300 (N_16300,N_16057,N_16025);
or U16301 (N_16301,N_16047,N_16068);
xor U16302 (N_16302,N_16034,N_16039);
nor U16303 (N_16303,N_16104,N_16134);
or U16304 (N_16304,N_16159,N_16040);
nor U16305 (N_16305,N_16032,N_16067);
and U16306 (N_16306,N_16115,N_16134);
nand U16307 (N_16307,N_16002,N_16144);
and U16308 (N_16308,N_16049,N_16078);
nand U16309 (N_16309,N_16155,N_16062);
nand U16310 (N_16310,N_16095,N_16103);
or U16311 (N_16311,N_16023,N_16126);
xor U16312 (N_16312,N_16041,N_16035);
nor U16313 (N_16313,N_16072,N_16158);
and U16314 (N_16314,N_16020,N_16009);
nand U16315 (N_16315,N_16129,N_16103);
xnor U16316 (N_16316,N_16104,N_16039);
xnor U16317 (N_16317,N_16076,N_16066);
and U16318 (N_16318,N_16136,N_16014);
xor U16319 (N_16319,N_16130,N_16121);
xor U16320 (N_16320,N_16161,N_16209);
xnor U16321 (N_16321,N_16234,N_16302);
xor U16322 (N_16322,N_16300,N_16168);
nand U16323 (N_16323,N_16272,N_16292);
xnor U16324 (N_16324,N_16180,N_16265);
nand U16325 (N_16325,N_16258,N_16224);
or U16326 (N_16326,N_16236,N_16166);
xnor U16327 (N_16327,N_16241,N_16288);
or U16328 (N_16328,N_16313,N_16193);
nand U16329 (N_16329,N_16256,N_16197);
or U16330 (N_16330,N_16246,N_16240);
and U16331 (N_16331,N_16231,N_16282);
xor U16332 (N_16332,N_16305,N_16195);
and U16333 (N_16333,N_16179,N_16283);
xnor U16334 (N_16334,N_16277,N_16307);
nand U16335 (N_16335,N_16296,N_16188);
or U16336 (N_16336,N_16306,N_16171);
and U16337 (N_16337,N_16235,N_16250);
and U16338 (N_16338,N_16278,N_16269);
nor U16339 (N_16339,N_16294,N_16257);
or U16340 (N_16340,N_16217,N_16252);
or U16341 (N_16341,N_16316,N_16230);
or U16342 (N_16342,N_16259,N_16215);
and U16343 (N_16343,N_16206,N_16167);
or U16344 (N_16344,N_16199,N_16196);
nand U16345 (N_16345,N_16309,N_16220);
nor U16346 (N_16346,N_16244,N_16263);
and U16347 (N_16347,N_16295,N_16284);
nor U16348 (N_16348,N_16249,N_16315);
xor U16349 (N_16349,N_16183,N_16191);
xor U16350 (N_16350,N_16226,N_16271);
and U16351 (N_16351,N_16312,N_16243);
or U16352 (N_16352,N_16237,N_16178);
and U16353 (N_16353,N_16318,N_16186);
and U16354 (N_16354,N_16164,N_16262);
xor U16355 (N_16355,N_16213,N_16205);
and U16356 (N_16356,N_16253,N_16297);
nor U16357 (N_16357,N_16293,N_16202);
xor U16358 (N_16358,N_16308,N_16163);
xnor U16359 (N_16359,N_16255,N_16317);
xnor U16360 (N_16360,N_16203,N_16176);
nand U16361 (N_16361,N_16212,N_16304);
nand U16362 (N_16362,N_16264,N_16273);
and U16363 (N_16363,N_16242,N_16267);
nand U16364 (N_16364,N_16221,N_16286);
nor U16365 (N_16365,N_16266,N_16268);
and U16366 (N_16366,N_16211,N_16208);
or U16367 (N_16367,N_16169,N_16239);
nand U16368 (N_16368,N_16160,N_16314);
or U16369 (N_16369,N_16172,N_16290);
nor U16370 (N_16370,N_16174,N_16173);
nor U16371 (N_16371,N_16192,N_16228);
xnor U16372 (N_16372,N_16216,N_16185);
or U16373 (N_16373,N_16170,N_16165);
or U16374 (N_16374,N_16210,N_16311);
nand U16375 (N_16375,N_16214,N_16184);
and U16376 (N_16376,N_16181,N_16245);
nor U16377 (N_16377,N_16177,N_16204);
or U16378 (N_16378,N_16247,N_16260);
xnor U16379 (N_16379,N_16248,N_16162);
nor U16380 (N_16380,N_16182,N_16189);
xor U16381 (N_16381,N_16198,N_16222);
xor U16382 (N_16382,N_16319,N_16251);
or U16383 (N_16383,N_16310,N_16285);
nor U16384 (N_16384,N_16287,N_16219);
or U16385 (N_16385,N_16232,N_16233);
nand U16386 (N_16386,N_16275,N_16223);
xor U16387 (N_16387,N_16207,N_16301);
or U16388 (N_16388,N_16194,N_16281);
nand U16389 (N_16389,N_16175,N_16190);
xor U16390 (N_16390,N_16225,N_16218);
and U16391 (N_16391,N_16229,N_16261);
and U16392 (N_16392,N_16299,N_16303);
and U16393 (N_16393,N_16289,N_16279);
xnor U16394 (N_16394,N_16238,N_16298);
and U16395 (N_16395,N_16270,N_16227);
or U16396 (N_16396,N_16201,N_16280);
nor U16397 (N_16397,N_16276,N_16200);
or U16398 (N_16398,N_16254,N_16274);
or U16399 (N_16399,N_16291,N_16187);
or U16400 (N_16400,N_16306,N_16293);
nor U16401 (N_16401,N_16213,N_16177);
xnor U16402 (N_16402,N_16166,N_16292);
or U16403 (N_16403,N_16215,N_16273);
xnor U16404 (N_16404,N_16300,N_16273);
xnor U16405 (N_16405,N_16306,N_16226);
nor U16406 (N_16406,N_16296,N_16281);
nor U16407 (N_16407,N_16317,N_16243);
xnor U16408 (N_16408,N_16183,N_16178);
xor U16409 (N_16409,N_16279,N_16187);
nand U16410 (N_16410,N_16208,N_16205);
xnor U16411 (N_16411,N_16185,N_16222);
nor U16412 (N_16412,N_16303,N_16317);
nand U16413 (N_16413,N_16188,N_16228);
nand U16414 (N_16414,N_16240,N_16203);
nand U16415 (N_16415,N_16295,N_16307);
nor U16416 (N_16416,N_16246,N_16269);
nor U16417 (N_16417,N_16281,N_16220);
or U16418 (N_16418,N_16221,N_16294);
and U16419 (N_16419,N_16209,N_16204);
nand U16420 (N_16420,N_16199,N_16250);
xnor U16421 (N_16421,N_16319,N_16318);
and U16422 (N_16422,N_16256,N_16245);
xnor U16423 (N_16423,N_16225,N_16273);
nand U16424 (N_16424,N_16214,N_16292);
xnor U16425 (N_16425,N_16258,N_16270);
nand U16426 (N_16426,N_16274,N_16186);
or U16427 (N_16427,N_16180,N_16189);
and U16428 (N_16428,N_16224,N_16196);
or U16429 (N_16429,N_16236,N_16297);
and U16430 (N_16430,N_16274,N_16227);
and U16431 (N_16431,N_16192,N_16161);
nor U16432 (N_16432,N_16163,N_16294);
xor U16433 (N_16433,N_16242,N_16295);
nor U16434 (N_16434,N_16274,N_16184);
or U16435 (N_16435,N_16294,N_16315);
nor U16436 (N_16436,N_16264,N_16202);
and U16437 (N_16437,N_16288,N_16231);
and U16438 (N_16438,N_16255,N_16183);
nor U16439 (N_16439,N_16183,N_16300);
nand U16440 (N_16440,N_16263,N_16297);
xor U16441 (N_16441,N_16287,N_16210);
and U16442 (N_16442,N_16204,N_16168);
xnor U16443 (N_16443,N_16244,N_16221);
and U16444 (N_16444,N_16277,N_16265);
or U16445 (N_16445,N_16168,N_16195);
xnor U16446 (N_16446,N_16260,N_16265);
xor U16447 (N_16447,N_16211,N_16195);
nand U16448 (N_16448,N_16235,N_16207);
nand U16449 (N_16449,N_16168,N_16221);
nand U16450 (N_16450,N_16194,N_16179);
and U16451 (N_16451,N_16170,N_16168);
nand U16452 (N_16452,N_16221,N_16305);
nor U16453 (N_16453,N_16319,N_16269);
or U16454 (N_16454,N_16191,N_16293);
and U16455 (N_16455,N_16315,N_16299);
and U16456 (N_16456,N_16291,N_16284);
or U16457 (N_16457,N_16208,N_16227);
and U16458 (N_16458,N_16249,N_16169);
or U16459 (N_16459,N_16167,N_16190);
and U16460 (N_16460,N_16187,N_16313);
and U16461 (N_16461,N_16214,N_16262);
and U16462 (N_16462,N_16268,N_16162);
or U16463 (N_16463,N_16279,N_16236);
and U16464 (N_16464,N_16251,N_16272);
and U16465 (N_16465,N_16230,N_16241);
and U16466 (N_16466,N_16221,N_16252);
nand U16467 (N_16467,N_16211,N_16237);
nor U16468 (N_16468,N_16313,N_16317);
and U16469 (N_16469,N_16194,N_16299);
nand U16470 (N_16470,N_16203,N_16227);
nor U16471 (N_16471,N_16280,N_16172);
nor U16472 (N_16472,N_16173,N_16292);
nand U16473 (N_16473,N_16298,N_16180);
or U16474 (N_16474,N_16260,N_16311);
or U16475 (N_16475,N_16270,N_16182);
nand U16476 (N_16476,N_16289,N_16266);
nor U16477 (N_16477,N_16292,N_16168);
nand U16478 (N_16478,N_16278,N_16319);
or U16479 (N_16479,N_16231,N_16280);
nand U16480 (N_16480,N_16439,N_16473);
xor U16481 (N_16481,N_16396,N_16364);
and U16482 (N_16482,N_16468,N_16463);
nand U16483 (N_16483,N_16345,N_16399);
nor U16484 (N_16484,N_16400,N_16437);
nand U16485 (N_16485,N_16394,N_16323);
or U16486 (N_16486,N_16344,N_16356);
nor U16487 (N_16487,N_16320,N_16431);
nand U16488 (N_16488,N_16448,N_16395);
or U16489 (N_16489,N_16409,N_16331);
xor U16490 (N_16490,N_16398,N_16350);
nor U16491 (N_16491,N_16430,N_16391);
and U16492 (N_16492,N_16421,N_16382);
nor U16493 (N_16493,N_16359,N_16434);
nor U16494 (N_16494,N_16371,N_16337);
and U16495 (N_16495,N_16466,N_16342);
and U16496 (N_16496,N_16328,N_16428);
nand U16497 (N_16497,N_16405,N_16377);
nor U16498 (N_16498,N_16464,N_16361);
and U16499 (N_16499,N_16392,N_16412);
and U16500 (N_16500,N_16449,N_16478);
nand U16501 (N_16501,N_16470,N_16322);
nor U16502 (N_16502,N_16378,N_16458);
nand U16503 (N_16503,N_16461,N_16414);
and U16504 (N_16504,N_16389,N_16455);
and U16505 (N_16505,N_16476,N_16452);
or U16506 (N_16506,N_16438,N_16333);
nand U16507 (N_16507,N_16354,N_16401);
and U16508 (N_16508,N_16404,N_16429);
or U16509 (N_16509,N_16424,N_16365);
nand U16510 (N_16510,N_16454,N_16366);
nand U16511 (N_16511,N_16479,N_16441);
xor U16512 (N_16512,N_16446,N_16471);
and U16513 (N_16513,N_16330,N_16386);
and U16514 (N_16514,N_16426,N_16335);
nor U16515 (N_16515,N_16406,N_16403);
xor U16516 (N_16516,N_16411,N_16450);
nand U16517 (N_16517,N_16447,N_16408);
nor U16518 (N_16518,N_16419,N_16423);
nand U16519 (N_16519,N_16397,N_16457);
or U16520 (N_16520,N_16334,N_16456);
nor U16521 (N_16521,N_16325,N_16376);
nor U16522 (N_16522,N_16341,N_16451);
nand U16523 (N_16523,N_16475,N_16368);
nor U16524 (N_16524,N_16353,N_16444);
nor U16525 (N_16525,N_16460,N_16418);
or U16526 (N_16526,N_16385,N_16357);
or U16527 (N_16527,N_16433,N_16349);
or U16528 (N_16528,N_16442,N_16375);
xor U16529 (N_16529,N_16329,N_16346);
and U16530 (N_16530,N_16427,N_16465);
nand U16531 (N_16531,N_16321,N_16372);
nand U16532 (N_16532,N_16435,N_16348);
nand U16533 (N_16533,N_16436,N_16415);
or U16534 (N_16534,N_16422,N_16467);
and U16535 (N_16535,N_16474,N_16445);
or U16536 (N_16536,N_16477,N_16388);
and U16537 (N_16537,N_16352,N_16360);
nand U16538 (N_16538,N_16432,N_16374);
and U16539 (N_16539,N_16355,N_16380);
or U16540 (N_16540,N_16407,N_16443);
nand U16541 (N_16541,N_16373,N_16416);
or U16542 (N_16542,N_16343,N_16340);
nand U16543 (N_16543,N_16338,N_16440);
nand U16544 (N_16544,N_16402,N_16383);
nor U16545 (N_16545,N_16351,N_16358);
nor U16546 (N_16546,N_16410,N_16425);
nand U16547 (N_16547,N_16379,N_16417);
and U16548 (N_16548,N_16420,N_16390);
or U16549 (N_16549,N_16362,N_16472);
and U16550 (N_16550,N_16363,N_16367);
and U16551 (N_16551,N_16381,N_16459);
or U16552 (N_16552,N_16469,N_16327);
and U16553 (N_16553,N_16332,N_16339);
xnor U16554 (N_16554,N_16347,N_16326);
or U16555 (N_16555,N_16393,N_16336);
nand U16556 (N_16556,N_16462,N_16453);
and U16557 (N_16557,N_16369,N_16324);
nand U16558 (N_16558,N_16384,N_16413);
and U16559 (N_16559,N_16370,N_16387);
xor U16560 (N_16560,N_16417,N_16430);
and U16561 (N_16561,N_16411,N_16439);
nand U16562 (N_16562,N_16463,N_16454);
xor U16563 (N_16563,N_16397,N_16434);
and U16564 (N_16564,N_16361,N_16410);
nand U16565 (N_16565,N_16372,N_16361);
nand U16566 (N_16566,N_16352,N_16415);
or U16567 (N_16567,N_16390,N_16476);
xor U16568 (N_16568,N_16442,N_16457);
or U16569 (N_16569,N_16392,N_16437);
or U16570 (N_16570,N_16343,N_16355);
xor U16571 (N_16571,N_16423,N_16449);
or U16572 (N_16572,N_16342,N_16363);
nand U16573 (N_16573,N_16428,N_16348);
or U16574 (N_16574,N_16387,N_16339);
nor U16575 (N_16575,N_16436,N_16402);
nand U16576 (N_16576,N_16463,N_16358);
xnor U16577 (N_16577,N_16460,N_16320);
nor U16578 (N_16578,N_16330,N_16378);
and U16579 (N_16579,N_16376,N_16437);
xnor U16580 (N_16580,N_16472,N_16457);
nor U16581 (N_16581,N_16422,N_16333);
and U16582 (N_16582,N_16468,N_16381);
xnor U16583 (N_16583,N_16354,N_16466);
nor U16584 (N_16584,N_16363,N_16446);
nor U16585 (N_16585,N_16479,N_16469);
and U16586 (N_16586,N_16421,N_16466);
nand U16587 (N_16587,N_16455,N_16422);
nor U16588 (N_16588,N_16440,N_16401);
nor U16589 (N_16589,N_16376,N_16351);
xor U16590 (N_16590,N_16454,N_16420);
nor U16591 (N_16591,N_16398,N_16447);
xnor U16592 (N_16592,N_16402,N_16422);
and U16593 (N_16593,N_16325,N_16442);
and U16594 (N_16594,N_16372,N_16427);
xor U16595 (N_16595,N_16394,N_16460);
nand U16596 (N_16596,N_16368,N_16382);
nor U16597 (N_16597,N_16335,N_16446);
and U16598 (N_16598,N_16406,N_16402);
nor U16599 (N_16599,N_16447,N_16361);
or U16600 (N_16600,N_16427,N_16453);
nor U16601 (N_16601,N_16450,N_16334);
nor U16602 (N_16602,N_16358,N_16433);
nor U16603 (N_16603,N_16401,N_16399);
or U16604 (N_16604,N_16375,N_16351);
or U16605 (N_16605,N_16345,N_16443);
xnor U16606 (N_16606,N_16330,N_16422);
or U16607 (N_16607,N_16470,N_16351);
xor U16608 (N_16608,N_16384,N_16456);
nand U16609 (N_16609,N_16339,N_16431);
nand U16610 (N_16610,N_16462,N_16327);
and U16611 (N_16611,N_16454,N_16361);
nor U16612 (N_16612,N_16335,N_16331);
and U16613 (N_16613,N_16330,N_16406);
or U16614 (N_16614,N_16470,N_16469);
nand U16615 (N_16615,N_16452,N_16341);
nor U16616 (N_16616,N_16405,N_16464);
or U16617 (N_16617,N_16343,N_16394);
nand U16618 (N_16618,N_16356,N_16465);
or U16619 (N_16619,N_16346,N_16401);
nand U16620 (N_16620,N_16466,N_16418);
xnor U16621 (N_16621,N_16384,N_16435);
nand U16622 (N_16622,N_16380,N_16411);
or U16623 (N_16623,N_16387,N_16455);
xnor U16624 (N_16624,N_16358,N_16321);
nor U16625 (N_16625,N_16413,N_16325);
nor U16626 (N_16626,N_16324,N_16342);
xnor U16627 (N_16627,N_16428,N_16457);
or U16628 (N_16628,N_16322,N_16423);
and U16629 (N_16629,N_16325,N_16336);
or U16630 (N_16630,N_16335,N_16431);
xnor U16631 (N_16631,N_16454,N_16358);
nand U16632 (N_16632,N_16441,N_16459);
xor U16633 (N_16633,N_16331,N_16353);
xor U16634 (N_16634,N_16392,N_16455);
nand U16635 (N_16635,N_16412,N_16469);
nand U16636 (N_16636,N_16460,N_16438);
and U16637 (N_16637,N_16442,N_16397);
xnor U16638 (N_16638,N_16384,N_16443);
nor U16639 (N_16639,N_16393,N_16425);
nand U16640 (N_16640,N_16555,N_16590);
or U16641 (N_16641,N_16603,N_16570);
xor U16642 (N_16642,N_16601,N_16502);
xnor U16643 (N_16643,N_16492,N_16559);
or U16644 (N_16644,N_16531,N_16523);
and U16645 (N_16645,N_16610,N_16627);
or U16646 (N_16646,N_16535,N_16625);
xnor U16647 (N_16647,N_16602,N_16534);
or U16648 (N_16648,N_16484,N_16600);
and U16649 (N_16649,N_16519,N_16529);
and U16650 (N_16650,N_16493,N_16591);
and U16651 (N_16651,N_16503,N_16631);
nor U16652 (N_16652,N_16541,N_16537);
nor U16653 (N_16653,N_16533,N_16510);
and U16654 (N_16654,N_16571,N_16540);
nand U16655 (N_16655,N_16482,N_16568);
nand U16656 (N_16656,N_16576,N_16536);
xnor U16657 (N_16657,N_16552,N_16528);
or U16658 (N_16658,N_16556,N_16544);
xnor U16659 (N_16659,N_16511,N_16551);
or U16660 (N_16660,N_16575,N_16614);
nor U16661 (N_16661,N_16562,N_16542);
or U16662 (N_16662,N_16596,N_16527);
or U16663 (N_16663,N_16525,N_16549);
nand U16664 (N_16664,N_16588,N_16632);
or U16665 (N_16665,N_16538,N_16530);
or U16666 (N_16666,N_16573,N_16558);
and U16667 (N_16667,N_16504,N_16619);
or U16668 (N_16668,N_16580,N_16597);
nand U16669 (N_16669,N_16506,N_16608);
nand U16670 (N_16670,N_16572,N_16498);
and U16671 (N_16671,N_16512,N_16637);
nand U16672 (N_16672,N_16481,N_16550);
xnor U16673 (N_16673,N_16574,N_16607);
nand U16674 (N_16674,N_16480,N_16606);
or U16675 (N_16675,N_16496,N_16638);
or U16676 (N_16676,N_16616,N_16626);
or U16677 (N_16677,N_16564,N_16622);
and U16678 (N_16678,N_16561,N_16560);
and U16679 (N_16679,N_16615,N_16505);
nand U16680 (N_16680,N_16557,N_16630);
and U16681 (N_16681,N_16524,N_16501);
or U16682 (N_16682,N_16584,N_16494);
and U16683 (N_16683,N_16599,N_16500);
nand U16684 (N_16684,N_16499,N_16515);
nor U16685 (N_16685,N_16553,N_16612);
nand U16686 (N_16686,N_16581,N_16563);
nor U16687 (N_16687,N_16629,N_16491);
xor U16688 (N_16688,N_16520,N_16633);
or U16689 (N_16689,N_16569,N_16583);
and U16690 (N_16690,N_16522,N_16617);
xor U16691 (N_16691,N_16628,N_16486);
nand U16692 (N_16692,N_16634,N_16636);
nand U16693 (N_16693,N_16490,N_16516);
and U16694 (N_16694,N_16548,N_16488);
and U16695 (N_16695,N_16620,N_16613);
or U16696 (N_16696,N_16497,N_16621);
nor U16697 (N_16697,N_16489,N_16566);
nand U16698 (N_16698,N_16539,N_16554);
and U16699 (N_16699,N_16485,N_16483);
nand U16700 (N_16700,N_16487,N_16495);
xnor U16701 (N_16701,N_16585,N_16577);
xor U16702 (N_16702,N_16639,N_16514);
or U16703 (N_16703,N_16578,N_16513);
nor U16704 (N_16704,N_16526,N_16509);
nand U16705 (N_16705,N_16507,N_16624);
nand U16706 (N_16706,N_16587,N_16592);
or U16707 (N_16707,N_16618,N_16579);
and U16708 (N_16708,N_16635,N_16586);
and U16709 (N_16709,N_16521,N_16593);
xnor U16710 (N_16710,N_16582,N_16595);
nor U16711 (N_16711,N_16589,N_16517);
nand U16712 (N_16712,N_16543,N_16598);
xor U16713 (N_16713,N_16532,N_16547);
nor U16714 (N_16714,N_16545,N_16611);
and U16715 (N_16715,N_16604,N_16623);
nor U16716 (N_16716,N_16565,N_16605);
nand U16717 (N_16717,N_16546,N_16594);
xor U16718 (N_16718,N_16609,N_16508);
xor U16719 (N_16719,N_16567,N_16518);
xnor U16720 (N_16720,N_16557,N_16529);
nor U16721 (N_16721,N_16631,N_16531);
and U16722 (N_16722,N_16578,N_16482);
and U16723 (N_16723,N_16567,N_16636);
nor U16724 (N_16724,N_16627,N_16505);
xnor U16725 (N_16725,N_16539,N_16521);
or U16726 (N_16726,N_16609,N_16512);
xnor U16727 (N_16727,N_16504,N_16595);
nor U16728 (N_16728,N_16580,N_16538);
nand U16729 (N_16729,N_16574,N_16617);
nor U16730 (N_16730,N_16534,N_16515);
or U16731 (N_16731,N_16526,N_16611);
and U16732 (N_16732,N_16503,N_16565);
nand U16733 (N_16733,N_16598,N_16510);
and U16734 (N_16734,N_16554,N_16569);
nand U16735 (N_16735,N_16605,N_16613);
nor U16736 (N_16736,N_16517,N_16592);
nor U16737 (N_16737,N_16597,N_16504);
nor U16738 (N_16738,N_16558,N_16622);
nand U16739 (N_16739,N_16489,N_16614);
or U16740 (N_16740,N_16631,N_16597);
and U16741 (N_16741,N_16534,N_16497);
and U16742 (N_16742,N_16628,N_16515);
nand U16743 (N_16743,N_16529,N_16606);
nand U16744 (N_16744,N_16554,N_16574);
xnor U16745 (N_16745,N_16616,N_16541);
xnor U16746 (N_16746,N_16572,N_16623);
or U16747 (N_16747,N_16498,N_16555);
xnor U16748 (N_16748,N_16521,N_16535);
nor U16749 (N_16749,N_16529,N_16534);
or U16750 (N_16750,N_16590,N_16481);
xor U16751 (N_16751,N_16494,N_16504);
and U16752 (N_16752,N_16494,N_16575);
xor U16753 (N_16753,N_16518,N_16585);
and U16754 (N_16754,N_16481,N_16519);
nor U16755 (N_16755,N_16587,N_16601);
and U16756 (N_16756,N_16480,N_16622);
nor U16757 (N_16757,N_16507,N_16497);
or U16758 (N_16758,N_16565,N_16593);
nand U16759 (N_16759,N_16609,N_16571);
nor U16760 (N_16760,N_16582,N_16578);
xor U16761 (N_16761,N_16611,N_16622);
xnor U16762 (N_16762,N_16507,N_16587);
nor U16763 (N_16763,N_16607,N_16596);
nand U16764 (N_16764,N_16626,N_16617);
or U16765 (N_16765,N_16566,N_16585);
nand U16766 (N_16766,N_16576,N_16581);
nor U16767 (N_16767,N_16619,N_16526);
or U16768 (N_16768,N_16510,N_16638);
nand U16769 (N_16769,N_16497,N_16569);
and U16770 (N_16770,N_16608,N_16480);
or U16771 (N_16771,N_16488,N_16543);
and U16772 (N_16772,N_16538,N_16550);
or U16773 (N_16773,N_16542,N_16616);
or U16774 (N_16774,N_16532,N_16570);
nand U16775 (N_16775,N_16566,N_16604);
or U16776 (N_16776,N_16532,N_16486);
xnor U16777 (N_16777,N_16582,N_16558);
nor U16778 (N_16778,N_16574,N_16623);
nand U16779 (N_16779,N_16528,N_16633);
nand U16780 (N_16780,N_16616,N_16617);
xnor U16781 (N_16781,N_16499,N_16501);
and U16782 (N_16782,N_16619,N_16530);
nand U16783 (N_16783,N_16554,N_16583);
or U16784 (N_16784,N_16485,N_16620);
xnor U16785 (N_16785,N_16528,N_16521);
nand U16786 (N_16786,N_16542,N_16529);
and U16787 (N_16787,N_16608,N_16595);
nand U16788 (N_16788,N_16541,N_16529);
and U16789 (N_16789,N_16606,N_16603);
and U16790 (N_16790,N_16633,N_16499);
and U16791 (N_16791,N_16544,N_16620);
xor U16792 (N_16792,N_16566,N_16628);
nor U16793 (N_16793,N_16544,N_16566);
and U16794 (N_16794,N_16485,N_16628);
nor U16795 (N_16795,N_16486,N_16564);
and U16796 (N_16796,N_16505,N_16555);
nor U16797 (N_16797,N_16592,N_16633);
nand U16798 (N_16798,N_16601,N_16539);
xor U16799 (N_16799,N_16595,N_16527);
nand U16800 (N_16800,N_16712,N_16790);
nand U16801 (N_16801,N_16747,N_16731);
and U16802 (N_16802,N_16703,N_16797);
nand U16803 (N_16803,N_16690,N_16663);
nor U16804 (N_16804,N_16683,N_16646);
nand U16805 (N_16805,N_16693,N_16798);
or U16806 (N_16806,N_16758,N_16732);
xor U16807 (N_16807,N_16686,N_16755);
xor U16808 (N_16808,N_16702,N_16741);
and U16809 (N_16809,N_16724,N_16651);
and U16810 (N_16810,N_16697,N_16761);
xnor U16811 (N_16811,N_16684,N_16753);
xnor U16812 (N_16812,N_16654,N_16767);
xnor U16813 (N_16813,N_16718,N_16783);
or U16814 (N_16814,N_16787,N_16656);
nor U16815 (N_16815,N_16773,N_16657);
and U16816 (N_16816,N_16766,N_16661);
xnor U16817 (N_16817,N_16682,N_16688);
or U16818 (N_16818,N_16770,N_16679);
nor U16819 (N_16819,N_16665,N_16645);
or U16820 (N_16820,N_16799,N_16739);
or U16821 (N_16821,N_16711,N_16659);
nor U16822 (N_16822,N_16658,N_16763);
nor U16823 (N_16823,N_16698,N_16784);
or U16824 (N_16824,N_16676,N_16650);
xor U16825 (N_16825,N_16716,N_16707);
nand U16826 (N_16826,N_16789,N_16653);
nor U16827 (N_16827,N_16668,N_16667);
or U16828 (N_16828,N_16719,N_16735);
and U16829 (N_16829,N_16779,N_16713);
nand U16830 (N_16830,N_16670,N_16700);
xnor U16831 (N_16831,N_16734,N_16788);
xnor U16832 (N_16832,N_16768,N_16647);
or U16833 (N_16833,N_16652,N_16742);
nand U16834 (N_16834,N_16733,N_16728);
xor U16835 (N_16835,N_16662,N_16776);
nand U16836 (N_16836,N_16648,N_16762);
and U16837 (N_16837,N_16705,N_16757);
or U16838 (N_16838,N_16714,N_16642);
nor U16839 (N_16839,N_16793,N_16640);
and U16840 (N_16840,N_16752,N_16738);
or U16841 (N_16841,N_16694,N_16730);
nor U16842 (N_16842,N_16796,N_16759);
nor U16843 (N_16843,N_16740,N_16764);
nand U16844 (N_16844,N_16775,N_16745);
nand U16845 (N_16845,N_16720,N_16710);
nand U16846 (N_16846,N_16737,N_16743);
or U16847 (N_16847,N_16715,N_16687);
and U16848 (N_16848,N_16721,N_16681);
and U16849 (N_16849,N_16795,N_16691);
and U16850 (N_16850,N_16680,N_16785);
or U16851 (N_16851,N_16781,N_16777);
and U16852 (N_16852,N_16655,N_16701);
and U16853 (N_16853,N_16751,N_16750);
nand U16854 (N_16854,N_16772,N_16699);
or U16855 (N_16855,N_16726,N_16671);
xnor U16856 (N_16856,N_16666,N_16774);
and U16857 (N_16857,N_16729,N_16760);
and U16858 (N_16858,N_16749,N_16660);
and U16859 (N_16859,N_16649,N_16669);
and U16860 (N_16860,N_16641,N_16725);
nand U16861 (N_16861,N_16746,N_16717);
nor U16862 (N_16862,N_16794,N_16673);
nor U16863 (N_16863,N_16672,N_16723);
or U16864 (N_16864,N_16689,N_16685);
nor U16865 (N_16865,N_16736,N_16782);
nand U16866 (N_16866,N_16722,N_16674);
or U16867 (N_16867,N_16696,N_16778);
and U16868 (N_16868,N_16695,N_16748);
and U16869 (N_16869,N_16678,N_16704);
and U16870 (N_16870,N_16708,N_16706);
nor U16871 (N_16871,N_16786,N_16643);
and U16872 (N_16872,N_16692,N_16792);
xnor U16873 (N_16873,N_16727,N_16709);
and U16874 (N_16874,N_16677,N_16754);
xnor U16875 (N_16875,N_16675,N_16765);
xor U16876 (N_16876,N_16756,N_16780);
nor U16877 (N_16877,N_16644,N_16769);
or U16878 (N_16878,N_16771,N_16744);
nor U16879 (N_16879,N_16664,N_16791);
xor U16880 (N_16880,N_16659,N_16692);
xor U16881 (N_16881,N_16724,N_16770);
or U16882 (N_16882,N_16689,N_16690);
and U16883 (N_16883,N_16792,N_16759);
and U16884 (N_16884,N_16692,N_16640);
nand U16885 (N_16885,N_16646,N_16673);
or U16886 (N_16886,N_16782,N_16786);
nand U16887 (N_16887,N_16753,N_16772);
nor U16888 (N_16888,N_16760,N_16682);
or U16889 (N_16889,N_16713,N_16745);
xor U16890 (N_16890,N_16760,N_16769);
nor U16891 (N_16891,N_16731,N_16671);
and U16892 (N_16892,N_16723,N_16742);
and U16893 (N_16893,N_16673,N_16692);
xor U16894 (N_16894,N_16778,N_16775);
or U16895 (N_16895,N_16693,N_16683);
nor U16896 (N_16896,N_16747,N_16653);
xnor U16897 (N_16897,N_16786,N_16659);
nand U16898 (N_16898,N_16649,N_16646);
xnor U16899 (N_16899,N_16645,N_16698);
and U16900 (N_16900,N_16671,N_16661);
or U16901 (N_16901,N_16701,N_16694);
nor U16902 (N_16902,N_16650,N_16722);
nor U16903 (N_16903,N_16778,N_16655);
nor U16904 (N_16904,N_16742,N_16690);
and U16905 (N_16905,N_16769,N_16652);
nor U16906 (N_16906,N_16766,N_16646);
or U16907 (N_16907,N_16769,N_16791);
xor U16908 (N_16908,N_16731,N_16785);
and U16909 (N_16909,N_16747,N_16720);
nand U16910 (N_16910,N_16696,N_16724);
xor U16911 (N_16911,N_16661,N_16694);
nor U16912 (N_16912,N_16769,N_16772);
nor U16913 (N_16913,N_16721,N_16727);
xnor U16914 (N_16914,N_16793,N_16649);
or U16915 (N_16915,N_16771,N_16675);
and U16916 (N_16916,N_16748,N_16769);
and U16917 (N_16917,N_16759,N_16753);
and U16918 (N_16918,N_16686,N_16729);
or U16919 (N_16919,N_16764,N_16654);
nor U16920 (N_16920,N_16693,N_16711);
nor U16921 (N_16921,N_16786,N_16761);
or U16922 (N_16922,N_16706,N_16765);
nand U16923 (N_16923,N_16655,N_16752);
nor U16924 (N_16924,N_16716,N_16726);
and U16925 (N_16925,N_16728,N_16648);
xnor U16926 (N_16926,N_16769,N_16740);
and U16927 (N_16927,N_16770,N_16745);
xnor U16928 (N_16928,N_16684,N_16667);
nand U16929 (N_16929,N_16700,N_16660);
nor U16930 (N_16930,N_16650,N_16729);
nand U16931 (N_16931,N_16783,N_16754);
xor U16932 (N_16932,N_16729,N_16655);
and U16933 (N_16933,N_16798,N_16737);
or U16934 (N_16934,N_16704,N_16787);
nand U16935 (N_16935,N_16732,N_16663);
xor U16936 (N_16936,N_16759,N_16770);
nand U16937 (N_16937,N_16671,N_16674);
or U16938 (N_16938,N_16720,N_16716);
nand U16939 (N_16939,N_16715,N_16763);
xor U16940 (N_16940,N_16715,N_16696);
and U16941 (N_16941,N_16640,N_16798);
nor U16942 (N_16942,N_16657,N_16687);
nand U16943 (N_16943,N_16642,N_16782);
or U16944 (N_16944,N_16739,N_16648);
nor U16945 (N_16945,N_16657,N_16778);
nor U16946 (N_16946,N_16645,N_16658);
nor U16947 (N_16947,N_16640,N_16722);
xor U16948 (N_16948,N_16767,N_16698);
and U16949 (N_16949,N_16668,N_16648);
xor U16950 (N_16950,N_16730,N_16653);
xor U16951 (N_16951,N_16695,N_16719);
nand U16952 (N_16952,N_16685,N_16702);
and U16953 (N_16953,N_16668,N_16708);
or U16954 (N_16954,N_16671,N_16787);
and U16955 (N_16955,N_16718,N_16685);
xor U16956 (N_16956,N_16755,N_16649);
nor U16957 (N_16957,N_16751,N_16737);
nand U16958 (N_16958,N_16692,N_16655);
nand U16959 (N_16959,N_16674,N_16786);
and U16960 (N_16960,N_16833,N_16932);
xor U16961 (N_16961,N_16817,N_16958);
xnor U16962 (N_16962,N_16863,N_16922);
or U16963 (N_16963,N_16944,N_16938);
nand U16964 (N_16964,N_16848,N_16930);
nor U16965 (N_16965,N_16891,N_16845);
nor U16966 (N_16966,N_16880,N_16933);
xor U16967 (N_16967,N_16837,N_16950);
nand U16968 (N_16968,N_16844,N_16810);
nand U16969 (N_16969,N_16923,N_16892);
nand U16970 (N_16970,N_16858,N_16947);
nor U16971 (N_16971,N_16818,N_16931);
and U16972 (N_16972,N_16905,N_16815);
and U16973 (N_16973,N_16806,N_16889);
nand U16974 (N_16974,N_16935,N_16926);
xor U16975 (N_16975,N_16825,N_16943);
and U16976 (N_16976,N_16803,N_16915);
nand U16977 (N_16977,N_16809,N_16812);
nand U16978 (N_16978,N_16827,N_16822);
or U16979 (N_16979,N_16885,N_16874);
and U16980 (N_16980,N_16940,N_16916);
and U16981 (N_16981,N_16949,N_16867);
nor U16982 (N_16982,N_16869,N_16925);
xor U16983 (N_16983,N_16824,N_16920);
xnor U16984 (N_16984,N_16904,N_16875);
nor U16985 (N_16985,N_16956,N_16828);
nor U16986 (N_16986,N_16829,N_16847);
and U16987 (N_16987,N_16886,N_16873);
xor U16988 (N_16988,N_16897,N_16850);
and U16989 (N_16989,N_16868,N_16865);
and U16990 (N_16990,N_16813,N_16842);
xnor U16991 (N_16991,N_16910,N_16801);
or U16992 (N_16992,N_16902,N_16857);
nor U16993 (N_16993,N_16859,N_16835);
and U16994 (N_16994,N_16898,N_16942);
nor U16995 (N_16995,N_16823,N_16860);
xor U16996 (N_16996,N_16854,N_16802);
xor U16997 (N_16997,N_16906,N_16929);
or U16998 (N_16998,N_16814,N_16821);
xor U16999 (N_16999,N_16901,N_16877);
nor U17000 (N_17000,N_16861,N_16918);
nand U17001 (N_17001,N_16952,N_16832);
nor U17002 (N_17002,N_16899,N_16917);
xnor U17003 (N_17003,N_16830,N_16941);
and U17004 (N_17004,N_16888,N_16911);
and U17005 (N_17005,N_16800,N_16834);
nand U17006 (N_17006,N_16881,N_16870);
xor U17007 (N_17007,N_16826,N_16909);
or U17008 (N_17008,N_16853,N_16890);
nand U17009 (N_17009,N_16807,N_16840);
xor U17010 (N_17010,N_16937,N_16883);
xnor U17011 (N_17011,N_16864,N_16913);
or U17012 (N_17012,N_16895,N_16862);
xnor U17013 (N_17013,N_16851,N_16804);
or U17014 (N_17014,N_16934,N_16939);
xnor U17015 (N_17015,N_16852,N_16887);
nand U17016 (N_17016,N_16831,N_16819);
and U17017 (N_17017,N_16808,N_16900);
nand U17018 (N_17018,N_16811,N_16953);
xor U17019 (N_17019,N_16876,N_16896);
and U17020 (N_17020,N_16856,N_16843);
xor U17021 (N_17021,N_16927,N_16882);
or U17022 (N_17022,N_16903,N_16841);
nor U17023 (N_17023,N_16849,N_16945);
nor U17024 (N_17024,N_16912,N_16951);
or U17025 (N_17025,N_16893,N_16838);
and U17026 (N_17026,N_16836,N_16907);
or U17027 (N_17027,N_16957,N_16928);
and U17028 (N_17028,N_16846,N_16884);
or U17029 (N_17029,N_16866,N_16955);
and U17030 (N_17030,N_16871,N_16879);
or U17031 (N_17031,N_16959,N_16914);
xnor U17032 (N_17032,N_16924,N_16919);
nand U17033 (N_17033,N_16872,N_16921);
xnor U17034 (N_17034,N_16855,N_16948);
nand U17035 (N_17035,N_16878,N_16820);
xnor U17036 (N_17036,N_16805,N_16816);
and U17037 (N_17037,N_16946,N_16936);
nand U17038 (N_17038,N_16908,N_16894);
or U17039 (N_17039,N_16954,N_16839);
nor U17040 (N_17040,N_16870,N_16894);
and U17041 (N_17041,N_16876,N_16881);
or U17042 (N_17042,N_16820,N_16874);
or U17043 (N_17043,N_16841,N_16945);
xnor U17044 (N_17044,N_16898,N_16894);
nand U17045 (N_17045,N_16835,N_16893);
and U17046 (N_17046,N_16942,N_16830);
and U17047 (N_17047,N_16886,N_16883);
and U17048 (N_17048,N_16945,N_16944);
and U17049 (N_17049,N_16914,N_16895);
and U17050 (N_17050,N_16846,N_16919);
and U17051 (N_17051,N_16804,N_16943);
or U17052 (N_17052,N_16939,N_16905);
and U17053 (N_17053,N_16809,N_16933);
or U17054 (N_17054,N_16943,N_16953);
xor U17055 (N_17055,N_16869,N_16837);
xor U17056 (N_17056,N_16887,N_16862);
nor U17057 (N_17057,N_16869,N_16829);
or U17058 (N_17058,N_16833,N_16805);
nor U17059 (N_17059,N_16842,N_16919);
xnor U17060 (N_17060,N_16939,N_16958);
xnor U17061 (N_17061,N_16947,N_16956);
nand U17062 (N_17062,N_16939,N_16898);
xor U17063 (N_17063,N_16823,N_16885);
or U17064 (N_17064,N_16821,N_16930);
nor U17065 (N_17065,N_16883,N_16800);
nand U17066 (N_17066,N_16871,N_16818);
or U17067 (N_17067,N_16904,N_16935);
nor U17068 (N_17068,N_16871,N_16825);
and U17069 (N_17069,N_16837,N_16876);
nand U17070 (N_17070,N_16945,N_16832);
xor U17071 (N_17071,N_16833,N_16947);
or U17072 (N_17072,N_16841,N_16951);
xnor U17073 (N_17073,N_16838,N_16817);
xor U17074 (N_17074,N_16943,N_16925);
and U17075 (N_17075,N_16896,N_16852);
and U17076 (N_17076,N_16804,N_16929);
nand U17077 (N_17077,N_16812,N_16861);
or U17078 (N_17078,N_16945,N_16865);
nand U17079 (N_17079,N_16865,N_16869);
xor U17080 (N_17080,N_16884,N_16814);
and U17081 (N_17081,N_16933,N_16863);
xor U17082 (N_17082,N_16929,N_16919);
nor U17083 (N_17083,N_16812,N_16822);
or U17084 (N_17084,N_16826,N_16829);
xor U17085 (N_17085,N_16929,N_16818);
or U17086 (N_17086,N_16887,N_16893);
xor U17087 (N_17087,N_16881,N_16891);
and U17088 (N_17088,N_16844,N_16837);
nor U17089 (N_17089,N_16822,N_16852);
or U17090 (N_17090,N_16948,N_16907);
nand U17091 (N_17091,N_16930,N_16956);
xnor U17092 (N_17092,N_16931,N_16894);
nor U17093 (N_17093,N_16949,N_16801);
and U17094 (N_17094,N_16907,N_16812);
nor U17095 (N_17095,N_16816,N_16923);
xor U17096 (N_17096,N_16911,N_16831);
xnor U17097 (N_17097,N_16887,N_16842);
or U17098 (N_17098,N_16822,N_16889);
or U17099 (N_17099,N_16833,N_16918);
and U17100 (N_17100,N_16924,N_16879);
or U17101 (N_17101,N_16918,N_16880);
and U17102 (N_17102,N_16824,N_16845);
or U17103 (N_17103,N_16931,N_16829);
nor U17104 (N_17104,N_16827,N_16878);
nand U17105 (N_17105,N_16918,N_16875);
nand U17106 (N_17106,N_16877,N_16875);
and U17107 (N_17107,N_16899,N_16901);
and U17108 (N_17108,N_16847,N_16949);
xor U17109 (N_17109,N_16910,N_16925);
nor U17110 (N_17110,N_16801,N_16880);
nand U17111 (N_17111,N_16815,N_16865);
xor U17112 (N_17112,N_16839,N_16838);
nand U17113 (N_17113,N_16828,N_16804);
nor U17114 (N_17114,N_16841,N_16856);
xnor U17115 (N_17115,N_16881,N_16807);
xor U17116 (N_17116,N_16830,N_16847);
xnor U17117 (N_17117,N_16839,N_16836);
and U17118 (N_17118,N_16883,N_16846);
or U17119 (N_17119,N_16913,N_16818);
xor U17120 (N_17120,N_17034,N_17017);
nand U17121 (N_17121,N_17070,N_16964);
nor U17122 (N_17122,N_17041,N_17069);
nand U17123 (N_17123,N_17046,N_16995);
or U17124 (N_17124,N_17038,N_17098);
nand U17125 (N_17125,N_16969,N_17044);
nand U17126 (N_17126,N_17092,N_17004);
or U17127 (N_17127,N_16991,N_17081);
and U17128 (N_17128,N_17049,N_17026);
xnor U17129 (N_17129,N_16998,N_16977);
nand U17130 (N_17130,N_17042,N_17007);
nor U17131 (N_17131,N_16961,N_17015);
or U17132 (N_17132,N_17060,N_17100);
nand U17133 (N_17133,N_17101,N_17108);
nand U17134 (N_17134,N_17110,N_17011);
and U17135 (N_17135,N_17102,N_16984);
or U17136 (N_17136,N_17056,N_17071);
and U17137 (N_17137,N_17024,N_17032);
and U17138 (N_17138,N_17096,N_17033);
xor U17139 (N_17139,N_17086,N_17112);
nor U17140 (N_17140,N_17019,N_17057);
xnor U17141 (N_17141,N_17021,N_16973);
or U17142 (N_17142,N_17012,N_17083);
nand U17143 (N_17143,N_17097,N_16994);
nand U17144 (N_17144,N_17115,N_17088);
and U17145 (N_17145,N_17059,N_16989);
nand U17146 (N_17146,N_17029,N_17107);
nand U17147 (N_17147,N_16986,N_16982);
nand U17148 (N_17148,N_17053,N_17077);
and U17149 (N_17149,N_17005,N_17073);
nor U17150 (N_17150,N_17063,N_17016);
nor U17151 (N_17151,N_17025,N_16983);
xnor U17152 (N_17152,N_17043,N_16960);
nand U17153 (N_17153,N_16978,N_17087);
nor U17154 (N_17154,N_17048,N_17091);
or U17155 (N_17155,N_16997,N_17013);
xnor U17156 (N_17156,N_17022,N_16963);
and U17157 (N_17157,N_17018,N_17076);
nand U17158 (N_17158,N_17027,N_16975);
or U17159 (N_17159,N_16967,N_17093);
xnor U17160 (N_17160,N_17020,N_16966);
or U17161 (N_17161,N_16985,N_16976);
xnor U17162 (N_17162,N_17037,N_16970);
or U17163 (N_17163,N_16972,N_17054);
or U17164 (N_17164,N_17062,N_17094);
nand U17165 (N_17165,N_17066,N_16993);
and U17166 (N_17166,N_16992,N_17014);
or U17167 (N_17167,N_17116,N_16968);
nand U17168 (N_17168,N_17010,N_17052);
nand U17169 (N_17169,N_17006,N_17009);
xnor U17170 (N_17170,N_17079,N_17105);
nor U17171 (N_17171,N_17035,N_17106);
nand U17172 (N_17172,N_17065,N_17109);
nand U17173 (N_17173,N_17082,N_17030);
and U17174 (N_17174,N_17068,N_16971);
and U17175 (N_17175,N_17113,N_17114);
or U17176 (N_17176,N_17084,N_17045);
or U17177 (N_17177,N_17078,N_17117);
and U17178 (N_17178,N_16987,N_17090);
or U17179 (N_17179,N_16979,N_17075);
nand U17180 (N_17180,N_17080,N_17040);
or U17181 (N_17181,N_17036,N_16996);
nand U17182 (N_17182,N_17002,N_16981);
or U17183 (N_17183,N_16990,N_16988);
nand U17184 (N_17184,N_17064,N_17072);
nand U17185 (N_17185,N_17095,N_17061);
xnor U17186 (N_17186,N_16974,N_17111);
and U17187 (N_17187,N_17055,N_17085);
xnor U17188 (N_17188,N_17067,N_17118);
and U17189 (N_17189,N_17058,N_17089);
or U17190 (N_17190,N_17104,N_17047);
nor U17191 (N_17191,N_17119,N_17099);
nand U17192 (N_17192,N_17074,N_17031);
xor U17193 (N_17193,N_17023,N_17051);
nor U17194 (N_17194,N_16999,N_17028);
and U17195 (N_17195,N_16962,N_17008);
xor U17196 (N_17196,N_16980,N_17003);
xnor U17197 (N_17197,N_16965,N_17103);
or U17198 (N_17198,N_17039,N_17000);
xor U17199 (N_17199,N_17050,N_17001);
xnor U17200 (N_17200,N_16986,N_17106);
xnor U17201 (N_17201,N_16975,N_17093);
and U17202 (N_17202,N_17112,N_17045);
and U17203 (N_17203,N_17025,N_17007);
nand U17204 (N_17204,N_17041,N_16970);
nor U17205 (N_17205,N_17065,N_17062);
nor U17206 (N_17206,N_17014,N_17042);
nand U17207 (N_17207,N_17028,N_17045);
and U17208 (N_17208,N_17089,N_17027);
or U17209 (N_17209,N_17107,N_17067);
xor U17210 (N_17210,N_17073,N_17088);
nand U17211 (N_17211,N_17100,N_16974);
nand U17212 (N_17212,N_17094,N_16987);
xor U17213 (N_17213,N_16980,N_17012);
and U17214 (N_17214,N_17112,N_17044);
and U17215 (N_17215,N_17012,N_16992);
and U17216 (N_17216,N_17055,N_17108);
and U17217 (N_17217,N_16975,N_17095);
nand U17218 (N_17218,N_16992,N_17041);
nand U17219 (N_17219,N_16989,N_17083);
nand U17220 (N_17220,N_17056,N_17093);
or U17221 (N_17221,N_17051,N_17045);
nor U17222 (N_17222,N_17074,N_17027);
nand U17223 (N_17223,N_17077,N_17073);
or U17224 (N_17224,N_16970,N_17082);
and U17225 (N_17225,N_16985,N_16999);
and U17226 (N_17226,N_16976,N_17009);
nor U17227 (N_17227,N_17033,N_16989);
nand U17228 (N_17228,N_16990,N_17031);
and U17229 (N_17229,N_17025,N_17004);
xor U17230 (N_17230,N_17087,N_16972);
xor U17231 (N_17231,N_17091,N_17011);
and U17232 (N_17232,N_17003,N_16969);
nor U17233 (N_17233,N_17028,N_16981);
nand U17234 (N_17234,N_16968,N_16999);
nor U17235 (N_17235,N_17014,N_17018);
xnor U17236 (N_17236,N_16960,N_16998);
or U17237 (N_17237,N_17070,N_17086);
xor U17238 (N_17238,N_16999,N_17070);
and U17239 (N_17239,N_17039,N_17065);
xor U17240 (N_17240,N_17020,N_17004);
nor U17241 (N_17241,N_17039,N_17008);
xor U17242 (N_17242,N_17047,N_17014);
xor U17243 (N_17243,N_16993,N_16966);
and U17244 (N_17244,N_17004,N_17032);
nor U17245 (N_17245,N_16964,N_17103);
or U17246 (N_17246,N_17045,N_17000);
xnor U17247 (N_17247,N_17041,N_17062);
nor U17248 (N_17248,N_17082,N_17078);
or U17249 (N_17249,N_17012,N_17093);
and U17250 (N_17250,N_17018,N_17069);
or U17251 (N_17251,N_17034,N_17043);
nor U17252 (N_17252,N_17081,N_16974);
nor U17253 (N_17253,N_16992,N_17007);
and U17254 (N_17254,N_16985,N_17041);
xnor U17255 (N_17255,N_17116,N_17010);
nor U17256 (N_17256,N_17114,N_17028);
and U17257 (N_17257,N_17059,N_17044);
xnor U17258 (N_17258,N_17080,N_16982);
or U17259 (N_17259,N_17113,N_17045);
nor U17260 (N_17260,N_17063,N_16964);
nand U17261 (N_17261,N_17061,N_17010);
nand U17262 (N_17262,N_17044,N_17045);
or U17263 (N_17263,N_17084,N_17092);
and U17264 (N_17264,N_17096,N_17113);
nand U17265 (N_17265,N_17046,N_16972);
xnor U17266 (N_17266,N_17117,N_16986);
and U17267 (N_17267,N_17109,N_17115);
or U17268 (N_17268,N_16968,N_16975);
or U17269 (N_17269,N_17068,N_17079);
xor U17270 (N_17270,N_16993,N_17103);
nor U17271 (N_17271,N_17078,N_17043);
nand U17272 (N_17272,N_17078,N_17091);
and U17273 (N_17273,N_16982,N_16998);
nor U17274 (N_17274,N_17067,N_17089);
nand U17275 (N_17275,N_16994,N_17011);
xor U17276 (N_17276,N_17075,N_17113);
nand U17277 (N_17277,N_17072,N_17047);
or U17278 (N_17278,N_17076,N_17100);
xor U17279 (N_17279,N_17081,N_16986);
xnor U17280 (N_17280,N_17263,N_17245);
or U17281 (N_17281,N_17220,N_17266);
nand U17282 (N_17282,N_17185,N_17257);
nor U17283 (N_17283,N_17188,N_17223);
and U17284 (N_17284,N_17249,N_17190);
or U17285 (N_17285,N_17224,N_17212);
xor U17286 (N_17286,N_17125,N_17217);
nand U17287 (N_17287,N_17161,N_17272);
nor U17288 (N_17288,N_17154,N_17186);
and U17289 (N_17289,N_17140,N_17153);
nor U17290 (N_17290,N_17127,N_17221);
nor U17291 (N_17291,N_17279,N_17129);
nor U17292 (N_17292,N_17218,N_17184);
and U17293 (N_17293,N_17171,N_17228);
nor U17294 (N_17294,N_17134,N_17260);
nor U17295 (N_17295,N_17145,N_17152);
nand U17296 (N_17296,N_17143,N_17169);
xnor U17297 (N_17297,N_17243,N_17165);
xnor U17298 (N_17298,N_17175,N_17122);
xnor U17299 (N_17299,N_17139,N_17240);
or U17300 (N_17300,N_17187,N_17268);
nand U17301 (N_17301,N_17180,N_17242);
nor U17302 (N_17302,N_17234,N_17237);
nor U17303 (N_17303,N_17162,N_17121);
nand U17304 (N_17304,N_17136,N_17276);
and U17305 (N_17305,N_17247,N_17201);
or U17306 (N_17306,N_17182,N_17199);
nor U17307 (N_17307,N_17213,N_17258);
xor U17308 (N_17308,N_17254,N_17216);
nand U17309 (N_17309,N_17274,N_17264);
or U17310 (N_17310,N_17196,N_17207);
nor U17311 (N_17311,N_17241,N_17225);
nand U17312 (N_17312,N_17183,N_17233);
xor U17313 (N_17313,N_17273,N_17177);
or U17314 (N_17314,N_17200,N_17230);
nand U17315 (N_17315,N_17146,N_17179);
xor U17316 (N_17316,N_17193,N_17229);
or U17317 (N_17317,N_17168,N_17194);
nor U17318 (N_17318,N_17151,N_17238);
nor U17319 (N_17319,N_17135,N_17141);
and U17320 (N_17320,N_17231,N_17251);
nor U17321 (N_17321,N_17176,N_17227);
nand U17322 (N_17322,N_17261,N_17239);
nor U17323 (N_17323,N_17178,N_17144);
nor U17324 (N_17324,N_17170,N_17157);
xor U17325 (N_17325,N_17275,N_17278);
or U17326 (N_17326,N_17204,N_17156);
nor U17327 (N_17327,N_17222,N_17211);
or U17328 (N_17328,N_17181,N_17205);
xnor U17329 (N_17329,N_17195,N_17214);
or U17330 (N_17330,N_17150,N_17209);
xor U17331 (N_17331,N_17202,N_17248);
or U17332 (N_17332,N_17166,N_17235);
nand U17333 (N_17333,N_17232,N_17277);
nand U17334 (N_17334,N_17206,N_17256);
nor U17335 (N_17335,N_17167,N_17215);
xnor U17336 (N_17336,N_17137,N_17131);
nor U17337 (N_17337,N_17133,N_17226);
nor U17338 (N_17338,N_17123,N_17158);
and U17339 (N_17339,N_17197,N_17148);
xor U17340 (N_17340,N_17126,N_17173);
nand U17341 (N_17341,N_17142,N_17203);
and U17342 (N_17342,N_17130,N_17269);
and U17343 (N_17343,N_17172,N_17163);
and U17344 (N_17344,N_17270,N_17192);
nand U17345 (N_17345,N_17253,N_17236);
nand U17346 (N_17346,N_17124,N_17246);
nor U17347 (N_17347,N_17128,N_17191);
and U17348 (N_17348,N_17208,N_17250);
and U17349 (N_17349,N_17132,N_17259);
and U17350 (N_17350,N_17159,N_17267);
or U17351 (N_17351,N_17160,N_17147);
and U17352 (N_17352,N_17198,N_17210);
xnor U17353 (N_17353,N_17244,N_17155);
xor U17354 (N_17354,N_17149,N_17265);
or U17355 (N_17355,N_17219,N_17271);
and U17356 (N_17356,N_17174,N_17189);
or U17357 (N_17357,N_17120,N_17138);
or U17358 (N_17358,N_17164,N_17262);
nand U17359 (N_17359,N_17255,N_17252);
or U17360 (N_17360,N_17157,N_17249);
nand U17361 (N_17361,N_17235,N_17171);
nand U17362 (N_17362,N_17279,N_17247);
xnor U17363 (N_17363,N_17219,N_17165);
and U17364 (N_17364,N_17234,N_17194);
xor U17365 (N_17365,N_17196,N_17148);
or U17366 (N_17366,N_17274,N_17123);
or U17367 (N_17367,N_17239,N_17273);
nor U17368 (N_17368,N_17192,N_17147);
nand U17369 (N_17369,N_17220,N_17138);
and U17370 (N_17370,N_17273,N_17259);
xor U17371 (N_17371,N_17228,N_17162);
and U17372 (N_17372,N_17218,N_17192);
or U17373 (N_17373,N_17246,N_17224);
nor U17374 (N_17374,N_17223,N_17277);
and U17375 (N_17375,N_17162,N_17225);
xor U17376 (N_17376,N_17145,N_17121);
nor U17377 (N_17377,N_17202,N_17240);
nor U17378 (N_17378,N_17241,N_17123);
nand U17379 (N_17379,N_17264,N_17127);
nand U17380 (N_17380,N_17271,N_17121);
and U17381 (N_17381,N_17269,N_17229);
or U17382 (N_17382,N_17172,N_17248);
nand U17383 (N_17383,N_17199,N_17148);
nor U17384 (N_17384,N_17278,N_17257);
xor U17385 (N_17385,N_17173,N_17147);
xor U17386 (N_17386,N_17133,N_17176);
or U17387 (N_17387,N_17128,N_17165);
xor U17388 (N_17388,N_17205,N_17278);
xor U17389 (N_17389,N_17249,N_17145);
xnor U17390 (N_17390,N_17250,N_17207);
or U17391 (N_17391,N_17272,N_17127);
nor U17392 (N_17392,N_17252,N_17213);
nor U17393 (N_17393,N_17175,N_17196);
and U17394 (N_17394,N_17271,N_17130);
and U17395 (N_17395,N_17255,N_17151);
nand U17396 (N_17396,N_17214,N_17231);
nor U17397 (N_17397,N_17146,N_17178);
xor U17398 (N_17398,N_17266,N_17248);
xnor U17399 (N_17399,N_17255,N_17190);
nand U17400 (N_17400,N_17173,N_17270);
nor U17401 (N_17401,N_17136,N_17259);
xnor U17402 (N_17402,N_17196,N_17143);
nor U17403 (N_17403,N_17227,N_17188);
and U17404 (N_17404,N_17233,N_17192);
or U17405 (N_17405,N_17178,N_17159);
and U17406 (N_17406,N_17204,N_17190);
or U17407 (N_17407,N_17199,N_17224);
or U17408 (N_17408,N_17154,N_17192);
nor U17409 (N_17409,N_17278,N_17166);
or U17410 (N_17410,N_17154,N_17190);
nor U17411 (N_17411,N_17132,N_17270);
and U17412 (N_17412,N_17180,N_17160);
nand U17413 (N_17413,N_17237,N_17260);
and U17414 (N_17414,N_17262,N_17150);
and U17415 (N_17415,N_17126,N_17207);
nor U17416 (N_17416,N_17153,N_17237);
or U17417 (N_17417,N_17187,N_17228);
xor U17418 (N_17418,N_17236,N_17212);
nand U17419 (N_17419,N_17140,N_17197);
nor U17420 (N_17420,N_17199,N_17248);
or U17421 (N_17421,N_17165,N_17257);
and U17422 (N_17422,N_17264,N_17195);
or U17423 (N_17423,N_17154,N_17153);
nor U17424 (N_17424,N_17229,N_17211);
xor U17425 (N_17425,N_17215,N_17162);
and U17426 (N_17426,N_17126,N_17233);
and U17427 (N_17427,N_17159,N_17163);
and U17428 (N_17428,N_17261,N_17255);
nand U17429 (N_17429,N_17185,N_17254);
xnor U17430 (N_17430,N_17130,N_17267);
and U17431 (N_17431,N_17251,N_17267);
nand U17432 (N_17432,N_17163,N_17213);
nand U17433 (N_17433,N_17172,N_17262);
nand U17434 (N_17434,N_17251,N_17229);
or U17435 (N_17435,N_17231,N_17184);
xnor U17436 (N_17436,N_17266,N_17166);
nand U17437 (N_17437,N_17264,N_17204);
and U17438 (N_17438,N_17172,N_17179);
nand U17439 (N_17439,N_17197,N_17132);
or U17440 (N_17440,N_17413,N_17381);
or U17441 (N_17441,N_17368,N_17291);
nor U17442 (N_17442,N_17281,N_17296);
nand U17443 (N_17443,N_17389,N_17285);
nor U17444 (N_17444,N_17283,N_17375);
or U17445 (N_17445,N_17377,N_17379);
nand U17446 (N_17446,N_17304,N_17350);
xnor U17447 (N_17447,N_17403,N_17391);
nor U17448 (N_17448,N_17367,N_17393);
xor U17449 (N_17449,N_17335,N_17373);
xor U17450 (N_17450,N_17394,N_17311);
xor U17451 (N_17451,N_17372,N_17351);
or U17452 (N_17452,N_17356,N_17321);
nor U17453 (N_17453,N_17429,N_17405);
and U17454 (N_17454,N_17435,N_17328);
nand U17455 (N_17455,N_17306,N_17342);
and U17456 (N_17456,N_17308,N_17385);
xor U17457 (N_17457,N_17301,N_17297);
nor U17458 (N_17458,N_17334,N_17417);
nor U17459 (N_17459,N_17387,N_17407);
nor U17460 (N_17460,N_17310,N_17353);
nand U17461 (N_17461,N_17298,N_17333);
and U17462 (N_17462,N_17420,N_17355);
xor U17463 (N_17463,N_17421,N_17300);
or U17464 (N_17464,N_17370,N_17439);
nand U17465 (N_17465,N_17320,N_17436);
nand U17466 (N_17466,N_17325,N_17292);
nor U17467 (N_17467,N_17343,N_17338);
nand U17468 (N_17468,N_17299,N_17388);
or U17469 (N_17469,N_17318,N_17347);
or U17470 (N_17470,N_17401,N_17314);
and U17471 (N_17471,N_17412,N_17319);
or U17472 (N_17472,N_17290,N_17424);
nand U17473 (N_17473,N_17348,N_17309);
and U17474 (N_17474,N_17426,N_17303);
nor U17475 (N_17475,N_17349,N_17400);
and U17476 (N_17476,N_17329,N_17336);
and U17477 (N_17477,N_17317,N_17427);
nor U17478 (N_17478,N_17295,N_17366);
or U17479 (N_17479,N_17418,N_17352);
xor U17480 (N_17480,N_17398,N_17378);
nand U17481 (N_17481,N_17331,N_17287);
and U17482 (N_17482,N_17410,N_17358);
and U17483 (N_17483,N_17392,N_17316);
nand U17484 (N_17484,N_17315,N_17432);
or U17485 (N_17485,N_17293,N_17425);
nand U17486 (N_17486,N_17288,N_17384);
nand U17487 (N_17487,N_17323,N_17402);
nand U17488 (N_17488,N_17344,N_17374);
nor U17489 (N_17489,N_17404,N_17433);
or U17490 (N_17490,N_17364,N_17289);
xor U17491 (N_17491,N_17322,N_17324);
nand U17492 (N_17492,N_17340,N_17302);
and U17493 (N_17493,N_17411,N_17341);
xnor U17494 (N_17494,N_17397,N_17345);
and U17495 (N_17495,N_17339,N_17359);
nor U17496 (N_17496,N_17313,N_17369);
nor U17497 (N_17497,N_17346,N_17337);
and U17498 (N_17498,N_17395,N_17365);
nand U17499 (N_17499,N_17371,N_17419);
or U17500 (N_17500,N_17360,N_17390);
and U17501 (N_17501,N_17286,N_17431);
and U17502 (N_17502,N_17414,N_17330);
and U17503 (N_17503,N_17423,N_17437);
or U17504 (N_17504,N_17280,N_17282);
and U17505 (N_17505,N_17428,N_17363);
or U17506 (N_17506,N_17332,N_17307);
and U17507 (N_17507,N_17284,N_17422);
nand U17508 (N_17508,N_17383,N_17399);
xnor U17509 (N_17509,N_17430,N_17396);
or U17510 (N_17510,N_17382,N_17326);
nand U17511 (N_17511,N_17361,N_17362);
nor U17512 (N_17512,N_17376,N_17434);
nand U17513 (N_17513,N_17354,N_17416);
nand U17514 (N_17514,N_17438,N_17312);
or U17515 (N_17515,N_17386,N_17415);
xnor U17516 (N_17516,N_17294,N_17408);
nand U17517 (N_17517,N_17357,N_17406);
nand U17518 (N_17518,N_17305,N_17409);
nor U17519 (N_17519,N_17327,N_17380);
and U17520 (N_17520,N_17410,N_17345);
nor U17521 (N_17521,N_17286,N_17401);
nand U17522 (N_17522,N_17416,N_17331);
xnor U17523 (N_17523,N_17402,N_17363);
or U17524 (N_17524,N_17301,N_17338);
and U17525 (N_17525,N_17320,N_17391);
and U17526 (N_17526,N_17324,N_17433);
or U17527 (N_17527,N_17363,N_17347);
xor U17528 (N_17528,N_17281,N_17375);
nand U17529 (N_17529,N_17340,N_17310);
nor U17530 (N_17530,N_17368,N_17378);
and U17531 (N_17531,N_17318,N_17304);
nand U17532 (N_17532,N_17339,N_17306);
or U17533 (N_17533,N_17285,N_17430);
nand U17534 (N_17534,N_17377,N_17372);
nand U17535 (N_17535,N_17350,N_17354);
or U17536 (N_17536,N_17418,N_17371);
and U17537 (N_17537,N_17356,N_17382);
nor U17538 (N_17538,N_17327,N_17397);
nand U17539 (N_17539,N_17344,N_17358);
or U17540 (N_17540,N_17366,N_17426);
nor U17541 (N_17541,N_17308,N_17317);
nand U17542 (N_17542,N_17310,N_17375);
or U17543 (N_17543,N_17422,N_17408);
xor U17544 (N_17544,N_17418,N_17318);
nor U17545 (N_17545,N_17348,N_17313);
nor U17546 (N_17546,N_17386,N_17372);
nand U17547 (N_17547,N_17425,N_17282);
nor U17548 (N_17548,N_17340,N_17335);
or U17549 (N_17549,N_17411,N_17283);
xnor U17550 (N_17550,N_17369,N_17321);
nor U17551 (N_17551,N_17431,N_17284);
or U17552 (N_17552,N_17427,N_17315);
nand U17553 (N_17553,N_17292,N_17284);
and U17554 (N_17554,N_17350,N_17317);
nor U17555 (N_17555,N_17309,N_17305);
nor U17556 (N_17556,N_17280,N_17377);
xor U17557 (N_17557,N_17425,N_17382);
or U17558 (N_17558,N_17421,N_17435);
or U17559 (N_17559,N_17373,N_17300);
xor U17560 (N_17560,N_17342,N_17417);
nand U17561 (N_17561,N_17432,N_17436);
xnor U17562 (N_17562,N_17408,N_17362);
and U17563 (N_17563,N_17359,N_17322);
nor U17564 (N_17564,N_17335,N_17388);
xnor U17565 (N_17565,N_17432,N_17394);
or U17566 (N_17566,N_17281,N_17311);
and U17567 (N_17567,N_17280,N_17367);
and U17568 (N_17568,N_17352,N_17307);
and U17569 (N_17569,N_17325,N_17392);
and U17570 (N_17570,N_17406,N_17411);
nand U17571 (N_17571,N_17423,N_17290);
nor U17572 (N_17572,N_17363,N_17280);
nand U17573 (N_17573,N_17414,N_17361);
or U17574 (N_17574,N_17312,N_17343);
nand U17575 (N_17575,N_17381,N_17343);
or U17576 (N_17576,N_17368,N_17420);
nor U17577 (N_17577,N_17384,N_17331);
xor U17578 (N_17578,N_17325,N_17367);
nand U17579 (N_17579,N_17433,N_17339);
nand U17580 (N_17580,N_17301,N_17328);
and U17581 (N_17581,N_17375,N_17348);
nor U17582 (N_17582,N_17283,N_17384);
or U17583 (N_17583,N_17374,N_17429);
or U17584 (N_17584,N_17375,N_17381);
or U17585 (N_17585,N_17325,N_17345);
and U17586 (N_17586,N_17359,N_17361);
nand U17587 (N_17587,N_17286,N_17329);
nor U17588 (N_17588,N_17345,N_17433);
or U17589 (N_17589,N_17344,N_17416);
nor U17590 (N_17590,N_17295,N_17321);
xor U17591 (N_17591,N_17402,N_17349);
nand U17592 (N_17592,N_17317,N_17398);
nand U17593 (N_17593,N_17306,N_17303);
nand U17594 (N_17594,N_17322,N_17349);
nor U17595 (N_17595,N_17355,N_17290);
nor U17596 (N_17596,N_17417,N_17369);
and U17597 (N_17597,N_17354,N_17439);
nand U17598 (N_17598,N_17408,N_17309);
xnor U17599 (N_17599,N_17391,N_17355);
or U17600 (N_17600,N_17500,N_17527);
or U17601 (N_17601,N_17590,N_17454);
and U17602 (N_17602,N_17502,N_17567);
and U17603 (N_17603,N_17518,N_17496);
xor U17604 (N_17604,N_17489,N_17447);
nand U17605 (N_17605,N_17503,N_17596);
nand U17606 (N_17606,N_17461,N_17533);
and U17607 (N_17607,N_17449,N_17467);
and U17608 (N_17608,N_17482,N_17547);
or U17609 (N_17609,N_17591,N_17480);
and U17610 (N_17610,N_17487,N_17508);
or U17611 (N_17611,N_17497,N_17501);
and U17612 (N_17612,N_17522,N_17520);
nand U17613 (N_17613,N_17490,N_17494);
or U17614 (N_17614,N_17488,N_17555);
xnor U17615 (N_17615,N_17452,N_17524);
and U17616 (N_17616,N_17478,N_17512);
nand U17617 (N_17617,N_17481,N_17541);
and U17618 (N_17618,N_17446,N_17571);
xor U17619 (N_17619,N_17580,N_17599);
and U17620 (N_17620,N_17577,N_17451);
xnor U17621 (N_17621,N_17462,N_17558);
and U17622 (N_17622,N_17566,N_17493);
or U17623 (N_17623,N_17573,N_17542);
nor U17624 (N_17624,N_17592,N_17455);
or U17625 (N_17625,N_17549,N_17450);
or U17626 (N_17626,N_17523,N_17597);
nor U17627 (N_17627,N_17507,N_17598);
and U17628 (N_17628,N_17594,N_17540);
or U17629 (N_17629,N_17546,N_17460);
nand U17630 (N_17630,N_17453,N_17543);
xor U17631 (N_17631,N_17544,N_17530);
xor U17632 (N_17632,N_17473,N_17560);
and U17633 (N_17633,N_17516,N_17463);
or U17634 (N_17634,N_17509,N_17554);
nor U17635 (N_17635,N_17528,N_17556);
or U17636 (N_17636,N_17525,N_17498);
and U17637 (N_17637,N_17588,N_17553);
and U17638 (N_17638,N_17484,N_17545);
nand U17639 (N_17639,N_17537,N_17583);
or U17640 (N_17640,N_17557,N_17476);
nand U17641 (N_17641,N_17539,N_17511);
or U17642 (N_17642,N_17477,N_17495);
nor U17643 (N_17643,N_17443,N_17526);
and U17644 (N_17644,N_17587,N_17468);
nor U17645 (N_17645,N_17506,N_17585);
and U17646 (N_17646,N_17538,N_17582);
nand U17647 (N_17647,N_17515,N_17562);
nand U17648 (N_17648,N_17465,N_17589);
xor U17649 (N_17649,N_17445,N_17513);
xor U17650 (N_17650,N_17505,N_17548);
xor U17651 (N_17651,N_17483,N_17442);
nor U17652 (N_17652,N_17440,N_17561);
or U17653 (N_17653,N_17534,N_17579);
or U17654 (N_17654,N_17536,N_17531);
or U17655 (N_17655,N_17471,N_17486);
xor U17656 (N_17656,N_17550,N_17575);
nor U17657 (N_17657,N_17485,N_17458);
nand U17658 (N_17658,N_17569,N_17459);
and U17659 (N_17659,N_17519,N_17535);
and U17660 (N_17660,N_17568,N_17586);
nor U17661 (N_17661,N_17584,N_17551);
nor U17662 (N_17662,N_17576,N_17514);
nor U17663 (N_17663,N_17472,N_17510);
and U17664 (N_17664,N_17504,N_17448);
xnor U17665 (N_17665,N_17529,N_17470);
xnor U17666 (N_17666,N_17574,N_17581);
xor U17667 (N_17667,N_17521,N_17469);
xor U17668 (N_17668,N_17564,N_17578);
nand U17669 (N_17669,N_17491,N_17456);
xor U17670 (N_17670,N_17593,N_17466);
xnor U17671 (N_17671,N_17492,N_17517);
nand U17672 (N_17672,N_17444,N_17475);
or U17673 (N_17673,N_17464,N_17559);
or U17674 (N_17674,N_17457,N_17563);
nor U17675 (N_17675,N_17595,N_17572);
nor U17676 (N_17676,N_17552,N_17499);
nand U17677 (N_17677,N_17565,N_17479);
nand U17678 (N_17678,N_17570,N_17474);
and U17679 (N_17679,N_17441,N_17532);
and U17680 (N_17680,N_17442,N_17475);
nand U17681 (N_17681,N_17471,N_17484);
and U17682 (N_17682,N_17460,N_17468);
or U17683 (N_17683,N_17535,N_17457);
and U17684 (N_17684,N_17457,N_17533);
or U17685 (N_17685,N_17553,N_17568);
nor U17686 (N_17686,N_17460,N_17531);
nor U17687 (N_17687,N_17539,N_17463);
or U17688 (N_17688,N_17533,N_17566);
nor U17689 (N_17689,N_17521,N_17447);
and U17690 (N_17690,N_17521,N_17445);
nand U17691 (N_17691,N_17522,N_17465);
xor U17692 (N_17692,N_17450,N_17532);
nor U17693 (N_17693,N_17440,N_17511);
nand U17694 (N_17694,N_17442,N_17477);
xnor U17695 (N_17695,N_17511,N_17463);
and U17696 (N_17696,N_17519,N_17548);
xor U17697 (N_17697,N_17568,N_17539);
or U17698 (N_17698,N_17498,N_17585);
nor U17699 (N_17699,N_17530,N_17527);
or U17700 (N_17700,N_17473,N_17547);
or U17701 (N_17701,N_17480,N_17479);
and U17702 (N_17702,N_17584,N_17483);
and U17703 (N_17703,N_17543,N_17472);
xnor U17704 (N_17704,N_17483,N_17486);
and U17705 (N_17705,N_17583,N_17460);
and U17706 (N_17706,N_17571,N_17472);
xnor U17707 (N_17707,N_17465,N_17554);
nor U17708 (N_17708,N_17547,N_17480);
and U17709 (N_17709,N_17509,N_17457);
nand U17710 (N_17710,N_17558,N_17499);
nor U17711 (N_17711,N_17516,N_17511);
xnor U17712 (N_17712,N_17584,N_17497);
xor U17713 (N_17713,N_17572,N_17464);
nand U17714 (N_17714,N_17593,N_17535);
nand U17715 (N_17715,N_17452,N_17529);
xnor U17716 (N_17716,N_17478,N_17535);
or U17717 (N_17717,N_17511,N_17595);
nand U17718 (N_17718,N_17445,N_17471);
and U17719 (N_17719,N_17462,N_17480);
and U17720 (N_17720,N_17490,N_17534);
xor U17721 (N_17721,N_17447,N_17480);
xnor U17722 (N_17722,N_17460,N_17515);
xnor U17723 (N_17723,N_17498,N_17559);
xnor U17724 (N_17724,N_17587,N_17551);
xor U17725 (N_17725,N_17444,N_17592);
nand U17726 (N_17726,N_17549,N_17526);
and U17727 (N_17727,N_17588,N_17569);
nor U17728 (N_17728,N_17598,N_17591);
or U17729 (N_17729,N_17485,N_17529);
nor U17730 (N_17730,N_17449,N_17475);
or U17731 (N_17731,N_17484,N_17508);
or U17732 (N_17732,N_17544,N_17574);
xor U17733 (N_17733,N_17518,N_17594);
or U17734 (N_17734,N_17519,N_17449);
or U17735 (N_17735,N_17504,N_17488);
nand U17736 (N_17736,N_17453,N_17535);
nor U17737 (N_17737,N_17455,N_17546);
or U17738 (N_17738,N_17582,N_17463);
or U17739 (N_17739,N_17569,N_17499);
or U17740 (N_17740,N_17555,N_17456);
and U17741 (N_17741,N_17572,N_17580);
and U17742 (N_17742,N_17479,N_17575);
or U17743 (N_17743,N_17592,N_17449);
or U17744 (N_17744,N_17577,N_17475);
nand U17745 (N_17745,N_17480,N_17573);
or U17746 (N_17746,N_17557,N_17457);
xor U17747 (N_17747,N_17510,N_17538);
nor U17748 (N_17748,N_17549,N_17599);
and U17749 (N_17749,N_17504,N_17575);
and U17750 (N_17750,N_17492,N_17538);
nand U17751 (N_17751,N_17493,N_17457);
or U17752 (N_17752,N_17470,N_17526);
nor U17753 (N_17753,N_17531,N_17555);
nor U17754 (N_17754,N_17511,N_17599);
and U17755 (N_17755,N_17583,N_17529);
and U17756 (N_17756,N_17472,N_17483);
nand U17757 (N_17757,N_17516,N_17514);
xnor U17758 (N_17758,N_17556,N_17509);
xnor U17759 (N_17759,N_17510,N_17509);
nand U17760 (N_17760,N_17736,N_17670);
nand U17761 (N_17761,N_17639,N_17717);
or U17762 (N_17762,N_17716,N_17606);
nand U17763 (N_17763,N_17650,N_17728);
and U17764 (N_17764,N_17757,N_17706);
xor U17765 (N_17765,N_17692,N_17647);
nand U17766 (N_17766,N_17707,N_17678);
or U17767 (N_17767,N_17636,N_17630);
and U17768 (N_17768,N_17617,N_17691);
xnor U17769 (N_17769,N_17608,N_17712);
and U17770 (N_17770,N_17690,N_17659);
nor U17771 (N_17771,N_17704,N_17623);
nand U17772 (N_17772,N_17665,N_17758);
nand U17773 (N_17773,N_17609,N_17641);
nor U17774 (N_17774,N_17601,N_17637);
or U17775 (N_17775,N_17616,N_17628);
or U17776 (N_17776,N_17677,N_17751);
xor U17777 (N_17777,N_17612,N_17705);
nand U17778 (N_17778,N_17696,N_17633);
xor U17779 (N_17779,N_17709,N_17687);
xor U17780 (N_17780,N_17664,N_17666);
xnor U17781 (N_17781,N_17721,N_17652);
or U17782 (N_17782,N_17607,N_17715);
and U17783 (N_17783,N_17626,N_17669);
xor U17784 (N_17784,N_17663,N_17725);
nand U17785 (N_17785,N_17688,N_17679);
and U17786 (N_17786,N_17681,N_17673);
nor U17787 (N_17787,N_17735,N_17632);
nor U17788 (N_17788,N_17600,N_17648);
xor U17789 (N_17789,N_17613,N_17610);
xor U17790 (N_17790,N_17711,N_17653);
and U17791 (N_17791,N_17631,N_17710);
or U17792 (N_17792,N_17729,N_17748);
nand U17793 (N_17793,N_17667,N_17733);
nor U17794 (N_17794,N_17702,N_17738);
nand U17795 (N_17795,N_17732,N_17635);
or U17796 (N_17796,N_17755,N_17720);
xor U17797 (N_17797,N_17682,N_17695);
nor U17798 (N_17798,N_17642,N_17689);
nor U17799 (N_17799,N_17743,N_17654);
or U17800 (N_17800,N_17744,N_17713);
nor U17801 (N_17801,N_17605,N_17656);
or U17802 (N_17802,N_17644,N_17620);
xor U17803 (N_17803,N_17741,N_17680);
and U17804 (N_17804,N_17730,N_17724);
xnor U17805 (N_17805,N_17657,N_17752);
nor U17806 (N_17806,N_17671,N_17756);
or U17807 (N_17807,N_17651,N_17753);
and U17808 (N_17808,N_17602,N_17655);
or U17809 (N_17809,N_17649,N_17629);
nand U17810 (N_17810,N_17684,N_17640);
nor U17811 (N_17811,N_17604,N_17634);
nand U17812 (N_17812,N_17615,N_17745);
xor U17813 (N_17813,N_17614,N_17723);
and U17814 (N_17814,N_17746,N_17718);
or U17815 (N_17815,N_17700,N_17672);
nand U17816 (N_17816,N_17611,N_17708);
nand U17817 (N_17817,N_17750,N_17737);
nor U17818 (N_17818,N_17683,N_17747);
xor U17819 (N_17819,N_17675,N_17749);
and U17820 (N_17820,N_17645,N_17638);
xor U17821 (N_17821,N_17739,N_17658);
and U17822 (N_17822,N_17703,N_17661);
nor U17823 (N_17823,N_17719,N_17627);
nand U17824 (N_17824,N_17618,N_17622);
or U17825 (N_17825,N_17603,N_17693);
and U17826 (N_17826,N_17619,N_17759);
and U17827 (N_17827,N_17685,N_17727);
nand U17828 (N_17828,N_17660,N_17699);
nor U17829 (N_17829,N_17621,N_17731);
or U17830 (N_17830,N_17714,N_17643);
xor U17831 (N_17831,N_17698,N_17676);
xor U17832 (N_17832,N_17726,N_17701);
xor U17833 (N_17833,N_17742,N_17734);
nand U17834 (N_17834,N_17668,N_17624);
nand U17835 (N_17835,N_17662,N_17754);
nand U17836 (N_17836,N_17674,N_17625);
nor U17837 (N_17837,N_17686,N_17694);
and U17838 (N_17838,N_17697,N_17740);
xnor U17839 (N_17839,N_17646,N_17722);
and U17840 (N_17840,N_17734,N_17701);
and U17841 (N_17841,N_17623,N_17697);
xnor U17842 (N_17842,N_17675,N_17635);
or U17843 (N_17843,N_17687,N_17625);
xnor U17844 (N_17844,N_17644,N_17660);
nor U17845 (N_17845,N_17736,N_17649);
or U17846 (N_17846,N_17675,N_17730);
nor U17847 (N_17847,N_17641,N_17714);
xnor U17848 (N_17848,N_17730,N_17635);
nor U17849 (N_17849,N_17600,N_17625);
nor U17850 (N_17850,N_17722,N_17674);
or U17851 (N_17851,N_17713,N_17667);
xor U17852 (N_17852,N_17699,N_17623);
nand U17853 (N_17853,N_17743,N_17662);
or U17854 (N_17854,N_17731,N_17724);
or U17855 (N_17855,N_17755,N_17630);
nor U17856 (N_17856,N_17734,N_17603);
or U17857 (N_17857,N_17678,N_17687);
nor U17858 (N_17858,N_17724,N_17654);
and U17859 (N_17859,N_17699,N_17694);
nand U17860 (N_17860,N_17695,N_17603);
nor U17861 (N_17861,N_17749,N_17672);
nand U17862 (N_17862,N_17617,N_17621);
or U17863 (N_17863,N_17642,N_17692);
and U17864 (N_17864,N_17745,N_17614);
nand U17865 (N_17865,N_17615,N_17710);
nor U17866 (N_17866,N_17639,N_17678);
and U17867 (N_17867,N_17722,N_17601);
xor U17868 (N_17868,N_17759,N_17660);
and U17869 (N_17869,N_17605,N_17607);
nand U17870 (N_17870,N_17621,N_17727);
nor U17871 (N_17871,N_17664,N_17711);
or U17872 (N_17872,N_17748,N_17718);
and U17873 (N_17873,N_17681,N_17708);
xnor U17874 (N_17874,N_17758,N_17618);
nand U17875 (N_17875,N_17669,N_17615);
or U17876 (N_17876,N_17745,N_17696);
xor U17877 (N_17877,N_17671,N_17706);
nor U17878 (N_17878,N_17709,N_17723);
nand U17879 (N_17879,N_17705,N_17649);
xnor U17880 (N_17880,N_17746,N_17675);
nand U17881 (N_17881,N_17659,N_17684);
nand U17882 (N_17882,N_17610,N_17646);
nor U17883 (N_17883,N_17602,N_17614);
xor U17884 (N_17884,N_17716,N_17633);
xor U17885 (N_17885,N_17665,N_17754);
nand U17886 (N_17886,N_17667,N_17684);
or U17887 (N_17887,N_17741,N_17704);
and U17888 (N_17888,N_17639,N_17660);
nor U17889 (N_17889,N_17609,N_17683);
and U17890 (N_17890,N_17665,N_17730);
nor U17891 (N_17891,N_17738,N_17622);
and U17892 (N_17892,N_17635,N_17611);
nor U17893 (N_17893,N_17628,N_17703);
xor U17894 (N_17894,N_17639,N_17700);
nor U17895 (N_17895,N_17700,N_17757);
or U17896 (N_17896,N_17753,N_17662);
or U17897 (N_17897,N_17654,N_17607);
nand U17898 (N_17898,N_17708,N_17639);
or U17899 (N_17899,N_17695,N_17719);
and U17900 (N_17900,N_17630,N_17655);
nor U17901 (N_17901,N_17720,N_17737);
nor U17902 (N_17902,N_17675,N_17688);
or U17903 (N_17903,N_17690,N_17717);
nand U17904 (N_17904,N_17726,N_17625);
and U17905 (N_17905,N_17679,N_17632);
nand U17906 (N_17906,N_17627,N_17620);
nor U17907 (N_17907,N_17631,N_17611);
xor U17908 (N_17908,N_17754,N_17705);
or U17909 (N_17909,N_17739,N_17713);
nor U17910 (N_17910,N_17739,N_17656);
nand U17911 (N_17911,N_17689,N_17722);
nand U17912 (N_17912,N_17750,N_17647);
nand U17913 (N_17913,N_17629,N_17683);
or U17914 (N_17914,N_17755,N_17732);
nor U17915 (N_17915,N_17612,N_17685);
nand U17916 (N_17916,N_17651,N_17664);
xnor U17917 (N_17917,N_17677,N_17737);
nand U17918 (N_17918,N_17717,N_17672);
and U17919 (N_17919,N_17726,N_17748);
and U17920 (N_17920,N_17784,N_17818);
or U17921 (N_17921,N_17826,N_17909);
nand U17922 (N_17922,N_17889,N_17894);
or U17923 (N_17923,N_17788,N_17882);
xnor U17924 (N_17924,N_17837,N_17854);
nand U17925 (N_17925,N_17883,N_17798);
xnor U17926 (N_17926,N_17845,N_17918);
nand U17927 (N_17927,N_17906,N_17876);
and U17928 (N_17928,N_17828,N_17783);
nor U17929 (N_17929,N_17851,N_17823);
and U17930 (N_17930,N_17901,N_17770);
nand U17931 (N_17931,N_17919,N_17916);
nand U17932 (N_17932,N_17833,N_17795);
or U17933 (N_17933,N_17879,N_17804);
and U17934 (N_17934,N_17820,N_17810);
xor U17935 (N_17935,N_17830,N_17864);
and U17936 (N_17936,N_17900,N_17819);
xnor U17937 (N_17937,N_17844,N_17785);
and U17938 (N_17938,N_17908,N_17842);
nand U17939 (N_17939,N_17777,N_17898);
or U17940 (N_17940,N_17791,N_17865);
xor U17941 (N_17941,N_17761,N_17884);
nor U17942 (N_17942,N_17829,N_17803);
xnor U17943 (N_17943,N_17780,N_17890);
nand U17944 (N_17944,N_17808,N_17872);
xnor U17945 (N_17945,N_17866,N_17775);
and U17946 (N_17946,N_17764,N_17895);
xnor U17947 (N_17947,N_17873,N_17805);
nor U17948 (N_17948,N_17911,N_17899);
and U17949 (N_17949,N_17847,N_17892);
xor U17950 (N_17950,N_17858,N_17796);
and U17951 (N_17951,N_17836,N_17812);
or U17952 (N_17952,N_17822,N_17886);
nor U17953 (N_17953,N_17806,N_17799);
or U17954 (N_17954,N_17834,N_17779);
and U17955 (N_17955,N_17850,N_17878);
nor U17956 (N_17956,N_17913,N_17902);
xnor U17957 (N_17957,N_17877,N_17825);
and U17958 (N_17958,N_17809,N_17915);
and U17959 (N_17959,N_17811,N_17824);
or U17960 (N_17960,N_17881,N_17793);
nor U17961 (N_17961,N_17766,N_17771);
or U17962 (N_17962,N_17885,N_17816);
and U17963 (N_17963,N_17838,N_17856);
nor U17964 (N_17964,N_17774,N_17807);
or U17965 (N_17965,N_17839,N_17853);
xor U17966 (N_17966,N_17813,N_17868);
xnor U17967 (N_17967,N_17801,N_17831);
xnor U17968 (N_17968,N_17843,N_17893);
nor U17969 (N_17969,N_17773,N_17817);
nand U17970 (N_17970,N_17763,N_17912);
nand U17971 (N_17971,N_17769,N_17914);
and U17972 (N_17972,N_17874,N_17790);
nand U17973 (N_17973,N_17888,N_17863);
or U17974 (N_17974,N_17910,N_17897);
xor U17975 (N_17975,N_17871,N_17841);
and U17976 (N_17976,N_17862,N_17767);
xnor U17977 (N_17977,N_17903,N_17896);
nor U17978 (N_17978,N_17870,N_17887);
nor U17979 (N_17979,N_17765,N_17789);
or U17980 (N_17980,N_17802,N_17800);
xnor U17981 (N_17981,N_17846,N_17760);
nand U17982 (N_17982,N_17797,N_17827);
and U17983 (N_17983,N_17787,N_17782);
nand U17984 (N_17984,N_17907,N_17905);
xor U17985 (N_17985,N_17861,N_17867);
nor U17986 (N_17986,N_17917,N_17778);
nor U17987 (N_17987,N_17786,N_17880);
xor U17988 (N_17988,N_17814,N_17857);
xnor U17989 (N_17989,N_17776,N_17891);
nor U17990 (N_17990,N_17762,N_17904);
and U17991 (N_17991,N_17869,N_17860);
nor U17992 (N_17992,N_17840,N_17815);
xnor U17993 (N_17993,N_17821,N_17768);
nor U17994 (N_17994,N_17848,N_17781);
and U17995 (N_17995,N_17859,N_17835);
nor U17996 (N_17996,N_17875,N_17852);
xor U17997 (N_17997,N_17772,N_17855);
and U17998 (N_17998,N_17794,N_17849);
nand U17999 (N_17999,N_17832,N_17792);
xor U18000 (N_18000,N_17781,N_17826);
and U18001 (N_18001,N_17801,N_17908);
nor U18002 (N_18002,N_17821,N_17797);
nor U18003 (N_18003,N_17910,N_17855);
nor U18004 (N_18004,N_17820,N_17811);
xor U18005 (N_18005,N_17915,N_17840);
nand U18006 (N_18006,N_17850,N_17838);
xnor U18007 (N_18007,N_17773,N_17846);
xor U18008 (N_18008,N_17826,N_17906);
or U18009 (N_18009,N_17834,N_17819);
xnor U18010 (N_18010,N_17893,N_17872);
or U18011 (N_18011,N_17787,N_17832);
xnor U18012 (N_18012,N_17858,N_17875);
nor U18013 (N_18013,N_17837,N_17834);
and U18014 (N_18014,N_17909,N_17900);
nor U18015 (N_18015,N_17801,N_17890);
xnor U18016 (N_18016,N_17808,N_17828);
and U18017 (N_18017,N_17844,N_17836);
xnor U18018 (N_18018,N_17806,N_17900);
nor U18019 (N_18019,N_17844,N_17814);
or U18020 (N_18020,N_17883,N_17774);
and U18021 (N_18021,N_17861,N_17787);
nand U18022 (N_18022,N_17845,N_17863);
or U18023 (N_18023,N_17803,N_17877);
and U18024 (N_18024,N_17861,N_17839);
xnor U18025 (N_18025,N_17880,N_17863);
nand U18026 (N_18026,N_17873,N_17903);
xnor U18027 (N_18027,N_17814,N_17872);
or U18028 (N_18028,N_17904,N_17799);
xor U18029 (N_18029,N_17813,N_17878);
xnor U18030 (N_18030,N_17785,N_17890);
nand U18031 (N_18031,N_17864,N_17857);
nor U18032 (N_18032,N_17864,N_17842);
nand U18033 (N_18033,N_17879,N_17782);
nand U18034 (N_18034,N_17823,N_17829);
nand U18035 (N_18035,N_17825,N_17900);
or U18036 (N_18036,N_17797,N_17906);
nand U18037 (N_18037,N_17917,N_17834);
nor U18038 (N_18038,N_17818,N_17761);
and U18039 (N_18039,N_17842,N_17811);
or U18040 (N_18040,N_17881,N_17790);
nor U18041 (N_18041,N_17850,N_17819);
nor U18042 (N_18042,N_17829,N_17789);
nand U18043 (N_18043,N_17898,N_17827);
nand U18044 (N_18044,N_17843,N_17763);
nand U18045 (N_18045,N_17798,N_17844);
or U18046 (N_18046,N_17801,N_17778);
nand U18047 (N_18047,N_17783,N_17851);
or U18048 (N_18048,N_17856,N_17817);
or U18049 (N_18049,N_17828,N_17880);
or U18050 (N_18050,N_17762,N_17812);
and U18051 (N_18051,N_17853,N_17766);
nand U18052 (N_18052,N_17866,N_17800);
and U18053 (N_18053,N_17830,N_17784);
or U18054 (N_18054,N_17849,N_17807);
and U18055 (N_18055,N_17915,N_17771);
nor U18056 (N_18056,N_17764,N_17768);
nor U18057 (N_18057,N_17871,N_17852);
xnor U18058 (N_18058,N_17832,N_17861);
xnor U18059 (N_18059,N_17914,N_17879);
or U18060 (N_18060,N_17866,N_17792);
or U18061 (N_18061,N_17828,N_17795);
xnor U18062 (N_18062,N_17916,N_17854);
nand U18063 (N_18063,N_17800,N_17796);
nand U18064 (N_18064,N_17784,N_17877);
xnor U18065 (N_18065,N_17852,N_17903);
nand U18066 (N_18066,N_17780,N_17893);
nand U18067 (N_18067,N_17872,N_17795);
nor U18068 (N_18068,N_17884,N_17899);
nor U18069 (N_18069,N_17887,N_17808);
xnor U18070 (N_18070,N_17861,N_17845);
or U18071 (N_18071,N_17882,N_17792);
nor U18072 (N_18072,N_17841,N_17870);
or U18073 (N_18073,N_17908,N_17782);
and U18074 (N_18074,N_17809,N_17760);
nand U18075 (N_18075,N_17854,N_17841);
nor U18076 (N_18076,N_17870,N_17764);
nor U18077 (N_18077,N_17761,N_17913);
nor U18078 (N_18078,N_17919,N_17877);
nand U18079 (N_18079,N_17914,N_17852);
xor U18080 (N_18080,N_17924,N_17961);
xor U18081 (N_18081,N_17978,N_17922);
nor U18082 (N_18082,N_17995,N_18029);
nor U18083 (N_18083,N_17998,N_17957);
nand U18084 (N_18084,N_18045,N_17987);
xnor U18085 (N_18085,N_18043,N_17942);
or U18086 (N_18086,N_17992,N_17980);
nor U18087 (N_18087,N_17936,N_18011);
nand U18088 (N_18088,N_17950,N_18009);
nand U18089 (N_18089,N_17968,N_18044);
xor U18090 (N_18090,N_18049,N_17958);
or U18091 (N_18091,N_18066,N_17990);
and U18092 (N_18092,N_17943,N_18027);
nand U18093 (N_18093,N_17974,N_18077);
and U18094 (N_18094,N_18040,N_18016);
or U18095 (N_18095,N_18006,N_18076);
nor U18096 (N_18096,N_17986,N_17929);
and U18097 (N_18097,N_18038,N_18053);
or U18098 (N_18098,N_18072,N_18050);
nand U18099 (N_18099,N_18014,N_17948);
xor U18100 (N_18100,N_17983,N_18051);
nor U18101 (N_18101,N_17933,N_17991);
or U18102 (N_18102,N_17930,N_18054);
or U18103 (N_18103,N_17952,N_17920);
nand U18104 (N_18104,N_18058,N_18039);
xor U18105 (N_18105,N_18060,N_18018);
or U18106 (N_18106,N_17994,N_17993);
and U18107 (N_18107,N_18033,N_17937);
xnor U18108 (N_18108,N_18057,N_17956);
nand U18109 (N_18109,N_17982,N_18069);
nor U18110 (N_18110,N_18059,N_18005);
nor U18111 (N_18111,N_17931,N_18065);
xnor U18112 (N_18112,N_18022,N_18001);
nand U18113 (N_18113,N_17947,N_17935);
nand U18114 (N_18114,N_18064,N_18015);
nand U18115 (N_18115,N_18048,N_17944);
xnor U18116 (N_18116,N_18010,N_18012);
and U18117 (N_18117,N_17939,N_17928);
xor U18118 (N_18118,N_17934,N_18078);
or U18119 (N_18119,N_17989,N_18028);
or U18120 (N_18120,N_17985,N_17945);
nor U18121 (N_18121,N_18056,N_18023);
and U18122 (N_18122,N_17964,N_18024);
xor U18123 (N_18123,N_17977,N_17938);
nand U18124 (N_18124,N_18032,N_17953);
xnor U18125 (N_18125,N_18073,N_17962);
nand U18126 (N_18126,N_17960,N_17997);
nand U18127 (N_18127,N_17951,N_17966);
or U18128 (N_18128,N_17925,N_18074);
xnor U18129 (N_18129,N_18000,N_18067);
xnor U18130 (N_18130,N_18025,N_17976);
nand U18131 (N_18131,N_18035,N_18004);
or U18132 (N_18132,N_17965,N_18047);
and U18133 (N_18133,N_17996,N_18046);
xnor U18134 (N_18134,N_17979,N_17926);
nor U18135 (N_18135,N_17975,N_18030);
and U18136 (N_18136,N_18042,N_17955);
or U18137 (N_18137,N_17969,N_18070);
nor U18138 (N_18138,N_18055,N_18007);
nand U18139 (N_18139,N_18021,N_17927);
nand U18140 (N_18140,N_18003,N_18034);
nor U18141 (N_18141,N_17988,N_17923);
nand U18142 (N_18142,N_18020,N_18052);
nor U18143 (N_18143,N_18031,N_17999);
nor U18144 (N_18144,N_18075,N_17954);
xor U18145 (N_18145,N_17973,N_18063);
xor U18146 (N_18146,N_18026,N_18041);
or U18147 (N_18147,N_17932,N_17970);
xnor U18148 (N_18148,N_18008,N_17921);
and U18149 (N_18149,N_17949,N_17984);
xnor U18150 (N_18150,N_17946,N_17940);
nor U18151 (N_18151,N_17972,N_17967);
nor U18152 (N_18152,N_18062,N_18079);
and U18153 (N_18153,N_18061,N_17963);
nand U18154 (N_18154,N_18071,N_18036);
and U18155 (N_18155,N_17971,N_17981);
nand U18156 (N_18156,N_18037,N_18068);
xor U18157 (N_18157,N_18017,N_17959);
xnor U18158 (N_18158,N_18013,N_17941);
xnor U18159 (N_18159,N_18019,N_18002);
or U18160 (N_18160,N_18066,N_17987);
nand U18161 (N_18161,N_17942,N_18061);
xor U18162 (N_18162,N_18003,N_18067);
nand U18163 (N_18163,N_18028,N_17979);
nor U18164 (N_18164,N_18041,N_18005);
or U18165 (N_18165,N_18068,N_17964);
nor U18166 (N_18166,N_17922,N_17988);
nand U18167 (N_18167,N_18001,N_17977);
and U18168 (N_18168,N_17924,N_17995);
and U18169 (N_18169,N_18037,N_18018);
xor U18170 (N_18170,N_17931,N_17955);
nor U18171 (N_18171,N_17925,N_18030);
and U18172 (N_18172,N_18053,N_18013);
xnor U18173 (N_18173,N_17974,N_17959);
nor U18174 (N_18174,N_18035,N_18007);
nand U18175 (N_18175,N_17969,N_17990);
nor U18176 (N_18176,N_17980,N_18051);
or U18177 (N_18177,N_18038,N_18014);
or U18178 (N_18178,N_17966,N_18051);
or U18179 (N_18179,N_17937,N_17970);
xor U18180 (N_18180,N_17988,N_17940);
or U18181 (N_18181,N_17966,N_17929);
nand U18182 (N_18182,N_18051,N_18067);
xor U18183 (N_18183,N_17974,N_17937);
nor U18184 (N_18184,N_17975,N_18006);
xnor U18185 (N_18185,N_18073,N_18054);
nand U18186 (N_18186,N_17981,N_18031);
nand U18187 (N_18187,N_17933,N_17936);
nor U18188 (N_18188,N_18058,N_18000);
nand U18189 (N_18189,N_18015,N_17985);
or U18190 (N_18190,N_17947,N_17933);
xor U18191 (N_18191,N_17994,N_18075);
nor U18192 (N_18192,N_18050,N_17944);
or U18193 (N_18193,N_17952,N_17955);
nor U18194 (N_18194,N_17974,N_17936);
nor U18195 (N_18195,N_17981,N_18041);
nor U18196 (N_18196,N_18009,N_17971);
nand U18197 (N_18197,N_18024,N_18073);
or U18198 (N_18198,N_18022,N_18028);
xnor U18199 (N_18199,N_17930,N_18033);
and U18200 (N_18200,N_17984,N_18052);
nand U18201 (N_18201,N_17942,N_18026);
and U18202 (N_18202,N_17934,N_18077);
xor U18203 (N_18203,N_17977,N_18068);
and U18204 (N_18204,N_17982,N_18017);
nor U18205 (N_18205,N_17935,N_17948);
nand U18206 (N_18206,N_18054,N_18028);
or U18207 (N_18207,N_17922,N_18064);
nand U18208 (N_18208,N_18007,N_17990);
or U18209 (N_18209,N_17928,N_17973);
xor U18210 (N_18210,N_18059,N_18032);
and U18211 (N_18211,N_17995,N_17996);
nor U18212 (N_18212,N_18007,N_17966);
nand U18213 (N_18213,N_18037,N_17969);
nor U18214 (N_18214,N_18015,N_18051);
nor U18215 (N_18215,N_17924,N_17945);
and U18216 (N_18216,N_17986,N_17923);
xor U18217 (N_18217,N_18019,N_17976);
or U18218 (N_18218,N_17969,N_18059);
nor U18219 (N_18219,N_18028,N_17930);
or U18220 (N_18220,N_18008,N_18060);
and U18221 (N_18221,N_17925,N_18065);
xor U18222 (N_18222,N_18056,N_18011);
nand U18223 (N_18223,N_17920,N_18029);
or U18224 (N_18224,N_17986,N_18030);
nand U18225 (N_18225,N_18073,N_17940);
nand U18226 (N_18226,N_18073,N_17997);
nand U18227 (N_18227,N_17965,N_17998);
or U18228 (N_18228,N_17977,N_18032);
or U18229 (N_18229,N_17984,N_17956);
or U18230 (N_18230,N_17927,N_17986);
or U18231 (N_18231,N_17958,N_18027);
xor U18232 (N_18232,N_17944,N_17948);
or U18233 (N_18233,N_17986,N_18064);
or U18234 (N_18234,N_17969,N_18036);
xor U18235 (N_18235,N_18029,N_18060);
or U18236 (N_18236,N_17946,N_17933);
xnor U18237 (N_18237,N_17969,N_18000);
nand U18238 (N_18238,N_18060,N_17976);
or U18239 (N_18239,N_18046,N_18041);
and U18240 (N_18240,N_18098,N_18208);
and U18241 (N_18241,N_18193,N_18147);
xor U18242 (N_18242,N_18214,N_18215);
xor U18243 (N_18243,N_18159,N_18239);
nand U18244 (N_18244,N_18126,N_18157);
xnor U18245 (N_18245,N_18174,N_18150);
and U18246 (N_18246,N_18109,N_18183);
nor U18247 (N_18247,N_18084,N_18105);
nor U18248 (N_18248,N_18235,N_18182);
xnor U18249 (N_18249,N_18082,N_18170);
xor U18250 (N_18250,N_18111,N_18094);
or U18251 (N_18251,N_18127,N_18232);
and U18252 (N_18252,N_18162,N_18196);
nand U18253 (N_18253,N_18176,N_18149);
xnor U18254 (N_18254,N_18224,N_18124);
and U18255 (N_18255,N_18095,N_18163);
and U18256 (N_18256,N_18188,N_18123);
nor U18257 (N_18257,N_18083,N_18093);
and U18258 (N_18258,N_18220,N_18230);
and U18259 (N_18259,N_18190,N_18142);
xor U18260 (N_18260,N_18089,N_18091);
and U18261 (N_18261,N_18146,N_18186);
and U18262 (N_18262,N_18228,N_18097);
or U18263 (N_18263,N_18227,N_18130);
and U18264 (N_18264,N_18134,N_18209);
xnor U18265 (N_18265,N_18202,N_18114);
or U18266 (N_18266,N_18087,N_18108);
and U18267 (N_18267,N_18191,N_18116);
xnor U18268 (N_18268,N_18184,N_18086);
nand U18269 (N_18269,N_18212,N_18198);
xor U18270 (N_18270,N_18177,N_18129);
nand U18271 (N_18271,N_18160,N_18166);
nand U18272 (N_18272,N_18122,N_18219);
nor U18273 (N_18273,N_18237,N_18136);
xor U18274 (N_18274,N_18236,N_18180);
nor U18275 (N_18275,N_18225,N_18164);
and U18276 (N_18276,N_18155,N_18156);
xnor U18277 (N_18277,N_18106,N_18113);
and U18278 (N_18278,N_18197,N_18102);
nor U18279 (N_18279,N_18195,N_18143);
xnor U18280 (N_18280,N_18119,N_18107);
xor U18281 (N_18281,N_18158,N_18213);
nand U18282 (N_18282,N_18238,N_18167);
xor U18283 (N_18283,N_18144,N_18226);
xnor U18284 (N_18284,N_18231,N_18148);
nor U18285 (N_18285,N_18117,N_18088);
and U18286 (N_18286,N_18175,N_18118);
xnor U18287 (N_18287,N_18194,N_18112);
nor U18288 (N_18288,N_18135,N_18218);
nor U18289 (N_18289,N_18168,N_18133);
nor U18290 (N_18290,N_18203,N_18090);
nor U18291 (N_18291,N_18181,N_18206);
nor U18292 (N_18292,N_18085,N_18178);
xnor U18293 (N_18293,N_18165,N_18145);
or U18294 (N_18294,N_18101,N_18125);
and U18295 (N_18295,N_18161,N_18233);
nand U18296 (N_18296,N_18140,N_18179);
nand U18297 (N_18297,N_18121,N_18120);
xor U18298 (N_18298,N_18110,N_18081);
xor U18299 (N_18299,N_18137,N_18173);
and U18300 (N_18300,N_18210,N_18216);
xnor U18301 (N_18301,N_18103,N_18096);
xnor U18302 (N_18302,N_18100,N_18234);
and U18303 (N_18303,N_18200,N_18207);
xnor U18304 (N_18304,N_18132,N_18222);
or U18305 (N_18305,N_18080,N_18115);
xnor U18306 (N_18306,N_18139,N_18169);
and U18307 (N_18307,N_18092,N_18099);
nand U18308 (N_18308,N_18128,N_18229);
or U18309 (N_18309,N_18211,N_18154);
xnor U18310 (N_18310,N_18221,N_18152);
xnor U18311 (N_18311,N_18205,N_18217);
nor U18312 (N_18312,N_18192,N_18187);
nor U18313 (N_18313,N_18171,N_18204);
nand U18314 (N_18314,N_18189,N_18153);
nor U18315 (N_18315,N_18185,N_18201);
xnor U18316 (N_18316,N_18131,N_18141);
and U18317 (N_18317,N_18151,N_18223);
nor U18318 (N_18318,N_18172,N_18138);
nor U18319 (N_18319,N_18199,N_18104);
and U18320 (N_18320,N_18157,N_18158);
nor U18321 (N_18321,N_18217,N_18166);
or U18322 (N_18322,N_18106,N_18092);
nand U18323 (N_18323,N_18235,N_18209);
nand U18324 (N_18324,N_18094,N_18081);
nand U18325 (N_18325,N_18114,N_18156);
and U18326 (N_18326,N_18108,N_18148);
or U18327 (N_18327,N_18115,N_18117);
nand U18328 (N_18328,N_18225,N_18101);
xor U18329 (N_18329,N_18210,N_18186);
nor U18330 (N_18330,N_18191,N_18225);
and U18331 (N_18331,N_18104,N_18083);
or U18332 (N_18332,N_18116,N_18095);
nand U18333 (N_18333,N_18238,N_18105);
nand U18334 (N_18334,N_18155,N_18173);
and U18335 (N_18335,N_18082,N_18083);
or U18336 (N_18336,N_18225,N_18088);
xnor U18337 (N_18337,N_18110,N_18093);
xor U18338 (N_18338,N_18093,N_18190);
nor U18339 (N_18339,N_18170,N_18161);
nand U18340 (N_18340,N_18106,N_18237);
and U18341 (N_18341,N_18225,N_18081);
nor U18342 (N_18342,N_18238,N_18226);
nor U18343 (N_18343,N_18209,N_18094);
and U18344 (N_18344,N_18100,N_18125);
nor U18345 (N_18345,N_18166,N_18095);
nand U18346 (N_18346,N_18186,N_18126);
and U18347 (N_18347,N_18137,N_18091);
xnor U18348 (N_18348,N_18199,N_18095);
nor U18349 (N_18349,N_18194,N_18124);
and U18350 (N_18350,N_18220,N_18214);
nor U18351 (N_18351,N_18231,N_18111);
nor U18352 (N_18352,N_18181,N_18133);
nor U18353 (N_18353,N_18205,N_18144);
nand U18354 (N_18354,N_18200,N_18131);
and U18355 (N_18355,N_18147,N_18126);
xor U18356 (N_18356,N_18233,N_18173);
or U18357 (N_18357,N_18108,N_18226);
nand U18358 (N_18358,N_18236,N_18158);
nor U18359 (N_18359,N_18212,N_18148);
nor U18360 (N_18360,N_18145,N_18223);
nand U18361 (N_18361,N_18116,N_18142);
and U18362 (N_18362,N_18080,N_18113);
or U18363 (N_18363,N_18111,N_18134);
nor U18364 (N_18364,N_18168,N_18084);
nand U18365 (N_18365,N_18082,N_18229);
and U18366 (N_18366,N_18111,N_18172);
nand U18367 (N_18367,N_18183,N_18090);
nand U18368 (N_18368,N_18186,N_18085);
and U18369 (N_18369,N_18118,N_18171);
nand U18370 (N_18370,N_18178,N_18187);
nand U18371 (N_18371,N_18142,N_18154);
or U18372 (N_18372,N_18162,N_18155);
xor U18373 (N_18373,N_18168,N_18127);
or U18374 (N_18374,N_18197,N_18109);
or U18375 (N_18375,N_18124,N_18139);
and U18376 (N_18376,N_18132,N_18202);
nor U18377 (N_18377,N_18217,N_18103);
nor U18378 (N_18378,N_18110,N_18091);
and U18379 (N_18379,N_18230,N_18103);
nand U18380 (N_18380,N_18178,N_18121);
nor U18381 (N_18381,N_18218,N_18228);
nor U18382 (N_18382,N_18096,N_18228);
nor U18383 (N_18383,N_18199,N_18111);
or U18384 (N_18384,N_18164,N_18214);
nor U18385 (N_18385,N_18191,N_18220);
or U18386 (N_18386,N_18163,N_18227);
nand U18387 (N_18387,N_18140,N_18155);
nor U18388 (N_18388,N_18128,N_18111);
nor U18389 (N_18389,N_18121,N_18152);
and U18390 (N_18390,N_18128,N_18085);
or U18391 (N_18391,N_18201,N_18133);
and U18392 (N_18392,N_18222,N_18131);
or U18393 (N_18393,N_18107,N_18147);
nand U18394 (N_18394,N_18176,N_18238);
nand U18395 (N_18395,N_18138,N_18161);
nand U18396 (N_18396,N_18153,N_18203);
nor U18397 (N_18397,N_18151,N_18142);
nor U18398 (N_18398,N_18178,N_18214);
xnor U18399 (N_18399,N_18233,N_18239);
xor U18400 (N_18400,N_18288,N_18280);
xnor U18401 (N_18401,N_18359,N_18241);
xnor U18402 (N_18402,N_18328,N_18341);
nand U18403 (N_18403,N_18388,N_18383);
nor U18404 (N_18404,N_18308,N_18346);
or U18405 (N_18405,N_18330,N_18264);
nand U18406 (N_18406,N_18278,N_18266);
or U18407 (N_18407,N_18309,N_18372);
and U18408 (N_18408,N_18327,N_18257);
or U18409 (N_18409,N_18331,N_18384);
or U18410 (N_18410,N_18281,N_18302);
and U18411 (N_18411,N_18333,N_18276);
and U18412 (N_18412,N_18377,N_18268);
xnor U18413 (N_18413,N_18378,N_18256);
and U18414 (N_18414,N_18303,N_18322);
nor U18415 (N_18415,N_18269,N_18368);
nor U18416 (N_18416,N_18299,N_18289);
xnor U18417 (N_18417,N_18332,N_18393);
nand U18418 (N_18418,N_18387,N_18274);
nand U18419 (N_18419,N_18389,N_18287);
nand U18420 (N_18420,N_18340,N_18248);
nand U18421 (N_18421,N_18381,N_18375);
nor U18422 (N_18422,N_18334,N_18360);
xnor U18423 (N_18423,N_18348,N_18324);
and U18424 (N_18424,N_18282,N_18295);
nand U18425 (N_18425,N_18316,N_18312);
or U18426 (N_18426,N_18323,N_18350);
or U18427 (N_18427,N_18321,N_18313);
nand U18428 (N_18428,N_18240,N_18272);
and U18429 (N_18429,N_18314,N_18292);
xor U18430 (N_18430,N_18335,N_18307);
nand U18431 (N_18431,N_18310,N_18349);
nor U18432 (N_18432,N_18365,N_18343);
nor U18433 (N_18433,N_18339,N_18277);
nor U18434 (N_18434,N_18270,N_18391);
or U18435 (N_18435,N_18263,N_18364);
and U18436 (N_18436,N_18338,N_18265);
xor U18437 (N_18437,N_18301,N_18311);
or U18438 (N_18438,N_18242,N_18394);
xor U18439 (N_18439,N_18261,N_18318);
and U18440 (N_18440,N_18345,N_18271);
or U18441 (N_18441,N_18247,N_18317);
xor U18442 (N_18442,N_18344,N_18279);
xor U18443 (N_18443,N_18275,N_18357);
xnor U18444 (N_18444,N_18351,N_18329);
xnor U18445 (N_18445,N_18315,N_18304);
or U18446 (N_18446,N_18260,N_18320);
nand U18447 (N_18447,N_18252,N_18379);
xnor U18448 (N_18448,N_18246,N_18397);
nand U18449 (N_18449,N_18366,N_18306);
nand U18450 (N_18450,N_18273,N_18291);
nor U18451 (N_18451,N_18262,N_18285);
xnor U18452 (N_18452,N_18258,N_18267);
nor U18453 (N_18453,N_18358,N_18298);
and U18454 (N_18454,N_18367,N_18290);
or U18455 (N_18455,N_18244,N_18385);
nor U18456 (N_18456,N_18392,N_18243);
xnor U18457 (N_18457,N_18370,N_18305);
or U18458 (N_18458,N_18380,N_18259);
nor U18459 (N_18459,N_18245,N_18250);
or U18460 (N_18460,N_18326,N_18337);
nand U18461 (N_18461,N_18353,N_18355);
and U18462 (N_18462,N_18374,N_18347);
nand U18463 (N_18463,N_18255,N_18373);
nand U18464 (N_18464,N_18356,N_18382);
nor U18465 (N_18465,N_18386,N_18376);
and U18466 (N_18466,N_18399,N_18293);
or U18467 (N_18467,N_18297,N_18319);
nand U18468 (N_18468,N_18254,N_18286);
or U18469 (N_18469,N_18390,N_18336);
and U18470 (N_18470,N_18249,N_18342);
nor U18471 (N_18471,N_18352,N_18294);
or U18472 (N_18472,N_18296,N_18251);
and U18473 (N_18473,N_18361,N_18369);
or U18474 (N_18474,N_18325,N_18371);
nor U18475 (N_18475,N_18396,N_18398);
xnor U18476 (N_18476,N_18283,N_18354);
nor U18477 (N_18477,N_18284,N_18253);
nor U18478 (N_18478,N_18363,N_18395);
nor U18479 (N_18479,N_18300,N_18362);
and U18480 (N_18480,N_18329,N_18249);
xor U18481 (N_18481,N_18368,N_18265);
xnor U18482 (N_18482,N_18310,N_18326);
or U18483 (N_18483,N_18369,N_18346);
nand U18484 (N_18484,N_18289,N_18380);
nand U18485 (N_18485,N_18266,N_18299);
nor U18486 (N_18486,N_18360,N_18389);
and U18487 (N_18487,N_18272,N_18387);
and U18488 (N_18488,N_18346,N_18327);
and U18489 (N_18489,N_18288,N_18297);
nor U18490 (N_18490,N_18313,N_18281);
nor U18491 (N_18491,N_18360,N_18291);
and U18492 (N_18492,N_18367,N_18322);
xnor U18493 (N_18493,N_18256,N_18364);
and U18494 (N_18494,N_18251,N_18367);
xor U18495 (N_18495,N_18307,N_18395);
xnor U18496 (N_18496,N_18266,N_18275);
or U18497 (N_18497,N_18388,N_18260);
nand U18498 (N_18498,N_18339,N_18320);
or U18499 (N_18499,N_18344,N_18394);
xor U18500 (N_18500,N_18256,N_18309);
xor U18501 (N_18501,N_18359,N_18372);
nor U18502 (N_18502,N_18283,N_18301);
and U18503 (N_18503,N_18291,N_18270);
xnor U18504 (N_18504,N_18383,N_18245);
nor U18505 (N_18505,N_18245,N_18387);
xor U18506 (N_18506,N_18376,N_18300);
and U18507 (N_18507,N_18351,N_18274);
nor U18508 (N_18508,N_18325,N_18343);
or U18509 (N_18509,N_18300,N_18379);
xnor U18510 (N_18510,N_18305,N_18350);
or U18511 (N_18511,N_18322,N_18363);
and U18512 (N_18512,N_18386,N_18309);
nand U18513 (N_18513,N_18289,N_18337);
and U18514 (N_18514,N_18338,N_18300);
nand U18515 (N_18515,N_18300,N_18299);
nand U18516 (N_18516,N_18337,N_18294);
or U18517 (N_18517,N_18366,N_18263);
nand U18518 (N_18518,N_18374,N_18250);
nand U18519 (N_18519,N_18246,N_18248);
xnor U18520 (N_18520,N_18302,N_18277);
xor U18521 (N_18521,N_18359,N_18316);
or U18522 (N_18522,N_18246,N_18305);
and U18523 (N_18523,N_18388,N_18337);
xor U18524 (N_18524,N_18357,N_18364);
and U18525 (N_18525,N_18300,N_18356);
or U18526 (N_18526,N_18321,N_18282);
or U18527 (N_18527,N_18325,N_18276);
nand U18528 (N_18528,N_18370,N_18314);
and U18529 (N_18529,N_18313,N_18357);
nor U18530 (N_18530,N_18386,N_18273);
xnor U18531 (N_18531,N_18376,N_18266);
or U18532 (N_18532,N_18322,N_18376);
xnor U18533 (N_18533,N_18380,N_18260);
or U18534 (N_18534,N_18266,N_18370);
and U18535 (N_18535,N_18372,N_18393);
xor U18536 (N_18536,N_18255,N_18306);
nor U18537 (N_18537,N_18369,N_18270);
and U18538 (N_18538,N_18337,N_18364);
nand U18539 (N_18539,N_18339,N_18372);
xor U18540 (N_18540,N_18394,N_18314);
or U18541 (N_18541,N_18251,N_18343);
or U18542 (N_18542,N_18344,N_18337);
nand U18543 (N_18543,N_18310,N_18284);
xor U18544 (N_18544,N_18256,N_18268);
xnor U18545 (N_18545,N_18248,N_18274);
or U18546 (N_18546,N_18383,N_18308);
nand U18547 (N_18547,N_18306,N_18394);
xnor U18548 (N_18548,N_18339,N_18332);
nand U18549 (N_18549,N_18383,N_18352);
xnor U18550 (N_18550,N_18297,N_18374);
or U18551 (N_18551,N_18367,N_18350);
and U18552 (N_18552,N_18269,N_18329);
and U18553 (N_18553,N_18274,N_18297);
or U18554 (N_18554,N_18295,N_18354);
xor U18555 (N_18555,N_18313,N_18284);
or U18556 (N_18556,N_18392,N_18244);
nor U18557 (N_18557,N_18249,N_18295);
or U18558 (N_18558,N_18330,N_18305);
and U18559 (N_18559,N_18272,N_18288);
nor U18560 (N_18560,N_18470,N_18489);
nand U18561 (N_18561,N_18523,N_18528);
nor U18562 (N_18562,N_18538,N_18477);
or U18563 (N_18563,N_18441,N_18439);
or U18564 (N_18564,N_18433,N_18501);
and U18565 (N_18565,N_18488,N_18485);
xor U18566 (N_18566,N_18494,N_18497);
xnor U18567 (N_18567,N_18437,N_18541);
and U18568 (N_18568,N_18504,N_18490);
nand U18569 (N_18569,N_18510,N_18434);
xnor U18570 (N_18570,N_18557,N_18495);
nor U18571 (N_18571,N_18507,N_18440);
xor U18572 (N_18572,N_18429,N_18438);
or U18573 (N_18573,N_18473,N_18403);
or U18574 (N_18574,N_18533,N_18454);
or U18575 (N_18575,N_18539,N_18475);
or U18576 (N_18576,N_18401,N_18478);
nor U18577 (N_18577,N_18524,N_18500);
or U18578 (N_18578,N_18416,N_18453);
xnor U18579 (N_18579,N_18554,N_18515);
and U18580 (N_18580,N_18444,N_18460);
nor U18581 (N_18581,N_18514,N_18542);
nor U18582 (N_18582,N_18531,N_18499);
xor U18583 (N_18583,N_18445,N_18476);
or U18584 (N_18584,N_18550,N_18412);
and U18585 (N_18585,N_18417,N_18456);
nor U18586 (N_18586,N_18431,N_18421);
and U18587 (N_18587,N_18509,N_18442);
or U18588 (N_18588,N_18452,N_18492);
nor U18589 (N_18589,N_18424,N_18483);
nor U18590 (N_18590,N_18411,N_18435);
nand U18591 (N_18591,N_18540,N_18546);
or U18592 (N_18592,N_18423,N_18508);
nand U18593 (N_18593,N_18487,N_18462);
and U18594 (N_18594,N_18425,N_18448);
xor U18595 (N_18595,N_18518,N_18420);
xnor U18596 (N_18596,N_18543,N_18547);
xnor U18597 (N_18597,N_18409,N_18471);
and U18598 (N_18598,N_18517,N_18468);
or U18599 (N_18599,N_18455,N_18534);
nor U18600 (N_18600,N_18402,N_18548);
or U18601 (N_18601,N_18505,N_18472);
and U18602 (N_18602,N_18426,N_18479);
xnor U18603 (N_18603,N_18559,N_18449);
or U18604 (N_18604,N_18418,N_18530);
and U18605 (N_18605,N_18466,N_18450);
or U18606 (N_18606,N_18451,N_18527);
or U18607 (N_18607,N_18410,N_18529);
nor U18608 (N_18608,N_18436,N_18408);
nand U18609 (N_18609,N_18467,N_18464);
nor U18610 (N_18610,N_18427,N_18443);
nor U18611 (N_18611,N_18521,N_18558);
and U18612 (N_18612,N_18545,N_18463);
or U18613 (N_18613,N_18498,N_18465);
xnor U18614 (N_18614,N_18549,N_18512);
or U18615 (N_18615,N_18493,N_18491);
xnor U18616 (N_18616,N_18486,N_18496);
nor U18617 (N_18617,N_18461,N_18459);
nor U18618 (N_18618,N_18519,N_18481);
or U18619 (N_18619,N_18511,N_18474);
nor U18620 (N_18620,N_18406,N_18553);
nand U18621 (N_18621,N_18551,N_18535);
and U18622 (N_18622,N_18480,N_18526);
or U18623 (N_18623,N_18428,N_18482);
and U18624 (N_18624,N_18404,N_18484);
xor U18625 (N_18625,N_18419,N_18414);
and U18626 (N_18626,N_18555,N_18405);
and U18627 (N_18627,N_18469,N_18532);
and U18628 (N_18628,N_18544,N_18536);
xnor U18629 (N_18629,N_18525,N_18516);
xor U18630 (N_18630,N_18503,N_18446);
xnor U18631 (N_18631,N_18407,N_18502);
or U18632 (N_18632,N_18413,N_18457);
and U18633 (N_18633,N_18400,N_18556);
and U18634 (N_18634,N_18506,N_18432);
nand U18635 (N_18635,N_18422,N_18537);
xnor U18636 (N_18636,N_18552,N_18415);
or U18637 (N_18637,N_18513,N_18458);
nor U18638 (N_18638,N_18447,N_18430);
xor U18639 (N_18639,N_18522,N_18520);
and U18640 (N_18640,N_18515,N_18417);
nor U18641 (N_18641,N_18413,N_18533);
nor U18642 (N_18642,N_18421,N_18533);
and U18643 (N_18643,N_18530,N_18543);
nand U18644 (N_18644,N_18495,N_18531);
nor U18645 (N_18645,N_18521,N_18473);
nand U18646 (N_18646,N_18406,N_18504);
or U18647 (N_18647,N_18448,N_18526);
or U18648 (N_18648,N_18505,N_18401);
nand U18649 (N_18649,N_18409,N_18510);
nor U18650 (N_18650,N_18444,N_18512);
nand U18651 (N_18651,N_18511,N_18485);
xnor U18652 (N_18652,N_18527,N_18489);
or U18653 (N_18653,N_18554,N_18403);
and U18654 (N_18654,N_18539,N_18433);
nand U18655 (N_18655,N_18550,N_18466);
or U18656 (N_18656,N_18485,N_18522);
and U18657 (N_18657,N_18548,N_18430);
nor U18658 (N_18658,N_18415,N_18468);
or U18659 (N_18659,N_18465,N_18505);
or U18660 (N_18660,N_18459,N_18514);
or U18661 (N_18661,N_18489,N_18412);
nand U18662 (N_18662,N_18494,N_18477);
or U18663 (N_18663,N_18431,N_18487);
and U18664 (N_18664,N_18486,N_18407);
or U18665 (N_18665,N_18490,N_18495);
or U18666 (N_18666,N_18495,N_18461);
xnor U18667 (N_18667,N_18511,N_18410);
nand U18668 (N_18668,N_18412,N_18504);
xor U18669 (N_18669,N_18512,N_18487);
xor U18670 (N_18670,N_18525,N_18404);
or U18671 (N_18671,N_18444,N_18527);
nand U18672 (N_18672,N_18486,N_18453);
xor U18673 (N_18673,N_18461,N_18423);
nor U18674 (N_18674,N_18509,N_18517);
and U18675 (N_18675,N_18486,N_18467);
and U18676 (N_18676,N_18451,N_18484);
and U18677 (N_18677,N_18554,N_18492);
nor U18678 (N_18678,N_18516,N_18488);
xor U18679 (N_18679,N_18556,N_18456);
xnor U18680 (N_18680,N_18555,N_18410);
nor U18681 (N_18681,N_18429,N_18478);
and U18682 (N_18682,N_18413,N_18439);
or U18683 (N_18683,N_18546,N_18532);
or U18684 (N_18684,N_18429,N_18500);
xnor U18685 (N_18685,N_18476,N_18512);
and U18686 (N_18686,N_18438,N_18407);
nor U18687 (N_18687,N_18444,N_18435);
nor U18688 (N_18688,N_18476,N_18468);
and U18689 (N_18689,N_18516,N_18415);
xor U18690 (N_18690,N_18520,N_18488);
or U18691 (N_18691,N_18452,N_18541);
or U18692 (N_18692,N_18503,N_18510);
nor U18693 (N_18693,N_18544,N_18538);
nand U18694 (N_18694,N_18506,N_18467);
or U18695 (N_18695,N_18519,N_18538);
xnor U18696 (N_18696,N_18409,N_18435);
or U18697 (N_18697,N_18463,N_18544);
and U18698 (N_18698,N_18512,N_18480);
nand U18699 (N_18699,N_18465,N_18425);
and U18700 (N_18700,N_18488,N_18432);
and U18701 (N_18701,N_18518,N_18484);
nor U18702 (N_18702,N_18496,N_18514);
and U18703 (N_18703,N_18422,N_18445);
and U18704 (N_18704,N_18418,N_18479);
and U18705 (N_18705,N_18541,N_18522);
nand U18706 (N_18706,N_18408,N_18456);
nand U18707 (N_18707,N_18514,N_18472);
and U18708 (N_18708,N_18529,N_18419);
nor U18709 (N_18709,N_18526,N_18410);
nor U18710 (N_18710,N_18492,N_18481);
nand U18711 (N_18711,N_18545,N_18522);
nand U18712 (N_18712,N_18526,N_18433);
nor U18713 (N_18713,N_18496,N_18524);
nor U18714 (N_18714,N_18537,N_18559);
or U18715 (N_18715,N_18504,N_18539);
xor U18716 (N_18716,N_18547,N_18459);
xor U18717 (N_18717,N_18424,N_18480);
or U18718 (N_18718,N_18538,N_18556);
nand U18719 (N_18719,N_18426,N_18527);
nand U18720 (N_18720,N_18594,N_18568);
and U18721 (N_18721,N_18701,N_18580);
and U18722 (N_18722,N_18563,N_18607);
nand U18723 (N_18723,N_18581,N_18679);
xor U18724 (N_18724,N_18565,N_18641);
xnor U18725 (N_18725,N_18617,N_18691);
xor U18726 (N_18726,N_18570,N_18684);
nand U18727 (N_18727,N_18595,N_18714);
nor U18728 (N_18728,N_18653,N_18708);
and U18729 (N_18729,N_18562,N_18611);
and U18730 (N_18730,N_18694,N_18602);
and U18731 (N_18731,N_18640,N_18699);
or U18732 (N_18732,N_18589,N_18591);
and U18733 (N_18733,N_18672,N_18671);
or U18734 (N_18734,N_18600,N_18709);
or U18735 (N_18735,N_18670,N_18576);
and U18736 (N_18736,N_18673,N_18706);
xor U18737 (N_18737,N_18662,N_18643);
or U18738 (N_18738,N_18719,N_18637);
or U18739 (N_18739,N_18590,N_18695);
or U18740 (N_18740,N_18598,N_18690);
nand U18741 (N_18741,N_18642,N_18711);
or U18742 (N_18742,N_18698,N_18561);
xor U18743 (N_18743,N_18603,N_18681);
nand U18744 (N_18744,N_18664,N_18682);
xor U18745 (N_18745,N_18717,N_18638);
nor U18746 (N_18746,N_18592,N_18585);
and U18747 (N_18747,N_18588,N_18703);
and U18748 (N_18748,N_18618,N_18574);
nand U18749 (N_18749,N_18601,N_18639);
or U18750 (N_18750,N_18658,N_18577);
and U18751 (N_18751,N_18606,N_18668);
or U18752 (N_18752,N_18584,N_18700);
and U18753 (N_18753,N_18655,N_18648);
or U18754 (N_18754,N_18620,N_18605);
nand U18755 (N_18755,N_18612,N_18685);
nor U18756 (N_18756,N_18627,N_18630);
nand U18757 (N_18757,N_18621,N_18710);
nor U18758 (N_18758,N_18659,N_18582);
and U18759 (N_18759,N_18674,N_18656);
xnor U18760 (N_18760,N_18610,N_18686);
and U18761 (N_18761,N_18677,N_18564);
nand U18762 (N_18762,N_18716,N_18705);
nand U18763 (N_18763,N_18634,N_18624);
or U18764 (N_18764,N_18608,N_18599);
and U18765 (N_18765,N_18693,N_18687);
xor U18766 (N_18766,N_18586,N_18704);
nor U18767 (N_18767,N_18667,N_18718);
xor U18768 (N_18768,N_18609,N_18587);
or U18769 (N_18769,N_18613,N_18615);
xnor U18770 (N_18770,N_18678,N_18669);
xor U18771 (N_18771,N_18632,N_18622);
nand U18772 (N_18772,N_18660,N_18665);
or U18773 (N_18773,N_18571,N_18629);
and U18774 (N_18774,N_18579,N_18623);
nor U18775 (N_18775,N_18707,N_18635);
and U18776 (N_18776,N_18647,N_18631);
nand U18777 (N_18777,N_18619,N_18593);
or U18778 (N_18778,N_18689,N_18697);
and U18779 (N_18779,N_18616,N_18572);
xnor U18780 (N_18780,N_18676,N_18569);
xor U18781 (N_18781,N_18652,N_18597);
nor U18782 (N_18782,N_18628,N_18696);
xor U18783 (N_18783,N_18566,N_18567);
xor U18784 (N_18784,N_18650,N_18560);
xnor U18785 (N_18785,N_18666,N_18575);
or U18786 (N_18786,N_18649,N_18625);
xor U18787 (N_18787,N_18646,N_18680);
nor U18788 (N_18788,N_18654,N_18636);
or U18789 (N_18789,N_18578,N_18657);
xor U18790 (N_18790,N_18715,N_18626);
or U18791 (N_18791,N_18604,N_18675);
nor U18792 (N_18792,N_18663,N_18583);
xnor U18793 (N_18793,N_18692,N_18573);
nor U18794 (N_18794,N_18644,N_18712);
xnor U18795 (N_18795,N_18614,N_18651);
nor U18796 (N_18796,N_18596,N_18702);
nand U18797 (N_18797,N_18688,N_18661);
and U18798 (N_18798,N_18645,N_18633);
and U18799 (N_18799,N_18713,N_18683);
and U18800 (N_18800,N_18573,N_18628);
nand U18801 (N_18801,N_18586,N_18570);
nand U18802 (N_18802,N_18577,N_18709);
nor U18803 (N_18803,N_18696,N_18706);
or U18804 (N_18804,N_18693,N_18627);
and U18805 (N_18805,N_18617,N_18710);
xnor U18806 (N_18806,N_18714,N_18569);
xnor U18807 (N_18807,N_18610,N_18617);
xor U18808 (N_18808,N_18576,N_18671);
or U18809 (N_18809,N_18693,N_18588);
nand U18810 (N_18810,N_18575,N_18627);
xor U18811 (N_18811,N_18591,N_18635);
nand U18812 (N_18812,N_18630,N_18574);
nand U18813 (N_18813,N_18575,N_18617);
or U18814 (N_18814,N_18717,N_18579);
nor U18815 (N_18815,N_18657,N_18718);
nand U18816 (N_18816,N_18560,N_18674);
nand U18817 (N_18817,N_18714,N_18711);
xor U18818 (N_18818,N_18695,N_18645);
or U18819 (N_18819,N_18583,N_18600);
xnor U18820 (N_18820,N_18660,N_18704);
and U18821 (N_18821,N_18680,N_18694);
and U18822 (N_18822,N_18586,N_18648);
xnor U18823 (N_18823,N_18597,N_18636);
nor U18824 (N_18824,N_18689,N_18626);
nor U18825 (N_18825,N_18659,N_18644);
nand U18826 (N_18826,N_18637,N_18718);
and U18827 (N_18827,N_18649,N_18680);
nand U18828 (N_18828,N_18588,N_18653);
nor U18829 (N_18829,N_18660,N_18611);
or U18830 (N_18830,N_18592,N_18717);
nand U18831 (N_18831,N_18601,N_18590);
or U18832 (N_18832,N_18711,N_18654);
xor U18833 (N_18833,N_18639,N_18719);
nor U18834 (N_18834,N_18709,N_18630);
and U18835 (N_18835,N_18675,N_18656);
nor U18836 (N_18836,N_18626,N_18662);
or U18837 (N_18837,N_18658,N_18585);
nand U18838 (N_18838,N_18649,N_18619);
and U18839 (N_18839,N_18598,N_18648);
nor U18840 (N_18840,N_18644,N_18717);
and U18841 (N_18841,N_18707,N_18718);
nand U18842 (N_18842,N_18647,N_18607);
xor U18843 (N_18843,N_18710,N_18612);
nand U18844 (N_18844,N_18614,N_18650);
nand U18845 (N_18845,N_18655,N_18635);
nor U18846 (N_18846,N_18645,N_18607);
xnor U18847 (N_18847,N_18610,N_18654);
or U18848 (N_18848,N_18708,N_18642);
nor U18849 (N_18849,N_18580,N_18611);
or U18850 (N_18850,N_18649,N_18610);
nand U18851 (N_18851,N_18642,N_18702);
nor U18852 (N_18852,N_18686,N_18645);
nor U18853 (N_18853,N_18706,N_18715);
or U18854 (N_18854,N_18653,N_18649);
nor U18855 (N_18855,N_18703,N_18685);
nor U18856 (N_18856,N_18572,N_18682);
or U18857 (N_18857,N_18641,N_18648);
and U18858 (N_18858,N_18574,N_18605);
and U18859 (N_18859,N_18579,N_18675);
and U18860 (N_18860,N_18624,N_18662);
nand U18861 (N_18861,N_18579,N_18700);
xor U18862 (N_18862,N_18605,N_18656);
xor U18863 (N_18863,N_18634,N_18626);
nor U18864 (N_18864,N_18718,N_18681);
nor U18865 (N_18865,N_18590,N_18669);
nand U18866 (N_18866,N_18699,N_18584);
nand U18867 (N_18867,N_18671,N_18597);
nor U18868 (N_18868,N_18573,N_18587);
nor U18869 (N_18869,N_18688,N_18601);
or U18870 (N_18870,N_18660,N_18568);
nand U18871 (N_18871,N_18613,N_18609);
nor U18872 (N_18872,N_18618,N_18702);
nor U18873 (N_18873,N_18651,N_18650);
and U18874 (N_18874,N_18656,N_18672);
nor U18875 (N_18875,N_18714,N_18680);
nor U18876 (N_18876,N_18717,N_18686);
xor U18877 (N_18877,N_18610,N_18600);
or U18878 (N_18878,N_18712,N_18560);
nor U18879 (N_18879,N_18703,N_18568);
or U18880 (N_18880,N_18802,N_18877);
and U18881 (N_18881,N_18821,N_18723);
nor U18882 (N_18882,N_18825,N_18733);
xnor U18883 (N_18883,N_18753,N_18792);
or U18884 (N_18884,N_18824,N_18818);
or U18885 (N_18885,N_18801,N_18836);
xor U18886 (N_18886,N_18768,N_18831);
and U18887 (N_18887,N_18845,N_18868);
and U18888 (N_18888,N_18752,N_18800);
nor U18889 (N_18889,N_18826,N_18813);
nor U18890 (N_18890,N_18832,N_18812);
xor U18891 (N_18891,N_18780,N_18808);
nand U18892 (N_18892,N_18823,N_18748);
nor U18893 (N_18893,N_18811,N_18771);
or U18894 (N_18894,N_18851,N_18775);
nand U18895 (N_18895,N_18849,N_18765);
and U18896 (N_18896,N_18805,N_18777);
xor U18897 (N_18897,N_18767,N_18782);
xnor U18898 (N_18898,N_18844,N_18827);
and U18899 (N_18899,N_18721,N_18864);
nand U18900 (N_18900,N_18817,N_18720);
and U18901 (N_18901,N_18839,N_18734);
xnor U18902 (N_18902,N_18758,N_18854);
nand U18903 (N_18903,N_18822,N_18742);
nand U18904 (N_18904,N_18786,N_18769);
nor U18905 (N_18905,N_18772,N_18755);
nor U18906 (N_18906,N_18814,N_18749);
nand U18907 (N_18907,N_18750,N_18874);
nor U18908 (N_18908,N_18858,N_18779);
xor U18909 (N_18909,N_18746,N_18762);
xor U18910 (N_18910,N_18724,N_18837);
or U18911 (N_18911,N_18840,N_18737);
nand U18912 (N_18912,N_18797,N_18731);
or U18913 (N_18913,N_18867,N_18859);
and U18914 (N_18914,N_18773,N_18744);
and U18915 (N_18915,N_18842,N_18873);
nor U18916 (N_18916,N_18804,N_18725);
nand U18917 (N_18917,N_18745,N_18810);
or U18918 (N_18918,N_18846,N_18794);
nor U18919 (N_18919,N_18870,N_18757);
nor U18920 (N_18920,N_18829,N_18739);
nor U18921 (N_18921,N_18788,N_18820);
or U18922 (N_18922,N_18789,N_18860);
nand U18923 (N_18923,N_18751,N_18806);
nor U18924 (N_18924,N_18759,N_18754);
and U18925 (N_18925,N_18878,N_18774);
xor U18926 (N_18926,N_18766,N_18830);
and U18927 (N_18927,N_18848,N_18726);
and U18928 (N_18928,N_18722,N_18841);
xnor U18929 (N_18929,N_18778,N_18798);
or U18930 (N_18930,N_18876,N_18727);
nor U18931 (N_18931,N_18843,N_18736);
nand U18932 (N_18932,N_18847,N_18855);
and U18933 (N_18933,N_18764,N_18795);
xor U18934 (N_18934,N_18828,N_18863);
nor U18935 (N_18935,N_18781,N_18871);
nand U18936 (N_18936,N_18735,N_18791);
and U18937 (N_18937,N_18732,N_18793);
and U18938 (N_18938,N_18856,N_18747);
and U18939 (N_18939,N_18852,N_18834);
xor U18940 (N_18940,N_18815,N_18853);
and U18941 (N_18941,N_18783,N_18743);
nor U18942 (N_18942,N_18838,N_18879);
xnor U18943 (N_18943,N_18819,N_18799);
or U18944 (N_18944,N_18875,N_18763);
nand U18945 (N_18945,N_18807,N_18740);
or U18946 (N_18946,N_18861,N_18729);
or U18947 (N_18947,N_18761,N_18730);
xor U18948 (N_18948,N_18866,N_18803);
nor U18949 (N_18949,N_18741,N_18857);
xnor U18950 (N_18950,N_18738,N_18785);
nor U18951 (N_18951,N_18728,N_18865);
nor U18952 (N_18952,N_18796,N_18862);
nor U18953 (N_18953,N_18809,N_18787);
nand U18954 (N_18954,N_18756,N_18816);
nor U18955 (N_18955,N_18784,N_18872);
xor U18956 (N_18956,N_18790,N_18835);
nand U18957 (N_18957,N_18776,N_18850);
or U18958 (N_18958,N_18760,N_18770);
xor U18959 (N_18959,N_18869,N_18833);
nand U18960 (N_18960,N_18790,N_18829);
nand U18961 (N_18961,N_18771,N_18765);
xor U18962 (N_18962,N_18776,N_18841);
or U18963 (N_18963,N_18860,N_18802);
or U18964 (N_18964,N_18863,N_18822);
or U18965 (N_18965,N_18873,N_18812);
xor U18966 (N_18966,N_18869,N_18730);
nand U18967 (N_18967,N_18823,N_18865);
xor U18968 (N_18968,N_18850,N_18780);
xor U18969 (N_18969,N_18847,N_18879);
or U18970 (N_18970,N_18772,N_18846);
or U18971 (N_18971,N_18853,N_18735);
xor U18972 (N_18972,N_18804,N_18827);
nand U18973 (N_18973,N_18875,N_18830);
xnor U18974 (N_18974,N_18827,N_18766);
xnor U18975 (N_18975,N_18871,N_18799);
nand U18976 (N_18976,N_18747,N_18729);
xnor U18977 (N_18977,N_18803,N_18795);
xor U18978 (N_18978,N_18778,N_18786);
nor U18979 (N_18979,N_18782,N_18802);
nor U18980 (N_18980,N_18754,N_18732);
nand U18981 (N_18981,N_18740,N_18850);
and U18982 (N_18982,N_18794,N_18770);
xor U18983 (N_18983,N_18795,N_18734);
and U18984 (N_18984,N_18728,N_18856);
and U18985 (N_18985,N_18766,N_18805);
nor U18986 (N_18986,N_18748,N_18822);
or U18987 (N_18987,N_18859,N_18749);
and U18988 (N_18988,N_18816,N_18736);
and U18989 (N_18989,N_18852,N_18768);
nor U18990 (N_18990,N_18829,N_18830);
xor U18991 (N_18991,N_18816,N_18811);
xor U18992 (N_18992,N_18792,N_18860);
nand U18993 (N_18993,N_18824,N_18770);
xnor U18994 (N_18994,N_18862,N_18792);
nor U18995 (N_18995,N_18870,N_18722);
and U18996 (N_18996,N_18784,N_18773);
nor U18997 (N_18997,N_18869,N_18780);
nand U18998 (N_18998,N_18814,N_18727);
or U18999 (N_18999,N_18844,N_18741);
xnor U19000 (N_19000,N_18840,N_18870);
or U19001 (N_19001,N_18823,N_18818);
xnor U19002 (N_19002,N_18720,N_18768);
nand U19003 (N_19003,N_18772,N_18727);
and U19004 (N_19004,N_18878,N_18835);
xnor U19005 (N_19005,N_18785,N_18823);
and U19006 (N_19006,N_18727,N_18860);
nor U19007 (N_19007,N_18870,N_18877);
and U19008 (N_19008,N_18868,N_18770);
and U19009 (N_19009,N_18770,N_18802);
nor U19010 (N_19010,N_18823,N_18820);
xnor U19011 (N_19011,N_18753,N_18840);
nor U19012 (N_19012,N_18770,N_18720);
nor U19013 (N_19013,N_18804,N_18869);
nand U19014 (N_19014,N_18738,N_18848);
nor U19015 (N_19015,N_18731,N_18785);
or U19016 (N_19016,N_18786,N_18738);
or U19017 (N_19017,N_18838,N_18825);
nor U19018 (N_19018,N_18803,N_18837);
nor U19019 (N_19019,N_18740,N_18865);
or U19020 (N_19020,N_18743,N_18856);
and U19021 (N_19021,N_18804,N_18816);
nand U19022 (N_19022,N_18834,N_18870);
and U19023 (N_19023,N_18818,N_18852);
xor U19024 (N_19024,N_18764,N_18807);
nand U19025 (N_19025,N_18731,N_18800);
and U19026 (N_19026,N_18821,N_18771);
nand U19027 (N_19027,N_18759,N_18767);
xor U19028 (N_19028,N_18788,N_18787);
nor U19029 (N_19029,N_18769,N_18820);
nand U19030 (N_19030,N_18812,N_18782);
nand U19031 (N_19031,N_18820,N_18774);
and U19032 (N_19032,N_18807,N_18842);
nand U19033 (N_19033,N_18771,N_18798);
xor U19034 (N_19034,N_18770,N_18787);
or U19035 (N_19035,N_18791,N_18856);
or U19036 (N_19036,N_18753,N_18816);
nor U19037 (N_19037,N_18732,N_18765);
nor U19038 (N_19038,N_18850,N_18802);
nor U19039 (N_19039,N_18807,N_18851);
xor U19040 (N_19040,N_18902,N_18988);
nand U19041 (N_19041,N_18893,N_19004);
xnor U19042 (N_19042,N_18930,N_19015);
nand U19043 (N_19043,N_18979,N_18960);
nand U19044 (N_19044,N_18994,N_18915);
and U19045 (N_19045,N_18973,N_19024);
or U19046 (N_19046,N_18952,N_18895);
nor U19047 (N_19047,N_18948,N_18937);
xnor U19048 (N_19048,N_19032,N_19020);
or U19049 (N_19049,N_18949,N_18891);
nor U19050 (N_19050,N_18968,N_18995);
nand U19051 (N_19051,N_18955,N_18999);
nand U19052 (N_19052,N_18890,N_18982);
or U19053 (N_19053,N_18980,N_19027);
and U19054 (N_19054,N_18958,N_18925);
nand U19055 (N_19055,N_18996,N_18887);
and U19056 (N_19056,N_18900,N_18899);
nor U19057 (N_19057,N_18991,N_18967);
or U19058 (N_19058,N_18880,N_19038);
xnor U19059 (N_19059,N_19022,N_18903);
or U19060 (N_19060,N_18928,N_18997);
xor U19061 (N_19061,N_18938,N_18916);
nand U19062 (N_19062,N_18907,N_19007);
or U19063 (N_19063,N_18953,N_18918);
and U19064 (N_19064,N_18888,N_18978);
or U19065 (N_19065,N_18909,N_19030);
nand U19066 (N_19066,N_18964,N_18970);
xnor U19067 (N_19067,N_18933,N_18976);
and U19068 (N_19068,N_18942,N_18983);
nand U19069 (N_19069,N_18946,N_18917);
and U19070 (N_19070,N_18969,N_18965);
or U19071 (N_19071,N_18950,N_19031);
and U19072 (N_19072,N_18919,N_18898);
nor U19073 (N_19073,N_18984,N_18981);
nand U19074 (N_19074,N_19039,N_18956);
or U19075 (N_19075,N_18911,N_18989);
and U19076 (N_19076,N_18894,N_19016);
xor U19077 (N_19077,N_18886,N_18954);
or U19078 (N_19078,N_18924,N_19014);
xor U19079 (N_19079,N_18987,N_18951);
or U19080 (N_19080,N_18962,N_18943);
xnor U19081 (N_19081,N_18905,N_18974);
or U19082 (N_19082,N_18977,N_18910);
nand U19083 (N_19083,N_18939,N_18944);
xnor U19084 (N_19084,N_18945,N_19028);
and U19085 (N_19085,N_18882,N_18957);
or U19086 (N_19086,N_19001,N_18998);
nand U19087 (N_19087,N_18885,N_19026);
nand U19088 (N_19088,N_18993,N_18961);
xnor U19089 (N_19089,N_19012,N_18883);
xor U19090 (N_19090,N_18947,N_19023);
xnor U19091 (N_19091,N_19000,N_19036);
nand U19092 (N_19092,N_18927,N_18941);
and U19093 (N_19093,N_19034,N_19018);
and U19094 (N_19094,N_18908,N_18921);
and U19095 (N_19095,N_18912,N_19029);
or U19096 (N_19096,N_18931,N_18922);
or U19097 (N_19097,N_19009,N_18990);
xor U19098 (N_19098,N_18940,N_19011);
and U19099 (N_19099,N_18901,N_18906);
and U19100 (N_19100,N_19037,N_18985);
nand U19101 (N_19101,N_19013,N_19019);
nor U19102 (N_19102,N_19010,N_18936);
nor U19103 (N_19103,N_19008,N_18966);
xnor U19104 (N_19104,N_18923,N_19017);
xnor U19105 (N_19105,N_19025,N_18881);
or U19106 (N_19106,N_18929,N_19035);
xnor U19107 (N_19107,N_19003,N_18932);
nor U19108 (N_19108,N_18992,N_18892);
nor U19109 (N_19109,N_18884,N_18904);
or U19110 (N_19110,N_18934,N_18975);
xnor U19111 (N_19111,N_18896,N_18959);
xnor U19112 (N_19112,N_19006,N_18926);
nand U19113 (N_19113,N_18914,N_18920);
nor U19114 (N_19114,N_18935,N_19033);
nand U19115 (N_19115,N_18889,N_18971);
xnor U19116 (N_19116,N_19021,N_18963);
nor U19117 (N_19117,N_18972,N_18913);
nor U19118 (N_19118,N_19002,N_18986);
nor U19119 (N_19119,N_19005,N_18897);
nand U19120 (N_19120,N_19012,N_18880);
or U19121 (N_19121,N_18903,N_19019);
or U19122 (N_19122,N_19006,N_18886);
nand U19123 (N_19123,N_18992,N_19015);
nor U19124 (N_19124,N_18928,N_18927);
nor U19125 (N_19125,N_18923,N_18942);
nor U19126 (N_19126,N_19017,N_18973);
nand U19127 (N_19127,N_18951,N_18916);
nand U19128 (N_19128,N_18986,N_18922);
or U19129 (N_19129,N_18950,N_18966);
or U19130 (N_19130,N_18930,N_18972);
xnor U19131 (N_19131,N_19031,N_18920);
or U19132 (N_19132,N_19026,N_19027);
nor U19133 (N_19133,N_18935,N_18884);
and U19134 (N_19134,N_18966,N_19022);
and U19135 (N_19135,N_18991,N_18997);
nor U19136 (N_19136,N_19024,N_18892);
nor U19137 (N_19137,N_18913,N_19028);
nand U19138 (N_19138,N_18997,N_18996);
nand U19139 (N_19139,N_18942,N_18995);
nand U19140 (N_19140,N_18936,N_18991);
nand U19141 (N_19141,N_18883,N_19015);
xnor U19142 (N_19142,N_18934,N_18962);
nor U19143 (N_19143,N_18904,N_18936);
xnor U19144 (N_19144,N_18958,N_18940);
or U19145 (N_19145,N_18894,N_19024);
or U19146 (N_19146,N_19016,N_18970);
xnor U19147 (N_19147,N_18896,N_18997);
nand U19148 (N_19148,N_18991,N_19039);
and U19149 (N_19149,N_18914,N_18966);
nor U19150 (N_19150,N_18926,N_18945);
and U19151 (N_19151,N_18891,N_18919);
nor U19152 (N_19152,N_18957,N_18913);
nor U19153 (N_19153,N_18918,N_18922);
nor U19154 (N_19154,N_18938,N_18888);
or U19155 (N_19155,N_18896,N_19037);
xnor U19156 (N_19156,N_18923,N_18881);
xor U19157 (N_19157,N_18943,N_18955);
and U19158 (N_19158,N_18946,N_18969);
xor U19159 (N_19159,N_19023,N_18935);
nor U19160 (N_19160,N_19034,N_18932);
and U19161 (N_19161,N_18944,N_18927);
nand U19162 (N_19162,N_18976,N_19020);
or U19163 (N_19163,N_18934,N_18982);
xor U19164 (N_19164,N_18931,N_19012);
nor U19165 (N_19165,N_18978,N_18936);
nand U19166 (N_19166,N_19036,N_18965);
and U19167 (N_19167,N_18892,N_19037);
nor U19168 (N_19168,N_18975,N_18903);
or U19169 (N_19169,N_18971,N_18945);
and U19170 (N_19170,N_18954,N_19033);
or U19171 (N_19171,N_18959,N_18991);
xor U19172 (N_19172,N_19034,N_18988);
nand U19173 (N_19173,N_19026,N_18946);
xnor U19174 (N_19174,N_18890,N_18948);
nor U19175 (N_19175,N_18941,N_19023);
nor U19176 (N_19176,N_19022,N_18963);
or U19177 (N_19177,N_19002,N_18891);
nand U19178 (N_19178,N_18980,N_18983);
xnor U19179 (N_19179,N_18980,N_18909);
nor U19180 (N_19180,N_18929,N_18892);
nand U19181 (N_19181,N_18939,N_18994);
nor U19182 (N_19182,N_18888,N_18924);
and U19183 (N_19183,N_19010,N_19017);
and U19184 (N_19184,N_19018,N_18891);
nand U19185 (N_19185,N_19038,N_18914);
and U19186 (N_19186,N_19000,N_18928);
xnor U19187 (N_19187,N_18929,N_19036);
nor U19188 (N_19188,N_19010,N_18881);
and U19189 (N_19189,N_18997,N_18917);
and U19190 (N_19190,N_19009,N_18892);
nand U19191 (N_19191,N_18995,N_19002);
or U19192 (N_19192,N_18896,N_18880);
nand U19193 (N_19193,N_18903,N_19030);
nand U19194 (N_19194,N_19000,N_19018);
and U19195 (N_19195,N_18983,N_18991);
xnor U19196 (N_19196,N_18981,N_18926);
and U19197 (N_19197,N_19031,N_18946);
or U19198 (N_19198,N_19003,N_18900);
xnor U19199 (N_19199,N_18990,N_19035);
nor U19200 (N_19200,N_19109,N_19108);
and U19201 (N_19201,N_19061,N_19173);
nand U19202 (N_19202,N_19127,N_19110);
or U19203 (N_19203,N_19074,N_19174);
and U19204 (N_19204,N_19097,N_19129);
xnor U19205 (N_19205,N_19182,N_19133);
nand U19206 (N_19206,N_19075,N_19164);
and U19207 (N_19207,N_19181,N_19073);
nor U19208 (N_19208,N_19086,N_19193);
xnor U19209 (N_19209,N_19145,N_19103);
xnor U19210 (N_19210,N_19112,N_19066);
nor U19211 (N_19211,N_19043,N_19091);
xnor U19212 (N_19212,N_19094,N_19084);
and U19213 (N_19213,N_19069,N_19160);
nand U19214 (N_19214,N_19158,N_19166);
xor U19215 (N_19215,N_19134,N_19096);
nand U19216 (N_19216,N_19046,N_19065);
nor U19217 (N_19217,N_19198,N_19183);
or U19218 (N_19218,N_19057,N_19076);
xnor U19219 (N_19219,N_19100,N_19104);
nor U19220 (N_19220,N_19184,N_19197);
xor U19221 (N_19221,N_19063,N_19171);
or U19222 (N_19222,N_19105,N_19044);
or U19223 (N_19223,N_19176,N_19187);
nor U19224 (N_19224,N_19153,N_19189);
nand U19225 (N_19225,N_19170,N_19142);
xnor U19226 (N_19226,N_19150,N_19119);
nor U19227 (N_19227,N_19120,N_19149);
nand U19228 (N_19228,N_19169,N_19121);
or U19229 (N_19229,N_19147,N_19122);
nor U19230 (N_19230,N_19054,N_19102);
xor U19231 (N_19231,N_19048,N_19131);
and U19232 (N_19232,N_19196,N_19154);
or U19233 (N_19233,N_19128,N_19168);
nand U19234 (N_19234,N_19049,N_19050);
nand U19235 (N_19235,N_19042,N_19088);
nor U19236 (N_19236,N_19070,N_19126);
nand U19237 (N_19237,N_19143,N_19056);
or U19238 (N_19238,N_19125,N_19079);
or U19239 (N_19239,N_19047,N_19045);
nand U19240 (N_19240,N_19188,N_19064);
or U19241 (N_19241,N_19067,N_19194);
nand U19242 (N_19242,N_19082,N_19078);
or U19243 (N_19243,N_19137,N_19068);
or U19244 (N_19244,N_19152,N_19186);
nand U19245 (N_19245,N_19124,N_19148);
xnor U19246 (N_19246,N_19113,N_19099);
xnor U19247 (N_19247,N_19191,N_19077);
nand U19248 (N_19248,N_19146,N_19195);
xor U19249 (N_19249,N_19060,N_19136);
xnor U19250 (N_19250,N_19175,N_19178);
nand U19251 (N_19251,N_19157,N_19165);
or U19252 (N_19252,N_19055,N_19138);
or U19253 (N_19253,N_19114,N_19163);
and U19254 (N_19254,N_19072,N_19144);
and U19255 (N_19255,N_19141,N_19058);
or U19256 (N_19256,N_19117,N_19130);
xnor U19257 (N_19257,N_19095,N_19085);
and U19258 (N_19258,N_19107,N_19090);
or U19259 (N_19259,N_19052,N_19083);
nor U19260 (N_19260,N_19159,N_19111);
and U19261 (N_19261,N_19081,N_19185);
nand U19262 (N_19262,N_19087,N_19155);
nor U19263 (N_19263,N_19089,N_19162);
nand U19264 (N_19264,N_19115,N_19190);
or U19265 (N_19265,N_19041,N_19139);
nand U19266 (N_19266,N_19172,N_19080);
nand U19267 (N_19267,N_19161,N_19151);
nand U19268 (N_19268,N_19116,N_19040);
nor U19269 (N_19269,N_19062,N_19192);
and U19270 (N_19270,N_19180,N_19071);
or U19271 (N_19271,N_19118,N_19132);
or U19272 (N_19272,N_19135,N_19177);
nor U19273 (N_19273,N_19101,N_19098);
or U19274 (N_19274,N_19093,N_19156);
xor U19275 (N_19275,N_19167,N_19179);
nand U19276 (N_19276,N_19106,N_19092);
or U19277 (N_19277,N_19053,N_19140);
xnor U19278 (N_19278,N_19051,N_19123);
nor U19279 (N_19279,N_19199,N_19059);
nand U19280 (N_19280,N_19054,N_19071);
and U19281 (N_19281,N_19060,N_19175);
or U19282 (N_19282,N_19151,N_19180);
or U19283 (N_19283,N_19068,N_19172);
nor U19284 (N_19284,N_19097,N_19136);
xor U19285 (N_19285,N_19068,N_19107);
nor U19286 (N_19286,N_19080,N_19110);
nor U19287 (N_19287,N_19199,N_19190);
nor U19288 (N_19288,N_19146,N_19182);
nor U19289 (N_19289,N_19061,N_19136);
and U19290 (N_19290,N_19132,N_19094);
and U19291 (N_19291,N_19130,N_19161);
and U19292 (N_19292,N_19128,N_19196);
xnor U19293 (N_19293,N_19175,N_19074);
nand U19294 (N_19294,N_19138,N_19157);
or U19295 (N_19295,N_19047,N_19146);
nand U19296 (N_19296,N_19177,N_19078);
nor U19297 (N_19297,N_19113,N_19152);
and U19298 (N_19298,N_19126,N_19091);
and U19299 (N_19299,N_19182,N_19063);
nand U19300 (N_19300,N_19043,N_19101);
nand U19301 (N_19301,N_19089,N_19123);
or U19302 (N_19302,N_19117,N_19182);
and U19303 (N_19303,N_19170,N_19041);
nand U19304 (N_19304,N_19144,N_19097);
or U19305 (N_19305,N_19106,N_19172);
or U19306 (N_19306,N_19155,N_19093);
nand U19307 (N_19307,N_19186,N_19139);
nand U19308 (N_19308,N_19048,N_19182);
and U19309 (N_19309,N_19117,N_19055);
and U19310 (N_19310,N_19042,N_19094);
nand U19311 (N_19311,N_19056,N_19057);
nand U19312 (N_19312,N_19183,N_19042);
and U19313 (N_19313,N_19045,N_19098);
and U19314 (N_19314,N_19156,N_19176);
or U19315 (N_19315,N_19080,N_19064);
nand U19316 (N_19316,N_19146,N_19138);
xnor U19317 (N_19317,N_19112,N_19152);
nor U19318 (N_19318,N_19058,N_19195);
and U19319 (N_19319,N_19120,N_19154);
nor U19320 (N_19320,N_19058,N_19118);
xor U19321 (N_19321,N_19102,N_19046);
and U19322 (N_19322,N_19112,N_19197);
and U19323 (N_19323,N_19148,N_19145);
and U19324 (N_19324,N_19064,N_19147);
or U19325 (N_19325,N_19173,N_19048);
nor U19326 (N_19326,N_19138,N_19151);
or U19327 (N_19327,N_19134,N_19165);
nor U19328 (N_19328,N_19056,N_19111);
nand U19329 (N_19329,N_19125,N_19056);
xnor U19330 (N_19330,N_19104,N_19189);
xor U19331 (N_19331,N_19118,N_19065);
xor U19332 (N_19332,N_19161,N_19148);
or U19333 (N_19333,N_19061,N_19163);
xnor U19334 (N_19334,N_19118,N_19114);
and U19335 (N_19335,N_19158,N_19048);
nand U19336 (N_19336,N_19153,N_19165);
xnor U19337 (N_19337,N_19146,N_19165);
or U19338 (N_19338,N_19079,N_19159);
or U19339 (N_19339,N_19175,N_19048);
nor U19340 (N_19340,N_19059,N_19089);
and U19341 (N_19341,N_19097,N_19040);
nand U19342 (N_19342,N_19189,N_19083);
nand U19343 (N_19343,N_19105,N_19137);
or U19344 (N_19344,N_19185,N_19066);
and U19345 (N_19345,N_19080,N_19117);
xor U19346 (N_19346,N_19118,N_19052);
and U19347 (N_19347,N_19079,N_19083);
and U19348 (N_19348,N_19099,N_19105);
xor U19349 (N_19349,N_19106,N_19087);
and U19350 (N_19350,N_19135,N_19115);
xor U19351 (N_19351,N_19055,N_19073);
xor U19352 (N_19352,N_19089,N_19192);
or U19353 (N_19353,N_19166,N_19048);
xnor U19354 (N_19354,N_19052,N_19070);
nand U19355 (N_19355,N_19099,N_19119);
and U19356 (N_19356,N_19114,N_19055);
or U19357 (N_19357,N_19041,N_19164);
nand U19358 (N_19358,N_19190,N_19092);
or U19359 (N_19359,N_19170,N_19191);
xor U19360 (N_19360,N_19299,N_19305);
xnor U19361 (N_19361,N_19226,N_19341);
xor U19362 (N_19362,N_19265,N_19204);
nand U19363 (N_19363,N_19202,N_19334);
nand U19364 (N_19364,N_19230,N_19242);
xnor U19365 (N_19365,N_19355,N_19319);
nor U19366 (N_19366,N_19336,N_19237);
and U19367 (N_19367,N_19288,N_19253);
and U19368 (N_19368,N_19248,N_19201);
nand U19369 (N_19369,N_19238,N_19272);
nor U19370 (N_19370,N_19313,N_19358);
and U19371 (N_19371,N_19261,N_19303);
and U19372 (N_19372,N_19219,N_19295);
or U19373 (N_19373,N_19267,N_19290);
nand U19374 (N_19374,N_19325,N_19220);
and U19375 (N_19375,N_19284,N_19281);
or U19376 (N_19376,N_19221,N_19274);
xnor U19377 (N_19377,N_19335,N_19214);
xnor U19378 (N_19378,N_19245,N_19251);
nand U19379 (N_19379,N_19208,N_19206);
nor U19380 (N_19380,N_19329,N_19279);
xnor U19381 (N_19381,N_19207,N_19282);
or U19382 (N_19382,N_19345,N_19225);
nand U19383 (N_19383,N_19353,N_19337);
and U19384 (N_19384,N_19234,N_19339);
nor U19385 (N_19385,N_19217,N_19269);
xnor U19386 (N_19386,N_19314,N_19354);
or U19387 (N_19387,N_19239,N_19293);
nand U19388 (N_19388,N_19338,N_19203);
nor U19389 (N_19389,N_19210,N_19250);
nand U19390 (N_19390,N_19256,N_19323);
nor U19391 (N_19391,N_19236,N_19312);
xnor U19392 (N_19392,N_19351,N_19356);
nor U19393 (N_19393,N_19324,N_19277);
and U19394 (N_19394,N_19212,N_19233);
nor U19395 (N_19395,N_19231,N_19307);
and U19396 (N_19396,N_19211,N_19322);
and U19397 (N_19397,N_19289,N_19241);
nand U19398 (N_19398,N_19342,N_19318);
xor U19399 (N_19399,N_19321,N_19213);
and U19400 (N_19400,N_19227,N_19301);
nand U19401 (N_19401,N_19232,N_19235);
and U19402 (N_19402,N_19352,N_19331);
or U19403 (N_19403,N_19209,N_19332);
xor U19404 (N_19404,N_19263,N_19287);
or U19405 (N_19405,N_19258,N_19268);
nand U19406 (N_19406,N_19346,N_19270);
xor U19407 (N_19407,N_19278,N_19283);
or U19408 (N_19408,N_19264,N_19326);
nor U19409 (N_19409,N_19349,N_19247);
xor U19410 (N_19410,N_19273,N_19229);
nor U19411 (N_19411,N_19259,N_19266);
and U19412 (N_19412,N_19347,N_19298);
xnor U19413 (N_19413,N_19275,N_19306);
or U19414 (N_19414,N_19308,N_19333);
nand U19415 (N_19415,N_19271,N_19340);
and U19416 (N_19416,N_19317,N_19276);
or U19417 (N_19417,N_19257,N_19228);
xor U19418 (N_19418,N_19244,N_19240);
and U19419 (N_19419,N_19254,N_19200);
or U19420 (N_19420,N_19311,N_19330);
and U19421 (N_19421,N_19310,N_19205);
xnor U19422 (N_19422,N_19222,N_19218);
xor U19423 (N_19423,N_19302,N_19294);
nor U19424 (N_19424,N_19343,N_19291);
nand U19425 (N_19425,N_19320,N_19350);
nand U19426 (N_19426,N_19285,N_19359);
or U19427 (N_19427,N_19255,N_19260);
nand U19428 (N_19428,N_19292,N_19280);
xnor U19429 (N_19429,N_19249,N_19224);
nand U19430 (N_19430,N_19300,N_19315);
and U19431 (N_19431,N_19286,N_19223);
nor U19432 (N_19432,N_19243,N_19262);
nor U19433 (N_19433,N_19328,N_19246);
xor U19434 (N_19434,N_19309,N_19316);
or U19435 (N_19435,N_19216,N_19348);
or U19436 (N_19436,N_19304,N_19357);
nor U19437 (N_19437,N_19344,N_19297);
and U19438 (N_19438,N_19296,N_19327);
xnor U19439 (N_19439,N_19215,N_19252);
and U19440 (N_19440,N_19248,N_19322);
and U19441 (N_19441,N_19322,N_19295);
xor U19442 (N_19442,N_19304,N_19231);
xor U19443 (N_19443,N_19259,N_19267);
nand U19444 (N_19444,N_19291,N_19270);
xor U19445 (N_19445,N_19220,N_19251);
or U19446 (N_19446,N_19321,N_19259);
nor U19447 (N_19447,N_19262,N_19350);
or U19448 (N_19448,N_19331,N_19274);
or U19449 (N_19449,N_19314,N_19253);
nor U19450 (N_19450,N_19249,N_19329);
xor U19451 (N_19451,N_19284,N_19298);
xnor U19452 (N_19452,N_19204,N_19317);
nor U19453 (N_19453,N_19239,N_19209);
nand U19454 (N_19454,N_19358,N_19300);
and U19455 (N_19455,N_19271,N_19259);
nand U19456 (N_19456,N_19263,N_19227);
nor U19457 (N_19457,N_19315,N_19344);
or U19458 (N_19458,N_19249,N_19256);
xor U19459 (N_19459,N_19282,N_19310);
xnor U19460 (N_19460,N_19290,N_19256);
or U19461 (N_19461,N_19271,N_19242);
or U19462 (N_19462,N_19352,N_19334);
nor U19463 (N_19463,N_19311,N_19278);
or U19464 (N_19464,N_19246,N_19215);
or U19465 (N_19465,N_19308,N_19254);
nand U19466 (N_19466,N_19341,N_19253);
nand U19467 (N_19467,N_19275,N_19245);
and U19468 (N_19468,N_19351,N_19286);
and U19469 (N_19469,N_19226,N_19329);
nand U19470 (N_19470,N_19299,N_19237);
or U19471 (N_19471,N_19206,N_19235);
or U19472 (N_19472,N_19263,N_19348);
xnor U19473 (N_19473,N_19322,N_19317);
and U19474 (N_19474,N_19311,N_19249);
nor U19475 (N_19475,N_19263,N_19299);
and U19476 (N_19476,N_19310,N_19351);
nor U19477 (N_19477,N_19215,N_19207);
nand U19478 (N_19478,N_19278,N_19242);
nor U19479 (N_19479,N_19311,N_19235);
or U19480 (N_19480,N_19258,N_19216);
nand U19481 (N_19481,N_19200,N_19333);
and U19482 (N_19482,N_19319,N_19295);
and U19483 (N_19483,N_19270,N_19238);
nand U19484 (N_19484,N_19239,N_19228);
and U19485 (N_19485,N_19255,N_19352);
and U19486 (N_19486,N_19317,N_19251);
nor U19487 (N_19487,N_19293,N_19201);
or U19488 (N_19488,N_19271,N_19277);
or U19489 (N_19489,N_19251,N_19272);
and U19490 (N_19490,N_19289,N_19330);
nor U19491 (N_19491,N_19317,N_19353);
xnor U19492 (N_19492,N_19205,N_19236);
and U19493 (N_19493,N_19287,N_19290);
or U19494 (N_19494,N_19278,N_19325);
xnor U19495 (N_19495,N_19303,N_19357);
or U19496 (N_19496,N_19279,N_19247);
and U19497 (N_19497,N_19291,N_19205);
nor U19498 (N_19498,N_19222,N_19283);
xor U19499 (N_19499,N_19255,N_19345);
and U19500 (N_19500,N_19291,N_19315);
nor U19501 (N_19501,N_19256,N_19339);
or U19502 (N_19502,N_19330,N_19280);
and U19503 (N_19503,N_19267,N_19221);
nor U19504 (N_19504,N_19331,N_19304);
xor U19505 (N_19505,N_19205,N_19235);
or U19506 (N_19506,N_19282,N_19336);
and U19507 (N_19507,N_19308,N_19352);
or U19508 (N_19508,N_19318,N_19279);
or U19509 (N_19509,N_19303,N_19283);
and U19510 (N_19510,N_19307,N_19347);
nor U19511 (N_19511,N_19284,N_19271);
nand U19512 (N_19512,N_19263,N_19261);
or U19513 (N_19513,N_19234,N_19300);
nor U19514 (N_19514,N_19207,N_19329);
nand U19515 (N_19515,N_19234,N_19219);
or U19516 (N_19516,N_19293,N_19332);
nor U19517 (N_19517,N_19291,N_19241);
nand U19518 (N_19518,N_19334,N_19314);
or U19519 (N_19519,N_19312,N_19255);
nand U19520 (N_19520,N_19517,N_19466);
xor U19521 (N_19521,N_19450,N_19360);
or U19522 (N_19522,N_19459,N_19444);
and U19523 (N_19523,N_19372,N_19514);
nor U19524 (N_19524,N_19430,N_19382);
and U19525 (N_19525,N_19417,N_19453);
or U19526 (N_19526,N_19463,N_19509);
xnor U19527 (N_19527,N_19394,N_19428);
or U19528 (N_19528,N_19454,N_19474);
nor U19529 (N_19529,N_19398,N_19456);
and U19530 (N_19530,N_19468,N_19470);
and U19531 (N_19531,N_19407,N_19479);
and U19532 (N_19532,N_19461,N_19501);
xor U19533 (N_19533,N_19410,N_19441);
nand U19534 (N_19534,N_19368,N_19469);
nor U19535 (N_19535,N_19375,N_19413);
nor U19536 (N_19536,N_19381,N_19478);
xnor U19537 (N_19537,N_19485,N_19452);
nand U19538 (N_19538,N_19486,N_19516);
xnor U19539 (N_19539,N_19405,N_19435);
xnor U19540 (N_19540,N_19391,N_19481);
or U19541 (N_19541,N_19439,N_19383);
or U19542 (N_19542,N_19484,N_19483);
nand U19543 (N_19543,N_19401,N_19473);
xnor U19544 (N_19544,N_19499,N_19460);
nor U19545 (N_19545,N_19457,N_19403);
and U19546 (N_19546,N_19385,N_19414);
nand U19547 (N_19547,N_19366,N_19511);
xnor U19548 (N_19548,N_19489,N_19418);
or U19549 (N_19549,N_19502,N_19379);
or U19550 (N_19550,N_19458,N_19507);
nand U19551 (N_19551,N_19378,N_19377);
nand U19552 (N_19552,N_19415,N_19402);
xnor U19553 (N_19553,N_19429,N_19362);
and U19554 (N_19554,N_19437,N_19373);
xnor U19555 (N_19555,N_19471,N_19467);
nand U19556 (N_19556,N_19393,N_19445);
nand U19557 (N_19557,N_19455,N_19475);
xor U19558 (N_19558,N_19423,N_19397);
or U19559 (N_19559,N_19361,N_19506);
and U19560 (N_19560,N_19493,N_19464);
nand U19561 (N_19561,N_19426,N_19477);
or U19562 (N_19562,N_19436,N_19370);
or U19563 (N_19563,N_19438,N_19496);
nand U19564 (N_19564,N_19490,N_19404);
xnor U19565 (N_19565,N_19421,N_19386);
nand U19566 (N_19566,N_19498,N_19446);
nor U19567 (N_19567,N_19491,N_19390);
xnor U19568 (N_19568,N_19519,N_19431);
and U19569 (N_19569,N_19364,N_19447);
nand U19570 (N_19570,N_19400,N_19424);
and U19571 (N_19571,N_19395,N_19416);
xnor U19572 (N_19572,N_19462,N_19449);
and U19573 (N_19573,N_19465,N_19488);
and U19574 (N_19574,N_19451,N_19505);
nor U19575 (N_19575,N_19518,N_19419);
nand U19576 (N_19576,N_19497,N_19433);
nor U19577 (N_19577,N_19411,N_19406);
nand U19578 (N_19578,N_19380,N_19442);
nand U19579 (N_19579,N_19503,N_19367);
xnor U19580 (N_19580,N_19384,N_19472);
nor U19581 (N_19581,N_19494,N_19369);
nor U19582 (N_19582,N_19508,N_19389);
xnor U19583 (N_19583,N_19392,N_19448);
or U19584 (N_19584,N_19440,N_19512);
or U19585 (N_19585,N_19482,N_19387);
nand U19586 (N_19586,N_19374,N_19408);
nor U19587 (N_19587,N_19432,N_19420);
or U19588 (N_19588,N_19480,N_19427);
nor U19589 (N_19589,N_19396,N_19365);
or U19590 (N_19590,N_19422,N_19376);
nor U19591 (N_19591,N_19409,N_19510);
nand U19592 (N_19592,N_19492,N_19388);
nor U19593 (N_19593,N_19434,N_19515);
and U19594 (N_19594,N_19425,N_19476);
or U19595 (N_19595,N_19363,N_19371);
and U19596 (N_19596,N_19500,N_19443);
nor U19597 (N_19597,N_19412,N_19487);
or U19598 (N_19598,N_19399,N_19495);
and U19599 (N_19599,N_19513,N_19504);
and U19600 (N_19600,N_19459,N_19458);
xnor U19601 (N_19601,N_19432,N_19477);
or U19602 (N_19602,N_19441,N_19427);
or U19603 (N_19603,N_19478,N_19405);
xor U19604 (N_19604,N_19476,N_19460);
and U19605 (N_19605,N_19381,N_19387);
xnor U19606 (N_19606,N_19408,N_19388);
nand U19607 (N_19607,N_19377,N_19375);
nor U19608 (N_19608,N_19511,N_19484);
xor U19609 (N_19609,N_19488,N_19454);
nand U19610 (N_19610,N_19490,N_19485);
nor U19611 (N_19611,N_19469,N_19422);
or U19612 (N_19612,N_19489,N_19401);
nor U19613 (N_19613,N_19415,N_19502);
nor U19614 (N_19614,N_19432,N_19413);
nor U19615 (N_19615,N_19424,N_19401);
nand U19616 (N_19616,N_19500,N_19482);
nor U19617 (N_19617,N_19406,N_19447);
nor U19618 (N_19618,N_19488,N_19374);
and U19619 (N_19619,N_19425,N_19460);
xor U19620 (N_19620,N_19402,N_19427);
or U19621 (N_19621,N_19386,N_19484);
nor U19622 (N_19622,N_19448,N_19504);
nor U19623 (N_19623,N_19363,N_19483);
or U19624 (N_19624,N_19405,N_19462);
or U19625 (N_19625,N_19490,N_19368);
nor U19626 (N_19626,N_19378,N_19506);
and U19627 (N_19627,N_19400,N_19379);
and U19628 (N_19628,N_19399,N_19508);
nor U19629 (N_19629,N_19494,N_19399);
or U19630 (N_19630,N_19366,N_19413);
or U19631 (N_19631,N_19360,N_19434);
nand U19632 (N_19632,N_19491,N_19392);
and U19633 (N_19633,N_19378,N_19448);
nand U19634 (N_19634,N_19495,N_19465);
and U19635 (N_19635,N_19414,N_19476);
and U19636 (N_19636,N_19432,N_19386);
xnor U19637 (N_19637,N_19413,N_19516);
and U19638 (N_19638,N_19499,N_19395);
xnor U19639 (N_19639,N_19409,N_19500);
nor U19640 (N_19640,N_19485,N_19398);
nand U19641 (N_19641,N_19429,N_19404);
and U19642 (N_19642,N_19420,N_19362);
xor U19643 (N_19643,N_19469,N_19451);
and U19644 (N_19644,N_19465,N_19429);
and U19645 (N_19645,N_19435,N_19505);
and U19646 (N_19646,N_19391,N_19416);
or U19647 (N_19647,N_19468,N_19484);
or U19648 (N_19648,N_19493,N_19381);
xor U19649 (N_19649,N_19503,N_19375);
nand U19650 (N_19650,N_19418,N_19371);
nor U19651 (N_19651,N_19396,N_19487);
nor U19652 (N_19652,N_19374,N_19360);
or U19653 (N_19653,N_19449,N_19466);
nand U19654 (N_19654,N_19386,N_19446);
or U19655 (N_19655,N_19394,N_19390);
and U19656 (N_19656,N_19451,N_19432);
nor U19657 (N_19657,N_19495,N_19500);
nand U19658 (N_19658,N_19490,N_19427);
nand U19659 (N_19659,N_19364,N_19482);
xnor U19660 (N_19660,N_19367,N_19391);
nor U19661 (N_19661,N_19478,N_19496);
xor U19662 (N_19662,N_19409,N_19471);
or U19663 (N_19663,N_19499,N_19458);
nand U19664 (N_19664,N_19362,N_19393);
nand U19665 (N_19665,N_19509,N_19372);
or U19666 (N_19666,N_19445,N_19518);
nor U19667 (N_19667,N_19478,N_19453);
or U19668 (N_19668,N_19395,N_19443);
or U19669 (N_19669,N_19411,N_19473);
and U19670 (N_19670,N_19518,N_19473);
xor U19671 (N_19671,N_19517,N_19385);
or U19672 (N_19672,N_19423,N_19508);
nor U19673 (N_19673,N_19496,N_19477);
and U19674 (N_19674,N_19429,N_19504);
xor U19675 (N_19675,N_19421,N_19428);
nor U19676 (N_19676,N_19511,N_19441);
and U19677 (N_19677,N_19457,N_19476);
nor U19678 (N_19678,N_19450,N_19436);
nor U19679 (N_19679,N_19384,N_19454);
nor U19680 (N_19680,N_19641,N_19529);
nand U19681 (N_19681,N_19645,N_19588);
or U19682 (N_19682,N_19647,N_19673);
or U19683 (N_19683,N_19571,N_19646);
and U19684 (N_19684,N_19604,N_19637);
or U19685 (N_19685,N_19547,N_19630);
nor U19686 (N_19686,N_19640,N_19525);
and U19687 (N_19687,N_19550,N_19603);
and U19688 (N_19688,N_19595,N_19590);
nand U19689 (N_19689,N_19643,N_19563);
or U19690 (N_19690,N_19530,N_19633);
xnor U19691 (N_19691,N_19629,N_19656);
and U19692 (N_19692,N_19545,N_19541);
and U19693 (N_19693,N_19522,N_19556);
xnor U19694 (N_19694,N_19533,N_19651);
xor U19695 (N_19695,N_19670,N_19674);
and U19696 (N_19696,N_19675,N_19679);
nor U19697 (N_19697,N_19628,N_19653);
nor U19698 (N_19698,N_19557,N_19622);
and U19699 (N_19699,N_19600,N_19583);
xnor U19700 (N_19700,N_19615,N_19672);
xnor U19701 (N_19701,N_19526,N_19542);
or U19702 (N_19702,N_19669,N_19598);
or U19703 (N_19703,N_19568,N_19671);
or U19704 (N_19704,N_19678,N_19562);
and U19705 (N_19705,N_19677,N_19574);
and U19706 (N_19706,N_19523,N_19607);
and U19707 (N_19707,N_19558,N_19618);
nand U19708 (N_19708,N_19614,N_19540);
xor U19709 (N_19709,N_19555,N_19577);
or U19710 (N_19710,N_19593,N_19619);
nand U19711 (N_19711,N_19642,N_19597);
nor U19712 (N_19712,N_19527,N_19548);
nand U19713 (N_19713,N_19602,N_19611);
xnor U19714 (N_19714,N_19639,N_19596);
or U19715 (N_19715,N_19528,N_19636);
nor U19716 (N_19716,N_19662,N_19538);
nand U19717 (N_19717,N_19564,N_19627);
nand U19718 (N_19718,N_19635,N_19632);
nand U19719 (N_19719,N_19581,N_19566);
or U19720 (N_19720,N_19665,N_19524);
nor U19721 (N_19721,N_19549,N_19544);
or U19722 (N_19722,N_19660,N_19658);
xor U19723 (N_19723,N_19573,N_19659);
xor U19724 (N_19724,N_19650,N_19521);
nand U19725 (N_19725,N_19559,N_19605);
nand U19726 (N_19726,N_19621,N_19536);
or U19727 (N_19727,N_19537,N_19613);
nand U19728 (N_19728,N_19617,N_19654);
or U19729 (N_19729,N_19584,N_19589);
or U19730 (N_19730,N_19610,N_19585);
and U19731 (N_19731,N_19520,N_19657);
nand U19732 (N_19732,N_19608,N_19664);
and U19733 (N_19733,N_19539,N_19543);
nor U19734 (N_19734,N_19638,N_19661);
xor U19735 (N_19735,N_19616,N_19572);
xnor U19736 (N_19736,N_19553,N_19592);
or U19737 (N_19737,N_19634,N_19631);
nor U19738 (N_19738,N_19569,N_19612);
or U19739 (N_19739,N_19531,N_19648);
and U19740 (N_19740,N_19580,N_19666);
or U19741 (N_19741,N_19606,N_19579);
nand U19742 (N_19742,N_19576,N_19552);
or U19743 (N_19743,N_19652,N_19554);
xnor U19744 (N_19744,N_19551,N_19575);
nand U19745 (N_19745,N_19570,N_19582);
xor U19746 (N_19746,N_19578,N_19668);
nand U19747 (N_19747,N_19586,N_19626);
or U19748 (N_19748,N_19644,N_19624);
nand U19749 (N_19749,N_19561,N_19655);
xor U19750 (N_19750,N_19594,N_19623);
nor U19751 (N_19751,N_19620,N_19565);
nand U19752 (N_19752,N_19601,N_19599);
nor U19753 (N_19753,N_19591,N_19649);
nand U19754 (N_19754,N_19567,N_19532);
xor U19755 (N_19755,N_19546,N_19560);
nand U19756 (N_19756,N_19534,N_19587);
nand U19757 (N_19757,N_19625,N_19676);
nand U19758 (N_19758,N_19609,N_19663);
nand U19759 (N_19759,N_19535,N_19667);
or U19760 (N_19760,N_19593,N_19625);
xnor U19761 (N_19761,N_19542,N_19630);
nand U19762 (N_19762,N_19577,N_19669);
nand U19763 (N_19763,N_19608,N_19607);
nand U19764 (N_19764,N_19568,N_19626);
and U19765 (N_19765,N_19603,N_19676);
or U19766 (N_19766,N_19536,N_19554);
nor U19767 (N_19767,N_19677,N_19537);
nor U19768 (N_19768,N_19629,N_19664);
nor U19769 (N_19769,N_19639,N_19647);
xnor U19770 (N_19770,N_19535,N_19656);
and U19771 (N_19771,N_19592,N_19673);
nand U19772 (N_19772,N_19549,N_19564);
or U19773 (N_19773,N_19656,N_19540);
nand U19774 (N_19774,N_19590,N_19565);
nand U19775 (N_19775,N_19676,N_19643);
or U19776 (N_19776,N_19673,N_19624);
nand U19777 (N_19777,N_19540,N_19671);
or U19778 (N_19778,N_19643,N_19523);
nor U19779 (N_19779,N_19648,N_19534);
or U19780 (N_19780,N_19654,N_19555);
nor U19781 (N_19781,N_19645,N_19674);
nor U19782 (N_19782,N_19570,N_19524);
or U19783 (N_19783,N_19585,N_19593);
xnor U19784 (N_19784,N_19558,N_19632);
or U19785 (N_19785,N_19616,N_19607);
nand U19786 (N_19786,N_19656,N_19586);
xnor U19787 (N_19787,N_19665,N_19548);
or U19788 (N_19788,N_19647,N_19537);
xnor U19789 (N_19789,N_19579,N_19627);
and U19790 (N_19790,N_19627,N_19567);
and U19791 (N_19791,N_19554,N_19601);
nor U19792 (N_19792,N_19619,N_19626);
xnor U19793 (N_19793,N_19578,N_19559);
or U19794 (N_19794,N_19673,N_19548);
xnor U19795 (N_19795,N_19530,N_19557);
and U19796 (N_19796,N_19589,N_19615);
nor U19797 (N_19797,N_19632,N_19586);
nor U19798 (N_19798,N_19619,N_19587);
nor U19799 (N_19799,N_19572,N_19622);
or U19800 (N_19800,N_19577,N_19578);
xnor U19801 (N_19801,N_19650,N_19537);
nor U19802 (N_19802,N_19629,N_19616);
nor U19803 (N_19803,N_19643,N_19582);
nor U19804 (N_19804,N_19660,N_19565);
nand U19805 (N_19805,N_19639,N_19598);
and U19806 (N_19806,N_19638,N_19564);
nor U19807 (N_19807,N_19593,N_19624);
or U19808 (N_19808,N_19674,N_19647);
nand U19809 (N_19809,N_19558,N_19568);
or U19810 (N_19810,N_19611,N_19521);
xnor U19811 (N_19811,N_19622,N_19605);
nor U19812 (N_19812,N_19641,N_19596);
nand U19813 (N_19813,N_19652,N_19642);
or U19814 (N_19814,N_19556,N_19592);
or U19815 (N_19815,N_19540,N_19552);
or U19816 (N_19816,N_19626,N_19529);
and U19817 (N_19817,N_19667,N_19564);
or U19818 (N_19818,N_19642,N_19623);
nand U19819 (N_19819,N_19625,N_19564);
nand U19820 (N_19820,N_19618,N_19635);
nand U19821 (N_19821,N_19668,N_19637);
or U19822 (N_19822,N_19528,N_19562);
xnor U19823 (N_19823,N_19542,N_19559);
nand U19824 (N_19824,N_19637,N_19643);
nor U19825 (N_19825,N_19522,N_19534);
or U19826 (N_19826,N_19586,N_19643);
nand U19827 (N_19827,N_19664,N_19644);
xnor U19828 (N_19828,N_19659,N_19529);
nor U19829 (N_19829,N_19667,N_19639);
nand U19830 (N_19830,N_19670,N_19522);
or U19831 (N_19831,N_19521,N_19545);
nor U19832 (N_19832,N_19629,N_19543);
nand U19833 (N_19833,N_19679,N_19582);
nand U19834 (N_19834,N_19527,N_19609);
and U19835 (N_19835,N_19650,N_19644);
nand U19836 (N_19836,N_19563,N_19537);
xor U19837 (N_19837,N_19679,N_19636);
or U19838 (N_19838,N_19541,N_19533);
nor U19839 (N_19839,N_19537,N_19541);
xnor U19840 (N_19840,N_19729,N_19701);
or U19841 (N_19841,N_19832,N_19805);
nand U19842 (N_19842,N_19827,N_19694);
nor U19843 (N_19843,N_19717,N_19738);
and U19844 (N_19844,N_19688,N_19782);
nor U19845 (N_19845,N_19806,N_19836);
and U19846 (N_19846,N_19820,N_19807);
xnor U19847 (N_19847,N_19801,N_19690);
nor U19848 (N_19848,N_19795,N_19734);
xor U19849 (N_19849,N_19753,N_19743);
nand U19850 (N_19850,N_19733,N_19839);
nor U19851 (N_19851,N_19787,N_19830);
nand U19852 (N_19852,N_19811,N_19714);
and U19853 (N_19853,N_19772,N_19808);
xor U19854 (N_19854,N_19755,N_19748);
nor U19855 (N_19855,N_19689,N_19725);
xnor U19856 (N_19856,N_19681,N_19696);
and U19857 (N_19857,N_19708,N_19726);
and U19858 (N_19858,N_19684,N_19797);
nor U19859 (N_19859,N_19828,N_19771);
and U19860 (N_19860,N_19803,N_19818);
or U19861 (N_19861,N_19686,N_19758);
xor U19862 (N_19862,N_19724,N_19815);
or U19863 (N_19863,N_19685,N_19826);
nor U19864 (N_19864,N_19773,N_19810);
nor U19865 (N_19865,N_19809,N_19796);
or U19866 (N_19866,N_19819,N_19756);
or U19867 (N_19867,N_19713,N_19709);
or U19868 (N_19868,N_19786,N_19728);
nor U19869 (N_19869,N_19765,N_19779);
xnor U19870 (N_19870,N_19760,N_19802);
nand U19871 (N_19871,N_19784,N_19700);
xnor U19872 (N_19872,N_19682,N_19792);
and U19873 (N_19873,N_19780,N_19835);
xnor U19874 (N_19874,N_19737,N_19716);
nor U19875 (N_19875,N_19798,N_19757);
and U19876 (N_19876,N_19752,N_19719);
xor U19877 (N_19877,N_19769,N_19829);
nor U19878 (N_19878,N_19777,N_19707);
or U19879 (N_19879,N_19804,N_19750);
or U19880 (N_19880,N_19762,N_19747);
and U19881 (N_19881,N_19739,N_19742);
xnor U19882 (N_19882,N_19764,N_19767);
or U19883 (N_19883,N_19781,N_19736);
or U19884 (N_19884,N_19823,N_19703);
and U19885 (N_19885,N_19821,N_19816);
and U19886 (N_19886,N_19741,N_19766);
nand U19887 (N_19887,N_19825,N_19794);
nand U19888 (N_19888,N_19822,N_19793);
and U19889 (N_19889,N_19727,N_19774);
nand U19890 (N_19890,N_19721,N_19761);
nor U19891 (N_19891,N_19702,N_19759);
nor U19892 (N_19892,N_19800,N_19776);
or U19893 (N_19893,N_19732,N_19812);
nor U19894 (N_19894,N_19710,N_19785);
xor U19895 (N_19895,N_19723,N_19744);
or U19896 (N_19896,N_19824,N_19837);
nor U19897 (N_19897,N_19680,N_19746);
nand U19898 (N_19898,N_19720,N_19778);
or U19899 (N_19899,N_19711,N_19789);
nor U19900 (N_19900,N_19788,N_19817);
or U19901 (N_19901,N_19691,N_19749);
or U19902 (N_19902,N_19763,N_19722);
xnor U19903 (N_19903,N_19783,N_19740);
nor U19904 (N_19904,N_19693,N_19692);
xor U19905 (N_19905,N_19754,N_19770);
nor U19906 (N_19906,N_19735,N_19705);
xnor U19907 (N_19907,N_19695,N_19768);
and U19908 (N_19908,N_19683,N_19799);
xor U19909 (N_19909,N_19704,N_19715);
or U19910 (N_19910,N_19791,N_19731);
nand U19911 (N_19911,N_19697,N_19751);
and U19912 (N_19912,N_19699,N_19813);
or U19913 (N_19913,N_19814,N_19745);
nand U19914 (N_19914,N_19831,N_19718);
xnor U19915 (N_19915,N_19698,N_19790);
nand U19916 (N_19916,N_19834,N_19838);
and U19917 (N_19917,N_19712,N_19706);
or U19918 (N_19918,N_19775,N_19833);
nor U19919 (N_19919,N_19730,N_19687);
xnor U19920 (N_19920,N_19733,N_19687);
and U19921 (N_19921,N_19770,N_19706);
and U19922 (N_19922,N_19681,N_19822);
or U19923 (N_19923,N_19752,N_19758);
or U19924 (N_19924,N_19812,N_19794);
nor U19925 (N_19925,N_19836,N_19829);
nand U19926 (N_19926,N_19797,N_19809);
and U19927 (N_19927,N_19801,N_19772);
xor U19928 (N_19928,N_19780,N_19814);
and U19929 (N_19929,N_19743,N_19829);
nor U19930 (N_19930,N_19752,N_19770);
nand U19931 (N_19931,N_19688,N_19834);
nand U19932 (N_19932,N_19815,N_19687);
and U19933 (N_19933,N_19804,N_19718);
nor U19934 (N_19934,N_19806,N_19812);
xor U19935 (N_19935,N_19824,N_19706);
nor U19936 (N_19936,N_19753,N_19748);
xor U19937 (N_19937,N_19754,N_19685);
or U19938 (N_19938,N_19727,N_19731);
and U19939 (N_19939,N_19784,N_19807);
nand U19940 (N_19940,N_19783,N_19743);
or U19941 (N_19941,N_19749,N_19712);
nand U19942 (N_19942,N_19800,N_19795);
nor U19943 (N_19943,N_19811,N_19728);
nor U19944 (N_19944,N_19709,N_19809);
nor U19945 (N_19945,N_19745,N_19712);
nor U19946 (N_19946,N_19720,N_19682);
xnor U19947 (N_19947,N_19775,N_19821);
nand U19948 (N_19948,N_19765,N_19762);
or U19949 (N_19949,N_19767,N_19739);
xor U19950 (N_19950,N_19792,N_19815);
xor U19951 (N_19951,N_19777,N_19804);
nand U19952 (N_19952,N_19764,N_19720);
and U19953 (N_19953,N_19728,N_19732);
xnor U19954 (N_19954,N_19725,N_19838);
or U19955 (N_19955,N_19722,N_19806);
xnor U19956 (N_19956,N_19740,N_19726);
or U19957 (N_19957,N_19725,N_19810);
nor U19958 (N_19958,N_19700,N_19686);
nand U19959 (N_19959,N_19683,N_19785);
and U19960 (N_19960,N_19716,N_19835);
or U19961 (N_19961,N_19762,N_19839);
nor U19962 (N_19962,N_19736,N_19697);
nor U19963 (N_19963,N_19776,N_19790);
and U19964 (N_19964,N_19749,N_19704);
xor U19965 (N_19965,N_19838,N_19825);
or U19966 (N_19966,N_19765,N_19758);
nand U19967 (N_19967,N_19721,N_19803);
nor U19968 (N_19968,N_19683,N_19831);
nor U19969 (N_19969,N_19814,N_19838);
xor U19970 (N_19970,N_19803,N_19707);
nor U19971 (N_19971,N_19783,N_19771);
nand U19972 (N_19972,N_19768,N_19778);
and U19973 (N_19973,N_19706,N_19816);
nor U19974 (N_19974,N_19818,N_19749);
xnor U19975 (N_19975,N_19800,N_19713);
nor U19976 (N_19976,N_19739,N_19685);
xor U19977 (N_19977,N_19704,N_19733);
xor U19978 (N_19978,N_19799,N_19727);
nand U19979 (N_19979,N_19811,N_19786);
nand U19980 (N_19980,N_19815,N_19768);
nor U19981 (N_19981,N_19781,N_19707);
nor U19982 (N_19982,N_19731,N_19806);
nand U19983 (N_19983,N_19712,N_19723);
nor U19984 (N_19984,N_19722,N_19790);
nor U19985 (N_19985,N_19832,N_19724);
nor U19986 (N_19986,N_19832,N_19837);
nand U19987 (N_19987,N_19766,N_19748);
and U19988 (N_19988,N_19718,N_19684);
nand U19989 (N_19989,N_19767,N_19729);
or U19990 (N_19990,N_19815,N_19812);
xor U19991 (N_19991,N_19789,N_19779);
or U19992 (N_19992,N_19791,N_19807);
or U19993 (N_19993,N_19795,N_19834);
or U19994 (N_19994,N_19772,N_19797);
or U19995 (N_19995,N_19766,N_19691);
or U19996 (N_19996,N_19795,N_19700);
or U19997 (N_19997,N_19716,N_19801);
nand U19998 (N_19998,N_19739,N_19704);
or U19999 (N_19999,N_19826,N_19691);
xnor UO_0 (O_0,N_19844,N_19955);
xnor UO_1 (O_1,N_19892,N_19933);
nand UO_2 (O_2,N_19919,N_19874);
and UO_3 (O_3,N_19918,N_19900);
nand UO_4 (O_4,N_19896,N_19932);
xor UO_5 (O_5,N_19886,N_19952);
or UO_6 (O_6,N_19897,N_19857);
and UO_7 (O_7,N_19969,N_19971);
nor UO_8 (O_8,N_19843,N_19945);
and UO_9 (O_9,N_19943,N_19986);
and UO_10 (O_10,N_19953,N_19873);
and UO_11 (O_11,N_19938,N_19976);
nor UO_12 (O_12,N_19987,N_19922);
and UO_13 (O_13,N_19927,N_19931);
or UO_14 (O_14,N_19921,N_19880);
and UO_15 (O_15,N_19942,N_19924);
or UO_16 (O_16,N_19860,N_19913);
xnor UO_17 (O_17,N_19840,N_19983);
and UO_18 (O_18,N_19962,N_19988);
xnor UO_19 (O_19,N_19889,N_19970);
or UO_20 (O_20,N_19887,N_19937);
or UO_21 (O_21,N_19862,N_19984);
nor UO_22 (O_22,N_19972,N_19966);
or UO_23 (O_23,N_19989,N_19968);
xnor UO_24 (O_24,N_19916,N_19948);
or UO_25 (O_25,N_19883,N_19910);
and UO_26 (O_26,N_19863,N_19930);
and UO_27 (O_27,N_19959,N_19894);
nand UO_28 (O_28,N_19929,N_19974);
or UO_29 (O_29,N_19923,N_19902);
or UO_30 (O_30,N_19977,N_19956);
nand UO_31 (O_31,N_19905,N_19973);
and UO_32 (O_32,N_19908,N_19865);
or UO_33 (O_33,N_19926,N_19841);
and UO_34 (O_34,N_19917,N_19994);
or UO_35 (O_35,N_19848,N_19847);
nand UO_36 (O_36,N_19884,N_19999);
and UO_37 (O_37,N_19911,N_19979);
xor UO_38 (O_38,N_19893,N_19998);
or UO_39 (O_39,N_19906,N_19855);
nor UO_40 (O_40,N_19996,N_19870);
or UO_41 (O_41,N_19990,N_19949);
or UO_42 (O_42,N_19914,N_19851);
or UO_43 (O_43,N_19842,N_19891);
xnor UO_44 (O_44,N_19872,N_19935);
xor UO_45 (O_45,N_19915,N_19876);
nand UO_46 (O_46,N_19868,N_19993);
nand UO_47 (O_47,N_19982,N_19944);
xor UO_48 (O_48,N_19980,N_19950);
or UO_49 (O_49,N_19985,N_19925);
nor UO_50 (O_50,N_19947,N_19849);
nand UO_51 (O_51,N_19853,N_19940);
nand UO_52 (O_52,N_19881,N_19899);
nand UO_53 (O_53,N_19920,N_19934);
nand UO_54 (O_54,N_19978,N_19936);
xnor UO_55 (O_55,N_19877,N_19845);
or UO_56 (O_56,N_19941,N_19854);
xor UO_57 (O_57,N_19975,N_19912);
or UO_58 (O_58,N_19939,N_19964);
xnor UO_59 (O_59,N_19928,N_19903);
xor UO_60 (O_60,N_19904,N_19869);
nor UO_61 (O_61,N_19957,N_19991);
nand UO_62 (O_62,N_19965,N_19846);
and UO_63 (O_63,N_19890,N_19954);
or UO_64 (O_64,N_19888,N_19879);
and UO_65 (O_65,N_19875,N_19909);
or UO_66 (O_66,N_19981,N_19967);
or UO_67 (O_67,N_19858,N_19861);
and UO_68 (O_68,N_19871,N_19885);
xor UO_69 (O_69,N_19907,N_19859);
nand UO_70 (O_70,N_19852,N_19856);
or UO_71 (O_71,N_19963,N_19867);
nor UO_72 (O_72,N_19901,N_19866);
xor UO_73 (O_73,N_19850,N_19895);
nand UO_74 (O_74,N_19951,N_19995);
or UO_75 (O_75,N_19898,N_19960);
and UO_76 (O_76,N_19946,N_19882);
nand UO_77 (O_77,N_19864,N_19961);
or UO_78 (O_78,N_19958,N_19878);
or UO_79 (O_79,N_19997,N_19992);
nor UO_80 (O_80,N_19984,N_19901);
nor UO_81 (O_81,N_19895,N_19966);
xor UO_82 (O_82,N_19909,N_19920);
nand UO_83 (O_83,N_19995,N_19957);
and UO_84 (O_84,N_19904,N_19906);
nor UO_85 (O_85,N_19938,N_19914);
xnor UO_86 (O_86,N_19871,N_19886);
or UO_87 (O_87,N_19934,N_19856);
and UO_88 (O_88,N_19965,N_19843);
and UO_89 (O_89,N_19868,N_19918);
or UO_90 (O_90,N_19979,N_19923);
nor UO_91 (O_91,N_19870,N_19866);
and UO_92 (O_92,N_19926,N_19910);
or UO_93 (O_93,N_19917,N_19993);
and UO_94 (O_94,N_19912,N_19959);
nor UO_95 (O_95,N_19938,N_19908);
or UO_96 (O_96,N_19963,N_19880);
nor UO_97 (O_97,N_19928,N_19884);
nand UO_98 (O_98,N_19972,N_19878);
nor UO_99 (O_99,N_19896,N_19935);
nand UO_100 (O_100,N_19993,N_19881);
or UO_101 (O_101,N_19962,N_19936);
or UO_102 (O_102,N_19963,N_19873);
xor UO_103 (O_103,N_19953,N_19901);
nand UO_104 (O_104,N_19902,N_19932);
and UO_105 (O_105,N_19889,N_19939);
nor UO_106 (O_106,N_19981,N_19941);
nor UO_107 (O_107,N_19983,N_19925);
or UO_108 (O_108,N_19846,N_19847);
or UO_109 (O_109,N_19953,N_19899);
nand UO_110 (O_110,N_19996,N_19958);
and UO_111 (O_111,N_19904,N_19860);
nand UO_112 (O_112,N_19884,N_19920);
nor UO_113 (O_113,N_19909,N_19949);
nor UO_114 (O_114,N_19924,N_19915);
and UO_115 (O_115,N_19969,N_19892);
and UO_116 (O_116,N_19901,N_19884);
nor UO_117 (O_117,N_19909,N_19867);
nor UO_118 (O_118,N_19910,N_19907);
xnor UO_119 (O_119,N_19885,N_19845);
or UO_120 (O_120,N_19998,N_19968);
nor UO_121 (O_121,N_19860,N_19900);
nor UO_122 (O_122,N_19920,N_19908);
nand UO_123 (O_123,N_19862,N_19857);
xor UO_124 (O_124,N_19890,N_19988);
xor UO_125 (O_125,N_19889,N_19854);
nand UO_126 (O_126,N_19863,N_19849);
nor UO_127 (O_127,N_19873,N_19983);
nor UO_128 (O_128,N_19971,N_19930);
xor UO_129 (O_129,N_19875,N_19965);
or UO_130 (O_130,N_19953,N_19866);
xnor UO_131 (O_131,N_19866,N_19920);
nor UO_132 (O_132,N_19871,N_19842);
and UO_133 (O_133,N_19873,N_19932);
or UO_134 (O_134,N_19923,N_19842);
or UO_135 (O_135,N_19869,N_19864);
nand UO_136 (O_136,N_19943,N_19993);
nand UO_137 (O_137,N_19966,N_19857);
and UO_138 (O_138,N_19848,N_19861);
nand UO_139 (O_139,N_19931,N_19966);
nor UO_140 (O_140,N_19894,N_19973);
nor UO_141 (O_141,N_19992,N_19972);
nor UO_142 (O_142,N_19959,N_19855);
or UO_143 (O_143,N_19921,N_19961);
or UO_144 (O_144,N_19966,N_19887);
xnor UO_145 (O_145,N_19983,N_19986);
nand UO_146 (O_146,N_19990,N_19978);
nor UO_147 (O_147,N_19927,N_19877);
nor UO_148 (O_148,N_19981,N_19976);
or UO_149 (O_149,N_19944,N_19903);
xnor UO_150 (O_150,N_19972,N_19924);
xnor UO_151 (O_151,N_19952,N_19905);
or UO_152 (O_152,N_19874,N_19862);
and UO_153 (O_153,N_19996,N_19851);
nand UO_154 (O_154,N_19856,N_19916);
xnor UO_155 (O_155,N_19972,N_19995);
nor UO_156 (O_156,N_19992,N_19910);
nor UO_157 (O_157,N_19966,N_19925);
or UO_158 (O_158,N_19876,N_19848);
nor UO_159 (O_159,N_19897,N_19848);
xor UO_160 (O_160,N_19940,N_19944);
or UO_161 (O_161,N_19910,N_19909);
and UO_162 (O_162,N_19867,N_19997);
nor UO_163 (O_163,N_19916,N_19947);
nand UO_164 (O_164,N_19934,N_19861);
nor UO_165 (O_165,N_19884,N_19930);
or UO_166 (O_166,N_19986,N_19913);
xnor UO_167 (O_167,N_19891,N_19921);
nand UO_168 (O_168,N_19972,N_19936);
or UO_169 (O_169,N_19918,N_19970);
xor UO_170 (O_170,N_19948,N_19877);
or UO_171 (O_171,N_19973,N_19884);
and UO_172 (O_172,N_19901,N_19987);
xor UO_173 (O_173,N_19964,N_19887);
and UO_174 (O_174,N_19900,N_19956);
nand UO_175 (O_175,N_19943,N_19996);
nor UO_176 (O_176,N_19905,N_19895);
xnor UO_177 (O_177,N_19880,N_19916);
nor UO_178 (O_178,N_19976,N_19987);
and UO_179 (O_179,N_19880,N_19855);
or UO_180 (O_180,N_19950,N_19919);
or UO_181 (O_181,N_19848,N_19853);
xor UO_182 (O_182,N_19951,N_19924);
nand UO_183 (O_183,N_19978,N_19935);
and UO_184 (O_184,N_19874,N_19905);
and UO_185 (O_185,N_19875,N_19880);
or UO_186 (O_186,N_19908,N_19861);
xnor UO_187 (O_187,N_19890,N_19952);
nor UO_188 (O_188,N_19895,N_19992);
nand UO_189 (O_189,N_19977,N_19965);
and UO_190 (O_190,N_19850,N_19886);
nor UO_191 (O_191,N_19873,N_19841);
xnor UO_192 (O_192,N_19875,N_19936);
xnor UO_193 (O_193,N_19970,N_19947);
or UO_194 (O_194,N_19884,N_19970);
nor UO_195 (O_195,N_19882,N_19974);
nor UO_196 (O_196,N_19909,N_19922);
or UO_197 (O_197,N_19946,N_19944);
or UO_198 (O_198,N_19953,N_19986);
nand UO_199 (O_199,N_19914,N_19961);
or UO_200 (O_200,N_19885,N_19877);
nand UO_201 (O_201,N_19902,N_19997);
xor UO_202 (O_202,N_19875,N_19941);
or UO_203 (O_203,N_19870,N_19953);
nor UO_204 (O_204,N_19874,N_19940);
nor UO_205 (O_205,N_19888,N_19980);
or UO_206 (O_206,N_19980,N_19918);
nor UO_207 (O_207,N_19871,N_19846);
and UO_208 (O_208,N_19934,N_19957);
xor UO_209 (O_209,N_19870,N_19975);
or UO_210 (O_210,N_19881,N_19978);
xor UO_211 (O_211,N_19976,N_19884);
xnor UO_212 (O_212,N_19865,N_19885);
nand UO_213 (O_213,N_19957,N_19971);
xor UO_214 (O_214,N_19890,N_19972);
and UO_215 (O_215,N_19917,N_19900);
xor UO_216 (O_216,N_19918,N_19842);
and UO_217 (O_217,N_19841,N_19894);
xnor UO_218 (O_218,N_19897,N_19972);
nand UO_219 (O_219,N_19867,N_19940);
xnor UO_220 (O_220,N_19998,N_19906);
nor UO_221 (O_221,N_19948,N_19870);
nand UO_222 (O_222,N_19843,N_19885);
xor UO_223 (O_223,N_19924,N_19911);
and UO_224 (O_224,N_19842,N_19956);
and UO_225 (O_225,N_19967,N_19925);
nor UO_226 (O_226,N_19880,N_19964);
nand UO_227 (O_227,N_19888,N_19983);
nand UO_228 (O_228,N_19890,N_19848);
and UO_229 (O_229,N_19888,N_19999);
xor UO_230 (O_230,N_19881,N_19866);
xor UO_231 (O_231,N_19865,N_19935);
nor UO_232 (O_232,N_19852,N_19951);
or UO_233 (O_233,N_19980,N_19880);
or UO_234 (O_234,N_19896,N_19906);
nor UO_235 (O_235,N_19912,N_19924);
or UO_236 (O_236,N_19900,N_19899);
nor UO_237 (O_237,N_19905,N_19861);
nand UO_238 (O_238,N_19865,N_19888);
nand UO_239 (O_239,N_19869,N_19897);
xnor UO_240 (O_240,N_19879,N_19942);
xnor UO_241 (O_241,N_19973,N_19937);
nand UO_242 (O_242,N_19861,N_19996);
or UO_243 (O_243,N_19867,N_19859);
xor UO_244 (O_244,N_19859,N_19882);
nand UO_245 (O_245,N_19877,N_19907);
and UO_246 (O_246,N_19921,N_19899);
and UO_247 (O_247,N_19943,N_19916);
nor UO_248 (O_248,N_19910,N_19881);
and UO_249 (O_249,N_19965,N_19898);
and UO_250 (O_250,N_19980,N_19913);
or UO_251 (O_251,N_19853,N_19864);
and UO_252 (O_252,N_19929,N_19946);
xnor UO_253 (O_253,N_19874,N_19964);
nand UO_254 (O_254,N_19870,N_19885);
nor UO_255 (O_255,N_19951,N_19863);
nand UO_256 (O_256,N_19985,N_19889);
or UO_257 (O_257,N_19970,N_19927);
xor UO_258 (O_258,N_19970,N_19890);
nor UO_259 (O_259,N_19846,N_19918);
or UO_260 (O_260,N_19902,N_19861);
or UO_261 (O_261,N_19959,N_19885);
nand UO_262 (O_262,N_19959,N_19843);
and UO_263 (O_263,N_19962,N_19983);
and UO_264 (O_264,N_19906,N_19869);
or UO_265 (O_265,N_19865,N_19951);
nand UO_266 (O_266,N_19855,N_19989);
nand UO_267 (O_267,N_19897,N_19888);
xnor UO_268 (O_268,N_19952,N_19993);
xor UO_269 (O_269,N_19986,N_19974);
nand UO_270 (O_270,N_19918,N_19869);
xnor UO_271 (O_271,N_19954,N_19875);
and UO_272 (O_272,N_19905,N_19970);
or UO_273 (O_273,N_19965,N_19971);
xnor UO_274 (O_274,N_19938,N_19939);
nor UO_275 (O_275,N_19878,N_19846);
and UO_276 (O_276,N_19855,N_19895);
nand UO_277 (O_277,N_19845,N_19869);
xnor UO_278 (O_278,N_19989,N_19892);
nand UO_279 (O_279,N_19918,N_19912);
xor UO_280 (O_280,N_19883,N_19948);
or UO_281 (O_281,N_19893,N_19986);
xor UO_282 (O_282,N_19966,N_19900);
nor UO_283 (O_283,N_19878,N_19976);
nor UO_284 (O_284,N_19951,N_19848);
xnor UO_285 (O_285,N_19988,N_19928);
nor UO_286 (O_286,N_19945,N_19938);
and UO_287 (O_287,N_19845,N_19911);
and UO_288 (O_288,N_19843,N_19954);
and UO_289 (O_289,N_19988,N_19849);
xnor UO_290 (O_290,N_19961,N_19876);
xor UO_291 (O_291,N_19931,N_19936);
xnor UO_292 (O_292,N_19860,N_19968);
nand UO_293 (O_293,N_19980,N_19902);
nor UO_294 (O_294,N_19847,N_19903);
nand UO_295 (O_295,N_19954,N_19970);
xnor UO_296 (O_296,N_19964,N_19894);
or UO_297 (O_297,N_19848,N_19844);
nor UO_298 (O_298,N_19972,N_19856);
and UO_299 (O_299,N_19960,N_19983);
xnor UO_300 (O_300,N_19976,N_19965);
or UO_301 (O_301,N_19982,N_19922);
or UO_302 (O_302,N_19945,N_19927);
nor UO_303 (O_303,N_19946,N_19976);
or UO_304 (O_304,N_19927,N_19998);
and UO_305 (O_305,N_19932,N_19848);
nand UO_306 (O_306,N_19965,N_19964);
nand UO_307 (O_307,N_19915,N_19920);
nand UO_308 (O_308,N_19923,N_19969);
nor UO_309 (O_309,N_19847,N_19953);
nor UO_310 (O_310,N_19932,N_19868);
or UO_311 (O_311,N_19915,N_19994);
and UO_312 (O_312,N_19941,N_19907);
xor UO_313 (O_313,N_19856,N_19994);
xnor UO_314 (O_314,N_19860,N_19928);
and UO_315 (O_315,N_19913,N_19957);
nor UO_316 (O_316,N_19952,N_19935);
xnor UO_317 (O_317,N_19992,N_19932);
and UO_318 (O_318,N_19930,N_19924);
nand UO_319 (O_319,N_19865,N_19953);
nor UO_320 (O_320,N_19850,N_19979);
or UO_321 (O_321,N_19989,N_19872);
nand UO_322 (O_322,N_19995,N_19947);
nand UO_323 (O_323,N_19891,N_19841);
or UO_324 (O_324,N_19986,N_19861);
or UO_325 (O_325,N_19840,N_19962);
or UO_326 (O_326,N_19868,N_19876);
xor UO_327 (O_327,N_19893,N_19884);
and UO_328 (O_328,N_19917,N_19954);
xnor UO_329 (O_329,N_19878,N_19892);
nand UO_330 (O_330,N_19881,N_19971);
and UO_331 (O_331,N_19974,N_19955);
or UO_332 (O_332,N_19863,N_19891);
and UO_333 (O_333,N_19946,N_19843);
and UO_334 (O_334,N_19908,N_19877);
xor UO_335 (O_335,N_19887,N_19968);
and UO_336 (O_336,N_19855,N_19922);
and UO_337 (O_337,N_19918,N_19845);
nand UO_338 (O_338,N_19860,N_19853);
or UO_339 (O_339,N_19919,N_19960);
and UO_340 (O_340,N_19910,N_19846);
or UO_341 (O_341,N_19948,N_19864);
nor UO_342 (O_342,N_19933,N_19966);
and UO_343 (O_343,N_19896,N_19986);
nor UO_344 (O_344,N_19983,N_19939);
or UO_345 (O_345,N_19867,N_19850);
and UO_346 (O_346,N_19918,N_19876);
and UO_347 (O_347,N_19871,N_19906);
nor UO_348 (O_348,N_19969,N_19921);
and UO_349 (O_349,N_19939,N_19999);
and UO_350 (O_350,N_19895,N_19988);
nand UO_351 (O_351,N_19933,N_19947);
nor UO_352 (O_352,N_19941,N_19945);
or UO_353 (O_353,N_19891,N_19857);
xnor UO_354 (O_354,N_19879,N_19868);
and UO_355 (O_355,N_19912,N_19840);
or UO_356 (O_356,N_19961,N_19954);
xnor UO_357 (O_357,N_19960,N_19950);
or UO_358 (O_358,N_19998,N_19896);
xor UO_359 (O_359,N_19878,N_19931);
or UO_360 (O_360,N_19913,N_19869);
nor UO_361 (O_361,N_19891,N_19911);
or UO_362 (O_362,N_19898,N_19874);
nand UO_363 (O_363,N_19930,N_19948);
xor UO_364 (O_364,N_19977,N_19914);
xor UO_365 (O_365,N_19975,N_19861);
and UO_366 (O_366,N_19968,N_19996);
nand UO_367 (O_367,N_19910,N_19914);
xnor UO_368 (O_368,N_19862,N_19953);
and UO_369 (O_369,N_19860,N_19862);
and UO_370 (O_370,N_19874,N_19963);
nand UO_371 (O_371,N_19960,N_19925);
xor UO_372 (O_372,N_19998,N_19841);
and UO_373 (O_373,N_19877,N_19913);
nor UO_374 (O_374,N_19885,N_19936);
xor UO_375 (O_375,N_19997,N_19989);
or UO_376 (O_376,N_19964,N_19901);
nor UO_377 (O_377,N_19975,N_19852);
or UO_378 (O_378,N_19911,N_19900);
xnor UO_379 (O_379,N_19878,N_19916);
nor UO_380 (O_380,N_19882,N_19850);
xnor UO_381 (O_381,N_19922,N_19961);
nor UO_382 (O_382,N_19913,N_19993);
or UO_383 (O_383,N_19927,N_19883);
nand UO_384 (O_384,N_19979,N_19952);
xnor UO_385 (O_385,N_19941,N_19924);
nand UO_386 (O_386,N_19853,N_19999);
nand UO_387 (O_387,N_19851,N_19956);
nand UO_388 (O_388,N_19872,N_19971);
and UO_389 (O_389,N_19886,N_19901);
or UO_390 (O_390,N_19886,N_19992);
xnor UO_391 (O_391,N_19951,N_19871);
or UO_392 (O_392,N_19956,N_19970);
nand UO_393 (O_393,N_19971,N_19857);
or UO_394 (O_394,N_19929,N_19865);
and UO_395 (O_395,N_19862,N_19900);
nand UO_396 (O_396,N_19982,N_19907);
nor UO_397 (O_397,N_19857,N_19843);
or UO_398 (O_398,N_19916,N_19926);
and UO_399 (O_399,N_19973,N_19860);
xor UO_400 (O_400,N_19900,N_19902);
nand UO_401 (O_401,N_19929,N_19940);
nor UO_402 (O_402,N_19998,N_19929);
and UO_403 (O_403,N_19971,N_19948);
nand UO_404 (O_404,N_19858,N_19845);
or UO_405 (O_405,N_19880,N_19960);
nand UO_406 (O_406,N_19864,N_19944);
or UO_407 (O_407,N_19948,N_19871);
and UO_408 (O_408,N_19906,N_19930);
nand UO_409 (O_409,N_19858,N_19875);
and UO_410 (O_410,N_19947,N_19938);
xor UO_411 (O_411,N_19961,N_19946);
nor UO_412 (O_412,N_19979,N_19909);
and UO_413 (O_413,N_19933,N_19940);
and UO_414 (O_414,N_19886,N_19910);
nand UO_415 (O_415,N_19997,N_19916);
or UO_416 (O_416,N_19860,N_19934);
or UO_417 (O_417,N_19908,N_19939);
or UO_418 (O_418,N_19872,N_19878);
xnor UO_419 (O_419,N_19982,N_19947);
xor UO_420 (O_420,N_19988,N_19853);
nor UO_421 (O_421,N_19895,N_19849);
nor UO_422 (O_422,N_19976,N_19841);
nand UO_423 (O_423,N_19841,N_19840);
xnor UO_424 (O_424,N_19907,N_19929);
xnor UO_425 (O_425,N_19942,N_19864);
and UO_426 (O_426,N_19950,N_19857);
nand UO_427 (O_427,N_19877,N_19911);
and UO_428 (O_428,N_19922,N_19885);
and UO_429 (O_429,N_19893,N_19982);
or UO_430 (O_430,N_19845,N_19972);
xnor UO_431 (O_431,N_19908,N_19869);
nor UO_432 (O_432,N_19985,N_19927);
or UO_433 (O_433,N_19953,N_19993);
or UO_434 (O_434,N_19971,N_19919);
xor UO_435 (O_435,N_19994,N_19965);
xnor UO_436 (O_436,N_19894,N_19846);
or UO_437 (O_437,N_19886,N_19927);
xor UO_438 (O_438,N_19868,N_19988);
nand UO_439 (O_439,N_19929,N_19976);
nor UO_440 (O_440,N_19984,N_19890);
and UO_441 (O_441,N_19877,N_19931);
nor UO_442 (O_442,N_19992,N_19904);
nand UO_443 (O_443,N_19861,N_19917);
nand UO_444 (O_444,N_19920,N_19897);
or UO_445 (O_445,N_19979,N_19862);
or UO_446 (O_446,N_19916,N_19894);
or UO_447 (O_447,N_19938,N_19951);
or UO_448 (O_448,N_19934,N_19873);
nor UO_449 (O_449,N_19939,N_19849);
nor UO_450 (O_450,N_19961,N_19920);
and UO_451 (O_451,N_19901,N_19896);
and UO_452 (O_452,N_19915,N_19916);
nand UO_453 (O_453,N_19897,N_19930);
nor UO_454 (O_454,N_19906,N_19899);
xor UO_455 (O_455,N_19921,N_19999);
or UO_456 (O_456,N_19956,N_19998);
nand UO_457 (O_457,N_19950,N_19974);
xnor UO_458 (O_458,N_19951,N_19926);
or UO_459 (O_459,N_19879,N_19964);
and UO_460 (O_460,N_19854,N_19947);
nand UO_461 (O_461,N_19840,N_19905);
nand UO_462 (O_462,N_19911,N_19919);
nand UO_463 (O_463,N_19953,N_19941);
nor UO_464 (O_464,N_19959,N_19872);
nor UO_465 (O_465,N_19954,N_19886);
nor UO_466 (O_466,N_19903,N_19935);
xor UO_467 (O_467,N_19964,N_19841);
nand UO_468 (O_468,N_19846,N_19916);
and UO_469 (O_469,N_19972,N_19895);
or UO_470 (O_470,N_19920,N_19972);
nor UO_471 (O_471,N_19849,N_19960);
nor UO_472 (O_472,N_19882,N_19926);
or UO_473 (O_473,N_19851,N_19859);
nand UO_474 (O_474,N_19859,N_19966);
and UO_475 (O_475,N_19855,N_19962);
nor UO_476 (O_476,N_19943,N_19927);
xnor UO_477 (O_477,N_19895,N_19981);
or UO_478 (O_478,N_19907,N_19857);
xnor UO_479 (O_479,N_19979,N_19998);
nor UO_480 (O_480,N_19931,N_19922);
and UO_481 (O_481,N_19952,N_19988);
or UO_482 (O_482,N_19942,N_19891);
nand UO_483 (O_483,N_19884,N_19954);
and UO_484 (O_484,N_19947,N_19885);
nand UO_485 (O_485,N_19980,N_19922);
xor UO_486 (O_486,N_19971,N_19927);
and UO_487 (O_487,N_19928,N_19924);
nor UO_488 (O_488,N_19997,N_19943);
nor UO_489 (O_489,N_19959,N_19888);
or UO_490 (O_490,N_19936,N_19864);
nand UO_491 (O_491,N_19938,N_19897);
xnor UO_492 (O_492,N_19841,N_19969);
xnor UO_493 (O_493,N_19851,N_19942);
xnor UO_494 (O_494,N_19923,N_19932);
nor UO_495 (O_495,N_19999,N_19972);
xor UO_496 (O_496,N_19993,N_19885);
nor UO_497 (O_497,N_19849,N_19888);
xor UO_498 (O_498,N_19927,N_19859);
nand UO_499 (O_499,N_19998,N_19942);
nor UO_500 (O_500,N_19914,N_19868);
nand UO_501 (O_501,N_19996,N_19964);
xnor UO_502 (O_502,N_19847,N_19914);
or UO_503 (O_503,N_19996,N_19972);
and UO_504 (O_504,N_19891,N_19953);
nand UO_505 (O_505,N_19871,N_19959);
nor UO_506 (O_506,N_19950,N_19993);
xor UO_507 (O_507,N_19957,N_19894);
nand UO_508 (O_508,N_19909,N_19997);
and UO_509 (O_509,N_19874,N_19910);
nand UO_510 (O_510,N_19936,N_19840);
nor UO_511 (O_511,N_19961,N_19968);
or UO_512 (O_512,N_19967,N_19888);
and UO_513 (O_513,N_19935,N_19846);
nand UO_514 (O_514,N_19897,N_19855);
nand UO_515 (O_515,N_19965,N_19860);
xnor UO_516 (O_516,N_19869,N_19899);
nor UO_517 (O_517,N_19975,N_19895);
or UO_518 (O_518,N_19969,N_19961);
and UO_519 (O_519,N_19986,N_19948);
or UO_520 (O_520,N_19877,N_19891);
and UO_521 (O_521,N_19980,N_19898);
nor UO_522 (O_522,N_19862,N_19962);
or UO_523 (O_523,N_19888,N_19964);
nor UO_524 (O_524,N_19853,N_19863);
or UO_525 (O_525,N_19972,N_19952);
or UO_526 (O_526,N_19899,N_19951);
xnor UO_527 (O_527,N_19996,N_19935);
nand UO_528 (O_528,N_19895,N_19861);
nand UO_529 (O_529,N_19967,N_19983);
and UO_530 (O_530,N_19998,N_19902);
or UO_531 (O_531,N_19912,N_19908);
or UO_532 (O_532,N_19920,N_19900);
nor UO_533 (O_533,N_19892,N_19911);
nor UO_534 (O_534,N_19885,N_19948);
or UO_535 (O_535,N_19912,N_19886);
xor UO_536 (O_536,N_19894,N_19851);
or UO_537 (O_537,N_19858,N_19977);
nand UO_538 (O_538,N_19965,N_19889);
and UO_539 (O_539,N_19979,N_19840);
nor UO_540 (O_540,N_19886,N_19889);
and UO_541 (O_541,N_19991,N_19914);
or UO_542 (O_542,N_19923,N_19922);
xor UO_543 (O_543,N_19925,N_19908);
nand UO_544 (O_544,N_19888,N_19986);
and UO_545 (O_545,N_19951,N_19850);
nand UO_546 (O_546,N_19987,N_19851);
nand UO_547 (O_547,N_19877,N_19882);
nor UO_548 (O_548,N_19901,N_19895);
nor UO_549 (O_549,N_19883,N_19842);
xor UO_550 (O_550,N_19939,N_19950);
and UO_551 (O_551,N_19879,N_19898);
or UO_552 (O_552,N_19992,N_19978);
nand UO_553 (O_553,N_19965,N_19850);
nand UO_554 (O_554,N_19970,N_19983);
nor UO_555 (O_555,N_19843,N_19898);
nand UO_556 (O_556,N_19854,N_19883);
xnor UO_557 (O_557,N_19843,N_19992);
or UO_558 (O_558,N_19892,N_19896);
or UO_559 (O_559,N_19964,N_19857);
and UO_560 (O_560,N_19950,N_19859);
or UO_561 (O_561,N_19875,N_19933);
and UO_562 (O_562,N_19966,N_19964);
and UO_563 (O_563,N_19847,N_19875);
xor UO_564 (O_564,N_19987,N_19917);
nor UO_565 (O_565,N_19860,N_19878);
nor UO_566 (O_566,N_19844,N_19969);
xor UO_567 (O_567,N_19854,N_19982);
xnor UO_568 (O_568,N_19963,N_19850);
nor UO_569 (O_569,N_19871,N_19882);
nand UO_570 (O_570,N_19843,N_19864);
or UO_571 (O_571,N_19933,N_19903);
and UO_572 (O_572,N_19989,N_19879);
nor UO_573 (O_573,N_19848,N_19933);
nor UO_574 (O_574,N_19946,N_19949);
nor UO_575 (O_575,N_19887,N_19998);
nand UO_576 (O_576,N_19923,N_19982);
and UO_577 (O_577,N_19863,N_19992);
or UO_578 (O_578,N_19915,N_19971);
nand UO_579 (O_579,N_19869,N_19993);
nor UO_580 (O_580,N_19985,N_19983);
and UO_581 (O_581,N_19999,N_19844);
nor UO_582 (O_582,N_19979,N_19901);
or UO_583 (O_583,N_19867,N_19995);
nor UO_584 (O_584,N_19906,N_19986);
or UO_585 (O_585,N_19962,N_19887);
or UO_586 (O_586,N_19901,N_19899);
or UO_587 (O_587,N_19996,N_19904);
and UO_588 (O_588,N_19902,N_19947);
nor UO_589 (O_589,N_19859,N_19915);
or UO_590 (O_590,N_19966,N_19865);
or UO_591 (O_591,N_19966,N_19890);
nor UO_592 (O_592,N_19882,N_19935);
nor UO_593 (O_593,N_19902,N_19898);
nand UO_594 (O_594,N_19884,N_19914);
or UO_595 (O_595,N_19972,N_19894);
or UO_596 (O_596,N_19949,N_19995);
or UO_597 (O_597,N_19857,N_19983);
nor UO_598 (O_598,N_19860,N_19989);
nor UO_599 (O_599,N_19905,N_19979);
nand UO_600 (O_600,N_19880,N_19866);
or UO_601 (O_601,N_19979,N_19929);
and UO_602 (O_602,N_19970,N_19843);
and UO_603 (O_603,N_19866,N_19941);
nand UO_604 (O_604,N_19909,N_19880);
or UO_605 (O_605,N_19972,N_19844);
xor UO_606 (O_606,N_19897,N_19935);
nor UO_607 (O_607,N_19901,N_19951);
and UO_608 (O_608,N_19982,N_19975);
and UO_609 (O_609,N_19878,N_19957);
and UO_610 (O_610,N_19906,N_19918);
nor UO_611 (O_611,N_19941,N_19958);
nand UO_612 (O_612,N_19897,N_19947);
and UO_613 (O_613,N_19937,N_19950);
or UO_614 (O_614,N_19950,N_19881);
nand UO_615 (O_615,N_19950,N_19972);
or UO_616 (O_616,N_19923,N_19945);
and UO_617 (O_617,N_19991,N_19941);
xor UO_618 (O_618,N_19868,N_19965);
nand UO_619 (O_619,N_19875,N_19931);
nand UO_620 (O_620,N_19930,N_19898);
or UO_621 (O_621,N_19872,N_19919);
xor UO_622 (O_622,N_19897,N_19998);
nor UO_623 (O_623,N_19934,N_19896);
or UO_624 (O_624,N_19969,N_19914);
or UO_625 (O_625,N_19899,N_19866);
nor UO_626 (O_626,N_19897,N_19963);
and UO_627 (O_627,N_19963,N_19853);
nor UO_628 (O_628,N_19886,N_19956);
nand UO_629 (O_629,N_19955,N_19858);
nor UO_630 (O_630,N_19851,N_19880);
xor UO_631 (O_631,N_19873,N_19864);
or UO_632 (O_632,N_19960,N_19924);
nor UO_633 (O_633,N_19904,N_19978);
or UO_634 (O_634,N_19841,N_19949);
xor UO_635 (O_635,N_19848,N_19925);
and UO_636 (O_636,N_19979,N_19965);
and UO_637 (O_637,N_19892,N_19877);
xor UO_638 (O_638,N_19919,N_19935);
or UO_639 (O_639,N_19949,N_19916);
and UO_640 (O_640,N_19861,N_19967);
xor UO_641 (O_641,N_19978,N_19922);
xnor UO_642 (O_642,N_19905,N_19975);
xnor UO_643 (O_643,N_19868,N_19941);
nand UO_644 (O_644,N_19962,N_19987);
nand UO_645 (O_645,N_19916,N_19993);
and UO_646 (O_646,N_19949,N_19884);
and UO_647 (O_647,N_19986,N_19930);
xnor UO_648 (O_648,N_19869,N_19932);
or UO_649 (O_649,N_19843,N_19861);
nor UO_650 (O_650,N_19924,N_19998);
or UO_651 (O_651,N_19901,N_19949);
nand UO_652 (O_652,N_19874,N_19994);
and UO_653 (O_653,N_19949,N_19871);
or UO_654 (O_654,N_19964,N_19871);
nor UO_655 (O_655,N_19954,N_19915);
and UO_656 (O_656,N_19941,N_19922);
nor UO_657 (O_657,N_19931,N_19857);
xor UO_658 (O_658,N_19899,N_19962);
and UO_659 (O_659,N_19924,N_19858);
nand UO_660 (O_660,N_19956,N_19938);
nor UO_661 (O_661,N_19965,N_19902);
xor UO_662 (O_662,N_19987,N_19885);
xnor UO_663 (O_663,N_19922,N_19888);
nand UO_664 (O_664,N_19875,N_19973);
nand UO_665 (O_665,N_19849,N_19938);
and UO_666 (O_666,N_19841,N_19872);
nor UO_667 (O_667,N_19877,N_19968);
nor UO_668 (O_668,N_19874,N_19872);
nor UO_669 (O_669,N_19858,N_19857);
nand UO_670 (O_670,N_19949,N_19891);
xor UO_671 (O_671,N_19903,N_19894);
and UO_672 (O_672,N_19881,N_19875);
nand UO_673 (O_673,N_19891,N_19936);
xnor UO_674 (O_674,N_19991,N_19899);
or UO_675 (O_675,N_19974,N_19920);
nor UO_676 (O_676,N_19896,N_19949);
nand UO_677 (O_677,N_19931,N_19862);
nor UO_678 (O_678,N_19935,N_19927);
nor UO_679 (O_679,N_19936,N_19860);
nand UO_680 (O_680,N_19954,N_19905);
nor UO_681 (O_681,N_19979,N_19989);
and UO_682 (O_682,N_19975,N_19889);
nor UO_683 (O_683,N_19987,N_19954);
or UO_684 (O_684,N_19923,N_19999);
nor UO_685 (O_685,N_19972,N_19938);
nand UO_686 (O_686,N_19937,N_19982);
nand UO_687 (O_687,N_19935,N_19891);
xnor UO_688 (O_688,N_19887,N_19912);
and UO_689 (O_689,N_19994,N_19946);
nand UO_690 (O_690,N_19875,N_19943);
and UO_691 (O_691,N_19978,N_19957);
and UO_692 (O_692,N_19990,N_19904);
nor UO_693 (O_693,N_19869,N_19960);
nand UO_694 (O_694,N_19860,N_19987);
nand UO_695 (O_695,N_19975,N_19948);
nand UO_696 (O_696,N_19944,N_19959);
or UO_697 (O_697,N_19876,N_19897);
or UO_698 (O_698,N_19863,N_19926);
or UO_699 (O_699,N_19942,N_19880);
nor UO_700 (O_700,N_19886,N_19945);
and UO_701 (O_701,N_19977,N_19852);
xor UO_702 (O_702,N_19959,N_19903);
and UO_703 (O_703,N_19855,N_19908);
and UO_704 (O_704,N_19859,N_19881);
and UO_705 (O_705,N_19862,N_19842);
and UO_706 (O_706,N_19925,N_19876);
and UO_707 (O_707,N_19886,N_19851);
and UO_708 (O_708,N_19993,N_19846);
nor UO_709 (O_709,N_19903,N_19925);
nor UO_710 (O_710,N_19843,N_19956);
nor UO_711 (O_711,N_19953,N_19981);
and UO_712 (O_712,N_19973,N_19890);
nor UO_713 (O_713,N_19904,N_19871);
and UO_714 (O_714,N_19876,N_19967);
xnor UO_715 (O_715,N_19963,N_19886);
nand UO_716 (O_716,N_19905,N_19977);
xor UO_717 (O_717,N_19861,N_19896);
or UO_718 (O_718,N_19936,N_19847);
xnor UO_719 (O_719,N_19998,N_19978);
nor UO_720 (O_720,N_19971,N_19858);
nand UO_721 (O_721,N_19985,N_19957);
and UO_722 (O_722,N_19915,N_19948);
xnor UO_723 (O_723,N_19899,N_19955);
nand UO_724 (O_724,N_19983,N_19893);
or UO_725 (O_725,N_19922,N_19871);
nor UO_726 (O_726,N_19872,N_19928);
nand UO_727 (O_727,N_19936,N_19908);
and UO_728 (O_728,N_19901,N_19954);
nand UO_729 (O_729,N_19847,N_19974);
nor UO_730 (O_730,N_19951,N_19963);
xor UO_731 (O_731,N_19880,N_19895);
and UO_732 (O_732,N_19876,N_19853);
nand UO_733 (O_733,N_19934,N_19972);
nand UO_734 (O_734,N_19955,N_19926);
or UO_735 (O_735,N_19867,N_19989);
nand UO_736 (O_736,N_19931,N_19872);
or UO_737 (O_737,N_19876,N_19858);
nand UO_738 (O_738,N_19958,N_19919);
xnor UO_739 (O_739,N_19912,N_19949);
or UO_740 (O_740,N_19870,N_19941);
nor UO_741 (O_741,N_19997,N_19954);
xor UO_742 (O_742,N_19863,N_19997);
nor UO_743 (O_743,N_19890,N_19957);
and UO_744 (O_744,N_19979,N_19933);
or UO_745 (O_745,N_19949,N_19980);
nor UO_746 (O_746,N_19948,N_19938);
nor UO_747 (O_747,N_19872,N_19857);
or UO_748 (O_748,N_19976,N_19853);
and UO_749 (O_749,N_19879,N_19858);
nand UO_750 (O_750,N_19985,N_19923);
nor UO_751 (O_751,N_19920,N_19871);
xnor UO_752 (O_752,N_19863,N_19865);
xor UO_753 (O_753,N_19863,N_19973);
nor UO_754 (O_754,N_19849,N_19951);
nand UO_755 (O_755,N_19882,N_19886);
xor UO_756 (O_756,N_19957,N_19993);
nor UO_757 (O_757,N_19970,N_19896);
or UO_758 (O_758,N_19991,N_19867);
or UO_759 (O_759,N_19897,N_19932);
nor UO_760 (O_760,N_19969,N_19981);
xnor UO_761 (O_761,N_19869,N_19939);
and UO_762 (O_762,N_19990,N_19912);
nor UO_763 (O_763,N_19892,N_19983);
xnor UO_764 (O_764,N_19930,N_19900);
and UO_765 (O_765,N_19858,N_19926);
nand UO_766 (O_766,N_19916,N_19859);
xnor UO_767 (O_767,N_19937,N_19925);
and UO_768 (O_768,N_19951,N_19947);
or UO_769 (O_769,N_19867,N_19939);
and UO_770 (O_770,N_19991,N_19944);
xor UO_771 (O_771,N_19922,N_19891);
and UO_772 (O_772,N_19945,N_19948);
xnor UO_773 (O_773,N_19955,N_19859);
and UO_774 (O_774,N_19926,N_19888);
nand UO_775 (O_775,N_19999,N_19886);
xor UO_776 (O_776,N_19890,N_19897);
and UO_777 (O_777,N_19985,N_19909);
nand UO_778 (O_778,N_19955,N_19896);
nor UO_779 (O_779,N_19987,N_19853);
nand UO_780 (O_780,N_19934,N_19999);
nor UO_781 (O_781,N_19965,N_19869);
xor UO_782 (O_782,N_19891,N_19995);
nor UO_783 (O_783,N_19945,N_19985);
and UO_784 (O_784,N_19840,N_19966);
xnor UO_785 (O_785,N_19996,N_19956);
nand UO_786 (O_786,N_19977,N_19986);
and UO_787 (O_787,N_19872,N_19859);
nand UO_788 (O_788,N_19894,N_19980);
nand UO_789 (O_789,N_19858,N_19911);
or UO_790 (O_790,N_19993,N_19948);
xnor UO_791 (O_791,N_19998,N_19900);
nand UO_792 (O_792,N_19953,N_19908);
xor UO_793 (O_793,N_19863,N_19886);
or UO_794 (O_794,N_19906,N_19932);
nand UO_795 (O_795,N_19931,N_19866);
xnor UO_796 (O_796,N_19955,N_19850);
nand UO_797 (O_797,N_19873,N_19879);
xor UO_798 (O_798,N_19992,N_19868);
or UO_799 (O_799,N_19971,N_19995);
or UO_800 (O_800,N_19842,N_19916);
nor UO_801 (O_801,N_19998,N_19976);
xor UO_802 (O_802,N_19992,N_19945);
xnor UO_803 (O_803,N_19896,N_19926);
xor UO_804 (O_804,N_19986,N_19844);
and UO_805 (O_805,N_19932,N_19891);
nand UO_806 (O_806,N_19972,N_19962);
nand UO_807 (O_807,N_19856,N_19869);
nand UO_808 (O_808,N_19927,N_19999);
nand UO_809 (O_809,N_19852,N_19936);
or UO_810 (O_810,N_19892,N_19948);
xor UO_811 (O_811,N_19890,N_19855);
nand UO_812 (O_812,N_19940,N_19888);
and UO_813 (O_813,N_19916,N_19841);
xor UO_814 (O_814,N_19977,N_19945);
and UO_815 (O_815,N_19856,N_19847);
or UO_816 (O_816,N_19981,N_19928);
and UO_817 (O_817,N_19960,N_19851);
xnor UO_818 (O_818,N_19861,N_19881);
nand UO_819 (O_819,N_19948,N_19908);
and UO_820 (O_820,N_19876,N_19956);
nand UO_821 (O_821,N_19900,N_19866);
or UO_822 (O_822,N_19840,N_19869);
nor UO_823 (O_823,N_19912,N_19890);
nor UO_824 (O_824,N_19999,N_19885);
xor UO_825 (O_825,N_19916,N_19899);
nand UO_826 (O_826,N_19857,N_19915);
nand UO_827 (O_827,N_19967,N_19897);
nor UO_828 (O_828,N_19953,N_19961);
nand UO_829 (O_829,N_19903,N_19905);
or UO_830 (O_830,N_19983,N_19890);
xnor UO_831 (O_831,N_19992,N_19994);
and UO_832 (O_832,N_19848,N_19898);
or UO_833 (O_833,N_19907,N_19893);
and UO_834 (O_834,N_19845,N_19982);
or UO_835 (O_835,N_19854,N_19959);
or UO_836 (O_836,N_19953,N_19912);
nand UO_837 (O_837,N_19955,N_19925);
and UO_838 (O_838,N_19856,N_19867);
nor UO_839 (O_839,N_19882,N_19885);
or UO_840 (O_840,N_19912,N_19931);
nand UO_841 (O_841,N_19940,N_19873);
xnor UO_842 (O_842,N_19992,N_19966);
nand UO_843 (O_843,N_19902,N_19967);
nor UO_844 (O_844,N_19873,N_19847);
nand UO_845 (O_845,N_19994,N_19925);
and UO_846 (O_846,N_19850,N_19861);
xnor UO_847 (O_847,N_19965,N_19852);
nor UO_848 (O_848,N_19959,N_19971);
and UO_849 (O_849,N_19949,N_19992);
nor UO_850 (O_850,N_19922,N_19906);
xor UO_851 (O_851,N_19971,N_19895);
or UO_852 (O_852,N_19845,N_19968);
nor UO_853 (O_853,N_19990,N_19968);
and UO_854 (O_854,N_19877,N_19840);
nor UO_855 (O_855,N_19941,N_19845);
and UO_856 (O_856,N_19845,N_19907);
nand UO_857 (O_857,N_19995,N_19984);
nor UO_858 (O_858,N_19988,N_19969);
nor UO_859 (O_859,N_19861,N_19910);
and UO_860 (O_860,N_19867,N_19994);
nand UO_861 (O_861,N_19867,N_19895);
xor UO_862 (O_862,N_19930,N_19939);
xnor UO_863 (O_863,N_19910,N_19906);
or UO_864 (O_864,N_19962,N_19891);
or UO_865 (O_865,N_19886,N_19853);
nand UO_866 (O_866,N_19979,N_19871);
nor UO_867 (O_867,N_19866,N_19852);
and UO_868 (O_868,N_19851,N_19964);
nor UO_869 (O_869,N_19874,N_19943);
and UO_870 (O_870,N_19890,N_19950);
nor UO_871 (O_871,N_19973,N_19948);
and UO_872 (O_872,N_19886,N_19933);
or UO_873 (O_873,N_19859,N_19900);
or UO_874 (O_874,N_19920,N_19861);
xnor UO_875 (O_875,N_19985,N_19978);
nand UO_876 (O_876,N_19934,N_19915);
xnor UO_877 (O_877,N_19907,N_19890);
or UO_878 (O_878,N_19873,N_19888);
nor UO_879 (O_879,N_19998,N_19955);
or UO_880 (O_880,N_19870,N_19875);
nor UO_881 (O_881,N_19921,N_19860);
xnor UO_882 (O_882,N_19889,N_19904);
xor UO_883 (O_883,N_19924,N_19904);
xor UO_884 (O_884,N_19907,N_19942);
nor UO_885 (O_885,N_19867,N_19982);
nor UO_886 (O_886,N_19928,N_19957);
nor UO_887 (O_887,N_19969,N_19911);
xnor UO_888 (O_888,N_19927,N_19979);
nand UO_889 (O_889,N_19940,N_19994);
nor UO_890 (O_890,N_19947,N_19959);
nor UO_891 (O_891,N_19902,N_19865);
and UO_892 (O_892,N_19909,N_19877);
nor UO_893 (O_893,N_19906,N_19924);
nand UO_894 (O_894,N_19907,N_19887);
or UO_895 (O_895,N_19951,N_19946);
nand UO_896 (O_896,N_19941,N_19960);
and UO_897 (O_897,N_19888,N_19951);
xnor UO_898 (O_898,N_19965,N_19957);
xor UO_899 (O_899,N_19909,N_19917);
xnor UO_900 (O_900,N_19845,N_19943);
xor UO_901 (O_901,N_19985,N_19862);
nand UO_902 (O_902,N_19893,N_19974);
nand UO_903 (O_903,N_19945,N_19910);
nand UO_904 (O_904,N_19961,N_19858);
or UO_905 (O_905,N_19853,N_19924);
xor UO_906 (O_906,N_19887,N_19926);
and UO_907 (O_907,N_19860,N_19855);
xnor UO_908 (O_908,N_19871,N_19870);
or UO_909 (O_909,N_19943,N_19862);
or UO_910 (O_910,N_19848,N_19995);
nor UO_911 (O_911,N_19881,N_19982);
xnor UO_912 (O_912,N_19942,N_19964);
nand UO_913 (O_913,N_19994,N_19858);
and UO_914 (O_914,N_19887,N_19915);
and UO_915 (O_915,N_19978,N_19993);
and UO_916 (O_916,N_19997,N_19984);
xnor UO_917 (O_917,N_19961,N_19964);
nand UO_918 (O_918,N_19950,N_19934);
or UO_919 (O_919,N_19969,N_19840);
or UO_920 (O_920,N_19843,N_19997);
or UO_921 (O_921,N_19904,N_19873);
or UO_922 (O_922,N_19865,N_19866);
nand UO_923 (O_923,N_19930,N_19853);
nand UO_924 (O_924,N_19892,N_19881);
nand UO_925 (O_925,N_19964,N_19925);
and UO_926 (O_926,N_19901,N_19860);
or UO_927 (O_927,N_19854,N_19927);
or UO_928 (O_928,N_19908,N_19960);
or UO_929 (O_929,N_19987,N_19911);
and UO_930 (O_930,N_19879,N_19886);
nor UO_931 (O_931,N_19882,N_19948);
nor UO_932 (O_932,N_19973,N_19927);
or UO_933 (O_933,N_19966,N_19868);
nor UO_934 (O_934,N_19931,N_19859);
nand UO_935 (O_935,N_19972,N_19862);
or UO_936 (O_936,N_19861,N_19950);
xor UO_937 (O_937,N_19865,N_19934);
xor UO_938 (O_938,N_19981,N_19960);
and UO_939 (O_939,N_19906,N_19985);
xnor UO_940 (O_940,N_19918,N_19954);
and UO_941 (O_941,N_19939,N_19966);
nand UO_942 (O_942,N_19996,N_19868);
nor UO_943 (O_943,N_19981,N_19905);
xnor UO_944 (O_944,N_19869,N_19933);
and UO_945 (O_945,N_19993,N_19920);
xnor UO_946 (O_946,N_19921,N_19985);
and UO_947 (O_947,N_19893,N_19847);
xnor UO_948 (O_948,N_19931,N_19993);
and UO_949 (O_949,N_19997,N_19934);
and UO_950 (O_950,N_19898,N_19927);
or UO_951 (O_951,N_19870,N_19865);
nand UO_952 (O_952,N_19889,N_19863);
xnor UO_953 (O_953,N_19889,N_19868);
xor UO_954 (O_954,N_19945,N_19908);
nor UO_955 (O_955,N_19932,N_19944);
nor UO_956 (O_956,N_19944,N_19956);
and UO_957 (O_957,N_19902,N_19926);
nand UO_958 (O_958,N_19907,N_19969);
and UO_959 (O_959,N_19909,N_19898);
or UO_960 (O_960,N_19886,N_19852);
or UO_961 (O_961,N_19909,N_19943);
nor UO_962 (O_962,N_19854,N_19903);
nand UO_963 (O_963,N_19935,N_19968);
or UO_964 (O_964,N_19944,N_19901);
or UO_965 (O_965,N_19865,N_19856);
nand UO_966 (O_966,N_19995,N_19853);
or UO_967 (O_967,N_19861,N_19963);
xor UO_968 (O_968,N_19989,N_19930);
nand UO_969 (O_969,N_19859,N_19883);
nand UO_970 (O_970,N_19902,N_19883);
or UO_971 (O_971,N_19957,N_19941);
or UO_972 (O_972,N_19910,N_19855);
or UO_973 (O_973,N_19959,N_19862);
and UO_974 (O_974,N_19990,N_19866);
xnor UO_975 (O_975,N_19898,N_19903);
nand UO_976 (O_976,N_19886,N_19958);
xor UO_977 (O_977,N_19850,N_19964);
nor UO_978 (O_978,N_19994,N_19930);
and UO_979 (O_979,N_19883,N_19987);
or UO_980 (O_980,N_19963,N_19902);
or UO_981 (O_981,N_19849,N_19980);
and UO_982 (O_982,N_19890,N_19880);
nand UO_983 (O_983,N_19937,N_19945);
nor UO_984 (O_984,N_19857,N_19949);
and UO_985 (O_985,N_19975,N_19867);
and UO_986 (O_986,N_19959,N_19875);
or UO_987 (O_987,N_19912,N_19849);
nor UO_988 (O_988,N_19870,N_19892);
nor UO_989 (O_989,N_19998,N_19934);
xor UO_990 (O_990,N_19889,N_19972);
nand UO_991 (O_991,N_19921,N_19930);
nor UO_992 (O_992,N_19856,N_19937);
or UO_993 (O_993,N_19888,N_19973);
and UO_994 (O_994,N_19951,N_19994);
and UO_995 (O_995,N_19890,N_19874);
nor UO_996 (O_996,N_19893,N_19977);
nor UO_997 (O_997,N_19963,N_19929);
and UO_998 (O_998,N_19856,N_19926);
nand UO_999 (O_999,N_19956,N_19925);
and UO_1000 (O_1000,N_19919,N_19892);
xnor UO_1001 (O_1001,N_19942,N_19949);
or UO_1002 (O_1002,N_19930,N_19937);
nand UO_1003 (O_1003,N_19966,N_19878);
nor UO_1004 (O_1004,N_19846,N_19956);
nor UO_1005 (O_1005,N_19992,N_19841);
nand UO_1006 (O_1006,N_19874,N_19948);
or UO_1007 (O_1007,N_19907,N_19950);
xor UO_1008 (O_1008,N_19951,N_19846);
and UO_1009 (O_1009,N_19901,N_19931);
nand UO_1010 (O_1010,N_19857,N_19903);
and UO_1011 (O_1011,N_19860,N_19977);
nor UO_1012 (O_1012,N_19981,N_19996);
nor UO_1013 (O_1013,N_19879,N_19930);
and UO_1014 (O_1014,N_19958,N_19877);
or UO_1015 (O_1015,N_19991,N_19873);
xnor UO_1016 (O_1016,N_19840,N_19906);
nand UO_1017 (O_1017,N_19999,N_19957);
nand UO_1018 (O_1018,N_19869,N_19992);
xnor UO_1019 (O_1019,N_19951,N_19959);
nor UO_1020 (O_1020,N_19861,N_19844);
xnor UO_1021 (O_1021,N_19853,N_19871);
and UO_1022 (O_1022,N_19893,N_19883);
nor UO_1023 (O_1023,N_19904,N_19958);
nor UO_1024 (O_1024,N_19979,N_19978);
nand UO_1025 (O_1025,N_19898,N_19886);
nand UO_1026 (O_1026,N_19935,N_19934);
and UO_1027 (O_1027,N_19866,N_19904);
nor UO_1028 (O_1028,N_19975,N_19871);
xor UO_1029 (O_1029,N_19870,N_19931);
nand UO_1030 (O_1030,N_19848,N_19952);
nand UO_1031 (O_1031,N_19921,N_19990);
or UO_1032 (O_1032,N_19998,N_19959);
nor UO_1033 (O_1033,N_19931,N_19971);
xor UO_1034 (O_1034,N_19957,N_19867);
or UO_1035 (O_1035,N_19897,N_19881);
or UO_1036 (O_1036,N_19990,N_19859);
and UO_1037 (O_1037,N_19976,N_19995);
or UO_1038 (O_1038,N_19987,N_19904);
nor UO_1039 (O_1039,N_19929,N_19899);
and UO_1040 (O_1040,N_19997,N_19990);
and UO_1041 (O_1041,N_19975,N_19891);
nor UO_1042 (O_1042,N_19914,N_19949);
and UO_1043 (O_1043,N_19848,N_19982);
nor UO_1044 (O_1044,N_19947,N_19901);
xor UO_1045 (O_1045,N_19849,N_19987);
nor UO_1046 (O_1046,N_19949,N_19948);
nand UO_1047 (O_1047,N_19845,N_19970);
xor UO_1048 (O_1048,N_19898,N_19989);
and UO_1049 (O_1049,N_19950,N_19913);
xor UO_1050 (O_1050,N_19983,N_19905);
and UO_1051 (O_1051,N_19915,N_19959);
nand UO_1052 (O_1052,N_19869,N_19878);
xnor UO_1053 (O_1053,N_19993,N_19878);
nand UO_1054 (O_1054,N_19867,N_19955);
nand UO_1055 (O_1055,N_19968,N_19905);
xnor UO_1056 (O_1056,N_19840,N_19950);
xor UO_1057 (O_1057,N_19974,N_19872);
or UO_1058 (O_1058,N_19898,N_19941);
xor UO_1059 (O_1059,N_19930,N_19909);
nor UO_1060 (O_1060,N_19897,N_19901);
nand UO_1061 (O_1061,N_19915,N_19847);
nor UO_1062 (O_1062,N_19867,N_19998);
xnor UO_1063 (O_1063,N_19869,N_19942);
nor UO_1064 (O_1064,N_19976,N_19863);
nor UO_1065 (O_1065,N_19934,N_19905);
nor UO_1066 (O_1066,N_19992,N_19894);
nor UO_1067 (O_1067,N_19918,N_19958);
xnor UO_1068 (O_1068,N_19976,N_19916);
and UO_1069 (O_1069,N_19886,N_19860);
xor UO_1070 (O_1070,N_19981,N_19851);
nor UO_1071 (O_1071,N_19942,N_19960);
xnor UO_1072 (O_1072,N_19877,N_19975);
nor UO_1073 (O_1073,N_19841,N_19993);
and UO_1074 (O_1074,N_19910,N_19966);
nor UO_1075 (O_1075,N_19892,N_19866);
xor UO_1076 (O_1076,N_19925,N_19852);
nand UO_1077 (O_1077,N_19860,N_19972);
nor UO_1078 (O_1078,N_19877,N_19934);
xnor UO_1079 (O_1079,N_19959,N_19997);
nor UO_1080 (O_1080,N_19898,N_19870);
nand UO_1081 (O_1081,N_19954,N_19994);
nand UO_1082 (O_1082,N_19862,N_19977);
and UO_1083 (O_1083,N_19990,N_19925);
and UO_1084 (O_1084,N_19979,N_19899);
or UO_1085 (O_1085,N_19915,N_19891);
xnor UO_1086 (O_1086,N_19888,N_19899);
xnor UO_1087 (O_1087,N_19984,N_19908);
and UO_1088 (O_1088,N_19970,N_19907);
or UO_1089 (O_1089,N_19975,N_19899);
nand UO_1090 (O_1090,N_19878,N_19956);
and UO_1091 (O_1091,N_19977,N_19959);
and UO_1092 (O_1092,N_19989,N_19884);
or UO_1093 (O_1093,N_19966,N_19862);
nor UO_1094 (O_1094,N_19932,N_19934);
and UO_1095 (O_1095,N_19891,N_19852);
or UO_1096 (O_1096,N_19994,N_19880);
nand UO_1097 (O_1097,N_19955,N_19866);
or UO_1098 (O_1098,N_19888,N_19862);
or UO_1099 (O_1099,N_19883,N_19907);
nor UO_1100 (O_1100,N_19891,N_19866);
or UO_1101 (O_1101,N_19880,N_19848);
and UO_1102 (O_1102,N_19959,N_19993);
and UO_1103 (O_1103,N_19922,N_19841);
nand UO_1104 (O_1104,N_19938,N_19925);
nor UO_1105 (O_1105,N_19996,N_19875);
or UO_1106 (O_1106,N_19872,N_19957);
xnor UO_1107 (O_1107,N_19930,N_19902);
nor UO_1108 (O_1108,N_19916,N_19945);
and UO_1109 (O_1109,N_19920,N_19888);
and UO_1110 (O_1110,N_19841,N_19986);
and UO_1111 (O_1111,N_19869,N_19873);
nor UO_1112 (O_1112,N_19860,N_19841);
nand UO_1113 (O_1113,N_19913,N_19896);
nand UO_1114 (O_1114,N_19846,N_19929);
nand UO_1115 (O_1115,N_19967,N_19997);
and UO_1116 (O_1116,N_19945,N_19844);
or UO_1117 (O_1117,N_19888,N_19961);
nor UO_1118 (O_1118,N_19877,N_19938);
nor UO_1119 (O_1119,N_19995,N_19934);
xor UO_1120 (O_1120,N_19870,N_19855);
nand UO_1121 (O_1121,N_19932,N_19978);
or UO_1122 (O_1122,N_19999,N_19960);
xor UO_1123 (O_1123,N_19977,N_19952);
and UO_1124 (O_1124,N_19993,N_19874);
xor UO_1125 (O_1125,N_19997,N_19887);
nor UO_1126 (O_1126,N_19915,N_19883);
xor UO_1127 (O_1127,N_19983,N_19871);
nand UO_1128 (O_1128,N_19891,N_19880);
xnor UO_1129 (O_1129,N_19944,N_19905);
nand UO_1130 (O_1130,N_19896,N_19859);
nor UO_1131 (O_1131,N_19843,N_19951);
xnor UO_1132 (O_1132,N_19904,N_19847);
nor UO_1133 (O_1133,N_19969,N_19877);
and UO_1134 (O_1134,N_19861,N_19998);
or UO_1135 (O_1135,N_19931,N_19915);
xor UO_1136 (O_1136,N_19840,N_19999);
xor UO_1137 (O_1137,N_19941,N_19857);
and UO_1138 (O_1138,N_19950,N_19965);
nor UO_1139 (O_1139,N_19841,N_19929);
nor UO_1140 (O_1140,N_19963,N_19916);
and UO_1141 (O_1141,N_19900,N_19923);
nand UO_1142 (O_1142,N_19881,N_19965);
xnor UO_1143 (O_1143,N_19986,N_19949);
or UO_1144 (O_1144,N_19850,N_19904);
xnor UO_1145 (O_1145,N_19928,N_19953);
nor UO_1146 (O_1146,N_19928,N_19855);
or UO_1147 (O_1147,N_19849,N_19926);
nand UO_1148 (O_1148,N_19953,N_19936);
or UO_1149 (O_1149,N_19942,N_19930);
nand UO_1150 (O_1150,N_19971,N_19860);
or UO_1151 (O_1151,N_19867,N_19937);
xnor UO_1152 (O_1152,N_19860,N_19894);
nand UO_1153 (O_1153,N_19975,N_19922);
nor UO_1154 (O_1154,N_19892,N_19915);
or UO_1155 (O_1155,N_19986,N_19957);
or UO_1156 (O_1156,N_19914,N_19960);
xnor UO_1157 (O_1157,N_19981,N_19862);
and UO_1158 (O_1158,N_19988,N_19881);
nand UO_1159 (O_1159,N_19913,N_19848);
nor UO_1160 (O_1160,N_19902,N_19977);
or UO_1161 (O_1161,N_19986,N_19970);
or UO_1162 (O_1162,N_19927,N_19948);
or UO_1163 (O_1163,N_19973,N_19915);
and UO_1164 (O_1164,N_19848,N_19917);
or UO_1165 (O_1165,N_19892,N_19853);
xnor UO_1166 (O_1166,N_19899,N_19964);
xnor UO_1167 (O_1167,N_19999,N_19986);
xor UO_1168 (O_1168,N_19994,N_19909);
and UO_1169 (O_1169,N_19915,N_19936);
nor UO_1170 (O_1170,N_19908,N_19928);
or UO_1171 (O_1171,N_19963,N_19894);
and UO_1172 (O_1172,N_19910,N_19952);
xor UO_1173 (O_1173,N_19996,N_19938);
and UO_1174 (O_1174,N_19939,N_19935);
nand UO_1175 (O_1175,N_19955,N_19975);
nand UO_1176 (O_1176,N_19867,N_19946);
nor UO_1177 (O_1177,N_19876,N_19864);
nand UO_1178 (O_1178,N_19914,N_19861);
and UO_1179 (O_1179,N_19901,N_19958);
xnor UO_1180 (O_1180,N_19877,N_19966);
or UO_1181 (O_1181,N_19917,N_19961);
or UO_1182 (O_1182,N_19982,N_19886);
nand UO_1183 (O_1183,N_19848,N_19935);
or UO_1184 (O_1184,N_19929,N_19870);
nor UO_1185 (O_1185,N_19840,N_19967);
nand UO_1186 (O_1186,N_19968,N_19894);
and UO_1187 (O_1187,N_19903,N_19879);
and UO_1188 (O_1188,N_19869,N_19853);
or UO_1189 (O_1189,N_19943,N_19935);
xor UO_1190 (O_1190,N_19976,N_19989);
xor UO_1191 (O_1191,N_19895,N_19856);
nor UO_1192 (O_1192,N_19960,N_19991);
and UO_1193 (O_1193,N_19950,N_19948);
nor UO_1194 (O_1194,N_19974,N_19926);
xnor UO_1195 (O_1195,N_19903,N_19887);
nand UO_1196 (O_1196,N_19899,N_19931);
and UO_1197 (O_1197,N_19911,N_19925);
nand UO_1198 (O_1198,N_19921,N_19937);
nor UO_1199 (O_1199,N_19923,N_19852);
nor UO_1200 (O_1200,N_19993,N_19975);
nand UO_1201 (O_1201,N_19985,N_19981);
nand UO_1202 (O_1202,N_19988,N_19918);
nor UO_1203 (O_1203,N_19954,N_19891);
nand UO_1204 (O_1204,N_19956,N_19919);
nand UO_1205 (O_1205,N_19909,N_19847);
xor UO_1206 (O_1206,N_19966,N_19981);
nand UO_1207 (O_1207,N_19889,N_19857);
nand UO_1208 (O_1208,N_19985,N_19916);
nor UO_1209 (O_1209,N_19912,N_19992);
xnor UO_1210 (O_1210,N_19977,N_19931);
xor UO_1211 (O_1211,N_19947,N_19911);
nand UO_1212 (O_1212,N_19998,N_19871);
and UO_1213 (O_1213,N_19925,N_19954);
nor UO_1214 (O_1214,N_19965,N_19954);
or UO_1215 (O_1215,N_19981,N_19890);
nand UO_1216 (O_1216,N_19915,N_19917);
and UO_1217 (O_1217,N_19962,N_19935);
or UO_1218 (O_1218,N_19993,N_19949);
nand UO_1219 (O_1219,N_19923,N_19909);
nand UO_1220 (O_1220,N_19969,N_19957);
nand UO_1221 (O_1221,N_19914,N_19841);
xor UO_1222 (O_1222,N_19964,N_19861);
or UO_1223 (O_1223,N_19965,N_19906);
xor UO_1224 (O_1224,N_19852,N_19871);
nand UO_1225 (O_1225,N_19893,N_19930);
nand UO_1226 (O_1226,N_19912,N_19997);
and UO_1227 (O_1227,N_19956,N_19937);
and UO_1228 (O_1228,N_19844,N_19932);
nand UO_1229 (O_1229,N_19941,N_19995);
xnor UO_1230 (O_1230,N_19929,N_19867);
nand UO_1231 (O_1231,N_19944,N_19920);
nand UO_1232 (O_1232,N_19902,N_19856);
nor UO_1233 (O_1233,N_19930,N_19978);
or UO_1234 (O_1234,N_19916,N_19898);
nor UO_1235 (O_1235,N_19932,N_19965);
xnor UO_1236 (O_1236,N_19877,N_19857);
and UO_1237 (O_1237,N_19934,N_19965);
xor UO_1238 (O_1238,N_19863,N_19920);
nor UO_1239 (O_1239,N_19906,N_19908);
nor UO_1240 (O_1240,N_19944,N_19875);
xnor UO_1241 (O_1241,N_19843,N_19926);
nand UO_1242 (O_1242,N_19943,N_19888);
nor UO_1243 (O_1243,N_19930,N_19993);
nor UO_1244 (O_1244,N_19982,N_19887);
and UO_1245 (O_1245,N_19885,N_19981);
or UO_1246 (O_1246,N_19998,N_19939);
xor UO_1247 (O_1247,N_19861,N_19863);
nor UO_1248 (O_1248,N_19960,N_19901);
nor UO_1249 (O_1249,N_19872,N_19984);
nand UO_1250 (O_1250,N_19932,N_19999);
nor UO_1251 (O_1251,N_19902,N_19846);
nand UO_1252 (O_1252,N_19971,N_19986);
xor UO_1253 (O_1253,N_19900,N_19950);
nand UO_1254 (O_1254,N_19863,N_19894);
xnor UO_1255 (O_1255,N_19896,N_19876);
xor UO_1256 (O_1256,N_19968,N_19873);
and UO_1257 (O_1257,N_19943,N_19933);
and UO_1258 (O_1258,N_19888,N_19855);
and UO_1259 (O_1259,N_19865,N_19999);
nand UO_1260 (O_1260,N_19990,N_19950);
nand UO_1261 (O_1261,N_19980,N_19858);
or UO_1262 (O_1262,N_19970,N_19851);
and UO_1263 (O_1263,N_19953,N_19861);
or UO_1264 (O_1264,N_19851,N_19847);
and UO_1265 (O_1265,N_19854,N_19857);
nor UO_1266 (O_1266,N_19974,N_19871);
nand UO_1267 (O_1267,N_19937,N_19866);
nand UO_1268 (O_1268,N_19896,N_19984);
or UO_1269 (O_1269,N_19921,N_19986);
nor UO_1270 (O_1270,N_19951,N_19956);
and UO_1271 (O_1271,N_19850,N_19840);
and UO_1272 (O_1272,N_19935,N_19883);
xor UO_1273 (O_1273,N_19985,N_19937);
or UO_1274 (O_1274,N_19969,N_19983);
nor UO_1275 (O_1275,N_19981,N_19936);
xor UO_1276 (O_1276,N_19990,N_19852);
nand UO_1277 (O_1277,N_19949,N_19972);
xor UO_1278 (O_1278,N_19846,N_19992);
or UO_1279 (O_1279,N_19855,N_19842);
xnor UO_1280 (O_1280,N_19979,N_19950);
or UO_1281 (O_1281,N_19873,N_19998);
nor UO_1282 (O_1282,N_19929,N_19955);
nor UO_1283 (O_1283,N_19943,N_19918);
xor UO_1284 (O_1284,N_19865,N_19855);
and UO_1285 (O_1285,N_19868,N_19881);
nand UO_1286 (O_1286,N_19848,N_19896);
nor UO_1287 (O_1287,N_19928,N_19901);
nor UO_1288 (O_1288,N_19970,N_19959);
nand UO_1289 (O_1289,N_19845,N_19908);
and UO_1290 (O_1290,N_19964,N_19998);
or UO_1291 (O_1291,N_19871,N_19921);
xor UO_1292 (O_1292,N_19925,N_19883);
xnor UO_1293 (O_1293,N_19955,N_19902);
or UO_1294 (O_1294,N_19935,N_19949);
nand UO_1295 (O_1295,N_19916,N_19920);
nand UO_1296 (O_1296,N_19937,N_19929);
or UO_1297 (O_1297,N_19970,N_19924);
and UO_1298 (O_1298,N_19864,N_19931);
or UO_1299 (O_1299,N_19882,N_19939);
nor UO_1300 (O_1300,N_19872,N_19842);
nor UO_1301 (O_1301,N_19928,N_19963);
nor UO_1302 (O_1302,N_19912,N_19927);
or UO_1303 (O_1303,N_19893,N_19901);
nand UO_1304 (O_1304,N_19973,N_19954);
or UO_1305 (O_1305,N_19944,N_19983);
nor UO_1306 (O_1306,N_19956,N_19860);
and UO_1307 (O_1307,N_19953,N_19955);
xnor UO_1308 (O_1308,N_19984,N_19979);
and UO_1309 (O_1309,N_19994,N_19949);
or UO_1310 (O_1310,N_19972,N_19963);
nor UO_1311 (O_1311,N_19885,N_19901);
or UO_1312 (O_1312,N_19889,N_19907);
nand UO_1313 (O_1313,N_19954,N_19897);
and UO_1314 (O_1314,N_19864,N_19981);
or UO_1315 (O_1315,N_19953,N_19897);
and UO_1316 (O_1316,N_19893,N_19973);
xor UO_1317 (O_1317,N_19933,N_19948);
or UO_1318 (O_1318,N_19920,N_19958);
and UO_1319 (O_1319,N_19867,N_19951);
xor UO_1320 (O_1320,N_19882,N_19851);
nand UO_1321 (O_1321,N_19882,N_19873);
xor UO_1322 (O_1322,N_19924,N_19989);
and UO_1323 (O_1323,N_19921,N_19894);
nor UO_1324 (O_1324,N_19953,N_19958);
xnor UO_1325 (O_1325,N_19992,N_19989);
and UO_1326 (O_1326,N_19885,N_19849);
and UO_1327 (O_1327,N_19842,N_19860);
xor UO_1328 (O_1328,N_19880,N_19868);
or UO_1329 (O_1329,N_19944,N_19904);
and UO_1330 (O_1330,N_19934,N_19874);
xnor UO_1331 (O_1331,N_19873,N_19984);
xor UO_1332 (O_1332,N_19965,N_19915);
nand UO_1333 (O_1333,N_19964,N_19993);
and UO_1334 (O_1334,N_19868,N_19842);
nor UO_1335 (O_1335,N_19998,N_19980);
nor UO_1336 (O_1336,N_19852,N_19997);
or UO_1337 (O_1337,N_19964,N_19883);
xor UO_1338 (O_1338,N_19841,N_19999);
and UO_1339 (O_1339,N_19917,N_19908);
nor UO_1340 (O_1340,N_19996,N_19872);
and UO_1341 (O_1341,N_19977,N_19843);
or UO_1342 (O_1342,N_19996,N_19910);
nand UO_1343 (O_1343,N_19941,N_19881);
and UO_1344 (O_1344,N_19969,N_19922);
or UO_1345 (O_1345,N_19848,N_19907);
nor UO_1346 (O_1346,N_19855,N_19898);
xor UO_1347 (O_1347,N_19898,N_19975);
and UO_1348 (O_1348,N_19975,N_19947);
xor UO_1349 (O_1349,N_19997,N_19862);
and UO_1350 (O_1350,N_19911,N_19852);
nor UO_1351 (O_1351,N_19852,N_19912);
nor UO_1352 (O_1352,N_19854,N_19864);
xnor UO_1353 (O_1353,N_19859,N_19984);
and UO_1354 (O_1354,N_19920,N_19983);
and UO_1355 (O_1355,N_19867,N_19996);
nor UO_1356 (O_1356,N_19875,N_19903);
nor UO_1357 (O_1357,N_19917,N_19898);
nand UO_1358 (O_1358,N_19970,N_19897);
nand UO_1359 (O_1359,N_19898,N_19873);
and UO_1360 (O_1360,N_19880,N_19950);
or UO_1361 (O_1361,N_19975,N_19962);
or UO_1362 (O_1362,N_19921,N_19900);
or UO_1363 (O_1363,N_19874,N_19907);
and UO_1364 (O_1364,N_19965,N_19888);
nor UO_1365 (O_1365,N_19946,N_19849);
nand UO_1366 (O_1366,N_19861,N_19878);
and UO_1367 (O_1367,N_19889,N_19990);
xor UO_1368 (O_1368,N_19930,N_19998);
nor UO_1369 (O_1369,N_19950,N_19851);
or UO_1370 (O_1370,N_19929,N_19888);
or UO_1371 (O_1371,N_19929,N_19901);
xnor UO_1372 (O_1372,N_19983,N_19945);
nand UO_1373 (O_1373,N_19951,N_19925);
nand UO_1374 (O_1374,N_19948,N_19936);
or UO_1375 (O_1375,N_19854,N_19976);
nor UO_1376 (O_1376,N_19958,N_19921);
nor UO_1377 (O_1377,N_19856,N_19991);
nand UO_1378 (O_1378,N_19947,N_19999);
nor UO_1379 (O_1379,N_19881,N_19916);
or UO_1380 (O_1380,N_19980,N_19989);
or UO_1381 (O_1381,N_19850,N_19952);
nand UO_1382 (O_1382,N_19858,N_19922);
xor UO_1383 (O_1383,N_19994,N_19919);
xnor UO_1384 (O_1384,N_19933,N_19909);
nor UO_1385 (O_1385,N_19906,N_19958);
xor UO_1386 (O_1386,N_19934,N_19952);
nor UO_1387 (O_1387,N_19938,N_19859);
or UO_1388 (O_1388,N_19840,N_19844);
nor UO_1389 (O_1389,N_19907,N_19938);
and UO_1390 (O_1390,N_19906,N_19945);
nor UO_1391 (O_1391,N_19992,N_19956);
nand UO_1392 (O_1392,N_19918,N_19853);
nand UO_1393 (O_1393,N_19931,N_19943);
nor UO_1394 (O_1394,N_19957,N_19984);
or UO_1395 (O_1395,N_19855,N_19968);
nor UO_1396 (O_1396,N_19976,N_19896);
nor UO_1397 (O_1397,N_19843,N_19845);
or UO_1398 (O_1398,N_19972,N_19883);
and UO_1399 (O_1399,N_19897,N_19902);
xnor UO_1400 (O_1400,N_19891,N_19855);
nor UO_1401 (O_1401,N_19903,N_19861);
and UO_1402 (O_1402,N_19904,N_19863);
nand UO_1403 (O_1403,N_19844,N_19909);
xor UO_1404 (O_1404,N_19875,N_19860);
and UO_1405 (O_1405,N_19913,N_19996);
nand UO_1406 (O_1406,N_19861,N_19840);
xor UO_1407 (O_1407,N_19949,N_19931);
xnor UO_1408 (O_1408,N_19966,N_19870);
xor UO_1409 (O_1409,N_19957,N_19883);
nor UO_1410 (O_1410,N_19891,N_19895);
xnor UO_1411 (O_1411,N_19959,N_19905);
nand UO_1412 (O_1412,N_19947,N_19890);
nor UO_1413 (O_1413,N_19891,N_19872);
and UO_1414 (O_1414,N_19990,N_19896);
nand UO_1415 (O_1415,N_19938,N_19889);
or UO_1416 (O_1416,N_19903,N_19916);
nor UO_1417 (O_1417,N_19916,N_19917);
or UO_1418 (O_1418,N_19930,N_19949);
nand UO_1419 (O_1419,N_19857,N_19994);
or UO_1420 (O_1420,N_19885,N_19950);
and UO_1421 (O_1421,N_19900,N_19988);
or UO_1422 (O_1422,N_19903,N_19868);
or UO_1423 (O_1423,N_19983,N_19963);
or UO_1424 (O_1424,N_19857,N_19894);
nand UO_1425 (O_1425,N_19945,N_19978);
or UO_1426 (O_1426,N_19936,N_19988);
nand UO_1427 (O_1427,N_19843,N_19849);
nor UO_1428 (O_1428,N_19991,N_19881);
xnor UO_1429 (O_1429,N_19903,N_19922);
and UO_1430 (O_1430,N_19925,N_19933);
or UO_1431 (O_1431,N_19997,N_19861);
xor UO_1432 (O_1432,N_19978,N_19974);
and UO_1433 (O_1433,N_19907,N_19992);
xor UO_1434 (O_1434,N_19969,N_19928);
or UO_1435 (O_1435,N_19942,N_19889);
nor UO_1436 (O_1436,N_19852,N_19978);
nand UO_1437 (O_1437,N_19866,N_19864);
and UO_1438 (O_1438,N_19889,N_19964);
xnor UO_1439 (O_1439,N_19893,N_19900);
or UO_1440 (O_1440,N_19945,N_19925);
or UO_1441 (O_1441,N_19917,N_19853);
nand UO_1442 (O_1442,N_19940,N_19939);
nand UO_1443 (O_1443,N_19854,N_19899);
xor UO_1444 (O_1444,N_19932,N_19919);
and UO_1445 (O_1445,N_19879,N_19938);
and UO_1446 (O_1446,N_19892,N_19912);
xnor UO_1447 (O_1447,N_19982,N_19935);
xor UO_1448 (O_1448,N_19888,N_19946);
xnor UO_1449 (O_1449,N_19888,N_19933);
xnor UO_1450 (O_1450,N_19929,N_19961);
nor UO_1451 (O_1451,N_19960,N_19967);
xnor UO_1452 (O_1452,N_19844,N_19903);
nand UO_1453 (O_1453,N_19978,N_19991);
and UO_1454 (O_1454,N_19886,N_19846);
and UO_1455 (O_1455,N_19922,N_19962);
nand UO_1456 (O_1456,N_19969,N_19990);
or UO_1457 (O_1457,N_19995,N_19909);
xor UO_1458 (O_1458,N_19846,N_19849);
nand UO_1459 (O_1459,N_19989,N_19925);
nand UO_1460 (O_1460,N_19940,N_19914);
and UO_1461 (O_1461,N_19940,N_19883);
nand UO_1462 (O_1462,N_19876,N_19912);
nor UO_1463 (O_1463,N_19866,N_19875);
xor UO_1464 (O_1464,N_19954,N_19898);
nor UO_1465 (O_1465,N_19911,N_19897);
xnor UO_1466 (O_1466,N_19883,N_19962);
nor UO_1467 (O_1467,N_19946,N_19940);
nor UO_1468 (O_1468,N_19886,N_19859);
nand UO_1469 (O_1469,N_19916,N_19852);
nor UO_1470 (O_1470,N_19875,N_19994);
nor UO_1471 (O_1471,N_19979,N_19898);
nor UO_1472 (O_1472,N_19845,N_19871);
nor UO_1473 (O_1473,N_19979,N_19842);
nand UO_1474 (O_1474,N_19845,N_19988);
nor UO_1475 (O_1475,N_19995,N_19843);
and UO_1476 (O_1476,N_19858,N_19912);
nand UO_1477 (O_1477,N_19919,N_19959);
and UO_1478 (O_1478,N_19942,N_19935);
nor UO_1479 (O_1479,N_19930,N_19963);
and UO_1480 (O_1480,N_19962,N_19980);
or UO_1481 (O_1481,N_19891,N_19941);
or UO_1482 (O_1482,N_19964,N_19878);
or UO_1483 (O_1483,N_19892,N_19991);
and UO_1484 (O_1484,N_19895,N_19886);
and UO_1485 (O_1485,N_19992,N_19896);
nand UO_1486 (O_1486,N_19842,N_19993);
or UO_1487 (O_1487,N_19990,N_19856);
and UO_1488 (O_1488,N_19999,N_19910);
nor UO_1489 (O_1489,N_19989,N_19946);
xor UO_1490 (O_1490,N_19989,N_19990);
nor UO_1491 (O_1491,N_19844,N_19917);
and UO_1492 (O_1492,N_19921,N_19947);
or UO_1493 (O_1493,N_19936,N_19855);
nor UO_1494 (O_1494,N_19957,N_19893);
or UO_1495 (O_1495,N_19876,N_19960);
or UO_1496 (O_1496,N_19955,N_19951);
nand UO_1497 (O_1497,N_19963,N_19955);
or UO_1498 (O_1498,N_19897,N_19887);
or UO_1499 (O_1499,N_19901,N_19887);
and UO_1500 (O_1500,N_19996,N_19849);
nand UO_1501 (O_1501,N_19944,N_19980);
and UO_1502 (O_1502,N_19917,N_19904);
or UO_1503 (O_1503,N_19963,N_19946);
xnor UO_1504 (O_1504,N_19920,N_19927);
or UO_1505 (O_1505,N_19869,N_19880);
xnor UO_1506 (O_1506,N_19993,N_19908);
nand UO_1507 (O_1507,N_19940,N_19982);
xor UO_1508 (O_1508,N_19992,N_19890);
and UO_1509 (O_1509,N_19942,N_19989);
nor UO_1510 (O_1510,N_19932,N_19945);
nor UO_1511 (O_1511,N_19878,N_19898);
or UO_1512 (O_1512,N_19950,N_19967);
nand UO_1513 (O_1513,N_19902,N_19866);
nor UO_1514 (O_1514,N_19859,N_19875);
xor UO_1515 (O_1515,N_19906,N_19914);
nand UO_1516 (O_1516,N_19944,N_19869);
or UO_1517 (O_1517,N_19965,N_19931);
or UO_1518 (O_1518,N_19887,N_19859);
nor UO_1519 (O_1519,N_19980,N_19975);
nor UO_1520 (O_1520,N_19935,N_19894);
or UO_1521 (O_1521,N_19959,N_19969);
nor UO_1522 (O_1522,N_19857,N_19961);
nand UO_1523 (O_1523,N_19845,N_19894);
or UO_1524 (O_1524,N_19918,N_19888);
or UO_1525 (O_1525,N_19913,N_19863);
nor UO_1526 (O_1526,N_19943,N_19863);
xnor UO_1527 (O_1527,N_19958,N_19978);
and UO_1528 (O_1528,N_19899,N_19864);
xor UO_1529 (O_1529,N_19993,N_19840);
or UO_1530 (O_1530,N_19997,N_19986);
xor UO_1531 (O_1531,N_19951,N_19922);
nand UO_1532 (O_1532,N_19954,N_19859);
and UO_1533 (O_1533,N_19854,N_19990);
nor UO_1534 (O_1534,N_19855,N_19974);
nor UO_1535 (O_1535,N_19976,N_19851);
or UO_1536 (O_1536,N_19883,N_19971);
nor UO_1537 (O_1537,N_19966,N_19881);
xnor UO_1538 (O_1538,N_19994,N_19964);
xnor UO_1539 (O_1539,N_19874,N_19861);
or UO_1540 (O_1540,N_19910,N_19879);
and UO_1541 (O_1541,N_19988,N_19887);
or UO_1542 (O_1542,N_19995,N_19969);
and UO_1543 (O_1543,N_19963,N_19868);
and UO_1544 (O_1544,N_19946,N_19847);
and UO_1545 (O_1545,N_19897,N_19894);
nand UO_1546 (O_1546,N_19961,N_19866);
and UO_1547 (O_1547,N_19945,N_19986);
nor UO_1548 (O_1548,N_19884,N_19916);
nand UO_1549 (O_1549,N_19872,N_19899);
and UO_1550 (O_1550,N_19954,N_19977);
xor UO_1551 (O_1551,N_19989,N_19953);
nor UO_1552 (O_1552,N_19943,N_19976);
nand UO_1553 (O_1553,N_19935,N_19966);
nor UO_1554 (O_1554,N_19869,N_19889);
nor UO_1555 (O_1555,N_19895,N_19846);
and UO_1556 (O_1556,N_19994,N_19850);
xnor UO_1557 (O_1557,N_19893,N_19947);
xor UO_1558 (O_1558,N_19875,N_19901);
nor UO_1559 (O_1559,N_19900,N_19896);
or UO_1560 (O_1560,N_19950,N_19966);
nor UO_1561 (O_1561,N_19869,N_19955);
nand UO_1562 (O_1562,N_19961,N_19983);
and UO_1563 (O_1563,N_19862,N_19894);
nor UO_1564 (O_1564,N_19993,N_19972);
xnor UO_1565 (O_1565,N_19902,N_19957);
xor UO_1566 (O_1566,N_19990,N_19928);
nand UO_1567 (O_1567,N_19870,N_19859);
nor UO_1568 (O_1568,N_19912,N_19991);
nor UO_1569 (O_1569,N_19923,N_19844);
nor UO_1570 (O_1570,N_19983,N_19965);
and UO_1571 (O_1571,N_19859,N_19979);
and UO_1572 (O_1572,N_19842,N_19850);
xor UO_1573 (O_1573,N_19998,N_19844);
or UO_1574 (O_1574,N_19932,N_19924);
nand UO_1575 (O_1575,N_19969,N_19859);
and UO_1576 (O_1576,N_19980,N_19947);
and UO_1577 (O_1577,N_19978,N_19981);
nand UO_1578 (O_1578,N_19960,N_19890);
xnor UO_1579 (O_1579,N_19898,N_19964);
and UO_1580 (O_1580,N_19991,N_19888);
and UO_1581 (O_1581,N_19876,N_19989);
nand UO_1582 (O_1582,N_19893,N_19975);
nor UO_1583 (O_1583,N_19959,N_19876);
and UO_1584 (O_1584,N_19924,N_19894);
xnor UO_1585 (O_1585,N_19983,N_19987);
and UO_1586 (O_1586,N_19859,N_19924);
nand UO_1587 (O_1587,N_19840,N_19976);
or UO_1588 (O_1588,N_19957,N_19849);
and UO_1589 (O_1589,N_19971,N_19892);
or UO_1590 (O_1590,N_19982,N_19972);
nand UO_1591 (O_1591,N_19879,N_19967);
nand UO_1592 (O_1592,N_19911,N_19996);
xor UO_1593 (O_1593,N_19968,N_19900);
nand UO_1594 (O_1594,N_19874,N_19850);
xor UO_1595 (O_1595,N_19989,N_19960);
or UO_1596 (O_1596,N_19957,N_19926);
xor UO_1597 (O_1597,N_19869,N_19956);
nor UO_1598 (O_1598,N_19910,N_19842);
and UO_1599 (O_1599,N_19869,N_19978);
or UO_1600 (O_1600,N_19926,N_19868);
nor UO_1601 (O_1601,N_19847,N_19889);
nor UO_1602 (O_1602,N_19860,N_19945);
nand UO_1603 (O_1603,N_19891,N_19860);
nand UO_1604 (O_1604,N_19908,N_19969);
nor UO_1605 (O_1605,N_19843,N_19848);
or UO_1606 (O_1606,N_19907,N_19960);
nor UO_1607 (O_1607,N_19885,N_19953);
xnor UO_1608 (O_1608,N_19857,N_19905);
and UO_1609 (O_1609,N_19877,N_19946);
xnor UO_1610 (O_1610,N_19868,N_19960);
or UO_1611 (O_1611,N_19920,N_19971);
xnor UO_1612 (O_1612,N_19942,N_19840);
nand UO_1613 (O_1613,N_19939,N_19982);
xor UO_1614 (O_1614,N_19894,N_19955);
and UO_1615 (O_1615,N_19924,N_19956);
xor UO_1616 (O_1616,N_19890,N_19978);
nor UO_1617 (O_1617,N_19940,N_19868);
or UO_1618 (O_1618,N_19881,N_19970);
nor UO_1619 (O_1619,N_19865,N_19988);
and UO_1620 (O_1620,N_19884,N_19855);
and UO_1621 (O_1621,N_19963,N_19855);
xnor UO_1622 (O_1622,N_19923,N_19926);
or UO_1623 (O_1623,N_19865,N_19921);
xnor UO_1624 (O_1624,N_19949,N_19960);
and UO_1625 (O_1625,N_19939,N_19858);
nor UO_1626 (O_1626,N_19840,N_19866);
nor UO_1627 (O_1627,N_19999,N_19895);
xor UO_1628 (O_1628,N_19971,N_19962);
and UO_1629 (O_1629,N_19955,N_19954);
or UO_1630 (O_1630,N_19960,N_19988);
nor UO_1631 (O_1631,N_19972,N_19978);
or UO_1632 (O_1632,N_19971,N_19897);
nor UO_1633 (O_1633,N_19868,N_19983);
xor UO_1634 (O_1634,N_19954,N_19876);
or UO_1635 (O_1635,N_19944,N_19896);
and UO_1636 (O_1636,N_19852,N_19878);
nand UO_1637 (O_1637,N_19947,N_19925);
or UO_1638 (O_1638,N_19879,N_19978);
nor UO_1639 (O_1639,N_19891,N_19978);
nor UO_1640 (O_1640,N_19973,N_19953);
xor UO_1641 (O_1641,N_19885,N_19991);
xor UO_1642 (O_1642,N_19976,N_19994);
nor UO_1643 (O_1643,N_19933,N_19863);
nor UO_1644 (O_1644,N_19874,N_19871);
nor UO_1645 (O_1645,N_19894,N_19908);
or UO_1646 (O_1646,N_19882,N_19840);
nand UO_1647 (O_1647,N_19930,N_19873);
nand UO_1648 (O_1648,N_19841,N_19879);
or UO_1649 (O_1649,N_19870,N_19974);
nand UO_1650 (O_1650,N_19993,N_19967);
xnor UO_1651 (O_1651,N_19887,N_19922);
or UO_1652 (O_1652,N_19978,N_19987);
xor UO_1653 (O_1653,N_19927,N_19847);
nand UO_1654 (O_1654,N_19974,N_19843);
xor UO_1655 (O_1655,N_19976,N_19928);
and UO_1656 (O_1656,N_19890,N_19998);
nand UO_1657 (O_1657,N_19853,N_19916);
nor UO_1658 (O_1658,N_19904,N_19970);
and UO_1659 (O_1659,N_19852,N_19926);
or UO_1660 (O_1660,N_19909,N_19856);
and UO_1661 (O_1661,N_19905,N_19957);
or UO_1662 (O_1662,N_19907,N_19935);
xor UO_1663 (O_1663,N_19972,N_19863);
nor UO_1664 (O_1664,N_19947,N_19853);
xnor UO_1665 (O_1665,N_19886,N_19942);
xor UO_1666 (O_1666,N_19978,N_19861);
xor UO_1667 (O_1667,N_19857,N_19865);
xnor UO_1668 (O_1668,N_19929,N_19997);
or UO_1669 (O_1669,N_19921,N_19903);
xnor UO_1670 (O_1670,N_19874,N_19925);
and UO_1671 (O_1671,N_19976,N_19949);
nor UO_1672 (O_1672,N_19999,N_19998);
or UO_1673 (O_1673,N_19977,N_19903);
nor UO_1674 (O_1674,N_19857,N_19932);
or UO_1675 (O_1675,N_19882,N_19890);
or UO_1676 (O_1676,N_19863,N_19966);
or UO_1677 (O_1677,N_19881,N_19985);
and UO_1678 (O_1678,N_19928,N_19866);
nor UO_1679 (O_1679,N_19998,N_19915);
nor UO_1680 (O_1680,N_19867,N_19882);
xnor UO_1681 (O_1681,N_19900,N_19924);
nand UO_1682 (O_1682,N_19939,N_19995);
nor UO_1683 (O_1683,N_19863,N_19919);
or UO_1684 (O_1684,N_19905,N_19907);
xor UO_1685 (O_1685,N_19917,N_19899);
xnor UO_1686 (O_1686,N_19915,N_19923);
nor UO_1687 (O_1687,N_19928,N_19929);
or UO_1688 (O_1688,N_19999,N_19848);
nand UO_1689 (O_1689,N_19959,N_19906);
xnor UO_1690 (O_1690,N_19895,N_19945);
xor UO_1691 (O_1691,N_19962,N_19906);
nor UO_1692 (O_1692,N_19852,N_19898);
xnor UO_1693 (O_1693,N_19921,N_19851);
and UO_1694 (O_1694,N_19916,N_19872);
xnor UO_1695 (O_1695,N_19874,N_19935);
nor UO_1696 (O_1696,N_19863,N_19961);
or UO_1697 (O_1697,N_19870,N_19895);
xor UO_1698 (O_1698,N_19929,N_19902);
nand UO_1699 (O_1699,N_19857,N_19868);
xnor UO_1700 (O_1700,N_19980,N_19903);
and UO_1701 (O_1701,N_19953,N_19996);
or UO_1702 (O_1702,N_19876,N_19847);
nand UO_1703 (O_1703,N_19850,N_19959);
xnor UO_1704 (O_1704,N_19985,N_19924);
nor UO_1705 (O_1705,N_19923,N_19957);
and UO_1706 (O_1706,N_19921,N_19864);
and UO_1707 (O_1707,N_19874,N_19855);
xnor UO_1708 (O_1708,N_19907,N_19867);
nor UO_1709 (O_1709,N_19961,N_19986);
and UO_1710 (O_1710,N_19912,N_19883);
and UO_1711 (O_1711,N_19842,N_19998);
and UO_1712 (O_1712,N_19885,N_19945);
xor UO_1713 (O_1713,N_19951,N_19905);
xnor UO_1714 (O_1714,N_19927,N_19942);
nor UO_1715 (O_1715,N_19851,N_19945);
nor UO_1716 (O_1716,N_19845,N_19840);
xor UO_1717 (O_1717,N_19954,N_19980);
nand UO_1718 (O_1718,N_19972,N_19909);
nor UO_1719 (O_1719,N_19987,N_19934);
nor UO_1720 (O_1720,N_19985,N_19891);
nand UO_1721 (O_1721,N_19846,N_19943);
xor UO_1722 (O_1722,N_19918,N_19948);
and UO_1723 (O_1723,N_19900,N_19840);
xnor UO_1724 (O_1724,N_19975,N_19979);
and UO_1725 (O_1725,N_19869,N_19995);
and UO_1726 (O_1726,N_19898,N_19858);
and UO_1727 (O_1727,N_19887,N_19919);
or UO_1728 (O_1728,N_19844,N_19851);
or UO_1729 (O_1729,N_19876,N_19974);
and UO_1730 (O_1730,N_19875,N_19863);
xor UO_1731 (O_1731,N_19918,N_19859);
nor UO_1732 (O_1732,N_19955,N_19964);
or UO_1733 (O_1733,N_19934,N_19938);
xnor UO_1734 (O_1734,N_19871,N_19978);
nand UO_1735 (O_1735,N_19883,N_19960);
nand UO_1736 (O_1736,N_19995,N_19913);
xor UO_1737 (O_1737,N_19911,N_19864);
xor UO_1738 (O_1738,N_19900,N_19984);
nor UO_1739 (O_1739,N_19982,N_19912);
xnor UO_1740 (O_1740,N_19938,N_19866);
or UO_1741 (O_1741,N_19872,N_19869);
nand UO_1742 (O_1742,N_19987,N_19948);
xor UO_1743 (O_1743,N_19922,N_19967);
or UO_1744 (O_1744,N_19894,N_19904);
xor UO_1745 (O_1745,N_19931,N_19900);
xnor UO_1746 (O_1746,N_19968,N_19895);
and UO_1747 (O_1747,N_19846,N_19948);
nand UO_1748 (O_1748,N_19990,N_19956);
nor UO_1749 (O_1749,N_19944,N_19938);
xnor UO_1750 (O_1750,N_19945,N_19848);
and UO_1751 (O_1751,N_19925,N_19872);
nand UO_1752 (O_1752,N_19988,N_19921);
nand UO_1753 (O_1753,N_19945,N_19976);
or UO_1754 (O_1754,N_19934,N_19907);
nor UO_1755 (O_1755,N_19859,N_19841);
nor UO_1756 (O_1756,N_19945,N_19930);
or UO_1757 (O_1757,N_19889,N_19846);
nand UO_1758 (O_1758,N_19945,N_19993);
nand UO_1759 (O_1759,N_19897,N_19975);
xor UO_1760 (O_1760,N_19956,N_19988);
or UO_1761 (O_1761,N_19912,N_19925);
nand UO_1762 (O_1762,N_19987,N_19875);
nor UO_1763 (O_1763,N_19874,N_19857);
or UO_1764 (O_1764,N_19914,N_19852);
or UO_1765 (O_1765,N_19997,N_19941);
or UO_1766 (O_1766,N_19992,N_19984);
nor UO_1767 (O_1767,N_19886,N_19977);
nand UO_1768 (O_1768,N_19941,N_19912);
and UO_1769 (O_1769,N_19848,N_19891);
nor UO_1770 (O_1770,N_19913,N_19862);
nand UO_1771 (O_1771,N_19850,N_19855);
nor UO_1772 (O_1772,N_19998,N_19973);
nor UO_1773 (O_1773,N_19923,N_19847);
and UO_1774 (O_1774,N_19878,N_19919);
and UO_1775 (O_1775,N_19852,N_19944);
nor UO_1776 (O_1776,N_19902,N_19840);
and UO_1777 (O_1777,N_19927,N_19840);
nor UO_1778 (O_1778,N_19874,N_19945);
xnor UO_1779 (O_1779,N_19965,N_19895);
nand UO_1780 (O_1780,N_19992,N_19980);
nor UO_1781 (O_1781,N_19993,N_19965);
nand UO_1782 (O_1782,N_19864,N_19969);
and UO_1783 (O_1783,N_19897,N_19995);
nand UO_1784 (O_1784,N_19887,N_19869);
nor UO_1785 (O_1785,N_19867,N_19950);
and UO_1786 (O_1786,N_19881,N_19871);
or UO_1787 (O_1787,N_19857,N_19929);
or UO_1788 (O_1788,N_19982,N_19981);
nand UO_1789 (O_1789,N_19975,N_19903);
or UO_1790 (O_1790,N_19896,N_19880);
or UO_1791 (O_1791,N_19889,N_19874);
nand UO_1792 (O_1792,N_19979,N_19845);
nand UO_1793 (O_1793,N_19958,N_19859);
nor UO_1794 (O_1794,N_19994,N_19847);
or UO_1795 (O_1795,N_19935,N_19895);
nor UO_1796 (O_1796,N_19910,N_19951);
and UO_1797 (O_1797,N_19930,N_19903);
and UO_1798 (O_1798,N_19886,N_19874);
nor UO_1799 (O_1799,N_19940,N_19886);
and UO_1800 (O_1800,N_19988,N_19939);
or UO_1801 (O_1801,N_19858,N_19895);
and UO_1802 (O_1802,N_19860,N_19962);
or UO_1803 (O_1803,N_19993,N_19981);
nor UO_1804 (O_1804,N_19908,N_19956);
or UO_1805 (O_1805,N_19929,N_19980);
nor UO_1806 (O_1806,N_19866,N_19940);
nand UO_1807 (O_1807,N_19903,N_19949);
and UO_1808 (O_1808,N_19953,N_19999);
and UO_1809 (O_1809,N_19853,N_19890);
or UO_1810 (O_1810,N_19924,N_19994);
and UO_1811 (O_1811,N_19890,N_19965);
xnor UO_1812 (O_1812,N_19893,N_19853);
and UO_1813 (O_1813,N_19865,N_19905);
and UO_1814 (O_1814,N_19888,N_19896);
nand UO_1815 (O_1815,N_19882,N_19891);
nand UO_1816 (O_1816,N_19927,N_19842);
and UO_1817 (O_1817,N_19847,N_19881);
nor UO_1818 (O_1818,N_19898,N_19996);
xor UO_1819 (O_1819,N_19997,N_19848);
and UO_1820 (O_1820,N_19900,N_19843);
or UO_1821 (O_1821,N_19899,N_19855);
nand UO_1822 (O_1822,N_19880,N_19905);
nand UO_1823 (O_1823,N_19955,N_19889);
and UO_1824 (O_1824,N_19876,N_19958);
or UO_1825 (O_1825,N_19933,N_19851);
nor UO_1826 (O_1826,N_19899,N_19882);
nor UO_1827 (O_1827,N_19896,N_19994);
nor UO_1828 (O_1828,N_19915,N_19996);
and UO_1829 (O_1829,N_19943,N_19973);
nor UO_1830 (O_1830,N_19951,N_19909);
or UO_1831 (O_1831,N_19938,N_19915);
xnor UO_1832 (O_1832,N_19859,N_19858);
and UO_1833 (O_1833,N_19930,N_19849);
nor UO_1834 (O_1834,N_19934,N_19864);
nand UO_1835 (O_1835,N_19897,N_19847);
xor UO_1836 (O_1836,N_19867,N_19915);
nand UO_1837 (O_1837,N_19981,N_19945);
nand UO_1838 (O_1838,N_19862,N_19907);
or UO_1839 (O_1839,N_19958,N_19860);
nor UO_1840 (O_1840,N_19891,N_19991);
and UO_1841 (O_1841,N_19992,N_19845);
nor UO_1842 (O_1842,N_19985,N_19938);
nor UO_1843 (O_1843,N_19849,N_19981);
and UO_1844 (O_1844,N_19845,N_19920);
and UO_1845 (O_1845,N_19891,N_19948);
and UO_1846 (O_1846,N_19858,N_19964);
nand UO_1847 (O_1847,N_19991,N_19976);
or UO_1848 (O_1848,N_19933,N_19866);
xor UO_1849 (O_1849,N_19961,N_19900);
or UO_1850 (O_1850,N_19904,N_19986);
xnor UO_1851 (O_1851,N_19905,N_19894);
and UO_1852 (O_1852,N_19933,N_19941);
xor UO_1853 (O_1853,N_19900,N_19901);
xor UO_1854 (O_1854,N_19871,N_19962);
or UO_1855 (O_1855,N_19945,N_19903);
nor UO_1856 (O_1856,N_19975,N_19914);
nand UO_1857 (O_1857,N_19949,N_19853);
nor UO_1858 (O_1858,N_19922,N_19927);
and UO_1859 (O_1859,N_19933,N_19938);
nor UO_1860 (O_1860,N_19844,N_19953);
xor UO_1861 (O_1861,N_19985,N_19928);
xor UO_1862 (O_1862,N_19936,N_19994);
and UO_1863 (O_1863,N_19880,N_19961);
nand UO_1864 (O_1864,N_19967,N_19944);
and UO_1865 (O_1865,N_19877,N_19905);
xor UO_1866 (O_1866,N_19852,N_19876);
and UO_1867 (O_1867,N_19913,N_19850);
nand UO_1868 (O_1868,N_19858,N_19883);
or UO_1869 (O_1869,N_19938,N_19895);
xnor UO_1870 (O_1870,N_19943,N_19963);
or UO_1871 (O_1871,N_19879,N_19893);
or UO_1872 (O_1872,N_19968,N_19936);
and UO_1873 (O_1873,N_19911,N_19902);
nand UO_1874 (O_1874,N_19859,N_19917);
or UO_1875 (O_1875,N_19955,N_19903);
nand UO_1876 (O_1876,N_19892,N_19859);
and UO_1877 (O_1877,N_19946,N_19979);
nand UO_1878 (O_1878,N_19851,N_19958);
xor UO_1879 (O_1879,N_19945,N_19915);
xor UO_1880 (O_1880,N_19934,N_19937);
nor UO_1881 (O_1881,N_19849,N_19990);
nand UO_1882 (O_1882,N_19974,N_19965);
nand UO_1883 (O_1883,N_19857,N_19886);
xnor UO_1884 (O_1884,N_19913,N_19861);
and UO_1885 (O_1885,N_19852,N_19993);
nand UO_1886 (O_1886,N_19880,N_19962);
or UO_1887 (O_1887,N_19903,N_19866);
nand UO_1888 (O_1888,N_19893,N_19943);
xor UO_1889 (O_1889,N_19921,N_19996);
and UO_1890 (O_1890,N_19861,N_19865);
and UO_1891 (O_1891,N_19866,N_19847);
or UO_1892 (O_1892,N_19881,N_19857);
xnor UO_1893 (O_1893,N_19969,N_19934);
xnor UO_1894 (O_1894,N_19875,N_19934);
and UO_1895 (O_1895,N_19956,N_19993);
nand UO_1896 (O_1896,N_19968,N_19840);
nor UO_1897 (O_1897,N_19978,N_19917);
nor UO_1898 (O_1898,N_19965,N_19968);
or UO_1899 (O_1899,N_19980,N_19933);
or UO_1900 (O_1900,N_19847,N_19860);
nor UO_1901 (O_1901,N_19934,N_19850);
nor UO_1902 (O_1902,N_19947,N_19983);
or UO_1903 (O_1903,N_19956,N_19895);
nor UO_1904 (O_1904,N_19873,N_19901);
xor UO_1905 (O_1905,N_19961,N_19975);
xor UO_1906 (O_1906,N_19884,N_19860);
and UO_1907 (O_1907,N_19925,N_19843);
xnor UO_1908 (O_1908,N_19920,N_19860);
xnor UO_1909 (O_1909,N_19841,N_19877);
xor UO_1910 (O_1910,N_19948,N_19901);
and UO_1911 (O_1911,N_19900,N_19852);
and UO_1912 (O_1912,N_19953,N_19933);
nand UO_1913 (O_1913,N_19970,N_19968);
xor UO_1914 (O_1914,N_19910,N_19938);
nor UO_1915 (O_1915,N_19931,N_19842);
xor UO_1916 (O_1916,N_19942,N_19919);
xor UO_1917 (O_1917,N_19864,N_19971);
nand UO_1918 (O_1918,N_19891,N_19898);
or UO_1919 (O_1919,N_19978,N_19873);
nand UO_1920 (O_1920,N_19952,N_19901);
nand UO_1921 (O_1921,N_19930,N_19935);
or UO_1922 (O_1922,N_19972,N_19923);
xor UO_1923 (O_1923,N_19993,N_19900);
nand UO_1924 (O_1924,N_19997,N_19842);
and UO_1925 (O_1925,N_19970,N_19926);
nor UO_1926 (O_1926,N_19872,N_19940);
xnor UO_1927 (O_1927,N_19847,N_19840);
xnor UO_1928 (O_1928,N_19858,N_19982);
and UO_1929 (O_1929,N_19876,N_19909);
and UO_1930 (O_1930,N_19865,N_19976);
xor UO_1931 (O_1931,N_19934,N_19964);
xor UO_1932 (O_1932,N_19857,N_19998);
or UO_1933 (O_1933,N_19988,N_19863);
nor UO_1934 (O_1934,N_19884,N_19971);
nand UO_1935 (O_1935,N_19989,N_19857);
or UO_1936 (O_1936,N_19897,N_19987);
xnor UO_1937 (O_1937,N_19862,N_19920);
xor UO_1938 (O_1938,N_19922,N_19876);
nor UO_1939 (O_1939,N_19883,N_19900);
nor UO_1940 (O_1940,N_19936,N_19922);
nand UO_1941 (O_1941,N_19958,N_19923);
nand UO_1942 (O_1942,N_19864,N_19983);
and UO_1943 (O_1943,N_19913,N_19956);
xnor UO_1944 (O_1944,N_19846,N_19978);
and UO_1945 (O_1945,N_19847,N_19959);
xnor UO_1946 (O_1946,N_19923,N_19959);
xor UO_1947 (O_1947,N_19882,N_19969);
nand UO_1948 (O_1948,N_19895,N_19857);
nor UO_1949 (O_1949,N_19984,N_19851);
xor UO_1950 (O_1950,N_19882,N_19916);
nor UO_1951 (O_1951,N_19993,N_19941);
nor UO_1952 (O_1952,N_19961,N_19913);
or UO_1953 (O_1953,N_19966,N_19855);
and UO_1954 (O_1954,N_19917,N_19882);
nand UO_1955 (O_1955,N_19999,N_19873);
or UO_1956 (O_1956,N_19966,N_19953);
and UO_1957 (O_1957,N_19896,N_19928);
nand UO_1958 (O_1958,N_19971,N_19899);
nand UO_1959 (O_1959,N_19880,N_19972);
and UO_1960 (O_1960,N_19854,N_19841);
xnor UO_1961 (O_1961,N_19895,N_19990);
nor UO_1962 (O_1962,N_19902,N_19914);
and UO_1963 (O_1963,N_19999,N_19870);
and UO_1964 (O_1964,N_19890,N_19850);
xor UO_1965 (O_1965,N_19890,N_19906);
nand UO_1966 (O_1966,N_19993,N_19924);
and UO_1967 (O_1967,N_19900,N_19945);
xnor UO_1968 (O_1968,N_19923,N_19884);
and UO_1969 (O_1969,N_19932,N_19916);
xnor UO_1970 (O_1970,N_19880,N_19912);
or UO_1971 (O_1971,N_19930,N_19877);
xor UO_1972 (O_1972,N_19954,N_19904);
or UO_1973 (O_1973,N_19976,N_19911);
or UO_1974 (O_1974,N_19967,N_19964);
and UO_1975 (O_1975,N_19840,N_19956);
and UO_1976 (O_1976,N_19980,N_19907);
nand UO_1977 (O_1977,N_19977,N_19992);
or UO_1978 (O_1978,N_19992,N_19880);
and UO_1979 (O_1979,N_19874,N_19974);
xor UO_1980 (O_1980,N_19960,N_19954);
or UO_1981 (O_1981,N_19988,N_19984);
and UO_1982 (O_1982,N_19937,N_19847);
nor UO_1983 (O_1983,N_19887,N_19850);
and UO_1984 (O_1984,N_19917,N_19884);
and UO_1985 (O_1985,N_19859,N_19876);
nor UO_1986 (O_1986,N_19862,N_19949);
and UO_1987 (O_1987,N_19857,N_19846);
nor UO_1988 (O_1988,N_19857,N_19978);
xnor UO_1989 (O_1989,N_19917,N_19845);
or UO_1990 (O_1990,N_19939,N_19884);
nor UO_1991 (O_1991,N_19995,N_19960);
nand UO_1992 (O_1992,N_19960,N_19935);
nor UO_1993 (O_1993,N_19949,N_19910);
nor UO_1994 (O_1994,N_19869,N_19954);
nand UO_1995 (O_1995,N_19999,N_19985);
and UO_1996 (O_1996,N_19851,N_19915);
or UO_1997 (O_1997,N_19872,N_19847);
xnor UO_1998 (O_1998,N_19909,N_19894);
nand UO_1999 (O_1999,N_19938,N_19975);
nand UO_2000 (O_2000,N_19862,N_19974);
nand UO_2001 (O_2001,N_19885,N_19918);
or UO_2002 (O_2002,N_19886,N_19984);
or UO_2003 (O_2003,N_19892,N_19847);
xnor UO_2004 (O_2004,N_19853,N_19928);
and UO_2005 (O_2005,N_19989,N_19993);
or UO_2006 (O_2006,N_19889,N_19902);
and UO_2007 (O_2007,N_19999,N_19964);
nor UO_2008 (O_2008,N_19956,N_19914);
xnor UO_2009 (O_2009,N_19963,N_19910);
or UO_2010 (O_2010,N_19944,N_19992);
and UO_2011 (O_2011,N_19908,N_19989);
or UO_2012 (O_2012,N_19936,N_19955);
nand UO_2013 (O_2013,N_19883,N_19921);
nand UO_2014 (O_2014,N_19889,N_19859);
nand UO_2015 (O_2015,N_19891,N_19925);
nand UO_2016 (O_2016,N_19883,N_19930);
or UO_2017 (O_2017,N_19918,N_19987);
nand UO_2018 (O_2018,N_19865,N_19924);
nor UO_2019 (O_2019,N_19902,N_19953);
nand UO_2020 (O_2020,N_19991,N_19896);
xnor UO_2021 (O_2021,N_19992,N_19941);
or UO_2022 (O_2022,N_19933,N_19912);
xor UO_2023 (O_2023,N_19966,N_19915);
nand UO_2024 (O_2024,N_19868,N_19845);
nand UO_2025 (O_2025,N_19910,N_19962);
and UO_2026 (O_2026,N_19903,N_19976);
xor UO_2027 (O_2027,N_19843,N_19863);
nand UO_2028 (O_2028,N_19900,N_19971);
xnor UO_2029 (O_2029,N_19965,N_19944);
xnor UO_2030 (O_2030,N_19942,N_19999);
nand UO_2031 (O_2031,N_19994,N_19859);
and UO_2032 (O_2032,N_19952,N_19876);
and UO_2033 (O_2033,N_19990,N_19972);
and UO_2034 (O_2034,N_19989,N_19959);
xor UO_2035 (O_2035,N_19975,N_19992);
xnor UO_2036 (O_2036,N_19899,N_19852);
and UO_2037 (O_2037,N_19862,N_19935);
and UO_2038 (O_2038,N_19840,N_19996);
xor UO_2039 (O_2039,N_19877,N_19979);
xnor UO_2040 (O_2040,N_19992,N_19930);
nor UO_2041 (O_2041,N_19915,N_19956);
xor UO_2042 (O_2042,N_19954,N_19850);
nand UO_2043 (O_2043,N_19958,N_19951);
nor UO_2044 (O_2044,N_19894,N_19927);
nor UO_2045 (O_2045,N_19942,N_19931);
nand UO_2046 (O_2046,N_19958,N_19957);
xnor UO_2047 (O_2047,N_19852,N_19939);
xor UO_2048 (O_2048,N_19932,N_19986);
or UO_2049 (O_2049,N_19909,N_19919);
xor UO_2050 (O_2050,N_19939,N_19921);
or UO_2051 (O_2051,N_19907,N_19892);
or UO_2052 (O_2052,N_19894,N_19847);
nor UO_2053 (O_2053,N_19913,N_19901);
or UO_2054 (O_2054,N_19853,N_19844);
or UO_2055 (O_2055,N_19990,N_19926);
nor UO_2056 (O_2056,N_19943,N_19850);
nor UO_2057 (O_2057,N_19998,N_19914);
or UO_2058 (O_2058,N_19887,N_19872);
xnor UO_2059 (O_2059,N_19884,N_19956);
xor UO_2060 (O_2060,N_19843,N_19940);
or UO_2061 (O_2061,N_19842,N_19930);
nand UO_2062 (O_2062,N_19940,N_19988);
nor UO_2063 (O_2063,N_19846,N_19852);
nand UO_2064 (O_2064,N_19988,N_19922);
nand UO_2065 (O_2065,N_19889,N_19918);
and UO_2066 (O_2066,N_19977,N_19995);
and UO_2067 (O_2067,N_19900,N_19847);
nor UO_2068 (O_2068,N_19949,N_19944);
nor UO_2069 (O_2069,N_19866,N_19845);
xnor UO_2070 (O_2070,N_19840,N_19985);
nor UO_2071 (O_2071,N_19876,N_19887);
and UO_2072 (O_2072,N_19962,N_19943);
nor UO_2073 (O_2073,N_19959,N_19964);
nor UO_2074 (O_2074,N_19987,N_19843);
or UO_2075 (O_2075,N_19860,N_19944);
nor UO_2076 (O_2076,N_19878,N_19893);
nor UO_2077 (O_2077,N_19960,N_19912);
xor UO_2078 (O_2078,N_19864,N_19903);
nand UO_2079 (O_2079,N_19893,N_19958);
and UO_2080 (O_2080,N_19872,N_19873);
nand UO_2081 (O_2081,N_19936,N_19943);
nor UO_2082 (O_2082,N_19848,N_19905);
or UO_2083 (O_2083,N_19920,N_19879);
and UO_2084 (O_2084,N_19962,N_19913);
or UO_2085 (O_2085,N_19887,N_19939);
nand UO_2086 (O_2086,N_19893,N_19944);
nor UO_2087 (O_2087,N_19889,N_19858);
nand UO_2088 (O_2088,N_19896,N_19884);
or UO_2089 (O_2089,N_19871,N_19893);
nand UO_2090 (O_2090,N_19853,N_19996);
nor UO_2091 (O_2091,N_19970,N_19874);
xnor UO_2092 (O_2092,N_19933,N_19853);
nor UO_2093 (O_2093,N_19903,N_19968);
or UO_2094 (O_2094,N_19960,N_19860);
or UO_2095 (O_2095,N_19914,N_19955);
nor UO_2096 (O_2096,N_19894,N_19971);
and UO_2097 (O_2097,N_19840,N_19932);
nor UO_2098 (O_2098,N_19904,N_19901);
or UO_2099 (O_2099,N_19998,N_19958);
xor UO_2100 (O_2100,N_19886,N_19955);
nor UO_2101 (O_2101,N_19922,N_19878);
nand UO_2102 (O_2102,N_19919,N_19920);
or UO_2103 (O_2103,N_19947,N_19991);
nor UO_2104 (O_2104,N_19955,N_19994);
or UO_2105 (O_2105,N_19898,N_19971);
nand UO_2106 (O_2106,N_19919,N_19987);
nand UO_2107 (O_2107,N_19986,N_19860);
xnor UO_2108 (O_2108,N_19983,N_19911);
and UO_2109 (O_2109,N_19931,N_19846);
nor UO_2110 (O_2110,N_19959,N_19863);
nor UO_2111 (O_2111,N_19952,N_19912);
nor UO_2112 (O_2112,N_19952,N_19997);
and UO_2113 (O_2113,N_19841,N_19913);
xnor UO_2114 (O_2114,N_19996,N_19902);
nor UO_2115 (O_2115,N_19886,N_19926);
or UO_2116 (O_2116,N_19961,N_19906);
xor UO_2117 (O_2117,N_19980,N_19976);
or UO_2118 (O_2118,N_19991,N_19841);
nor UO_2119 (O_2119,N_19874,N_19893);
nand UO_2120 (O_2120,N_19875,N_19951);
xnor UO_2121 (O_2121,N_19955,N_19949);
nor UO_2122 (O_2122,N_19938,N_19874);
nand UO_2123 (O_2123,N_19908,N_19940);
nand UO_2124 (O_2124,N_19972,N_19874);
or UO_2125 (O_2125,N_19922,N_19914);
and UO_2126 (O_2126,N_19881,N_19851);
nor UO_2127 (O_2127,N_19914,N_19952);
nand UO_2128 (O_2128,N_19950,N_19908);
and UO_2129 (O_2129,N_19918,N_19913);
and UO_2130 (O_2130,N_19941,N_19974);
or UO_2131 (O_2131,N_19970,N_19957);
xor UO_2132 (O_2132,N_19910,N_19925);
nand UO_2133 (O_2133,N_19931,N_19996);
and UO_2134 (O_2134,N_19894,N_19947);
nor UO_2135 (O_2135,N_19900,N_19958);
nand UO_2136 (O_2136,N_19858,N_19844);
nor UO_2137 (O_2137,N_19882,N_19967);
nand UO_2138 (O_2138,N_19976,N_19918);
nand UO_2139 (O_2139,N_19979,N_19968);
or UO_2140 (O_2140,N_19904,N_19849);
or UO_2141 (O_2141,N_19916,N_19986);
nor UO_2142 (O_2142,N_19861,N_19866);
nor UO_2143 (O_2143,N_19891,N_19986);
xnor UO_2144 (O_2144,N_19931,N_19863);
xor UO_2145 (O_2145,N_19854,N_19892);
nand UO_2146 (O_2146,N_19954,N_19922);
xor UO_2147 (O_2147,N_19929,N_19996);
nor UO_2148 (O_2148,N_19969,N_19904);
and UO_2149 (O_2149,N_19942,N_19916);
nor UO_2150 (O_2150,N_19940,N_19877);
nand UO_2151 (O_2151,N_19996,N_19965);
and UO_2152 (O_2152,N_19999,N_19883);
nand UO_2153 (O_2153,N_19926,N_19933);
nor UO_2154 (O_2154,N_19966,N_19954);
and UO_2155 (O_2155,N_19980,N_19936);
nor UO_2156 (O_2156,N_19981,N_19959);
or UO_2157 (O_2157,N_19989,N_19988);
and UO_2158 (O_2158,N_19976,N_19973);
nor UO_2159 (O_2159,N_19845,N_19998);
and UO_2160 (O_2160,N_19990,N_19868);
nor UO_2161 (O_2161,N_19861,N_19938);
and UO_2162 (O_2162,N_19845,N_19874);
and UO_2163 (O_2163,N_19882,N_19997);
nand UO_2164 (O_2164,N_19917,N_19842);
or UO_2165 (O_2165,N_19876,N_19924);
nand UO_2166 (O_2166,N_19895,N_19980);
nand UO_2167 (O_2167,N_19973,N_19939);
or UO_2168 (O_2168,N_19915,N_19877);
nand UO_2169 (O_2169,N_19933,N_19931);
xor UO_2170 (O_2170,N_19931,N_19956);
xnor UO_2171 (O_2171,N_19942,N_19937);
nand UO_2172 (O_2172,N_19977,N_19928);
nand UO_2173 (O_2173,N_19949,N_19917);
nand UO_2174 (O_2174,N_19875,N_19872);
and UO_2175 (O_2175,N_19876,N_19962);
and UO_2176 (O_2176,N_19862,N_19890);
and UO_2177 (O_2177,N_19982,N_19965);
nor UO_2178 (O_2178,N_19961,N_19999);
xnor UO_2179 (O_2179,N_19852,N_19974);
nand UO_2180 (O_2180,N_19861,N_19987);
nand UO_2181 (O_2181,N_19873,N_19874);
or UO_2182 (O_2182,N_19995,N_19968);
nand UO_2183 (O_2183,N_19889,N_19986);
nand UO_2184 (O_2184,N_19967,N_19969);
xnor UO_2185 (O_2185,N_19952,N_19855);
nor UO_2186 (O_2186,N_19891,N_19908);
xor UO_2187 (O_2187,N_19957,N_19857);
and UO_2188 (O_2188,N_19950,N_19958);
or UO_2189 (O_2189,N_19993,N_19907);
nor UO_2190 (O_2190,N_19857,N_19946);
and UO_2191 (O_2191,N_19877,N_19880);
xor UO_2192 (O_2192,N_19890,N_19991);
or UO_2193 (O_2193,N_19888,N_19939);
nand UO_2194 (O_2194,N_19847,N_19898);
or UO_2195 (O_2195,N_19890,N_19985);
xnor UO_2196 (O_2196,N_19853,N_19950);
nand UO_2197 (O_2197,N_19844,N_19913);
nand UO_2198 (O_2198,N_19862,N_19939);
or UO_2199 (O_2199,N_19940,N_19911);
nor UO_2200 (O_2200,N_19876,N_19955);
and UO_2201 (O_2201,N_19909,N_19929);
xnor UO_2202 (O_2202,N_19882,N_19941);
or UO_2203 (O_2203,N_19986,N_19963);
nor UO_2204 (O_2204,N_19911,N_19872);
and UO_2205 (O_2205,N_19932,N_19956);
or UO_2206 (O_2206,N_19911,N_19868);
or UO_2207 (O_2207,N_19950,N_19884);
nor UO_2208 (O_2208,N_19956,N_19952);
nor UO_2209 (O_2209,N_19991,N_19970);
or UO_2210 (O_2210,N_19939,N_19919);
and UO_2211 (O_2211,N_19895,N_19914);
and UO_2212 (O_2212,N_19862,N_19934);
nand UO_2213 (O_2213,N_19895,N_19932);
nor UO_2214 (O_2214,N_19895,N_19841);
nand UO_2215 (O_2215,N_19950,N_19943);
nand UO_2216 (O_2216,N_19967,N_19956);
and UO_2217 (O_2217,N_19968,N_19841);
and UO_2218 (O_2218,N_19854,N_19901);
xnor UO_2219 (O_2219,N_19958,N_19852);
and UO_2220 (O_2220,N_19916,N_19912);
nor UO_2221 (O_2221,N_19884,N_19866);
xnor UO_2222 (O_2222,N_19937,N_19855);
nand UO_2223 (O_2223,N_19854,N_19996);
and UO_2224 (O_2224,N_19926,N_19998);
nand UO_2225 (O_2225,N_19915,N_19888);
nand UO_2226 (O_2226,N_19989,N_19928);
nand UO_2227 (O_2227,N_19908,N_19964);
nor UO_2228 (O_2228,N_19855,N_19935);
nand UO_2229 (O_2229,N_19873,N_19941);
nor UO_2230 (O_2230,N_19947,N_19996);
nand UO_2231 (O_2231,N_19962,N_19957);
and UO_2232 (O_2232,N_19849,N_19883);
or UO_2233 (O_2233,N_19929,N_19951);
nor UO_2234 (O_2234,N_19872,N_19904);
nor UO_2235 (O_2235,N_19866,N_19841);
and UO_2236 (O_2236,N_19993,N_19970);
and UO_2237 (O_2237,N_19909,N_19869);
and UO_2238 (O_2238,N_19975,N_19991);
nand UO_2239 (O_2239,N_19845,N_19971);
xnor UO_2240 (O_2240,N_19844,N_19849);
and UO_2241 (O_2241,N_19996,N_19857);
and UO_2242 (O_2242,N_19929,N_19956);
or UO_2243 (O_2243,N_19895,N_19896);
xor UO_2244 (O_2244,N_19912,N_19864);
and UO_2245 (O_2245,N_19986,N_19912);
xnor UO_2246 (O_2246,N_19981,N_19910);
and UO_2247 (O_2247,N_19996,N_19977);
or UO_2248 (O_2248,N_19910,N_19955);
nor UO_2249 (O_2249,N_19974,N_19954);
nor UO_2250 (O_2250,N_19858,N_19904);
nor UO_2251 (O_2251,N_19891,N_19968);
and UO_2252 (O_2252,N_19868,N_19844);
and UO_2253 (O_2253,N_19877,N_19888);
nor UO_2254 (O_2254,N_19931,N_19960);
and UO_2255 (O_2255,N_19846,N_19968);
nand UO_2256 (O_2256,N_19911,N_19875);
nor UO_2257 (O_2257,N_19901,N_19892);
xnor UO_2258 (O_2258,N_19971,N_19882);
or UO_2259 (O_2259,N_19943,N_19980);
xor UO_2260 (O_2260,N_19950,N_19941);
or UO_2261 (O_2261,N_19919,N_19888);
nand UO_2262 (O_2262,N_19966,N_19914);
or UO_2263 (O_2263,N_19981,N_19917);
nor UO_2264 (O_2264,N_19936,N_19933);
xor UO_2265 (O_2265,N_19938,N_19930);
nand UO_2266 (O_2266,N_19958,N_19844);
nand UO_2267 (O_2267,N_19842,N_19982);
and UO_2268 (O_2268,N_19977,N_19853);
nor UO_2269 (O_2269,N_19909,N_19969);
xor UO_2270 (O_2270,N_19960,N_19902);
and UO_2271 (O_2271,N_19895,N_19876);
and UO_2272 (O_2272,N_19898,N_19992);
nor UO_2273 (O_2273,N_19857,N_19908);
and UO_2274 (O_2274,N_19972,N_19884);
xnor UO_2275 (O_2275,N_19845,N_19942);
nand UO_2276 (O_2276,N_19961,N_19848);
or UO_2277 (O_2277,N_19953,N_19859);
xnor UO_2278 (O_2278,N_19970,N_19908);
nor UO_2279 (O_2279,N_19925,N_19897);
xor UO_2280 (O_2280,N_19946,N_19887);
nand UO_2281 (O_2281,N_19905,N_19862);
nor UO_2282 (O_2282,N_19946,N_19967);
nand UO_2283 (O_2283,N_19954,N_19907);
and UO_2284 (O_2284,N_19917,N_19995);
and UO_2285 (O_2285,N_19943,N_19867);
nand UO_2286 (O_2286,N_19928,N_19923);
nor UO_2287 (O_2287,N_19974,N_19842);
or UO_2288 (O_2288,N_19952,N_19927);
xnor UO_2289 (O_2289,N_19857,N_19851);
or UO_2290 (O_2290,N_19962,N_19967);
nand UO_2291 (O_2291,N_19960,N_19976);
nor UO_2292 (O_2292,N_19953,N_19841);
and UO_2293 (O_2293,N_19924,N_19995);
xnor UO_2294 (O_2294,N_19894,N_19901);
and UO_2295 (O_2295,N_19869,N_19974);
nor UO_2296 (O_2296,N_19935,N_19932);
xor UO_2297 (O_2297,N_19867,N_19976);
nor UO_2298 (O_2298,N_19885,N_19929);
nand UO_2299 (O_2299,N_19952,N_19882);
nor UO_2300 (O_2300,N_19953,N_19918);
and UO_2301 (O_2301,N_19993,N_19915);
nand UO_2302 (O_2302,N_19996,N_19980);
and UO_2303 (O_2303,N_19871,N_19941);
nor UO_2304 (O_2304,N_19914,N_19875);
or UO_2305 (O_2305,N_19981,N_19951);
or UO_2306 (O_2306,N_19859,N_19974);
and UO_2307 (O_2307,N_19865,N_19933);
nor UO_2308 (O_2308,N_19934,N_19897);
nand UO_2309 (O_2309,N_19859,N_19929);
nor UO_2310 (O_2310,N_19892,N_19942);
and UO_2311 (O_2311,N_19859,N_19970);
nor UO_2312 (O_2312,N_19912,N_19899);
and UO_2313 (O_2313,N_19840,N_19872);
nand UO_2314 (O_2314,N_19856,N_19861);
nand UO_2315 (O_2315,N_19930,N_19932);
nand UO_2316 (O_2316,N_19843,N_19936);
xnor UO_2317 (O_2317,N_19893,N_19970);
or UO_2318 (O_2318,N_19962,N_19912);
xnor UO_2319 (O_2319,N_19959,N_19916);
and UO_2320 (O_2320,N_19982,N_19983);
nor UO_2321 (O_2321,N_19968,N_19955);
xor UO_2322 (O_2322,N_19861,N_19891);
and UO_2323 (O_2323,N_19977,N_19937);
and UO_2324 (O_2324,N_19986,N_19934);
nand UO_2325 (O_2325,N_19898,N_19910);
xnor UO_2326 (O_2326,N_19927,N_19863);
nand UO_2327 (O_2327,N_19912,N_19841);
nand UO_2328 (O_2328,N_19978,N_19894);
or UO_2329 (O_2329,N_19898,N_19982);
or UO_2330 (O_2330,N_19995,N_19973);
or UO_2331 (O_2331,N_19929,N_19844);
or UO_2332 (O_2332,N_19880,N_19892);
xnor UO_2333 (O_2333,N_19888,N_19852);
and UO_2334 (O_2334,N_19849,N_19958);
nor UO_2335 (O_2335,N_19955,N_19870);
xnor UO_2336 (O_2336,N_19919,N_19877);
or UO_2337 (O_2337,N_19888,N_19884);
or UO_2338 (O_2338,N_19910,N_19997);
xor UO_2339 (O_2339,N_19965,N_19921);
or UO_2340 (O_2340,N_19971,N_19917);
xnor UO_2341 (O_2341,N_19972,N_19931);
and UO_2342 (O_2342,N_19914,N_19964);
nor UO_2343 (O_2343,N_19889,N_19974);
and UO_2344 (O_2344,N_19976,N_19927);
xnor UO_2345 (O_2345,N_19995,N_19876);
nand UO_2346 (O_2346,N_19921,N_19975);
xor UO_2347 (O_2347,N_19844,N_19984);
nand UO_2348 (O_2348,N_19880,N_19984);
nand UO_2349 (O_2349,N_19856,N_19947);
nand UO_2350 (O_2350,N_19909,N_19958);
nor UO_2351 (O_2351,N_19846,N_19923);
xnor UO_2352 (O_2352,N_19967,N_19951);
xor UO_2353 (O_2353,N_19979,N_19843);
or UO_2354 (O_2354,N_19913,N_19883);
or UO_2355 (O_2355,N_19919,N_19995);
xor UO_2356 (O_2356,N_19986,N_19962);
nor UO_2357 (O_2357,N_19892,N_19869);
nand UO_2358 (O_2358,N_19864,N_19957);
xor UO_2359 (O_2359,N_19958,N_19976);
nand UO_2360 (O_2360,N_19988,N_19976);
nor UO_2361 (O_2361,N_19902,N_19895);
xnor UO_2362 (O_2362,N_19873,N_19850);
nor UO_2363 (O_2363,N_19979,N_19872);
xor UO_2364 (O_2364,N_19953,N_19920);
or UO_2365 (O_2365,N_19939,N_19885);
xnor UO_2366 (O_2366,N_19873,N_19942);
nand UO_2367 (O_2367,N_19876,N_19886);
xor UO_2368 (O_2368,N_19850,N_19851);
nand UO_2369 (O_2369,N_19872,N_19997);
nor UO_2370 (O_2370,N_19870,N_19857);
xor UO_2371 (O_2371,N_19946,N_19991);
nand UO_2372 (O_2372,N_19876,N_19856);
nor UO_2373 (O_2373,N_19944,N_19979);
or UO_2374 (O_2374,N_19874,N_19923);
and UO_2375 (O_2375,N_19938,N_19992);
and UO_2376 (O_2376,N_19972,N_19980);
and UO_2377 (O_2377,N_19879,N_19915);
nor UO_2378 (O_2378,N_19933,N_19952);
and UO_2379 (O_2379,N_19962,N_19865);
xor UO_2380 (O_2380,N_19918,N_19945);
nand UO_2381 (O_2381,N_19875,N_19921);
or UO_2382 (O_2382,N_19983,N_19957);
nand UO_2383 (O_2383,N_19955,N_19864);
nand UO_2384 (O_2384,N_19876,N_19881);
and UO_2385 (O_2385,N_19966,N_19852);
xnor UO_2386 (O_2386,N_19904,N_19878);
nor UO_2387 (O_2387,N_19960,N_19970);
xnor UO_2388 (O_2388,N_19884,N_19842);
xor UO_2389 (O_2389,N_19948,N_19992);
or UO_2390 (O_2390,N_19954,N_19976);
xor UO_2391 (O_2391,N_19846,N_19960);
nand UO_2392 (O_2392,N_19887,N_19877);
or UO_2393 (O_2393,N_19910,N_19991);
nor UO_2394 (O_2394,N_19986,N_19935);
or UO_2395 (O_2395,N_19926,N_19931);
nor UO_2396 (O_2396,N_19905,N_19922);
or UO_2397 (O_2397,N_19913,N_19968);
or UO_2398 (O_2398,N_19974,N_19996);
nand UO_2399 (O_2399,N_19981,N_19875);
nand UO_2400 (O_2400,N_19887,N_19861);
and UO_2401 (O_2401,N_19944,N_19931);
xnor UO_2402 (O_2402,N_19995,N_19881);
nor UO_2403 (O_2403,N_19963,N_19927);
nand UO_2404 (O_2404,N_19900,N_19864);
and UO_2405 (O_2405,N_19923,N_19995);
or UO_2406 (O_2406,N_19878,N_19890);
and UO_2407 (O_2407,N_19934,N_19892);
nor UO_2408 (O_2408,N_19924,N_19844);
nor UO_2409 (O_2409,N_19841,N_19963);
nand UO_2410 (O_2410,N_19991,N_19862);
and UO_2411 (O_2411,N_19935,N_19890);
nor UO_2412 (O_2412,N_19850,N_19847);
nor UO_2413 (O_2413,N_19975,N_19971);
nor UO_2414 (O_2414,N_19862,N_19847);
nor UO_2415 (O_2415,N_19948,N_19998);
and UO_2416 (O_2416,N_19976,N_19842);
nor UO_2417 (O_2417,N_19858,N_19965);
nor UO_2418 (O_2418,N_19930,N_19865);
xor UO_2419 (O_2419,N_19945,N_19880);
nor UO_2420 (O_2420,N_19865,N_19875);
nand UO_2421 (O_2421,N_19964,N_19923);
nor UO_2422 (O_2422,N_19939,N_19994);
and UO_2423 (O_2423,N_19858,N_19975);
nand UO_2424 (O_2424,N_19939,N_19978);
xnor UO_2425 (O_2425,N_19985,N_19848);
or UO_2426 (O_2426,N_19856,N_19905);
nand UO_2427 (O_2427,N_19880,N_19993);
and UO_2428 (O_2428,N_19898,N_19867);
nor UO_2429 (O_2429,N_19912,N_19930);
nor UO_2430 (O_2430,N_19922,N_19892);
and UO_2431 (O_2431,N_19880,N_19946);
nor UO_2432 (O_2432,N_19980,N_19893);
xor UO_2433 (O_2433,N_19983,N_19909);
nand UO_2434 (O_2434,N_19902,N_19940);
xnor UO_2435 (O_2435,N_19889,N_19931);
nand UO_2436 (O_2436,N_19890,N_19977);
nand UO_2437 (O_2437,N_19998,N_19933);
or UO_2438 (O_2438,N_19996,N_19951);
nor UO_2439 (O_2439,N_19860,N_19899);
nor UO_2440 (O_2440,N_19963,N_19950);
nor UO_2441 (O_2441,N_19886,N_19909);
nor UO_2442 (O_2442,N_19919,N_19915);
or UO_2443 (O_2443,N_19987,N_19876);
or UO_2444 (O_2444,N_19972,N_19946);
and UO_2445 (O_2445,N_19966,N_19842);
nand UO_2446 (O_2446,N_19966,N_19995);
nor UO_2447 (O_2447,N_19911,N_19934);
xnor UO_2448 (O_2448,N_19890,N_19872);
nor UO_2449 (O_2449,N_19869,N_19854);
nand UO_2450 (O_2450,N_19925,N_19953);
xor UO_2451 (O_2451,N_19879,N_19917);
xor UO_2452 (O_2452,N_19929,N_19960);
nor UO_2453 (O_2453,N_19931,N_19856);
or UO_2454 (O_2454,N_19864,N_19878);
or UO_2455 (O_2455,N_19914,N_19990);
and UO_2456 (O_2456,N_19972,N_19879);
and UO_2457 (O_2457,N_19915,N_19843);
nand UO_2458 (O_2458,N_19921,N_19881);
xor UO_2459 (O_2459,N_19868,N_19954);
nor UO_2460 (O_2460,N_19877,N_19895);
or UO_2461 (O_2461,N_19893,N_19978);
or UO_2462 (O_2462,N_19878,N_19885);
or UO_2463 (O_2463,N_19921,N_19997);
nand UO_2464 (O_2464,N_19952,N_19967);
and UO_2465 (O_2465,N_19886,N_19890);
and UO_2466 (O_2466,N_19993,N_19906);
xor UO_2467 (O_2467,N_19998,N_19907);
xor UO_2468 (O_2468,N_19968,N_19975);
and UO_2469 (O_2469,N_19927,N_19902);
or UO_2470 (O_2470,N_19967,N_19850);
and UO_2471 (O_2471,N_19990,N_19880);
and UO_2472 (O_2472,N_19884,N_19977);
xor UO_2473 (O_2473,N_19869,N_19929);
and UO_2474 (O_2474,N_19997,N_19944);
nand UO_2475 (O_2475,N_19977,N_19883);
xnor UO_2476 (O_2476,N_19975,N_19958);
xor UO_2477 (O_2477,N_19844,N_19920);
and UO_2478 (O_2478,N_19988,N_19875);
or UO_2479 (O_2479,N_19989,N_19853);
xnor UO_2480 (O_2480,N_19947,N_19870);
and UO_2481 (O_2481,N_19939,N_19840);
xnor UO_2482 (O_2482,N_19912,N_19855);
nand UO_2483 (O_2483,N_19968,N_19954);
or UO_2484 (O_2484,N_19931,N_19882);
or UO_2485 (O_2485,N_19844,N_19936);
and UO_2486 (O_2486,N_19968,N_19896);
nor UO_2487 (O_2487,N_19978,N_19856);
and UO_2488 (O_2488,N_19925,N_19929);
xor UO_2489 (O_2489,N_19997,N_19970);
or UO_2490 (O_2490,N_19986,N_19854);
xor UO_2491 (O_2491,N_19931,N_19874);
and UO_2492 (O_2492,N_19916,N_19999);
or UO_2493 (O_2493,N_19883,N_19891);
or UO_2494 (O_2494,N_19854,N_19868);
nor UO_2495 (O_2495,N_19959,N_19945);
nand UO_2496 (O_2496,N_19899,N_19958);
nor UO_2497 (O_2497,N_19883,N_19936);
nor UO_2498 (O_2498,N_19876,N_19971);
or UO_2499 (O_2499,N_19927,N_19950);
endmodule