module basic_1000_10000_1500_2_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5002,N_5004,N_5005,N_5006,N_5007,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5020,N_5021,N_5022,N_5027,N_5029,N_5030,N_5031,N_5034,N_5036,N_5040,N_5041,N_5043,N_5044,N_5045,N_5046,N_5047,N_5051,N_5052,N_5053,N_5056,N_5057,N_5059,N_5063,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5074,N_5075,N_5081,N_5085,N_5086,N_5087,N_5088,N_5089,N_5092,N_5093,N_5095,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5107,N_5108,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5117,N_5120,N_5121,N_5122,N_5124,N_5125,N_5126,N_5128,N_5130,N_5131,N_5132,N_5133,N_5134,N_5136,N_5137,N_5139,N_5140,N_5145,N_5146,N_5147,N_5149,N_5150,N_5155,N_5156,N_5158,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5168,N_5169,N_5170,N_5172,N_5175,N_5178,N_5180,N_5182,N_5183,N_5185,N_5187,N_5188,N_5192,N_5195,N_5197,N_5198,N_5199,N_5200,N_5202,N_5205,N_5207,N_5209,N_5212,N_5214,N_5217,N_5219,N_5222,N_5224,N_5227,N_5228,N_5229,N_5231,N_5232,N_5233,N_5248,N_5249,N_5251,N_5252,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5263,N_5265,N_5267,N_5268,N_5269,N_5271,N_5274,N_5277,N_5279,N_5280,N_5281,N_5284,N_5287,N_5289,N_5290,N_5291,N_5292,N_5293,N_5296,N_5297,N_5298,N_5300,N_5301,N_5302,N_5303,N_5304,N_5306,N_5308,N_5311,N_5313,N_5315,N_5316,N_5320,N_5321,N_5323,N_5325,N_5328,N_5330,N_5331,N_5333,N_5335,N_5336,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5345,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5354,N_5355,N_5356,N_5360,N_5362,N_5363,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5373,N_5374,N_5376,N_5379,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5392,N_5393,N_5396,N_5397,N_5399,N_5403,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5414,N_5415,N_5416,N_5420,N_5421,N_5422,N_5424,N_5425,N_5426,N_5427,N_5428,N_5430,N_5431,N_5432,N_5433,N_5434,N_5436,N_5437,N_5438,N_5440,N_5443,N_5444,N_5445,N_5446,N_5453,N_5455,N_5456,N_5458,N_5459,N_5461,N_5464,N_5465,N_5467,N_5468,N_5469,N_5472,N_5475,N_5477,N_5478,N_5479,N_5482,N_5483,N_5484,N_5485,N_5486,N_5489,N_5492,N_5493,N_5495,N_5497,N_5498,N_5501,N_5505,N_5507,N_5508,N_5509,N_5512,N_5513,N_5514,N_5515,N_5518,N_5520,N_5522,N_5525,N_5526,N_5527,N_5528,N_5529,N_5534,N_5535,N_5536,N_5537,N_5539,N_5545,N_5546,N_5547,N_5549,N_5550,N_5553,N_5554,N_5556,N_5558,N_5559,N_5561,N_5566,N_5567,N_5568,N_5569,N_5571,N_5572,N_5575,N_5576,N_5577,N_5580,N_5581,N_5583,N_5584,N_5585,N_5586,N_5591,N_5593,N_5595,N_5596,N_5598,N_5599,N_5600,N_5601,N_5602,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5614,N_5615,N_5617,N_5618,N_5620,N_5621,N_5622,N_5623,N_5629,N_5631,N_5633,N_5634,N_5636,N_5638,N_5639,N_5640,N_5641,N_5642,N_5644,N_5648,N_5649,N_5650,N_5651,N_5653,N_5654,N_5656,N_5657,N_5658,N_5659,N_5661,N_5662,N_5663,N_5666,N_5667,N_5668,N_5670,N_5671,N_5673,N_5674,N_5675,N_5677,N_5678,N_5680,N_5681,N_5683,N_5684,N_5685,N_5688,N_5690,N_5691,N_5693,N_5696,N_5698,N_5700,N_5701,N_5702,N_5703,N_5706,N_5707,N_5708,N_5709,N_5710,N_5712,N_5716,N_5719,N_5721,N_5723,N_5724,N_5725,N_5727,N_5729,N_5732,N_5733,N_5734,N_5735,N_5736,N_5738,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5748,N_5749,N_5750,N_5751,N_5753,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5763,N_5765,N_5769,N_5770,N_5771,N_5773,N_5774,N_5779,N_5780,N_5783,N_5787,N_5788,N_5793,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5803,N_5805,N_5807,N_5809,N_5810,N_5812,N_5813,N_5814,N_5815,N_5817,N_5819,N_5820,N_5822,N_5824,N_5826,N_5827,N_5830,N_5831,N_5832,N_5834,N_5836,N_5837,N_5838,N_5839,N_5841,N_5842,N_5843,N_5844,N_5845,N_5847,N_5851,N_5852,N_5853,N_5854,N_5856,N_5857,N_5858,N_5859,N_5860,N_5862,N_5863,N_5866,N_5867,N_5869,N_5870,N_5871,N_5873,N_5875,N_5876,N_5877,N_5879,N_5881,N_5883,N_5884,N_5885,N_5888,N_5893,N_5894,N_5895,N_5896,N_5898,N_5900,N_5901,N_5902,N_5903,N_5904,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5915,N_5917,N_5923,N_5924,N_5925,N_5926,N_5928,N_5929,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5939,N_5940,N_5941,N_5942,N_5944,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5955,N_5956,N_5958,N_5959,N_5962,N_5963,N_5965,N_5966,N_5967,N_5968,N_5969,N_5971,N_5972,N_5973,N_5974,N_5975,N_5977,N_5978,N_5980,N_5982,N_5984,N_5985,N_5986,N_5987,N_5988,N_5990,N_5991,N_5992,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6004,N_6005,N_6010,N_6015,N_6016,N_6019,N_6020,N_6021,N_6023,N_6025,N_6026,N_6028,N_6029,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6040,N_6041,N_6042,N_6043,N_6046,N_6047,N_6048,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6058,N_6059,N_6060,N_6065,N_6066,N_6067,N_6070,N_6071,N_6072,N_6073,N_6076,N_6077,N_6078,N_6080,N_6082,N_6083,N_6085,N_6089,N_6091,N_6093,N_6094,N_6095,N_6096,N_6099,N_6100,N_6101,N_6102,N_6104,N_6105,N_6108,N_6109,N_6110,N_6111,N_6113,N_6115,N_6116,N_6118,N_6122,N_6123,N_6125,N_6126,N_6128,N_6130,N_6131,N_6134,N_6135,N_6136,N_6137,N_6138,N_6140,N_6142,N_6145,N_6146,N_6147,N_6148,N_6149,N_6153,N_6156,N_6158,N_6162,N_6163,N_6164,N_6166,N_6169,N_6171,N_6173,N_6175,N_6176,N_6177,N_6181,N_6183,N_6185,N_6186,N_6188,N_6190,N_6191,N_6193,N_6194,N_6195,N_6196,N_6198,N_6200,N_6203,N_6204,N_6207,N_6208,N_6209,N_6212,N_6213,N_6214,N_6216,N_6218,N_6219,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6234,N_6235,N_6236,N_6238,N_6239,N_6241,N_6243,N_6244,N_6246,N_6247,N_6248,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6258,N_6260,N_6261,N_6262,N_6263,N_6266,N_6267,N_6268,N_6269,N_6270,N_6272,N_6273,N_6274,N_6275,N_6276,N_6279,N_6281,N_6282,N_6283,N_6285,N_6286,N_6287,N_6288,N_6290,N_6292,N_6294,N_6295,N_6296,N_6297,N_6299,N_6302,N_6304,N_6305,N_6306,N_6308,N_6309,N_6313,N_6314,N_6317,N_6319,N_6320,N_6322,N_6323,N_6326,N_6328,N_6332,N_6334,N_6335,N_6336,N_6338,N_6341,N_6345,N_6347,N_6348,N_6349,N_6350,N_6351,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6360,N_6364,N_6365,N_6368,N_6369,N_6374,N_6375,N_6376,N_6378,N_6379,N_6381,N_6382,N_6388,N_6389,N_6391,N_6393,N_6394,N_6397,N_6398,N_6399,N_6402,N_6404,N_6405,N_6407,N_6408,N_6409,N_6415,N_6419,N_6420,N_6421,N_6422,N_6425,N_6427,N_6428,N_6430,N_6431,N_6432,N_6433,N_6434,N_6436,N_6437,N_6441,N_6443,N_6445,N_6449,N_6450,N_6451,N_6452,N_6453,N_6455,N_6457,N_6459,N_6460,N_6461,N_6462,N_6464,N_6465,N_6466,N_6468,N_6472,N_6473,N_6475,N_6478,N_6479,N_6480,N_6481,N_6483,N_6485,N_6486,N_6490,N_6491,N_6492,N_6493,N_6495,N_6497,N_6498,N_6499,N_6500,N_6501,N_6503,N_6505,N_6507,N_6509,N_6510,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6520,N_6521,N_6525,N_6526,N_6529,N_6531,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6563,N_6565,N_6567,N_6569,N_6570,N_6572,N_6574,N_6575,N_6576,N_6577,N_6580,N_6581,N_6582,N_6584,N_6585,N_6586,N_6588,N_6590,N_6592,N_6595,N_6596,N_6597,N_6599,N_6600,N_6601,N_6602,N_6603,N_6605,N_6606,N_6607,N_6613,N_6616,N_6618,N_6619,N_6620,N_6622,N_6624,N_6627,N_6628,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6642,N_6644,N_6645,N_6650,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6665,N_6666,N_6668,N_6670,N_6671,N_6673,N_6674,N_6675,N_6677,N_6680,N_6682,N_6685,N_6687,N_6689,N_6691,N_6692,N_6695,N_6696,N_6698,N_6700,N_6703,N_6704,N_6705,N_6706,N_6708,N_6709,N_6710,N_6712,N_6714,N_6716,N_6718,N_6721,N_6722,N_6723,N_6724,N_6725,N_6727,N_6728,N_6729,N_6730,N_6732,N_6733,N_6736,N_6738,N_6739,N_6742,N_6745,N_6747,N_6748,N_6750,N_6751,N_6753,N_6756,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6769,N_6770,N_6771,N_6774,N_6775,N_6776,N_6779,N_6780,N_6781,N_6785,N_6787,N_6788,N_6789,N_6791,N_6792,N_6794,N_6797,N_6798,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6809,N_6810,N_6811,N_6812,N_6815,N_6817,N_6819,N_6820,N_6821,N_6823,N_6824,N_6827,N_6828,N_6829,N_6831,N_6832,N_6833,N_6834,N_6839,N_6840,N_6841,N_6842,N_6843,N_6847,N_6848,N_6852,N_6853,N_6854,N_6855,N_6856,N_6858,N_6861,N_6862,N_6865,N_6868,N_6870,N_6871,N_6872,N_6873,N_6874,N_6877,N_6880,N_6883,N_6884,N_6889,N_6890,N_6896,N_6899,N_6900,N_6903,N_6904,N_6905,N_6906,N_6908,N_6909,N_6910,N_6911,N_6913,N_6914,N_6916,N_6917,N_6921,N_6922,N_6923,N_6927,N_6929,N_6931,N_6932,N_6936,N_6937,N_6939,N_6943,N_6944,N_6947,N_6948,N_6950,N_6951,N_6955,N_6957,N_6958,N_6959,N_6960,N_6962,N_6963,N_6964,N_6965,N_6966,N_6968,N_6969,N_6972,N_6974,N_6975,N_6976,N_6978,N_6981,N_6982,N_6983,N_6984,N_6985,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6996,N_6997,N_6998,N_6999,N_7004,N_7005,N_7008,N_7009,N_7011,N_7013,N_7016,N_7017,N_7018,N_7020,N_7022,N_7023,N_7024,N_7025,N_7027,N_7030,N_7031,N_7032,N_7033,N_7035,N_7036,N_7037,N_7040,N_7041,N_7042,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7055,N_7057,N_7058,N_7059,N_7061,N_7064,N_7065,N_7068,N_7072,N_7074,N_7079,N_7080,N_7082,N_7083,N_7085,N_7087,N_7089,N_7090,N_7092,N_7094,N_7095,N_7097,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7118,N_7119,N_7120,N_7121,N_7124,N_7129,N_7131,N_7132,N_7133,N_7134,N_7135,N_7137,N_7139,N_7143,N_7144,N_7150,N_7151,N_7152,N_7155,N_7157,N_7158,N_7164,N_7166,N_7168,N_7169,N_7171,N_7172,N_7173,N_7177,N_7178,N_7179,N_7181,N_7182,N_7184,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7194,N_7197,N_7198,N_7199,N_7200,N_7202,N_7203,N_7204,N_7205,N_7206,N_7209,N_7211,N_7212,N_7213,N_7214,N_7216,N_7219,N_7220,N_7221,N_7222,N_7224,N_7227,N_7229,N_7230,N_7233,N_7234,N_7235,N_7236,N_7237,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7247,N_7248,N_7249,N_7250,N_7253,N_7254,N_7255,N_7257,N_7258,N_7259,N_7261,N_7265,N_7267,N_7268,N_7269,N_7271,N_7273,N_7274,N_7275,N_7277,N_7279,N_7281,N_7284,N_7285,N_7286,N_7289,N_7291,N_7292,N_7295,N_7296,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7305,N_7309,N_7310,N_7314,N_7315,N_7317,N_7320,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7330,N_7331,N_7333,N_7334,N_7336,N_7337,N_7338,N_7339,N_7341,N_7342,N_7343,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7355,N_7356,N_7359,N_7361,N_7362,N_7363,N_7366,N_7368,N_7369,N_7372,N_7373,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7383,N_7384,N_7385,N_7387,N_7388,N_7390,N_7392,N_7393,N_7397,N_7398,N_7401,N_7402,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7412,N_7413,N_7414,N_7415,N_7416,N_7418,N_7419,N_7420,N_7422,N_7423,N_7425,N_7428,N_7429,N_7430,N_7432,N_7433,N_7434,N_7436,N_7437,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7448,N_7450,N_7451,N_7452,N_7453,N_7460,N_7462,N_7465,N_7467,N_7468,N_7469,N_7470,N_7472,N_7473,N_7475,N_7477,N_7480,N_7481,N_7482,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7495,N_7497,N_7503,N_7507,N_7509,N_7510,N_7514,N_7515,N_7516,N_7517,N_7518,N_7521,N_7523,N_7524,N_7527,N_7528,N_7529,N_7531,N_7532,N_7534,N_7536,N_7537,N_7538,N_7539,N_7540,N_7542,N_7543,N_7545,N_7547,N_7548,N_7550,N_7553,N_7554,N_7556,N_7557,N_7560,N_7562,N_7563,N_7565,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7576,N_7577,N_7578,N_7581,N_7583,N_7585,N_7586,N_7587,N_7588,N_7589,N_7591,N_7592,N_7594,N_7595,N_7597,N_7598,N_7599,N_7602,N_7603,N_7604,N_7607,N_7609,N_7610,N_7611,N_7613,N_7614,N_7617,N_7618,N_7621,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7635,N_7636,N_7637,N_7638,N_7639,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7651,N_7652,N_7653,N_7654,N_7657,N_7658,N_7660,N_7662,N_7663,N_7664,N_7666,N_7668,N_7670,N_7671,N_7672,N_7673,N_7675,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7701,N_7702,N_7703,N_7704,N_7705,N_7708,N_7709,N_7711,N_7713,N_7714,N_7715,N_7717,N_7718,N_7720,N_7726,N_7728,N_7730,N_7732,N_7734,N_7736,N_7737,N_7738,N_7744,N_7745,N_7746,N_7747,N_7750,N_7751,N_7753,N_7754,N_7755,N_7758,N_7760,N_7761,N_7762,N_7763,N_7766,N_7769,N_7772,N_7773,N_7775,N_7777,N_7779,N_7780,N_7781,N_7783,N_7785,N_7786,N_7787,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7797,N_7799,N_7802,N_7803,N_7805,N_7807,N_7809,N_7810,N_7811,N_7814,N_7815,N_7819,N_7820,N_7821,N_7824,N_7825,N_7827,N_7828,N_7830,N_7836,N_7837,N_7838,N_7839,N_7842,N_7843,N_7844,N_7846,N_7849,N_7850,N_7851,N_7855,N_7856,N_7858,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7869,N_7870,N_7871,N_7873,N_7874,N_7876,N_7878,N_7879,N_7881,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7899,N_7901,N_7903,N_7907,N_7908,N_7909,N_7911,N_7912,N_7916,N_7917,N_7918,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7932,N_7934,N_7936,N_7937,N_7938,N_7939,N_7945,N_7946,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7957,N_7958,N_7959,N_7961,N_7964,N_7967,N_7968,N_7969,N_7974,N_7976,N_7977,N_7979,N_7980,N_7983,N_7985,N_7986,N_7987,N_7988,N_7989,N_7992,N_7995,N_7996,N_7998,N_7999,N_8000,N_8004,N_8005,N_8010,N_8012,N_8013,N_8017,N_8018,N_8019,N_8023,N_8024,N_8025,N_8026,N_8028,N_8029,N_8030,N_8031,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8044,N_8045,N_8046,N_8047,N_8048,N_8050,N_8052,N_8053,N_8054,N_8055,N_8056,N_8058,N_8059,N_8061,N_8063,N_8064,N_8065,N_8066,N_8067,N_8069,N_8070,N_8071,N_8075,N_8076,N_8079,N_8080,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8094,N_8095,N_8096,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8105,N_8106,N_8107,N_8108,N_8110,N_8113,N_8114,N_8115,N_8118,N_8119,N_8120,N_8122,N_8123,N_8124,N_8125,N_8126,N_8128,N_8129,N_8130,N_8131,N_8133,N_8134,N_8136,N_8137,N_8138,N_8139,N_8140,N_8143,N_8144,N_8146,N_8147,N_8148,N_8152,N_8153,N_8154,N_8155,N_8159,N_8160,N_8162,N_8166,N_8167,N_8168,N_8170,N_8173,N_8174,N_8176,N_8181,N_8184,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8194,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8209,N_8211,N_8214,N_8216,N_8218,N_8219,N_8221,N_8227,N_8232,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8246,N_8248,N_8250,N_8251,N_8252,N_8253,N_8254,N_8256,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8268,N_8269,N_8271,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8281,N_8282,N_8283,N_8285,N_8286,N_8287,N_8288,N_8289,N_8291,N_8293,N_8296,N_8298,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8309,N_8311,N_8312,N_8313,N_8314,N_8316,N_8317,N_8318,N_8319,N_8321,N_8322,N_8325,N_8326,N_8329,N_8330,N_8332,N_8334,N_8335,N_8336,N_8340,N_8341,N_8342,N_8344,N_8345,N_8348,N_8349,N_8353,N_8354,N_8355,N_8356,N_8358,N_8360,N_8364,N_8366,N_8368,N_8371,N_8374,N_8377,N_8378,N_8381,N_8385,N_8386,N_8388,N_8389,N_8394,N_8395,N_8396,N_8398,N_8399,N_8400,N_8401,N_8402,N_8404,N_8405,N_8406,N_8408,N_8409,N_8410,N_8411,N_8414,N_8415,N_8416,N_8417,N_8419,N_8421,N_8422,N_8424,N_8425,N_8428,N_8429,N_8431,N_8432,N_8433,N_8436,N_8437,N_8439,N_8441,N_8442,N_8443,N_8444,N_8446,N_8449,N_8450,N_8452,N_8454,N_8455,N_8457,N_8458,N_8459,N_8460,N_8461,N_8463,N_8465,N_8467,N_8468,N_8472,N_8475,N_8476,N_8477,N_8478,N_8479,N_8482,N_8485,N_8487,N_8489,N_8491,N_8492,N_8496,N_8497,N_8498,N_8499,N_8500,N_8506,N_8509,N_8510,N_8512,N_8514,N_8515,N_8517,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8529,N_8530,N_8532,N_8533,N_8535,N_8538,N_8541,N_8544,N_8546,N_8550,N_8551,N_8553,N_8555,N_8556,N_8561,N_8562,N_8570,N_8572,N_8573,N_8576,N_8577,N_8578,N_8579,N_8580,N_8585,N_8586,N_8587,N_8592,N_8593,N_8596,N_8599,N_8600,N_8601,N_8604,N_8609,N_8611,N_8613,N_8614,N_8615,N_8618,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8631,N_8634,N_8636,N_8637,N_8639,N_8640,N_8641,N_8642,N_8645,N_8646,N_8647,N_8649,N_8652,N_8654,N_8655,N_8657,N_8658,N_8659,N_8661,N_8662,N_8663,N_8665,N_8667,N_8670,N_8671,N_8673,N_8675,N_8676,N_8680,N_8681,N_8683,N_8684,N_8686,N_8688,N_8689,N_8690,N_8691,N_8693,N_8694,N_8695,N_8697,N_8698,N_8699,N_8701,N_8702,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8712,N_8715,N_8717,N_8719,N_8720,N_8726,N_8727,N_8728,N_8731,N_8733,N_8734,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8749,N_8750,N_8752,N_8753,N_8754,N_8756,N_8757,N_8758,N_8762,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8772,N_8774,N_8775,N_8776,N_8779,N_8780,N_8781,N_8782,N_8783,N_8785,N_8786,N_8788,N_8790,N_8794,N_8795,N_8797,N_8798,N_8799,N_8800,N_8802,N_8804,N_8805,N_8807,N_8809,N_8813,N_8814,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8826,N_8829,N_8830,N_8834,N_8835,N_8836,N_8837,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8851,N_8855,N_8857,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8868,N_8870,N_8872,N_8874,N_8877,N_8878,N_8879,N_8881,N_8883,N_8885,N_8886,N_8887,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8899,N_8900,N_8901,N_8902,N_8906,N_8907,N_8911,N_8912,N_8916,N_8918,N_8919,N_8921,N_8922,N_8923,N_8924,N_8925,N_8927,N_8928,N_8930,N_8934,N_8935,N_8939,N_8942,N_8944,N_8945,N_8947,N_8949,N_8950,N_8951,N_8952,N_8955,N_8956,N_8960,N_8961,N_8962,N_8963,N_8964,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8980,N_8981,N_8983,N_8986,N_8990,N_8991,N_8994,N_8995,N_8996,N_8997,N_8998,N_9000,N_9002,N_9003,N_9004,N_9006,N_9007,N_9010,N_9011,N_9012,N_9013,N_9015,N_9017,N_9018,N_9019,N_9020,N_9021,N_9023,N_9024,N_9025,N_9028,N_9029,N_9030,N_9031,N_9036,N_9038,N_9039,N_9040,N_9041,N_9043,N_9044,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9054,N_9056,N_9057,N_9058,N_9059,N_9061,N_9062,N_9064,N_9065,N_9067,N_9068,N_9071,N_9072,N_9074,N_9076,N_9078,N_9079,N_9080,N_9081,N_9083,N_9085,N_9087,N_9090,N_9092,N_9093,N_9095,N_9096,N_9097,N_9098,N_9099,N_9101,N_9102,N_9103,N_9105,N_9106,N_9109,N_9111,N_9112,N_9114,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9129,N_9131,N_9132,N_9135,N_9136,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9153,N_9154,N_9155,N_9157,N_9159,N_9161,N_9163,N_9167,N_9169,N_9170,N_9175,N_9176,N_9177,N_9178,N_9179,N_9181,N_9182,N_9183,N_9184,N_9187,N_9190,N_9193,N_9195,N_9197,N_9198,N_9199,N_9202,N_9204,N_9205,N_9207,N_9208,N_9209,N_9212,N_9213,N_9214,N_9217,N_9219,N_9220,N_9221,N_9222,N_9228,N_9229,N_9231,N_9232,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9243,N_9244,N_9245,N_9247,N_9249,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9264,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9283,N_9285,N_9287,N_9288,N_9289,N_9294,N_9295,N_9296,N_9300,N_9303,N_9304,N_9307,N_9308,N_9310,N_9311,N_9312,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9325,N_9326,N_9328,N_9329,N_9331,N_9333,N_9334,N_9338,N_9339,N_9342,N_9343,N_9344,N_9345,N_9347,N_9348,N_9350,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9359,N_9360,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9371,N_9373,N_9374,N_9375,N_9376,N_9378,N_9379,N_9381,N_9386,N_9387,N_9389,N_9390,N_9392,N_9393,N_9394,N_9395,N_9397,N_9398,N_9399,N_9402,N_9403,N_9404,N_9405,N_9406,N_9408,N_9409,N_9412,N_9413,N_9416,N_9417,N_9418,N_9420,N_9421,N_9422,N_9425,N_9426,N_9428,N_9429,N_9430,N_9432,N_9434,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9448,N_9450,N_9452,N_9455,N_9456,N_9457,N_9458,N_9461,N_9462,N_9463,N_9464,N_9465,N_9467,N_9469,N_9471,N_9473,N_9474,N_9475,N_9476,N_9478,N_9483,N_9484,N_9486,N_9487,N_9489,N_9491,N_9493,N_9495,N_9496,N_9497,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9512,N_9513,N_9515,N_9517,N_9519,N_9520,N_9521,N_9522,N_9524,N_9527,N_9529,N_9531,N_9533,N_9534,N_9535,N_9536,N_9537,N_9539,N_9541,N_9542,N_9543,N_9548,N_9549,N_9551,N_9552,N_9554,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9564,N_9566,N_9572,N_9574,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9587,N_9589,N_9591,N_9594,N_9595,N_9596,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9605,N_9606,N_9607,N_9609,N_9611,N_9612,N_9613,N_9616,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9644,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9660,N_9662,N_9663,N_9664,N_9666,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9679,N_9680,N_9681,N_9683,N_9684,N_9686,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9698,N_9700,N_9702,N_9703,N_9705,N_9707,N_9708,N_9709,N_9711,N_9712,N_9713,N_9715,N_9716,N_9720,N_9722,N_9724,N_9727,N_9728,N_9729,N_9730,N_9731,N_9734,N_9735,N_9739,N_9742,N_9744,N_9745,N_9746,N_9748,N_9749,N_9751,N_9752,N_9753,N_9759,N_9761,N_9763,N_9764,N_9766,N_9767,N_9768,N_9770,N_9773,N_9775,N_9776,N_9777,N_9778,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9787,N_9788,N_9789,N_9790,N_9792,N_9793,N_9795,N_9796,N_9798,N_9801,N_9806,N_9807,N_9808,N_9812,N_9814,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9823,N_9824,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9833,N_9835,N_9836,N_9840,N_9842,N_9845,N_9848,N_9849,N_9850,N_9852,N_9853,N_9854,N_9855,N_9861,N_9862,N_9864,N_9865,N_9866,N_9867,N_9868,N_9874,N_9876,N_9877,N_9880,N_9881,N_9883,N_9886,N_9887,N_9889,N_9890,N_9893,N_9896,N_9897,N_9900,N_9901,N_9906,N_9908,N_9909,N_9910,N_9911,N_9914,N_9916,N_9918,N_9921,N_9922,N_9926,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9936,N_9939,N_9941,N_9946,N_9947,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9959,N_9960,N_9961,N_9963,N_9964,N_9965,N_9966,N_9970,N_9972,N_9973,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9984,N_9985,N_9988,N_9989,N_9990,N_9995,N_9997,N_9998,N_9999;
or U0 (N_0,In_575,In_853);
and U1 (N_1,In_914,In_507);
and U2 (N_2,In_186,In_585);
nand U3 (N_3,In_735,In_114);
nand U4 (N_4,In_763,In_97);
nand U5 (N_5,In_627,In_330);
or U6 (N_6,In_551,In_443);
or U7 (N_7,In_506,In_749);
and U8 (N_8,In_728,In_11);
nand U9 (N_9,In_98,In_458);
nor U10 (N_10,In_435,In_845);
and U11 (N_11,In_319,In_215);
and U12 (N_12,In_717,In_648);
xor U13 (N_13,In_838,In_349);
xor U14 (N_14,In_850,In_398);
or U15 (N_15,In_290,In_108);
nor U16 (N_16,In_940,In_988);
and U17 (N_17,In_689,In_158);
nand U18 (N_18,In_391,In_746);
nor U19 (N_19,In_467,In_217);
or U20 (N_20,In_273,In_166);
nor U21 (N_21,In_979,In_687);
or U22 (N_22,In_255,In_296);
nand U23 (N_23,In_906,In_780);
xor U24 (N_24,In_250,In_303);
nand U25 (N_25,In_21,In_457);
nor U26 (N_26,In_710,In_346);
or U27 (N_27,In_269,In_619);
nor U28 (N_28,In_495,In_995);
nand U29 (N_29,In_563,In_220);
and U30 (N_30,In_82,In_697);
or U31 (N_31,In_417,In_422);
and U32 (N_32,In_676,In_253);
or U33 (N_33,In_700,In_726);
nand U34 (N_34,In_858,In_798);
or U35 (N_35,In_187,In_712);
nand U36 (N_36,In_786,In_447);
nand U37 (N_37,In_883,In_565);
nor U38 (N_38,In_571,In_970);
or U39 (N_39,In_863,In_913);
nand U40 (N_40,In_386,In_56);
and U41 (N_41,In_51,In_288);
nor U42 (N_42,In_315,In_229);
and U43 (N_43,In_93,In_668);
or U44 (N_44,In_76,In_441);
nand U45 (N_45,In_163,In_372);
nor U46 (N_46,In_63,In_946);
or U47 (N_47,In_891,In_626);
nor U48 (N_48,In_823,In_607);
nand U49 (N_49,In_399,In_478);
and U50 (N_50,In_683,In_459);
nand U51 (N_51,In_87,In_910);
and U52 (N_52,In_953,In_201);
nand U53 (N_53,In_453,In_722);
nand U54 (N_54,In_942,In_895);
nor U55 (N_55,In_72,In_715);
and U56 (N_56,In_91,In_742);
and U57 (N_57,In_353,In_524);
nor U58 (N_58,In_941,In_831);
nand U59 (N_59,In_170,In_385);
or U60 (N_60,In_111,In_112);
and U61 (N_61,In_643,In_909);
nand U62 (N_62,In_699,In_981);
and U63 (N_63,In_813,In_358);
and U64 (N_64,In_937,In_38);
nand U65 (N_65,In_44,In_123);
and U66 (N_66,In_90,In_471);
or U67 (N_67,In_88,In_233);
nor U68 (N_68,In_768,In_963);
or U69 (N_69,In_598,In_541);
nand U70 (N_70,In_679,In_367);
nor U71 (N_71,In_390,In_511);
nand U72 (N_72,In_164,In_868);
nand U73 (N_73,In_53,In_420);
and U74 (N_74,In_802,In_282);
nor U75 (N_75,In_355,In_204);
and U76 (N_76,In_211,In_968);
or U77 (N_77,In_176,In_101);
or U78 (N_78,In_415,In_787);
and U79 (N_79,In_528,In_210);
and U80 (N_80,In_789,In_948);
nor U81 (N_81,In_128,In_359);
nor U82 (N_82,In_394,In_505);
nand U83 (N_83,In_335,In_960);
and U84 (N_84,In_446,In_851);
or U85 (N_85,In_852,In_522);
nand U86 (N_86,In_487,In_543);
or U87 (N_87,In_587,In_915);
or U88 (N_88,In_939,In_998);
nand U89 (N_89,In_148,In_804);
or U90 (N_90,In_835,In_468);
or U91 (N_91,In_957,In_232);
nor U92 (N_92,In_149,In_413);
or U93 (N_93,In_493,In_212);
nor U94 (N_94,In_83,In_143);
or U95 (N_95,In_388,In_50);
and U96 (N_96,In_442,In_199);
and U97 (N_97,In_664,In_558);
or U98 (N_98,In_281,In_252);
or U99 (N_99,In_411,In_969);
nand U100 (N_100,In_188,In_757);
and U101 (N_101,In_280,In_449);
nand U102 (N_102,In_736,In_228);
or U103 (N_103,In_698,In_864);
nor U104 (N_104,In_124,In_959);
and U105 (N_105,In_274,In_974);
nor U106 (N_106,In_284,In_2);
and U107 (N_107,In_729,In_387);
nand U108 (N_108,In_251,In_965);
and U109 (N_109,In_438,In_616);
and U110 (N_110,In_337,In_613);
or U111 (N_111,In_494,In_535);
and U112 (N_112,In_33,In_918);
nor U113 (N_113,In_944,In_748);
or U114 (N_114,In_539,In_999);
and U115 (N_115,In_404,In_557);
nor U116 (N_116,In_134,In_336);
nand U117 (N_117,In_907,In_426);
nor U118 (N_118,In_136,In_191);
and U119 (N_119,In_66,In_16);
nand U120 (N_120,In_295,In_892);
nor U121 (N_121,In_32,In_964);
and U122 (N_122,In_833,In_455);
or U123 (N_123,In_520,In_120);
nor U124 (N_124,In_238,In_949);
nor U125 (N_125,In_65,In_327);
and U126 (N_126,In_671,In_793);
and U127 (N_127,In_560,In_854);
and U128 (N_128,In_466,In_80);
nor U129 (N_129,In_380,In_828);
or U130 (N_130,In_107,In_633);
and U131 (N_131,In_23,In_921);
or U132 (N_132,In_206,In_890);
or U133 (N_133,In_876,In_339);
nor U134 (N_134,In_423,In_778);
nor U135 (N_135,In_92,In_834);
and U136 (N_136,In_405,In_923);
or U137 (N_137,In_272,In_71);
and U138 (N_138,In_977,In_313);
nand U139 (N_139,In_256,In_922);
and U140 (N_140,In_967,In_917);
nand U141 (N_141,In_397,In_69);
nand U142 (N_142,In_860,In_925);
nor U143 (N_143,In_160,In_642);
nand U144 (N_144,In_46,In_951);
nor U145 (N_145,In_434,In_73);
nor U146 (N_146,In_733,In_461);
nand U147 (N_147,In_580,In_983);
and U148 (N_148,In_325,In_481);
nor U149 (N_149,In_504,In_5);
nor U150 (N_150,In_317,In_817);
or U151 (N_151,In_975,In_617);
nor U152 (N_152,In_432,In_376);
nand U153 (N_153,In_234,In_573);
nor U154 (N_154,In_591,In_456);
nor U155 (N_155,In_695,In_329);
or U156 (N_156,In_118,In_338);
nand U157 (N_157,In_27,In_589);
or U158 (N_158,In_138,In_875);
nor U159 (N_159,In_320,In_58);
nor U160 (N_160,In_95,In_360);
nand U161 (N_161,In_155,In_127);
nand U162 (N_162,In_846,In_418);
nand U163 (N_163,In_930,In_6);
or U164 (N_164,In_324,In_132);
or U165 (N_165,In_830,In_905);
or U166 (N_166,In_427,In_862);
nand U167 (N_167,In_214,In_609);
nand U168 (N_168,In_744,In_908);
nand U169 (N_169,In_570,In_1);
or U170 (N_170,In_472,In_774);
nand U171 (N_171,In_685,In_276);
nor U172 (N_172,In_821,In_248);
or U173 (N_173,In_646,In_634);
nand U174 (N_174,In_615,In_96);
nand U175 (N_175,In_486,In_22);
nand U176 (N_176,In_696,In_393);
or U177 (N_177,In_601,In_309);
nor U178 (N_178,In_644,In_952);
nor U179 (N_179,In_612,In_622);
and U180 (N_180,In_167,In_488);
nand U181 (N_181,In_738,In_556);
or U182 (N_182,In_990,In_168);
and U183 (N_183,In_829,In_719);
xnor U184 (N_184,In_430,In_750);
or U185 (N_185,In_912,In_564);
or U186 (N_186,In_364,In_165);
nor U187 (N_187,In_377,In_986);
or U188 (N_188,In_992,In_670);
or U189 (N_189,In_278,In_812);
and U190 (N_190,In_826,In_523);
and U191 (N_191,In_597,In_265);
nand U192 (N_192,In_103,In_533);
and U193 (N_193,In_402,In_231);
nor U194 (N_194,In_966,In_752);
nand U195 (N_195,In_635,In_920);
nor U196 (N_196,In_824,In_770);
and U197 (N_197,In_242,In_903);
nor U198 (N_198,In_326,In_395);
and U199 (N_199,In_614,In_703);
nand U200 (N_200,In_623,In_125);
or U201 (N_201,In_929,In_153);
or U202 (N_202,In_663,In_785);
and U203 (N_203,In_344,In_832);
nor U204 (N_204,In_972,In_348);
and U205 (N_205,In_655,In_68);
xnor U206 (N_206,In_224,In_869);
and U207 (N_207,In_790,In_305);
and U208 (N_208,In_536,In_263);
and U209 (N_209,In_352,In_285);
and U210 (N_210,In_665,In_734);
or U211 (N_211,In_289,In_482);
nand U212 (N_212,In_209,In_254);
and U213 (N_213,In_600,In_428);
or U214 (N_214,In_791,In_608);
and U215 (N_215,In_261,In_463);
or U216 (N_216,In_421,In_958);
nor U217 (N_217,In_436,In_678);
nand U218 (N_218,In_307,In_800);
and U219 (N_219,In_842,In_259);
and U220 (N_220,In_70,In_611);
nor U221 (N_221,In_861,In_137);
nor U222 (N_222,In_870,In_89);
nand U223 (N_223,In_424,In_777);
nor U224 (N_224,In_796,In_709);
nor U225 (N_225,In_61,In_419);
or U226 (N_226,In_216,In_566);
and U227 (N_227,In_682,In_521);
or U228 (N_228,In_904,In_691);
nand U229 (N_229,In_287,In_886);
nand U230 (N_230,In_947,In_596);
nand U231 (N_231,In_878,In_175);
or U232 (N_232,In_310,In_450);
and U233 (N_233,In_501,In_818);
nand U234 (N_234,In_694,In_808);
nand U235 (N_235,In_816,In_246);
or U236 (N_236,In_270,In_680);
nand U237 (N_237,In_532,In_384);
nor U238 (N_238,In_445,In_340);
nor U239 (N_239,In_140,In_485);
or U240 (N_240,In_116,In_29);
and U241 (N_241,In_652,In_797);
nand U242 (N_242,In_500,In_859);
nor U243 (N_243,In_145,In_462);
nor U244 (N_244,In_12,In_131);
and U245 (N_245,In_807,In_630);
or U246 (N_246,In_993,In_515);
nand U247 (N_247,In_584,In_286);
xor U248 (N_248,In_213,In_559);
and U249 (N_249,In_311,In_782);
or U250 (N_250,In_332,In_721);
or U251 (N_251,In_299,In_230);
nor U252 (N_252,In_102,In_433);
and U253 (N_253,In_581,In_529);
or U254 (N_254,In_882,In_328);
nor U255 (N_255,In_931,In_264);
nor U256 (N_256,In_100,In_512);
and U257 (N_257,In_971,In_751);
nor U258 (N_258,In_727,In_576);
nor U259 (N_259,In_582,In_599);
and U260 (N_260,In_901,In_341);
or U261 (N_261,In_962,In_221);
and U262 (N_262,In_756,In_516);
nor U263 (N_263,In_141,In_400);
and U264 (N_264,In_258,In_74);
xnor U265 (N_265,In_15,In_654);
or U266 (N_266,In_45,In_954);
nor U267 (N_267,In_677,In_110);
nor U268 (N_268,In_479,In_241);
nor U269 (N_269,In_379,In_498);
nand U270 (N_270,In_115,In_55);
or U271 (N_271,In_26,In_179);
nand U272 (N_272,In_249,In_126);
xor U273 (N_273,In_193,In_189);
nand U274 (N_274,In_840,In_531);
or U275 (N_275,In_753,In_545);
nor U276 (N_276,In_59,In_933);
and U277 (N_277,In_991,In_17);
or U278 (N_278,In_629,In_718);
and U279 (N_279,In_898,In_13);
and U280 (N_280,In_927,In_156);
or U281 (N_281,In_19,In_595);
nor U282 (N_282,In_809,In_740);
or U283 (N_283,In_620,In_347);
nor U284 (N_284,In_78,In_688);
nor U285 (N_285,In_416,In_350);
nand U286 (N_286,In_378,In_171);
and U287 (N_287,In_874,In_976);
and U288 (N_288,In_227,In_173);
nand U289 (N_289,In_534,In_820);
or U290 (N_290,In_638,In_631);
nor U291 (N_291,In_881,In_119);
nor U292 (N_292,In_574,In_579);
nor U293 (N_293,In_469,In_928);
or U294 (N_294,In_117,In_547);
and U295 (N_295,In_705,In_867);
and U296 (N_296,In_99,In_916);
nand U297 (N_297,In_490,In_489);
or U298 (N_298,In_105,In_414);
nand U299 (N_299,In_381,In_444);
and U300 (N_300,In_184,In_980);
or U301 (N_301,In_244,In_109);
and U302 (N_302,In_20,In_7);
and U303 (N_303,In_316,In_900);
nor U304 (N_304,In_185,In_121);
and U305 (N_305,In_130,In_849);
nand U306 (N_306,In_182,In_375);
and U307 (N_307,In_464,In_950);
xor U308 (N_308,In_739,In_262);
nor U309 (N_309,In_645,In_650);
and U310 (N_310,In_621,In_667);
or U311 (N_311,In_767,In_602);
or U312 (N_312,In_568,In_815);
nor U313 (N_313,In_491,In_538);
and U314 (N_314,In_361,In_25);
nand U315 (N_315,In_803,In_159);
nand U316 (N_316,In_509,In_301);
and U317 (N_317,In_162,In_885);
and U318 (N_318,In_431,In_297);
and U319 (N_319,In_139,In_819);
and U320 (N_320,In_773,In_30);
and U321 (N_321,In_877,In_24);
nor U322 (N_322,In_673,In_871);
or U323 (N_323,In_605,In_527);
nand U324 (N_324,In_144,In_439);
xor U325 (N_325,In_169,In_354);
and U326 (N_326,In_425,In_106);
or U327 (N_327,In_784,In_686);
nand U328 (N_328,In_366,In_866);
nand U329 (N_329,In_542,In_460);
nand U330 (N_330,In_496,In_825);
or U331 (N_331,In_692,In_291);
and U332 (N_332,In_530,In_334);
or U333 (N_333,In_492,In_219);
and U334 (N_334,In_934,In_708);
nand U335 (N_335,In_454,In_172);
nand U336 (N_336,In_779,In_195);
nand U337 (N_337,In_755,In_122);
or U338 (N_338,In_382,In_267);
nor U339 (N_339,In_268,In_806);
nand U340 (N_340,In_572,In_14);
and U341 (N_341,In_639,In_625);
or U342 (N_342,In_245,In_503);
xor U343 (N_343,In_470,In_776);
and U344 (N_344,In_856,In_389);
and U345 (N_345,In_684,In_476);
and U346 (N_346,In_997,In_919);
nor U347 (N_347,In_401,In_226);
or U348 (N_348,In_60,In_77);
nor U349 (N_349,In_658,In_693);
or U350 (N_350,In_28,In_847);
and U351 (N_351,In_603,In_312);
nor U352 (N_352,In_129,In_984);
and U353 (N_353,In_661,In_150);
xnor U354 (N_354,In_3,In_762);
and U355 (N_355,In_514,In_844);
and U356 (N_356,In_298,In_766);
or U357 (N_357,In_437,In_562);
and U358 (N_358,In_938,In_180);
and U359 (N_359,In_943,In_896);
xnor U360 (N_360,In_429,In_978);
and U361 (N_361,In_932,In_146);
xor U362 (N_362,In_894,In_183);
and U363 (N_363,In_333,In_588);
nand U364 (N_364,In_865,In_314);
or U365 (N_365,In_151,In_198);
and U366 (N_366,In_300,In_279);
and U367 (N_367,In_519,In_653);
nor U368 (N_368,In_257,In_292);
or U369 (N_369,In_54,In_769);
or U370 (N_370,In_872,In_569);
or U371 (N_371,In_304,In_578);
and U372 (N_372,In_660,In_36);
and U373 (N_373,In_544,In_765);
nand U374 (N_374,In_202,In_0);
nor U375 (N_375,In_716,In_371);
and U376 (N_376,In_935,In_142);
nand U377 (N_377,In_302,In_656);
nor U378 (N_378,In_618,In_239);
nor U379 (N_379,In_711,In_363);
or U380 (N_380,In_540,In_440);
or U381 (N_381,In_731,In_795);
and U382 (N_382,In_659,In_982);
or U383 (N_383,In_794,In_537);
nor U384 (N_384,In_640,In_57);
xor U385 (N_385,In_37,In_518);
nor U386 (N_386,In_758,In_702);
nor U387 (N_387,In_247,In_567);
nand U388 (N_388,In_35,In_357);
or U389 (N_389,In_410,In_737);
nor U390 (N_390,In_887,In_724);
xor U391 (N_391,In_743,In_848);
nor U392 (N_392,In_266,In_190);
nand U393 (N_393,In_104,In_331);
nand U394 (N_394,In_499,In_720);
nor U395 (N_395,In_893,In_508);
and U396 (N_396,In_836,In_884);
and U397 (N_397,In_647,In_178);
or U398 (N_398,In_636,In_662);
nand U399 (N_399,In_632,In_392);
nor U400 (N_400,In_672,In_275);
nor U401 (N_401,In_889,In_873);
nor U402 (N_402,In_465,In_628);
nor U403 (N_403,In_801,In_985);
nand U404 (N_404,In_549,In_85);
nand U405 (N_405,In_356,In_152);
nor U406 (N_406,In_81,In_62);
or U407 (N_407,In_577,In_84);
nor U408 (N_408,In_207,In_480);
nor U409 (N_409,In_723,In_75);
and U410 (N_410,In_713,In_181);
nand U411 (N_411,In_792,In_936);
and U412 (N_412,In_8,In_745);
and U413 (N_413,In_203,In_177);
or U414 (N_414,In_318,In_383);
and U415 (N_415,In_225,In_94);
nor U416 (N_416,In_448,In_771);
nor U417 (N_417,In_759,In_624);
or U418 (N_418,In_641,In_374);
xor U419 (N_419,In_553,In_725);
nand U420 (N_420,In_994,In_474);
nand U421 (N_421,In_49,In_9);
or U422 (N_422,In_64,In_675);
or U423 (N_423,In_218,In_47);
nand U424 (N_424,In_961,In_52);
nand U425 (N_425,In_322,In_681);
nand U426 (N_426,In_194,In_606);
and U427 (N_427,In_406,In_788);
nor U428 (N_428,In_10,In_747);
nor U429 (N_429,In_714,In_513);
nand U430 (N_430,In_732,In_365);
nor U431 (N_431,In_483,In_517);
nand U432 (N_432,In_34,In_706);
or U433 (N_433,In_526,In_197);
nor U434 (N_434,In_987,In_911);
nor U435 (N_435,In_837,In_761);
and U436 (N_436,In_154,In_554);
nand U437 (N_437,In_586,In_924);
or U438 (N_438,In_637,In_649);
and U439 (N_439,In_18,In_237);
or U440 (N_440,In_555,In_955);
and U441 (N_441,In_855,In_510);
nand U442 (N_442,In_666,In_926);
xor U443 (N_443,In_475,In_772);
nand U444 (N_444,In_39,In_996);
and U445 (N_445,In_306,In_4);
nor U446 (N_446,In_408,In_822);
and U447 (N_447,In_451,In_373);
and U448 (N_448,In_989,In_283);
or U449 (N_449,In_502,In_561);
nand U450 (N_450,In_814,In_764);
or U451 (N_451,In_811,In_208);
and U452 (N_452,In_396,In_293);
nand U453 (N_453,In_321,In_308);
and U454 (N_454,In_839,In_42);
and U455 (N_455,In_552,In_161);
nor U456 (N_456,In_741,In_235);
nor U457 (N_457,In_192,In_857);
and U458 (N_458,In_590,In_452);
nor U459 (N_459,In_651,In_323);
or U460 (N_460,In_704,In_370);
nand U461 (N_461,In_945,In_412);
nand U462 (N_462,In_200,In_657);
nor U463 (N_463,In_48,In_113);
and U464 (N_464,In_477,In_754);
nor U465 (N_465,In_174,In_236);
nand U466 (N_466,In_196,In_583);
nor U467 (N_467,In_604,In_294);
or U468 (N_468,In_805,In_147);
or U469 (N_469,In_674,In_690);
or U470 (N_470,In_888,In_799);
nor U471 (N_471,In_133,In_973);
and U472 (N_472,In_956,In_902);
or U473 (N_473,In_730,In_86);
nand U474 (N_474,In_222,In_707);
or U475 (N_475,In_409,In_223);
nor U476 (N_476,In_31,In_781);
and U477 (N_477,In_592,In_67);
or U478 (N_478,In_701,In_473);
nand U479 (N_479,In_525,In_342);
or U480 (N_480,In_843,In_550);
and U481 (N_481,In_407,In_594);
or U482 (N_482,In_157,In_345);
and U483 (N_483,In_548,In_240);
nand U484 (N_484,In_775,In_205);
or U485 (N_485,In_593,In_841);
nand U486 (N_486,In_135,In_827);
nand U487 (N_487,In_669,In_43);
and U488 (N_488,In_343,In_783);
nand U489 (N_489,In_271,In_897);
and U490 (N_490,In_546,In_368);
and U491 (N_491,In_899,In_484);
nor U492 (N_492,In_760,In_362);
nor U493 (N_493,In_880,In_403);
nand U494 (N_494,In_610,In_351);
nand U495 (N_495,In_810,In_497);
and U496 (N_496,In_79,In_277);
and U497 (N_497,In_260,In_369);
and U498 (N_498,In_879,In_243);
nand U499 (N_499,In_40,In_41);
or U500 (N_500,In_252,In_873);
nor U501 (N_501,In_221,In_836);
and U502 (N_502,In_164,In_789);
or U503 (N_503,In_638,In_360);
nor U504 (N_504,In_699,In_765);
and U505 (N_505,In_514,In_557);
or U506 (N_506,In_970,In_851);
nand U507 (N_507,In_621,In_597);
nor U508 (N_508,In_42,In_442);
nor U509 (N_509,In_141,In_240);
and U510 (N_510,In_964,In_602);
nor U511 (N_511,In_326,In_792);
and U512 (N_512,In_179,In_89);
nand U513 (N_513,In_304,In_794);
and U514 (N_514,In_748,In_89);
or U515 (N_515,In_996,In_892);
nand U516 (N_516,In_184,In_561);
nand U517 (N_517,In_44,In_604);
xor U518 (N_518,In_521,In_409);
nand U519 (N_519,In_162,In_337);
nand U520 (N_520,In_274,In_607);
nor U521 (N_521,In_73,In_326);
nor U522 (N_522,In_854,In_228);
xnor U523 (N_523,In_351,In_20);
and U524 (N_524,In_13,In_187);
and U525 (N_525,In_132,In_192);
or U526 (N_526,In_892,In_448);
and U527 (N_527,In_716,In_476);
nor U528 (N_528,In_846,In_687);
or U529 (N_529,In_474,In_841);
or U530 (N_530,In_214,In_775);
or U531 (N_531,In_775,In_323);
or U532 (N_532,In_418,In_725);
and U533 (N_533,In_585,In_498);
or U534 (N_534,In_733,In_801);
and U535 (N_535,In_304,In_929);
nor U536 (N_536,In_153,In_203);
and U537 (N_537,In_318,In_66);
or U538 (N_538,In_204,In_983);
nand U539 (N_539,In_724,In_391);
nand U540 (N_540,In_236,In_540);
nand U541 (N_541,In_618,In_766);
nor U542 (N_542,In_461,In_927);
nor U543 (N_543,In_42,In_879);
and U544 (N_544,In_696,In_126);
xor U545 (N_545,In_92,In_192);
nor U546 (N_546,In_411,In_724);
xnor U547 (N_547,In_690,In_903);
nor U548 (N_548,In_74,In_29);
nand U549 (N_549,In_756,In_695);
nor U550 (N_550,In_372,In_732);
and U551 (N_551,In_227,In_376);
or U552 (N_552,In_94,In_186);
nor U553 (N_553,In_328,In_286);
and U554 (N_554,In_1,In_843);
and U555 (N_555,In_321,In_342);
nor U556 (N_556,In_702,In_513);
nor U557 (N_557,In_106,In_487);
xor U558 (N_558,In_792,In_285);
nand U559 (N_559,In_293,In_710);
or U560 (N_560,In_305,In_624);
or U561 (N_561,In_341,In_430);
and U562 (N_562,In_986,In_721);
and U563 (N_563,In_47,In_644);
nor U564 (N_564,In_768,In_839);
or U565 (N_565,In_500,In_335);
or U566 (N_566,In_304,In_52);
nor U567 (N_567,In_328,In_235);
nand U568 (N_568,In_567,In_902);
and U569 (N_569,In_515,In_485);
xor U570 (N_570,In_747,In_971);
and U571 (N_571,In_830,In_121);
nor U572 (N_572,In_944,In_513);
and U573 (N_573,In_572,In_516);
or U574 (N_574,In_897,In_930);
or U575 (N_575,In_216,In_410);
nor U576 (N_576,In_55,In_215);
xnor U577 (N_577,In_616,In_533);
nor U578 (N_578,In_323,In_854);
nor U579 (N_579,In_706,In_67);
nor U580 (N_580,In_111,In_576);
or U581 (N_581,In_223,In_914);
nor U582 (N_582,In_65,In_52);
nand U583 (N_583,In_995,In_876);
and U584 (N_584,In_747,In_206);
or U585 (N_585,In_564,In_950);
nor U586 (N_586,In_853,In_840);
nor U587 (N_587,In_340,In_777);
nand U588 (N_588,In_695,In_859);
nor U589 (N_589,In_995,In_109);
and U590 (N_590,In_976,In_31);
and U591 (N_591,In_607,In_29);
or U592 (N_592,In_515,In_60);
nand U593 (N_593,In_239,In_826);
or U594 (N_594,In_700,In_935);
or U595 (N_595,In_239,In_61);
or U596 (N_596,In_827,In_379);
and U597 (N_597,In_781,In_872);
nand U598 (N_598,In_882,In_116);
and U599 (N_599,In_980,In_323);
or U600 (N_600,In_817,In_323);
nand U601 (N_601,In_559,In_182);
nand U602 (N_602,In_241,In_344);
or U603 (N_603,In_536,In_143);
and U604 (N_604,In_214,In_298);
nor U605 (N_605,In_704,In_84);
nand U606 (N_606,In_165,In_460);
and U607 (N_607,In_970,In_740);
or U608 (N_608,In_160,In_672);
and U609 (N_609,In_821,In_857);
and U610 (N_610,In_728,In_635);
nor U611 (N_611,In_219,In_462);
nor U612 (N_612,In_711,In_335);
nand U613 (N_613,In_327,In_76);
and U614 (N_614,In_261,In_643);
nor U615 (N_615,In_938,In_472);
xnor U616 (N_616,In_168,In_282);
nor U617 (N_617,In_924,In_488);
and U618 (N_618,In_635,In_291);
xnor U619 (N_619,In_908,In_530);
and U620 (N_620,In_629,In_260);
and U621 (N_621,In_944,In_530);
nor U622 (N_622,In_944,In_630);
and U623 (N_623,In_503,In_226);
nor U624 (N_624,In_62,In_187);
nand U625 (N_625,In_205,In_883);
nor U626 (N_626,In_312,In_925);
or U627 (N_627,In_309,In_128);
nand U628 (N_628,In_534,In_446);
and U629 (N_629,In_374,In_593);
nor U630 (N_630,In_654,In_510);
and U631 (N_631,In_752,In_881);
nand U632 (N_632,In_772,In_313);
or U633 (N_633,In_342,In_947);
or U634 (N_634,In_648,In_692);
and U635 (N_635,In_271,In_426);
nand U636 (N_636,In_638,In_907);
or U637 (N_637,In_273,In_975);
or U638 (N_638,In_621,In_728);
and U639 (N_639,In_378,In_744);
nand U640 (N_640,In_686,In_85);
or U641 (N_641,In_814,In_218);
nand U642 (N_642,In_616,In_152);
nor U643 (N_643,In_883,In_148);
and U644 (N_644,In_319,In_747);
or U645 (N_645,In_82,In_780);
and U646 (N_646,In_788,In_343);
nand U647 (N_647,In_397,In_271);
nand U648 (N_648,In_526,In_820);
or U649 (N_649,In_455,In_63);
nand U650 (N_650,In_52,In_647);
nand U651 (N_651,In_876,In_247);
and U652 (N_652,In_811,In_32);
nor U653 (N_653,In_361,In_388);
nor U654 (N_654,In_222,In_84);
or U655 (N_655,In_38,In_706);
and U656 (N_656,In_549,In_421);
nor U657 (N_657,In_3,In_283);
or U658 (N_658,In_190,In_667);
nand U659 (N_659,In_171,In_405);
xor U660 (N_660,In_770,In_457);
or U661 (N_661,In_659,In_46);
nor U662 (N_662,In_903,In_9);
and U663 (N_663,In_654,In_657);
nor U664 (N_664,In_119,In_977);
or U665 (N_665,In_272,In_590);
nor U666 (N_666,In_701,In_239);
nor U667 (N_667,In_691,In_836);
nand U668 (N_668,In_399,In_604);
nand U669 (N_669,In_983,In_413);
or U670 (N_670,In_661,In_309);
and U671 (N_671,In_561,In_565);
nor U672 (N_672,In_25,In_566);
nor U673 (N_673,In_792,In_264);
or U674 (N_674,In_119,In_360);
or U675 (N_675,In_719,In_894);
or U676 (N_676,In_655,In_129);
or U677 (N_677,In_472,In_155);
and U678 (N_678,In_599,In_760);
nand U679 (N_679,In_591,In_911);
nor U680 (N_680,In_55,In_931);
xor U681 (N_681,In_763,In_288);
nor U682 (N_682,In_374,In_556);
nand U683 (N_683,In_399,In_350);
and U684 (N_684,In_896,In_406);
and U685 (N_685,In_546,In_963);
nor U686 (N_686,In_841,In_658);
nor U687 (N_687,In_256,In_818);
nand U688 (N_688,In_526,In_511);
nor U689 (N_689,In_983,In_78);
nand U690 (N_690,In_665,In_618);
nor U691 (N_691,In_537,In_405);
nor U692 (N_692,In_265,In_217);
nand U693 (N_693,In_677,In_531);
nor U694 (N_694,In_263,In_842);
nor U695 (N_695,In_367,In_757);
nand U696 (N_696,In_819,In_940);
nand U697 (N_697,In_623,In_999);
or U698 (N_698,In_596,In_759);
nand U699 (N_699,In_919,In_918);
and U700 (N_700,In_929,In_964);
nor U701 (N_701,In_25,In_874);
nor U702 (N_702,In_548,In_639);
and U703 (N_703,In_551,In_832);
and U704 (N_704,In_684,In_686);
xnor U705 (N_705,In_521,In_816);
or U706 (N_706,In_629,In_791);
nand U707 (N_707,In_526,In_819);
or U708 (N_708,In_847,In_465);
or U709 (N_709,In_98,In_357);
and U710 (N_710,In_614,In_180);
nor U711 (N_711,In_208,In_4);
xor U712 (N_712,In_729,In_434);
nand U713 (N_713,In_799,In_720);
nand U714 (N_714,In_982,In_750);
and U715 (N_715,In_317,In_439);
nand U716 (N_716,In_132,In_778);
nand U717 (N_717,In_38,In_613);
nor U718 (N_718,In_353,In_368);
nand U719 (N_719,In_26,In_277);
or U720 (N_720,In_865,In_143);
and U721 (N_721,In_508,In_502);
and U722 (N_722,In_722,In_317);
nand U723 (N_723,In_97,In_657);
nand U724 (N_724,In_61,In_741);
nor U725 (N_725,In_917,In_306);
or U726 (N_726,In_981,In_112);
or U727 (N_727,In_587,In_271);
and U728 (N_728,In_739,In_270);
nor U729 (N_729,In_78,In_472);
nand U730 (N_730,In_841,In_72);
or U731 (N_731,In_733,In_789);
or U732 (N_732,In_420,In_604);
nor U733 (N_733,In_666,In_19);
and U734 (N_734,In_754,In_968);
nor U735 (N_735,In_979,In_946);
and U736 (N_736,In_751,In_956);
and U737 (N_737,In_144,In_781);
or U738 (N_738,In_328,In_306);
or U739 (N_739,In_772,In_78);
or U740 (N_740,In_728,In_690);
nand U741 (N_741,In_903,In_445);
and U742 (N_742,In_650,In_812);
and U743 (N_743,In_555,In_89);
or U744 (N_744,In_441,In_359);
or U745 (N_745,In_644,In_532);
nor U746 (N_746,In_189,In_446);
nor U747 (N_747,In_546,In_405);
and U748 (N_748,In_95,In_336);
nand U749 (N_749,In_988,In_82);
nor U750 (N_750,In_425,In_568);
nor U751 (N_751,In_760,In_247);
and U752 (N_752,In_137,In_773);
nor U753 (N_753,In_45,In_562);
nor U754 (N_754,In_912,In_460);
or U755 (N_755,In_361,In_212);
or U756 (N_756,In_32,In_384);
nor U757 (N_757,In_384,In_587);
nand U758 (N_758,In_474,In_24);
or U759 (N_759,In_754,In_616);
nand U760 (N_760,In_819,In_12);
and U761 (N_761,In_415,In_137);
nor U762 (N_762,In_266,In_206);
or U763 (N_763,In_772,In_669);
and U764 (N_764,In_483,In_319);
nor U765 (N_765,In_429,In_783);
nor U766 (N_766,In_613,In_355);
nand U767 (N_767,In_727,In_45);
nand U768 (N_768,In_741,In_681);
nor U769 (N_769,In_684,In_789);
nand U770 (N_770,In_77,In_100);
nand U771 (N_771,In_287,In_884);
or U772 (N_772,In_119,In_98);
nor U773 (N_773,In_97,In_516);
nand U774 (N_774,In_505,In_526);
or U775 (N_775,In_972,In_940);
nor U776 (N_776,In_661,In_397);
and U777 (N_777,In_7,In_869);
nor U778 (N_778,In_528,In_670);
nor U779 (N_779,In_673,In_935);
nor U780 (N_780,In_229,In_48);
nor U781 (N_781,In_843,In_838);
or U782 (N_782,In_260,In_688);
nor U783 (N_783,In_433,In_744);
nand U784 (N_784,In_862,In_743);
nor U785 (N_785,In_861,In_534);
nor U786 (N_786,In_470,In_201);
nor U787 (N_787,In_103,In_398);
or U788 (N_788,In_115,In_857);
nor U789 (N_789,In_850,In_235);
and U790 (N_790,In_621,In_751);
nand U791 (N_791,In_301,In_396);
or U792 (N_792,In_259,In_703);
nor U793 (N_793,In_560,In_553);
nand U794 (N_794,In_723,In_742);
nor U795 (N_795,In_299,In_990);
or U796 (N_796,In_284,In_872);
nand U797 (N_797,In_679,In_275);
nor U798 (N_798,In_994,In_683);
nand U799 (N_799,In_0,In_84);
and U800 (N_800,In_814,In_291);
nor U801 (N_801,In_243,In_330);
xor U802 (N_802,In_320,In_804);
nand U803 (N_803,In_7,In_130);
or U804 (N_804,In_125,In_863);
nor U805 (N_805,In_438,In_869);
nand U806 (N_806,In_585,In_518);
nor U807 (N_807,In_552,In_283);
or U808 (N_808,In_475,In_270);
nor U809 (N_809,In_460,In_847);
nand U810 (N_810,In_575,In_326);
nor U811 (N_811,In_6,In_681);
nand U812 (N_812,In_579,In_802);
nand U813 (N_813,In_831,In_328);
and U814 (N_814,In_225,In_575);
nand U815 (N_815,In_302,In_417);
nand U816 (N_816,In_466,In_395);
and U817 (N_817,In_31,In_138);
and U818 (N_818,In_592,In_916);
and U819 (N_819,In_972,In_586);
nor U820 (N_820,In_552,In_920);
or U821 (N_821,In_224,In_544);
nand U822 (N_822,In_506,In_924);
nand U823 (N_823,In_207,In_441);
nor U824 (N_824,In_623,In_116);
nor U825 (N_825,In_317,In_398);
nor U826 (N_826,In_150,In_779);
or U827 (N_827,In_964,In_583);
xor U828 (N_828,In_63,In_775);
nand U829 (N_829,In_719,In_582);
nand U830 (N_830,In_974,In_898);
and U831 (N_831,In_175,In_101);
and U832 (N_832,In_908,In_208);
or U833 (N_833,In_202,In_498);
nor U834 (N_834,In_502,In_38);
and U835 (N_835,In_529,In_935);
nor U836 (N_836,In_623,In_279);
or U837 (N_837,In_914,In_41);
and U838 (N_838,In_515,In_353);
nand U839 (N_839,In_45,In_340);
or U840 (N_840,In_14,In_140);
and U841 (N_841,In_808,In_561);
nand U842 (N_842,In_738,In_747);
nor U843 (N_843,In_315,In_675);
and U844 (N_844,In_640,In_821);
nand U845 (N_845,In_273,In_656);
or U846 (N_846,In_231,In_529);
or U847 (N_847,In_886,In_997);
nand U848 (N_848,In_39,In_828);
nand U849 (N_849,In_558,In_289);
nor U850 (N_850,In_962,In_377);
nor U851 (N_851,In_133,In_577);
nand U852 (N_852,In_354,In_200);
nor U853 (N_853,In_571,In_257);
and U854 (N_854,In_230,In_305);
or U855 (N_855,In_956,In_995);
or U856 (N_856,In_245,In_67);
or U857 (N_857,In_665,In_549);
or U858 (N_858,In_1,In_912);
nand U859 (N_859,In_750,In_220);
xnor U860 (N_860,In_398,In_899);
and U861 (N_861,In_646,In_653);
nor U862 (N_862,In_395,In_433);
nand U863 (N_863,In_367,In_248);
xnor U864 (N_864,In_786,In_531);
nor U865 (N_865,In_922,In_718);
or U866 (N_866,In_124,In_866);
nand U867 (N_867,In_272,In_984);
or U868 (N_868,In_29,In_318);
nand U869 (N_869,In_279,In_951);
or U870 (N_870,In_657,In_105);
or U871 (N_871,In_365,In_651);
and U872 (N_872,In_897,In_671);
nand U873 (N_873,In_484,In_110);
nand U874 (N_874,In_570,In_770);
and U875 (N_875,In_247,In_899);
or U876 (N_876,In_560,In_166);
and U877 (N_877,In_921,In_831);
nor U878 (N_878,In_922,In_910);
and U879 (N_879,In_183,In_386);
or U880 (N_880,In_872,In_467);
or U881 (N_881,In_585,In_812);
nor U882 (N_882,In_515,In_663);
and U883 (N_883,In_826,In_633);
nand U884 (N_884,In_427,In_508);
and U885 (N_885,In_363,In_735);
and U886 (N_886,In_374,In_389);
and U887 (N_887,In_203,In_274);
nor U888 (N_888,In_345,In_756);
nand U889 (N_889,In_513,In_436);
nand U890 (N_890,In_112,In_97);
nor U891 (N_891,In_528,In_792);
and U892 (N_892,In_279,In_967);
nor U893 (N_893,In_15,In_908);
and U894 (N_894,In_55,In_784);
xnor U895 (N_895,In_256,In_825);
or U896 (N_896,In_686,In_450);
nand U897 (N_897,In_135,In_878);
nand U898 (N_898,In_671,In_759);
or U899 (N_899,In_961,In_226);
nor U900 (N_900,In_27,In_454);
and U901 (N_901,In_726,In_126);
and U902 (N_902,In_582,In_293);
or U903 (N_903,In_127,In_266);
and U904 (N_904,In_732,In_42);
nand U905 (N_905,In_91,In_999);
and U906 (N_906,In_643,In_105);
nor U907 (N_907,In_320,In_598);
nor U908 (N_908,In_347,In_759);
nor U909 (N_909,In_783,In_517);
nand U910 (N_910,In_772,In_566);
or U911 (N_911,In_454,In_648);
and U912 (N_912,In_850,In_781);
nor U913 (N_913,In_685,In_768);
nand U914 (N_914,In_432,In_167);
nor U915 (N_915,In_651,In_33);
and U916 (N_916,In_950,In_818);
nand U917 (N_917,In_922,In_618);
and U918 (N_918,In_94,In_66);
and U919 (N_919,In_938,In_980);
xor U920 (N_920,In_503,In_855);
nand U921 (N_921,In_732,In_533);
and U922 (N_922,In_696,In_405);
and U923 (N_923,In_160,In_403);
nand U924 (N_924,In_258,In_760);
nand U925 (N_925,In_575,In_878);
and U926 (N_926,In_932,In_277);
nor U927 (N_927,In_125,In_43);
nand U928 (N_928,In_691,In_895);
nand U929 (N_929,In_805,In_168);
and U930 (N_930,In_768,In_212);
nor U931 (N_931,In_827,In_377);
or U932 (N_932,In_661,In_198);
nand U933 (N_933,In_868,In_712);
nor U934 (N_934,In_819,In_241);
or U935 (N_935,In_398,In_329);
nand U936 (N_936,In_44,In_131);
nor U937 (N_937,In_991,In_718);
or U938 (N_938,In_748,In_395);
and U939 (N_939,In_175,In_928);
nand U940 (N_940,In_551,In_915);
nor U941 (N_941,In_304,In_157);
nor U942 (N_942,In_436,In_841);
nand U943 (N_943,In_173,In_88);
nor U944 (N_944,In_9,In_59);
and U945 (N_945,In_468,In_875);
nor U946 (N_946,In_512,In_222);
or U947 (N_947,In_386,In_108);
xnor U948 (N_948,In_793,In_877);
and U949 (N_949,In_144,In_727);
and U950 (N_950,In_717,In_716);
and U951 (N_951,In_94,In_146);
nor U952 (N_952,In_686,In_582);
nor U953 (N_953,In_66,In_485);
nor U954 (N_954,In_577,In_99);
or U955 (N_955,In_709,In_820);
or U956 (N_956,In_506,In_470);
nand U957 (N_957,In_719,In_967);
or U958 (N_958,In_21,In_680);
and U959 (N_959,In_465,In_520);
and U960 (N_960,In_64,In_689);
and U961 (N_961,In_100,In_442);
nor U962 (N_962,In_343,In_679);
and U963 (N_963,In_793,In_26);
or U964 (N_964,In_362,In_865);
nand U965 (N_965,In_903,In_401);
nand U966 (N_966,In_679,In_608);
nor U967 (N_967,In_897,In_606);
nand U968 (N_968,In_174,In_719);
nand U969 (N_969,In_255,In_211);
nor U970 (N_970,In_878,In_933);
nand U971 (N_971,In_939,In_10);
or U972 (N_972,In_3,In_465);
or U973 (N_973,In_464,In_902);
nand U974 (N_974,In_693,In_584);
xnor U975 (N_975,In_335,In_643);
or U976 (N_976,In_433,In_270);
nor U977 (N_977,In_24,In_669);
or U978 (N_978,In_718,In_712);
or U979 (N_979,In_456,In_754);
nor U980 (N_980,In_257,In_483);
or U981 (N_981,In_822,In_402);
and U982 (N_982,In_851,In_828);
and U983 (N_983,In_300,In_281);
and U984 (N_984,In_22,In_992);
nand U985 (N_985,In_359,In_258);
and U986 (N_986,In_39,In_139);
nand U987 (N_987,In_656,In_877);
and U988 (N_988,In_148,In_740);
nand U989 (N_989,In_336,In_121);
nand U990 (N_990,In_77,In_170);
or U991 (N_991,In_17,In_951);
nor U992 (N_992,In_248,In_906);
and U993 (N_993,In_724,In_305);
and U994 (N_994,In_989,In_456);
nor U995 (N_995,In_560,In_588);
and U996 (N_996,In_728,In_969);
or U997 (N_997,In_678,In_213);
or U998 (N_998,In_167,In_198);
nand U999 (N_999,In_552,In_22);
nor U1000 (N_1000,In_840,In_684);
and U1001 (N_1001,In_570,In_152);
and U1002 (N_1002,In_283,In_108);
nand U1003 (N_1003,In_825,In_646);
nor U1004 (N_1004,In_905,In_76);
nor U1005 (N_1005,In_446,In_872);
or U1006 (N_1006,In_397,In_872);
and U1007 (N_1007,In_760,In_821);
nor U1008 (N_1008,In_778,In_629);
or U1009 (N_1009,In_812,In_158);
nor U1010 (N_1010,In_252,In_467);
nor U1011 (N_1011,In_989,In_40);
or U1012 (N_1012,In_577,In_770);
and U1013 (N_1013,In_661,In_767);
and U1014 (N_1014,In_577,In_554);
nor U1015 (N_1015,In_706,In_8);
nor U1016 (N_1016,In_133,In_417);
and U1017 (N_1017,In_942,In_502);
or U1018 (N_1018,In_853,In_33);
and U1019 (N_1019,In_784,In_905);
nor U1020 (N_1020,In_566,In_590);
nor U1021 (N_1021,In_870,In_981);
or U1022 (N_1022,In_505,In_81);
or U1023 (N_1023,In_789,In_981);
nand U1024 (N_1024,In_526,In_165);
and U1025 (N_1025,In_990,In_947);
and U1026 (N_1026,In_359,In_885);
or U1027 (N_1027,In_500,In_613);
or U1028 (N_1028,In_291,In_952);
and U1029 (N_1029,In_19,In_928);
nand U1030 (N_1030,In_418,In_406);
nand U1031 (N_1031,In_453,In_59);
or U1032 (N_1032,In_111,In_944);
or U1033 (N_1033,In_491,In_685);
or U1034 (N_1034,In_145,In_665);
or U1035 (N_1035,In_542,In_493);
nand U1036 (N_1036,In_807,In_799);
and U1037 (N_1037,In_816,In_647);
xor U1038 (N_1038,In_446,In_732);
or U1039 (N_1039,In_812,In_999);
and U1040 (N_1040,In_765,In_353);
and U1041 (N_1041,In_140,In_38);
nand U1042 (N_1042,In_153,In_550);
nor U1043 (N_1043,In_894,In_0);
and U1044 (N_1044,In_259,In_911);
and U1045 (N_1045,In_404,In_111);
and U1046 (N_1046,In_184,In_714);
and U1047 (N_1047,In_218,In_738);
nand U1048 (N_1048,In_484,In_24);
or U1049 (N_1049,In_415,In_952);
nor U1050 (N_1050,In_626,In_879);
or U1051 (N_1051,In_838,In_620);
and U1052 (N_1052,In_807,In_357);
nor U1053 (N_1053,In_322,In_409);
nand U1054 (N_1054,In_79,In_197);
and U1055 (N_1055,In_684,In_699);
nand U1056 (N_1056,In_3,In_79);
nand U1057 (N_1057,In_182,In_56);
and U1058 (N_1058,In_858,In_98);
nor U1059 (N_1059,In_766,In_365);
nand U1060 (N_1060,In_720,In_801);
and U1061 (N_1061,In_852,In_754);
nor U1062 (N_1062,In_141,In_839);
nand U1063 (N_1063,In_282,In_993);
or U1064 (N_1064,In_193,In_965);
or U1065 (N_1065,In_676,In_747);
nor U1066 (N_1066,In_3,In_586);
or U1067 (N_1067,In_725,In_942);
nor U1068 (N_1068,In_88,In_175);
nand U1069 (N_1069,In_931,In_493);
and U1070 (N_1070,In_174,In_116);
and U1071 (N_1071,In_246,In_945);
or U1072 (N_1072,In_264,In_914);
and U1073 (N_1073,In_932,In_87);
and U1074 (N_1074,In_483,In_796);
nor U1075 (N_1075,In_100,In_179);
or U1076 (N_1076,In_336,In_588);
nor U1077 (N_1077,In_730,In_61);
or U1078 (N_1078,In_321,In_924);
nor U1079 (N_1079,In_919,In_142);
nand U1080 (N_1080,In_367,In_361);
or U1081 (N_1081,In_802,In_475);
and U1082 (N_1082,In_983,In_560);
and U1083 (N_1083,In_995,In_632);
and U1084 (N_1084,In_878,In_983);
and U1085 (N_1085,In_494,In_957);
nor U1086 (N_1086,In_734,In_518);
nand U1087 (N_1087,In_221,In_714);
nor U1088 (N_1088,In_406,In_910);
xnor U1089 (N_1089,In_717,In_462);
nor U1090 (N_1090,In_296,In_876);
nand U1091 (N_1091,In_128,In_495);
nor U1092 (N_1092,In_845,In_363);
xnor U1093 (N_1093,In_389,In_18);
nor U1094 (N_1094,In_810,In_635);
or U1095 (N_1095,In_736,In_460);
or U1096 (N_1096,In_655,In_668);
or U1097 (N_1097,In_978,In_589);
nor U1098 (N_1098,In_510,In_336);
and U1099 (N_1099,In_6,In_830);
nor U1100 (N_1100,In_486,In_338);
and U1101 (N_1101,In_992,In_610);
nor U1102 (N_1102,In_371,In_53);
nand U1103 (N_1103,In_859,In_515);
and U1104 (N_1104,In_41,In_26);
and U1105 (N_1105,In_71,In_492);
or U1106 (N_1106,In_58,In_862);
nor U1107 (N_1107,In_34,In_627);
or U1108 (N_1108,In_553,In_529);
and U1109 (N_1109,In_981,In_539);
nor U1110 (N_1110,In_973,In_52);
or U1111 (N_1111,In_602,In_751);
and U1112 (N_1112,In_53,In_244);
or U1113 (N_1113,In_393,In_917);
nor U1114 (N_1114,In_748,In_112);
and U1115 (N_1115,In_311,In_756);
and U1116 (N_1116,In_600,In_852);
or U1117 (N_1117,In_86,In_414);
and U1118 (N_1118,In_281,In_993);
nand U1119 (N_1119,In_50,In_755);
and U1120 (N_1120,In_547,In_853);
nor U1121 (N_1121,In_664,In_535);
or U1122 (N_1122,In_245,In_62);
nand U1123 (N_1123,In_845,In_15);
nand U1124 (N_1124,In_421,In_166);
or U1125 (N_1125,In_308,In_580);
and U1126 (N_1126,In_631,In_822);
nand U1127 (N_1127,In_682,In_305);
nor U1128 (N_1128,In_629,In_798);
nand U1129 (N_1129,In_949,In_538);
or U1130 (N_1130,In_726,In_928);
nor U1131 (N_1131,In_210,In_906);
or U1132 (N_1132,In_34,In_450);
nor U1133 (N_1133,In_261,In_538);
and U1134 (N_1134,In_478,In_692);
or U1135 (N_1135,In_54,In_518);
and U1136 (N_1136,In_858,In_439);
and U1137 (N_1137,In_695,In_70);
nor U1138 (N_1138,In_674,In_112);
or U1139 (N_1139,In_642,In_480);
nand U1140 (N_1140,In_882,In_933);
nor U1141 (N_1141,In_151,In_737);
and U1142 (N_1142,In_8,In_458);
nor U1143 (N_1143,In_730,In_287);
nand U1144 (N_1144,In_983,In_816);
nor U1145 (N_1145,In_982,In_35);
or U1146 (N_1146,In_634,In_124);
nor U1147 (N_1147,In_409,In_144);
or U1148 (N_1148,In_556,In_375);
nor U1149 (N_1149,In_883,In_345);
and U1150 (N_1150,In_688,In_49);
nand U1151 (N_1151,In_913,In_536);
or U1152 (N_1152,In_879,In_208);
and U1153 (N_1153,In_943,In_444);
xnor U1154 (N_1154,In_918,In_728);
and U1155 (N_1155,In_15,In_311);
and U1156 (N_1156,In_963,In_955);
and U1157 (N_1157,In_239,In_891);
nand U1158 (N_1158,In_956,In_997);
nor U1159 (N_1159,In_558,In_320);
and U1160 (N_1160,In_702,In_919);
or U1161 (N_1161,In_562,In_862);
or U1162 (N_1162,In_151,In_999);
nand U1163 (N_1163,In_305,In_684);
xor U1164 (N_1164,In_340,In_496);
nor U1165 (N_1165,In_522,In_734);
or U1166 (N_1166,In_306,In_950);
nor U1167 (N_1167,In_688,In_269);
nand U1168 (N_1168,In_96,In_965);
nor U1169 (N_1169,In_237,In_335);
or U1170 (N_1170,In_379,In_250);
or U1171 (N_1171,In_631,In_96);
nand U1172 (N_1172,In_683,In_493);
nor U1173 (N_1173,In_690,In_491);
and U1174 (N_1174,In_812,In_2);
nand U1175 (N_1175,In_960,In_546);
nor U1176 (N_1176,In_941,In_826);
or U1177 (N_1177,In_870,In_68);
nand U1178 (N_1178,In_503,In_589);
and U1179 (N_1179,In_762,In_724);
and U1180 (N_1180,In_78,In_618);
nand U1181 (N_1181,In_396,In_151);
or U1182 (N_1182,In_28,In_133);
and U1183 (N_1183,In_398,In_158);
nor U1184 (N_1184,In_801,In_718);
nand U1185 (N_1185,In_232,In_940);
or U1186 (N_1186,In_90,In_278);
or U1187 (N_1187,In_705,In_769);
and U1188 (N_1188,In_833,In_161);
or U1189 (N_1189,In_288,In_29);
nand U1190 (N_1190,In_496,In_213);
nor U1191 (N_1191,In_323,In_434);
or U1192 (N_1192,In_628,In_983);
or U1193 (N_1193,In_87,In_844);
nor U1194 (N_1194,In_143,In_208);
xor U1195 (N_1195,In_604,In_996);
nand U1196 (N_1196,In_393,In_233);
and U1197 (N_1197,In_808,In_576);
nand U1198 (N_1198,In_247,In_253);
and U1199 (N_1199,In_138,In_63);
and U1200 (N_1200,In_386,In_696);
or U1201 (N_1201,In_695,In_885);
or U1202 (N_1202,In_359,In_44);
and U1203 (N_1203,In_216,In_524);
nor U1204 (N_1204,In_3,In_838);
nor U1205 (N_1205,In_541,In_588);
nand U1206 (N_1206,In_632,In_641);
nand U1207 (N_1207,In_86,In_301);
nand U1208 (N_1208,In_239,In_574);
nor U1209 (N_1209,In_665,In_747);
or U1210 (N_1210,In_403,In_276);
or U1211 (N_1211,In_53,In_817);
nand U1212 (N_1212,In_982,In_629);
nand U1213 (N_1213,In_272,In_940);
nand U1214 (N_1214,In_732,In_913);
or U1215 (N_1215,In_73,In_550);
xor U1216 (N_1216,In_692,In_60);
nand U1217 (N_1217,In_37,In_370);
and U1218 (N_1218,In_609,In_747);
nor U1219 (N_1219,In_816,In_166);
or U1220 (N_1220,In_904,In_217);
nand U1221 (N_1221,In_659,In_150);
and U1222 (N_1222,In_257,In_538);
and U1223 (N_1223,In_255,In_922);
and U1224 (N_1224,In_756,In_64);
xor U1225 (N_1225,In_850,In_644);
and U1226 (N_1226,In_644,In_792);
or U1227 (N_1227,In_861,In_503);
and U1228 (N_1228,In_928,In_529);
and U1229 (N_1229,In_808,In_498);
nand U1230 (N_1230,In_784,In_177);
and U1231 (N_1231,In_566,In_163);
nand U1232 (N_1232,In_139,In_620);
or U1233 (N_1233,In_345,In_493);
or U1234 (N_1234,In_879,In_598);
nor U1235 (N_1235,In_427,In_47);
or U1236 (N_1236,In_860,In_52);
nand U1237 (N_1237,In_751,In_201);
and U1238 (N_1238,In_801,In_361);
and U1239 (N_1239,In_553,In_523);
or U1240 (N_1240,In_24,In_741);
xnor U1241 (N_1241,In_736,In_422);
xor U1242 (N_1242,In_511,In_547);
and U1243 (N_1243,In_902,In_165);
nand U1244 (N_1244,In_329,In_840);
and U1245 (N_1245,In_704,In_286);
and U1246 (N_1246,In_373,In_468);
and U1247 (N_1247,In_388,In_71);
nand U1248 (N_1248,In_876,In_366);
or U1249 (N_1249,In_24,In_393);
or U1250 (N_1250,In_515,In_591);
and U1251 (N_1251,In_51,In_165);
or U1252 (N_1252,In_333,In_376);
nand U1253 (N_1253,In_873,In_771);
nor U1254 (N_1254,In_314,In_885);
and U1255 (N_1255,In_355,In_123);
nand U1256 (N_1256,In_25,In_421);
or U1257 (N_1257,In_948,In_876);
nor U1258 (N_1258,In_760,In_366);
nand U1259 (N_1259,In_756,In_979);
or U1260 (N_1260,In_611,In_966);
nand U1261 (N_1261,In_632,In_128);
or U1262 (N_1262,In_914,In_691);
nor U1263 (N_1263,In_26,In_66);
nor U1264 (N_1264,In_479,In_361);
and U1265 (N_1265,In_56,In_857);
or U1266 (N_1266,In_536,In_191);
and U1267 (N_1267,In_338,In_787);
and U1268 (N_1268,In_148,In_696);
and U1269 (N_1269,In_207,In_80);
and U1270 (N_1270,In_164,In_573);
and U1271 (N_1271,In_528,In_171);
nor U1272 (N_1272,In_608,In_756);
nor U1273 (N_1273,In_821,In_132);
or U1274 (N_1274,In_801,In_898);
nor U1275 (N_1275,In_946,In_272);
or U1276 (N_1276,In_496,In_521);
and U1277 (N_1277,In_782,In_516);
or U1278 (N_1278,In_544,In_827);
nor U1279 (N_1279,In_85,In_721);
nor U1280 (N_1280,In_729,In_169);
or U1281 (N_1281,In_60,In_51);
and U1282 (N_1282,In_181,In_334);
and U1283 (N_1283,In_228,In_474);
nor U1284 (N_1284,In_20,In_365);
xnor U1285 (N_1285,In_635,In_516);
nand U1286 (N_1286,In_65,In_402);
and U1287 (N_1287,In_585,In_391);
and U1288 (N_1288,In_769,In_244);
nand U1289 (N_1289,In_30,In_160);
and U1290 (N_1290,In_830,In_649);
nor U1291 (N_1291,In_566,In_237);
nand U1292 (N_1292,In_823,In_751);
nand U1293 (N_1293,In_429,In_781);
or U1294 (N_1294,In_962,In_978);
or U1295 (N_1295,In_60,In_980);
nand U1296 (N_1296,In_234,In_664);
nor U1297 (N_1297,In_215,In_685);
or U1298 (N_1298,In_30,In_924);
nor U1299 (N_1299,In_177,In_877);
or U1300 (N_1300,In_426,In_16);
nand U1301 (N_1301,In_135,In_838);
nand U1302 (N_1302,In_957,In_383);
or U1303 (N_1303,In_347,In_515);
nor U1304 (N_1304,In_91,In_69);
nor U1305 (N_1305,In_629,In_610);
nor U1306 (N_1306,In_909,In_428);
nand U1307 (N_1307,In_86,In_136);
nor U1308 (N_1308,In_210,In_959);
and U1309 (N_1309,In_628,In_607);
nand U1310 (N_1310,In_499,In_162);
and U1311 (N_1311,In_470,In_2);
and U1312 (N_1312,In_455,In_749);
or U1313 (N_1313,In_554,In_711);
or U1314 (N_1314,In_200,In_176);
or U1315 (N_1315,In_851,In_12);
nand U1316 (N_1316,In_431,In_718);
nor U1317 (N_1317,In_867,In_99);
or U1318 (N_1318,In_365,In_556);
nor U1319 (N_1319,In_480,In_318);
and U1320 (N_1320,In_258,In_110);
nor U1321 (N_1321,In_951,In_36);
or U1322 (N_1322,In_941,In_331);
nor U1323 (N_1323,In_686,In_221);
nand U1324 (N_1324,In_980,In_45);
xnor U1325 (N_1325,In_63,In_773);
nand U1326 (N_1326,In_766,In_249);
or U1327 (N_1327,In_552,In_786);
or U1328 (N_1328,In_236,In_989);
nor U1329 (N_1329,In_493,In_592);
nor U1330 (N_1330,In_910,In_355);
or U1331 (N_1331,In_455,In_541);
nand U1332 (N_1332,In_503,In_670);
and U1333 (N_1333,In_309,In_416);
nor U1334 (N_1334,In_322,In_161);
and U1335 (N_1335,In_401,In_905);
and U1336 (N_1336,In_858,In_947);
or U1337 (N_1337,In_214,In_97);
nor U1338 (N_1338,In_294,In_77);
nand U1339 (N_1339,In_917,In_946);
nor U1340 (N_1340,In_887,In_425);
or U1341 (N_1341,In_330,In_852);
nor U1342 (N_1342,In_312,In_134);
nand U1343 (N_1343,In_566,In_805);
nand U1344 (N_1344,In_582,In_103);
nand U1345 (N_1345,In_84,In_369);
nor U1346 (N_1346,In_50,In_692);
nor U1347 (N_1347,In_138,In_602);
nand U1348 (N_1348,In_130,In_538);
and U1349 (N_1349,In_765,In_223);
nand U1350 (N_1350,In_935,In_655);
and U1351 (N_1351,In_769,In_127);
or U1352 (N_1352,In_227,In_841);
nand U1353 (N_1353,In_113,In_554);
or U1354 (N_1354,In_995,In_886);
nand U1355 (N_1355,In_719,In_307);
or U1356 (N_1356,In_291,In_859);
nor U1357 (N_1357,In_339,In_472);
or U1358 (N_1358,In_877,In_440);
nand U1359 (N_1359,In_657,In_882);
nor U1360 (N_1360,In_138,In_676);
nand U1361 (N_1361,In_672,In_152);
or U1362 (N_1362,In_795,In_139);
nor U1363 (N_1363,In_981,In_656);
or U1364 (N_1364,In_311,In_483);
nor U1365 (N_1365,In_630,In_753);
nor U1366 (N_1366,In_179,In_718);
or U1367 (N_1367,In_441,In_669);
nand U1368 (N_1368,In_710,In_316);
or U1369 (N_1369,In_626,In_877);
and U1370 (N_1370,In_816,In_787);
nand U1371 (N_1371,In_829,In_987);
nand U1372 (N_1372,In_335,In_915);
or U1373 (N_1373,In_470,In_51);
nor U1374 (N_1374,In_729,In_782);
and U1375 (N_1375,In_639,In_937);
nor U1376 (N_1376,In_806,In_455);
nor U1377 (N_1377,In_479,In_608);
xnor U1378 (N_1378,In_600,In_638);
or U1379 (N_1379,In_947,In_23);
nand U1380 (N_1380,In_231,In_661);
nand U1381 (N_1381,In_130,In_401);
xor U1382 (N_1382,In_781,In_462);
or U1383 (N_1383,In_318,In_838);
and U1384 (N_1384,In_790,In_609);
nor U1385 (N_1385,In_353,In_188);
nor U1386 (N_1386,In_723,In_399);
or U1387 (N_1387,In_289,In_171);
and U1388 (N_1388,In_293,In_874);
nand U1389 (N_1389,In_856,In_546);
or U1390 (N_1390,In_481,In_53);
or U1391 (N_1391,In_797,In_315);
or U1392 (N_1392,In_626,In_565);
nor U1393 (N_1393,In_823,In_723);
and U1394 (N_1394,In_631,In_513);
xnor U1395 (N_1395,In_45,In_731);
nand U1396 (N_1396,In_581,In_755);
and U1397 (N_1397,In_782,In_310);
nor U1398 (N_1398,In_774,In_87);
nand U1399 (N_1399,In_491,In_622);
nor U1400 (N_1400,In_850,In_363);
and U1401 (N_1401,In_318,In_223);
nand U1402 (N_1402,In_194,In_641);
and U1403 (N_1403,In_15,In_446);
nand U1404 (N_1404,In_739,In_722);
nor U1405 (N_1405,In_557,In_184);
or U1406 (N_1406,In_174,In_102);
nor U1407 (N_1407,In_48,In_111);
or U1408 (N_1408,In_732,In_492);
nor U1409 (N_1409,In_979,In_419);
nor U1410 (N_1410,In_763,In_543);
or U1411 (N_1411,In_135,In_681);
or U1412 (N_1412,In_181,In_290);
xnor U1413 (N_1413,In_455,In_127);
or U1414 (N_1414,In_706,In_559);
nor U1415 (N_1415,In_809,In_796);
nor U1416 (N_1416,In_647,In_863);
or U1417 (N_1417,In_370,In_518);
nand U1418 (N_1418,In_217,In_346);
nor U1419 (N_1419,In_702,In_427);
or U1420 (N_1420,In_962,In_132);
nor U1421 (N_1421,In_394,In_342);
nor U1422 (N_1422,In_22,In_942);
nand U1423 (N_1423,In_654,In_387);
or U1424 (N_1424,In_233,In_714);
nor U1425 (N_1425,In_252,In_158);
nor U1426 (N_1426,In_456,In_235);
nor U1427 (N_1427,In_290,In_925);
and U1428 (N_1428,In_374,In_411);
nor U1429 (N_1429,In_164,In_489);
nand U1430 (N_1430,In_32,In_37);
nand U1431 (N_1431,In_682,In_320);
and U1432 (N_1432,In_825,In_490);
nand U1433 (N_1433,In_174,In_696);
nor U1434 (N_1434,In_779,In_205);
or U1435 (N_1435,In_743,In_772);
nor U1436 (N_1436,In_756,In_592);
xnor U1437 (N_1437,In_762,In_833);
nor U1438 (N_1438,In_544,In_591);
and U1439 (N_1439,In_808,In_555);
or U1440 (N_1440,In_606,In_224);
nand U1441 (N_1441,In_51,In_948);
or U1442 (N_1442,In_473,In_657);
nor U1443 (N_1443,In_197,In_769);
or U1444 (N_1444,In_478,In_137);
or U1445 (N_1445,In_165,In_643);
nand U1446 (N_1446,In_427,In_573);
or U1447 (N_1447,In_832,In_494);
nand U1448 (N_1448,In_815,In_179);
nand U1449 (N_1449,In_232,In_684);
or U1450 (N_1450,In_274,In_223);
or U1451 (N_1451,In_287,In_303);
nor U1452 (N_1452,In_231,In_124);
xnor U1453 (N_1453,In_14,In_204);
nand U1454 (N_1454,In_658,In_790);
and U1455 (N_1455,In_860,In_534);
or U1456 (N_1456,In_429,In_396);
nand U1457 (N_1457,In_224,In_86);
nand U1458 (N_1458,In_311,In_240);
nor U1459 (N_1459,In_100,In_482);
nand U1460 (N_1460,In_663,In_253);
nor U1461 (N_1461,In_637,In_745);
nand U1462 (N_1462,In_564,In_120);
nor U1463 (N_1463,In_611,In_398);
nand U1464 (N_1464,In_900,In_345);
and U1465 (N_1465,In_129,In_628);
or U1466 (N_1466,In_361,In_825);
or U1467 (N_1467,In_538,In_115);
and U1468 (N_1468,In_270,In_870);
or U1469 (N_1469,In_134,In_419);
nand U1470 (N_1470,In_710,In_481);
nor U1471 (N_1471,In_246,In_82);
xor U1472 (N_1472,In_500,In_729);
and U1473 (N_1473,In_206,In_644);
nor U1474 (N_1474,In_705,In_701);
nand U1475 (N_1475,In_509,In_964);
or U1476 (N_1476,In_725,In_195);
and U1477 (N_1477,In_5,In_183);
or U1478 (N_1478,In_959,In_117);
nand U1479 (N_1479,In_94,In_427);
nand U1480 (N_1480,In_390,In_933);
nor U1481 (N_1481,In_513,In_619);
xnor U1482 (N_1482,In_374,In_459);
nor U1483 (N_1483,In_697,In_617);
or U1484 (N_1484,In_607,In_638);
nand U1485 (N_1485,In_219,In_249);
nor U1486 (N_1486,In_766,In_742);
and U1487 (N_1487,In_231,In_60);
nand U1488 (N_1488,In_567,In_70);
nor U1489 (N_1489,In_954,In_611);
and U1490 (N_1490,In_478,In_63);
nand U1491 (N_1491,In_543,In_276);
xnor U1492 (N_1492,In_560,In_382);
nor U1493 (N_1493,In_747,In_751);
and U1494 (N_1494,In_699,In_139);
nor U1495 (N_1495,In_47,In_930);
nor U1496 (N_1496,In_684,In_951);
or U1497 (N_1497,In_766,In_967);
or U1498 (N_1498,In_636,In_708);
xor U1499 (N_1499,In_520,In_882);
and U1500 (N_1500,In_984,In_641);
nand U1501 (N_1501,In_826,In_725);
nand U1502 (N_1502,In_694,In_227);
or U1503 (N_1503,In_318,In_297);
and U1504 (N_1504,In_385,In_615);
nand U1505 (N_1505,In_839,In_506);
or U1506 (N_1506,In_44,In_304);
nor U1507 (N_1507,In_5,In_286);
or U1508 (N_1508,In_485,In_446);
nand U1509 (N_1509,In_763,In_915);
and U1510 (N_1510,In_882,In_833);
and U1511 (N_1511,In_837,In_996);
nand U1512 (N_1512,In_276,In_33);
nand U1513 (N_1513,In_320,In_214);
nand U1514 (N_1514,In_280,In_42);
nand U1515 (N_1515,In_993,In_373);
or U1516 (N_1516,In_683,In_119);
nand U1517 (N_1517,In_967,In_609);
and U1518 (N_1518,In_688,In_410);
and U1519 (N_1519,In_160,In_155);
nand U1520 (N_1520,In_50,In_630);
nor U1521 (N_1521,In_20,In_289);
nor U1522 (N_1522,In_799,In_553);
or U1523 (N_1523,In_153,In_855);
or U1524 (N_1524,In_528,In_37);
nand U1525 (N_1525,In_717,In_225);
nand U1526 (N_1526,In_29,In_650);
and U1527 (N_1527,In_93,In_663);
nand U1528 (N_1528,In_61,In_432);
or U1529 (N_1529,In_550,In_457);
or U1530 (N_1530,In_936,In_187);
nand U1531 (N_1531,In_137,In_979);
and U1532 (N_1532,In_269,In_945);
nand U1533 (N_1533,In_687,In_629);
or U1534 (N_1534,In_542,In_497);
and U1535 (N_1535,In_108,In_729);
or U1536 (N_1536,In_254,In_820);
or U1537 (N_1537,In_958,In_743);
and U1538 (N_1538,In_172,In_343);
nor U1539 (N_1539,In_563,In_521);
or U1540 (N_1540,In_256,In_441);
or U1541 (N_1541,In_58,In_158);
nor U1542 (N_1542,In_344,In_6);
nand U1543 (N_1543,In_973,In_278);
or U1544 (N_1544,In_636,In_993);
nand U1545 (N_1545,In_143,In_304);
nand U1546 (N_1546,In_295,In_579);
and U1547 (N_1547,In_848,In_471);
nand U1548 (N_1548,In_105,In_745);
or U1549 (N_1549,In_787,In_199);
nor U1550 (N_1550,In_344,In_729);
and U1551 (N_1551,In_597,In_37);
or U1552 (N_1552,In_853,In_798);
or U1553 (N_1553,In_818,In_865);
and U1554 (N_1554,In_97,In_973);
nand U1555 (N_1555,In_359,In_331);
and U1556 (N_1556,In_657,In_426);
and U1557 (N_1557,In_322,In_215);
or U1558 (N_1558,In_286,In_18);
nor U1559 (N_1559,In_502,In_780);
or U1560 (N_1560,In_996,In_447);
nand U1561 (N_1561,In_711,In_606);
and U1562 (N_1562,In_417,In_726);
and U1563 (N_1563,In_457,In_531);
nor U1564 (N_1564,In_267,In_991);
and U1565 (N_1565,In_232,In_333);
nor U1566 (N_1566,In_50,In_516);
and U1567 (N_1567,In_120,In_278);
and U1568 (N_1568,In_508,In_753);
nor U1569 (N_1569,In_80,In_903);
and U1570 (N_1570,In_48,In_290);
and U1571 (N_1571,In_603,In_183);
nand U1572 (N_1572,In_655,In_660);
or U1573 (N_1573,In_518,In_661);
nor U1574 (N_1574,In_531,In_583);
and U1575 (N_1575,In_350,In_568);
nand U1576 (N_1576,In_350,In_525);
and U1577 (N_1577,In_241,In_940);
or U1578 (N_1578,In_848,In_263);
nor U1579 (N_1579,In_654,In_64);
or U1580 (N_1580,In_805,In_159);
and U1581 (N_1581,In_875,In_63);
and U1582 (N_1582,In_721,In_505);
and U1583 (N_1583,In_907,In_478);
and U1584 (N_1584,In_265,In_884);
nor U1585 (N_1585,In_769,In_961);
and U1586 (N_1586,In_645,In_777);
nand U1587 (N_1587,In_67,In_780);
and U1588 (N_1588,In_524,In_415);
nor U1589 (N_1589,In_520,In_741);
nor U1590 (N_1590,In_433,In_507);
or U1591 (N_1591,In_637,In_715);
nor U1592 (N_1592,In_920,In_77);
xor U1593 (N_1593,In_317,In_402);
nand U1594 (N_1594,In_454,In_685);
nand U1595 (N_1595,In_2,In_827);
and U1596 (N_1596,In_237,In_202);
and U1597 (N_1597,In_889,In_305);
nand U1598 (N_1598,In_803,In_645);
xor U1599 (N_1599,In_91,In_684);
or U1600 (N_1600,In_849,In_162);
nand U1601 (N_1601,In_199,In_3);
nand U1602 (N_1602,In_721,In_249);
or U1603 (N_1603,In_660,In_471);
nand U1604 (N_1604,In_299,In_654);
nor U1605 (N_1605,In_735,In_471);
xor U1606 (N_1606,In_193,In_868);
nor U1607 (N_1607,In_519,In_49);
or U1608 (N_1608,In_11,In_173);
or U1609 (N_1609,In_505,In_533);
nand U1610 (N_1610,In_219,In_624);
and U1611 (N_1611,In_671,In_605);
nor U1612 (N_1612,In_580,In_663);
or U1613 (N_1613,In_558,In_184);
nor U1614 (N_1614,In_525,In_951);
or U1615 (N_1615,In_431,In_405);
nand U1616 (N_1616,In_631,In_28);
nand U1617 (N_1617,In_681,In_977);
and U1618 (N_1618,In_340,In_215);
nand U1619 (N_1619,In_169,In_885);
nand U1620 (N_1620,In_451,In_439);
xnor U1621 (N_1621,In_642,In_703);
nor U1622 (N_1622,In_788,In_737);
nor U1623 (N_1623,In_765,In_41);
and U1624 (N_1624,In_400,In_843);
nand U1625 (N_1625,In_916,In_837);
nor U1626 (N_1626,In_305,In_787);
nand U1627 (N_1627,In_192,In_375);
and U1628 (N_1628,In_638,In_581);
nand U1629 (N_1629,In_605,In_961);
nand U1630 (N_1630,In_779,In_620);
nor U1631 (N_1631,In_384,In_38);
nand U1632 (N_1632,In_852,In_294);
and U1633 (N_1633,In_998,In_976);
or U1634 (N_1634,In_89,In_285);
or U1635 (N_1635,In_252,In_776);
nand U1636 (N_1636,In_525,In_748);
or U1637 (N_1637,In_548,In_728);
xnor U1638 (N_1638,In_472,In_816);
nor U1639 (N_1639,In_81,In_46);
nor U1640 (N_1640,In_88,In_31);
and U1641 (N_1641,In_455,In_49);
nand U1642 (N_1642,In_495,In_447);
and U1643 (N_1643,In_493,In_492);
or U1644 (N_1644,In_853,In_740);
nand U1645 (N_1645,In_951,In_600);
nor U1646 (N_1646,In_177,In_693);
nand U1647 (N_1647,In_203,In_752);
nand U1648 (N_1648,In_143,In_105);
nor U1649 (N_1649,In_915,In_580);
nor U1650 (N_1650,In_46,In_202);
or U1651 (N_1651,In_439,In_170);
and U1652 (N_1652,In_401,In_664);
or U1653 (N_1653,In_996,In_762);
nand U1654 (N_1654,In_35,In_364);
and U1655 (N_1655,In_246,In_472);
nand U1656 (N_1656,In_593,In_343);
nor U1657 (N_1657,In_283,In_893);
and U1658 (N_1658,In_44,In_704);
or U1659 (N_1659,In_586,In_86);
nand U1660 (N_1660,In_974,In_736);
nor U1661 (N_1661,In_740,In_215);
nand U1662 (N_1662,In_627,In_497);
nor U1663 (N_1663,In_246,In_858);
or U1664 (N_1664,In_38,In_885);
nand U1665 (N_1665,In_347,In_557);
or U1666 (N_1666,In_114,In_960);
and U1667 (N_1667,In_266,In_764);
nor U1668 (N_1668,In_115,In_122);
and U1669 (N_1669,In_56,In_894);
and U1670 (N_1670,In_308,In_29);
nor U1671 (N_1671,In_566,In_903);
nand U1672 (N_1672,In_32,In_195);
and U1673 (N_1673,In_454,In_595);
or U1674 (N_1674,In_617,In_666);
nor U1675 (N_1675,In_476,In_135);
and U1676 (N_1676,In_796,In_145);
nor U1677 (N_1677,In_65,In_129);
and U1678 (N_1678,In_247,In_237);
or U1679 (N_1679,In_928,In_545);
nand U1680 (N_1680,In_254,In_701);
nand U1681 (N_1681,In_185,In_218);
nand U1682 (N_1682,In_199,In_808);
nor U1683 (N_1683,In_646,In_349);
or U1684 (N_1684,In_580,In_300);
nor U1685 (N_1685,In_173,In_455);
or U1686 (N_1686,In_646,In_366);
nand U1687 (N_1687,In_725,In_234);
or U1688 (N_1688,In_535,In_246);
nand U1689 (N_1689,In_634,In_217);
or U1690 (N_1690,In_492,In_755);
nor U1691 (N_1691,In_379,In_377);
nor U1692 (N_1692,In_210,In_934);
nand U1693 (N_1693,In_302,In_676);
or U1694 (N_1694,In_933,In_85);
nand U1695 (N_1695,In_567,In_202);
nor U1696 (N_1696,In_108,In_440);
nand U1697 (N_1697,In_233,In_126);
and U1698 (N_1698,In_284,In_637);
xnor U1699 (N_1699,In_976,In_946);
nor U1700 (N_1700,In_528,In_198);
or U1701 (N_1701,In_756,In_802);
nor U1702 (N_1702,In_622,In_601);
nand U1703 (N_1703,In_669,In_302);
nor U1704 (N_1704,In_924,In_169);
nand U1705 (N_1705,In_929,In_410);
and U1706 (N_1706,In_694,In_10);
and U1707 (N_1707,In_368,In_192);
nand U1708 (N_1708,In_145,In_113);
nor U1709 (N_1709,In_635,In_720);
and U1710 (N_1710,In_57,In_702);
or U1711 (N_1711,In_717,In_630);
nand U1712 (N_1712,In_106,In_59);
and U1713 (N_1713,In_67,In_400);
or U1714 (N_1714,In_14,In_946);
nor U1715 (N_1715,In_190,In_812);
nand U1716 (N_1716,In_345,In_453);
and U1717 (N_1717,In_313,In_399);
or U1718 (N_1718,In_842,In_865);
nor U1719 (N_1719,In_555,In_857);
nor U1720 (N_1720,In_368,In_2);
and U1721 (N_1721,In_573,In_5);
or U1722 (N_1722,In_618,In_232);
or U1723 (N_1723,In_28,In_431);
and U1724 (N_1724,In_382,In_773);
nor U1725 (N_1725,In_48,In_883);
or U1726 (N_1726,In_525,In_259);
nand U1727 (N_1727,In_456,In_605);
or U1728 (N_1728,In_423,In_800);
nor U1729 (N_1729,In_372,In_393);
nor U1730 (N_1730,In_29,In_732);
nand U1731 (N_1731,In_687,In_566);
nor U1732 (N_1732,In_516,In_418);
nand U1733 (N_1733,In_271,In_932);
or U1734 (N_1734,In_186,In_832);
nand U1735 (N_1735,In_610,In_438);
nand U1736 (N_1736,In_952,In_927);
nor U1737 (N_1737,In_299,In_439);
or U1738 (N_1738,In_629,In_630);
or U1739 (N_1739,In_118,In_270);
or U1740 (N_1740,In_778,In_242);
nor U1741 (N_1741,In_965,In_239);
nand U1742 (N_1742,In_981,In_152);
and U1743 (N_1743,In_316,In_156);
nand U1744 (N_1744,In_348,In_239);
nor U1745 (N_1745,In_648,In_2);
and U1746 (N_1746,In_736,In_91);
nand U1747 (N_1747,In_307,In_410);
nand U1748 (N_1748,In_565,In_559);
nand U1749 (N_1749,In_21,In_473);
nor U1750 (N_1750,In_287,In_297);
and U1751 (N_1751,In_458,In_558);
and U1752 (N_1752,In_689,In_171);
nor U1753 (N_1753,In_863,In_644);
nand U1754 (N_1754,In_801,In_550);
or U1755 (N_1755,In_367,In_722);
nor U1756 (N_1756,In_438,In_932);
nor U1757 (N_1757,In_728,In_303);
and U1758 (N_1758,In_72,In_552);
and U1759 (N_1759,In_178,In_654);
nand U1760 (N_1760,In_348,In_808);
or U1761 (N_1761,In_41,In_422);
nand U1762 (N_1762,In_910,In_948);
nor U1763 (N_1763,In_632,In_793);
and U1764 (N_1764,In_447,In_907);
or U1765 (N_1765,In_356,In_202);
nor U1766 (N_1766,In_813,In_999);
nand U1767 (N_1767,In_237,In_505);
and U1768 (N_1768,In_116,In_123);
and U1769 (N_1769,In_480,In_157);
and U1770 (N_1770,In_970,In_897);
and U1771 (N_1771,In_806,In_769);
and U1772 (N_1772,In_931,In_922);
xor U1773 (N_1773,In_372,In_131);
and U1774 (N_1774,In_615,In_691);
nand U1775 (N_1775,In_563,In_687);
or U1776 (N_1776,In_422,In_423);
nor U1777 (N_1777,In_695,In_836);
and U1778 (N_1778,In_649,In_937);
nand U1779 (N_1779,In_717,In_688);
nand U1780 (N_1780,In_547,In_908);
and U1781 (N_1781,In_522,In_816);
and U1782 (N_1782,In_578,In_615);
xnor U1783 (N_1783,In_844,In_239);
nor U1784 (N_1784,In_731,In_445);
and U1785 (N_1785,In_75,In_430);
nand U1786 (N_1786,In_874,In_395);
nand U1787 (N_1787,In_702,In_266);
and U1788 (N_1788,In_564,In_927);
nand U1789 (N_1789,In_956,In_119);
nor U1790 (N_1790,In_64,In_518);
and U1791 (N_1791,In_209,In_258);
and U1792 (N_1792,In_185,In_764);
or U1793 (N_1793,In_691,In_807);
nor U1794 (N_1794,In_875,In_433);
nor U1795 (N_1795,In_599,In_794);
and U1796 (N_1796,In_366,In_269);
nand U1797 (N_1797,In_643,In_93);
and U1798 (N_1798,In_260,In_804);
or U1799 (N_1799,In_559,In_103);
nor U1800 (N_1800,In_592,In_939);
nor U1801 (N_1801,In_974,In_691);
nand U1802 (N_1802,In_690,In_632);
nor U1803 (N_1803,In_371,In_912);
and U1804 (N_1804,In_121,In_253);
or U1805 (N_1805,In_801,In_457);
or U1806 (N_1806,In_534,In_473);
or U1807 (N_1807,In_619,In_842);
nor U1808 (N_1808,In_252,In_919);
nor U1809 (N_1809,In_789,In_935);
nand U1810 (N_1810,In_621,In_249);
nand U1811 (N_1811,In_204,In_781);
and U1812 (N_1812,In_351,In_980);
nor U1813 (N_1813,In_184,In_542);
and U1814 (N_1814,In_134,In_904);
nand U1815 (N_1815,In_220,In_286);
or U1816 (N_1816,In_751,In_863);
and U1817 (N_1817,In_944,In_823);
or U1818 (N_1818,In_789,In_480);
or U1819 (N_1819,In_912,In_217);
nor U1820 (N_1820,In_109,In_745);
nor U1821 (N_1821,In_98,In_525);
nor U1822 (N_1822,In_751,In_569);
and U1823 (N_1823,In_269,In_800);
and U1824 (N_1824,In_546,In_845);
xor U1825 (N_1825,In_251,In_753);
nand U1826 (N_1826,In_765,In_292);
or U1827 (N_1827,In_503,In_741);
or U1828 (N_1828,In_952,In_280);
xor U1829 (N_1829,In_17,In_521);
xnor U1830 (N_1830,In_89,In_577);
nand U1831 (N_1831,In_885,In_60);
and U1832 (N_1832,In_371,In_482);
and U1833 (N_1833,In_860,In_518);
nor U1834 (N_1834,In_438,In_714);
nand U1835 (N_1835,In_730,In_396);
nand U1836 (N_1836,In_464,In_575);
or U1837 (N_1837,In_485,In_511);
nand U1838 (N_1838,In_158,In_38);
nand U1839 (N_1839,In_458,In_531);
and U1840 (N_1840,In_904,In_533);
nand U1841 (N_1841,In_83,In_235);
nand U1842 (N_1842,In_53,In_974);
and U1843 (N_1843,In_129,In_92);
nand U1844 (N_1844,In_392,In_705);
nand U1845 (N_1845,In_12,In_361);
nor U1846 (N_1846,In_104,In_499);
or U1847 (N_1847,In_174,In_538);
xor U1848 (N_1848,In_960,In_856);
and U1849 (N_1849,In_63,In_941);
and U1850 (N_1850,In_536,In_961);
nor U1851 (N_1851,In_370,In_485);
nand U1852 (N_1852,In_47,In_977);
nor U1853 (N_1853,In_677,In_556);
nor U1854 (N_1854,In_111,In_562);
and U1855 (N_1855,In_33,In_901);
nand U1856 (N_1856,In_96,In_243);
and U1857 (N_1857,In_125,In_134);
nand U1858 (N_1858,In_579,In_166);
nand U1859 (N_1859,In_110,In_444);
or U1860 (N_1860,In_369,In_885);
or U1861 (N_1861,In_896,In_82);
and U1862 (N_1862,In_327,In_388);
nand U1863 (N_1863,In_975,In_78);
nor U1864 (N_1864,In_739,In_870);
nand U1865 (N_1865,In_552,In_716);
or U1866 (N_1866,In_332,In_876);
and U1867 (N_1867,In_67,In_657);
and U1868 (N_1868,In_329,In_121);
nand U1869 (N_1869,In_573,In_672);
nor U1870 (N_1870,In_933,In_520);
nand U1871 (N_1871,In_105,In_29);
xnor U1872 (N_1872,In_443,In_572);
or U1873 (N_1873,In_33,In_333);
and U1874 (N_1874,In_562,In_183);
and U1875 (N_1875,In_981,In_755);
and U1876 (N_1876,In_268,In_994);
nor U1877 (N_1877,In_470,In_474);
or U1878 (N_1878,In_935,In_517);
nand U1879 (N_1879,In_11,In_698);
nand U1880 (N_1880,In_138,In_844);
nor U1881 (N_1881,In_692,In_452);
nand U1882 (N_1882,In_179,In_299);
and U1883 (N_1883,In_936,In_924);
nor U1884 (N_1884,In_869,In_730);
and U1885 (N_1885,In_833,In_259);
nand U1886 (N_1886,In_145,In_965);
nand U1887 (N_1887,In_570,In_669);
nand U1888 (N_1888,In_185,In_711);
or U1889 (N_1889,In_264,In_1);
or U1890 (N_1890,In_196,In_222);
and U1891 (N_1891,In_270,In_640);
and U1892 (N_1892,In_698,In_962);
nor U1893 (N_1893,In_642,In_599);
nor U1894 (N_1894,In_280,In_134);
nor U1895 (N_1895,In_806,In_518);
and U1896 (N_1896,In_733,In_966);
or U1897 (N_1897,In_509,In_933);
nand U1898 (N_1898,In_489,In_817);
and U1899 (N_1899,In_798,In_259);
or U1900 (N_1900,In_26,In_122);
and U1901 (N_1901,In_74,In_794);
and U1902 (N_1902,In_684,In_452);
nand U1903 (N_1903,In_540,In_674);
nand U1904 (N_1904,In_664,In_759);
or U1905 (N_1905,In_956,In_577);
nand U1906 (N_1906,In_212,In_70);
nand U1907 (N_1907,In_806,In_314);
nor U1908 (N_1908,In_326,In_36);
and U1909 (N_1909,In_378,In_948);
nand U1910 (N_1910,In_540,In_569);
nand U1911 (N_1911,In_603,In_160);
nor U1912 (N_1912,In_293,In_494);
nor U1913 (N_1913,In_726,In_616);
nand U1914 (N_1914,In_601,In_441);
and U1915 (N_1915,In_669,In_304);
and U1916 (N_1916,In_783,In_201);
or U1917 (N_1917,In_422,In_846);
or U1918 (N_1918,In_143,In_45);
xor U1919 (N_1919,In_414,In_662);
nand U1920 (N_1920,In_321,In_819);
nor U1921 (N_1921,In_253,In_711);
nor U1922 (N_1922,In_287,In_43);
nand U1923 (N_1923,In_950,In_763);
nor U1924 (N_1924,In_201,In_599);
and U1925 (N_1925,In_482,In_269);
nand U1926 (N_1926,In_941,In_590);
nand U1927 (N_1927,In_393,In_722);
nor U1928 (N_1928,In_987,In_606);
or U1929 (N_1929,In_71,In_270);
or U1930 (N_1930,In_971,In_705);
or U1931 (N_1931,In_530,In_355);
or U1932 (N_1932,In_431,In_748);
or U1933 (N_1933,In_695,In_328);
and U1934 (N_1934,In_378,In_309);
and U1935 (N_1935,In_92,In_993);
nor U1936 (N_1936,In_649,In_978);
xor U1937 (N_1937,In_525,In_563);
or U1938 (N_1938,In_802,In_36);
nand U1939 (N_1939,In_57,In_303);
nand U1940 (N_1940,In_828,In_145);
nor U1941 (N_1941,In_774,In_869);
nor U1942 (N_1942,In_314,In_591);
or U1943 (N_1943,In_77,In_536);
or U1944 (N_1944,In_862,In_690);
and U1945 (N_1945,In_572,In_383);
or U1946 (N_1946,In_10,In_925);
or U1947 (N_1947,In_793,In_547);
nand U1948 (N_1948,In_791,In_484);
nor U1949 (N_1949,In_971,In_179);
nor U1950 (N_1950,In_755,In_966);
and U1951 (N_1951,In_337,In_211);
and U1952 (N_1952,In_264,In_725);
or U1953 (N_1953,In_3,In_940);
nand U1954 (N_1954,In_413,In_130);
nor U1955 (N_1955,In_212,In_627);
or U1956 (N_1956,In_155,In_252);
nor U1957 (N_1957,In_245,In_928);
and U1958 (N_1958,In_61,In_171);
or U1959 (N_1959,In_128,In_771);
xor U1960 (N_1960,In_145,In_189);
and U1961 (N_1961,In_674,In_937);
nor U1962 (N_1962,In_684,In_890);
nand U1963 (N_1963,In_248,In_510);
nand U1964 (N_1964,In_783,In_956);
and U1965 (N_1965,In_840,In_551);
and U1966 (N_1966,In_10,In_186);
or U1967 (N_1967,In_885,In_276);
or U1968 (N_1968,In_124,In_333);
xnor U1969 (N_1969,In_115,In_669);
nor U1970 (N_1970,In_415,In_848);
nor U1971 (N_1971,In_396,In_407);
nor U1972 (N_1972,In_994,In_166);
or U1973 (N_1973,In_916,In_248);
or U1974 (N_1974,In_389,In_60);
nor U1975 (N_1975,In_781,In_384);
and U1976 (N_1976,In_912,In_377);
nand U1977 (N_1977,In_40,In_876);
nor U1978 (N_1978,In_271,In_14);
or U1979 (N_1979,In_511,In_785);
and U1980 (N_1980,In_27,In_825);
and U1981 (N_1981,In_995,In_479);
nand U1982 (N_1982,In_244,In_473);
nor U1983 (N_1983,In_917,In_910);
or U1984 (N_1984,In_110,In_841);
nand U1985 (N_1985,In_399,In_690);
nand U1986 (N_1986,In_630,In_833);
nor U1987 (N_1987,In_28,In_683);
nand U1988 (N_1988,In_589,In_471);
nor U1989 (N_1989,In_306,In_59);
or U1990 (N_1990,In_201,In_303);
and U1991 (N_1991,In_625,In_45);
nor U1992 (N_1992,In_607,In_561);
nor U1993 (N_1993,In_376,In_791);
nor U1994 (N_1994,In_698,In_208);
and U1995 (N_1995,In_232,In_713);
or U1996 (N_1996,In_173,In_436);
or U1997 (N_1997,In_8,In_132);
nand U1998 (N_1998,In_76,In_966);
or U1999 (N_1999,In_513,In_520);
nand U2000 (N_2000,In_814,In_123);
or U2001 (N_2001,In_613,In_356);
and U2002 (N_2002,In_811,In_668);
and U2003 (N_2003,In_515,In_308);
or U2004 (N_2004,In_868,In_348);
and U2005 (N_2005,In_790,In_804);
nand U2006 (N_2006,In_159,In_533);
nor U2007 (N_2007,In_626,In_779);
nand U2008 (N_2008,In_980,In_582);
or U2009 (N_2009,In_349,In_731);
or U2010 (N_2010,In_241,In_213);
or U2011 (N_2011,In_343,In_324);
and U2012 (N_2012,In_449,In_848);
nor U2013 (N_2013,In_253,In_778);
and U2014 (N_2014,In_286,In_298);
or U2015 (N_2015,In_672,In_921);
nand U2016 (N_2016,In_341,In_210);
nand U2017 (N_2017,In_630,In_631);
or U2018 (N_2018,In_818,In_634);
nand U2019 (N_2019,In_389,In_190);
nand U2020 (N_2020,In_757,In_514);
or U2021 (N_2021,In_437,In_700);
nor U2022 (N_2022,In_367,In_451);
or U2023 (N_2023,In_642,In_221);
nor U2024 (N_2024,In_851,In_896);
or U2025 (N_2025,In_6,In_691);
nor U2026 (N_2026,In_247,In_219);
nand U2027 (N_2027,In_95,In_724);
or U2028 (N_2028,In_616,In_991);
nand U2029 (N_2029,In_192,In_396);
and U2030 (N_2030,In_649,In_229);
nand U2031 (N_2031,In_843,In_390);
nor U2032 (N_2032,In_271,In_291);
xnor U2033 (N_2033,In_0,In_33);
and U2034 (N_2034,In_341,In_808);
nand U2035 (N_2035,In_846,In_83);
or U2036 (N_2036,In_232,In_513);
nor U2037 (N_2037,In_818,In_466);
and U2038 (N_2038,In_365,In_788);
nand U2039 (N_2039,In_932,In_4);
nor U2040 (N_2040,In_795,In_514);
nor U2041 (N_2041,In_9,In_282);
or U2042 (N_2042,In_547,In_566);
or U2043 (N_2043,In_655,In_468);
nor U2044 (N_2044,In_460,In_465);
or U2045 (N_2045,In_864,In_36);
and U2046 (N_2046,In_583,In_349);
nand U2047 (N_2047,In_490,In_122);
nand U2048 (N_2048,In_549,In_321);
nand U2049 (N_2049,In_453,In_992);
xnor U2050 (N_2050,In_872,In_439);
or U2051 (N_2051,In_599,In_826);
nor U2052 (N_2052,In_67,In_128);
and U2053 (N_2053,In_916,In_68);
or U2054 (N_2054,In_11,In_763);
and U2055 (N_2055,In_710,In_741);
and U2056 (N_2056,In_527,In_442);
or U2057 (N_2057,In_3,In_556);
xor U2058 (N_2058,In_107,In_388);
or U2059 (N_2059,In_953,In_716);
nand U2060 (N_2060,In_981,In_360);
nor U2061 (N_2061,In_70,In_656);
or U2062 (N_2062,In_772,In_798);
nor U2063 (N_2063,In_754,In_887);
nand U2064 (N_2064,In_846,In_952);
or U2065 (N_2065,In_734,In_883);
or U2066 (N_2066,In_579,In_397);
nand U2067 (N_2067,In_206,In_830);
or U2068 (N_2068,In_645,In_755);
and U2069 (N_2069,In_300,In_900);
and U2070 (N_2070,In_716,In_681);
nand U2071 (N_2071,In_6,In_504);
and U2072 (N_2072,In_988,In_837);
and U2073 (N_2073,In_698,In_769);
or U2074 (N_2074,In_963,In_207);
nand U2075 (N_2075,In_817,In_218);
nor U2076 (N_2076,In_880,In_563);
and U2077 (N_2077,In_244,In_653);
nand U2078 (N_2078,In_63,In_134);
nand U2079 (N_2079,In_229,In_517);
nor U2080 (N_2080,In_674,In_859);
nor U2081 (N_2081,In_767,In_713);
or U2082 (N_2082,In_825,In_126);
nor U2083 (N_2083,In_523,In_692);
or U2084 (N_2084,In_281,In_117);
or U2085 (N_2085,In_33,In_457);
nand U2086 (N_2086,In_10,In_181);
and U2087 (N_2087,In_548,In_549);
or U2088 (N_2088,In_712,In_415);
or U2089 (N_2089,In_133,In_698);
nor U2090 (N_2090,In_339,In_572);
nor U2091 (N_2091,In_981,In_762);
or U2092 (N_2092,In_544,In_930);
nor U2093 (N_2093,In_564,In_845);
and U2094 (N_2094,In_504,In_443);
and U2095 (N_2095,In_340,In_475);
nand U2096 (N_2096,In_583,In_83);
nor U2097 (N_2097,In_761,In_257);
and U2098 (N_2098,In_109,In_722);
nand U2099 (N_2099,In_747,In_488);
and U2100 (N_2100,In_139,In_306);
and U2101 (N_2101,In_854,In_241);
and U2102 (N_2102,In_805,In_745);
and U2103 (N_2103,In_901,In_398);
and U2104 (N_2104,In_218,In_613);
nand U2105 (N_2105,In_712,In_843);
and U2106 (N_2106,In_0,In_46);
and U2107 (N_2107,In_184,In_369);
and U2108 (N_2108,In_232,In_768);
nor U2109 (N_2109,In_841,In_839);
or U2110 (N_2110,In_326,In_986);
nor U2111 (N_2111,In_264,In_627);
nor U2112 (N_2112,In_434,In_154);
and U2113 (N_2113,In_261,In_627);
nand U2114 (N_2114,In_102,In_349);
and U2115 (N_2115,In_402,In_311);
or U2116 (N_2116,In_598,In_695);
nor U2117 (N_2117,In_303,In_598);
nor U2118 (N_2118,In_519,In_138);
and U2119 (N_2119,In_770,In_474);
xnor U2120 (N_2120,In_505,In_777);
nor U2121 (N_2121,In_124,In_739);
and U2122 (N_2122,In_33,In_719);
xor U2123 (N_2123,In_211,In_283);
nor U2124 (N_2124,In_870,In_482);
and U2125 (N_2125,In_601,In_730);
or U2126 (N_2126,In_114,In_313);
or U2127 (N_2127,In_194,In_518);
nor U2128 (N_2128,In_285,In_245);
or U2129 (N_2129,In_292,In_158);
and U2130 (N_2130,In_159,In_668);
nor U2131 (N_2131,In_92,In_649);
or U2132 (N_2132,In_750,In_103);
nand U2133 (N_2133,In_433,In_225);
nand U2134 (N_2134,In_260,In_816);
nor U2135 (N_2135,In_435,In_109);
or U2136 (N_2136,In_974,In_720);
nor U2137 (N_2137,In_642,In_770);
or U2138 (N_2138,In_511,In_572);
or U2139 (N_2139,In_91,In_306);
nand U2140 (N_2140,In_681,In_410);
or U2141 (N_2141,In_157,In_309);
nand U2142 (N_2142,In_258,In_345);
nor U2143 (N_2143,In_602,In_615);
nand U2144 (N_2144,In_226,In_310);
or U2145 (N_2145,In_25,In_828);
nor U2146 (N_2146,In_384,In_208);
or U2147 (N_2147,In_582,In_653);
nand U2148 (N_2148,In_351,In_311);
and U2149 (N_2149,In_461,In_457);
or U2150 (N_2150,In_756,In_707);
nor U2151 (N_2151,In_650,In_698);
and U2152 (N_2152,In_825,In_451);
xnor U2153 (N_2153,In_734,In_856);
nand U2154 (N_2154,In_751,In_969);
nand U2155 (N_2155,In_565,In_608);
and U2156 (N_2156,In_229,In_820);
nor U2157 (N_2157,In_598,In_657);
nand U2158 (N_2158,In_726,In_263);
nand U2159 (N_2159,In_758,In_461);
nor U2160 (N_2160,In_528,In_684);
or U2161 (N_2161,In_134,In_522);
nand U2162 (N_2162,In_440,In_175);
nor U2163 (N_2163,In_539,In_615);
nor U2164 (N_2164,In_291,In_379);
nand U2165 (N_2165,In_493,In_844);
nor U2166 (N_2166,In_897,In_479);
and U2167 (N_2167,In_264,In_970);
nand U2168 (N_2168,In_416,In_136);
nor U2169 (N_2169,In_679,In_347);
nor U2170 (N_2170,In_11,In_609);
or U2171 (N_2171,In_317,In_653);
or U2172 (N_2172,In_551,In_151);
nor U2173 (N_2173,In_863,In_907);
and U2174 (N_2174,In_214,In_265);
nand U2175 (N_2175,In_831,In_612);
and U2176 (N_2176,In_792,In_730);
nor U2177 (N_2177,In_921,In_898);
and U2178 (N_2178,In_127,In_448);
nand U2179 (N_2179,In_892,In_833);
nand U2180 (N_2180,In_525,In_565);
or U2181 (N_2181,In_198,In_985);
nand U2182 (N_2182,In_32,In_337);
nand U2183 (N_2183,In_353,In_317);
and U2184 (N_2184,In_668,In_152);
nor U2185 (N_2185,In_857,In_921);
and U2186 (N_2186,In_427,In_659);
nor U2187 (N_2187,In_308,In_678);
and U2188 (N_2188,In_607,In_975);
or U2189 (N_2189,In_124,In_606);
nor U2190 (N_2190,In_408,In_400);
nand U2191 (N_2191,In_124,In_895);
nand U2192 (N_2192,In_375,In_118);
and U2193 (N_2193,In_861,In_524);
xnor U2194 (N_2194,In_592,In_933);
nand U2195 (N_2195,In_316,In_914);
nand U2196 (N_2196,In_836,In_420);
nand U2197 (N_2197,In_440,In_245);
and U2198 (N_2198,In_618,In_321);
or U2199 (N_2199,In_508,In_421);
nor U2200 (N_2200,In_940,In_458);
and U2201 (N_2201,In_138,In_947);
nand U2202 (N_2202,In_69,In_422);
nand U2203 (N_2203,In_854,In_41);
nand U2204 (N_2204,In_342,In_970);
and U2205 (N_2205,In_542,In_444);
and U2206 (N_2206,In_529,In_76);
nand U2207 (N_2207,In_72,In_933);
nand U2208 (N_2208,In_102,In_183);
nand U2209 (N_2209,In_904,In_578);
or U2210 (N_2210,In_679,In_956);
nand U2211 (N_2211,In_410,In_232);
nor U2212 (N_2212,In_32,In_724);
nor U2213 (N_2213,In_376,In_291);
and U2214 (N_2214,In_935,In_954);
nand U2215 (N_2215,In_621,In_188);
or U2216 (N_2216,In_381,In_495);
and U2217 (N_2217,In_205,In_656);
or U2218 (N_2218,In_923,In_195);
nand U2219 (N_2219,In_882,In_794);
or U2220 (N_2220,In_704,In_393);
nand U2221 (N_2221,In_714,In_627);
and U2222 (N_2222,In_927,In_185);
or U2223 (N_2223,In_873,In_760);
nand U2224 (N_2224,In_316,In_138);
or U2225 (N_2225,In_70,In_561);
and U2226 (N_2226,In_125,In_154);
nor U2227 (N_2227,In_491,In_351);
xor U2228 (N_2228,In_75,In_109);
nand U2229 (N_2229,In_14,In_755);
and U2230 (N_2230,In_898,In_265);
nand U2231 (N_2231,In_366,In_282);
or U2232 (N_2232,In_220,In_521);
nor U2233 (N_2233,In_476,In_23);
nor U2234 (N_2234,In_735,In_366);
or U2235 (N_2235,In_254,In_881);
nor U2236 (N_2236,In_825,In_679);
or U2237 (N_2237,In_32,In_513);
xor U2238 (N_2238,In_29,In_564);
or U2239 (N_2239,In_12,In_750);
nand U2240 (N_2240,In_371,In_500);
nor U2241 (N_2241,In_101,In_328);
or U2242 (N_2242,In_960,In_198);
nand U2243 (N_2243,In_216,In_368);
or U2244 (N_2244,In_346,In_55);
and U2245 (N_2245,In_38,In_277);
nand U2246 (N_2246,In_680,In_754);
nand U2247 (N_2247,In_200,In_104);
and U2248 (N_2248,In_723,In_720);
and U2249 (N_2249,In_15,In_774);
nand U2250 (N_2250,In_335,In_401);
or U2251 (N_2251,In_170,In_171);
or U2252 (N_2252,In_159,In_829);
and U2253 (N_2253,In_43,In_446);
and U2254 (N_2254,In_703,In_268);
and U2255 (N_2255,In_611,In_542);
nand U2256 (N_2256,In_469,In_272);
and U2257 (N_2257,In_545,In_455);
nor U2258 (N_2258,In_355,In_663);
or U2259 (N_2259,In_35,In_15);
and U2260 (N_2260,In_40,In_84);
nor U2261 (N_2261,In_448,In_259);
and U2262 (N_2262,In_452,In_813);
and U2263 (N_2263,In_912,In_319);
or U2264 (N_2264,In_618,In_464);
or U2265 (N_2265,In_592,In_862);
nor U2266 (N_2266,In_178,In_40);
nand U2267 (N_2267,In_147,In_88);
nor U2268 (N_2268,In_121,In_715);
or U2269 (N_2269,In_584,In_385);
or U2270 (N_2270,In_732,In_669);
nor U2271 (N_2271,In_410,In_378);
and U2272 (N_2272,In_362,In_460);
or U2273 (N_2273,In_382,In_76);
or U2274 (N_2274,In_86,In_105);
xor U2275 (N_2275,In_764,In_886);
and U2276 (N_2276,In_114,In_631);
nor U2277 (N_2277,In_125,In_503);
nand U2278 (N_2278,In_566,In_166);
or U2279 (N_2279,In_688,In_24);
nor U2280 (N_2280,In_711,In_546);
nand U2281 (N_2281,In_514,In_87);
or U2282 (N_2282,In_473,In_845);
or U2283 (N_2283,In_586,In_851);
nand U2284 (N_2284,In_295,In_69);
nand U2285 (N_2285,In_31,In_912);
and U2286 (N_2286,In_430,In_424);
and U2287 (N_2287,In_764,In_202);
nor U2288 (N_2288,In_942,In_151);
nand U2289 (N_2289,In_277,In_448);
nand U2290 (N_2290,In_997,In_186);
nor U2291 (N_2291,In_410,In_60);
and U2292 (N_2292,In_723,In_568);
nor U2293 (N_2293,In_303,In_297);
nor U2294 (N_2294,In_442,In_360);
and U2295 (N_2295,In_986,In_840);
and U2296 (N_2296,In_230,In_42);
nand U2297 (N_2297,In_641,In_771);
nor U2298 (N_2298,In_545,In_624);
and U2299 (N_2299,In_395,In_41);
nand U2300 (N_2300,In_936,In_149);
nor U2301 (N_2301,In_843,In_680);
nand U2302 (N_2302,In_77,In_503);
or U2303 (N_2303,In_734,In_793);
nand U2304 (N_2304,In_275,In_689);
and U2305 (N_2305,In_443,In_370);
or U2306 (N_2306,In_451,In_274);
nand U2307 (N_2307,In_72,In_399);
xnor U2308 (N_2308,In_802,In_311);
and U2309 (N_2309,In_655,In_993);
or U2310 (N_2310,In_617,In_368);
nand U2311 (N_2311,In_463,In_695);
or U2312 (N_2312,In_355,In_650);
or U2313 (N_2313,In_504,In_836);
nand U2314 (N_2314,In_922,In_992);
or U2315 (N_2315,In_975,In_717);
and U2316 (N_2316,In_574,In_885);
or U2317 (N_2317,In_523,In_386);
or U2318 (N_2318,In_61,In_311);
nor U2319 (N_2319,In_121,In_376);
and U2320 (N_2320,In_147,In_311);
or U2321 (N_2321,In_668,In_548);
nor U2322 (N_2322,In_319,In_601);
nor U2323 (N_2323,In_561,In_212);
nor U2324 (N_2324,In_710,In_112);
nor U2325 (N_2325,In_358,In_650);
and U2326 (N_2326,In_891,In_849);
and U2327 (N_2327,In_294,In_419);
nand U2328 (N_2328,In_651,In_247);
nor U2329 (N_2329,In_793,In_628);
or U2330 (N_2330,In_674,In_110);
xnor U2331 (N_2331,In_662,In_236);
or U2332 (N_2332,In_447,In_491);
and U2333 (N_2333,In_10,In_437);
nor U2334 (N_2334,In_773,In_269);
or U2335 (N_2335,In_528,In_235);
or U2336 (N_2336,In_845,In_926);
xnor U2337 (N_2337,In_849,In_287);
and U2338 (N_2338,In_80,In_72);
nor U2339 (N_2339,In_493,In_245);
and U2340 (N_2340,In_853,In_894);
nand U2341 (N_2341,In_430,In_204);
or U2342 (N_2342,In_951,In_835);
nor U2343 (N_2343,In_460,In_800);
and U2344 (N_2344,In_574,In_385);
nor U2345 (N_2345,In_204,In_628);
or U2346 (N_2346,In_630,In_701);
and U2347 (N_2347,In_742,In_101);
nand U2348 (N_2348,In_800,In_385);
nand U2349 (N_2349,In_29,In_840);
nor U2350 (N_2350,In_258,In_9);
nor U2351 (N_2351,In_956,In_985);
nor U2352 (N_2352,In_330,In_139);
xor U2353 (N_2353,In_616,In_387);
nand U2354 (N_2354,In_349,In_406);
nand U2355 (N_2355,In_445,In_866);
nand U2356 (N_2356,In_186,In_749);
or U2357 (N_2357,In_221,In_597);
and U2358 (N_2358,In_979,In_103);
or U2359 (N_2359,In_288,In_911);
nand U2360 (N_2360,In_106,In_496);
nor U2361 (N_2361,In_403,In_186);
nor U2362 (N_2362,In_356,In_149);
and U2363 (N_2363,In_567,In_83);
nor U2364 (N_2364,In_795,In_695);
nand U2365 (N_2365,In_467,In_44);
and U2366 (N_2366,In_629,In_651);
and U2367 (N_2367,In_515,In_76);
nor U2368 (N_2368,In_469,In_390);
and U2369 (N_2369,In_930,In_290);
nand U2370 (N_2370,In_936,In_229);
or U2371 (N_2371,In_179,In_572);
nor U2372 (N_2372,In_625,In_448);
nand U2373 (N_2373,In_248,In_172);
and U2374 (N_2374,In_533,In_31);
nand U2375 (N_2375,In_41,In_590);
and U2376 (N_2376,In_215,In_201);
or U2377 (N_2377,In_220,In_467);
nor U2378 (N_2378,In_237,In_903);
or U2379 (N_2379,In_987,In_11);
nor U2380 (N_2380,In_564,In_135);
nor U2381 (N_2381,In_141,In_984);
nand U2382 (N_2382,In_372,In_693);
nor U2383 (N_2383,In_780,In_315);
nor U2384 (N_2384,In_718,In_796);
nor U2385 (N_2385,In_236,In_525);
nor U2386 (N_2386,In_312,In_480);
or U2387 (N_2387,In_342,In_6);
or U2388 (N_2388,In_530,In_648);
and U2389 (N_2389,In_152,In_564);
nand U2390 (N_2390,In_913,In_934);
and U2391 (N_2391,In_199,In_446);
xor U2392 (N_2392,In_481,In_447);
and U2393 (N_2393,In_625,In_33);
or U2394 (N_2394,In_926,In_956);
xnor U2395 (N_2395,In_347,In_975);
nand U2396 (N_2396,In_869,In_746);
or U2397 (N_2397,In_493,In_300);
and U2398 (N_2398,In_660,In_206);
and U2399 (N_2399,In_284,In_727);
nor U2400 (N_2400,In_321,In_118);
and U2401 (N_2401,In_325,In_860);
nand U2402 (N_2402,In_180,In_973);
and U2403 (N_2403,In_961,In_358);
nand U2404 (N_2404,In_585,In_926);
or U2405 (N_2405,In_785,In_19);
nand U2406 (N_2406,In_169,In_905);
nand U2407 (N_2407,In_138,In_534);
nor U2408 (N_2408,In_38,In_466);
nor U2409 (N_2409,In_355,In_543);
nand U2410 (N_2410,In_771,In_943);
nor U2411 (N_2411,In_825,In_165);
or U2412 (N_2412,In_962,In_939);
nor U2413 (N_2413,In_794,In_884);
and U2414 (N_2414,In_473,In_530);
nor U2415 (N_2415,In_446,In_664);
nand U2416 (N_2416,In_136,In_221);
or U2417 (N_2417,In_850,In_283);
and U2418 (N_2418,In_730,In_976);
nor U2419 (N_2419,In_181,In_434);
or U2420 (N_2420,In_393,In_118);
and U2421 (N_2421,In_588,In_700);
nand U2422 (N_2422,In_469,In_442);
nand U2423 (N_2423,In_818,In_134);
or U2424 (N_2424,In_746,In_847);
nand U2425 (N_2425,In_996,In_559);
nand U2426 (N_2426,In_836,In_343);
nor U2427 (N_2427,In_600,In_40);
nand U2428 (N_2428,In_604,In_867);
and U2429 (N_2429,In_228,In_599);
and U2430 (N_2430,In_6,In_687);
and U2431 (N_2431,In_729,In_78);
or U2432 (N_2432,In_927,In_574);
and U2433 (N_2433,In_651,In_126);
and U2434 (N_2434,In_726,In_347);
nand U2435 (N_2435,In_688,In_962);
nor U2436 (N_2436,In_445,In_724);
or U2437 (N_2437,In_414,In_373);
or U2438 (N_2438,In_745,In_876);
nor U2439 (N_2439,In_323,In_83);
nor U2440 (N_2440,In_1,In_828);
nor U2441 (N_2441,In_397,In_582);
or U2442 (N_2442,In_843,In_359);
and U2443 (N_2443,In_933,In_527);
nand U2444 (N_2444,In_748,In_691);
or U2445 (N_2445,In_609,In_581);
nor U2446 (N_2446,In_463,In_631);
or U2447 (N_2447,In_207,In_121);
nand U2448 (N_2448,In_802,In_744);
and U2449 (N_2449,In_629,In_194);
and U2450 (N_2450,In_844,In_641);
nor U2451 (N_2451,In_830,In_868);
or U2452 (N_2452,In_745,In_693);
xor U2453 (N_2453,In_517,In_466);
nand U2454 (N_2454,In_784,In_206);
and U2455 (N_2455,In_3,In_2);
nor U2456 (N_2456,In_115,In_357);
or U2457 (N_2457,In_147,In_909);
and U2458 (N_2458,In_667,In_487);
or U2459 (N_2459,In_8,In_882);
or U2460 (N_2460,In_293,In_774);
nand U2461 (N_2461,In_606,In_666);
nor U2462 (N_2462,In_821,In_305);
nor U2463 (N_2463,In_942,In_282);
or U2464 (N_2464,In_535,In_802);
or U2465 (N_2465,In_722,In_46);
and U2466 (N_2466,In_283,In_436);
or U2467 (N_2467,In_574,In_539);
and U2468 (N_2468,In_471,In_835);
and U2469 (N_2469,In_655,In_680);
or U2470 (N_2470,In_792,In_215);
nand U2471 (N_2471,In_425,In_340);
nor U2472 (N_2472,In_947,In_294);
nand U2473 (N_2473,In_239,In_933);
nor U2474 (N_2474,In_2,In_474);
nor U2475 (N_2475,In_112,In_659);
or U2476 (N_2476,In_697,In_454);
and U2477 (N_2477,In_110,In_524);
or U2478 (N_2478,In_650,In_189);
or U2479 (N_2479,In_35,In_856);
nor U2480 (N_2480,In_653,In_198);
or U2481 (N_2481,In_817,In_970);
nand U2482 (N_2482,In_606,In_84);
nand U2483 (N_2483,In_838,In_611);
or U2484 (N_2484,In_326,In_287);
or U2485 (N_2485,In_970,In_778);
nand U2486 (N_2486,In_606,In_86);
nor U2487 (N_2487,In_702,In_806);
and U2488 (N_2488,In_593,In_972);
nor U2489 (N_2489,In_591,In_897);
and U2490 (N_2490,In_425,In_720);
nand U2491 (N_2491,In_196,In_981);
nand U2492 (N_2492,In_431,In_533);
nor U2493 (N_2493,In_87,In_249);
or U2494 (N_2494,In_509,In_549);
and U2495 (N_2495,In_281,In_126);
or U2496 (N_2496,In_927,In_452);
or U2497 (N_2497,In_486,In_424);
and U2498 (N_2498,In_770,In_158);
and U2499 (N_2499,In_626,In_159);
nor U2500 (N_2500,In_64,In_842);
nor U2501 (N_2501,In_734,In_220);
nand U2502 (N_2502,In_431,In_605);
nor U2503 (N_2503,In_573,In_254);
nand U2504 (N_2504,In_805,In_688);
nor U2505 (N_2505,In_490,In_795);
nor U2506 (N_2506,In_420,In_3);
and U2507 (N_2507,In_547,In_348);
and U2508 (N_2508,In_950,In_704);
nand U2509 (N_2509,In_389,In_84);
nand U2510 (N_2510,In_287,In_910);
nor U2511 (N_2511,In_47,In_828);
nor U2512 (N_2512,In_312,In_65);
nor U2513 (N_2513,In_945,In_943);
nand U2514 (N_2514,In_995,In_714);
nor U2515 (N_2515,In_961,In_573);
or U2516 (N_2516,In_254,In_588);
nor U2517 (N_2517,In_726,In_176);
nand U2518 (N_2518,In_833,In_287);
nor U2519 (N_2519,In_520,In_457);
nand U2520 (N_2520,In_52,In_327);
xor U2521 (N_2521,In_926,In_539);
and U2522 (N_2522,In_300,In_989);
and U2523 (N_2523,In_95,In_249);
and U2524 (N_2524,In_764,In_178);
or U2525 (N_2525,In_499,In_148);
nand U2526 (N_2526,In_378,In_83);
or U2527 (N_2527,In_727,In_299);
and U2528 (N_2528,In_951,In_371);
and U2529 (N_2529,In_39,In_273);
or U2530 (N_2530,In_446,In_699);
or U2531 (N_2531,In_528,In_750);
and U2532 (N_2532,In_321,In_803);
and U2533 (N_2533,In_261,In_773);
and U2534 (N_2534,In_133,In_953);
nand U2535 (N_2535,In_873,In_717);
nand U2536 (N_2536,In_219,In_19);
nor U2537 (N_2537,In_197,In_37);
or U2538 (N_2538,In_25,In_432);
or U2539 (N_2539,In_529,In_395);
or U2540 (N_2540,In_171,In_702);
or U2541 (N_2541,In_23,In_356);
nand U2542 (N_2542,In_492,In_246);
nand U2543 (N_2543,In_110,In_580);
and U2544 (N_2544,In_248,In_85);
or U2545 (N_2545,In_721,In_346);
nor U2546 (N_2546,In_259,In_69);
and U2547 (N_2547,In_110,In_980);
or U2548 (N_2548,In_924,In_980);
and U2549 (N_2549,In_910,In_312);
and U2550 (N_2550,In_538,In_356);
nor U2551 (N_2551,In_508,In_524);
and U2552 (N_2552,In_667,In_739);
nor U2553 (N_2553,In_977,In_570);
nor U2554 (N_2554,In_123,In_633);
or U2555 (N_2555,In_114,In_43);
or U2556 (N_2556,In_933,In_553);
nand U2557 (N_2557,In_633,In_528);
or U2558 (N_2558,In_535,In_548);
or U2559 (N_2559,In_889,In_817);
nand U2560 (N_2560,In_239,In_957);
nor U2561 (N_2561,In_776,In_465);
nand U2562 (N_2562,In_111,In_826);
or U2563 (N_2563,In_274,In_507);
and U2564 (N_2564,In_757,In_509);
nor U2565 (N_2565,In_25,In_286);
or U2566 (N_2566,In_314,In_171);
or U2567 (N_2567,In_16,In_916);
nand U2568 (N_2568,In_169,In_871);
nor U2569 (N_2569,In_966,In_218);
or U2570 (N_2570,In_738,In_563);
or U2571 (N_2571,In_77,In_692);
or U2572 (N_2572,In_891,In_30);
and U2573 (N_2573,In_902,In_336);
or U2574 (N_2574,In_83,In_416);
and U2575 (N_2575,In_666,In_272);
nor U2576 (N_2576,In_778,In_514);
and U2577 (N_2577,In_228,In_278);
nor U2578 (N_2578,In_576,In_7);
nor U2579 (N_2579,In_772,In_830);
and U2580 (N_2580,In_45,In_148);
nand U2581 (N_2581,In_380,In_231);
and U2582 (N_2582,In_142,In_643);
and U2583 (N_2583,In_442,In_137);
and U2584 (N_2584,In_550,In_937);
nor U2585 (N_2585,In_211,In_918);
and U2586 (N_2586,In_122,In_443);
nand U2587 (N_2587,In_629,In_673);
nand U2588 (N_2588,In_120,In_938);
nor U2589 (N_2589,In_301,In_24);
nor U2590 (N_2590,In_655,In_912);
nor U2591 (N_2591,In_977,In_877);
nor U2592 (N_2592,In_221,In_365);
nor U2593 (N_2593,In_954,In_35);
xnor U2594 (N_2594,In_615,In_318);
nand U2595 (N_2595,In_928,In_200);
nand U2596 (N_2596,In_446,In_46);
and U2597 (N_2597,In_179,In_78);
and U2598 (N_2598,In_318,In_823);
and U2599 (N_2599,In_273,In_341);
nor U2600 (N_2600,In_81,In_352);
and U2601 (N_2601,In_709,In_589);
nand U2602 (N_2602,In_706,In_842);
or U2603 (N_2603,In_400,In_826);
xnor U2604 (N_2604,In_324,In_573);
or U2605 (N_2605,In_887,In_257);
and U2606 (N_2606,In_597,In_969);
nand U2607 (N_2607,In_486,In_477);
nand U2608 (N_2608,In_871,In_544);
xor U2609 (N_2609,In_662,In_610);
and U2610 (N_2610,In_135,In_736);
and U2611 (N_2611,In_65,In_960);
nor U2612 (N_2612,In_248,In_496);
and U2613 (N_2613,In_4,In_773);
nor U2614 (N_2614,In_863,In_63);
or U2615 (N_2615,In_694,In_640);
nand U2616 (N_2616,In_245,In_529);
nor U2617 (N_2617,In_846,In_790);
or U2618 (N_2618,In_23,In_828);
nor U2619 (N_2619,In_151,In_390);
and U2620 (N_2620,In_262,In_878);
nand U2621 (N_2621,In_117,In_752);
xor U2622 (N_2622,In_30,In_484);
nor U2623 (N_2623,In_677,In_670);
nor U2624 (N_2624,In_859,In_868);
or U2625 (N_2625,In_567,In_412);
and U2626 (N_2626,In_486,In_854);
and U2627 (N_2627,In_953,In_622);
or U2628 (N_2628,In_354,In_811);
nand U2629 (N_2629,In_924,In_358);
or U2630 (N_2630,In_235,In_961);
and U2631 (N_2631,In_217,In_579);
nand U2632 (N_2632,In_824,In_895);
or U2633 (N_2633,In_396,In_915);
nand U2634 (N_2634,In_316,In_139);
nand U2635 (N_2635,In_102,In_321);
or U2636 (N_2636,In_227,In_738);
and U2637 (N_2637,In_372,In_578);
nand U2638 (N_2638,In_743,In_495);
or U2639 (N_2639,In_465,In_724);
nor U2640 (N_2640,In_923,In_710);
nand U2641 (N_2641,In_690,In_544);
and U2642 (N_2642,In_217,In_820);
nor U2643 (N_2643,In_901,In_443);
or U2644 (N_2644,In_300,In_182);
nor U2645 (N_2645,In_297,In_751);
and U2646 (N_2646,In_726,In_301);
and U2647 (N_2647,In_342,In_407);
or U2648 (N_2648,In_365,In_887);
nand U2649 (N_2649,In_727,In_329);
nand U2650 (N_2650,In_117,In_408);
or U2651 (N_2651,In_951,In_68);
and U2652 (N_2652,In_281,In_957);
nand U2653 (N_2653,In_577,In_19);
and U2654 (N_2654,In_88,In_880);
nor U2655 (N_2655,In_641,In_792);
xnor U2656 (N_2656,In_515,In_997);
nand U2657 (N_2657,In_454,In_945);
nor U2658 (N_2658,In_9,In_269);
and U2659 (N_2659,In_310,In_435);
and U2660 (N_2660,In_283,In_930);
nor U2661 (N_2661,In_14,In_857);
nand U2662 (N_2662,In_757,In_638);
and U2663 (N_2663,In_315,In_847);
xnor U2664 (N_2664,In_950,In_239);
nand U2665 (N_2665,In_906,In_640);
and U2666 (N_2666,In_978,In_35);
or U2667 (N_2667,In_978,In_597);
and U2668 (N_2668,In_86,In_917);
and U2669 (N_2669,In_730,In_91);
xor U2670 (N_2670,In_158,In_223);
and U2671 (N_2671,In_843,In_495);
or U2672 (N_2672,In_334,In_461);
and U2673 (N_2673,In_718,In_78);
and U2674 (N_2674,In_747,In_688);
nor U2675 (N_2675,In_237,In_68);
and U2676 (N_2676,In_250,In_286);
nor U2677 (N_2677,In_194,In_282);
nor U2678 (N_2678,In_428,In_415);
nor U2679 (N_2679,In_38,In_409);
and U2680 (N_2680,In_19,In_830);
nor U2681 (N_2681,In_857,In_897);
and U2682 (N_2682,In_673,In_572);
and U2683 (N_2683,In_976,In_766);
and U2684 (N_2684,In_673,In_323);
nor U2685 (N_2685,In_922,In_945);
nor U2686 (N_2686,In_266,In_790);
and U2687 (N_2687,In_228,In_951);
nand U2688 (N_2688,In_319,In_569);
nand U2689 (N_2689,In_916,In_624);
or U2690 (N_2690,In_805,In_934);
and U2691 (N_2691,In_367,In_844);
nand U2692 (N_2692,In_799,In_268);
or U2693 (N_2693,In_509,In_983);
nor U2694 (N_2694,In_869,In_580);
nor U2695 (N_2695,In_282,In_606);
nand U2696 (N_2696,In_675,In_120);
nor U2697 (N_2697,In_495,In_34);
or U2698 (N_2698,In_71,In_217);
nand U2699 (N_2699,In_141,In_462);
nor U2700 (N_2700,In_956,In_635);
nand U2701 (N_2701,In_710,In_936);
nand U2702 (N_2702,In_204,In_900);
xor U2703 (N_2703,In_339,In_877);
nor U2704 (N_2704,In_284,In_203);
nor U2705 (N_2705,In_482,In_390);
or U2706 (N_2706,In_822,In_912);
nor U2707 (N_2707,In_134,In_218);
nor U2708 (N_2708,In_567,In_610);
or U2709 (N_2709,In_609,In_924);
and U2710 (N_2710,In_337,In_820);
and U2711 (N_2711,In_114,In_653);
nor U2712 (N_2712,In_540,In_58);
nor U2713 (N_2713,In_365,In_691);
and U2714 (N_2714,In_949,In_126);
or U2715 (N_2715,In_455,In_506);
and U2716 (N_2716,In_642,In_887);
nand U2717 (N_2717,In_703,In_104);
and U2718 (N_2718,In_403,In_613);
and U2719 (N_2719,In_559,In_65);
nand U2720 (N_2720,In_853,In_619);
nor U2721 (N_2721,In_43,In_554);
nor U2722 (N_2722,In_393,In_763);
nand U2723 (N_2723,In_721,In_13);
nor U2724 (N_2724,In_944,In_628);
nor U2725 (N_2725,In_199,In_597);
nand U2726 (N_2726,In_263,In_841);
nor U2727 (N_2727,In_812,In_189);
nor U2728 (N_2728,In_712,In_532);
or U2729 (N_2729,In_710,In_625);
and U2730 (N_2730,In_669,In_389);
nor U2731 (N_2731,In_910,In_224);
nor U2732 (N_2732,In_406,In_515);
or U2733 (N_2733,In_341,In_390);
nor U2734 (N_2734,In_638,In_261);
and U2735 (N_2735,In_572,In_23);
xor U2736 (N_2736,In_509,In_770);
or U2737 (N_2737,In_193,In_351);
or U2738 (N_2738,In_670,In_869);
nand U2739 (N_2739,In_141,In_814);
nand U2740 (N_2740,In_9,In_251);
and U2741 (N_2741,In_111,In_782);
nor U2742 (N_2742,In_564,In_110);
nor U2743 (N_2743,In_196,In_472);
nand U2744 (N_2744,In_998,In_581);
and U2745 (N_2745,In_703,In_208);
nand U2746 (N_2746,In_558,In_546);
nand U2747 (N_2747,In_744,In_619);
nor U2748 (N_2748,In_755,In_237);
or U2749 (N_2749,In_741,In_471);
and U2750 (N_2750,In_632,In_853);
or U2751 (N_2751,In_439,In_810);
nor U2752 (N_2752,In_1,In_265);
nand U2753 (N_2753,In_383,In_938);
nor U2754 (N_2754,In_893,In_472);
and U2755 (N_2755,In_784,In_871);
and U2756 (N_2756,In_552,In_941);
nand U2757 (N_2757,In_933,In_120);
and U2758 (N_2758,In_431,In_545);
and U2759 (N_2759,In_231,In_305);
and U2760 (N_2760,In_499,In_630);
and U2761 (N_2761,In_557,In_219);
or U2762 (N_2762,In_820,In_886);
and U2763 (N_2763,In_656,In_858);
nor U2764 (N_2764,In_684,In_991);
nor U2765 (N_2765,In_10,In_24);
nor U2766 (N_2766,In_586,In_841);
xor U2767 (N_2767,In_129,In_31);
or U2768 (N_2768,In_748,In_255);
nor U2769 (N_2769,In_264,In_468);
nand U2770 (N_2770,In_972,In_279);
or U2771 (N_2771,In_858,In_42);
and U2772 (N_2772,In_158,In_603);
nand U2773 (N_2773,In_724,In_475);
and U2774 (N_2774,In_438,In_848);
nor U2775 (N_2775,In_306,In_543);
and U2776 (N_2776,In_186,In_25);
or U2777 (N_2777,In_713,In_340);
nor U2778 (N_2778,In_15,In_764);
nor U2779 (N_2779,In_412,In_639);
and U2780 (N_2780,In_92,In_694);
nand U2781 (N_2781,In_24,In_813);
and U2782 (N_2782,In_591,In_620);
or U2783 (N_2783,In_873,In_782);
and U2784 (N_2784,In_423,In_966);
nor U2785 (N_2785,In_777,In_222);
and U2786 (N_2786,In_856,In_911);
or U2787 (N_2787,In_404,In_206);
nand U2788 (N_2788,In_173,In_473);
nor U2789 (N_2789,In_677,In_885);
and U2790 (N_2790,In_660,In_66);
nand U2791 (N_2791,In_342,In_27);
nor U2792 (N_2792,In_841,In_229);
nor U2793 (N_2793,In_207,In_195);
nand U2794 (N_2794,In_48,In_776);
nand U2795 (N_2795,In_893,In_176);
or U2796 (N_2796,In_61,In_358);
and U2797 (N_2797,In_435,In_617);
nor U2798 (N_2798,In_988,In_936);
and U2799 (N_2799,In_176,In_488);
and U2800 (N_2800,In_241,In_694);
and U2801 (N_2801,In_483,In_651);
nor U2802 (N_2802,In_973,In_602);
nand U2803 (N_2803,In_939,In_680);
nor U2804 (N_2804,In_511,In_23);
and U2805 (N_2805,In_993,In_345);
nand U2806 (N_2806,In_560,In_192);
xnor U2807 (N_2807,In_817,In_349);
and U2808 (N_2808,In_439,In_471);
nand U2809 (N_2809,In_174,In_697);
or U2810 (N_2810,In_904,In_335);
nand U2811 (N_2811,In_925,In_813);
nand U2812 (N_2812,In_123,In_55);
nor U2813 (N_2813,In_207,In_392);
nor U2814 (N_2814,In_602,In_3);
or U2815 (N_2815,In_380,In_296);
and U2816 (N_2816,In_586,In_525);
nor U2817 (N_2817,In_543,In_60);
nor U2818 (N_2818,In_49,In_956);
nand U2819 (N_2819,In_945,In_103);
nand U2820 (N_2820,In_197,In_881);
or U2821 (N_2821,In_571,In_344);
nand U2822 (N_2822,In_559,In_528);
nor U2823 (N_2823,In_409,In_691);
and U2824 (N_2824,In_769,In_738);
or U2825 (N_2825,In_417,In_838);
or U2826 (N_2826,In_719,In_202);
nand U2827 (N_2827,In_821,In_496);
and U2828 (N_2828,In_613,In_275);
or U2829 (N_2829,In_167,In_729);
nand U2830 (N_2830,In_607,In_820);
nor U2831 (N_2831,In_447,In_398);
nor U2832 (N_2832,In_173,In_513);
and U2833 (N_2833,In_465,In_932);
nor U2834 (N_2834,In_879,In_698);
or U2835 (N_2835,In_629,In_721);
nor U2836 (N_2836,In_204,In_634);
xor U2837 (N_2837,In_528,In_173);
and U2838 (N_2838,In_31,In_587);
nor U2839 (N_2839,In_76,In_394);
and U2840 (N_2840,In_268,In_269);
nor U2841 (N_2841,In_552,In_499);
or U2842 (N_2842,In_92,In_599);
nand U2843 (N_2843,In_508,In_989);
nand U2844 (N_2844,In_466,In_33);
nand U2845 (N_2845,In_939,In_433);
and U2846 (N_2846,In_543,In_80);
nand U2847 (N_2847,In_341,In_18);
and U2848 (N_2848,In_961,In_872);
nor U2849 (N_2849,In_228,In_846);
and U2850 (N_2850,In_63,In_660);
and U2851 (N_2851,In_601,In_837);
and U2852 (N_2852,In_610,In_445);
nor U2853 (N_2853,In_62,In_566);
nand U2854 (N_2854,In_221,In_127);
xnor U2855 (N_2855,In_266,In_340);
nor U2856 (N_2856,In_947,In_328);
or U2857 (N_2857,In_620,In_459);
or U2858 (N_2858,In_28,In_92);
or U2859 (N_2859,In_391,In_265);
or U2860 (N_2860,In_950,In_624);
or U2861 (N_2861,In_454,In_219);
or U2862 (N_2862,In_570,In_119);
nor U2863 (N_2863,In_550,In_586);
nand U2864 (N_2864,In_678,In_967);
and U2865 (N_2865,In_447,In_341);
nor U2866 (N_2866,In_910,In_534);
nor U2867 (N_2867,In_388,In_572);
nand U2868 (N_2868,In_647,In_59);
or U2869 (N_2869,In_859,In_624);
nor U2870 (N_2870,In_298,In_879);
nand U2871 (N_2871,In_258,In_26);
or U2872 (N_2872,In_368,In_813);
or U2873 (N_2873,In_156,In_876);
nand U2874 (N_2874,In_740,In_344);
or U2875 (N_2875,In_118,In_993);
xor U2876 (N_2876,In_316,In_981);
nor U2877 (N_2877,In_914,In_526);
xnor U2878 (N_2878,In_376,In_478);
nand U2879 (N_2879,In_222,In_90);
nand U2880 (N_2880,In_843,In_356);
and U2881 (N_2881,In_60,In_935);
or U2882 (N_2882,In_483,In_535);
nor U2883 (N_2883,In_545,In_475);
nor U2884 (N_2884,In_229,In_63);
or U2885 (N_2885,In_679,In_803);
and U2886 (N_2886,In_481,In_760);
nand U2887 (N_2887,In_132,In_771);
nand U2888 (N_2888,In_720,In_418);
nor U2889 (N_2889,In_107,In_498);
or U2890 (N_2890,In_442,In_213);
nand U2891 (N_2891,In_644,In_864);
or U2892 (N_2892,In_412,In_287);
or U2893 (N_2893,In_969,In_530);
nor U2894 (N_2894,In_814,In_650);
nand U2895 (N_2895,In_608,In_713);
or U2896 (N_2896,In_452,In_2);
nand U2897 (N_2897,In_481,In_299);
or U2898 (N_2898,In_581,In_970);
or U2899 (N_2899,In_353,In_842);
nand U2900 (N_2900,In_407,In_768);
xor U2901 (N_2901,In_459,In_88);
or U2902 (N_2902,In_422,In_55);
nand U2903 (N_2903,In_720,In_479);
nor U2904 (N_2904,In_828,In_292);
or U2905 (N_2905,In_139,In_296);
nor U2906 (N_2906,In_789,In_330);
and U2907 (N_2907,In_485,In_83);
nand U2908 (N_2908,In_556,In_339);
or U2909 (N_2909,In_566,In_485);
nor U2910 (N_2910,In_259,In_468);
nand U2911 (N_2911,In_993,In_394);
and U2912 (N_2912,In_963,In_857);
nand U2913 (N_2913,In_67,In_169);
or U2914 (N_2914,In_376,In_278);
nand U2915 (N_2915,In_430,In_779);
or U2916 (N_2916,In_25,In_255);
or U2917 (N_2917,In_181,In_397);
nor U2918 (N_2918,In_297,In_705);
or U2919 (N_2919,In_641,In_788);
nand U2920 (N_2920,In_845,In_879);
nand U2921 (N_2921,In_540,In_939);
xnor U2922 (N_2922,In_616,In_676);
nor U2923 (N_2923,In_17,In_852);
or U2924 (N_2924,In_681,In_978);
nor U2925 (N_2925,In_852,In_390);
nand U2926 (N_2926,In_690,In_27);
nand U2927 (N_2927,In_436,In_373);
or U2928 (N_2928,In_325,In_875);
or U2929 (N_2929,In_731,In_333);
nor U2930 (N_2930,In_950,In_898);
and U2931 (N_2931,In_573,In_874);
and U2932 (N_2932,In_616,In_0);
nor U2933 (N_2933,In_48,In_423);
nand U2934 (N_2934,In_474,In_410);
and U2935 (N_2935,In_559,In_816);
or U2936 (N_2936,In_148,In_235);
or U2937 (N_2937,In_606,In_662);
nor U2938 (N_2938,In_358,In_842);
or U2939 (N_2939,In_961,In_610);
nand U2940 (N_2940,In_827,In_89);
or U2941 (N_2941,In_279,In_807);
nand U2942 (N_2942,In_867,In_855);
and U2943 (N_2943,In_728,In_21);
and U2944 (N_2944,In_214,In_198);
or U2945 (N_2945,In_117,In_165);
xnor U2946 (N_2946,In_747,In_119);
and U2947 (N_2947,In_148,In_981);
nand U2948 (N_2948,In_369,In_984);
or U2949 (N_2949,In_5,In_609);
nor U2950 (N_2950,In_524,In_99);
nand U2951 (N_2951,In_699,In_741);
nor U2952 (N_2952,In_177,In_713);
nand U2953 (N_2953,In_811,In_749);
nand U2954 (N_2954,In_19,In_27);
nand U2955 (N_2955,In_850,In_45);
or U2956 (N_2956,In_168,In_256);
and U2957 (N_2957,In_384,In_435);
nor U2958 (N_2958,In_406,In_463);
or U2959 (N_2959,In_820,In_367);
nor U2960 (N_2960,In_317,In_307);
or U2961 (N_2961,In_331,In_605);
nand U2962 (N_2962,In_695,In_599);
nand U2963 (N_2963,In_671,In_835);
and U2964 (N_2964,In_621,In_340);
xor U2965 (N_2965,In_423,In_962);
nor U2966 (N_2966,In_805,In_910);
or U2967 (N_2967,In_874,In_288);
nor U2968 (N_2968,In_912,In_921);
nor U2969 (N_2969,In_989,In_457);
and U2970 (N_2970,In_188,In_665);
nor U2971 (N_2971,In_833,In_163);
and U2972 (N_2972,In_285,In_45);
or U2973 (N_2973,In_302,In_603);
nand U2974 (N_2974,In_646,In_7);
or U2975 (N_2975,In_163,In_293);
nand U2976 (N_2976,In_276,In_206);
nand U2977 (N_2977,In_79,In_328);
nor U2978 (N_2978,In_588,In_575);
nor U2979 (N_2979,In_656,In_160);
nand U2980 (N_2980,In_667,In_423);
or U2981 (N_2981,In_189,In_638);
and U2982 (N_2982,In_498,In_635);
and U2983 (N_2983,In_28,In_731);
or U2984 (N_2984,In_398,In_386);
nor U2985 (N_2985,In_124,In_696);
nor U2986 (N_2986,In_692,In_78);
nor U2987 (N_2987,In_512,In_573);
or U2988 (N_2988,In_869,In_262);
or U2989 (N_2989,In_797,In_569);
and U2990 (N_2990,In_170,In_484);
nand U2991 (N_2991,In_400,In_442);
nand U2992 (N_2992,In_770,In_759);
and U2993 (N_2993,In_955,In_645);
and U2994 (N_2994,In_686,In_139);
nand U2995 (N_2995,In_889,In_222);
and U2996 (N_2996,In_223,In_162);
nand U2997 (N_2997,In_763,In_562);
nor U2998 (N_2998,In_891,In_787);
and U2999 (N_2999,In_589,In_507);
nand U3000 (N_3000,In_255,In_162);
or U3001 (N_3001,In_336,In_600);
and U3002 (N_3002,In_55,In_593);
nor U3003 (N_3003,In_777,In_588);
nand U3004 (N_3004,In_210,In_957);
nand U3005 (N_3005,In_264,In_753);
and U3006 (N_3006,In_234,In_405);
nor U3007 (N_3007,In_135,In_537);
nand U3008 (N_3008,In_112,In_107);
nand U3009 (N_3009,In_298,In_386);
xnor U3010 (N_3010,In_688,In_979);
or U3011 (N_3011,In_515,In_99);
xor U3012 (N_3012,In_397,In_696);
nor U3013 (N_3013,In_383,In_581);
and U3014 (N_3014,In_238,In_833);
and U3015 (N_3015,In_541,In_533);
and U3016 (N_3016,In_76,In_270);
nand U3017 (N_3017,In_20,In_568);
nor U3018 (N_3018,In_730,In_784);
or U3019 (N_3019,In_755,In_904);
nor U3020 (N_3020,In_351,In_353);
nand U3021 (N_3021,In_834,In_688);
nand U3022 (N_3022,In_971,In_375);
nor U3023 (N_3023,In_907,In_59);
and U3024 (N_3024,In_148,In_262);
nor U3025 (N_3025,In_370,In_82);
and U3026 (N_3026,In_852,In_512);
nor U3027 (N_3027,In_140,In_757);
and U3028 (N_3028,In_923,In_902);
xor U3029 (N_3029,In_615,In_773);
or U3030 (N_3030,In_196,In_674);
nand U3031 (N_3031,In_793,In_888);
nor U3032 (N_3032,In_666,In_167);
and U3033 (N_3033,In_153,In_711);
nor U3034 (N_3034,In_77,In_105);
nor U3035 (N_3035,In_951,In_264);
or U3036 (N_3036,In_587,In_268);
nand U3037 (N_3037,In_539,In_963);
or U3038 (N_3038,In_843,In_653);
nand U3039 (N_3039,In_192,In_829);
and U3040 (N_3040,In_57,In_114);
or U3041 (N_3041,In_520,In_63);
nand U3042 (N_3042,In_96,In_921);
nor U3043 (N_3043,In_770,In_455);
nand U3044 (N_3044,In_241,In_274);
nor U3045 (N_3045,In_634,In_294);
nand U3046 (N_3046,In_394,In_141);
nor U3047 (N_3047,In_487,In_773);
nor U3048 (N_3048,In_721,In_995);
nor U3049 (N_3049,In_262,In_223);
and U3050 (N_3050,In_827,In_679);
and U3051 (N_3051,In_661,In_149);
and U3052 (N_3052,In_807,In_970);
or U3053 (N_3053,In_256,In_232);
and U3054 (N_3054,In_133,In_553);
or U3055 (N_3055,In_673,In_671);
or U3056 (N_3056,In_716,In_344);
or U3057 (N_3057,In_277,In_911);
or U3058 (N_3058,In_246,In_610);
nand U3059 (N_3059,In_644,In_649);
or U3060 (N_3060,In_843,In_850);
or U3061 (N_3061,In_108,In_284);
or U3062 (N_3062,In_514,In_978);
nor U3063 (N_3063,In_414,In_150);
nor U3064 (N_3064,In_424,In_855);
nor U3065 (N_3065,In_364,In_650);
nand U3066 (N_3066,In_263,In_189);
and U3067 (N_3067,In_825,In_378);
or U3068 (N_3068,In_606,In_44);
nand U3069 (N_3069,In_676,In_141);
xor U3070 (N_3070,In_15,In_392);
nand U3071 (N_3071,In_499,In_53);
or U3072 (N_3072,In_637,In_946);
and U3073 (N_3073,In_744,In_113);
nand U3074 (N_3074,In_775,In_280);
nor U3075 (N_3075,In_245,In_479);
nand U3076 (N_3076,In_852,In_166);
or U3077 (N_3077,In_142,In_734);
or U3078 (N_3078,In_718,In_345);
nand U3079 (N_3079,In_31,In_164);
or U3080 (N_3080,In_784,In_631);
nand U3081 (N_3081,In_174,In_507);
or U3082 (N_3082,In_241,In_72);
nand U3083 (N_3083,In_233,In_761);
nor U3084 (N_3084,In_398,In_393);
and U3085 (N_3085,In_977,In_803);
nor U3086 (N_3086,In_874,In_133);
and U3087 (N_3087,In_745,In_139);
xnor U3088 (N_3088,In_154,In_549);
and U3089 (N_3089,In_886,In_701);
and U3090 (N_3090,In_925,In_131);
or U3091 (N_3091,In_611,In_687);
nand U3092 (N_3092,In_323,In_928);
nor U3093 (N_3093,In_361,In_814);
and U3094 (N_3094,In_856,In_896);
nor U3095 (N_3095,In_923,In_300);
nand U3096 (N_3096,In_481,In_550);
or U3097 (N_3097,In_694,In_716);
nand U3098 (N_3098,In_28,In_88);
nand U3099 (N_3099,In_864,In_7);
and U3100 (N_3100,In_196,In_374);
or U3101 (N_3101,In_894,In_454);
nand U3102 (N_3102,In_402,In_217);
nor U3103 (N_3103,In_87,In_330);
and U3104 (N_3104,In_743,In_98);
nor U3105 (N_3105,In_59,In_414);
or U3106 (N_3106,In_279,In_997);
nor U3107 (N_3107,In_321,In_674);
nand U3108 (N_3108,In_959,In_352);
nand U3109 (N_3109,In_401,In_662);
nor U3110 (N_3110,In_564,In_372);
or U3111 (N_3111,In_108,In_696);
nand U3112 (N_3112,In_220,In_438);
or U3113 (N_3113,In_207,In_241);
nand U3114 (N_3114,In_357,In_996);
nor U3115 (N_3115,In_628,In_706);
nand U3116 (N_3116,In_109,In_782);
and U3117 (N_3117,In_345,In_82);
nor U3118 (N_3118,In_724,In_623);
or U3119 (N_3119,In_508,In_747);
and U3120 (N_3120,In_15,In_159);
or U3121 (N_3121,In_977,In_2);
nand U3122 (N_3122,In_970,In_805);
and U3123 (N_3123,In_871,In_681);
or U3124 (N_3124,In_633,In_257);
and U3125 (N_3125,In_347,In_808);
nor U3126 (N_3126,In_546,In_672);
or U3127 (N_3127,In_123,In_230);
or U3128 (N_3128,In_233,In_394);
and U3129 (N_3129,In_619,In_919);
nand U3130 (N_3130,In_964,In_590);
nand U3131 (N_3131,In_822,In_403);
or U3132 (N_3132,In_409,In_78);
and U3133 (N_3133,In_110,In_468);
or U3134 (N_3134,In_336,In_901);
or U3135 (N_3135,In_973,In_192);
and U3136 (N_3136,In_930,In_961);
nand U3137 (N_3137,In_302,In_98);
nor U3138 (N_3138,In_774,In_590);
nor U3139 (N_3139,In_815,In_620);
or U3140 (N_3140,In_949,In_792);
and U3141 (N_3141,In_886,In_786);
and U3142 (N_3142,In_119,In_796);
or U3143 (N_3143,In_511,In_515);
nand U3144 (N_3144,In_829,In_377);
nand U3145 (N_3145,In_434,In_245);
nor U3146 (N_3146,In_423,In_402);
nor U3147 (N_3147,In_68,In_459);
nand U3148 (N_3148,In_234,In_773);
nor U3149 (N_3149,In_47,In_792);
or U3150 (N_3150,In_759,In_471);
and U3151 (N_3151,In_935,In_547);
nand U3152 (N_3152,In_634,In_233);
xnor U3153 (N_3153,In_395,In_115);
and U3154 (N_3154,In_396,In_743);
nand U3155 (N_3155,In_810,In_139);
nor U3156 (N_3156,In_442,In_942);
and U3157 (N_3157,In_665,In_452);
or U3158 (N_3158,In_837,In_493);
nor U3159 (N_3159,In_432,In_147);
nor U3160 (N_3160,In_439,In_486);
nand U3161 (N_3161,In_447,In_925);
and U3162 (N_3162,In_203,In_272);
or U3163 (N_3163,In_232,In_218);
or U3164 (N_3164,In_297,In_955);
nand U3165 (N_3165,In_854,In_708);
nor U3166 (N_3166,In_558,In_482);
or U3167 (N_3167,In_170,In_765);
or U3168 (N_3168,In_290,In_851);
or U3169 (N_3169,In_639,In_325);
nand U3170 (N_3170,In_97,In_767);
nor U3171 (N_3171,In_101,In_122);
nand U3172 (N_3172,In_158,In_1);
and U3173 (N_3173,In_294,In_19);
nand U3174 (N_3174,In_832,In_351);
or U3175 (N_3175,In_837,In_233);
and U3176 (N_3176,In_827,In_834);
and U3177 (N_3177,In_856,In_422);
and U3178 (N_3178,In_997,In_547);
nand U3179 (N_3179,In_615,In_529);
xor U3180 (N_3180,In_117,In_389);
or U3181 (N_3181,In_740,In_554);
or U3182 (N_3182,In_578,In_3);
nand U3183 (N_3183,In_2,In_63);
and U3184 (N_3184,In_836,In_597);
or U3185 (N_3185,In_797,In_767);
nand U3186 (N_3186,In_481,In_577);
and U3187 (N_3187,In_296,In_71);
and U3188 (N_3188,In_830,In_425);
and U3189 (N_3189,In_377,In_619);
and U3190 (N_3190,In_283,In_544);
nand U3191 (N_3191,In_422,In_338);
nor U3192 (N_3192,In_807,In_393);
nor U3193 (N_3193,In_575,In_737);
nor U3194 (N_3194,In_785,In_638);
nor U3195 (N_3195,In_352,In_185);
nor U3196 (N_3196,In_681,In_266);
or U3197 (N_3197,In_582,In_481);
nor U3198 (N_3198,In_68,In_1);
or U3199 (N_3199,In_754,In_121);
or U3200 (N_3200,In_595,In_434);
or U3201 (N_3201,In_470,In_315);
nor U3202 (N_3202,In_751,In_528);
and U3203 (N_3203,In_189,In_545);
nor U3204 (N_3204,In_932,In_694);
nand U3205 (N_3205,In_573,In_334);
nand U3206 (N_3206,In_474,In_616);
nand U3207 (N_3207,In_263,In_449);
and U3208 (N_3208,In_626,In_9);
nand U3209 (N_3209,In_677,In_359);
and U3210 (N_3210,In_419,In_256);
and U3211 (N_3211,In_863,In_506);
nor U3212 (N_3212,In_171,In_388);
xor U3213 (N_3213,In_595,In_709);
nor U3214 (N_3214,In_882,In_869);
nand U3215 (N_3215,In_436,In_433);
nor U3216 (N_3216,In_399,In_143);
nand U3217 (N_3217,In_715,In_65);
nand U3218 (N_3218,In_574,In_389);
and U3219 (N_3219,In_108,In_263);
and U3220 (N_3220,In_326,In_399);
nand U3221 (N_3221,In_377,In_501);
and U3222 (N_3222,In_761,In_657);
nor U3223 (N_3223,In_125,In_946);
or U3224 (N_3224,In_628,In_338);
and U3225 (N_3225,In_803,In_31);
xnor U3226 (N_3226,In_613,In_827);
or U3227 (N_3227,In_363,In_617);
nand U3228 (N_3228,In_409,In_125);
nand U3229 (N_3229,In_32,In_633);
and U3230 (N_3230,In_368,In_401);
or U3231 (N_3231,In_146,In_330);
nand U3232 (N_3232,In_36,In_680);
nand U3233 (N_3233,In_598,In_489);
nor U3234 (N_3234,In_786,In_74);
and U3235 (N_3235,In_215,In_193);
nor U3236 (N_3236,In_102,In_32);
nand U3237 (N_3237,In_383,In_486);
nand U3238 (N_3238,In_912,In_606);
or U3239 (N_3239,In_244,In_589);
nand U3240 (N_3240,In_970,In_526);
nor U3241 (N_3241,In_662,In_238);
nand U3242 (N_3242,In_606,In_408);
nand U3243 (N_3243,In_154,In_205);
or U3244 (N_3244,In_407,In_458);
nor U3245 (N_3245,In_611,In_61);
and U3246 (N_3246,In_178,In_955);
and U3247 (N_3247,In_471,In_425);
nor U3248 (N_3248,In_269,In_578);
or U3249 (N_3249,In_521,In_205);
or U3250 (N_3250,In_704,In_233);
and U3251 (N_3251,In_10,In_983);
nor U3252 (N_3252,In_733,In_520);
xnor U3253 (N_3253,In_424,In_727);
nor U3254 (N_3254,In_112,In_487);
and U3255 (N_3255,In_710,In_811);
and U3256 (N_3256,In_374,In_965);
nand U3257 (N_3257,In_749,In_228);
nor U3258 (N_3258,In_142,In_890);
and U3259 (N_3259,In_137,In_633);
or U3260 (N_3260,In_480,In_657);
nor U3261 (N_3261,In_184,In_897);
nand U3262 (N_3262,In_190,In_173);
nand U3263 (N_3263,In_587,In_925);
and U3264 (N_3264,In_44,In_20);
nand U3265 (N_3265,In_172,In_467);
and U3266 (N_3266,In_723,In_637);
or U3267 (N_3267,In_733,In_947);
and U3268 (N_3268,In_886,In_975);
or U3269 (N_3269,In_759,In_698);
nand U3270 (N_3270,In_187,In_23);
nor U3271 (N_3271,In_148,In_656);
or U3272 (N_3272,In_258,In_676);
or U3273 (N_3273,In_48,In_722);
nand U3274 (N_3274,In_504,In_683);
or U3275 (N_3275,In_484,In_595);
or U3276 (N_3276,In_212,In_41);
xor U3277 (N_3277,In_693,In_619);
nor U3278 (N_3278,In_1,In_259);
nor U3279 (N_3279,In_315,In_12);
nor U3280 (N_3280,In_383,In_592);
nor U3281 (N_3281,In_233,In_944);
or U3282 (N_3282,In_380,In_703);
and U3283 (N_3283,In_821,In_830);
and U3284 (N_3284,In_974,In_356);
nand U3285 (N_3285,In_816,In_467);
nand U3286 (N_3286,In_528,In_770);
or U3287 (N_3287,In_701,In_524);
nand U3288 (N_3288,In_946,In_275);
nor U3289 (N_3289,In_265,In_55);
and U3290 (N_3290,In_904,In_337);
or U3291 (N_3291,In_737,In_891);
and U3292 (N_3292,In_736,In_375);
or U3293 (N_3293,In_648,In_823);
and U3294 (N_3294,In_379,In_347);
or U3295 (N_3295,In_139,In_841);
and U3296 (N_3296,In_527,In_493);
or U3297 (N_3297,In_382,In_408);
and U3298 (N_3298,In_351,In_894);
nor U3299 (N_3299,In_349,In_986);
nor U3300 (N_3300,In_811,In_40);
and U3301 (N_3301,In_619,In_251);
or U3302 (N_3302,In_501,In_601);
and U3303 (N_3303,In_449,In_334);
nand U3304 (N_3304,In_341,In_454);
nand U3305 (N_3305,In_65,In_95);
or U3306 (N_3306,In_742,In_619);
nand U3307 (N_3307,In_890,In_335);
nand U3308 (N_3308,In_509,In_676);
and U3309 (N_3309,In_721,In_806);
and U3310 (N_3310,In_609,In_416);
nor U3311 (N_3311,In_631,In_734);
and U3312 (N_3312,In_113,In_802);
and U3313 (N_3313,In_952,In_964);
or U3314 (N_3314,In_6,In_908);
nand U3315 (N_3315,In_875,In_947);
nand U3316 (N_3316,In_298,In_630);
nor U3317 (N_3317,In_756,In_417);
and U3318 (N_3318,In_146,In_138);
or U3319 (N_3319,In_988,In_836);
and U3320 (N_3320,In_819,In_963);
and U3321 (N_3321,In_794,In_247);
or U3322 (N_3322,In_655,In_592);
nand U3323 (N_3323,In_234,In_46);
and U3324 (N_3324,In_320,In_584);
nor U3325 (N_3325,In_72,In_548);
nand U3326 (N_3326,In_311,In_442);
nor U3327 (N_3327,In_584,In_386);
and U3328 (N_3328,In_818,In_28);
nand U3329 (N_3329,In_539,In_69);
nor U3330 (N_3330,In_364,In_186);
and U3331 (N_3331,In_545,In_925);
and U3332 (N_3332,In_162,In_631);
and U3333 (N_3333,In_567,In_738);
nor U3334 (N_3334,In_748,In_835);
and U3335 (N_3335,In_632,In_413);
nand U3336 (N_3336,In_914,In_350);
or U3337 (N_3337,In_448,In_269);
nor U3338 (N_3338,In_380,In_92);
nand U3339 (N_3339,In_99,In_636);
xor U3340 (N_3340,In_399,In_520);
or U3341 (N_3341,In_351,In_228);
nor U3342 (N_3342,In_988,In_941);
or U3343 (N_3343,In_367,In_4);
and U3344 (N_3344,In_360,In_570);
or U3345 (N_3345,In_399,In_588);
nor U3346 (N_3346,In_94,In_940);
nand U3347 (N_3347,In_856,In_348);
nand U3348 (N_3348,In_482,In_20);
nand U3349 (N_3349,In_416,In_620);
and U3350 (N_3350,In_972,In_553);
and U3351 (N_3351,In_505,In_185);
nand U3352 (N_3352,In_809,In_75);
nor U3353 (N_3353,In_766,In_350);
nand U3354 (N_3354,In_570,In_375);
or U3355 (N_3355,In_68,In_151);
xnor U3356 (N_3356,In_173,In_213);
nand U3357 (N_3357,In_199,In_295);
or U3358 (N_3358,In_729,In_455);
or U3359 (N_3359,In_598,In_758);
or U3360 (N_3360,In_657,In_829);
nor U3361 (N_3361,In_479,In_543);
nand U3362 (N_3362,In_199,In_347);
nor U3363 (N_3363,In_870,In_391);
nand U3364 (N_3364,In_871,In_989);
or U3365 (N_3365,In_578,In_497);
xor U3366 (N_3366,In_754,In_672);
nand U3367 (N_3367,In_209,In_518);
and U3368 (N_3368,In_388,In_267);
nand U3369 (N_3369,In_6,In_276);
nand U3370 (N_3370,In_405,In_150);
nand U3371 (N_3371,In_522,In_109);
or U3372 (N_3372,In_122,In_714);
or U3373 (N_3373,In_472,In_919);
and U3374 (N_3374,In_678,In_898);
or U3375 (N_3375,In_61,In_737);
or U3376 (N_3376,In_778,In_996);
nor U3377 (N_3377,In_492,In_889);
nor U3378 (N_3378,In_464,In_145);
nor U3379 (N_3379,In_8,In_522);
and U3380 (N_3380,In_92,In_829);
or U3381 (N_3381,In_184,In_19);
or U3382 (N_3382,In_804,In_891);
nor U3383 (N_3383,In_486,In_817);
nor U3384 (N_3384,In_656,In_550);
nor U3385 (N_3385,In_943,In_58);
and U3386 (N_3386,In_973,In_783);
nor U3387 (N_3387,In_581,In_663);
or U3388 (N_3388,In_949,In_892);
nand U3389 (N_3389,In_769,In_580);
nand U3390 (N_3390,In_531,In_528);
or U3391 (N_3391,In_82,In_922);
or U3392 (N_3392,In_348,In_275);
or U3393 (N_3393,In_238,In_630);
nor U3394 (N_3394,In_681,In_662);
nand U3395 (N_3395,In_424,In_500);
nor U3396 (N_3396,In_201,In_838);
nor U3397 (N_3397,In_517,In_25);
and U3398 (N_3398,In_58,In_568);
or U3399 (N_3399,In_355,In_855);
and U3400 (N_3400,In_906,In_899);
nor U3401 (N_3401,In_537,In_930);
or U3402 (N_3402,In_703,In_55);
nor U3403 (N_3403,In_118,In_517);
or U3404 (N_3404,In_795,In_173);
xnor U3405 (N_3405,In_773,In_113);
or U3406 (N_3406,In_755,In_626);
or U3407 (N_3407,In_692,In_63);
nor U3408 (N_3408,In_603,In_347);
nor U3409 (N_3409,In_811,In_450);
nor U3410 (N_3410,In_500,In_145);
or U3411 (N_3411,In_510,In_374);
and U3412 (N_3412,In_803,In_892);
nor U3413 (N_3413,In_194,In_981);
xnor U3414 (N_3414,In_743,In_180);
and U3415 (N_3415,In_16,In_308);
nor U3416 (N_3416,In_961,In_308);
and U3417 (N_3417,In_506,In_567);
and U3418 (N_3418,In_982,In_65);
nand U3419 (N_3419,In_677,In_339);
or U3420 (N_3420,In_94,In_800);
or U3421 (N_3421,In_56,In_650);
nor U3422 (N_3422,In_277,In_146);
nor U3423 (N_3423,In_771,In_841);
or U3424 (N_3424,In_660,In_45);
or U3425 (N_3425,In_52,In_192);
and U3426 (N_3426,In_310,In_757);
and U3427 (N_3427,In_793,In_975);
or U3428 (N_3428,In_865,In_573);
nor U3429 (N_3429,In_382,In_128);
and U3430 (N_3430,In_685,In_803);
xnor U3431 (N_3431,In_557,In_447);
nor U3432 (N_3432,In_529,In_984);
and U3433 (N_3433,In_20,In_518);
and U3434 (N_3434,In_970,In_62);
nand U3435 (N_3435,In_878,In_658);
nor U3436 (N_3436,In_179,In_987);
xnor U3437 (N_3437,In_639,In_469);
nand U3438 (N_3438,In_405,In_963);
nor U3439 (N_3439,In_45,In_822);
nand U3440 (N_3440,In_170,In_264);
and U3441 (N_3441,In_553,In_365);
and U3442 (N_3442,In_782,In_408);
nand U3443 (N_3443,In_309,In_347);
and U3444 (N_3444,In_712,In_858);
nor U3445 (N_3445,In_394,In_590);
or U3446 (N_3446,In_60,In_59);
nand U3447 (N_3447,In_29,In_835);
or U3448 (N_3448,In_552,In_824);
nor U3449 (N_3449,In_307,In_313);
or U3450 (N_3450,In_645,In_273);
or U3451 (N_3451,In_211,In_577);
or U3452 (N_3452,In_664,In_285);
and U3453 (N_3453,In_722,In_220);
and U3454 (N_3454,In_436,In_773);
nand U3455 (N_3455,In_90,In_360);
or U3456 (N_3456,In_875,In_114);
nand U3457 (N_3457,In_89,In_115);
and U3458 (N_3458,In_57,In_929);
and U3459 (N_3459,In_964,In_857);
and U3460 (N_3460,In_417,In_300);
or U3461 (N_3461,In_454,In_49);
or U3462 (N_3462,In_907,In_81);
nand U3463 (N_3463,In_835,In_905);
or U3464 (N_3464,In_40,In_947);
nand U3465 (N_3465,In_125,In_109);
xnor U3466 (N_3466,In_373,In_209);
and U3467 (N_3467,In_550,In_165);
nand U3468 (N_3468,In_776,In_493);
and U3469 (N_3469,In_690,In_733);
and U3470 (N_3470,In_422,In_453);
and U3471 (N_3471,In_712,In_578);
or U3472 (N_3472,In_3,In_300);
and U3473 (N_3473,In_207,In_552);
and U3474 (N_3474,In_285,In_269);
nor U3475 (N_3475,In_530,In_676);
or U3476 (N_3476,In_281,In_466);
or U3477 (N_3477,In_521,In_491);
or U3478 (N_3478,In_386,In_891);
nand U3479 (N_3479,In_873,In_255);
xor U3480 (N_3480,In_955,In_658);
and U3481 (N_3481,In_660,In_861);
nand U3482 (N_3482,In_560,In_806);
or U3483 (N_3483,In_696,In_520);
nor U3484 (N_3484,In_570,In_120);
or U3485 (N_3485,In_44,In_377);
or U3486 (N_3486,In_313,In_471);
nand U3487 (N_3487,In_556,In_95);
nor U3488 (N_3488,In_392,In_584);
nand U3489 (N_3489,In_591,In_218);
and U3490 (N_3490,In_159,In_630);
nor U3491 (N_3491,In_961,In_542);
nor U3492 (N_3492,In_48,In_957);
and U3493 (N_3493,In_641,In_731);
or U3494 (N_3494,In_572,In_521);
nand U3495 (N_3495,In_469,In_567);
and U3496 (N_3496,In_251,In_524);
or U3497 (N_3497,In_925,In_200);
or U3498 (N_3498,In_284,In_952);
nor U3499 (N_3499,In_354,In_730);
or U3500 (N_3500,In_125,In_794);
and U3501 (N_3501,In_123,In_877);
nand U3502 (N_3502,In_446,In_47);
xnor U3503 (N_3503,In_405,In_0);
nand U3504 (N_3504,In_695,In_959);
nor U3505 (N_3505,In_374,In_779);
nand U3506 (N_3506,In_216,In_347);
nand U3507 (N_3507,In_365,In_276);
and U3508 (N_3508,In_527,In_135);
or U3509 (N_3509,In_338,In_546);
nand U3510 (N_3510,In_267,In_531);
or U3511 (N_3511,In_738,In_275);
or U3512 (N_3512,In_203,In_473);
or U3513 (N_3513,In_468,In_432);
nand U3514 (N_3514,In_911,In_268);
xor U3515 (N_3515,In_195,In_987);
nand U3516 (N_3516,In_221,In_680);
and U3517 (N_3517,In_720,In_284);
and U3518 (N_3518,In_752,In_484);
nand U3519 (N_3519,In_176,In_483);
xnor U3520 (N_3520,In_903,In_859);
nor U3521 (N_3521,In_974,In_175);
nor U3522 (N_3522,In_473,In_703);
nor U3523 (N_3523,In_705,In_855);
xnor U3524 (N_3524,In_937,In_433);
and U3525 (N_3525,In_567,In_138);
nand U3526 (N_3526,In_265,In_261);
nor U3527 (N_3527,In_442,In_58);
or U3528 (N_3528,In_926,In_977);
nor U3529 (N_3529,In_507,In_936);
nor U3530 (N_3530,In_786,In_250);
xnor U3531 (N_3531,In_236,In_574);
nand U3532 (N_3532,In_548,In_915);
and U3533 (N_3533,In_407,In_904);
or U3534 (N_3534,In_60,In_266);
and U3535 (N_3535,In_585,In_791);
nor U3536 (N_3536,In_118,In_541);
nand U3537 (N_3537,In_865,In_862);
nor U3538 (N_3538,In_551,In_498);
and U3539 (N_3539,In_599,In_193);
or U3540 (N_3540,In_435,In_562);
nand U3541 (N_3541,In_266,In_978);
or U3542 (N_3542,In_120,In_846);
nand U3543 (N_3543,In_692,In_980);
nand U3544 (N_3544,In_163,In_120);
and U3545 (N_3545,In_202,In_717);
nor U3546 (N_3546,In_528,In_330);
and U3547 (N_3547,In_52,In_715);
nand U3548 (N_3548,In_695,In_701);
or U3549 (N_3549,In_982,In_501);
nand U3550 (N_3550,In_262,In_234);
or U3551 (N_3551,In_802,In_725);
or U3552 (N_3552,In_125,In_769);
or U3553 (N_3553,In_702,In_959);
nand U3554 (N_3554,In_129,In_263);
or U3555 (N_3555,In_922,In_557);
nor U3556 (N_3556,In_12,In_931);
nand U3557 (N_3557,In_828,In_942);
or U3558 (N_3558,In_678,In_788);
and U3559 (N_3559,In_436,In_465);
or U3560 (N_3560,In_914,In_256);
nand U3561 (N_3561,In_109,In_147);
nor U3562 (N_3562,In_453,In_287);
xor U3563 (N_3563,In_245,In_168);
nand U3564 (N_3564,In_965,In_947);
or U3565 (N_3565,In_641,In_935);
nand U3566 (N_3566,In_886,In_221);
or U3567 (N_3567,In_999,In_87);
or U3568 (N_3568,In_74,In_643);
and U3569 (N_3569,In_897,In_837);
or U3570 (N_3570,In_945,In_875);
or U3571 (N_3571,In_234,In_386);
or U3572 (N_3572,In_24,In_860);
and U3573 (N_3573,In_543,In_842);
or U3574 (N_3574,In_72,In_289);
or U3575 (N_3575,In_79,In_767);
or U3576 (N_3576,In_599,In_917);
or U3577 (N_3577,In_134,In_607);
nor U3578 (N_3578,In_632,In_346);
or U3579 (N_3579,In_916,In_100);
xor U3580 (N_3580,In_915,In_746);
and U3581 (N_3581,In_680,In_287);
nand U3582 (N_3582,In_864,In_477);
and U3583 (N_3583,In_198,In_64);
or U3584 (N_3584,In_626,In_433);
or U3585 (N_3585,In_283,In_711);
nor U3586 (N_3586,In_983,In_523);
nand U3587 (N_3587,In_897,In_278);
or U3588 (N_3588,In_552,In_619);
xor U3589 (N_3589,In_903,In_536);
nor U3590 (N_3590,In_11,In_516);
xor U3591 (N_3591,In_813,In_860);
nand U3592 (N_3592,In_916,In_844);
nand U3593 (N_3593,In_718,In_278);
or U3594 (N_3594,In_718,In_781);
or U3595 (N_3595,In_968,In_395);
or U3596 (N_3596,In_505,In_39);
or U3597 (N_3597,In_998,In_621);
nand U3598 (N_3598,In_603,In_500);
nor U3599 (N_3599,In_954,In_808);
or U3600 (N_3600,In_777,In_731);
nor U3601 (N_3601,In_239,In_236);
and U3602 (N_3602,In_148,In_320);
nor U3603 (N_3603,In_496,In_635);
nand U3604 (N_3604,In_15,In_990);
and U3605 (N_3605,In_566,In_273);
xor U3606 (N_3606,In_356,In_508);
and U3607 (N_3607,In_980,In_451);
and U3608 (N_3608,In_697,In_262);
nand U3609 (N_3609,In_344,In_972);
nor U3610 (N_3610,In_11,In_511);
nor U3611 (N_3611,In_394,In_605);
or U3612 (N_3612,In_954,In_96);
or U3613 (N_3613,In_622,In_597);
nor U3614 (N_3614,In_50,In_861);
nand U3615 (N_3615,In_805,In_874);
nand U3616 (N_3616,In_209,In_972);
or U3617 (N_3617,In_44,In_820);
or U3618 (N_3618,In_630,In_744);
nand U3619 (N_3619,In_505,In_273);
nor U3620 (N_3620,In_785,In_564);
nand U3621 (N_3621,In_39,In_829);
nand U3622 (N_3622,In_944,In_563);
and U3623 (N_3623,In_943,In_430);
nor U3624 (N_3624,In_128,In_992);
or U3625 (N_3625,In_628,In_384);
and U3626 (N_3626,In_91,In_415);
nand U3627 (N_3627,In_560,In_224);
nand U3628 (N_3628,In_869,In_852);
nand U3629 (N_3629,In_413,In_544);
and U3630 (N_3630,In_993,In_385);
or U3631 (N_3631,In_132,In_558);
nor U3632 (N_3632,In_119,In_691);
nor U3633 (N_3633,In_768,In_653);
nor U3634 (N_3634,In_233,In_873);
and U3635 (N_3635,In_182,In_460);
and U3636 (N_3636,In_199,In_502);
nor U3637 (N_3637,In_238,In_13);
or U3638 (N_3638,In_161,In_285);
nor U3639 (N_3639,In_497,In_996);
or U3640 (N_3640,In_476,In_509);
and U3641 (N_3641,In_367,In_439);
nand U3642 (N_3642,In_115,In_772);
nor U3643 (N_3643,In_324,In_440);
nor U3644 (N_3644,In_388,In_22);
nand U3645 (N_3645,In_804,In_808);
nand U3646 (N_3646,In_511,In_264);
nor U3647 (N_3647,In_255,In_640);
or U3648 (N_3648,In_432,In_489);
nor U3649 (N_3649,In_684,In_946);
nor U3650 (N_3650,In_349,In_288);
nor U3651 (N_3651,In_782,In_17);
nor U3652 (N_3652,In_76,In_373);
or U3653 (N_3653,In_671,In_380);
nor U3654 (N_3654,In_788,In_401);
and U3655 (N_3655,In_456,In_948);
and U3656 (N_3656,In_513,In_567);
or U3657 (N_3657,In_823,In_548);
or U3658 (N_3658,In_992,In_83);
and U3659 (N_3659,In_59,In_751);
nor U3660 (N_3660,In_892,In_927);
and U3661 (N_3661,In_577,In_421);
or U3662 (N_3662,In_206,In_121);
or U3663 (N_3663,In_645,In_455);
and U3664 (N_3664,In_607,In_96);
or U3665 (N_3665,In_383,In_227);
or U3666 (N_3666,In_574,In_768);
nand U3667 (N_3667,In_302,In_51);
and U3668 (N_3668,In_169,In_745);
and U3669 (N_3669,In_849,In_182);
or U3670 (N_3670,In_767,In_811);
and U3671 (N_3671,In_523,In_327);
nor U3672 (N_3672,In_450,In_23);
nand U3673 (N_3673,In_881,In_976);
nand U3674 (N_3674,In_90,In_785);
nor U3675 (N_3675,In_145,In_657);
and U3676 (N_3676,In_494,In_323);
or U3677 (N_3677,In_636,In_121);
nand U3678 (N_3678,In_686,In_248);
xor U3679 (N_3679,In_8,In_600);
or U3680 (N_3680,In_847,In_528);
or U3681 (N_3681,In_119,In_777);
or U3682 (N_3682,In_939,In_32);
and U3683 (N_3683,In_250,In_389);
nor U3684 (N_3684,In_417,In_459);
nand U3685 (N_3685,In_578,In_229);
and U3686 (N_3686,In_944,In_469);
xnor U3687 (N_3687,In_288,In_784);
and U3688 (N_3688,In_420,In_69);
or U3689 (N_3689,In_247,In_936);
nor U3690 (N_3690,In_592,In_251);
or U3691 (N_3691,In_591,In_30);
nor U3692 (N_3692,In_597,In_558);
and U3693 (N_3693,In_843,In_399);
and U3694 (N_3694,In_940,In_345);
or U3695 (N_3695,In_953,In_819);
nor U3696 (N_3696,In_671,In_728);
nand U3697 (N_3697,In_105,In_989);
or U3698 (N_3698,In_956,In_858);
nor U3699 (N_3699,In_380,In_878);
and U3700 (N_3700,In_352,In_750);
nor U3701 (N_3701,In_330,In_107);
and U3702 (N_3702,In_135,In_2);
and U3703 (N_3703,In_448,In_959);
or U3704 (N_3704,In_541,In_99);
nor U3705 (N_3705,In_593,In_186);
or U3706 (N_3706,In_556,In_49);
nand U3707 (N_3707,In_415,In_658);
and U3708 (N_3708,In_433,In_237);
and U3709 (N_3709,In_37,In_304);
or U3710 (N_3710,In_669,In_846);
and U3711 (N_3711,In_425,In_357);
nor U3712 (N_3712,In_222,In_711);
or U3713 (N_3713,In_285,In_900);
or U3714 (N_3714,In_823,In_145);
and U3715 (N_3715,In_180,In_912);
and U3716 (N_3716,In_118,In_28);
nand U3717 (N_3717,In_676,In_188);
xnor U3718 (N_3718,In_799,In_39);
nand U3719 (N_3719,In_297,In_324);
nor U3720 (N_3720,In_745,In_51);
and U3721 (N_3721,In_385,In_899);
nand U3722 (N_3722,In_82,In_657);
and U3723 (N_3723,In_425,In_711);
or U3724 (N_3724,In_451,In_764);
nand U3725 (N_3725,In_176,In_102);
nand U3726 (N_3726,In_859,In_657);
or U3727 (N_3727,In_9,In_174);
nor U3728 (N_3728,In_435,In_684);
nand U3729 (N_3729,In_487,In_392);
and U3730 (N_3730,In_783,In_241);
nor U3731 (N_3731,In_754,In_346);
and U3732 (N_3732,In_459,In_678);
or U3733 (N_3733,In_690,In_153);
and U3734 (N_3734,In_378,In_773);
nand U3735 (N_3735,In_486,In_405);
nor U3736 (N_3736,In_480,In_47);
nor U3737 (N_3737,In_161,In_746);
nand U3738 (N_3738,In_324,In_438);
nor U3739 (N_3739,In_138,In_181);
and U3740 (N_3740,In_260,In_608);
or U3741 (N_3741,In_89,In_3);
nor U3742 (N_3742,In_653,In_761);
nor U3743 (N_3743,In_243,In_941);
nor U3744 (N_3744,In_198,In_589);
nand U3745 (N_3745,In_41,In_653);
nor U3746 (N_3746,In_111,In_258);
nand U3747 (N_3747,In_127,In_280);
nor U3748 (N_3748,In_269,In_39);
nor U3749 (N_3749,In_714,In_351);
or U3750 (N_3750,In_105,In_878);
and U3751 (N_3751,In_968,In_932);
and U3752 (N_3752,In_888,In_733);
or U3753 (N_3753,In_16,In_206);
nor U3754 (N_3754,In_491,In_501);
or U3755 (N_3755,In_776,In_885);
or U3756 (N_3756,In_709,In_30);
nand U3757 (N_3757,In_823,In_433);
nor U3758 (N_3758,In_959,In_823);
nor U3759 (N_3759,In_878,In_840);
nor U3760 (N_3760,In_237,In_177);
or U3761 (N_3761,In_510,In_791);
or U3762 (N_3762,In_860,In_730);
or U3763 (N_3763,In_767,In_91);
nand U3764 (N_3764,In_851,In_302);
or U3765 (N_3765,In_485,In_533);
nand U3766 (N_3766,In_618,In_992);
or U3767 (N_3767,In_332,In_241);
or U3768 (N_3768,In_532,In_305);
or U3769 (N_3769,In_612,In_854);
nor U3770 (N_3770,In_480,In_851);
or U3771 (N_3771,In_408,In_751);
and U3772 (N_3772,In_433,In_172);
nand U3773 (N_3773,In_704,In_461);
nand U3774 (N_3774,In_997,In_471);
or U3775 (N_3775,In_287,In_33);
nand U3776 (N_3776,In_689,In_78);
nand U3777 (N_3777,In_127,In_780);
or U3778 (N_3778,In_909,In_65);
nor U3779 (N_3779,In_288,In_778);
nor U3780 (N_3780,In_858,In_911);
nand U3781 (N_3781,In_355,In_539);
and U3782 (N_3782,In_693,In_686);
and U3783 (N_3783,In_709,In_713);
nor U3784 (N_3784,In_338,In_173);
and U3785 (N_3785,In_712,In_256);
nand U3786 (N_3786,In_939,In_960);
or U3787 (N_3787,In_563,In_768);
nand U3788 (N_3788,In_794,In_439);
and U3789 (N_3789,In_934,In_141);
nor U3790 (N_3790,In_469,In_858);
nor U3791 (N_3791,In_322,In_863);
nand U3792 (N_3792,In_986,In_873);
nand U3793 (N_3793,In_428,In_193);
nor U3794 (N_3794,In_24,In_184);
nand U3795 (N_3795,In_790,In_445);
and U3796 (N_3796,In_923,In_976);
nor U3797 (N_3797,In_90,In_869);
and U3798 (N_3798,In_839,In_968);
or U3799 (N_3799,In_397,In_63);
and U3800 (N_3800,In_705,In_121);
and U3801 (N_3801,In_543,In_547);
nor U3802 (N_3802,In_259,In_869);
nor U3803 (N_3803,In_68,In_351);
nand U3804 (N_3804,In_920,In_996);
or U3805 (N_3805,In_561,In_898);
and U3806 (N_3806,In_580,In_152);
or U3807 (N_3807,In_45,In_443);
nor U3808 (N_3808,In_847,In_419);
nor U3809 (N_3809,In_329,In_234);
or U3810 (N_3810,In_211,In_40);
and U3811 (N_3811,In_724,In_310);
or U3812 (N_3812,In_577,In_744);
or U3813 (N_3813,In_223,In_305);
or U3814 (N_3814,In_298,In_314);
nand U3815 (N_3815,In_894,In_819);
nand U3816 (N_3816,In_710,In_538);
nand U3817 (N_3817,In_964,In_569);
nor U3818 (N_3818,In_177,In_212);
or U3819 (N_3819,In_953,In_442);
or U3820 (N_3820,In_644,In_121);
or U3821 (N_3821,In_820,In_43);
or U3822 (N_3822,In_184,In_70);
nor U3823 (N_3823,In_345,In_110);
or U3824 (N_3824,In_645,In_699);
or U3825 (N_3825,In_569,In_205);
and U3826 (N_3826,In_861,In_630);
nand U3827 (N_3827,In_872,In_646);
nor U3828 (N_3828,In_623,In_74);
and U3829 (N_3829,In_478,In_510);
and U3830 (N_3830,In_866,In_197);
nor U3831 (N_3831,In_58,In_454);
nor U3832 (N_3832,In_732,In_803);
nor U3833 (N_3833,In_593,In_460);
nand U3834 (N_3834,In_588,In_305);
or U3835 (N_3835,In_434,In_960);
nand U3836 (N_3836,In_363,In_216);
nand U3837 (N_3837,In_189,In_236);
nand U3838 (N_3838,In_543,In_421);
nand U3839 (N_3839,In_771,In_423);
and U3840 (N_3840,In_764,In_74);
nor U3841 (N_3841,In_884,In_180);
nor U3842 (N_3842,In_390,In_187);
or U3843 (N_3843,In_684,In_429);
and U3844 (N_3844,In_304,In_438);
nor U3845 (N_3845,In_907,In_133);
xor U3846 (N_3846,In_240,In_212);
nand U3847 (N_3847,In_43,In_605);
nor U3848 (N_3848,In_263,In_691);
nand U3849 (N_3849,In_841,In_137);
or U3850 (N_3850,In_184,In_945);
or U3851 (N_3851,In_631,In_824);
nor U3852 (N_3852,In_516,In_445);
nor U3853 (N_3853,In_895,In_451);
or U3854 (N_3854,In_387,In_492);
nor U3855 (N_3855,In_719,In_607);
and U3856 (N_3856,In_482,In_275);
nor U3857 (N_3857,In_550,In_811);
nand U3858 (N_3858,In_666,In_314);
nor U3859 (N_3859,In_351,In_602);
nand U3860 (N_3860,In_998,In_422);
or U3861 (N_3861,In_887,In_683);
nand U3862 (N_3862,In_567,In_525);
and U3863 (N_3863,In_716,In_765);
xor U3864 (N_3864,In_535,In_412);
nand U3865 (N_3865,In_720,In_252);
nand U3866 (N_3866,In_123,In_675);
nor U3867 (N_3867,In_315,In_769);
or U3868 (N_3868,In_41,In_360);
nand U3869 (N_3869,In_746,In_619);
nand U3870 (N_3870,In_571,In_954);
nand U3871 (N_3871,In_383,In_728);
nor U3872 (N_3872,In_372,In_106);
and U3873 (N_3873,In_531,In_49);
nand U3874 (N_3874,In_965,In_167);
nand U3875 (N_3875,In_508,In_875);
or U3876 (N_3876,In_774,In_335);
nand U3877 (N_3877,In_604,In_865);
nand U3878 (N_3878,In_997,In_826);
or U3879 (N_3879,In_620,In_111);
and U3880 (N_3880,In_423,In_967);
or U3881 (N_3881,In_981,In_658);
nand U3882 (N_3882,In_564,In_162);
or U3883 (N_3883,In_330,In_979);
or U3884 (N_3884,In_543,In_71);
or U3885 (N_3885,In_338,In_957);
and U3886 (N_3886,In_383,In_87);
and U3887 (N_3887,In_585,In_567);
xor U3888 (N_3888,In_826,In_955);
and U3889 (N_3889,In_812,In_256);
and U3890 (N_3890,In_836,In_869);
or U3891 (N_3891,In_756,In_713);
and U3892 (N_3892,In_987,In_543);
or U3893 (N_3893,In_948,In_510);
nand U3894 (N_3894,In_428,In_262);
or U3895 (N_3895,In_65,In_679);
nor U3896 (N_3896,In_702,In_815);
nand U3897 (N_3897,In_914,In_762);
nand U3898 (N_3898,In_459,In_515);
nand U3899 (N_3899,In_674,In_459);
nor U3900 (N_3900,In_769,In_156);
nor U3901 (N_3901,In_850,In_428);
and U3902 (N_3902,In_573,In_725);
nand U3903 (N_3903,In_783,In_339);
nor U3904 (N_3904,In_978,In_472);
nor U3905 (N_3905,In_886,In_732);
or U3906 (N_3906,In_509,In_858);
and U3907 (N_3907,In_909,In_75);
or U3908 (N_3908,In_12,In_620);
or U3909 (N_3909,In_342,In_706);
nor U3910 (N_3910,In_469,In_537);
nor U3911 (N_3911,In_930,In_693);
or U3912 (N_3912,In_305,In_584);
nand U3913 (N_3913,In_465,In_835);
or U3914 (N_3914,In_50,In_512);
nand U3915 (N_3915,In_54,In_952);
nand U3916 (N_3916,In_958,In_602);
nor U3917 (N_3917,In_90,In_900);
nand U3918 (N_3918,In_770,In_583);
and U3919 (N_3919,In_873,In_595);
nand U3920 (N_3920,In_254,In_812);
or U3921 (N_3921,In_501,In_187);
and U3922 (N_3922,In_923,In_359);
or U3923 (N_3923,In_217,In_254);
nand U3924 (N_3924,In_189,In_857);
nor U3925 (N_3925,In_454,In_237);
nand U3926 (N_3926,In_570,In_256);
nand U3927 (N_3927,In_192,In_573);
and U3928 (N_3928,In_230,In_167);
nand U3929 (N_3929,In_360,In_237);
and U3930 (N_3930,In_172,In_798);
nor U3931 (N_3931,In_107,In_130);
and U3932 (N_3932,In_390,In_862);
or U3933 (N_3933,In_762,In_477);
and U3934 (N_3934,In_244,In_906);
nor U3935 (N_3935,In_175,In_348);
or U3936 (N_3936,In_695,In_746);
and U3937 (N_3937,In_815,In_822);
nor U3938 (N_3938,In_401,In_204);
or U3939 (N_3939,In_906,In_774);
and U3940 (N_3940,In_708,In_87);
or U3941 (N_3941,In_52,In_731);
nand U3942 (N_3942,In_306,In_594);
and U3943 (N_3943,In_185,In_476);
nand U3944 (N_3944,In_127,In_897);
or U3945 (N_3945,In_486,In_794);
and U3946 (N_3946,In_937,In_957);
and U3947 (N_3947,In_800,In_894);
nor U3948 (N_3948,In_788,In_964);
and U3949 (N_3949,In_935,In_970);
nand U3950 (N_3950,In_20,In_224);
nor U3951 (N_3951,In_735,In_154);
or U3952 (N_3952,In_931,In_861);
or U3953 (N_3953,In_131,In_299);
xor U3954 (N_3954,In_922,In_68);
and U3955 (N_3955,In_911,In_590);
and U3956 (N_3956,In_948,In_986);
and U3957 (N_3957,In_885,In_507);
nand U3958 (N_3958,In_405,In_615);
or U3959 (N_3959,In_593,In_152);
or U3960 (N_3960,In_947,In_250);
or U3961 (N_3961,In_367,In_546);
and U3962 (N_3962,In_79,In_440);
nor U3963 (N_3963,In_245,In_953);
nor U3964 (N_3964,In_91,In_96);
and U3965 (N_3965,In_717,In_333);
or U3966 (N_3966,In_214,In_624);
and U3967 (N_3967,In_501,In_306);
and U3968 (N_3968,In_841,In_557);
nand U3969 (N_3969,In_276,In_958);
and U3970 (N_3970,In_792,In_183);
or U3971 (N_3971,In_112,In_924);
or U3972 (N_3972,In_690,In_225);
or U3973 (N_3973,In_577,In_74);
and U3974 (N_3974,In_156,In_5);
nand U3975 (N_3975,In_740,In_598);
xnor U3976 (N_3976,In_561,In_598);
xnor U3977 (N_3977,In_165,In_594);
and U3978 (N_3978,In_8,In_231);
or U3979 (N_3979,In_502,In_610);
and U3980 (N_3980,In_514,In_668);
or U3981 (N_3981,In_453,In_914);
nand U3982 (N_3982,In_479,In_307);
nand U3983 (N_3983,In_492,In_720);
nor U3984 (N_3984,In_149,In_410);
xnor U3985 (N_3985,In_297,In_480);
or U3986 (N_3986,In_957,In_417);
and U3987 (N_3987,In_867,In_740);
and U3988 (N_3988,In_425,In_888);
and U3989 (N_3989,In_932,In_918);
nor U3990 (N_3990,In_508,In_583);
and U3991 (N_3991,In_386,In_84);
or U3992 (N_3992,In_523,In_816);
and U3993 (N_3993,In_56,In_205);
and U3994 (N_3994,In_418,In_577);
nor U3995 (N_3995,In_228,In_225);
or U3996 (N_3996,In_522,In_340);
nand U3997 (N_3997,In_430,In_662);
or U3998 (N_3998,In_227,In_902);
nor U3999 (N_3999,In_540,In_292);
and U4000 (N_4000,In_800,In_29);
and U4001 (N_4001,In_503,In_496);
and U4002 (N_4002,In_696,In_712);
or U4003 (N_4003,In_233,In_356);
nand U4004 (N_4004,In_548,In_812);
and U4005 (N_4005,In_465,In_238);
and U4006 (N_4006,In_719,In_429);
nand U4007 (N_4007,In_746,In_95);
nor U4008 (N_4008,In_251,In_464);
xor U4009 (N_4009,In_396,In_38);
and U4010 (N_4010,In_842,In_56);
nand U4011 (N_4011,In_12,In_782);
nand U4012 (N_4012,In_687,In_641);
or U4013 (N_4013,In_854,In_398);
nand U4014 (N_4014,In_24,In_67);
nor U4015 (N_4015,In_741,In_852);
and U4016 (N_4016,In_913,In_946);
or U4017 (N_4017,In_994,In_891);
nand U4018 (N_4018,In_490,In_15);
nor U4019 (N_4019,In_751,In_968);
or U4020 (N_4020,In_22,In_275);
and U4021 (N_4021,In_250,In_19);
nor U4022 (N_4022,In_53,In_293);
nand U4023 (N_4023,In_276,In_209);
nor U4024 (N_4024,In_146,In_254);
xnor U4025 (N_4025,In_92,In_5);
and U4026 (N_4026,In_37,In_274);
nand U4027 (N_4027,In_644,In_906);
and U4028 (N_4028,In_521,In_571);
or U4029 (N_4029,In_274,In_520);
nand U4030 (N_4030,In_502,In_251);
or U4031 (N_4031,In_620,In_748);
or U4032 (N_4032,In_866,In_348);
nor U4033 (N_4033,In_536,In_426);
xor U4034 (N_4034,In_37,In_296);
nand U4035 (N_4035,In_686,In_237);
and U4036 (N_4036,In_11,In_369);
nor U4037 (N_4037,In_747,In_225);
nor U4038 (N_4038,In_818,In_146);
or U4039 (N_4039,In_737,In_523);
or U4040 (N_4040,In_150,In_846);
nor U4041 (N_4041,In_868,In_677);
or U4042 (N_4042,In_99,In_915);
and U4043 (N_4043,In_123,In_811);
nand U4044 (N_4044,In_99,In_291);
xnor U4045 (N_4045,In_155,In_223);
nor U4046 (N_4046,In_763,In_153);
or U4047 (N_4047,In_181,In_386);
nand U4048 (N_4048,In_517,In_256);
nand U4049 (N_4049,In_892,In_828);
nand U4050 (N_4050,In_550,In_181);
and U4051 (N_4051,In_78,In_597);
xnor U4052 (N_4052,In_940,In_390);
or U4053 (N_4053,In_789,In_204);
nor U4054 (N_4054,In_61,In_776);
or U4055 (N_4055,In_673,In_516);
nor U4056 (N_4056,In_937,In_272);
nor U4057 (N_4057,In_200,In_82);
or U4058 (N_4058,In_949,In_429);
and U4059 (N_4059,In_107,In_20);
and U4060 (N_4060,In_832,In_55);
nand U4061 (N_4061,In_369,In_327);
nand U4062 (N_4062,In_48,In_349);
nor U4063 (N_4063,In_441,In_65);
and U4064 (N_4064,In_308,In_236);
nor U4065 (N_4065,In_521,In_670);
nor U4066 (N_4066,In_684,In_716);
nor U4067 (N_4067,In_18,In_587);
nor U4068 (N_4068,In_496,In_157);
nor U4069 (N_4069,In_790,In_330);
nand U4070 (N_4070,In_78,In_174);
or U4071 (N_4071,In_9,In_503);
nor U4072 (N_4072,In_826,In_257);
nand U4073 (N_4073,In_599,In_218);
nand U4074 (N_4074,In_723,In_54);
or U4075 (N_4075,In_836,In_473);
and U4076 (N_4076,In_70,In_729);
and U4077 (N_4077,In_134,In_729);
or U4078 (N_4078,In_508,In_889);
and U4079 (N_4079,In_511,In_400);
and U4080 (N_4080,In_581,In_44);
xnor U4081 (N_4081,In_699,In_781);
or U4082 (N_4082,In_164,In_335);
nand U4083 (N_4083,In_95,In_62);
or U4084 (N_4084,In_681,In_471);
or U4085 (N_4085,In_769,In_400);
nand U4086 (N_4086,In_936,In_4);
nor U4087 (N_4087,In_767,In_995);
or U4088 (N_4088,In_354,In_381);
and U4089 (N_4089,In_439,In_92);
and U4090 (N_4090,In_319,In_15);
and U4091 (N_4091,In_163,In_329);
and U4092 (N_4092,In_106,In_280);
and U4093 (N_4093,In_812,In_187);
nand U4094 (N_4094,In_412,In_705);
nand U4095 (N_4095,In_969,In_726);
or U4096 (N_4096,In_840,In_879);
or U4097 (N_4097,In_429,In_785);
nand U4098 (N_4098,In_466,In_361);
and U4099 (N_4099,In_103,In_157);
nor U4100 (N_4100,In_64,In_303);
xnor U4101 (N_4101,In_777,In_755);
nand U4102 (N_4102,In_658,In_742);
nand U4103 (N_4103,In_793,In_642);
or U4104 (N_4104,In_454,In_90);
nand U4105 (N_4105,In_659,In_0);
or U4106 (N_4106,In_889,In_607);
or U4107 (N_4107,In_58,In_985);
and U4108 (N_4108,In_254,In_468);
nand U4109 (N_4109,In_3,In_583);
nor U4110 (N_4110,In_682,In_512);
nand U4111 (N_4111,In_763,In_191);
or U4112 (N_4112,In_62,In_354);
and U4113 (N_4113,In_180,In_18);
or U4114 (N_4114,In_451,In_610);
and U4115 (N_4115,In_462,In_579);
xor U4116 (N_4116,In_178,In_889);
and U4117 (N_4117,In_25,In_480);
nand U4118 (N_4118,In_60,In_408);
nand U4119 (N_4119,In_348,In_217);
and U4120 (N_4120,In_96,In_998);
or U4121 (N_4121,In_220,In_6);
nor U4122 (N_4122,In_989,In_446);
nor U4123 (N_4123,In_104,In_556);
nor U4124 (N_4124,In_698,In_319);
nand U4125 (N_4125,In_392,In_106);
or U4126 (N_4126,In_281,In_80);
and U4127 (N_4127,In_127,In_728);
nand U4128 (N_4128,In_357,In_660);
nand U4129 (N_4129,In_154,In_46);
xnor U4130 (N_4130,In_435,In_291);
nor U4131 (N_4131,In_979,In_774);
nand U4132 (N_4132,In_554,In_621);
and U4133 (N_4133,In_542,In_310);
or U4134 (N_4134,In_966,In_679);
or U4135 (N_4135,In_387,In_471);
xor U4136 (N_4136,In_162,In_710);
nand U4137 (N_4137,In_838,In_427);
nand U4138 (N_4138,In_371,In_110);
nor U4139 (N_4139,In_730,In_950);
nand U4140 (N_4140,In_131,In_264);
nor U4141 (N_4141,In_940,In_931);
nor U4142 (N_4142,In_483,In_498);
nand U4143 (N_4143,In_41,In_191);
nand U4144 (N_4144,In_611,In_980);
or U4145 (N_4145,In_630,In_628);
and U4146 (N_4146,In_46,In_276);
xor U4147 (N_4147,In_904,In_697);
or U4148 (N_4148,In_639,In_669);
nand U4149 (N_4149,In_770,In_624);
and U4150 (N_4150,In_827,In_241);
nand U4151 (N_4151,In_807,In_900);
or U4152 (N_4152,In_271,In_51);
and U4153 (N_4153,In_326,In_128);
or U4154 (N_4154,In_750,In_596);
nand U4155 (N_4155,In_381,In_426);
nand U4156 (N_4156,In_91,In_584);
or U4157 (N_4157,In_135,In_624);
or U4158 (N_4158,In_824,In_130);
and U4159 (N_4159,In_200,In_867);
nor U4160 (N_4160,In_163,In_78);
nand U4161 (N_4161,In_482,In_166);
or U4162 (N_4162,In_284,In_853);
or U4163 (N_4163,In_361,In_659);
and U4164 (N_4164,In_119,In_14);
and U4165 (N_4165,In_879,In_975);
xnor U4166 (N_4166,In_307,In_565);
and U4167 (N_4167,In_745,In_99);
or U4168 (N_4168,In_746,In_687);
nand U4169 (N_4169,In_310,In_452);
nand U4170 (N_4170,In_870,In_520);
or U4171 (N_4171,In_619,In_186);
and U4172 (N_4172,In_43,In_60);
or U4173 (N_4173,In_817,In_217);
or U4174 (N_4174,In_149,In_530);
or U4175 (N_4175,In_297,In_746);
and U4176 (N_4176,In_279,In_304);
nor U4177 (N_4177,In_232,In_607);
nor U4178 (N_4178,In_67,In_298);
or U4179 (N_4179,In_184,In_965);
and U4180 (N_4180,In_251,In_515);
nand U4181 (N_4181,In_844,In_526);
nand U4182 (N_4182,In_366,In_0);
or U4183 (N_4183,In_703,In_554);
xnor U4184 (N_4184,In_702,In_421);
and U4185 (N_4185,In_807,In_300);
nor U4186 (N_4186,In_929,In_743);
and U4187 (N_4187,In_153,In_608);
nand U4188 (N_4188,In_238,In_849);
or U4189 (N_4189,In_271,In_819);
or U4190 (N_4190,In_587,In_144);
nor U4191 (N_4191,In_350,In_549);
nand U4192 (N_4192,In_182,In_188);
nand U4193 (N_4193,In_161,In_555);
nor U4194 (N_4194,In_826,In_761);
nand U4195 (N_4195,In_753,In_534);
or U4196 (N_4196,In_408,In_580);
nor U4197 (N_4197,In_867,In_382);
nand U4198 (N_4198,In_158,In_912);
nand U4199 (N_4199,In_304,In_33);
or U4200 (N_4200,In_514,In_273);
nor U4201 (N_4201,In_824,In_282);
and U4202 (N_4202,In_929,In_145);
nand U4203 (N_4203,In_25,In_936);
and U4204 (N_4204,In_745,In_421);
nand U4205 (N_4205,In_490,In_529);
nand U4206 (N_4206,In_261,In_954);
nor U4207 (N_4207,In_393,In_315);
nand U4208 (N_4208,In_200,In_482);
and U4209 (N_4209,In_811,In_342);
and U4210 (N_4210,In_538,In_311);
and U4211 (N_4211,In_711,In_400);
or U4212 (N_4212,In_580,In_400);
and U4213 (N_4213,In_832,In_453);
nand U4214 (N_4214,In_150,In_992);
or U4215 (N_4215,In_289,In_318);
nor U4216 (N_4216,In_748,In_269);
or U4217 (N_4217,In_149,In_551);
nor U4218 (N_4218,In_67,In_643);
or U4219 (N_4219,In_196,In_578);
and U4220 (N_4220,In_35,In_635);
or U4221 (N_4221,In_100,In_522);
nor U4222 (N_4222,In_856,In_307);
nor U4223 (N_4223,In_328,In_264);
and U4224 (N_4224,In_424,In_463);
nand U4225 (N_4225,In_109,In_662);
nand U4226 (N_4226,In_994,In_584);
nand U4227 (N_4227,In_677,In_482);
or U4228 (N_4228,In_741,In_325);
nor U4229 (N_4229,In_210,In_305);
nor U4230 (N_4230,In_100,In_360);
and U4231 (N_4231,In_49,In_122);
nor U4232 (N_4232,In_544,In_789);
nor U4233 (N_4233,In_107,In_738);
xor U4234 (N_4234,In_454,In_199);
nand U4235 (N_4235,In_709,In_699);
nand U4236 (N_4236,In_42,In_800);
nor U4237 (N_4237,In_582,In_120);
nor U4238 (N_4238,In_837,In_932);
and U4239 (N_4239,In_636,In_110);
or U4240 (N_4240,In_570,In_647);
or U4241 (N_4241,In_379,In_882);
or U4242 (N_4242,In_12,In_344);
and U4243 (N_4243,In_841,In_539);
nand U4244 (N_4244,In_417,In_380);
or U4245 (N_4245,In_490,In_47);
and U4246 (N_4246,In_358,In_913);
nand U4247 (N_4247,In_654,In_75);
and U4248 (N_4248,In_548,In_44);
nand U4249 (N_4249,In_945,In_67);
and U4250 (N_4250,In_938,In_391);
nand U4251 (N_4251,In_226,In_253);
and U4252 (N_4252,In_723,In_654);
and U4253 (N_4253,In_828,In_694);
nand U4254 (N_4254,In_619,In_844);
nor U4255 (N_4255,In_583,In_488);
nor U4256 (N_4256,In_659,In_232);
or U4257 (N_4257,In_743,In_549);
nand U4258 (N_4258,In_900,In_124);
or U4259 (N_4259,In_872,In_685);
nor U4260 (N_4260,In_642,In_866);
nand U4261 (N_4261,In_691,In_759);
nand U4262 (N_4262,In_597,In_110);
nor U4263 (N_4263,In_178,In_632);
or U4264 (N_4264,In_545,In_391);
nor U4265 (N_4265,In_881,In_241);
and U4266 (N_4266,In_74,In_711);
and U4267 (N_4267,In_789,In_920);
nand U4268 (N_4268,In_254,In_857);
nand U4269 (N_4269,In_836,In_999);
nand U4270 (N_4270,In_652,In_269);
and U4271 (N_4271,In_165,In_76);
and U4272 (N_4272,In_11,In_484);
and U4273 (N_4273,In_213,In_3);
nand U4274 (N_4274,In_288,In_237);
nor U4275 (N_4275,In_907,In_350);
nand U4276 (N_4276,In_153,In_179);
xnor U4277 (N_4277,In_908,In_649);
nor U4278 (N_4278,In_390,In_927);
nor U4279 (N_4279,In_697,In_428);
nand U4280 (N_4280,In_82,In_180);
or U4281 (N_4281,In_891,In_869);
nand U4282 (N_4282,In_620,In_172);
and U4283 (N_4283,In_637,In_160);
nor U4284 (N_4284,In_320,In_523);
or U4285 (N_4285,In_856,In_809);
nor U4286 (N_4286,In_457,In_135);
nor U4287 (N_4287,In_609,In_475);
and U4288 (N_4288,In_606,In_294);
nand U4289 (N_4289,In_917,In_911);
or U4290 (N_4290,In_729,In_580);
and U4291 (N_4291,In_931,In_515);
and U4292 (N_4292,In_636,In_650);
and U4293 (N_4293,In_168,In_221);
nand U4294 (N_4294,In_82,In_439);
and U4295 (N_4295,In_716,In_432);
and U4296 (N_4296,In_518,In_12);
nor U4297 (N_4297,In_968,In_270);
nor U4298 (N_4298,In_135,In_867);
and U4299 (N_4299,In_882,In_20);
and U4300 (N_4300,In_542,In_363);
nand U4301 (N_4301,In_515,In_215);
and U4302 (N_4302,In_496,In_420);
or U4303 (N_4303,In_249,In_396);
and U4304 (N_4304,In_572,In_17);
nand U4305 (N_4305,In_869,In_89);
and U4306 (N_4306,In_40,In_307);
nand U4307 (N_4307,In_693,In_41);
nand U4308 (N_4308,In_700,In_809);
or U4309 (N_4309,In_969,In_839);
nor U4310 (N_4310,In_463,In_525);
and U4311 (N_4311,In_40,In_681);
nor U4312 (N_4312,In_640,In_105);
and U4313 (N_4313,In_389,In_623);
nand U4314 (N_4314,In_885,In_576);
and U4315 (N_4315,In_944,In_100);
nor U4316 (N_4316,In_247,In_722);
and U4317 (N_4317,In_323,In_636);
or U4318 (N_4318,In_741,In_356);
nand U4319 (N_4319,In_909,In_735);
or U4320 (N_4320,In_365,In_601);
nor U4321 (N_4321,In_890,In_779);
or U4322 (N_4322,In_861,In_631);
nand U4323 (N_4323,In_445,In_566);
or U4324 (N_4324,In_107,In_598);
nor U4325 (N_4325,In_379,In_246);
nand U4326 (N_4326,In_339,In_965);
and U4327 (N_4327,In_192,In_398);
nor U4328 (N_4328,In_218,In_80);
nand U4329 (N_4329,In_248,In_762);
nand U4330 (N_4330,In_648,In_102);
nor U4331 (N_4331,In_586,In_457);
and U4332 (N_4332,In_344,In_892);
nand U4333 (N_4333,In_323,In_531);
or U4334 (N_4334,In_871,In_437);
nor U4335 (N_4335,In_923,In_174);
nand U4336 (N_4336,In_502,In_879);
nand U4337 (N_4337,In_607,In_534);
nor U4338 (N_4338,In_137,In_987);
or U4339 (N_4339,In_6,In_947);
or U4340 (N_4340,In_92,In_644);
or U4341 (N_4341,In_990,In_931);
nor U4342 (N_4342,In_955,In_72);
nand U4343 (N_4343,In_98,In_118);
or U4344 (N_4344,In_832,In_588);
or U4345 (N_4345,In_771,In_677);
nand U4346 (N_4346,In_729,In_566);
or U4347 (N_4347,In_573,In_199);
or U4348 (N_4348,In_549,In_491);
or U4349 (N_4349,In_699,In_316);
nand U4350 (N_4350,In_741,In_969);
and U4351 (N_4351,In_635,In_864);
and U4352 (N_4352,In_71,In_499);
nand U4353 (N_4353,In_172,In_542);
and U4354 (N_4354,In_342,In_723);
or U4355 (N_4355,In_213,In_195);
or U4356 (N_4356,In_925,In_544);
and U4357 (N_4357,In_807,In_621);
nor U4358 (N_4358,In_180,In_548);
or U4359 (N_4359,In_974,In_112);
nor U4360 (N_4360,In_440,In_227);
nor U4361 (N_4361,In_517,In_519);
and U4362 (N_4362,In_324,In_855);
nor U4363 (N_4363,In_275,In_333);
or U4364 (N_4364,In_19,In_36);
or U4365 (N_4365,In_399,In_485);
nor U4366 (N_4366,In_146,In_763);
or U4367 (N_4367,In_877,In_235);
nand U4368 (N_4368,In_743,In_710);
or U4369 (N_4369,In_476,In_355);
and U4370 (N_4370,In_591,In_687);
and U4371 (N_4371,In_781,In_928);
or U4372 (N_4372,In_322,In_543);
or U4373 (N_4373,In_747,In_12);
nor U4374 (N_4374,In_884,In_93);
or U4375 (N_4375,In_996,In_809);
nand U4376 (N_4376,In_762,In_217);
or U4377 (N_4377,In_8,In_78);
nand U4378 (N_4378,In_5,In_823);
nand U4379 (N_4379,In_63,In_585);
nor U4380 (N_4380,In_141,In_23);
nor U4381 (N_4381,In_335,In_216);
nand U4382 (N_4382,In_468,In_288);
or U4383 (N_4383,In_694,In_231);
or U4384 (N_4384,In_62,In_954);
or U4385 (N_4385,In_14,In_324);
and U4386 (N_4386,In_970,In_964);
and U4387 (N_4387,In_801,In_472);
and U4388 (N_4388,In_0,In_196);
and U4389 (N_4389,In_861,In_979);
nor U4390 (N_4390,In_278,In_431);
nor U4391 (N_4391,In_4,In_947);
nor U4392 (N_4392,In_90,In_148);
nand U4393 (N_4393,In_99,In_398);
and U4394 (N_4394,In_598,In_424);
xor U4395 (N_4395,In_185,In_828);
and U4396 (N_4396,In_526,In_632);
or U4397 (N_4397,In_201,In_573);
and U4398 (N_4398,In_855,In_1);
nand U4399 (N_4399,In_221,In_971);
nand U4400 (N_4400,In_736,In_746);
or U4401 (N_4401,In_723,In_645);
and U4402 (N_4402,In_609,In_676);
nor U4403 (N_4403,In_501,In_981);
xnor U4404 (N_4404,In_283,In_67);
and U4405 (N_4405,In_863,In_375);
nor U4406 (N_4406,In_731,In_803);
nor U4407 (N_4407,In_591,In_140);
nor U4408 (N_4408,In_742,In_544);
nor U4409 (N_4409,In_48,In_884);
nor U4410 (N_4410,In_3,In_68);
and U4411 (N_4411,In_801,In_963);
and U4412 (N_4412,In_100,In_39);
nand U4413 (N_4413,In_539,In_58);
nor U4414 (N_4414,In_593,In_921);
and U4415 (N_4415,In_45,In_472);
and U4416 (N_4416,In_713,In_536);
and U4417 (N_4417,In_71,In_64);
xnor U4418 (N_4418,In_62,In_863);
and U4419 (N_4419,In_240,In_250);
and U4420 (N_4420,In_792,In_51);
and U4421 (N_4421,In_556,In_771);
nand U4422 (N_4422,In_181,In_715);
nand U4423 (N_4423,In_617,In_289);
or U4424 (N_4424,In_298,In_7);
or U4425 (N_4425,In_819,In_749);
nand U4426 (N_4426,In_254,In_797);
or U4427 (N_4427,In_676,In_733);
nor U4428 (N_4428,In_374,In_360);
nor U4429 (N_4429,In_890,In_808);
and U4430 (N_4430,In_303,In_160);
nor U4431 (N_4431,In_759,In_639);
or U4432 (N_4432,In_808,In_935);
or U4433 (N_4433,In_129,In_846);
and U4434 (N_4434,In_440,In_271);
and U4435 (N_4435,In_921,In_855);
or U4436 (N_4436,In_978,In_387);
and U4437 (N_4437,In_401,In_449);
or U4438 (N_4438,In_552,In_482);
and U4439 (N_4439,In_196,In_207);
or U4440 (N_4440,In_116,In_799);
nand U4441 (N_4441,In_433,In_513);
or U4442 (N_4442,In_630,In_24);
and U4443 (N_4443,In_560,In_90);
and U4444 (N_4444,In_934,In_137);
and U4445 (N_4445,In_647,In_990);
nor U4446 (N_4446,In_115,In_203);
nand U4447 (N_4447,In_926,In_396);
nor U4448 (N_4448,In_397,In_980);
or U4449 (N_4449,In_323,In_523);
nand U4450 (N_4450,In_274,In_412);
and U4451 (N_4451,In_420,In_385);
nand U4452 (N_4452,In_3,In_397);
nand U4453 (N_4453,In_635,In_543);
and U4454 (N_4454,In_28,In_667);
and U4455 (N_4455,In_181,In_141);
and U4456 (N_4456,In_245,In_580);
nand U4457 (N_4457,In_264,In_266);
nand U4458 (N_4458,In_203,In_463);
nand U4459 (N_4459,In_92,In_143);
nor U4460 (N_4460,In_228,In_304);
or U4461 (N_4461,In_727,In_232);
or U4462 (N_4462,In_649,In_855);
nand U4463 (N_4463,In_779,In_602);
nor U4464 (N_4464,In_961,In_95);
nor U4465 (N_4465,In_174,In_850);
or U4466 (N_4466,In_0,In_108);
or U4467 (N_4467,In_112,In_956);
nor U4468 (N_4468,In_951,In_215);
or U4469 (N_4469,In_398,In_728);
nand U4470 (N_4470,In_262,In_60);
nor U4471 (N_4471,In_807,In_792);
nor U4472 (N_4472,In_27,In_318);
or U4473 (N_4473,In_322,In_611);
and U4474 (N_4474,In_692,In_800);
nand U4475 (N_4475,In_80,In_246);
and U4476 (N_4476,In_814,In_414);
and U4477 (N_4477,In_874,In_460);
or U4478 (N_4478,In_22,In_567);
or U4479 (N_4479,In_686,In_959);
and U4480 (N_4480,In_567,In_582);
nor U4481 (N_4481,In_872,In_406);
and U4482 (N_4482,In_804,In_246);
nand U4483 (N_4483,In_478,In_792);
and U4484 (N_4484,In_622,In_898);
or U4485 (N_4485,In_133,In_662);
nor U4486 (N_4486,In_84,In_796);
or U4487 (N_4487,In_85,In_884);
nor U4488 (N_4488,In_678,In_584);
nor U4489 (N_4489,In_668,In_97);
nand U4490 (N_4490,In_37,In_368);
xnor U4491 (N_4491,In_866,In_686);
and U4492 (N_4492,In_864,In_647);
nor U4493 (N_4493,In_188,In_171);
nor U4494 (N_4494,In_568,In_942);
and U4495 (N_4495,In_923,In_220);
nand U4496 (N_4496,In_830,In_829);
nor U4497 (N_4497,In_709,In_164);
and U4498 (N_4498,In_130,In_992);
and U4499 (N_4499,In_416,In_714);
nor U4500 (N_4500,In_111,In_28);
and U4501 (N_4501,In_866,In_253);
nand U4502 (N_4502,In_450,In_28);
or U4503 (N_4503,In_312,In_46);
nor U4504 (N_4504,In_755,In_290);
nand U4505 (N_4505,In_936,In_38);
and U4506 (N_4506,In_776,In_417);
or U4507 (N_4507,In_782,In_207);
or U4508 (N_4508,In_668,In_953);
xor U4509 (N_4509,In_727,In_41);
nor U4510 (N_4510,In_396,In_625);
and U4511 (N_4511,In_452,In_261);
and U4512 (N_4512,In_682,In_508);
or U4513 (N_4513,In_306,In_985);
nand U4514 (N_4514,In_744,In_421);
nor U4515 (N_4515,In_665,In_305);
xnor U4516 (N_4516,In_819,In_584);
nor U4517 (N_4517,In_702,In_92);
or U4518 (N_4518,In_931,In_377);
and U4519 (N_4519,In_326,In_687);
nand U4520 (N_4520,In_799,In_168);
nor U4521 (N_4521,In_199,In_697);
or U4522 (N_4522,In_208,In_627);
or U4523 (N_4523,In_890,In_795);
nor U4524 (N_4524,In_975,In_846);
and U4525 (N_4525,In_323,In_879);
nor U4526 (N_4526,In_163,In_919);
and U4527 (N_4527,In_250,In_446);
and U4528 (N_4528,In_140,In_150);
xnor U4529 (N_4529,In_181,In_821);
or U4530 (N_4530,In_405,In_770);
and U4531 (N_4531,In_686,In_820);
nor U4532 (N_4532,In_670,In_599);
nand U4533 (N_4533,In_935,In_563);
or U4534 (N_4534,In_543,In_454);
or U4535 (N_4535,In_147,In_541);
or U4536 (N_4536,In_550,In_84);
xnor U4537 (N_4537,In_239,In_848);
nand U4538 (N_4538,In_565,In_128);
nor U4539 (N_4539,In_704,In_101);
nand U4540 (N_4540,In_826,In_86);
nor U4541 (N_4541,In_165,In_308);
nand U4542 (N_4542,In_99,In_700);
nor U4543 (N_4543,In_306,In_179);
or U4544 (N_4544,In_402,In_937);
nand U4545 (N_4545,In_755,In_609);
nor U4546 (N_4546,In_918,In_89);
nor U4547 (N_4547,In_349,In_452);
and U4548 (N_4548,In_771,In_986);
or U4549 (N_4549,In_341,In_642);
or U4550 (N_4550,In_13,In_379);
and U4551 (N_4551,In_167,In_388);
and U4552 (N_4552,In_479,In_737);
or U4553 (N_4553,In_529,In_286);
nor U4554 (N_4554,In_570,In_13);
and U4555 (N_4555,In_364,In_264);
and U4556 (N_4556,In_70,In_792);
nor U4557 (N_4557,In_509,In_999);
nand U4558 (N_4558,In_525,In_320);
or U4559 (N_4559,In_677,In_804);
or U4560 (N_4560,In_170,In_382);
and U4561 (N_4561,In_993,In_292);
and U4562 (N_4562,In_704,In_108);
or U4563 (N_4563,In_604,In_119);
nand U4564 (N_4564,In_184,In_202);
nor U4565 (N_4565,In_539,In_580);
and U4566 (N_4566,In_147,In_505);
or U4567 (N_4567,In_112,In_150);
nor U4568 (N_4568,In_445,In_177);
and U4569 (N_4569,In_525,In_507);
nand U4570 (N_4570,In_627,In_794);
and U4571 (N_4571,In_967,In_185);
and U4572 (N_4572,In_447,In_544);
and U4573 (N_4573,In_457,In_833);
nand U4574 (N_4574,In_502,In_614);
nor U4575 (N_4575,In_717,In_992);
nor U4576 (N_4576,In_406,In_27);
and U4577 (N_4577,In_101,In_597);
and U4578 (N_4578,In_607,In_570);
nand U4579 (N_4579,In_865,In_520);
nand U4580 (N_4580,In_935,In_91);
or U4581 (N_4581,In_610,In_684);
or U4582 (N_4582,In_317,In_789);
nand U4583 (N_4583,In_638,In_987);
nor U4584 (N_4584,In_555,In_892);
nand U4585 (N_4585,In_437,In_736);
nand U4586 (N_4586,In_386,In_438);
nand U4587 (N_4587,In_188,In_410);
nand U4588 (N_4588,In_170,In_199);
nor U4589 (N_4589,In_219,In_283);
nand U4590 (N_4590,In_623,In_104);
or U4591 (N_4591,In_448,In_696);
nor U4592 (N_4592,In_117,In_925);
and U4593 (N_4593,In_409,In_471);
nor U4594 (N_4594,In_51,In_408);
nand U4595 (N_4595,In_196,In_127);
or U4596 (N_4596,In_189,In_541);
or U4597 (N_4597,In_663,In_926);
nor U4598 (N_4598,In_611,In_468);
nand U4599 (N_4599,In_658,In_980);
nand U4600 (N_4600,In_924,In_182);
xnor U4601 (N_4601,In_590,In_311);
nor U4602 (N_4602,In_677,In_573);
nand U4603 (N_4603,In_63,In_734);
nand U4604 (N_4604,In_354,In_729);
and U4605 (N_4605,In_401,In_950);
nor U4606 (N_4606,In_858,In_880);
nor U4607 (N_4607,In_88,In_900);
or U4608 (N_4608,In_96,In_605);
nor U4609 (N_4609,In_326,In_53);
or U4610 (N_4610,In_474,In_170);
nor U4611 (N_4611,In_848,In_332);
and U4612 (N_4612,In_681,In_488);
and U4613 (N_4613,In_3,In_671);
nor U4614 (N_4614,In_876,In_672);
nand U4615 (N_4615,In_812,In_259);
nand U4616 (N_4616,In_744,In_402);
nor U4617 (N_4617,In_806,In_708);
and U4618 (N_4618,In_694,In_734);
and U4619 (N_4619,In_533,In_835);
nand U4620 (N_4620,In_899,In_925);
and U4621 (N_4621,In_718,In_490);
nand U4622 (N_4622,In_905,In_171);
nand U4623 (N_4623,In_677,In_401);
nand U4624 (N_4624,In_340,In_499);
and U4625 (N_4625,In_14,In_276);
or U4626 (N_4626,In_572,In_745);
nor U4627 (N_4627,In_875,In_183);
and U4628 (N_4628,In_231,In_997);
nor U4629 (N_4629,In_486,In_201);
nor U4630 (N_4630,In_46,In_319);
and U4631 (N_4631,In_675,In_957);
and U4632 (N_4632,In_615,In_977);
nor U4633 (N_4633,In_136,In_849);
or U4634 (N_4634,In_985,In_146);
and U4635 (N_4635,In_69,In_501);
nor U4636 (N_4636,In_201,In_166);
nand U4637 (N_4637,In_907,In_736);
nor U4638 (N_4638,In_931,In_945);
nor U4639 (N_4639,In_863,In_744);
and U4640 (N_4640,In_457,In_219);
nor U4641 (N_4641,In_583,In_110);
nand U4642 (N_4642,In_169,In_434);
and U4643 (N_4643,In_241,In_189);
nor U4644 (N_4644,In_138,In_177);
or U4645 (N_4645,In_195,In_605);
nand U4646 (N_4646,In_765,In_207);
nor U4647 (N_4647,In_302,In_917);
or U4648 (N_4648,In_608,In_700);
and U4649 (N_4649,In_58,In_604);
nand U4650 (N_4650,In_451,In_494);
and U4651 (N_4651,In_769,In_742);
and U4652 (N_4652,In_353,In_770);
xnor U4653 (N_4653,In_313,In_987);
or U4654 (N_4654,In_308,In_521);
nor U4655 (N_4655,In_955,In_351);
nor U4656 (N_4656,In_257,In_842);
xor U4657 (N_4657,In_418,In_230);
nand U4658 (N_4658,In_631,In_304);
nand U4659 (N_4659,In_113,In_685);
nand U4660 (N_4660,In_850,In_857);
and U4661 (N_4661,In_902,In_816);
and U4662 (N_4662,In_754,In_556);
nor U4663 (N_4663,In_752,In_865);
or U4664 (N_4664,In_875,In_814);
nor U4665 (N_4665,In_98,In_27);
or U4666 (N_4666,In_880,In_176);
nand U4667 (N_4667,In_549,In_553);
and U4668 (N_4668,In_467,In_802);
xor U4669 (N_4669,In_407,In_842);
and U4670 (N_4670,In_862,In_268);
and U4671 (N_4671,In_454,In_684);
and U4672 (N_4672,In_320,In_432);
nor U4673 (N_4673,In_808,In_649);
and U4674 (N_4674,In_444,In_864);
and U4675 (N_4675,In_623,In_289);
or U4676 (N_4676,In_540,In_87);
or U4677 (N_4677,In_302,In_761);
nor U4678 (N_4678,In_474,In_834);
and U4679 (N_4679,In_107,In_305);
nand U4680 (N_4680,In_105,In_876);
and U4681 (N_4681,In_848,In_325);
nor U4682 (N_4682,In_931,In_260);
or U4683 (N_4683,In_241,In_578);
and U4684 (N_4684,In_671,In_732);
nand U4685 (N_4685,In_149,In_793);
and U4686 (N_4686,In_331,In_645);
and U4687 (N_4687,In_573,In_85);
and U4688 (N_4688,In_630,In_730);
xnor U4689 (N_4689,In_174,In_393);
nor U4690 (N_4690,In_494,In_313);
nand U4691 (N_4691,In_893,In_242);
nor U4692 (N_4692,In_559,In_994);
nor U4693 (N_4693,In_36,In_795);
or U4694 (N_4694,In_289,In_212);
or U4695 (N_4695,In_272,In_614);
nand U4696 (N_4696,In_980,In_801);
or U4697 (N_4697,In_694,In_576);
nor U4698 (N_4698,In_145,In_543);
nor U4699 (N_4699,In_878,In_489);
and U4700 (N_4700,In_64,In_750);
nand U4701 (N_4701,In_227,In_67);
nand U4702 (N_4702,In_401,In_104);
nand U4703 (N_4703,In_741,In_486);
or U4704 (N_4704,In_756,In_767);
nor U4705 (N_4705,In_296,In_123);
nor U4706 (N_4706,In_151,In_590);
and U4707 (N_4707,In_304,In_960);
or U4708 (N_4708,In_858,In_134);
or U4709 (N_4709,In_836,In_274);
nor U4710 (N_4710,In_670,In_737);
xnor U4711 (N_4711,In_909,In_522);
nor U4712 (N_4712,In_724,In_331);
nor U4713 (N_4713,In_258,In_891);
nand U4714 (N_4714,In_385,In_745);
xor U4715 (N_4715,In_462,In_539);
and U4716 (N_4716,In_848,In_551);
nor U4717 (N_4717,In_410,In_760);
and U4718 (N_4718,In_83,In_367);
nand U4719 (N_4719,In_830,In_870);
nor U4720 (N_4720,In_825,In_983);
nand U4721 (N_4721,In_53,In_552);
nor U4722 (N_4722,In_685,In_546);
and U4723 (N_4723,In_177,In_489);
xnor U4724 (N_4724,In_576,In_25);
nor U4725 (N_4725,In_579,In_913);
or U4726 (N_4726,In_697,In_366);
nor U4727 (N_4727,In_871,In_241);
or U4728 (N_4728,In_964,In_278);
or U4729 (N_4729,In_789,In_218);
and U4730 (N_4730,In_316,In_148);
or U4731 (N_4731,In_454,In_824);
nand U4732 (N_4732,In_84,In_902);
xnor U4733 (N_4733,In_259,In_386);
or U4734 (N_4734,In_94,In_130);
or U4735 (N_4735,In_797,In_820);
or U4736 (N_4736,In_998,In_916);
nor U4737 (N_4737,In_45,In_669);
or U4738 (N_4738,In_684,In_51);
nand U4739 (N_4739,In_432,In_10);
or U4740 (N_4740,In_108,In_612);
or U4741 (N_4741,In_548,In_926);
or U4742 (N_4742,In_812,In_764);
and U4743 (N_4743,In_659,In_571);
nor U4744 (N_4744,In_96,In_364);
nor U4745 (N_4745,In_946,In_3);
nor U4746 (N_4746,In_719,In_230);
nor U4747 (N_4747,In_35,In_269);
or U4748 (N_4748,In_396,In_783);
nand U4749 (N_4749,In_187,In_60);
or U4750 (N_4750,In_566,In_486);
or U4751 (N_4751,In_999,In_900);
nor U4752 (N_4752,In_165,In_877);
or U4753 (N_4753,In_923,In_568);
or U4754 (N_4754,In_302,In_319);
nor U4755 (N_4755,In_401,In_351);
or U4756 (N_4756,In_351,In_770);
nand U4757 (N_4757,In_458,In_302);
or U4758 (N_4758,In_670,In_337);
and U4759 (N_4759,In_94,In_789);
nor U4760 (N_4760,In_448,In_869);
nand U4761 (N_4761,In_848,In_309);
nor U4762 (N_4762,In_867,In_668);
nor U4763 (N_4763,In_560,In_320);
or U4764 (N_4764,In_733,In_31);
nor U4765 (N_4765,In_868,In_304);
nor U4766 (N_4766,In_384,In_506);
or U4767 (N_4767,In_745,In_268);
and U4768 (N_4768,In_736,In_823);
xor U4769 (N_4769,In_69,In_452);
nand U4770 (N_4770,In_757,In_483);
nand U4771 (N_4771,In_993,In_828);
nand U4772 (N_4772,In_597,In_457);
nor U4773 (N_4773,In_166,In_26);
and U4774 (N_4774,In_639,In_407);
nand U4775 (N_4775,In_565,In_691);
nand U4776 (N_4776,In_56,In_324);
nand U4777 (N_4777,In_587,In_205);
xor U4778 (N_4778,In_586,In_464);
or U4779 (N_4779,In_725,In_109);
or U4780 (N_4780,In_554,In_905);
nor U4781 (N_4781,In_200,In_689);
nand U4782 (N_4782,In_585,In_993);
nand U4783 (N_4783,In_770,In_452);
nor U4784 (N_4784,In_839,In_340);
and U4785 (N_4785,In_136,In_60);
or U4786 (N_4786,In_847,In_661);
or U4787 (N_4787,In_920,In_849);
and U4788 (N_4788,In_458,In_650);
nand U4789 (N_4789,In_929,In_812);
nor U4790 (N_4790,In_279,In_434);
and U4791 (N_4791,In_491,In_596);
nand U4792 (N_4792,In_693,In_64);
or U4793 (N_4793,In_815,In_89);
nor U4794 (N_4794,In_352,In_172);
nand U4795 (N_4795,In_717,In_154);
and U4796 (N_4796,In_134,In_394);
nor U4797 (N_4797,In_458,In_433);
or U4798 (N_4798,In_841,In_389);
or U4799 (N_4799,In_464,In_850);
nand U4800 (N_4800,In_66,In_963);
nor U4801 (N_4801,In_715,In_159);
nor U4802 (N_4802,In_965,In_515);
and U4803 (N_4803,In_536,In_228);
and U4804 (N_4804,In_443,In_446);
or U4805 (N_4805,In_984,In_463);
nor U4806 (N_4806,In_788,In_499);
nand U4807 (N_4807,In_806,In_323);
or U4808 (N_4808,In_810,In_584);
and U4809 (N_4809,In_976,In_188);
or U4810 (N_4810,In_16,In_77);
nor U4811 (N_4811,In_277,In_977);
and U4812 (N_4812,In_526,In_25);
or U4813 (N_4813,In_371,In_860);
nor U4814 (N_4814,In_269,In_987);
and U4815 (N_4815,In_136,In_4);
nor U4816 (N_4816,In_51,In_725);
xor U4817 (N_4817,In_651,In_618);
and U4818 (N_4818,In_281,In_963);
nand U4819 (N_4819,In_174,In_170);
and U4820 (N_4820,In_823,In_925);
nor U4821 (N_4821,In_767,In_376);
and U4822 (N_4822,In_0,In_18);
and U4823 (N_4823,In_25,In_615);
nand U4824 (N_4824,In_104,In_847);
nand U4825 (N_4825,In_948,In_660);
nor U4826 (N_4826,In_636,In_221);
and U4827 (N_4827,In_183,In_248);
nand U4828 (N_4828,In_42,In_269);
and U4829 (N_4829,In_408,In_115);
nor U4830 (N_4830,In_551,In_904);
nor U4831 (N_4831,In_187,In_82);
nand U4832 (N_4832,In_271,In_729);
and U4833 (N_4833,In_716,In_37);
and U4834 (N_4834,In_471,In_249);
nor U4835 (N_4835,In_489,In_41);
nand U4836 (N_4836,In_382,In_200);
nand U4837 (N_4837,In_847,In_624);
or U4838 (N_4838,In_329,In_781);
nor U4839 (N_4839,In_986,In_615);
or U4840 (N_4840,In_939,In_705);
nor U4841 (N_4841,In_508,In_192);
nor U4842 (N_4842,In_690,In_898);
nand U4843 (N_4843,In_252,In_273);
nand U4844 (N_4844,In_182,In_933);
or U4845 (N_4845,In_290,In_84);
or U4846 (N_4846,In_956,In_512);
or U4847 (N_4847,In_693,In_494);
nor U4848 (N_4848,In_133,In_889);
or U4849 (N_4849,In_991,In_449);
nand U4850 (N_4850,In_35,In_403);
nand U4851 (N_4851,In_48,In_164);
or U4852 (N_4852,In_655,In_762);
nor U4853 (N_4853,In_19,In_951);
or U4854 (N_4854,In_874,In_745);
and U4855 (N_4855,In_573,In_0);
or U4856 (N_4856,In_827,In_501);
and U4857 (N_4857,In_246,In_92);
or U4858 (N_4858,In_989,In_64);
nor U4859 (N_4859,In_428,In_125);
and U4860 (N_4860,In_747,In_682);
nand U4861 (N_4861,In_681,In_131);
and U4862 (N_4862,In_275,In_876);
and U4863 (N_4863,In_320,In_622);
nor U4864 (N_4864,In_548,In_101);
and U4865 (N_4865,In_561,In_390);
nor U4866 (N_4866,In_782,In_656);
nor U4867 (N_4867,In_422,In_812);
and U4868 (N_4868,In_892,In_497);
nor U4869 (N_4869,In_868,In_313);
nand U4870 (N_4870,In_604,In_202);
nand U4871 (N_4871,In_730,In_128);
nand U4872 (N_4872,In_167,In_653);
and U4873 (N_4873,In_988,In_763);
xor U4874 (N_4874,In_822,In_338);
or U4875 (N_4875,In_900,In_657);
or U4876 (N_4876,In_200,In_950);
nor U4877 (N_4877,In_987,In_655);
nor U4878 (N_4878,In_462,In_956);
or U4879 (N_4879,In_557,In_716);
nand U4880 (N_4880,In_961,In_311);
or U4881 (N_4881,In_269,In_37);
and U4882 (N_4882,In_535,In_468);
or U4883 (N_4883,In_883,In_132);
and U4884 (N_4884,In_508,In_995);
nand U4885 (N_4885,In_860,In_450);
or U4886 (N_4886,In_509,In_815);
nand U4887 (N_4887,In_698,In_325);
and U4888 (N_4888,In_308,In_524);
and U4889 (N_4889,In_231,In_897);
and U4890 (N_4890,In_240,In_456);
nor U4891 (N_4891,In_883,In_244);
nor U4892 (N_4892,In_550,In_953);
nand U4893 (N_4893,In_873,In_71);
nor U4894 (N_4894,In_296,In_355);
and U4895 (N_4895,In_625,In_497);
or U4896 (N_4896,In_153,In_649);
nand U4897 (N_4897,In_624,In_11);
nand U4898 (N_4898,In_865,In_718);
and U4899 (N_4899,In_864,In_766);
nor U4900 (N_4900,In_200,In_941);
nand U4901 (N_4901,In_218,In_751);
nand U4902 (N_4902,In_736,In_279);
or U4903 (N_4903,In_532,In_39);
nor U4904 (N_4904,In_574,In_777);
nand U4905 (N_4905,In_542,In_352);
or U4906 (N_4906,In_12,In_428);
or U4907 (N_4907,In_673,In_341);
and U4908 (N_4908,In_113,In_379);
or U4909 (N_4909,In_101,In_703);
nor U4910 (N_4910,In_336,In_156);
and U4911 (N_4911,In_409,In_335);
nor U4912 (N_4912,In_263,In_990);
nor U4913 (N_4913,In_383,In_114);
and U4914 (N_4914,In_964,In_15);
nor U4915 (N_4915,In_117,In_953);
or U4916 (N_4916,In_939,In_805);
or U4917 (N_4917,In_40,In_450);
or U4918 (N_4918,In_487,In_461);
nor U4919 (N_4919,In_349,In_335);
and U4920 (N_4920,In_108,In_117);
nor U4921 (N_4921,In_609,In_809);
nor U4922 (N_4922,In_893,In_813);
or U4923 (N_4923,In_523,In_33);
or U4924 (N_4924,In_781,In_163);
nor U4925 (N_4925,In_920,In_365);
nand U4926 (N_4926,In_232,In_700);
and U4927 (N_4927,In_711,In_955);
or U4928 (N_4928,In_642,In_832);
and U4929 (N_4929,In_141,In_54);
nor U4930 (N_4930,In_625,In_912);
nand U4931 (N_4931,In_500,In_575);
nor U4932 (N_4932,In_642,In_977);
or U4933 (N_4933,In_323,In_242);
xnor U4934 (N_4934,In_701,In_655);
and U4935 (N_4935,In_650,In_684);
nor U4936 (N_4936,In_596,In_710);
or U4937 (N_4937,In_212,In_860);
nor U4938 (N_4938,In_540,In_373);
nor U4939 (N_4939,In_322,In_484);
xor U4940 (N_4940,In_313,In_275);
or U4941 (N_4941,In_563,In_614);
or U4942 (N_4942,In_160,In_939);
or U4943 (N_4943,In_493,In_174);
nor U4944 (N_4944,In_682,In_40);
nor U4945 (N_4945,In_673,In_921);
or U4946 (N_4946,In_861,In_247);
and U4947 (N_4947,In_601,In_584);
nor U4948 (N_4948,In_936,In_325);
and U4949 (N_4949,In_350,In_911);
and U4950 (N_4950,In_216,In_562);
or U4951 (N_4951,In_918,In_318);
and U4952 (N_4952,In_878,In_218);
and U4953 (N_4953,In_300,In_216);
and U4954 (N_4954,In_909,In_543);
nor U4955 (N_4955,In_47,In_471);
or U4956 (N_4956,In_905,In_206);
nor U4957 (N_4957,In_837,In_961);
nor U4958 (N_4958,In_948,In_782);
and U4959 (N_4959,In_730,In_8);
nor U4960 (N_4960,In_781,In_749);
nand U4961 (N_4961,In_85,In_648);
nand U4962 (N_4962,In_884,In_69);
nand U4963 (N_4963,In_434,In_580);
or U4964 (N_4964,In_124,In_412);
and U4965 (N_4965,In_93,In_656);
nand U4966 (N_4966,In_754,In_69);
nand U4967 (N_4967,In_977,In_881);
nand U4968 (N_4968,In_57,In_466);
nand U4969 (N_4969,In_600,In_560);
nor U4970 (N_4970,In_892,In_666);
nand U4971 (N_4971,In_752,In_352);
and U4972 (N_4972,In_200,In_852);
nand U4973 (N_4973,In_947,In_967);
or U4974 (N_4974,In_679,In_167);
nand U4975 (N_4975,In_392,In_973);
nor U4976 (N_4976,In_729,In_187);
nand U4977 (N_4977,In_299,In_8);
nor U4978 (N_4978,In_534,In_547);
xor U4979 (N_4979,In_210,In_466);
nor U4980 (N_4980,In_402,In_97);
nor U4981 (N_4981,In_42,In_641);
nand U4982 (N_4982,In_573,In_438);
nor U4983 (N_4983,In_866,In_488);
and U4984 (N_4984,In_482,In_951);
nand U4985 (N_4985,In_956,In_551);
or U4986 (N_4986,In_967,In_177);
nand U4987 (N_4987,In_239,In_521);
or U4988 (N_4988,In_405,In_899);
nor U4989 (N_4989,In_989,In_483);
and U4990 (N_4990,In_41,In_613);
nand U4991 (N_4991,In_455,In_935);
and U4992 (N_4992,In_547,In_919);
nor U4993 (N_4993,In_673,In_18);
or U4994 (N_4994,In_483,In_778);
nor U4995 (N_4995,In_261,In_966);
nand U4996 (N_4996,In_637,In_217);
and U4997 (N_4997,In_574,In_613);
and U4998 (N_4998,In_126,In_851);
and U4999 (N_4999,In_583,In_737);
and U5000 (N_5000,N_670,N_440);
nand U5001 (N_5001,N_861,N_4864);
nand U5002 (N_5002,N_1386,N_525);
nand U5003 (N_5003,N_842,N_608);
xor U5004 (N_5004,N_1573,N_1029);
nor U5005 (N_5005,N_2359,N_4227);
or U5006 (N_5006,N_3421,N_4940);
nor U5007 (N_5007,N_1815,N_2570);
and U5008 (N_5008,N_1022,N_3127);
nor U5009 (N_5009,N_4011,N_3411);
nand U5010 (N_5010,N_2583,N_4030);
nand U5011 (N_5011,N_3743,N_4352);
or U5012 (N_5012,N_961,N_3613);
and U5013 (N_5013,N_3279,N_1725);
nand U5014 (N_5014,N_1073,N_3822);
nand U5015 (N_5015,N_2466,N_2900);
or U5016 (N_5016,N_4466,N_323);
nand U5017 (N_5017,N_2920,N_2602);
nand U5018 (N_5018,N_1647,N_1788);
nand U5019 (N_5019,N_3886,N_3044);
and U5020 (N_5020,N_4076,N_1496);
nand U5021 (N_5021,N_420,N_4526);
nand U5022 (N_5022,N_4586,N_4226);
or U5023 (N_5023,N_3794,N_3269);
and U5024 (N_5024,N_2671,N_1095);
and U5025 (N_5025,N_3379,N_522);
or U5026 (N_5026,N_773,N_2899);
and U5027 (N_5027,N_343,N_4023);
nand U5028 (N_5028,N_3109,N_455);
and U5029 (N_5029,N_689,N_878);
or U5030 (N_5030,N_602,N_2950);
nor U5031 (N_5031,N_3071,N_1538);
or U5032 (N_5032,N_3740,N_3157);
and U5033 (N_5033,N_4900,N_1049);
xor U5034 (N_5034,N_726,N_3492);
or U5035 (N_5035,N_1949,N_4158);
xor U5036 (N_5036,N_2263,N_845);
nand U5037 (N_5037,N_3659,N_2474);
nor U5038 (N_5038,N_4349,N_3891);
and U5039 (N_5039,N_180,N_4284);
xor U5040 (N_5040,N_460,N_4052);
and U5041 (N_5041,N_2635,N_1075);
and U5042 (N_5042,N_4140,N_1714);
nand U5043 (N_5043,N_4827,N_792);
nor U5044 (N_5044,N_4620,N_2180);
nand U5045 (N_5045,N_874,N_2021);
nor U5046 (N_5046,N_4272,N_3208);
or U5047 (N_5047,N_2267,N_4340);
or U5048 (N_5048,N_644,N_294);
and U5049 (N_5049,N_3679,N_2731);
and U5050 (N_5050,N_4175,N_3329);
nor U5051 (N_5051,N_4631,N_4582);
nor U5052 (N_5052,N_2047,N_4339);
and U5053 (N_5053,N_1456,N_2553);
xnor U5054 (N_5054,N_950,N_4539);
or U5055 (N_5055,N_4596,N_3398);
or U5056 (N_5056,N_4671,N_3161);
or U5057 (N_5057,N_1971,N_2578);
nor U5058 (N_5058,N_2092,N_938);
nor U5059 (N_5059,N_1378,N_2242);
nor U5060 (N_5060,N_4004,N_2998);
xor U5061 (N_5061,N_554,N_2879);
and U5062 (N_5062,N_4040,N_3002);
nor U5063 (N_5063,N_779,N_733);
nor U5064 (N_5064,N_926,N_905);
nor U5065 (N_5065,N_4522,N_2455);
or U5066 (N_5066,N_1369,N_4492);
and U5067 (N_5067,N_4960,N_669);
nor U5068 (N_5068,N_4171,N_3923);
or U5069 (N_5069,N_251,N_506);
and U5070 (N_5070,N_645,N_2364);
or U5071 (N_5071,N_3505,N_3133);
or U5072 (N_5072,N_1899,N_434);
nand U5073 (N_5073,N_4774,N_1636);
nor U5074 (N_5074,N_3456,N_2017);
and U5075 (N_5075,N_2418,N_3339);
nand U5076 (N_5076,N_379,N_916);
nor U5077 (N_5077,N_383,N_1986);
and U5078 (N_5078,N_3995,N_3872);
xnor U5079 (N_5079,N_83,N_4648);
nor U5080 (N_5080,N_1206,N_1021);
nor U5081 (N_5081,N_4686,N_2307);
and U5082 (N_5082,N_632,N_2807);
nand U5083 (N_5083,N_781,N_204);
nand U5084 (N_5084,N_841,N_3299);
or U5085 (N_5085,N_3388,N_4353);
nand U5086 (N_5086,N_4371,N_4881);
or U5087 (N_5087,N_4921,N_3930);
and U5088 (N_5088,N_1025,N_2110);
nor U5089 (N_5089,N_1295,N_1625);
and U5090 (N_5090,N_247,N_4232);
or U5091 (N_5091,N_3196,N_1287);
nor U5092 (N_5092,N_4738,N_4326);
or U5093 (N_5093,N_529,N_3014);
or U5094 (N_5094,N_576,N_807);
nor U5095 (N_5095,N_1885,N_2736);
xnor U5096 (N_5096,N_413,N_4788);
nor U5097 (N_5097,N_3833,N_4649);
or U5098 (N_5098,N_1972,N_1964);
nand U5099 (N_5099,N_226,N_2618);
nor U5100 (N_5100,N_1474,N_4816);
nand U5101 (N_5101,N_557,N_93);
or U5102 (N_5102,N_4278,N_1979);
nand U5103 (N_5103,N_3934,N_3455);
or U5104 (N_5104,N_2986,N_3340);
xor U5105 (N_5105,N_2095,N_3675);
and U5106 (N_5106,N_109,N_4263);
or U5107 (N_5107,N_3371,N_604);
nand U5108 (N_5108,N_2321,N_1070);
and U5109 (N_5109,N_2526,N_3596);
and U5110 (N_5110,N_2171,N_4305);
nor U5111 (N_5111,N_3181,N_1341);
nand U5112 (N_5112,N_1896,N_2908);
nor U5113 (N_5113,N_1939,N_3314);
or U5114 (N_5114,N_268,N_1605);
nand U5115 (N_5115,N_550,N_1257);
and U5116 (N_5116,N_1463,N_955);
nor U5117 (N_5117,N_3972,N_1064);
and U5118 (N_5118,N_1806,N_3107);
nor U5119 (N_5119,N_1084,N_2015);
and U5120 (N_5120,N_4018,N_1786);
or U5121 (N_5121,N_1513,N_1054);
xor U5122 (N_5122,N_4786,N_1012);
nand U5123 (N_5123,N_4715,N_2211);
xor U5124 (N_5124,N_1439,N_1619);
and U5125 (N_5125,N_3331,N_1348);
nand U5126 (N_5126,N_1805,N_3801);
xor U5127 (N_5127,N_2724,N_3300);
or U5128 (N_5128,N_3650,N_4877);
or U5129 (N_5129,N_1111,N_1442);
nand U5130 (N_5130,N_4022,N_3311);
nor U5131 (N_5131,N_3984,N_3325);
nor U5132 (N_5132,N_873,N_4693);
nor U5133 (N_5133,N_3457,N_940);
and U5134 (N_5134,N_1580,N_2616);
or U5135 (N_5135,N_3427,N_3548);
nor U5136 (N_5136,N_556,N_130);
or U5137 (N_5137,N_3174,N_4830);
and U5138 (N_5138,N_4945,N_1934);
and U5139 (N_5139,N_2245,N_3106);
or U5140 (N_5140,N_4682,N_3194);
or U5141 (N_5141,N_4652,N_2980);
nand U5142 (N_5142,N_2140,N_794);
nand U5143 (N_5143,N_4447,N_2801);
nand U5144 (N_5144,N_692,N_3045);
nand U5145 (N_5145,N_2363,N_2974);
nor U5146 (N_5146,N_2719,N_2195);
nor U5147 (N_5147,N_4880,N_1825);
or U5148 (N_5148,N_3628,N_4432);
xor U5149 (N_5149,N_3423,N_3054);
or U5150 (N_5150,N_680,N_2342);
nand U5151 (N_5151,N_1796,N_1418);
or U5152 (N_5152,N_3125,N_3495);
xnor U5153 (N_5153,N_4510,N_2210);
nand U5154 (N_5154,N_2790,N_3330);
or U5155 (N_5155,N_1326,N_1682);
xnor U5156 (N_5156,N_891,N_3324);
nand U5157 (N_5157,N_1950,N_3232);
nand U5158 (N_5158,N_3584,N_4903);
and U5159 (N_5159,N_2942,N_1485);
and U5160 (N_5160,N_1723,N_577);
and U5161 (N_5161,N_4930,N_4707);
or U5162 (N_5162,N_2885,N_969);
or U5163 (N_5163,N_4251,N_3531);
and U5164 (N_5164,N_3023,N_4219);
nand U5165 (N_5165,N_3342,N_2068);
nor U5166 (N_5166,N_2415,N_2820);
nand U5167 (N_5167,N_4071,N_2361);
nand U5168 (N_5168,N_1650,N_2038);
nand U5169 (N_5169,N_3394,N_4116);
or U5170 (N_5170,N_988,N_2381);
and U5171 (N_5171,N_472,N_3674);
xor U5172 (N_5172,N_3895,N_1771);
nand U5173 (N_5173,N_1931,N_1334);
nand U5174 (N_5174,N_1288,N_380);
nand U5175 (N_5175,N_1171,N_1921);
and U5176 (N_5176,N_3908,N_2059);
nor U5177 (N_5177,N_3770,N_2251);
nand U5178 (N_5178,N_3224,N_3449);
nor U5179 (N_5179,N_4836,N_759);
and U5180 (N_5180,N_1976,N_1307);
and U5181 (N_5181,N_1905,N_4568);
nor U5182 (N_5182,N_4919,N_3926);
and U5183 (N_5183,N_519,N_1944);
and U5184 (N_5184,N_2535,N_3665);
or U5185 (N_5185,N_3301,N_3074);
and U5186 (N_5186,N_3825,N_4828);
or U5187 (N_5187,N_1562,N_889);
nand U5188 (N_5188,N_4292,N_3386);
and U5189 (N_5189,N_3927,N_2883);
and U5190 (N_5190,N_2521,N_4107);
nor U5191 (N_5191,N_1205,N_4750);
nor U5192 (N_5192,N_4080,N_672);
or U5193 (N_5193,N_1933,N_1669);
or U5194 (N_5194,N_3618,N_1457);
nand U5195 (N_5195,N_886,N_4431);
nand U5196 (N_5196,N_4405,N_30);
nor U5197 (N_5197,N_4096,N_720);
or U5198 (N_5198,N_2437,N_4275);
nor U5199 (N_5199,N_360,N_4119);
nor U5200 (N_5200,N_4527,N_4303);
or U5201 (N_5201,N_3088,N_3429);
nand U5202 (N_5202,N_2413,N_666);
nor U5203 (N_5203,N_403,N_3861);
and U5204 (N_5204,N_4013,N_1429);
nand U5205 (N_5205,N_1795,N_4240);
nand U5206 (N_5206,N_2964,N_4056);
nand U5207 (N_5207,N_4058,N_444);
xor U5208 (N_5208,N_1594,N_3186);
or U5209 (N_5209,N_1421,N_162);
nor U5210 (N_5210,N_816,N_3152);
or U5211 (N_5211,N_1768,N_1278);
or U5212 (N_5212,N_3462,N_2912);
nand U5213 (N_5213,N_4411,N_755);
or U5214 (N_5214,N_2104,N_637);
and U5215 (N_5215,N_1048,N_3624);
nand U5216 (N_5216,N_2617,N_2734);
nand U5217 (N_5217,N_4289,N_2254);
or U5218 (N_5218,N_1104,N_4815);
and U5219 (N_5219,N_3222,N_482);
or U5220 (N_5220,N_1291,N_2276);
nor U5221 (N_5221,N_3017,N_863);
nand U5222 (N_5222,N_4656,N_744);
nand U5223 (N_5223,N_1058,N_948);
or U5224 (N_5224,N_2491,N_4832);
and U5225 (N_5225,N_3263,N_1602);
nor U5226 (N_5226,N_3562,N_1557);
nor U5227 (N_5227,N_4533,N_2056);
nor U5228 (N_5228,N_4768,N_2769);
nand U5229 (N_5229,N_2141,N_2405);
nor U5230 (N_5230,N_4100,N_171);
and U5231 (N_5231,N_4986,N_77);
and U5232 (N_5232,N_4714,N_2718);
nor U5233 (N_5233,N_2226,N_3787);
and U5234 (N_5234,N_4325,N_4237);
or U5235 (N_5235,N_2377,N_1253);
and U5236 (N_5236,N_4350,N_804);
nand U5237 (N_5237,N_3571,N_2194);
nor U5238 (N_5238,N_2914,N_376);
nand U5239 (N_5239,N_797,N_1910);
nor U5240 (N_5240,N_933,N_502);
xnor U5241 (N_5241,N_15,N_2090);
nor U5242 (N_5242,N_4535,N_3996);
and U5243 (N_5243,N_3922,N_1583);
and U5244 (N_5244,N_4366,N_4760);
or U5245 (N_5245,N_4034,N_711);
nor U5246 (N_5246,N_1843,N_815);
and U5247 (N_5247,N_4271,N_2128);
nand U5248 (N_5248,N_3589,N_4488);
xnor U5249 (N_5249,N_1898,N_2153);
and U5250 (N_5250,N_2600,N_593);
or U5251 (N_5251,N_1087,N_1559);
and U5252 (N_5252,N_2743,N_4451);
or U5253 (N_5253,N_1269,N_3382);
or U5254 (N_5254,N_4994,N_2449);
nand U5255 (N_5255,N_4127,N_2637);
and U5256 (N_5256,N_4010,N_1614);
and U5257 (N_5257,N_501,N_2096);
nor U5258 (N_5258,N_2881,N_4295);
or U5259 (N_5259,N_2597,N_2776);
and U5260 (N_5260,N_600,N_4988);
or U5261 (N_5261,N_1545,N_337);
nor U5262 (N_5262,N_2246,N_698);
or U5263 (N_5263,N_3982,N_2833);
nor U5264 (N_5264,N_3018,N_3254);
nand U5265 (N_5265,N_1314,N_3215);
nand U5266 (N_5266,N_1027,N_47);
and U5267 (N_5267,N_989,N_784);
and U5268 (N_5268,N_3315,N_4701);
and U5269 (N_5269,N_4798,N_4770);
nand U5270 (N_5270,N_316,N_2465);
or U5271 (N_5271,N_1592,N_503);
and U5272 (N_5272,N_2329,N_617);
nor U5273 (N_5273,N_2990,N_1229);
nor U5274 (N_5274,N_4509,N_4708);
and U5275 (N_5275,N_3491,N_433);
nand U5276 (N_5276,N_124,N_4874);
nor U5277 (N_5277,N_230,N_536);
nor U5278 (N_5278,N_3910,N_900);
and U5279 (N_5279,N_4905,N_1435);
or U5280 (N_5280,N_2030,N_3737);
or U5281 (N_5281,N_2199,N_3508);
or U5282 (N_5282,N_2518,N_1623);
nand U5283 (N_5283,N_1320,N_4440);
nand U5284 (N_5284,N_2621,N_1081);
nor U5285 (N_5285,N_3425,N_320);
nand U5286 (N_5286,N_4646,N_4664);
and U5287 (N_5287,N_2882,N_2829);
nor U5288 (N_5288,N_1517,N_936);
nand U5289 (N_5289,N_2072,N_3065);
and U5290 (N_5290,N_3566,N_4429);
nor U5291 (N_5291,N_613,N_4500);
and U5292 (N_5292,N_3093,N_2784);
and U5293 (N_5293,N_2164,N_3707);
nand U5294 (N_5294,N_88,N_1544);
or U5295 (N_5295,N_1695,N_350);
and U5296 (N_5296,N_4070,N_586);
nor U5297 (N_5297,N_1710,N_963);
nor U5298 (N_5298,N_3079,N_2483);
and U5299 (N_5299,N_172,N_4977);
nor U5300 (N_5300,N_627,N_3755);
nor U5301 (N_5301,N_3063,N_1493);
nand U5302 (N_5302,N_1373,N_4476);
nand U5303 (N_5303,N_763,N_1415);
xnor U5304 (N_5304,N_2277,N_4655);
or U5305 (N_5305,N_1036,N_872);
nor U5306 (N_5306,N_546,N_647);
and U5307 (N_5307,N_1826,N_3086);
nand U5308 (N_5308,N_2304,N_817);
nand U5309 (N_5309,N_4464,N_147);
nand U5310 (N_5310,N_3209,N_859);
nor U5311 (N_5311,N_4389,N_3916);
or U5312 (N_5312,N_1394,N_4525);
nor U5313 (N_5313,N_2855,N_1915);
and U5314 (N_5314,N_3575,N_4658);
or U5315 (N_5315,N_1762,N_1280);
or U5316 (N_5316,N_3460,N_377);
nor U5317 (N_5317,N_354,N_2634);
nand U5318 (N_5318,N_3585,N_4966);
or U5319 (N_5319,N_2065,N_3332);
or U5320 (N_5320,N_2149,N_351);
nor U5321 (N_5321,N_3645,N_4223);
or U5322 (N_5322,N_2120,N_1683);
nor U5323 (N_5323,N_3070,N_3742);
nand U5324 (N_5324,N_2118,N_2275);
or U5325 (N_5325,N_1338,N_2752);
nand U5326 (N_5326,N_651,N_1362);
nand U5327 (N_5327,N_611,N_4101);
nand U5328 (N_5328,N_1000,N_6);
and U5329 (N_5329,N_599,N_3990);
nand U5330 (N_5330,N_3101,N_4700);
nand U5331 (N_5331,N_4797,N_1638);
and U5332 (N_5332,N_696,N_4743);
and U5333 (N_5333,N_3466,N_4911);
and U5334 (N_5334,N_777,N_363);
nand U5335 (N_5335,N_995,N_4357);
or U5336 (N_5336,N_4494,N_1574);
nand U5337 (N_5337,N_4270,N_879);
nand U5338 (N_5338,N_2334,N_4996);
and U5339 (N_5339,N_3954,N_4266);
and U5340 (N_5340,N_2709,N_4072);
or U5341 (N_5341,N_1207,N_4122);
or U5342 (N_5342,N_1134,N_3780);
and U5343 (N_5343,N_236,N_2442);
and U5344 (N_5344,N_4862,N_753);
nand U5345 (N_5345,N_2571,N_4785);
or U5346 (N_5346,N_1617,N_3234);
and U5347 (N_5347,N_424,N_4194);
nor U5348 (N_5348,N_3971,N_1407);
nand U5349 (N_5349,N_4471,N_3574);
nor U5350 (N_5350,N_4917,N_2003);
nor U5351 (N_5351,N_76,N_3616);
and U5352 (N_5352,N_2421,N_2667);
and U5353 (N_5353,N_3733,N_3876);
and U5354 (N_5354,N_1697,N_4987);
or U5355 (N_5355,N_2266,N_2259);
nor U5356 (N_5356,N_2704,N_1286);
and U5357 (N_5357,N_4989,N_523);
nor U5358 (N_5358,N_3087,N_4078);
nor U5359 (N_5359,N_4360,N_3376);
and U5360 (N_5360,N_3956,N_2992);
nor U5361 (N_5361,N_3431,N_3728);
nor U5362 (N_5362,N_4433,N_4048);
nor U5363 (N_5363,N_2702,N_1561);
and U5364 (N_5364,N_619,N_237);
nand U5365 (N_5365,N_2086,N_1423);
nand U5366 (N_5366,N_1046,N_3128);
or U5367 (N_5367,N_4687,N_2726);
xor U5368 (N_5368,N_3994,N_2604);
and U5369 (N_5369,N_2585,N_9);
nand U5370 (N_5370,N_210,N_3841);
or U5371 (N_5371,N_4291,N_2649);
nand U5372 (N_5372,N_4578,N_2411);
xor U5373 (N_5373,N_2087,N_3179);
or U5374 (N_5374,N_4667,N_2335);
and U5375 (N_5375,N_4944,N_3461);
and U5376 (N_5376,N_4810,N_2630);
and U5377 (N_5377,N_1310,N_2219);
nand U5378 (N_5378,N_1700,N_3626);
or U5379 (N_5379,N_1651,N_2803);
or U5380 (N_5380,N_998,N_2520);
nand U5381 (N_5381,N_4739,N_2642);
nor U5382 (N_5382,N_2579,N_3621);
nor U5383 (N_5383,N_2052,N_3005);
nand U5384 (N_5384,N_3166,N_3677);
nand U5385 (N_5385,N_2260,N_3920);
and U5386 (N_5386,N_1686,N_3625);
or U5387 (N_5387,N_3808,N_3030);
nor U5388 (N_5388,N_877,N_4901);
nand U5389 (N_5389,N_4089,N_3448);
and U5390 (N_5390,N_1879,N_400);
nand U5391 (N_5391,N_2429,N_397);
nand U5392 (N_5392,N_1904,N_305);
xnor U5393 (N_5393,N_3700,N_3802);
nand U5394 (N_5394,N_4221,N_1735);
and U5395 (N_5395,N_394,N_402);
nor U5396 (N_5396,N_156,N_3655);
nor U5397 (N_5397,N_3167,N_4534);
nor U5398 (N_5398,N_3043,N_3577);
or U5399 (N_5399,N_1005,N_4245);
nor U5400 (N_5400,N_921,N_1869);
nand U5401 (N_5401,N_2979,N_762);
xor U5402 (N_5402,N_2692,N_2447);
nor U5403 (N_5403,N_791,N_612);
or U5404 (N_5404,N_4675,N_2176);
nor U5405 (N_5405,N_55,N_2683);
xor U5406 (N_5406,N_685,N_2515);
and U5407 (N_5407,N_1398,N_463);
xor U5408 (N_5408,N_111,N_3893);
nand U5409 (N_5409,N_2395,N_1542);
and U5410 (N_5410,N_1586,N_2101);
or U5411 (N_5411,N_2108,N_947);
or U5412 (N_5412,N_1279,N_4281);
nand U5413 (N_5413,N_2775,N_2541);
or U5414 (N_5414,N_4430,N_4602);
nor U5415 (N_5415,N_2143,N_1756);
nand U5416 (N_5416,N_946,N_4422);
nor U5417 (N_5417,N_4393,N_2410);
nand U5418 (N_5418,N_1618,N_29);
nand U5419 (N_5419,N_3986,N_3229);
and U5420 (N_5420,N_3378,N_3593);
or U5421 (N_5421,N_1590,N_1648);
nand U5422 (N_5422,N_119,N_4133);
and U5423 (N_5423,N_3878,N_184);
and U5424 (N_5424,N_1096,N_3527);
nor U5425 (N_5425,N_2419,N_1951);
nor U5426 (N_5426,N_2984,N_3695);
or U5427 (N_5427,N_3006,N_925);
and U5428 (N_5428,N_4834,N_509);
nand U5429 (N_5429,N_303,N_4141);
or U5430 (N_5430,N_984,N_2737);
nor U5431 (N_5431,N_2448,N_4933);
xnor U5432 (N_5432,N_1681,N_4699);
nand U5433 (N_5433,N_823,N_2186);
or U5434 (N_5434,N_1876,N_4028);
nor U5435 (N_5435,N_2102,N_3525);
nand U5436 (N_5436,N_721,N_4290);
and U5437 (N_5437,N_2590,N_134);
nand U5438 (N_5438,N_709,N_3009);
and U5439 (N_5439,N_3284,N_3957);
nor U5440 (N_5440,N_3355,N_4593);
or U5441 (N_5441,N_3955,N_2050);
and U5442 (N_5442,N_235,N_1006);
or U5443 (N_5443,N_741,N_3744);
and U5444 (N_5444,N_2244,N_4676);
nor U5445 (N_5445,N_2297,N_1906);
and U5446 (N_5446,N_396,N_3680);
and U5447 (N_5447,N_3966,N_4479);
or U5448 (N_5448,N_1220,N_2404);
and U5449 (N_5449,N_332,N_1626);
and U5450 (N_5450,N_2556,N_3228);
nand U5451 (N_5451,N_2063,N_567);
nand U5452 (N_5452,N_1168,N_3931);
nand U5453 (N_5453,N_1114,N_48);
xor U5454 (N_5454,N_2177,N_73);
nor U5455 (N_5455,N_2677,N_788);
nand U5456 (N_5456,N_4484,N_157);
and U5457 (N_5457,N_1615,N_228);
xor U5458 (N_5458,N_4206,N_100);
nand U5459 (N_5459,N_530,N_1852);
and U5460 (N_5460,N_1100,N_642);
and U5461 (N_5461,N_1039,N_258);
or U5462 (N_5462,N_2866,N_826);
and U5463 (N_5463,N_1599,N_2945);
or U5464 (N_5464,N_1881,N_2033);
nand U5465 (N_5465,N_1042,N_50);
nor U5466 (N_5466,N_1913,N_3310);
nor U5467 (N_5467,N_2686,N_2774);
or U5468 (N_5468,N_581,N_3795);
or U5469 (N_5469,N_2581,N_1502);
nor U5470 (N_5470,N_4347,N_2392);
and U5471 (N_5471,N_2792,N_1841);
and U5472 (N_5472,N_3641,N_866);
nor U5473 (N_5473,N_3843,N_3558);
or U5474 (N_5474,N_1477,N_3012);
or U5475 (N_5475,N_1312,N_2968);
and U5476 (N_5476,N_3413,N_4553);
or U5477 (N_5477,N_3520,N_1044);
xnor U5478 (N_5478,N_3271,N_3555);
nor U5479 (N_5479,N_1136,N_1322);
and U5480 (N_5480,N_618,N_699);
or U5481 (N_5481,N_467,N_959);
nor U5482 (N_5482,N_148,N_3983);
nor U5483 (N_5483,N_1736,N_2427);
xnor U5484 (N_5484,N_1764,N_1577);
or U5485 (N_5485,N_3809,N_385);
nor U5486 (N_5486,N_390,N_2158);
nand U5487 (N_5487,N_3711,N_795);
or U5488 (N_5488,N_1313,N_4195);
or U5489 (N_5489,N_1309,N_2548);
or U5490 (N_5490,N_4095,N_2640);
nor U5491 (N_5491,N_3467,N_1713);
and U5492 (N_5492,N_3115,N_1185);
and U5493 (N_5493,N_2779,N_2391);
nor U5494 (N_5494,N_4514,N_956);
nor U5495 (N_5495,N_3536,N_2196);
nor U5496 (N_5496,N_2814,N_3225);
or U5497 (N_5497,N_4261,N_2894);
or U5498 (N_5498,N_4801,N_1347);
nand U5499 (N_5499,N_952,N_628);
and U5500 (N_5500,N_117,N_4752);
nor U5501 (N_5501,N_1807,N_1704);
and U5502 (N_5502,N_799,N_2229);
xnor U5503 (N_5503,N_479,N_4617);
and U5504 (N_5504,N_3220,N_4265);
nor U5505 (N_5505,N_819,N_2388);
and U5506 (N_5506,N_287,N_1056);
or U5507 (N_5507,N_4971,N_4294);
nand U5508 (N_5508,N_2408,N_4477);
xor U5509 (N_5509,N_4401,N_3257);
nand U5510 (N_5510,N_3410,N_4870);
and U5511 (N_5511,N_3673,N_41);
nor U5512 (N_5512,N_408,N_1645);
or U5513 (N_5513,N_3162,N_471);
or U5514 (N_5514,N_3104,N_2438);
nand U5515 (N_5515,N_2288,N_4322);
nand U5516 (N_5516,N_2167,N_1450);
nand U5517 (N_5517,N_3451,N_2362);
or U5518 (N_5518,N_2272,N_2664);
or U5519 (N_5519,N_478,N_2511);
nor U5520 (N_5520,N_2477,N_4659);
nor U5521 (N_5521,N_2155,N_3717);
and U5522 (N_5522,N_4599,N_2893);
and U5523 (N_5523,N_3281,N_4633);
and U5524 (N_5524,N_1147,N_3476);
and U5525 (N_5525,N_4210,N_1196);
nand U5526 (N_5526,N_4624,N_658);
nand U5527 (N_5527,N_3977,N_1148);
nand U5528 (N_5528,N_1678,N_3146);
and U5529 (N_5529,N_2016,N_4073);
or U5530 (N_5530,N_1115,N_4865);
nand U5531 (N_5531,N_4097,N_200);
and U5532 (N_5532,N_3050,N_4638);
nor U5533 (N_5533,N_3374,N_4812);
or U5534 (N_5534,N_962,N_1302);
nor U5535 (N_5535,N_2930,N_4254);
nor U5536 (N_5536,N_1032,N_2647);
nand U5537 (N_5537,N_3535,N_114);
or U5538 (N_5538,N_1685,N_1726);
nand U5539 (N_5539,N_1020,N_3860);
and U5540 (N_5540,N_3218,N_3151);
nand U5541 (N_5541,N_549,N_2076);
or U5542 (N_5542,N_2516,N_2591);
and U5543 (N_5543,N_1998,N_803);
nor U5544 (N_5544,N_3275,N_1866);
or U5545 (N_5545,N_1716,N_1449);
and U5546 (N_5546,N_897,N_4528);
nand U5547 (N_5547,N_3119,N_4092);
nor U5548 (N_5548,N_4630,N_1729);
nand U5549 (N_5549,N_1299,N_4626);
nor U5550 (N_5550,N_3580,N_3392);
or U5551 (N_5551,N_4588,N_2049);
nor U5552 (N_5552,N_4601,N_4531);
and U5553 (N_5553,N_1479,N_3885);
and U5554 (N_5554,N_90,N_4168);
and U5555 (N_5555,N_578,N_4969);
nor U5556 (N_5556,N_2707,N_3671);
nand U5557 (N_5557,N_1067,N_227);
xor U5558 (N_5558,N_1470,N_1422);
nand U5559 (N_5559,N_1874,N_4420);
nor U5560 (N_5560,N_2946,N_2653);
and U5561 (N_5561,N_4981,N_2542);
nor U5562 (N_5562,N_107,N_1606);
xor U5563 (N_5563,N_3259,N_4167);
and U5564 (N_5564,N_589,N_4385);
and U5565 (N_5565,N_284,N_631);
or U5566 (N_5566,N_4821,N_3796);
nand U5567 (N_5567,N_1186,N_2223);
or U5568 (N_5568,N_1521,N_2973);
nor U5569 (N_5569,N_1294,N_520);
and U5570 (N_5570,N_89,N_518);
or U5571 (N_5571,N_3136,N_673);
and U5572 (N_5572,N_2215,N_4651);
and U5573 (N_5573,N_3066,N_223);
nand U5574 (N_5574,N_1177,N_4787);
or U5575 (N_5575,N_4691,N_1433);
or U5576 (N_5576,N_583,N_4591);
or U5577 (N_5577,N_2057,N_3918);
nand U5578 (N_5578,N_653,N_3091);
nand U5579 (N_5579,N_2549,N_1978);
nor U5580 (N_5580,N_4382,N_2357);
nor U5581 (N_5581,N_3176,N_212);
xor U5582 (N_5582,N_1935,N_1652);
nand U5583 (N_5583,N_2636,N_2374);
nor U5584 (N_5584,N_2145,N_3295);
nand U5585 (N_5585,N_4991,N_3480);
or U5586 (N_5586,N_1842,N_3458);
nand U5587 (N_5587,N_4543,N_3612);
nand U5588 (N_5588,N_3243,N_3682);
and U5589 (N_5589,N_4328,N_667);
or U5590 (N_5590,N_3945,N_1245);
nand U5591 (N_5591,N_2875,N_2133);
or U5592 (N_5592,N_2943,N_2432);
nand U5593 (N_5593,N_2903,N_2770);
nand U5594 (N_5594,N_2778,N_2848);
nor U5595 (N_5595,N_2838,N_362);
or U5596 (N_5596,N_1535,N_2661);
nor U5597 (N_5597,N_1878,N_431);
nor U5598 (N_5598,N_972,N_361);
nand U5599 (N_5599,N_3816,N_2963);
nor U5600 (N_5600,N_2358,N_1043);
or U5601 (N_5601,N_1687,N_1350);
and U5602 (N_5602,N_3953,N_3375);
nor U5603 (N_5603,N_417,N_1443);
and U5604 (N_5604,N_2918,N_2231);
or U5605 (N_5605,N_661,N_4419);
or U5606 (N_5606,N_4443,N_4457);
and U5607 (N_5607,N_2996,N_1717);
or U5608 (N_5608,N_4825,N_4508);
nand U5609 (N_5609,N_2496,N_3697);
or U5610 (N_5610,N_4852,N_2338);
or U5611 (N_5611,N_217,N_1159);
or U5612 (N_5612,N_1598,N_3960);
nor U5613 (N_5613,N_4005,N_603);
nand U5614 (N_5614,N_3468,N_4009);
and U5615 (N_5615,N_3766,N_775);
and U5616 (N_5616,N_3373,N_4939);
or U5617 (N_5617,N_3871,N_2070);
nand U5618 (N_5618,N_4321,N_4502);
nand U5619 (N_5619,N_286,N_3190);
or U5620 (N_5620,N_1514,N_1529);
and U5621 (N_5621,N_918,N_3142);
and U5622 (N_5622,N_4470,N_2004);
and U5623 (N_5623,N_4958,N_3020);
and U5624 (N_5624,N_1706,N_1352);
nand U5625 (N_5625,N_4125,N_2507);
nand U5626 (N_5626,N_4678,N_369);
or U5627 (N_5627,N_307,N_1211);
or U5628 (N_5628,N_4657,N_1116);
or U5629 (N_5629,N_4400,N_2048);
or U5630 (N_5630,N_1737,N_4085);
nand U5631 (N_5631,N_322,N_1464);
and U5632 (N_5632,N_4885,N_2166);
or U5633 (N_5633,N_3894,N_2714);
and U5634 (N_5634,N_1332,N_4038);
or U5635 (N_5635,N_1497,N_2499);
or U5636 (N_5636,N_929,N_3975);
nor U5637 (N_5637,N_1263,N_414);
nor U5638 (N_5638,N_3173,N_2749);
or U5639 (N_5639,N_3204,N_4308);
nand U5640 (N_5640,N_152,N_1246);
nor U5641 (N_5641,N_504,N_2999);
or U5642 (N_5642,N_1641,N_4209);
nor U5643 (N_5643,N_243,N_1649);
nand U5644 (N_5644,N_4282,N_2925);
nor U5645 (N_5645,N_1092,N_3266);
nor U5646 (N_5646,N_329,N_3967);
nor U5647 (N_5647,N_1488,N_242);
nand U5648 (N_5648,N_3929,N_2601);
nor U5649 (N_5649,N_2075,N_2293);
or U5650 (N_5650,N_3244,N_3719);
nand U5651 (N_5651,N_710,N_3068);
nand U5652 (N_5652,N_3741,N_1797);
and U5653 (N_5653,N_3493,N_3924);
nand U5654 (N_5654,N_585,N_2722);
nand U5655 (N_5655,N_1845,N_4268);
nand U5656 (N_5656,N_2904,N_3776);
nor U5657 (N_5657,N_3372,N_2459);
and U5658 (N_5658,N_1568,N_1865);
nor U5659 (N_5659,N_33,N_4615);
nor U5660 (N_5660,N_4449,N_1639);
and U5661 (N_5661,N_32,N_2485);
or U5662 (N_5662,N_2609,N_3543);
and U5663 (N_5663,N_1877,N_263);
and U5664 (N_5664,N_919,N_774);
or U5665 (N_5665,N_1604,N_367);
and U5666 (N_5666,N_4923,N_2623);
and U5667 (N_5667,N_452,N_2660);
or U5668 (N_5668,N_4929,N_1501);
or U5669 (N_5669,N_1772,N_2378);
nor U5670 (N_5670,N_1632,N_3367);
and U5671 (N_5671,N_4137,N_4894);
and U5672 (N_5672,N_1816,N_3438);
nor U5673 (N_5673,N_686,N_1621);
and U5674 (N_5674,N_2758,N_1640);
or U5675 (N_5675,N_3615,N_1509);
and U5676 (N_5676,N_2385,N_1767);
nor U5677 (N_5677,N_2537,N_1368);
nor U5678 (N_5678,N_2690,N_4468);
or U5679 (N_5679,N_4592,N_3784);
or U5680 (N_5680,N_4993,N_2586);
or U5681 (N_5681,N_1451,N_1549);
and U5682 (N_5682,N_2569,N_1197);
nor U5683 (N_5683,N_2536,N_3643);
nand U5684 (N_5684,N_1530,N_1703);
nor U5685 (N_5685,N_4696,N_3414);
nand U5686 (N_5686,N_187,N_1977);
and U5687 (N_5687,N_1321,N_1727);
or U5688 (N_5688,N_3203,N_4461);
nor U5689 (N_5689,N_1522,N_4276);
and U5690 (N_5690,N_2529,N_3387);
nor U5691 (N_5691,N_1643,N_652);
or U5692 (N_5692,N_2232,N_3932);
nand U5693 (N_5693,N_58,N_2313);
and U5694 (N_5694,N_1753,N_2123);
and U5695 (N_5695,N_565,N_3976);
xnor U5696 (N_5696,N_2937,N_1731);
nand U5697 (N_5697,N_3552,N_3758);
and U5698 (N_5698,N_4444,N_3851);
or U5699 (N_5699,N_4804,N_2039);
and U5700 (N_5700,N_3882,N_4513);
and U5701 (N_5701,N_17,N_2037);
and U5702 (N_5702,N_849,N_3517);
or U5703 (N_5703,N_3137,N_2933);
or U5704 (N_5704,N_3869,N_922);
and U5705 (N_5705,N_1188,N_3735);
or U5706 (N_5706,N_4735,N_1553);
nor U5707 (N_5707,N_757,N_4517);
or U5708 (N_5708,N_4584,N_4581);
nor U5709 (N_5709,N_513,N_3642);
nand U5710 (N_5710,N_220,N_1459);
nand U5711 (N_5711,N_697,N_3482);
nor U5712 (N_5712,N_3933,N_1163);
nor U5713 (N_5713,N_1133,N_2907);
nand U5714 (N_5714,N_4462,N_3964);
nand U5715 (N_5715,N_4015,N_931);
or U5716 (N_5716,N_3293,N_1218);
and U5717 (N_5717,N_3528,N_1637);
and U5718 (N_5718,N_1388,N_308);
or U5719 (N_5719,N_170,N_324);
and U5720 (N_5720,N_4594,N_3828);
nor U5721 (N_5721,N_1794,N_1399);
and U5722 (N_5722,N_1264,N_1983);
and U5723 (N_5723,N_703,N_1980);
nor U5724 (N_5724,N_1252,N_3405);
nor U5725 (N_5725,N_847,N_1853);
or U5726 (N_5726,N_175,N_1506);
nand U5727 (N_5727,N_3904,N_416);
or U5728 (N_5728,N_3917,N_4579);
or U5729 (N_5729,N_1354,N_118);
nor U5730 (N_5730,N_2822,N_3401);
nand U5731 (N_5731,N_1323,N_262);
nand U5732 (N_5732,N_338,N_4067);
nand U5733 (N_5733,N_4532,N_827);
and U5734 (N_5734,N_2227,N_2936);
nand U5735 (N_5735,N_2988,N_1550);
and U5736 (N_5736,N_776,N_1860);
and U5737 (N_5737,N_4394,N_3036);
or U5738 (N_5738,N_4064,N_4355);
or U5739 (N_5739,N_445,N_4050);
nand U5740 (N_5740,N_1578,N_1244);
or U5741 (N_5741,N_4571,N_2967);
nand U5742 (N_5742,N_1482,N_1664);
or U5743 (N_5743,N_4956,N_3646);
or U5744 (N_5744,N_641,N_2292);
and U5745 (N_5745,N_4925,N_635);
nor U5746 (N_5746,N_4060,N_4627);
nor U5747 (N_5747,N_4980,N_2960);
nor U5748 (N_5748,N_3046,N_1827);
nand U5749 (N_5749,N_1144,N_4441);
nand U5750 (N_5750,N_4765,N_735);
nand U5751 (N_5751,N_2759,N_3255);
xor U5752 (N_5752,N_4952,N_2041);
nand U5753 (N_5753,N_2464,N_2910);
or U5754 (N_5754,N_927,N_2058);
xnor U5755 (N_5755,N_4613,N_1201);
and U5756 (N_5756,N_3350,N_722);
nand U5757 (N_5757,N_4747,N_2587);
or U5758 (N_5758,N_932,N_179);
nand U5759 (N_5759,N_401,N_1015);
and U5760 (N_5760,N_1884,N_4390);
xnor U5761 (N_5761,N_3370,N_4843);
or U5762 (N_5762,N_4277,N_1374);
and U5763 (N_5763,N_2175,N_915);
and U5764 (N_5764,N_3721,N_705);
nand U5765 (N_5765,N_1847,N_3890);
and U5766 (N_5766,N_488,N_2517);
and U5767 (N_5767,N_4814,N_3951);
or U5768 (N_5768,N_2222,N_197);
or U5769 (N_5769,N_2216,N_3587);
xnor U5770 (N_5770,N_4231,N_428);
nor U5771 (N_5771,N_2504,N_2658);
nor U5772 (N_5772,N_643,N_2809);
nor U5773 (N_5773,N_140,N_3959);
or U5774 (N_5774,N_3829,N_2859);
nand U5775 (N_5775,N_3051,N_355);
and U5776 (N_5776,N_1393,N_3384);
nor U5777 (N_5777,N_1658,N_4907);
or U5778 (N_5778,N_3592,N_2319);
nor U5779 (N_5779,N_120,N_3336);
and U5780 (N_5780,N_2610,N_3205);
or U5781 (N_5781,N_2512,N_4345);
or U5782 (N_5782,N_4483,N_3231);
and U5783 (N_5783,N_2261,N_2249);
or U5784 (N_5784,N_1183,N_650);
and U5785 (N_5785,N_2080,N_295);
nor U5786 (N_5786,N_855,N_4998);
or U5787 (N_5787,N_1071,N_1146);
or U5788 (N_5788,N_543,N_4216);
or U5789 (N_5789,N_4949,N_4161);
xnor U5790 (N_5790,N_3276,N_2837);
nor U5791 (N_5791,N_2234,N_4398);
nand U5792 (N_5792,N_2795,N_958);
or U5793 (N_5793,N_4802,N_3919);
nand U5794 (N_5794,N_71,N_1342);
or U5795 (N_5795,N_387,N_4916);
nand U5796 (N_5796,N_2981,N_1142);
nor U5797 (N_5797,N_1803,N_384);
nand U5798 (N_5798,N_3022,N_4712);
and U5799 (N_5799,N_913,N_2489);
or U5800 (N_5800,N_137,N_4955);
or U5801 (N_5801,N_281,N_2400);
and U5802 (N_5802,N_110,N_3428);
nor U5803 (N_5803,N_3745,N_2846);
nor U5804 (N_5804,N_1646,N_4215);
nor U5805 (N_5805,N_4529,N_2116);
or U5806 (N_5806,N_2476,N_3781);
nand U5807 (N_5807,N_917,N_391);
nand U5808 (N_5808,N_2557,N_1883);
nand U5809 (N_5809,N_3660,N_3473);
or U5810 (N_5810,N_4622,N_1452);
xnor U5811 (N_5811,N_606,N_443);
and U5812 (N_5812,N_2870,N_2977);
or U5813 (N_5813,N_4159,N_1504);
or U5814 (N_5814,N_3412,N_2151);
or U5815 (N_5815,N_2798,N_4554);
or U5816 (N_5816,N_4758,N_3806);
nor U5817 (N_5817,N_3902,N_3950);
or U5818 (N_5818,N_1591,N_1982);
or U5819 (N_5819,N_2425,N_451);
nor U5820 (N_5820,N_4279,N_2627);
and U5821 (N_5821,N_4906,N_3867);
nor U5822 (N_5822,N_3360,N_3546);
nor U5823 (N_5823,N_2451,N_3447);
nand U5824 (N_5824,N_2603,N_1657);
nand U5825 (N_5825,N_193,N_3148);
nor U5826 (N_5826,N_4452,N_2106);
nor U5827 (N_5827,N_3139,N_801);
nor U5828 (N_5828,N_2555,N_1595);
xnor U5829 (N_5829,N_1219,N_978);
and U5830 (N_5830,N_1329,N_1563);
nor U5831 (N_5831,N_1708,N_4224);
nand U5832 (N_5832,N_2212,N_389);
or U5833 (N_5833,N_1920,N_4115);
and U5834 (N_5834,N_2721,N_4031);
nand U5835 (N_5835,N_1798,N_4948);
nand U5836 (N_5836,N_1787,N_500);
nand U5837 (N_5837,N_987,N_2927);
or U5838 (N_5838,N_4518,N_3058);
nor U5839 (N_5839,N_254,N_671);
and U5840 (N_5840,N_4635,N_4927);
or U5841 (N_5841,N_2446,N_712);
or U5842 (N_5842,N_3441,N_336);
or U5843 (N_5843,N_2285,N_205);
nor U5844 (N_5844,N_3541,N_1536);
nand U5845 (N_5845,N_3442,N_2652);
and U5846 (N_5846,N_4868,N_1106);
or U5847 (N_5847,N_638,N_2450);
nor U5848 (N_5848,N_4790,N_168);
nor U5849 (N_5849,N_368,N_3025);
or U5850 (N_5850,N_1867,N_2582);
or U5851 (N_5851,N_2024,N_1601);
nor U5852 (N_5852,N_1769,N_4453);
xnor U5853 (N_5853,N_524,N_684);
or U5854 (N_5854,N_2457,N_1164);
or U5855 (N_5855,N_4163,N_108);
or U5856 (N_5856,N_3481,N_1870);
or U5857 (N_5857,N_435,N_2802);
nor U5858 (N_5858,N_4415,N_331);
nor U5859 (N_5859,N_2097,N_514);
nand U5860 (N_5860,N_3488,N_3150);
and U5861 (N_5861,N_4829,N_694);
nor U5862 (N_5862,N_2804,N_769);
or U5863 (N_5863,N_2892,N_3153);
nand U5864 (N_5864,N_4725,N_977);
and U5865 (N_5865,N_3754,N_3568);
nand U5866 (N_5866,N_3812,N_4332);
nand U5867 (N_5867,N_4972,N_4561);
nand U5868 (N_5868,N_496,N_2132);
or U5869 (N_5869,N_2463,N_1633);
or U5870 (N_5870,N_4336,N_2924);
nor U5871 (N_5871,N_3811,N_2800);
nand U5872 (N_5872,N_3094,N_1083);
nor U5873 (N_5873,N_3941,N_3875);
nor U5874 (N_5874,N_477,N_190);
nand U5875 (N_5875,N_1519,N_2680);
nor U5876 (N_5876,N_2628,N_4260);
nand U5877 (N_5877,N_2827,N_4074);
nand U5878 (N_5878,N_3212,N_1864);
and U5879 (N_5879,N_2139,N_4564);
or U5880 (N_5880,N_4170,N_3765);
and U5881 (N_5881,N_1543,N_1730);
nand U5882 (N_5882,N_1026,N_640);
and U5883 (N_5883,N_4840,N_2713);
nand U5884 (N_5884,N_2327,N_4808);
or U5885 (N_5885,N_2595,N_2066);
nand U5886 (N_5886,N_4235,N_3515);
nand U5887 (N_5887,N_1539,N_1565);
nand U5888 (N_5888,N_317,N_3704);
nand U5889 (N_5889,N_470,N_2771);
or U5890 (N_5890,N_1235,N_4565);
and U5891 (N_5891,N_3010,N_4753);
or U5892 (N_5892,N_2823,N_3129);
nand U5893 (N_5893,N_3647,N_405);
nand U5894 (N_5894,N_2412,N_3767);
nand U5895 (N_5895,N_1340,N_1260);
and U5896 (N_5896,N_2939,N_314);
and U5897 (N_5897,N_4811,N_2742);
or U5898 (N_5898,N_3944,N_3270);
nor U5899 (N_5899,N_3319,N_2326);
and U5900 (N_5900,N_266,N_4799);
and U5901 (N_5901,N_2842,N_2162);
nor U5902 (N_5902,N_4103,N_72);
nor U5903 (N_5903,N_3506,N_2852);
or U5904 (N_5904,N_4979,N_353);
nor U5905 (N_5905,N_2527,N_4511);
or U5906 (N_5906,N_3003,N_2589);
nor U5907 (N_5907,N_790,N_1349);
and U5908 (N_5908,N_2901,N_219);
or U5909 (N_5909,N_4104,N_1372);
nand U5910 (N_5910,N_2531,N_4866);
or U5911 (N_5911,N_3099,N_3246);
nor U5912 (N_5912,N_2876,N_834);
nor U5913 (N_5913,N_2256,N_2645);
and U5914 (N_5914,N_3631,N_2631);
or U5915 (N_5915,N_2931,N_4106);
or U5916 (N_5916,N_4128,N_3985);
nor U5917 (N_5917,N_4143,N_2519);
or U5918 (N_5918,N_1965,N_2012);
nor U5919 (N_5919,N_437,N_2812);
and U5920 (N_5920,N_4759,N_4619);
nand U5921 (N_5921,N_283,N_1711);
and U5922 (N_5922,N_2868,N_3588);
and U5923 (N_5923,N_2741,N_808);
and U5924 (N_5924,N_2813,N_4365);
nand U5925 (N_5925,N_2237,N_4467);
nand U5926 (N_5926,N_2916,N_4007);
nand U5927 (N_5927,N_1566,N_4873);
or U5928 (N_5928,N_348,N_4213);
nor U5929 (N_5929,N_275,N_2403);
and U5930 (N_5930,N_2192,N_4192);
nor U5931 (N_5931,N_4567,N_1076);
and U5932 (N_5932,N_1465,N_1137);
nand U5933 (N_5933,N_870,N_321);
and U5934 (N_5934,N_2218,N_1135);
nand U5935 (N_5935,N_3549,N_568);
nor U5936 (N_5936,N_683,N_1165);
or U5937 (N_5937,N_3513,N_2989);
nor U5938 (N_5938,N_1941,N_2291);
or U5939 (N_5939,N_327,N_655);
nand U5940 (N_5940,N_787,N_1241);
nand U5941 (N_5941,N_3242,N_3261);
and U5942 (N_5942,N_1110,N_1284);
or U5943 (N_5943,N_798,N_867);
nand U5944 (N_5944,N_3771,N_3559);
nand U5945 (N_5945,N_1019,N_4142);
and U5946 (N_5946,N_570,N_2010);
and U5947 (N_5947,N_1057,N_1339);
nor U5948 (N_5948,N_786,N_534);
nand U5949 (N_5949,N_4249,N_1773);
nand U5950 (N_5950,N_4683,N_3683);
and U5951 (N_5951,N_2502,N_2170);
nand U5952 (N_5952,N_1089,N_4130);
or U5953 (N_5953,N_4229,N_4861);
nand U5954 (N_5954,N_10,N_1486);
xnor U5955 (N_5955,N_3262,N_668);
xnor U5956 (N_5956,N_3518,N_3789);
and U5957 (N_5957,N_740,N_2310);
nor U5958 (N_5958,N_2761,N_346);
and U5959 (N_5959,N_4110,N_4138);
or U5960 (N_5960,N_4166,N_3946);
and U5961 (N_5961,N_1367,N_4435);
nand U5962 (N_5962,N_3834,N_4805);
nor U5963 (N_5963,N_4362,N_3888);
nand U5964 (N_5964,N_116,N_4800);
or U5965 (N_5965,N_2240,N_2157);
nor U5966 (N_5966,N_2188,N_1033);
nand U5967 (N_5967,N_3501,N_4121);
nand U5968 (N_5968,N_1118,N_4144);
or U5969 (N_5969,N_1981,N_4705);
nor U5970 (N_5970,N_4672,N_1077);
nand U5971 (N_5971,N_3440,N_1335);
nor U5972 (N_5972,N_2632,N_113);
and U5973 (N_5973,N_3526,N_4117);
nand U5974 (N_5974,N_1490,N_4459);
and U5975 (N_5975,N_3661,N_192);
and U5976 (N_5976,N_4255,N_8);
and U5977 (N_5977,N_843,N_3866);
and U5978 (N_5978,N_392,N_3143);
nand U5979 (N_5979,N_3634,N_2161);
xor U5980 (N_5980,N_4795,N_850);
or U5981 (N_5981,N_515,N_4690);
nand U5982 (N_5982,N_1776,N_1426);
and U5983 (N_5983,N_3622,N_447);
and U5984 (N_5984,N_3800,N_865);
nor U5985 (N_5985,N_2278,N_4490);
or U5986 (N_5986,N_3237,N_4487);
and U5987 (N_5987,N_1045,N_3563);
and U5988 (N_5988,N_4947,N_1780);
and U5989 (N_5989,N_2847,N_2898);
nand U5990 (N_5990,N_4299,N_3083);
or U5991 (N_5991,N_3570,N_53);
or U5992 (N_5992,N_3317,N_772);
nand U5993 (N_5993,N_3598,N_3979);
and U5994 (N_5994,N_4181,N_4098);
nand U5995 (N_5995,N_1627,N_3385);
nor U5996 (N_5996,N_3859,N_4806);
and U5997 (N_5997,N_3282,N_3337);
nor U5998 (N_5998,N_2406,N_2567);
and U5999 (N_5999,N_2560,N_1065);
nand U6000 (N_6000,N_4819,N_1059);
nor U6001 (N_6001,N_2498,N_2679);
nor U6002 (N_6002,N_986,N_1379);
and U6003 (N_6003,N_2320,N_997);
nor U6004 (N_6004,N_3443,N_3033);
xnor U6005 (N_6005,N_1385,N_1909);
nand U6006 (N_6006,N_4875,N_150);
nand U6007 (N_6007,N_1740,N_954);
and U6008 (N_6008,N_1460,N_3049);
or U6009 (N_6009,N_3652,N_1656);
or U6010 (N_6010,N_1419,N_4932);
or U6011 (N_6011,N_3471,N_4724);
nor U6012 (N_6012,N_4670,N_4773);
or U6013 (N_6013,N_2074,N_1149);
and U6014 (N_6014,N_3052,N_4679);
or U6015 (N_6015,N_2350,N_3821);
and U6016 (N_6016,N_747,N_1917);
and U6017 (N_6017,N_1957,N_2544);
or U6018 (N_6018,N_4536,N_708);
nor U6019 (N_6019,N_2009,N_3848);
and U6020 (N_6020,N_765,N_1290);
nor U6021 (N_6021,N_3318,N_2568);
and U6022 (N_6022,N_3512,N_1754);
or U6023 (N_6023,N_1225,N_4334);
nor U6024 (N_6024,N_3619,N_1849);
or U6025 (N_6025,N_4309,N_2791);
and U6026 (N_6026,N_3939,N_1858);
and U6027 (N_6027,N_3790,N_4306);
and U6028 (N_6028,N_4236,N_2505);
and U6029 (N_6029,N_876,N_1396);
nand U6030 (N_6030,N_1217,N_3783);
nor U6031 (N_6031,N_4642,N_2994);
nor U6032 (N_6032,N_3095,N_3576);
or U6033 (N_6033,N_789,N_704);
or U6034 (N_6034,N_3444,N_1158);
nand U6035 (N_6035,N_1696,N_2040);
and U6036 (N_6036,N_4220,N_4751);
nor U6037 (N_6037,N_3430,N_115);
nor U6038 (N_6038,N_3069,N_4892);
or U6039 (N_6039,N_2129,N_45);
nor U6040 (N_6040,N_3445,N_2328);
or U6041 (N_6041,N_580,N_780);
nor U6042 (N_6042,N_4485,N_2019);
or U6043 (N_6043,N_858,N_4639);
or U6044 (N_6044,N_3306,N_3692);
nor U6045 (N_6045,N_2699,N_3832);
nor U6046 (N_6046,N_2452,N_2873);
and U6047 (N_6047,N_1868,N_102);
nor U6048 (N_6048,N_3486,N_4838);
and U6049 (N_6049,N_4388,N_2426);
nand U6050 (N_6050,N_4974,N_1113);
or U6051 (N_6051,N_4965,N_2243);
nor U6052 (N_6052,N_4134,N_2174);
or U6053 (N_6053,N_2733,N_768);
nand U6054 (N_6054,N_1960,N_1454);
or U6055 (N_6055,N_3053,N_498);
and U6056 (N_6056,N_1175,N_494);
nor U6057 (N_6057,N_4661,N_4086);
nor U6058 (N_6058,N_3067,N_99);
nor U6059 (N_6059,N_4211,N_887);
xor U6060 (N_6060,N_52,N_1819);
and U6061 (N_6061,N_1761,N_4942);
and U6062 (N_6062,N_246,N_382);
or U6063 (N_6063,N_2592,N_2137);
xor U6064 (N_6064,N_4898,N_4222);
and U6065 (N_6065,N_1037,N_2085);
or U6066 (N_6066,N_2178,N_2299);
nor U6067 (N_6067,N_770,N_1480);
or U6068 (N_6068,N_2760,N_1887);
or U6069 (N_6069,N_3840,N_4285);
nor U6070 (N_6070,N_1674,N_1346);
and U6071 (N_6071,N_4363,N_1663);
nor U6072 (N_6072,N_1475,N_144);
nor U6073 (N_6073,N_4611,N_4726);
and U6074 (N_6074,N_2732,N_3669);
nor U6075 (N_6075,N_75,N_4109);
nand U6076 (N_6076,N_3658,N_3322);
nor U6077 (N_6077,N_767,N_4537);
or U6078 (N_6078,N_375,N_1808);
nand U6079 (N_6079,N_4698,N_3901);
or U6080 (N_6080,N_1208,N_3892);
nor U6081 (N_6081,N_3842,N_2189);
nor U6082 (N_6082,N_64,N_4469);
and U6083 (N_6083,N_1141,N_1635);
or U6084 (N_6084,N_4310,N_750);
nor U6085 (N_6085,N_2169,N_3611);
nor U6086 (N_6086,N_1337,N_153);
nor U6087 (N_6087,N_4287,N_127);
or U6088 (N_6088,N_4164,N_928);
xnor U6089 (N_6089,N_3507,N_2230);
nor U6090 (N_6090,N_3235,N_2422);
nand U6091 (N_6091,N_3873,N_4027);
and U6092 (N_6092,N_4503,N_2046);
nand U6093 (N_6093,N_884,N_1985);
or U6094 (N_6094,N_4558,N_3609);
nand U6095 (N_6095,N_4976,N_3948);
nor U6096 (N_6096,N_2572,N_2399);
or U6097 (N_6097,N_527,N_2387);
nor U6098 (N_6098,N_1120,N_4381);
or U6099 (N_6099,N_2672,N_1259);
or U6100 (N_6100,N_1859,N_2322);
and U6101 (N_6101,N_3498,N_3391);
or U6102 (N_6102,N_4556,N_454);
or U6103 (N_6103,N_1129,N_3499);
and U6104 (N_6104,N_2701,N_57);
nand U6105 (N_6105,N_4688,N_1272);
nand U6106 (N_6106,N_4205,N_2727);
nand U6107 (N_6107,N_2416,N_1431);
or U6108 (N_6108,N_2303,N_3560);
and U6109 (N_6109,N_4418,N_1318);
or U6110 (N_6110,N_1961,N_2349);
nand U6111 (N_6111,N_256,N_3572);
nand U6112 (N_6112,N_182,N_3144);
nor U6113 (N_6113,N_3327,N_138);
nor U6114 (N_6114,N_1610,N_2874);
and U6115 (N_6115,N_3756,N_4162);
nor U6116 (N_6116,N_2159,N_796);
and U6117 (N_6117,N_1763,N_4608);
and U6118 (N_6118,N_3221,N_2552);
or U6119 (N_6119,N_991,N_238);
or U6120 (N_6120,N_202,N_4425);
and U6121 (N_6121,N_4997,N_2858);
or U6122 (N_6122,N_3197,N_2928);
or U6123 (N_6123,N_2115,N_2947);
xor U6124 (N_6124,N_2205,N_4406);
xnor U6125 (N_6125,N_2131,N_1882);
nand U6126 (N_6126,N_4845,N_1461);
nor U6127 (N_6127,N_4741,N_1301);
nor U6128 (N_6128,N_1467,N_347);
or U6129 (N_6129,N_2957,N_3001);
nand U6130 (N_6130,N_1821,N_1390);
or U6131 (N_6131,N_1282,N_754);
and U6132 (N_6132,N_1534,N_2315);
or U6133 (N_6133,N_564,N_82);
or U6134 (N_6134,N_1181,N_1487);
nor U6135 (N_6135,N_4954,N_62);
nand U6136 (N_6136,N_4754,N_4065);
nor U6137 (N_6137,N_1889,N_760);
nand U6138 (N_6138,N_3192,N_3307);
and U6139 (N_6139,N_2995,N_2264);
and U6140 (N_6140,N_1300,N_1838);
and U6141 (N_6141,N_4450,N_2889);
nand U6142 (N_6142,N_4204,N_1823);
and U6143 (N_6143,N_2369,N_2700);
or U6144 (N_6144,N_695,N_885);
nand U6145 (N_6145,N_199,N_1414);
or U6146 (N_6146,N_2523,N_4051);
or U6147 (N_6147,N_4603,N_1293);
nor U6148 (N_6148,N_3701,N_3729);
or U6149 (N_6149,N_729,N_1995);
nor U6150 (N_6150,N_3236,N_3489);
nor U6151 (N_6151,N_1481,N_2146);
nand U6152 (N_6152,N_2124,N_3019);
and U6153 (N_6153,N_3544,N_4225);
and U6154 (N_6154,N_3550,N_1430);
nor U6155 (N_6155,N_4203,N_4607);
nor U6156 (N_6156,N_624,N_1210);
or U6157 (N_6157,N_2287,N_2915);
or U6158 (N_6158,N_4928,N_2147);
or U6159 (N_6159,N_893,N_1131);
nor U6160 (N_6160,N_74,N_3814);
nand U6161 (N_6161,N_2815,N_3216);
or U6162 (N_6162,N_4423,N_723);
nor U6163 (N_6163,N_4681,N_4147);
or U6164 (N_6164,N_232,N_2331);
or U6165 (N_6165,N_822,N_2130);
or U6166 (N_6166,N_4574,N_1400);
or U6167 (N_6167,N_3241,N_1728);
and U6168 (N_6168,N_2958,N_3418);
nor U6169 (N_6169,N_1721,N_871);
and U6170 (N_6170,N_4807,N_1172);
xor U6171 (N_6171,N_2864,N_1953);
nor U6172 (N_6172,N_1234,N_3824);
or U6173 (N_6173,N_2472,N_143);
or U6174 (N_6174,N_1533,N_4304);
or U6175 (N_6175,N_923,N_1068);
nand U6176 (N_6176,N_207,N_4734);
and U6177 (N_6177,N_3664,N_1109);
nand U6178 (N_6178,N_492,N_1540);
and U6179 (N_6179,N_3008,N_992);
or U6180 (N_6180,N_2316,N_3870);
nand U6181 (N_6181,N_352,N_1836);
or U6182 (N_6182,N_1828,N_155);
and U6183 (N_6183,N_364,N_1653);
nand U6184 (N_6184,N_3712,N_1166);
nand U6185 (N_6185,N_1105,N_1178);
or U6186 (N_6186,N_1182,N_734);
and U6187 (N_6187,N_4820,N_3597);
nor U6188 (N_6188,N_746,N_1670);
and U6189 (N_6189,N_4606,N_902);
and U6190 (N_6190,N_4634,N_4320);
or U6191 (N_6191,N_4026,N_562);
or U6192 (N_6192,N_552,N_85);
nand U6193 (N_6193,N_1192,N_3724);
or U6194 (N_6194,N_681,N_4803);
nor U6195 (N_6195,N_2135,N_2190);
nor U6196 (N_6196,N_1180,N_4364);
nand U6197 (N_6197,N_3928,N_1722);
or U6198 (N_6198,N_1938,N_3267);
nand U6199 (N_6199,N_575,N_1666);
and U6200 (N_6200,N_3556,N_3793);
and U6201 (N_6201,N_448,N_2283);
nand U6202 (N_6202,N_3348,N_1930);
and U6203 (N_6203,N_2093,N_2768);
nand U6204 (N_6204,N_4132,N_4897);
nand U6205 (N_6205,N_1189,N_2860);
nand U6206 (N_6206,N_3042,N_930);
or U6207 (N_6207,N_837,N_2890);
xnor U6208 (N_6208,N_4063,N_4438);
nand U6209 (N_6209,N_2856,N_1273);
or U6210 (N_6210,N_4179,N_3898);
or U6211 (N_6211,N_1863,N_3059);
nand U6212 (N_6212,N_4784,N_3111);
or U6213 (N_6213,N_4757,N_3778);
and U6214 (N_6214,N_2919,N_4075);
nor U6215 (N_6215,N_3112,N_1676);
and U6216 (N_6216,N_3981,N_3230);
and U6217 (N_6217,N_1364,N_4293);
or U6218 (N_6218,N_1101,N_4037);
xor U6219 (N_6219,N_1677,N_2832);
or U6220 (N_6220,N_185,N_2853);
nor U6221 (N_6221,N_3238,N_4505);
nor U6222 (N_6222,N_2337,N_1062);
nor U6223 (N_6223,N_2000,N_1508);
nor U6224 (N_6224,N_2747,N_4684);
nand U6225 (N_6225,N_1952,N_2648);
nor U6226 (N_6226,N_4376,N_3132);
nand U6227 (N_6227,N_1954,N_224);
and U6228 (N_6228,N_3013,N_289);
nor U6229 (N_6229,N_3573,N_3595);
nand U6230 (N_6230,N_1942,N_846);
or U6231 (N_6231,N_2201,N_1660);
or U6232 (N_6232,N_944,N_2797);
nor U6233 (N_6233,N_2533,N_3678);
or U6234 (N_6234,N_1799,N_3648);
nor U6235 (N_6235,N_1612,N_2828);
nand U6236 (N_6236,N_2160,N_4732);
and U6237 (N_6237,N_1715,N_1155);
nand U6238 (N_6238,N_418,N_2740);
or U6239 (N_6239,N_1829,N_1013);
and U6240 (N_6240,N_4154,N_4036);
nand U6241 (N_6241,N_1055,N_3732);
nand U6242 (N_6242,N_4520,N_3640);
or U6243 (N_6243,N_1004,N_248);
nor U6244 (N_6244,N_3474,N_2078);
nand U6245 (N_6245,N_634,N_3047);
nand U6246 (N_6246,N_1473,N_489);
nand U6247 (N_6247,N_1611,N_1395);
or U6248 (N_6248,N_1634,N_393);
nand U6249 (N_6249,N_3987,N_4920);
nor U6250 (N_6250,N_4274,N_2032);
nor U6251 (N_6251,N_4061,N_540);
nand U6252 (N_6252,N_2509,N_3308);
or U6253 (N_6253,N_4902,N_2398);
nor U6254 (N_6254,N_3547,N_3061);
nand U6255 (N_6255,N_468,N_2869);
nand U6256 (N_6256,N_3199,N_1236);
and U6257 (N_6257,N_821,N_299);
nand U6258 (N_6258,N_1351,N_4723);
and U6259 (N_6259,N_4424,N_1525);
xor U6260 (N_6260,N_4359,N_3620);
nor U6261 (N_6261,N_3846,N_590);
or U6262 (N_6262,N_1503,N_4456);
and U6263 (N_6263,N_2861,N_4372);
or U6264 (N_6264,N_2906,N_1325);
nor U6265 (N_6265,N_2029,N_2987);
nor U6266 (N_6266,N_2681,N_4506);
nand U6267 (N_6267,N_91,N_2877);
nor U6268 (N_6268,N_1308,N_2694);
or U6269 (N_6269,N_3937,N_2710);
nor U6270 (N_6270,N_4889,N_2878);
and U6271 (N_6271,N_3265,N_4288);
nor U6272 (N_6272,N_4298,N_456);
nor U6273 (N_6273,N_2420,N_1620);
and U6274 (N_6274,N_3381,N_409);
or U6275 (N_6275,N_290,N_2109);
or U6276 (N_6276,N_1662,N_1028);
and U6277 (N_6277,N_1793,N_270);
and U6278 (N_6278,N_2467,N_1607);
nor U6279 (N_6279,N_1239,N_2911);
and U6280 (N_6280,N_890,N_914);
or U6281 (N_6281,N_4748,N_2341);
or U6282 (N_6282,N_1956,N_3639);
and U6283 (N_6283,N_829,N_4313);
and U6284 (N_6284,N_785,N_3122);
and U6285 (N_6285,N_167,N_1427);
and U6286 (N_6286,N_2252,N_3696);
and U6287 (N_6287,N_189,N_1989);
nand U6288 (N_6288,N_1720,N_429);
nand U6289 (N_6289,N_2550,N_3478);
and U6290 (N_6290,N_2441,N_3138);
nor U6291 (N_6291,N_2112,N_484);
nor U6292 (N_6292,N_4957,N_1052);
or U6293 (N_6293,N_756,N_3463);
or U6294 (N_6294,N_2644,N_3909);
or U6295 (N_6295,N_2384,N_4045);
nand U6296 (N_6296,N_3402,N_84);
nand U6297 (N_6297,N_3569,N_4772);
or U6298 (N_6298,N_20,N_2107);
nand U6299 (N_6299,N_980,N_610);
and U6300 (N_6300,N_2302,N_838);
nand U6301 (N_6301,N_2824,N_3903);
nor U6302 (N_6302,N_1872,N_3426);
or U6303 (N_6303,N_4344,N_4079);
nand U6304 (N_6304,N_2841,N_982);
or U6305 (N_6305,N_4926,N_1785);
or U6306 (N_6306,N_1891,N_3565);
nor U6307 (N_6307,N_441,N_4331);
nor U6308 (N_6308,N_1251,N_1990);
nand U6309 (N_6309,N_532,N_1187);
nor U6310 (N_6310,N_4191,N_2006);
or U6311 (N_6311,N_4609,N_2454);
nor U6312 (N_6312,N_1770,N_4604);
and U6313 (N_6313,N_272,N_3599);
xor U6314 (N_6314,N_3768,N_1918);
nand U6315 (N_6315,N_4146,N_1122);
nor U6316 (N_6316,N_4207,N_1370);
and U6317 (N_6317,N_1531,N_4891);
or U6318 (N_6318,N_3377,N_1834);
nor U6319 (N_6319,N_3108,N_2298);
and U6320 (N_6320,N_4316,N_4296);
and U6321 (N_6321,N_1086,N_169);
and U6322 (N_6322,N_3533,N_1227);
nor U6323 (N_6323,N_2561,N_1719);
nor U6324 (N_6324,N_4434,N_3746);
nor U6325 (N_6325,N_3510,N_3424);
nor U6326 (N_6326,N_4950,N_3720);
or U6327 (N_6327,N_311,N_3623);
and U6328 (N_6328,N_3797,N_545);
or U6329 (N_6329,N_388,N_3291);
or U6330 (N_6330,N_1215,N_888);
xor U6331 (N_6331,N_1824,N_23);
or U6332 (N_6332,N_1691,N_4995);
or U6333 (N_6333,N_4888,N_3786);
nand U6334 (N_6334,N_1174,N_2785);
or U6335 (N_6335,N_942,N_3118);
and U6336 (N_6336,N_2127,N_1671);
xnor U6337 (N_6337,N_3459,N_491);
or U6338 (N_6338,N_2684,N_344);
and U6339 (N_6339,N_1237,N_340);
and U6340 (N_6340,N_2799,N_1448);
or U6341 (N_6341,N_133,N_312);
or U6342 (N_6342,N_521,N_4428);
nor U6343 (N_6343,N_2554,N_2236);
nand U6344 (N_6344,N_1690,N_730);
nand U6345 (N_6345,N_4087,N_4641);
or U6346 (N_6346,N_3073,N_691);
nor U6347 (N_6347,N_1381,N_646);
nand U6348 (N_6348,N_4677,N_1739);
and U6349 (N_6349,N_1673,N_1063);
nand U6350 (N_6350,N_1476,N_4124);
or U6351 (N_6351,N_3368,N_3989);
and U6352 (N_6352,N_4922,N_4961);
or U6353 (N_6353,N_2073,N_3248);
and U6354 (N_6354,N_2840,N_4066);
xnor U6355 (N_6355,N_2789,N_2651);
and U6356 (N_6356,N_3352,N_3245);
and U6357 (N_6357,N_4465,N_3247);
nor U6358 (N_6358,N_1047,N_3168);
and U6359 (N_6359,N_1191,N_881);
or U6360 (N_6360,N_4139,N_4959);
nand U6361 (N_6361,N_1546,N_2280);
or U6362 (N_6362,N_4020,N_341);
nor U6363 (N_6363,N_2669,N_3804);
nand U6364 (N_6364,N_1751,N_4504);
and U6365 (N_6365,N_3214,N_3718);
nand U6366 (N_6366,N_422,N_3503);
and U6367 (N_6367,N_319,N_840);
and U6368 (N_6368,N_579,N_4177);
and U6369 (N_6369,N_2344,N_1420);
and U6370 (N_6370,N_3304,N_908);
nor U6371 (N_6371,N_1371,N_558);
or U6372 (N_6372,N_4937,N_296);
or U6373 (N_6373,N_971,N_3178);
nor U6374 (N_6374,N_2423,N_566);
nor U6375 (N_6375,N_657,N_551);
nand U6376 (N_6376,N_3364,N_1014);
and U6377 (N_6377,N_3617,N_2565);
xnor U6378 (N_6378,N_3130,N_253);
and U6379 (N_6379,N_883,N_339);
and U6380 (N_6380,N_880,N_4650);
nand U6381 (N_6381,N_4918,N_1124);
or U6382 (N_6382,N_2013,N_3433);
or U6383 (N_6383,N_2825,N_664);
nor U6384 (N_6384,N_1023,N_2481);
and U6385 (N_6385,N_901,N_3862);
nand U6386 (N_6386,N_2687,N_4123);
nor U6387 (N_6387,N_1195,N_1505);
or U6388 (N_6388,N_2148,N_2835);
nand U6389 (N_6389,N_3913,N_830);
nand U6390 (N_6390,N_2528,N_3343);
or U6391 (N_6391,N_3253,N_2270);
nor U6392 (N_6392,N_2750,N_825);
nor U6393 (N_6393,N_1231,N_906);
nor U6394 (N_6394,N_3494,N_1974);
nor U6395 (N_6395,N_2314,N_1699);
xnor U6396 (N_6396,N_4246,N_4521);
nand U6397 (N_6397,N_97,N_3561);
and U6398 (N_6398,N_1190,N_2575);
nor U6399 (N_6399,N_3857,N_4155);
nor U6400 (N_6400,N_293,N_2253);
nand U6401 (N_6401,N_87,N_1305);
or U6402 (N_6402,N_2896,N_3752);
and U6403 (N_6403,N_399,N_4569);
or U6404 (N_6404,N_2007,N_158);
or U6405 (N_6405,N_4689,N_4695);
nor U6406 (N_6406,N_3048,N_3629);
or U6407 (N_6407,N_177,N_3912);
nand U6408 (N_6408,N_4936,N_1927);
and U6409 (N_6409,N_4951,N_828);
nor U6410 (N_6410,N_146,N_2318);
xnor U6411 (N_6411,N_44,N_2917);
and U6412 (N_6412,N_3349,N_1945);
xor U6413 (N_6413,N_13,N_4848);
or U6414 (N_6414,N_4711,N_4573);
nand U6415 (N_6415,N_3351,N_1777);
xor U6416 (N_6416,N_2333,N_3827);
xor U6417 (N_6417,N_4160,N_3830);
and U6418 (N_6418,N_2678,N_1556);
xnor U6419 (N_6419,N_2208,N_2390);
nor U6420 (N_6420,N_309,N_2488);
and U6421 (N_6421,N_3880,N_3436);
or U6422 (N_6422,N_1281,N_4244);
nand U6423 (N_6423,N_4846,N_439);
nand U6424 (N_6424,N_19,N_1922);
nand U6425 (N_6425,N_3970,N_2250);
nor U6426 (N_6426,N_1397,N_559);
xnor U6427 (N_6427,N_848,N_1198);
nor U6428 (N_6428,N_366,N_2053);
and U6429 (N_6429,N_3470,N_584);
nand U6430 (N_6430,N_1873,N_3905);
nand U6431 (N_6431,N_24,N_2207);
or U6432 (N_6432,N_244,N_3187);
nand U6433 (N_6433,N_4230,N_538);
nor U6434 (N_6434,N_2430,N_4713);
nand U6435 (N_6435,N_1091,N_3542);
or U6436 (N_6436,N_4367,N_1009);
and U6437 (N_6437,N_1038,N_4402);
and U6438 (N_6438,N_3826,N_2360);
and U6439 (N_6439,N_3201,N_560);
or U6440 (N_6440,N_3529,N_2424);
nand U6441 (N_6441,N_2443,N_442);
nor U6442 (N_6442,N_4775,N_2394);
nor U6443 (N_6443,N_2389,N_4934);
nor U6444 (N_6444,N_4426,N_937);
and U6445 (N_6445,N_3578,N_4348);
nand U6446 (N_6446,N_2484,N_4823);
nand U6447 (N_6447,N_2035,N_4335);
or U6448 (N_6448,N_1285,N_2487);
nor U6449 (N_6449,N_4575,N_3123);
xor U6450 (N_6450,N_2938,N_2985);
nand U6451 (N_6451,N_1996,N_4896);
and U6452 (N_6452,N_3277,N_1925);
or U6453 (N_6453,N_3991,N_2577);
or U6454 (N_6454,N_1994,N_4680);
nor U6455 (N_6455,N_2045,N_4482);
nand U6456 (N_6456,N_1126,N_1030);
nor U6457 (N_6457,N_1923,N_3509);
or U6458 (N_6458,N_3739,N_3747);
nor U6459 (N_6459,N_1850,N_4016);
nand U6460 (N_6460,N_800,N_2844);
or U6461 (N_6461,N_3608,N_3450);
or U6462 (N_6462,N_3141,N_1520);
nand U6463 (N_6463,N_2055,N_1436);
or U6464 (N_6464,N_3523,N_4029);
nor U6465 (N_6465,N_1428,N_2633);
or U6466 (N_6466,N_4217,N_3110);
and U6467 (N_6467,N_3335,N_2471);
nor U6468 (N_6468,N_4408,N_3551);
and U6469 (N_6469,N_3713,N_2643);
nor U6470 (N_6470,N_495,N_4135);
and U6471 (N_6471,N_1571,N_818);
nor U6472 (N_6472,N_282,N_2184);
nand U6473 (N_6473,N_4563,N_1661);
nor U6474 (N_6474,N_60,N_2382);
and U6475 (N_6475,N_4755,N_3792);
and U6476 (N_6476,N_3114,N_649);
or U6477 (N_6477,N_1929,N_345);
or U6478 (N_6478,N_31,N_1523);
nor U6479 (N_6479,N_2034,N_4566);
and U6480 (N_6480,N_2596,N_1176);
nor U6481 (N_6481,N_1589,N_1222);
nand U6482 (N_6482,N_2002,N_2891);
and U6483 (N_6483,N_782,N_3819);
nor U6484 (N_6484,N_2729,N_1855);
nor U6485 (N_6485,N_4333,N_3252);
nor U6486 (N_6486,N_410,N_3164);
nand U6487 (N_6487,N_3485,N_2786);
nor U6488 (N_6488,N_3736,N_724);
nor U6489 (N_6489,N_54,N_2079);
or U6490 (N_6490,N_70,N_3341);
or U6491 (N_6491,N_3847,N_505);
or U6492 (N_6492,N_4983,N_4685);
nor U6493 (N_6493,N_4228,N_2365);
nand U6494 (N_6494,N_2744,N_1471);
and U6495 (N_6495,N_3206,N_2935);
nor U6496 (N_6496,N_3539,N_4585);
nor U6497 (N_6497,N_101,N_1093);
nand U6498 (N_6498,N_4384,N_3709);
or U6499 (N_6499,N_824,N_2300);
nand U6500 (N_6500,N_1125,N_325);
nor U6501 (N_6501,N_3969,N_2343);
and U6502 (N_6502,N_2431,N_2764);
and U6503 (N_6503,N_1382,N_1975);
or U6504 (N_6504,N_2913,N_3);
nor U6505 (N_6505,N_4557,N_2932);
or U6506 (N_6506,N_1090,N_4703);
and U6507 (N_6507,N_3303,N_4872);
and U6508 (N_6508,N_4151,N_3251);
or U6509 (N_6509,N_4198,N_4025);
or U6510 (N_6510,N_3538,N_2594);
or U6511 (N_6511,N_896,N_2546);
and U6512 (N_6512,N_3887,N_2366);
nand U6513 (N_6513,N_3772,N_1781);
nand U6514 (N_6514,N_4481,N_1999);
nand U6515 (N_6515,N_965,N_4369);
and U6516 (N_6516,N_2027,N_4436);
and U6517 (N_6517,N_3785,N_3845);
or U6518 (N_6518,N_2880,N_4091);
nand U6519 (N_6519,N_2001,N_820);
nor U6520 (N_6520,N_2089,N_3540);
or U6521 (N_6521,N_374,N_3264);
nand U6522 (N_6522,N_2473,N_4412);
nand U6523 (N_6523,N_2286,N_1791);
xor U6524 (N_6524,N_2206,N_183);
and U6525 (N_6525,N_2204,N_2182);
and U6526 (N_6526,N_485,N_3121);
nor U6527 (N_6527,N_1066,N_993);
and U6528 (N_6528,N_1810,N_2982);
and U6529 (N_6529,N_161,N_1492);
or U6530 (N_6530,N_1622,N_4257);
and U6531 (N_6531,N_4702,N_2325);
or U6532 (N_6532,N_1630,N_1315);
nor U6533 (N_6533,N_1822,N_1812);
or U6534 (N_6534,N_1080,N_2629);
xnor U6535 (N_6535,N_1383,N_1050);
and U6536 (N_6536,N_854,N_2951);
and U6537 (N_6537,N_2453,N_486);
nor U6538 (N_6538,N_3759,N_4968);
nor U6539 (N_6539,N_1069,N_3415);
nor U6540 (N_6540,N_2606,N_1034);
or U6541 (N_6541,N_4391,N_1169);
or U6542 (N_6542,N_2668,N_3195);
nand U6543 (N_6543,N_3714,N_4666);
or U6544 (N_6544,N_690,N_2613);
and U6545 (N_6545,N_3156,N_3484);
nor U6546 (N_6546,N_4736,N_510);
and U6547 (N_6547,N_3773,N_3026);
nor U6548 (N_6548,N_2676,N_2113);
or U6549 (N_6549,N_3292,N_3334);
or U6550 (N_6550,N_555,N_1900);
nor U6551 (N_6551,N_597,N_215);
and U6552 (N_6552,N_4486,N_404);
and U6553 (N_6553,N_990,N_274);
nand U6554 (N_6554,N_2172,N_605);
nor U6555 (N_6555,N_2444,N_2854);
or U6556 (N_6556,N_3899,N_2163);
or U6557 (N_6557,N_2062,N_3591);
and U6558 (N_6558,N_0,N_1528);
nand U6559 (N_6559,N_4495,N_1328);
and U6560 (N_6560,N_1345,N_1404);
and U6561 (N_6561,N_904,N_3511);
and U6562 (N_6562,N_1911,N_693);
nor U6563 (N_6563,N_4545,N_1024);
or U6564 (N_6564,N_3154,N_2969);
or U6565 (N_6565,N_259,N_2084);
and U6566 (N_6566,N_2345,N_2373);
nand U6567 (N_6567,N_1987,N_1079);
and U6568 (N_6568,N_743,N_851);
nor U6569 (N_6569,N_2375,N_3782);
and U6570 (N_6570,N_3686,N_3273);
or U6571 (N_6571,N_2336,N_2839);
or U6572 (N_6572,N_4694,N_1888);
and U6573 (N_6573,N_4044,N_326);
or U6574 (N_6574,N_1311,N_3530);
nand U6575 (N_6575,N_1432,N_2372);
nand U6576 (N_6576,N_2185,N_1758);
nand U6577 (N_6577,N_280,N_2434);
or U6578 (N_6578,N_4480,N_3649);
or U6579 (N_6579,N_736,N_3553);
and U6580 (N_6580,N_4643,N_2042);
and U6581 (N_6581,N_43,N_4253);
nand U6582 (N_6582,N_1391,N_357);
nor U6583 (N_6583,N_2717,N_678);
nand U6584 (N_6584,N_2168,N_1303);
and U6585 (N_6585,N_2367,N_4039);
nor U6586 (N_6586,N_4042,N_2970);
or U6587 (N_6587,N_1466,N_1745);
nor U6588 (N_6588,N_166,N_4190);
nand U6589 (N_6589,N_3420,N_2574);
nand U6590 (N_6590,N_3582,N_4129);
nand U6591 (N_6591,N_4395,N_4946);
or U6592 (N_6592,N_480,N_4612);
and U6593 (N_6593,N_2923,N_3594);
nor U6594 (N_6594,N_1327,N_2067);
or U6595 (N_6595,N_3534,N_4577);
nand U6596 (N_6596,N_415,N_4407);
or U6597 (N_6597,N_4833,N_4497);
or U6598 (N_6598,N_2689,N_3389);
nor U6599 (N_6599,N_2751,N_1733);
nand U6600 (N_6600,N_4202,N_1007);
or U6601 (N_6601,N_1800,N_1484);
or U6602 (N_6602,N_1844,N_934);
or U6603 (N_6603,N_1412,N_2268);
nand U6604 (N_6604,N_1002,N_2682);
or U6605 (N_6605,N_1527,N_675);
and U6606 (N_6606,N_3483,N_436);
xor U6607 (N_6607,N_2656,N_1233);
nor U6608 (N_6608,N_1255,N_1880);
or U6609 (N_6609,N_719,N_996);
and U6610 (N_6610,N_4610,N_967);
nand U6611 (N_6611,N_2121,N_3239);
nand U6612 (N_6612,N_1967,N_4413);
nor U6613 (N_6613,N_630,N_1319);
nand U6614 (N_6614,N_2414,N_2247);
or U6615 (N_6615,N_3397,N_4938);
nor U6616 (N_6616,N_425,N_3853);
nor U6617 (N_6617,N_3354,N_1204);
nor U6618 (N_6618,N_507,N_2311);
and U6619 (N_6619,N_3632,N_2064);
nand U6620 (N_6620,N_4307,N_1672);
xor U6621 (N_6621,N_4887,N_994);
or U6622 (N_6622,N_3799,N_4182);
or U6623 (N_6623,N_3815,N_2117);
nor U6624 (N_6624,N_4744,N_1894);
nor U6625 (N_6625,N_2539,N_1732);
nand U6626 (N_6626,N_1139,N_3803);
and U6627 (N_6627,N_1667,N_2712);
nand U6628 (N_6628,N_4286,N_3889);
nor U6629 (N_6629,N_3863,N_2284);
or U6630 (N_6630,N_4992,N_252);
or U6631 (N_6631,N_12,N_214);
nand U6632 (N_6632,N_4908,N_2486);
and U6633 (N_6633,N_623,N_78);
or U6634 (N_6634,N_4501,N_663);
nand U6635 (N_6635,N_1469,N_1250);
nor U6636 (N_6636,N_139,N_4185);
nand U6637 (N_6637,N_3716,N_68);
nand U6638 (N_6638,N_4475,N_56);
and U6639 (N_6639,N_2796,N_2547);
nor U6640 (N_6640,N_2605,N_2886);
nor U6641 (N_6641,N_4853,N_758);
nor U6642 (N_6642,N_2781,N_2011);
xor U6643 (N_6643,N_3943,N_3998);
nor U6644 (N_6644,N_3406,N_607);
nand U6645 (N_6645,N_1515,N_3500);
and U6646 (N_6646,N_3453,N_2510);
nand U6647 (N_6647,N_2983,N_2941);
and U6648 (N_6648,N_4262,N_216);
or U6649 (N_6649,N_2402,N_3024);
or U6650 (N_6650,N_4351,N_4201);
nor U6651 (N_6651,N_1053,N_2545);
nand U6652 (N_6652,N_3997,N_474);
nand U6653 (N_6653,N_59,N_2014);
nand U6654 (N_6654,N_4442,N_4731);
nor U6655 (N_6655,N_3286,N_2279);
nand U6656 (N_6656,N_4199,N_1051);
nand U6657 (N_6657,N_3852,N_4033);
nand U6658 (N_6658,N_3738,N_2962);
nand U6659 (N_6659,N_98,N_1389);
nor U6660 (N_6660,N_3313,N_229);
and U6661 (N_6661,N_66,N_2088);
nand U6662 (N_6662,N_3163,N_4111);
and U6663 (N_6663,N_831,N_449);
nor U6664 (N_6664,N_4841,N_4301);
or U6665 (N_6665,N_1802,N_1107);
nor U6666 (N_6666,N_512,N_1098);
nor U6667 (N_6667,N_2843,N_535);
nor U6668 (N_6668,N_2183,N_1216);
and U6669 (N_6669,N_2508,N_2850);
and U6670 (N_6670,N_1570,N_1003);
or U6671 (N_6671,N_149,N_864);
and U6672 (N_6672,N_3606,N_3532);
nand U6673 (N_6673,N_2730,N_4189);
xor U6674 (N_6674,N_4914,N_4822);
nor U6675 (N_6675,N_1988,N_4653);
or U6676 (N_6676,N_4002,N_713);
nor U6677 (N_6677,N_4319,N_3416);
and U6678 (N_6678,N_2674,N_1060);
nor U6679 (N_6679,N_196,N_1194);
nand U6680 (N_6680,N_1085,N_4377);
xnor U6681 (N_6681,N_1438,N_2144);
and U6682 (N_6682,N_4742,N_4771);
and U6683 (N_6683,N_1214,N_3874);
nand U6684 (N_6684,N_2787,N_2593);
nand U6685 (N_6685,N_973,N_195);
nor U6686 (N_6686,N_4077,N_4783);
and U6687 (N_6687,N_1440,N_4153);
or U6688 (N_6688,N_4414,N_4745);
nand U6689 (N_6689,N_22,N_245);
nand U6690 (N_6690,N_1755,N_3663);
and U6691 (N_6691,N_2497,N_682);
or U6692 (N_6692,N_2573,N_3395);
or U6693 (N_6693,N_3662,N_4837);
and U6694 (N_6694,N_395,N_1861);
xnor U6695 (N_6695,N_3323,N_3116);
nor U6696 (N_6696,N_3124,N_4776);
or U6697 (N_6697,N_3497,N_1008);
nor U6698 (N_6698,N_3973,N_3684);
nand U6699 (N_6699,N_1963,N_945);
xor U6700 (N_6700,N_1901,N_26);
nand U6701 (N_6701,N_1102,N_625);
nor U6702 (N_6702,N_716,N_4962);
xnor U6703 (N_6703,N_3250,N_2238);
nand U6704 (N_6704,N_4580,N_1103);
xor U6705 (N_6705,N_3614,N_601);
nand U6706 (N_6706,N_483,N_2295);
or U6707 (N_6707,N_2043,N_462);
and U6708 (N_6708,N_4587,N_1145);
or U6709 (N_6709,N_2756,N_4985);
nand U6710 (N_6710,N_2755,N_2895);
nor U6711 (N_6711,N_4756,N_2339);
and U6712 (N_6712,N_438,N_2309);
or U6713 (N_6713,N_1871,N_2563);
and U6714 (N_6714,N_1892,N_2953);
nor U6715 (N_6715,N_4267,N_4084);
nand U6716 (N_6716,N_4014,N_1078);
or U6717 (N_6717,N_1597,N_839);
nor U6718 (N_6718,N_3798,N_356);
nor U6719 (N_6719,N_3681,N_3868);
nand U6720 (N_6720,N_2580,N_4530);
or U6721 (N_6721,N_2872,N_4463);
nor U6722 (N_6722,N_1576,N_516);
or U6723 (N_6723,N_1912,N_39);
nand U6724 (N_6724,N_2817,N_1242);
or U6725 (N_6725,N_3725,N_208);
and U6726 (N_6726,N_676,N_1001);
nand U6727 (N_6727,N_1784,N_4550);
or U6728 (N_6728,N_7,N_706);
or U6729 (N_6729,N_964,N_4975);
nand U6730 (N_6730,N_132,N_3408);
nor U6731 (N_6731,N_301,N_2152);
nand U6732 (N_6732,N_2991,N_2765);
nor U6733 (N_6733,N_3477,N_1437);
and U6734 (N_6734,N_4629,N_378);
nor U6735 (N_6735,N_539,N_1919);
nand U6736 (N_6736,N_1790,N_2098);
or U6737 (N_6737,N_2301,N_738);
nand U6738 (N_6738,N_2978,N_656);
nand U6739 (N_6739,N_1167,N_4835);
nor U6740 (N_6740,N_912,N_3502);
and U6741 (N_6741,N_3791,N_3961);
nand U6742 (N_6742,N_4006,N_2479);
nor U6743 (N_6743,N_3579,N_92);
and U6744 (N_6744,N_3055,N_2094);
and U6745 (N_6745,N_1356,N_1363);
nand U6746 (N_6746,N_4697,N_2902);
xor U6747 (N_6747,N_1317,N_426);
nand U6748 (N_6748,N_406,N_188);
nand U6749 (N_6749,N_4269,N_209);
nand U6750 (N_6750,N_1628,N_3654);
and U6751 (N_6751,N_639,N_63);
nand U6752 (N_6752,N_3911,N_2965);
nand U6753 (N_6753,N_2500,N_4148);
and U6754 (N_6754,N_2782,N_2371);
and U6755 (N_6755,N_1712,N_178);
nor U6756 (N_6756,N_4499,N_3708);
and U6757 (N_6757,N_4778,N_2598);
or U6758 (N_6758,N_4105,N_493);
and U6759 (N_6759,N_37,N_3472);
nand U6760 (N_6760,N_3399,N_636);
nor U6761 (N_6761,N_3879,N_3702);
nor U6762 (N_6762,N_1603,N_1384);
nand U6763 (N_6763,N_701,N_3864);
xor U6764 (N_6764,N_1809,N_4157);
or U6765 (N_6765,N_4458,N_79);
and U6766 (N_6766,N_1804,N_40);
and U6767 (N_6767,N_2036,N_1775);
and U6768 (N_6768,N_2209,N_677);
nor U6769 (N_6769,N_1608,N_1616);
and U6770 (N_6770,N_4233,N_1966);
and U6771 (N_6771,N_1970,N_2625);
and U6772 (N_6772,N_2018,N_715);
or U6773 (N_6773,N_1857,N_1958);
or U6774 (N_6774,N_2214,N_2745);
nand U6775 (N_6775,N_1365,N_1018);
nor U6776 (N_6776,N_4445,N_3949);
and U6777 (N_6777,N_1040,N_2783);
or U6778 (N_6778,N_4315,N_4041);
nor U6779 (N_6779,N_4055,N_909);
and U6780 (N_6780,N_3504,N_4709);
and U6781 (N_6781,N_3131,N_1243);
and U6782 (N_6782,N_1893,N_136);
and U6783 (N_6783,N_1262,N_731);
nand U6784 (N_6784,N_4817,N_2922);
and U6785 (N_6785,N_1344,N_154);
nor U6786 (N_6786,N_3312,N_2794);
and U6787 (N_6787,N_596,N_1783);
nor U6788 (N_6788,N_751,N_1718);
nand U6789 (N_6789,N_4258,N_4791);
nor U6790 (N_6790,N_2220,N_3407);
nor U6791 (N_6791,N_3519,N_2993);
nor U6792 (N_6792,N_4184,N_3333);
and U6793 (N_6793,N_315,N_1668);
or U6794 (N_6794,N_4640,N_3272);
nor U6795 (N_6795,N_2588,N_1173);
and U6796 (N_6796,N_358,N_2241);
nand U6797 (N_6797,N_1835,N_1094);
nand U6798 (N_6798,N_1154,N_1444);
nand U6799 (N_6799,N_869,N_3698);
nor U6800 (N_6800,N_4730,N_732);
and U6801 (N_6801,N_2083,N_547);
or U6802 (N_6802,N_2125,N_3835);
and U6803 (N_6803,N_752,N_3607);
xor U6804 (N_6804,N_2069,N_3363);
nand U6805 (N_6805,N_3240,N_1408);
and U6806 (N_6806,N_4008,N_4059);
or U6807 (N_6807,N_1702,N_2696);
or U6808 (N_6808,N_811,N_4172);
nor U6809 (N_6809,N_3731,N_2540);
and U6810 (N_6810,N_104,N_4196);
nor U6811 (N_6811,N_1268,N_450);
and U6812 (N_6812,N_3855,N_582);
nand U6813 (N_6813,N_2200,N_1760);
and U6814 (N_6814,N_2478,N_633);
or U6815 (N_6815,N_240,N_1541);
nand U6816 (N_6816,N_2949,N_4710);
or U6817 (N_6817,N_3710,N_1213);
or U6818 (N_6818,N_3060,N_2323);
nor U6819 (N_6819,N_4855,N_975);
nand U6820 (N_6820,N_2458,N_3963);
and U6821 (N_6821,N_3690,N_412);
nor U6822 (N_6822,N_4904,N_4493);
or U6823 (N_6823,N_4238,N_2688);
nor U6824 (N_6824,N_4323,N_3165);
nand U6825 (N_6825,N_135,N_4890);
and U6826 (N_6826,N_1588,N_481);
nand U6827 (N_6827,N_4409,N_1903);
or U6828 (N_6828,N_1491,N_1483);
or U6829 (N_6829,N_1,N_4032);
and U6830 (N_6830,N_2558,N_2060);
nand U6831 (N_6831,N_3858,N_3726);
nor U6832 (N_6832,N_702,N_4197);
nand U6833 (N_6833,N_3249,N_1524);
or U6834 (N_6834,N_4343,N_4380);
nor U6835 (N_6835,N_159,N_458);
nor U6836 (N_6836,N_1698,N_1447);
nor U6837 (N_6837,N_1613,N_533);
or U6838 (N_6838,N_125,N_1744);
nand U6839 (N_6839,N_951,N_812);
nor U6840 (N_6840,N_4647,N_4970);
nand U6841 (N_6841,N_2022,N_2506);
and U6842 (N_6842,N_1261,N_3636);
and U6843 (N_6843,N_2608,N_4551);
and U6844 (N_6844,N_687,N_572);
or U6845 (N_6845,N_2665,N_4035);
nor U6846 (N_6846,N_160,N_3390);
nor U6847 (N_6847,N_4931,N_3283);
and U6848 (N_6848,N_806,N_4373);
and U6849 (N_6849,N_1946,N_517);
nand U6850 (N_6850,N_27,N_4346);
nand U6851 (N_6851,N_3935,N_3219);
and U6852 (N_6852,N_4416,N_122);
or U6853 (N_6853,N_2551,N_1424);
or U6854 (N_6854,N_3980,N_1184);
or U6855 (N_6855,N_4273,N_4542);
and U6856 (N_6856,N_1358,N_3469);
and U6857 (N_6857,N_4069,N_809);
and U6858 (N_6858,N_4718,N_3037);
nor U6859 (N_6859,N_1560,N_3422);
nand U6860 (N_6860,N_1693,N_1600);
or U6861 (N_6861,N_1017,N_727);
nor U6862 (N_6862,N_2213,N_2897);
xor U6863 (N_6863,N_3062,N_3188);
and U6864 (N_6864,N_2492,N_2620);
or U6865 (N_6865,N_1694,N_142);
and U6866 (N_6866,N_1406,N_3638);
nor U6867 (N_6867,N_2233,N_4093);
nand U6868 (N_6868,N_4856,N_2934);
and U6869 (N_6869,N_3490,N_4673);
and U6870 (N_6870,N_1232,N_1907);
nand U6871 (N_6871,N_4186,N_2576);
or U6872 (N_6872,N_1277,N_3865);
and U6873 (N_6873,N_4000,N_882);
nand U6874 (N_6874,N_1665,N_3158);
and U6875 (N_6875,N_2772,N_3760);
or U6876 (N_6876,N_4439,N_4910);
nand U6877 (N_6877,N_3734,N_852);
nor U6878 (N_6878,N_2948,N_4963);
and U6879 (N_6879,N_1631,N_381);
xor U6880 (N_6880,N_2808,N_3974);
nand U6881 (N_6881,N_1360,N_1274);
nand U6882 (N_6882,N_4193,N_4234);
and U6883 (N_6883,N_957,N_2766);
nand U6884 (N_6884,N_1552,N_3685);
nor U6885 (N_6885,N_4572,N_3604);
or U6886 (N_6886,N_1468,N_802);
nor U6887 (N_6887,N_3183,N_3380);
nor U6888 (N_6888,N_3140,N_970);
nand U6889 (N_6889,N_4283,N_2026);
and U6890 (N_6890,N_2693,N_4379);
nand U6891 (N_6891,N_3644,N_3357);
nor U6892 (N_6892,N_1558,N_2753);
and U6893 (N_6893,N_1119,N_3328);
xnor U6894 (N_6894,N_3653,N_2821);
nor U6895 (N_6895,N_1811,N_700);
and U6896 (N_6896,N_745,N_2655);
nand U6897 (N_6897,N_2495,N_1265);
xnor U6898 (N_6898,N_3633,N_250);
or U6899 (N_6899,N_2470,N_4826);
nand U6900 (N_6900,N_297,N_903);
or U6901 (N_6901,N_4737,N_476);
nand U6902 (N_6902,N_4764,N_3805);
nor U6903 (N_6903,N_3393,N_4187);
nand U6904 (N_6904,N_1993,N_4169);
or U6905 (N_6905,N_4358,N_94);
nand U6906 (N_6906,N_1516,N_4329);
and U6907 (N_6907,N_1624,N_4628);
xor U6908 (N_6908,N_3968,N_4165);
nand U6909 (N_6909,N_4583,N_3227);
or U6910 (N_6910,N_4978,N_1581);
or U6911 (N_6911,N_1991,N_2865);
nand U6912 (N_6912,N_2887,N_2805);
or U6913 (N_6913,N_279,N_3635);
or U6914 (N_6914,N_3189,N_2224);
nand U6915 (N_6915,N_51,N_4562);
and U6916 (N_6916,N_3211,N_911);
nor U6917 (N_6917,N_953,N_3699);
nand U6918 (N_6918,N_3210,N_941);
nor U6919 (N_6919,N_3035,N_3149);
and U6920 (N_6920,N_1959,N_1128);
nor U6921 (N_6921,N_3185,N_333);
xnor U6922 (N_6922,N_4049,N_4448);
or U6923 (N_6923,N_3881,N_1655);
nor U6924 (N_6924,N_544,N_3285);
nand U6925 (N_6925,N_1304,N_65);
and U6926 (N_6926,N_3298,N_261);
nor U6927 (N_6927,N_4354,N_206);
nand U6928 (N_6928,N_1532,N_4704);
and U6929 (N_6929,N_342,N_3028);
nor U6930 (N_6930,N_1224,N_3434);
nor U6931 (N_6931,N_4386,N_1392);
and U6932 (N_6932,N_2136,N_2156);
and U6933 (N_6933,N_2221,N_563);
nand U6934 (N_6934,N_1248,N_4605);
or U6935 (N_6935,N_1276,N_2972);
nand U6936 (N_6936,N_561,N_1948);
or U6937 (N_6937,N_28,N_2317);
xor U6938 (N_6938,N_4941,N_1943);
or U6939 (N_6939,N_4478,N_2530);
and U6940 (N_6940,N_1593,N_3942);
or U6941 (N_6941,N_2607,N_86);
and U6942 (N_6942,N_749,N_665);
nor U6943 (N_6943,N_469,N_907);
and U6944 (N_6944,N_69,N_2831);
and U6945 (N_6945,N_1266,N_276);
and U6946 (N_6946,N_4669,N_1582);
or U6947 (N_6947,N_1757,N_1199);
and U6948 (N_6948,N_1226,N_2239);
and U6949 (N_6949,N_3788,N_4973);
and U6950 (N_6950,N_3938,N_1596);
nor U6951 (N_6951,N_1283,N_3610);
xor U6952 (N_6952,N_1748,N_4733);
nand U6953 (N_6953,N_1256,N_4794);
and U6954 (N_6954,N_2691,N_3105);
nand U6955 (N_6955,N_4851,N_267);
nand U6956 (N_6956,N_2657,N_2269);
nand U6957 (N_6957,N_1537,N_3077);
nor U6958 (N_6958,N_2119,N_2355);
nor U6959 (N_6959,N_1832,N_748);
nand U6960 (N_6960,N_3554,N_1848);
and U6961 (N_6961,N_3896,N_1212);
and U6962 (N_6962,N_4300,N_2871);
xnor U6963 (N_6963,N_2020,N_860);
nand U6964 (N_6964,N_3807,N_1817);
and U6965 (N_6965,N_4370,N_2005);
nand U6966 (N_6966,N_4884,N_3135);
nand U6967 (N_6967,N_2435,N_1830);
or U6968 (N_6968,N_2462,N_1157);
nand U6969 (N_6969,N_176,N_4849);
or U6970 (N_6970,N_771,N_688);
nor U6971 (N_6971,N_3921,N_659);
nand U6972 (N_6972,N_2952,N_2863);
or U6973 (N_6973,N_1292,N_4644);
nor U6974 (N_6974,N_3316,N_1117);
nor U6975 (N_6975,N_3836,N_310);
or U6976 (N_6976,N_1099,N_1061);
and U6977 (N_6977,N_306,N_718);
nor U6978 (N_6978,N_1579,N_1584);
and U6979 (N_6979,N_761,N_553);
nor U6980 (N_6980,N_3727,N_3027);
nand U6981 (N_6981,N_1296,N_1962);
and U6982 (N_6982,N_609,N_225);
or U6983 (N_6983,N_4632,N_537);
and U6984 (N_6984,N_2265,N_1820);
nand U6985 (N_6985,N_2954,N_4781);
or U6986 (N_6986,N_241,N_4264);
nor U6987 (N_6987,N_4053,N_4068);
nand U6988 (N_6988,N_2675,N_4054);
nor U6989 (N_6989,N_2475,N_2780);
and U6990 (N_6990,N_1644,N_1353);
or U6991 (N_6991,N_4081,N_38);
nor U6992 (N_6992,N_2105,N_3213);
or U6993 (N_6993,N_1916,N_2725);
or U6994 (N_6994,N_427,N_1160);
and U6995 (N_6995,N_3774,N_4924);
nor U6996 (N_6996,N_2845,N_1441);
nand U6997 (N_6997,N_4512,N_2225);
and U6998 (N_6998,N_1692,N_3810);
nand U6999 (N_6999,N_4421,N_3084);
xor U7000 (N_7000,N_3603,N_2439);
or U7001 (N_7001,N_3169,N_145);
nand U7002 (N_7002,N_4717,N_2111);
nand U7003 (N_7003,N_2308,N_2646);
nor U7004 (N_7004,N_2626,N_4188);
nand U7005 (N_7005,N_2262,N_1782);
nor U7006 (N_7006,N_4507,N_35);
or U7007 (N_7007,N_2716,N_4212);
nor U7008 (N_7008,N_1403,N_3280);
or U7009 (N_7009,N_3769,N_1072);
nand U7010 (N_7010,N_1228,N_2956);
or U7011 (N_7011,N_291,N_3290);
nand U7012 (N_7012,N_4813,N_3439);
nand U7013 (N_7013,N_626,N_2619);
and U7014 (N_7014,N_3403,N_4552);
and U7015 (N_7015,N_2054,N_129);
or U7016 (N_7016,N_1973,N_277);
nand U7017 (N_7017,N_1011,N_2461);
nor U7018 (N_7018,N_2273,N_4540);
nor U7019 (N_7019,N_1801,N_2393);
nand U7020 (N_7020,N_3813,N_2997);
nor U7021 (N_7021,N_80,N_1707);
and U7022 (N_7022,N_2961,N_2584);
nand U7023 (N_7023,N_4882,N_1908);
or U7024 (N_7024,N_3191,N_1267);
or U7025 (N_7025,N_1161,N_1223);
xor U7026 (N_7026,N_1779,N_2921);
nand U7027 (N_7027,N_2612,N_3962);
and U7028 (N_7028,N_1629,N_1701);
nand U7029 (N_7029,N_2670,N_349);
or U7030 (N_7030,N_1675,N_3757);
and U7031 (N_7031,N_999,N_163);
nor U7032 (N_7032,N_3011,N_3113);
or U7033 (N_7033,N_1569,N_2179);
or U7034 (N_7034,N_3082,N_249);
or U7035 (N_7035,N_3207,N_411);
and U7036 (N_7036,N_398,N_3581);
or U7037 (N_7037,N_3906,N_4943);
or U7038 (N_7038,N_2099,N_3762);
nor U7039 (N_7039,N_2289,N_573);
nor U7040 (N_7040,N_4102,N_1992);
nand U7041 (N_7041,N_131,N_3703);
and U7042 (N_7042,N_3586,N_4114);
nand U7043 (N_7043,N_34,N_3041);
and U7044 (N_7044,N_2501,N_1401);
nor U7045 (N_7045,N_4895,N_430);
and U7046 (N_7046,N_3404,N_2353);
nor U7047 (N_7047,N_508,N_4623);
or U7048 (N_7048,N_3321,N_1275);
or U7049 (N_7049,N_3258,N_3365);
nor U7050 (N_7050,N_3417,N_497);
and U7051 (N_7051,N_42,N_1818);
nand U7052 (N_7052,N_1375,N_2641);
or U7053 (N_7053,N_974,N_3817);
and U7054 (N_7054,N_3400,N_4589);
nor U7055 (N_7055,N_3302,N_3170);
nor U7056 (N_7056,N_3820,N_674);
nor U7057 (N_7057,N_2294,N_1238);
nor U7058 (N_7058,N_981,N_4200);
and U7059 (N_7059,N_4570,N_2401);
nor U7060 (N_7060,N_4883,N_18);
nand U7061 (N_7061,N_4719,N_2103);
nor U7062 (N_7062,N_4524,N_1792);
nor U7063 (N_7063,N_766,N_3839);
nor U7064 (N_7064,N_271,N_2746);
and U7065 (N_7065,N_4782,N_4120);
nand U7066 (N_7066,N_1752,N_2165);
nand U7067 (N_7067,N_3831,N_335);
or U7068 (N_7068,N_1705,N_1202);
or U7069 (N_7069,N_1510,N_1152);
nand U7070 (N_7070,N_3854,N_4809);
and U7071 (N_7071,N_1411,N_300);
xor U7072 (N_7072,N_3627,N_2008);
and U7073 (N_7073,N_4472,N_4847);
and U7074 (N_7074,N_234,N_4538);
or U7075 (N_7075,N_106,N_1659);
and U7076 (N_7076,N_1886,N_1831);
nor U7077 (N_7077,N_3007,N_1789);
and U7078 (N_7078,N_386,N_4330);
and U7079 (N_7079,N_407,N_844);
nor U7080 (N_7080,N_4555,N_4311);
nand U7081 (N_7081,N_511,N_1010);
nor U7082 (N_7082,N_2134,N_4636);
nor U7083 (N_7083,N_1846,N_1416);
nor U7084 (N_7084,N_1446,N_1316);
nor U7085 (N_7085,N_3914,N_2114);
or U7086 (N_7086,N_4692,N_4886);
nand U7087 (N_7087,N_3089,N_2433);
or U7088 (N_7088,N_2025,N_4879);
or U7089 (N_7089,N_1405,N_2370);
or U7090 (N_7090,N_4854,N_2940);
nand U7091 (N_7091,N_4208,N_2330);
nor U7092 (N_7092,N_2217,N_419);
nand U7093 (N_7093,N_1498,N_4516);
and U7094 (N_7094,N_1130,N_292);
and U7095 (N_7095,N_3557,N_4280);
nand U7096 (N_7096,N_3730,N_662);
nand U7097 (N_7097,N_4824,N_4454);
xnor U7098 (N_7098,N_2971,N_3096);
nand U7099 (N_7099,N_2274,N_3452);
or U7100 (N_7100,N_2929,N_2816);
nand U7101 (N_7101,N_2884,N_1413);
and U7102 (N_7102,N_2044,N_1526);
and U7103 (N_7103,N_81,N_1458);
and U7104 (N_7104,N_2888,N_1749);
nor U7105 (N_7105,N_725,N_203);
or U7106 (N_7106,N_2023,N_1759);
or U7107 (N_7107,N_3090,N_1336);
or U7108 (N_7108,N_264,N_4548);
and U7109 (N_7109,N_3289,N_457);
nand U7110 (N_7110,N_592,N_265);
and U7111 (N_7111,N_4576,N_4019);
and U7112 (N_7112,N_2380,N_112);
or U7113 (N_7113,N_4616,N_4796);
and U7114 (N_7114,N_4876,N_4145);
nand U7115 (N_7115,N_2663,N_1377);
nand U7116 (N_7116,N_3925,N_2851);
nand U7117 (N_7117,N_1679,N_490);
and U7118 (N_7118,N_4024,N_985);
nor U7119 (N_7119,N_4915,N_3761);
and U7120 (N_7120,N_3691,N_1108);
nor U7121 (N_7121,N_1499,N_2757);
nor U7122 (N_7122,N_2197,N_2258);
or U7123 (N_7123,N_1548,N_2834);
nand U7124 (N_7124,N_1969,N_4239);
and U7125 (N_7125,N_814,N_164);
or U7126 (N_7126,N_11,N_334);
or U7127 (N_7127,N_3651,N_96);
and U7128 (N_7128,N_1741,N_4523);
or U7129 (N_7129,N_2793,N_14);
nand U7130 (N_7130,N_1333,N_4660);
nor U7131 (N_7131,N_298,N_4597);
and U7132 (N_7132,N_123,N_4863);
nand U7133 (N_7133,N_2564,N_2622);
and U7134 (N_7134,N_4108,N_2296);
nand U7135 (N_7135,N_2659,N_3435);
or U7136 (N_7136,N_1814,N_1724);
nand U7137 (N_7137,N_3748,N_328);
nor U7138 (N_7138,N_3076,N_2356);
and U7139 (N_7139,N_1200,N_1221);
or U7140 (N_7140,N_4600,N_3172);
xor U7141 (N_7141,N_3159,N_3524);
or U7142 (N_7142,N_4017,N_4174);
or U7143 (N_7143,N_3419,N_3751);
nand U7144 (N_7144,N_1551,N_128);
xnor U7145 (N_7145,N_4099,N_4893);
nand U7146 (N_7146,N_853,N_598);
and U7147 (N_7147,N_1138,N_1249);
xnor U7148 (N_7148,N_1445,N_3021);
or U7149 (N_7149,N_3777,N_1575);
nor U7150 (N_7150,N_3465,N_2407);
or U7151 (N_7151,N_1774,N_4706);
xnor U7152 (N_7152,N_4547,N_2255);
nand U7153 (N_7153,N_1331,N_856);
nand U7154 (N_7154,N_4113,N_3268);
nand U7155 (N_7155,N_3479,N_141);
and U7156 (N_7156,N_3198,N_2650);
or U7157 (N_7157,N_2513,N_1547);
nand U7158 (N_7158,N_1402,N_3992);
nand U7159 (N_7159,N_421,N_2396);
xor U7160 (N_7160,N_2379,N_3676);
nor U7161 (N_7161,N_3032,N_574);
nand U7162 (N_7162,N_4083,N_1297);
or U7163 (N_7163,N_4728,N_5);
nand U7164 (N_7164,N_3564,N_2723);
nand U7165 (N_7165,N_660,N_273);
nand U7166 (N_7166,N_1895,N_3600);
or U7167 (N_7167,N_373,N_3383);
nor U7168 (N_7168,N_1875,N_2228);
and U7169 (N_7169,N_4793,N_499);
nor U7170 (N_7170,N_3369,N_810);
nor U7171 (N_7171,N_1689,N_1495);
or U7172 (N_7172,N_3296,N_371);
nor U7173 (N_7173,N_898,N_939);
and U7174 (N_7174,N_4844,N_25);
or U7175 (N_7175,N_4729,N_2615);
nand U7176 (N_7176,N_3464,N_3171);
and U7177 (N_7177,N_49,N_1684);
nand U7178 (N_7178,N_1489,N_461);
nor U7179 (N_7179,N_1984,N_2711);
or U7180 (N_7180,N_2386,N_778);
and U7181 (N_7181,N_920,N_569);
nor U7182 (N_7182,N_1778,N_2436);
xor U7183 (N_7183,N_3126,N_1500);
or U7184 (N_7184,N_2061,N_3446);
nand U7185 (N_7185,N_3715,N_1511);
or U7186 (N_7186,N_2193,N_621);
and U7187 (N_7187,N_4392,N_4722);
or U7188 (N_7188,N_2720,N_4126);
xnor U7189 (N_7189,N_571,N_4342);
nand U7190 (N_7190,N_173,N_1518);
and U7191 (N_7191,N_4598,N_1031);
or U7192 (N_7192,N_2417,N_3081);
nor U7193 (N_7193,N_4046,N_622);
or U7194 (N_7194,N_4242,N_1856);
nor U7195 (N_7195,N_3705,N_4356);
or U7196 (N_7196,N_4437,N_1567);
and U7197 (N_7197,N_4850,N_943);
and U7198 (N_7198,N_3670,N_4136);
and U7199 (N_7199,N_3396,N_2409);
nor U7200 (N_7200,N_2857,N_4780);
or U7201 (N_7201,N_1193,N_464);
nor U7202 (N_7202,N_3072,N_4909);
nand U7203 (N_7203,N_4446,N_1298);
or U7204 (N_7204,N_1041,N_3175);
and U7205 (N_7205,N_3779,N_892);
nand U7206 (N_7206,N_2248,N_4403);
and U7207 (N_7207,N_46,N_4913);
nor U7208 (N_7208,N_2810,N_1587);
nand U7209 (N_7209,N_2081,N_4869);
and U7210 (N_7210,N_3260,N_3347);
or U7211 (N_7211,N_910,N_4515);
or U7212 (N_7212,N_2767,N_3907);
or U7213 (N_7213,N_2332,N_1851);
nand U7214 (N_7214,N_3668,N_4549);
or U7215 (N_7215,N_3672,N_2909);
nand U7216 (N_7216,N_1074,N_1410);
nand U7217 (N_7217,N_1247,N_1968);
nor U7218 (N_7218,N_2460,N_3723);
nor U7219 (N_7219,N_181,N_222);
nand U7220 (N_7220,N_3437,N_1112);
and U7221 (N_7221,N_3877,N_1472);
or U7222 (N_7222,N_2685,N_4455);
nand U7223 (N_7223,N_3223,N_3537);
nor U7224 (N_7224,N_3749,N_3850);
or U7225 (N_7225,N_3092,N_4621);
and U7226 (N_7226,N_3993,N_1097);
and U7227 (N_7227,N_2703,N_4427);
and U7228 (N_7228,N_4792,N_1016);
or U7229 (N_7229,N_2819,N_4878);
xnor U7230 (N_7230,N_3117,N_4618);
or U7231 (N_7231,N_648,N_1642);
nand U7232 (N_7232,N_4546,N_2494);
nor U7233 (N_7233,N_805,N_2708);
or U7234 (N_7234,N_3029,N_3722);
nor U7235 (N_7235,N_2469,N_4397);
or U7236 (N_7236,N_3958,N_3287);
nor U7237 (N_7237,N_2524,N_4982);
and U7238 (N_7238,N_591,N_1833);
nand U7239 (N_7239,N_4062,N_3078);
xnor U7240 (N_7240,N_3015,N_4763);
nand U7241 (N_7241,N_1766,N_4082);
nand U7242 (N_7242,N_4318,N_707);
nor U7243 (N_7243,N_4595,N_1897);
and U7244 (N_7244,N_3764,N_1839);
nand U7245 (N_7245,N_1355,N_3356);
and U7246 (N_7246,N_1932,N_4001);
nor U7247 (N_7247,N_2126,N_4314);
nand U7248 (N_7248,N_3823,N_3305);
and U7249 (N_7249,N_3775,N_4218);
and U7250 (N_7250,N_4489,N_4491);
and U7251 (N_7251,N_1254,N_793);
or U7252 (N_7252,N_3849,N_4859);
and U7253 (N_7253,N_1230,N_4871);
nand U7254 (N_7254,N_2849,N_1554);
nor U7255 (N_7255,N_151,N_3256);
nor U7256 (N_7256,N_4374,N_2154);
nor U7257 (N_7257,N_4857,N_2071);
nor U7258 (N_7258,N_302,N_4662);
and U7259 (N_7259,N_3999,N_2534);
or U7260 (N_7260,N_2955,N_3409);
or U7261 (N_7261,N_2351,N_4247);
or U7262 (N_7262,N_3039,N_239);
and U7263 (N_7263,N_2482,N_466);
and U7264 (N_7264,N_231,N_4043);
nand U7265 (N_7265,N_475,N_3180);
or U7266 (N_7266,N_3338,N_3134);
and U7267 (N_7267,N_2290,N_2490);
nand U7268 (N_7268,N_620,N_2493);
nor U7269 (N_7269,N_1734,N_4716);
or U7270 (N_7270,N_3075,N_4749);
nor U7271 (N_7271,N_3359,N_3097);
nor U7272 (N_7272,N_4248,N_2376);
and U7273 (N_7273,N_16,N_3432);
nor U7274 (N_7274,N_1271,N_3602);
nor U7275 (N_7275,N_4183,N_2187);
or U7276 (N_7276,N_1455,N_4214);
and U7277 (N_7277,N_3288,N_976);
nor U7278 (N_7278,N_4614,N_3666);
and U7279 (N_7279,N_2480,N_1854);
nand U7280 (N_7280,N_1162,N_1746);
nand U7281 (N_7281,N_833,N_3217);
nand U7282 (N_7282,N_2728,N_260);
and U7283 (N_7283,N_4252,N_3193);
nor U7284 (N_7284,N_1955,N_288);
nand U7285 (N_7285,N_1688,N_257);
nor U7286 (N_7286,N_4,N_764);
nor U7287 (N_7287,N_4740,N_3345);
nor U7288 (N_7288,N_3344,N_1366);
nand U7289 (N_7289,N_1742,N_4256);
or U7290 (N_7290,N_531,N_4990);
nor U7291 (N_7291,N_3100,N_4625);
or U7292 (N_7292,N_4152,N_3274);
or U7293 (N_7293,N_2428,N_3667);
or U7294 (N_7294,N_1709,N_2257);
nor U7295 (N_7295,N_1555,N_4766);
and U7296 (N_7296,N_1680,N_594);
nand U7297 (N_7297,N_3120,N_191);
or U7298 (N_7298,N_1151,N_1914);
and U7299 (N_7299,N_1357,N_1837);
and U7300 (N_7300,N_278,N_960);
and U7301 (N_7301,N_3583,N_2532);
nor U7302 (N_7302,N_1387,N_1179);
nor U7303 (N_7303,N_4341,N_4118);
xnor U7304 (N_7304,N_1434,N_1937);
and U7305 (N_7305,N_3689,N_588);
nor U7306 (N_7306,N_3496,N_3753);
and U7307 (N_7307,N_3936,N_3818);
or U7308 (N_7308,N_3516,N_4541);
nand U7309 (N_7309,N_4953,N_67);
nand U7310 (N_7310,N_2762,N_4496);
nor U7311 (N_7311,N_542,N_2282);
and U7312 (N_7312,N_2566,N_2562);
or U7313 (N_7313,N_4668,N_3694);
nor U7314 (N_7314,N_2383,N_4180);
or U7315 (N_7315,N_4338,N_218);
nor U7316 (N_7316,N_4012,N_2468);
and U7317 (N_7317,N_1150,N_4250);
nand U7318 (N_7318,N_2638,N_4779);
nand U7319 (N_7319,N_3155,N_2944);
nor U7320 (N_7320,N_2976,N_1494);
and U7321 (N_7321,N_895,N_1654);
nor U7322 (N_7322,N_2051,N_186);
xor U7323 (N_7323,N_2203,N_4935);
nor U7324 (N_7324,N_1997,N_4721);
or U7325 (N_7325,N_1936,N_654);
nand U7326 (N_7326,N_2077,N_1750);
xor U7327 (N_7327,N_3057,N_4777);
nor U7328 (N_7328,N_2826,N_2281);
nand U7329 (N_7329,N_836,N_2666);
or U7330 (N_7330,N_3763,N_3545);
nand U7331 (N_7331,N_739,N_2198);
and U7332 (N_7332,N_3475,N_717);
or U7333 (N_7333,N_2440,N_614);
or U7334 (N_7334,N_4094,N_2306);
nor U7335 (N_7335,N_4243,N_4378);
nor U7336 (N_7336,N_1928,N_4156);
or U7337 (N_7337,N_4460,N_4860);
nor U7338 (N_7338,N_3838,N_213);
and U7339 (N_7339,N_2599,N_3947);
and U7340 (N_7340,N_4410,N_3358);
nor U7341 (N_7341,N_979,N_2662);
nor U7342 (N_7342,N_3031,N_2312);
nor U7343 (N_7343,N_2,N_2191);
nand U7344 (N_7344,N_2559,N_4047);
nand U7345 (N_7345,N_3160,N_2705);
xor U7346 (N_7346,N_875,N_4112);
nand U7347 (N_7347,N_1409,N_2867);
nor U7348 (N_7348,N_1425,N_2503);
nor U7349 (N_7349,N_3567,N_4590);
nor U7350 (N_7350,N_194,N_3098);
nor U7351 (N_7351,N_1572,N_61);
or U7352 (N_7352,N_2738,N_2324);
nor U7353 (N_7353,N_3182,N_3514);
nor U7354 (N_7354,N_1924,N_1747);
nand U7355 (N_7355,N_3601,N_3297);
and U7356 (N_7356,N_679,N_359);
nor U7357 (N_7357,N_2181,N_4150);
nand U7358 (N_7358,N_2340,N_4637);
and U7359 (N_7359,N_2150,N_4727);
and U7360 (N_7360,N_4387,N_211);
nor U7361 (N_7361,N_2082,N_330);
nor U7362 (N_7362,N_3326,N_370);
and U7363 (N_7363,N_2811,N_4867);
and U7364 (N_7364,N_4399,N_318);
nand U7365 (N_7365,N_4176,N_1324);
nor U7366 (N_7366,N_2673,N_4984);
or U7367 (N_7367,N_3145,N_423);
nand U7368 (N_7368,N_2445,N_2754);
or U7369 (N_7369,N_4057,N_2031);
xor U7370 (N_7370,N_783,N_174);
or U7371 (N_7371,N_2654,N_4312);
nand U7372 (N_7372,N_2695,N_4241);
nor U7373 (N_7373,N_728,N_4762);
nand U7374 (N_7374,N_1417,N_3361);
or U7375 (N_7375,N_526,N_4361);
nor U7376 (N_7376,N_473,N_1289);
and U7377 (N_7377,N_1088,N_2966);
nand U7378 (N_7378,N_1121,N_857);
or U7379 (N_7379,N_1123,N_4769);
and U7380 (N_7380,N_21,N_1462);
or U7381 (N_7381,N_1890,N_233);
nor U7382 (N_7382,N_742,N_899);
and U7383 (N_7383,N_3004,N_2706);
and U7384 (N_7384,N_36,N_2522);
and U7385 (N_7385,N_221,N_2347);
nor U7386 (N_7386,N_4746,N_3353);
nor U7387 (N_7387,N_1153,N_4474);
nor U7388 (N_7388,N_4964,N_4088);
and U7389 (N_7389,N_2788,N_4021);
nor U7390 (N_7390,N_3040,N_95);
or U7391 (N_7391,N_2397,N_3657);
nand U7392 (N_7392,N_1947,N_1156);
and U7393 (N_7393,N_1813,N_4654);
and U7394 (N_7394,N_4396,N_2142);
or U7395 (N_7395,N_3064,N_966);
nand U7396 (N_7396,N_832,N_3750);
and U7397 (N_7397,N_3102,N_1127);
or U7398 (N_7398,N_4178,N_2525);
nor U7399 (N_7399,N_1270,N_1240);
or U7400 (N_7400,N_3884,N_3278);
or U7401 (N_7401,N_3952,N_2354);
nor U7402 (N_7402,N_4417,N_3988);
and U7403 (N_7403,N_465,N_4337);
nand U7404 (N_7404,N_4839,N_3080);
or U7405 (N_7405,N_587,N_2639);
or U7406 (N_7406,N_1209,N_3038);
and U7407 (N_7407,N_4498,N_3900);
nor U7408 (N_7408,N_3034,N_2777);
or U7409 (N_7409,N_3837,N_4720);
or U7410 (N_7410,N_4967,N_737);
nor U7411 (N_7411,N_3487,N_3362);
nand U7412 (N_7412,N_968,N_3294);
nor U7413 (N_7413,N_1082,N_4375);
nand U7414 (N_7414,N_3522,N_1940);
or U7415 (N_7415,N_4368,N_1140);
or U7416 (N_7416,N_2305,N_4404);
nor U7417 (N_7417,N_446,N_3897);
and U7418 (N_7418,N_2100,N_201);
and U7419 (N_7419,N_285,N_2352);
nand U7420 (N_7420,N_2830,N_2368);
nor U7421 (N_7421,N_4560,N_3521);
nor U7422 (N_7422,N_4473,N_3056);
nor U7423 (N_7423,N_453,N_2905);
and U7424 (N_7424,N_1478,N_1512);
or U7425 (N_7425,N_2862,N_3320);
nand U7426 (N_7426,N_459,N_165);
nand U7427 (N_7427,N_3605,N_4131);
nand U7428 (N_7428,N_3309,N_3883);
nand U7429 (N_7429,N_4818,N_3687);
nor U7430 (N_7430,N_304,N_2697);
nand U7431 (N_7431,N_983,N_1380);
or U7432 (N_7432,N_3637,N_1926);
nand U7433 (N_7433,N_3147,N_2818);
and U7434 (N_7434,N_528,N_1258);
nor U7435 (N_7435,N_4761,N_3085);
nand U7436 (N_7436,N_4259,N_3202);
and U7437 (N_7437,N_3016,N_3454);
nand U7438 (N_7438,N_3103,N_2202);
nor U7439 (N_7439,N_2735,N_105);
nor U7440 (N_7440,N_3226,N_813);
and U7441 (N_7441,N_3177,N_313);
nor U7442 (N_7442,N_2975,N_1203);
or U7443 (N_7443,N_868,N_4149);
nor U7444 (N_7444,N_3656,N_4383);
nand U7445 (N_7445,N_121,N_1840);
or U7446 (N_7446,N_1609,N_2763);
or U7447 (N_7447,N_862,N_835);
xnor U7448 (N_7448,N_1564,N_2138);
and U7449 (N_7449,N_1507,N_2514);
nand U7450 (N_7450,N_4645,N_1143);
or U7451 (N_7451,N_2748,N_372);
nor U7452 (N_7452,N_103,N_4665);
nor U7453 (N_7453,N_629,N_935);
nor U7454 (N_7454,N_1376,N_1343);
nor U7455 (N_7455,N_1035,N_2028);
nand U7456 (N_7456,N_4173,N_615);
nor U7457 (N_7457,N_1359,N_4663);
nand U7458 (N_7458,N_269,N_4327);
nand U7459 (N_7459,N_2091,N_894);
nor U7460 (N_7460,N_2235,N_4674);
nor U7461 (N_7461,N_714,N_2173);
xor U7462 (N_7462,N_1743,N_1765);
and U7463 (N_7463,N_3844,N_4003);
or U7464 (N_7464,N_4324,N_4858);
nor U7465 (N_7465,N_2122,N_1170);
nor U7466 (N_7466,N_1132,N_4544);
nor U7467 (N_7467,N_548,N_4842);
and U7468 (N_7468,N_432,N_541);
nor U7469 (N_7469,N_4789,N_1862);
nor U7470 (N_7470,N_3630,N_2715);
nand U7471 (N_7471,N_616,N_2456);
and U7472 (N_7472,N_2348,N_4831);
or U7473 (N_7473,N_1330,N_2698);
and U7474 (N_7474,N_4559,N_3590);
nor U7475 (N_7475,N_4912,N_2836);
nor U7476 (N_7476,N_3688,N_595);
or U7477 (N_7477,N_4767,N_3965);
xor U7478 (N_7478,N_2739,N_3915);
and U7479 (N_7479,N_3000,N_4999);
or U7480 (N_7480,N_2926,N_3940);
nand U7481 (N_7481,N_3233,N_1361);
nand U7482 (N_7482,N_4519,N_3184);
xnor U7483 (N_7483,N_365,N_3366);
nor U7484 (N_7484,N_2271,N_1453);
and U7485 (N_7485,N_1738,N_198);
or U7486 (N_7486,N_924,N_3346);
and U7487 (N_7487,N_3200,N_1585);
or U7488 (N_7488,N_3693,N_2806);
or U7489 (N_7489,N_487,N_255);
nor U7490 (N_7490,N_949,N_3706);
or U7491 (N_7491,N_2543,N_2959);
or U7492 (N_7492,N_2346,N_2624);
nor U7493 (N_7493,N_4090,N_1306);
and U7494 (N_7494,N_4297,N_2614);
and U7495 (N_7495,N_2611,N_2538);
nor U7496 (N_7496,N_126,N_4302);
and U7497 (N_7497,N_2773,N_1902);
or U7498 (N_7498,N_4899,N_3856);
and U7499 (N_7499,N_4317,N_3978);
nor U7500 (N_7500,N_1454,N_3433);
nand U7501 (N_7501,N_4924,N_624);
nand U7502 (N_7502,N_3490,N_3237);
or U7503 (N_7503,N_3945,N_4408);
nand U7504 (N_7504,N_1189,N_2650);
nand U7505 (N_7505,N_3039,N_3149);
nor U7506 (N_7506,N_3475,N_2010);
nand U7507 (N_7507,N_152,N_1278);
and U7508 (N_7508,N_609,N_1390);
nand U7509 (N_7509,N_395,N_3694);
or U7510 (N_7510,N_1687,N_1371);
nor U7511 (N_7511,N_3106,N_2805);
nor U7512 (N_7512,N_2210,N_1169);
or U7513 (N_7513,N_1043,N_4274);
or U7514 (N_7514,N_2150,N_4186);
and U7515 (N_7515,N_1393,N_3809);
nand U7516 (N_7516,N_1196,N_2513);
xnor U7517 (N_7517,N_1379,N_765);
nor U7518 (N_7518,N_3841,N_3917);
and U7519 (N_7519,N_2087,N_901);
nor U7520 (N_7520,N_4713,N_1712);
nand U7521 (N_7521,N_2460,N_624);
or U7522 (N_7522,N_1100,N_1789);
nor U7523 (N_7523,N_609,N_319);
and U7524 (N_7524,N_1436,N_855);
nand U7525 (N_7525,N_815,N_4465);
and U7526 (N_7526,N_4542,N_4815);
nor U7527 (N_7527,N_1434,N_2988);
nor U7528 (N_7528,N_3972,N_4744);
xnor U7529 (N_7529,N_3888,N_3516);
nand U7530 (N_7530,N_554,N_4409);
or U7531 (N_7531,N_3287,N_949);
nand U7532 (N_7532,N_3431,N_4114);
nand U7533 (N_7533,N_521,N_379);
nor U7534 (N_7534,N_4599,N_1818);
nor U7535 (N_7535,N_1978,N_4334);
and U7536 (N_7536,N_1308,N_1454);
and U7537 (N_7537,N_1818,N_2117);
or U7538 (N_7538,N_4814,N_2624);
nand U7539 (N_7539,N_1014,N_2281);
nand U7540 (N_7540,N_1151,N_770);
or U7541 (N_7541,N_1996,N_3241);
nor U7542 (N_7542,N_1573,N_4570);
nor U7543 (N_7543,N_4745,N_932);
or U7544 (N_7544,N_3768,N_4796);
nand U7545 (N_7545,N_506,N_1223);
or U7546 (N_7546,N_3249,N_1424);
nor U7547 (N_7547,N_4418,N_2112);
and U7548 (N_7548,N_3317,N_2819);
nor U7549 (N_7549,N_469,N_2063);
or U7550 (N_7550,N_2397,N_3662);
xnor U7551 (N_7551,N_4535,N_2734);
xnor U7552 (N_7552,N_1864,N_4918);
or U7553 (N_7553,N_4614,N_1215);
or U7554 (N_7554,N_1109,N_1474);
nand U7555 (N_7555,N_4406,N_1846);
nor U7556 (N_7556,N_3980,N_1216);
nor U7557 (N_7557,N_385,N_301);
nor U7558 (N_7558,N_4978,N_4385);
xnor U7559 (N_7559,N_4357,N_2971);
nor U7560 (N_7560,N_830,N_2309);
or U7561 (N_7561,N_1583,N_677);
nor U7562 (N_7562,N_4379,N_2330);
nand U7563 (N_7563,N_2110,N_456);
nor U7564 (N_7564,N_3445,N_1918);
nand U7565 (N_7565,N_3533,N_1605);
and U7566 (N_7566,N_4105,N_4524);
nor U7567 (N_7567,N_3747,N_3936);
nand U7568 (N_7568,N_1532,N_534);
nand U7569 (N_7569,N_2269,N_492);
nand U7570 (N_7570,N_706,N_544);
nand U7571 (N_7571,N_2170,N_585);
nor U7572 (N_7572,N_71,N_992);
nand U7573 (N_7573,N_519,N_4118);
nand U7574 (N_7574,N_3532,N_199);
nand U7575 (N_7575,N_3869,N_4160);
nand U7576 (N_7576,N_1156,N_779);
or U7577 (N_7577,N_444,N_4640);
nor U7578 (N_7578,N_4180,N_3382);
nor U7579 (N_7579,N_1302,N_3583);
nand U7580 (N_7580,N_3421,N_498);
nor U7581 (N_7581,N_4565,N_1757);
or U7582 (N_7582,N_2949,N_407);
nor U7583 (N_7583,N_3987,N_3185);
nor U7584 (N_7584,N_1400,N_4831);
nand U7585 (N_7585,N_474,N_2465);
xnor U7586 (N_7586,N_1597,N_2470);
nor U7587 (N_7587,N_2440,N_1204);
nor U7588 (N_7588,N_4184,N_36);
nor U7589 (N_7589,N_4249,N_21);
nor U7590 (N_7590,N_782,N_50);
xnor U7591 (N_7591,N_2635,N_616);
nor U7592 (N_7592,N_472,N_2566);
or U7593 (N_7593,N_293,N_4989);
and U7594 (N_7594,N_448,N_2710);
nor U7595 (N_7595,N_4779,N_2261);
nand U7596 (N_7596,N_3214,N_1027);
xnor U7597 (N_7597,N_2987,N_4446);
nor U7598 (N_7598,N_3890,N_3037);
nand U7599 (N_7599,N_2190,N_3509);
nand U7600 (N_7600,N_2328,N_703);
nand U7601 (N_7601,N_3842,N_1076);
or U7602 (N_7602,N_3371,N_1718);
nand U7603 (N_7603,N_4325,N_463);
and U7604 (N_7604,N_2499,N_1577);
nand U7605 (N_7605,N_2801,N_451);
or U7606 (N_7606,N_2131,N_302);
nor U7607 (N_7607,N_148,N_347);
nand U7608 (N_7608,N_2744,N_4295);
or U7609 (N_7609,N_1062,N_2122);
or U7610 (N_7610,N_2865,N_852);
nand U7611 (N_7611,N_1159,N_902);
nand U7612 (N_7612,N_966,N_4334);
and U7613 (N_7613,N_2936,N_308);
and U7614 (N_7614,N_383,N_122);
nand U7615 (N_7615,N_2848,N_4138);
nor U7616 (N_7616,N_3988,N_4085);
nor U7617 (N_7617,N_613,N_3126);
nand U7618 (N_7618,N_20,N_1134);
or U7619 (N_7619,N_4242,N_2585);
nand U7620 (N_7620,N_1694,N_4713);
or U7621 (N_7621,N_515,N_4659);
or U7622 (N_7622,N_2108,N_3995);
nand U7623 (N_7623,N_4118,N_3409);
nor U7624 (N_7624,N_769,N_655);
nor U7625 (N_7625,N_4195,N_2883);
nor U7626 (N_7626,N_4419,N_4146);
or U7627 (N_7627,N_3270,N_2392);
or U7628 (N_7628,N_3410,N_2138);
nand U7629 (N_7629,N_2883,N_2908);
nand U7630 (N_7630,N_3143,N_2451);
nor U7631 (N_7631,N_4650,N_2131);
or U7632 (N_7632,N_3174,N_2764);
nand U7633 (N_7633,N_4979,N_2320);
nand U7634 (N_7634,N_1535,N_82);
or U7635 (N_7635,N_3894,N_2602);
nand U7636 (N_7636,N_2990,N_2911);
and U7637 (N_7637,N_4279,N_845);
nor U7638 (N_7638,N_179,N_2587);
nor U7639 (N_7639,N_3900,N_4295);
xor U7640 (N_7640,N_1505,N_2554);
or U7641 (N_7641,N_2873,N_2626);
xnor U7642 (N_7642,N_940,N_3381);
and U7643 (N_7643,N_4355,N_3906);
and U7644 (N_7644,N_1400,N_680);
nand U7645 (N_7645,N_1315,N_696);
nor U7646 (N_7646,N_4053,N_2317);
nor U7647 (N_7647,N_29,N_701);
or U7648 (N_7648,N_4033,N_1877);
nor U7649 (N_7649,N_4675,N_424);
nand U7650 (N_7650,N_728,N_4172);
nand U7651 (N_7651,N_1697,N_2425);
or U7652 (N_7652,N_544,N_2642);
nand U7653 (N_7653,N_3753,N_996);
and U7654 (N_7654,N_3864,N_870);
xor U7655 (N_7655,N_4987,N_4832);
xnor U7656 (N_7656,N_4310,N_11);
nand U7657 (N_7657,N_1149,N_1860);
or U7658 (N_7658,N_4041,N_4997);
or U7659 (N_7659,N_2448,N_4012);
or U7660 (N_7660,N_4931,N_3365);
nand U7661 (N_7661,N_1630,N_749);
or U7662 (N_7662,N_3211,N_1915);
and U7663 (N_7663,N_2610,N_2478);
or U7664 (N_7664,N_2517,N_1347);
or U7665 (N_7665,N_2163,N_513);
nor U7666 (N_7666,N_2785,N_4643);
nor U7667 (N_7667,N_3275,N_3822);
nand U7668 (N_7668,N_4769,N_4592);
nand U7669 (N_7669,N_2285,N_2333);
nand U7670 (N_7670,N_3530,N_3165);
or U7671 (N_7671,N_4880,N_787);
nor U7672 (N_7672,N_1260,N_1440);
nand U7673 (N_7673,N_1436,N_53);
and U7674 (N_7674,N_4246,N_1060);
xnor U7675 (N_7675,N_3596,N_475);
nor U7676 (N_7676,N_3057,N_3123);
or U7677 (N_7677,N_4606,N_1183);
or U7678 (N_7678,N_2998,N_1506);
and U7679 (N_7679,N_3006,N_761);
or U7680 (N_7680,N_544,N_153);
or U7681 (N_7681,N_1532,N_4680);
nor U7682 (N_7682,N_1761,N_3765);
and U7683 (N_7683,N_4613,N_2225);
xor U7684 (N_7684,N_2795,N_1212);
xor U7685 (N_7685,N_1146,N_1814);
or U7686 (N_7686,N_920,N_3248);
or U7687 (N_7687,N_2767,N_1852);
and U7688 (N_7688,N_1037,N_4326);
and U7689 (N_7689,N_2037,N_3269);
nor U7690 (N_7690,N_2049,N_3017);
and U7691 (N_7691,N_3042,N_132);
or U7692 (N_7692,N_539,N_1154);
or U7693 (N_7693,N_3708,N_1775);
nand U7694 (N_7694,N_4723,N_2962);
xnor U7695 (N_7695,N_1414,N_4552);
nand U7696 (N_7696,N_2964,N_1303);
nor U7697 (N_7697,N_3141,N_4509);
nand U7698 (N_7698,N_3501,N_2074);
nor U7699 (N_7699,N_934,N_940);
nand U7700 (N_7700,N_4176,N_2714);
or U7701 (N_7701,N_920,N_1887);
or U7702 (N_7702,N_4571,N_3364);
nand U7703 (N_7703,N_2409,N_233);
nor U7704 (N_7704,N_2218,N_1412);
nor U7705 (N_7705,N_1086,N_648);
nand U7706 (N_7706,N_3378,N_1537);
nand U7707 (N_7707,N_1934,N_2762);
nand U7708 (N_7708,N_3706,N_2338);
and U7709 (N_7709,N_4054,N_745);
nand U7710 (N_7710,N_3304,N_3482);
nand U7711 (N_7711,N_3114,N_2427);
nand U7712 (N_7712,N_3599,N_3960);
nand U7713 (N_7713,N_921,N_3393);
and U7714 (N_7714,N_2468,N_1483);
or U7715 (N_7715,N_3236,N_1752);
or U7716 (N_7716,N_2361,N_3274);
nand U7717 (N_7717,N_1387,N_2577);
nand U7718 (N_7718,N_1830,N_367);
nor U7719 (N_7719,N_699,N_1511);
or U7720 (N_7720,N_4745,N_4280);
nor U7721 (N_7721,N_4173,N_4139);
and U7722 (N_7722,N_2079,N_3917);
nand U7723 (N_7723,N_3339,N_399);
or U7724 (N_7724,N_2118,N_319);
nand U7725 (N_7725,N_3172,N_2352);
and U7726 (N_7726,N_32,N_2728);
and U7727 (N_7727,N_3877,N_1230);
or U7728 (N_7728,N_2802,N_1056);
or U7729 (N_7729,N_4610,N_473);
nor U7730 (N_7730,N_4838,N_659);
nand U7731 (N_7731,N_3795,N_3884);
nor U7732 (N_7732,N_2976,N_4496);
nor U7733 (N_7733,N_4110,N_1827);
and U7734 (N_7734,N_2798,N_30);
or U7735 (N_7735,N_3840,N_4933);
or U7736 (N_7736,N_3036,N_2013);
nor U7737 (N_7737,N_2306,N_2785);
nor U7738 (N_7738,N_1541,N_3343);
nor U7739 (N_7739,N_3716,N_4525);
or U7740 (N_7740,N_686,N_2138);
or U7741 (N_7741,N_418,N_3575);
and U7742 (N_7742,N_2007,N_1887);
nand U7743 (N_7743,N_4625,N_2588);
nor U7744 (N_7744,N_2846,N_3459);
or U7745 (N_7745,N_3305,N_1147);
nand U7746 (N_7746,N_4866,N_2180);
nor U7747 (N_7747,N_2948,N_2897);
and U7748 (N_7748,N_183,N_2251);
or U7749 (N_7749,N_848,N_4075);
or U7750 (N_7750,N_643,N_3101);
and U7751 (N_7751,N_3379,N_4142);
nand U7752 (N_7752,N_871,N_1007);
or U7753 (N_7753,N_2728,N_4259);
nand U7754 (N_7754,N_3427,N_1246);
and U7755 (N_7755,N_1041,N_59);
nand U7756 (N_7756,N_2368,N_1396);
nand U7757 (N_7757,N_1202,N_95);
nand U7758 (N_7758,N_2382,N_487);
and U7759 (N_7759,N_1320,N_1765);
nor U7760 (N_7760,N_2687,N_3796);
and U7761 (N_7761,N_1093,N_3007);
or U7762 (N_7762,N_562,N_3451);
nand U7763 (N_7763,N_2039,N_3474);
nor U7764 (N_7764,N_623,N_773);
nor U7765 (N_7765,N_2215,N_895);
and U7766 (N_7766,N_1509,N_267);
and U7767 (N_7767,N_2868,N_773);
and U7768 (N_7768,N_347,N_384);
and U7769 (N_7769,N_4606,N_1378);
nand U7770 (N_7770,N_3844,N_3535);
xnor U7771 (N_7771,N_2846,N_2715);
or U7772 (N_7772,N_517,N_316);
nand U7773 (N_7773,N_4969,N_4274);
and U7774 (N_7774,N_2146,N_3225);
or U7775 (N_7775,N_1456,N_2373);
nor U7776 (N_7776,N_1962,N_1410);
nand U7777 (N_7777,N_4933,N_950);
and U7778 (N_7778,N_2136,N_4725);
nor U7779 (N_7779,N_3918,N_1779);
nor U7780 (N_7780,N_20,N_1944);
nor U7781 (N_7781,N_783,N_1642);
nand U7782 (N_7782,N_2811,N_4588);
or U7783 (N_7783,N_2205,N_4506);
nor U7784 (N_7784,N_2530,N_3289);
nand U7785 (N_7785,N_3281,N_1257);
and U7786 (N_7786,N_3928,N_3051);
nand U7787 (N_7787,N_3336,N_2807);
and U7788 (N_7788,N_3032,N_4296);
or U7789 (N_7789,N_171,N_689);
and U7790 (N_7790,N_3048,N_1257);
nand U7791 (N_7791,N_82,N_1030);
nor U7792 (N_7792,N_119,N_2795);
or U7793 (N_7793,N_2673,N_4324);
nand U7794 (N_7794,N_638,N_2151);
and U7795 (N_7795,N_886,N_199);
nor U7796 (N_7796,N_2801,N_2182);
nor U7797 (N_7797,N_1172,N_4403);
or U7798 (N_7798,N_4888,N_3798);
and U7799 (N_7799,N_1182,N_3703);
nand U7800 (N_7800,N_3462,N_801);
and U7801 (N_7801,N_4490,N_979);
or U7802 (N_7802,N_63,N_1437);
and U7803 (N_7803,N_2366,N_1914);
or U7804 (N_7804,N_2073,N_386);
nand U7805 (N_7805,N_3523,N_4958);
or U7806 (N_7806,N_1212,N_1611);
nor U7807 (N_7807,N_2111,N_2038);
and U7808 (N_7808,N_2548,N_1490);
and U7809 (N_7809,N_4826,N_527);
and U7810 (N_7810,N_1043,N_696);
and U7811 (N_7811,N_2895,N_3359);
nand U7812 (N_7812,N_3403,N_1307);
nor U7813 (N_7813,N_1316,N_3950);
and U7814 (N_7814,N_4219,N_923);
nor U7815 (N_7815,N_770,N_3880);
xnor U7816 (N_7816,N_2555,N_1141);
nand U7817 (N_7817,N_276,N_2217);
nor U7818 (N_7818,N_3933,N_3423);
nand U7819 (N_7819,N_3032,N_3678);
nand U7820 (N_7820,N_4158,N_136);
nand U7821 (N_7821,N_2823,N_2299);
nand U7822 (N_7822,N_404,N_4808);
nand U7823 (N_7823,N_234,N_4689);
and U7824 (N_7824,N_4812,N_314);
nand U7825 (N_7825,N_2969,N_4123);
and U7826 (N_7826,N_1190,N_3942);
or U7827 (N_7827,N_4744,N_544);
and U7828 (N_7828,N_3991,N_1159);
and U7829 (N_7829,N_623,N_1696);
or U7830 (N_7830,N_2411,N_2002);
nand U7831 (N_7831,N_792,N_3182);
or U7832 (N_7832,N_4310,N_4432);
nor U7833 (N_7833,N_1721,N_2484);
nand U7834 (N_7834,N_4,N_2269);
nand U7835 (N_7835,N_4917,N_878);
nor U7836 (N_7836,N_2323,N_2843);
nand U7837 (N_7837,N_4771,N_1261);
and U7838 (N_7838,N_2646,N_4553);
and U7839 (N_7839,N_2084,N_4906);
or U7840 (N_7840,N_2540,N_4916);
nor U7841 (N_7841,N_1710,N_2461);
and U7842 (N_7842,N_1606,N_4037);
nor U7843 (N_7843,N_3703,N_2517);
and U7844 (N_7844,N_3609,N_1896);
and U7845 (N_7845,N_2285,N_2374);
or U7846 (N_7846,N_1241,N_1781);
xnor U7847 (N_7847,N_727,N_1091);
nand U7848 (N_7848,N_3259,N_3257);
xnor U7849 (N_7849,N_212,N_1307);
and U7850 (N_7850,N_2636,N_1673);
or U7851 (N_7851,N_1370,N_4189);
or U7852 (N_7852,N_2257,N_1867);
nand U7853 (N_7853,N_4589,N_3875);
xor U7854 (N_7854,N_4231,N_2857);
or U7855 (N_7855,N_4532,N_2726);
nand U7856 (N_7856,N_3153,N_1909);
nand U7857 (N_7857,N_1846,N_1491);
and U7858 (N_7858,N_2577,N_203);
or U7859 (N_7859,N_1368,N_4709);
and U7860 (N_7860,N_4689,N_3638);
nand U7861 (N_7861,N_3872,N_2077);
nor U7862 (N_7862,N_4229,N_207);
and U7863 (N_7863,N_2690,N_1334);
nor U7864 (N_7864,N_1055,N_4596);
nand U7865 (N_7865,N_2015,N_1668);
nor U7866 (N_7866,N_3221,N_952);
nor U7867 (N_7867,N_3183,N_2824);
nor U7868 (N_7868,N_838,N_958);
nor U7869 (N_7869,N_3360,N_3947);
and U7870 (N_7870,N_742,N_4705);
xor U7871 (N_7871,N_4642,N_440);
nand U7872 (N_7872,N_2936,N_876);
nor U7873 (N_7873,N_2403,N_2838);
or U7874 (N_7874,N_2316,N_696);
nor U7875 (N_7875,N_1972,N_4934);
nand U7876 (N_7876,N_960,N_842);
nand U7877 (N_7877,N_1240,N_3038);
nor U7878 (N_7878,N_2703,N_3576);
nor U7879 (N_7879,N_1484,N_1047);
or U7880 (N_7880,N_1113,N_1325);
nor U7881 (N_7881,N_3405,N_4399);
xnor U7882 (N_7882,N_3353,N_4275);
and U7883 (N_7883,N_3831,N_4675);
and U7884 (N_7884,N_1717,N_4370);
and U7885 (N_7885,N_3987,N_1027);
or U7886 (N_7886,N_1870,N_380);
xnor U7887 (N_7887,N_3176,N_2784);
and U7888 (N_7888,N_200,N_4557);
nand U7889 (N_7889,N_2596,N_3841);
or U7890 (N_7890,N_2560,N_2502);
nand U7891 (N_7891,N_2425,N_2763);
nor U7892 (N_7892,N_3313,N_2055);
nor U7893 (N_7893,N_3082,N_848);
nor U7894 (N_7894,N_2254,N_3299);
and U7895 (N_7895,N_2607,N_2895);
or U7896 (N_7896,N_3092,N_4362);
nor U7897 (N_7897,N_2536,N_3711);
xnor U7898 (N_7898,N_3781,N_4192);
nor U7899 (N_7899,N_3387,N_2969);
nor U7900 (N_7900,N_4623,N_3840);
nand U7901 (N_7901,N_2748,N_853);
and U7902 (N_7902,N_1975,N_4666);
or U7903 (N_7903,N_4187,N_3128);
nand U7904 (N_7904,N_625,N_143);
nor U7905 (N_7905,N_4836,N_3118);
and U7906 (N_7906,N_461,N_4586);
nor U7907 (N_7907,N_4621,N_2219);
nor U7908 (N_7908,N_2489,N_1204);
and U7909 (N_7909,N_2895,N_2847);
and U7910 (N_7910,N_2313,N_1314);
or U7911 (N_7911,N_4414,N_2319);
or U7912 (N_7912,N_3257,N_2214);
nor U7913 (N_7913,N_2361,N_12);
or U7914 (N_7914,N_3718,N_2196);
or U7915 (N_7915,N_4625,N_334);
nor U7916 (N_7916,N_4327,N_3386);
or U7917 (N_7917,N_3664,N_398);
nor U7918 (N_7918,N_3872,N_437);
nand U7919 (N_7919,N_847,N_1477);
nor U7920 (N_7920,N_2413,N_1472);
xor U7921 (N_7921,N_4710,N_3645);
nand U7922 (N_7922,N_4604,N_1175);
and U7923 (N_7923,N_1899,N_2870);
or U7924 (N_7924,N_4139,N_1247);
or U7925 (N_7925,N_3688,N_2129);
nand U7926 (N_7926,N_761,N_2750);
xnor U7927 (N_7927,N_3698,N_1386);
nand U7928 (N_7928,N_1293,N_1991);
nor U7929 (N_7929,N_1117,N_1256);
or U7930 (N_7930,N_2461,N_1686);
and U7931 (N_7931,N_1902,N_4461);
nor U7932 (N_7932,N_2983,N_726);
and U7933 (N_7933,N_2582,N_1364);
xnor U7934 (N_7934,N_3567,N_1724);
nand U7935 (N_7935,N_2017,N_1476);
or U7936 (N_7936,N_1514,N_1960);
nand U7937 (N_7937,N_1391,N_532);
and U7938 (N_7938,N_2540,N_1204);
nand U7939 (N_7939,N_4922,N_437);
or U7940 (N_7940,N_439,N_4903);
and U7941 (N_7941,N_2464,N_2542);
nor U7942 (N_7942,N_1939,N_3750);
xnor U7943 (N_7943,N_2905,N_4995);
nand U7944 (N_7944,N_2532,N_118);
nor U7945 (N_7945,N_531,N_1688);
nor U7946 (N_7946,N_3400,N_4464);
nand U7947 (N_7947,N_2184,N_1092);
or U7948 (N_7948,N_3011,N_993);
and U7949 (N_7949,N_2778,N_2552);
nand U7950 (N_7950,N_138,N_1611);
and U7951 (N_7951,N_2530,N_2076);
or U7952 (N_7952,N_2508,N_383);
or U7953 (N_7953,N_3338,N_3397);
nor U7954 (N_7954,N_4496,N_74);
and U7955 (N_7955,N_3052,N_2192);
or U7956 (N_7956,N_1130,N_1528);
and U7957 (N_7957,N_2104,N_3008);
nor U7958 (N_7958,N_4288,N_2175);
nor U7959 (N_7959,N_4248,N_4802);
and U7960 (N_7960,N_884,N_446);
nand U7961 (N_7961,N_4774,N_2926);
nor U7962 (N_7962,N_4736,N_4549);
or U7963 (N_7963,N_3590,N_2227);
and U7964 (N_7964,N_4054,N_3832);
nand U7965 (N_7965,N_823,N_1612);
nand U7966 (N_7966,N_3023,N_3118);
xnor U7967 (N_7967,N_1841,N_3999);
nor U7968 (N_7968,N_1466,N_2749);
nand U7969 (N_7969,N_3188,N_4018);
nor U7970 (N_7970,N_1063,N_4667);
and U7971 (N_7971,N_3584,N_1880);
and U7972 (N_7972,N_2497,N_3711);
or U7973 (N_7973,N_4949,N_81);
and U7974 (N_7974,N_1601,N_1588);
or U7975 (N_7975,N_4678,N_3433);
and U7976 (N_7976,N_4478,N_1646);
or U7977 (N_7977,N_2061,N_3891);
and U7978 (N_7978,N_247,N_1557);
nor U7979 (N_7979,N_2713,N_4677);
nor U7980 (N_7980,N_2906,N_4416);
nand U7981 (N_7981,N_4646,N_4289);
nor U7982 (N_7982,N_2935,N_2274);
or U7983 (N_7983,N_3526,N_1317);
or U7984 (N_7984,N_805,N_3213);
nand U7985 (N_7985,N_1142,N_1283);
and U7986 (N_7986,N_4283,N_2287);
nand U7987 (N_7987,N_667,N_2142);
nand U7988 (N_7988,N_318,N_4593);
nor U7989 (N_7989,N_2300,N_1086);
and U7990 (N_7990,N_3099,N_2397);
nand U7991 (N_7991,N_3840,N_3003);
or U7992 (N_7992,N_1,N_24);
nand U7993 (N_7993,N_197,N_4086);
or U7994 (N_7994,N_1522,N_229);
or U7995 (N_7995,N_3976,N_577);
nor U7996 (N_7996,N_3139,N_751);
nand U7997 (N_7997,N_4681,N_3358);
or U7998 (N_7998,N_1941,N_1362);
nor U7999 (N_7999,N_2293,N_37);
and U8000 (N_8000,N_1462,N_3313);
and U8001 (N_8001,N_2951,N_3501);
nand U8002 (N_8002,N_4935,N_2130);
or U8003 (N_8003,N_4459,N_2209);
or U8004 (N_8004,N_4919,N_3322);
or U8005 (N_8005,N_2890,N_4066);
and U8006 (N_8006,N_4558,N_4736);
nand U8007 (N_8007,N_4917,N_2060);
nand U8008 (N_8008,N_3834,N_4592);
or U8009 (N_8009,N_3028,N_501);
and U8010 (N_8010,N_1440,N_3548);
nand U8011 (N_8011,N_1490,N_1552);
or U8012 (N_8012,N_2970,N_1442);
or U8013 (N_8013,N_1902,N_3748);
or U8014 (N_8014,N_2889,N_3486);
and U8015 (N_8015,N_2967,N_4440);
nand U8016 (N_8016,N_3008,N_3713);
and U8017 (N_8017,N_928,N_2531);
and U8018 (N_8018,N_4311,N_4968);
nand U8019 (N_8019,N_1974,N_3468);
nand U8020 (N_8020,N_2308,N_3526);
nand U8021 (N_8021,N_4449,N_94);
and U8022 (N_8022,N_4538,N_1695);
and U8023 (N_8023,N_2379,N_4174);
nand U8024 (N_8024,N_1921,N_1949);
nand U8025 (N_8025,N_2817,N_3992);
and U8026 (N_8026,N_990,N_4161);
or U8027 (N_8027,N_1772,N_1280);
nand U8028 (N_8028,N_3818,N_1967);
nand U8029 (N_8029,N_3666,N_2564);
or U8030 (N_8030,N_3935,N_2315);
or U8031 (N_8031,N_2336,N_825);
nand U8032 (N_8032,N_4807,N_1994);
xnor U8033 (N_8033,N_1521,N_4284);
nor U8034 (N_8034,N_1034,N_1283);
or U8035 (N_8035,N_971,N_2208);
nor U8036 (N_8036,N_4115,N_61);
nor U8037 (N_8037,N_1550,N_4220);
and U8038 (N_8038,N_3327,N_3889);
nand U8039 (N_8039,N_1173,N_1676);
and U8040 (N_8040,N_1913,N_1736);
nand U8041 (N_8041,N_4619,N_2622);
nor U8042 (N_8042,N_3322,N_3033);
and U8043 (N_8043,N_479,N_2284);
and U8044 (N_8044,N_2769,N_4576);
or U8045 (N_8045,N_1224,N_3112);
nand U8046 (N_8046,N_813,N_2097);
and U8047 (N_8047,N_3250,N_4610);
nand U8048 (N_8048,N_3176,N_3071);
or U8049 (N_8049,N_2682,N_3151);
and U8050 (N_8050,N_500,N_217);
nor U8051 (N_8051,N_4698,N_1503);
and U8052 (N_8052,N_1987,N_3254);
and U8053 (N_8053,N_335,N_2337);
nand U8054 (N_8054,N_4221,N_2545);
or U8055 (N_8055,N_4995,N_2605);
xor U8056 (N_8056,N_484,N_1150);
nand U8057 (N_8057,N_1389,N_4592);
or U8058 (N_8058,N_1304,N_487);
and U8059 (N_8059,N_473,N_1624);
or U8060 (N_8060,N_1134,N_1465);
and U8061 (N_8061,N_4157,N_4093);
and U8062 (N_8062,N_314,N_955);
or U8063 (N_8063,N_3834,N_4493);
nand U8064 (N_8064,N_1600,N_4961);
nor U8065 (N_8065,N_4360,N_1439);
and U8066 (N_8066,N_2752,N_1691);
nor U8067 (N_8067,N_4710,N_815);
nand U8068 (N_8068,N_228,N_868);
and U8069 (N_8069,N_1296,N_3363);
nand U8070 (N_8070,N_2890,N_4241);
or U8071 (N_8071,N_141,N_1924);
nand U8072 (N_8072,N_3722,N_3088);
and U8073 (N_8073,N_3470,N_4737);
nand U8074 (N_8074,N_3291,N_4018);
xnor U8075 (N_8075,N_2637,N_1464);
and U8076 (N_8076,N_2337,N_2799);
and U8077 (N_8077,N_3506,N_4421);
nor U8078 (N_8078,N_1954,N_2263);
nor U8079 (N_8079,N_2900,N_2119);
nor U8080 (N_8080,N_3687,N_2571);
or U8081 (N_8081,N_3001,N_4887);
nand U8082 (N_8082,N_4633,N_3853);
or U8083 (N_8083,N_2526,N_4708);
or U8084 (N_8084,N_4095,N_2030);
nand U8085 (N_8085,N_2553,N_1468);
or U8086 (N_8086,N_1638,N_2557);
and U8087 (N_8087,N_3386,N_1773);
nor U8088 (N_8088,N_3898,N_4303);
and U8089 (N_8089,N_1948,N_3731);
or U8090 (N_8090,N_2374,N_2963);
nor U8091 (N_8091,N_2207,N_4231);
nor U8092 (N_8092,N_2593,N_4825);
nor U8093 (N_8093,N_907,N_4489);
and U8094 (N_8094,N_1592,N_1496);
or U8095 (N_8095,N_4682,N_4674);
or U8096 (N_8096,N_3991,N_2605);
or U8097 (N_8097,N_3904,N_93);
nor U8098 (N_8098,N_2852,N_1968);
or U8099 (N_8099,N_218,N_1115);
and U8100 (N_8100,N_2815,N_2335);
and U8101 (N_8101,N_3646,N_2077);
nand U8102 (N_8102,N_4908,N_3023);
and U8103 (N_8103,N_4246,N_2453);
or U8104 (N_8104,N_408,N_3667);
and U8105 (N_8105,N_1534,N_1105);
and U8106 (N_8106,N_598,N_2701);
and U8107 (N_8107,N_542,N_393);
nor U8108 (N_8108,N_4008,N_1226);
and U8109 (N_8109,N_2161,N_2402);
nor U8110 (N_8110,N_278,N_3565);
nor U8111 (N_8111,N_4653,N_1715);
or U8112 (N_8112,N_4254,N_1347);
nand U8113 (N_8113,N_4993,N_164);
nand U8114 (N_8114,N_1543,N_570);
or U8115 (N_8115,N_1976,N_975);
nand U8116 (N_8116,N_379,N_647);
or U8117 (N_8117,N_807,N_132);
nor U8118 (N_8118,N_2668,N_3977);
or U8119 (N_8119,N_3185,N_4356);
nand U8120 (N_8120,N_3476,N_4575);
nand U8121 (N_8121,N_2155,N_420);
nand U8122 (N_8122,N_1052,N_4787);
nor U8123 (N_8123,N_2691,N_3477);
and U8124 (N_8124,N_2140,N_3725);
and U8125 (N_8125,N_2041,N_3759);
and U8126 (N_8126,N_3480,N_3900);
nor U8127 (N_8127,N_1661,N_1012);
or U8128 (N_8128,N_1970,N_4444);
and U8129 (N_8129,N_1321,N_2918);
nor U8130 (N_8130,N_3615,N_3381);
nor U8131 (N_8131,N_2122,N_1603);
nand U8132 (N_8132,N_1692,N_1989);
or U8133 (N_8133,N_1236,N_4447);
and U8134 (N_8134,N_1867,N_3078);
or U8135 (N_8135,N_4446,N_3735);
nor U8136 (N_8136,N_887,N_4626);
nor U8137 (N_8137,N_3117,N_207);
nand U8138 (N_8138,N_754,N_4232);
nor U8139 (N_8139,N_3783,N_4482);
and U8140 (N_8140,N_2043,N_3166);
and U8141 (N_8141,N_725,N_1024);
nor U8142 (N_8142,N_3919,N_4379);
or U8143 (N_8143,N_697,N_4949);
xnor U8144 (N_8144,N_716,N_1219);
nor U8145 (N_8145,N_3985,N_2071);
nor U8146 (N_8146,N_4089,N_71);
nand U8147 (N_8147,N_4126,N_2588);
and U8148 (N_8148,N_2678,N_2787);
nor U8149 (N_8149,N_461,N_3716);
or U8150 (N_8150,N_3232,N_850);
and U8151 (N_8151,N_3697,N_4634);
nor U8152 (N_8152,N_1579,N_4891);
and U8153 (N_8153,N_999,N_865);
and U8154 (N_8154,N_2129,N_2229);
nor U8155 (N_8155,N_4434,N_2419);
nand U8156 (N_8156,N_2257,N_2288);
and U8157 (N_8157,N_1820,N_4191);
or U8158 (N_8158,N_2654,N_1442);
or U8159 (N_8159,N_4038,N_226);
nand U8160 (N_8160,N_3257,N_122);
nor U8161 (N_8161,N_4279,N_3248);
nand U8162 (N_8162,N_1305,N_3145);
nand U8163 (N_8163,N_4068,N_2875);
nor U8164 (N_8164,N_1203,N_3017);
or U8165 (N_8165,N_219,N_158);
nand U8166 (N_8166,N_41,N_2795);
nand U8167 (N_8167,N_3111,N_2150);
or U8168 (N_8168,N_4532,N_2557);
or U8169 (N_8169,N_2195,N_3675);
nand U8170 (N_8170,N_2031,N_4340);
or U8171 (N_8171,N_2116,N_3817);
nor U8172 (N_8172,N_2759,N_1425);
nand U8173 (N_8173,N_2163,N_4428);
nand U8174 (N_8174,N_2146,N_4437);
or U8175 (N_8175,N_4833,N_4419);
nand U8176 (N_8176,N_1093,N_1503);
or U8177 (N_8177,N_1594,N_2433);
or U8178 (N_8178,N_2086,N_3933);
nand U8179 (N_8179,N_4846,N_1508);
nor U8180 (N_8180,N_2587,N_1116);
nor U8181 (N_8181,N_1299,N_2120);
or U8182 (N_8182,N_111,N_3733);
or U8183 (N_8183,N_2966,N_2480);
nand U8184 (N_8184,N_795,N_1869);
nor U8185 (N_8185,N_4931,N_4255);
or U8186 (N_8186,N_2343,N_4431);
or U8187 (N_8187,N_3732,N_4514);
nor U8188 (N_8188,N_1546,N_2826);
nor U8189 (N_8189,N_2166,N_1212);
nand U8190 (N_8190,N_3712,N_3353);
nor U8191 (N_8191,N_1778,N_2460);
or U8192 (N_8192,N_3965,N_706);
nor U8193 (N_8193,N_1924,N_2049);
nor U8194 (N_8194,N_4235,N_729);
or U8195 (N_8195,N_1165,N_4664);
nor U8196 (N_8196,N_2084,N_2337);
or U8197 (N_8197,N_4572,N_4392);
and U8198 (N_8198,N_202,N_838);
and U8199 (N_8199,N_1155,N_1466);
nor U8200 (N_8200,N_4841,N_3580);
nand U8201 (N_8201,N_793,N_3363);
and U8202 (N_8202,N_3825,N_2454);
nor U8203 (N_8203,N_3680,N_4499);
nand U8204 (N_8204,N_991,N_2840);
or U8205 (N_8205,N_2828,N_4176);
and U8206 (N_8206,N_1888,N_4592);
or U8207 (N_8207,N_517,N_3183);
or U8208 (N_8208,N_1360,N_4583);
and U8209 (N_8209,N_57,N_297);
nand U8210 (N_8210,N_1727,N_1336);
and U8211 (N_8211,N_4635,N_2077);
or U8212 (N_8212,N_1614,N_2407);
and U8213 (N_8213,N_2340,N_3955);
nand U8214 (N_8214,N_652,N_3054);
nor U8215 (N_8215,N_2,N_4013);
nor U8216 (N_8216,N_703,N_4180);
nand U8217 (N_8217,N_3796,N_950);
xnor U8218 (N_8218,N_4192,N_691);
and U8219 (N_8219,N_1204,N_2503);
nand U8220 (N_8220,N_3150,N_3396);
or U8221 (N_8221,N_1081,N_2230);
nor U8222 (N_8222,N_378,N_492);
or U8223 (N_8223,N_327,N_4473);
or U8224 (N_8224,N_1261,N_3341);
and U8225 (N_8225,N_1656,N_2991);
and U8226 (N_8226,N_3795,N_2169);
nand U8227 (N_8227,N_2466,N_755);
xor U8228 (N_8228,N_3416,N_3304);
nor U8229 (N_8229,N_4925,N_1476);
nor U8230 (N_8230,N_4657,N_3907);
nand U8231 (N_8231,N_1241,N_4801);
or U8232 (N_8232,N_14,N_3499);
nor U8233 (N_8233,N_3132,N_1589);
nor U8234 (N_8234,N_2723,N_784);
nand U8235 (N_8235,N_2416,N_3843);
or U8236 (N_8236,N_3619,N_3685);
nand U8237 (N_8237,N_2659,N_535);
and U8238 (N_8238,N_4955,N_299);
nand U8239 (N_8239,N_3450,N_1775);
nor U8240 (N_8240,N_4034,N_1829);
nand U8241 (N_8241,N_4723,N_3873);
nand U8242 (N_8242,N_980,N_217);
and U8243 (N_8243,N_1040,N_2869);
or U8244 (N_8244,N_3393,N_85);
nand U8245 (N_8245,N_3335,N_1567);
and U8246 (N_8246,N_1470,N_4595);
nand U8247 (N_8247,N_3547,N_692);
nand U8248 (N_8248,N_4530,N_1552);
nand U8249 (N_8249,N_4255,N_1381);
nor U8250 (N_8250,N_867,N_3049);
nor U8251 (N_8251,N_2183,N_4686);
or U8252 (N_8252,N_4587,N_1249);
nor U8253 (N_8253,N_2083,N_1432);
nand U8254 (N_8254,N_131,N_2327);
and U8255 (N_8255,N_2450,N_303);
and U8256 (N_8256,N_4917,N_687);
nand U8257 (N_8257,N_4873,N_428);
or U8258 (N_8258,N_2880,N_2592);
nand U8259 (N_8259,N_3654,N_361);
nor U8260 (N_8260,N_4272,N_5);
nor U8261 (N_8261,N_1466,N_4195);
nor U8262 (N_8262,N_2487,N_3002);
nor U8263 (N_8263,N_194,N_2468);
or U8264 (N_8264,N_4691,N_238);
nor U8265 (N_8265,N_4138,N_2467);
or U8266 (N_8266,N_4671,N_3552);
nor U8267 (N_8267,N_1043,N_4077);
nor U8268 (N_8268,N_642,N_1721);
and U8269 (N_8269,N_1012,N_1516);
and U8270 (N_8270,N_1601,N_2837);
nand U8271 (N_8271,N_4669,N_1787);
and U8272 (N_8272,N_83,N_5);
nand U8273 (N_8273,N_4595,N_3449);
and U8274 (N_8274,N_4110,N_1482);
or U8275 (N_8275,N_1137,N_1115);
nor U8276 (N_8276,N_1585,N_2035);
or U8277 (N_8277,N_181,N_834);
or U8278 (N_8278,N_1844,N_3693);
and U8279 (N_8279,N_4486,N_2538);
nor U8280 (N_8280,N_2118,N_1763);
nand U8281 (N_8281,N_2937,N_3163);
nand U8282 (N_8282,N_335,N_2523);
and U8283 (N_8283,N_3492,N_4644);
nand U8284 (N_8284,N_2833,N_2393);
or U8285 (N_8285,N_678,N_803);
xor U8286 (N_8286,N_2502,N_2256);
nand U8287 (N_8287,N_4559,N_4422);
and U8288 (N_8288,N_1664,N_3937);
nand U8289 (N_8289,N_3419,N_1806);
nand U8290 (N_8290,N_4810,N_3577);
nand U8291 (N_8291,N_2056,N_4997);
or U8292 (N_8292,N_17,N_3932);
nor U8293 (N_8293,N_2295,N_1601);
or U8294 (N_8294,N_744,N_3880);
nor U8295 (N_8295,N_4229,N_1059);
nand U8296 (N_8296,N_4097,N_4775);
or U8297 (N_8297,N_2453,N_2386);
and U8298 (N_8298,N_3144,N_1639);
nand U8299 (N_8299,N_2741,N_4952);
and U8300 (N_8300,N_4678,N_4053);
and U8301 (N_8301,N_3672,N_3785);
or U8302 (N_8302,N_1168,N_802);
or U8303 (N_8303,N_4831,N_1992);
and U8304 (N_8304,N_179,N_2817);
nor U8305 (N_8305,N_4857,N_4389);
nor U8306 (N_8306,N_145,N_3713);
nor U8307 (N_8307,N_4169,N_2979);
nor U8308 (N_8308,N_886,N_3286);
nand U8309 (N_8309,N_3675,N_3406);
or U8310 (N_8310,N_2282,N_158);
nand U8311 (N_8311,N_1565,N_1934);
nor U8312 (N_8312,N_2179,N_2119);
and U8313 (N_8313,N_159,N_811);
nor U8314 (N_8314,N_1493,N_3227);
nor U8315 (N_8315,N_3357,N_1);
or U8316 (N_8316,N_2818,N_1837);
nor U8317 (N_8317,N_4221,N_3472);
and U8318 (N_8318,N_2301,N_3783);
nand U8319 (N_8319,N_647,N_2309);
nor U8320 (N_8320,N_2284,N_1718);
nand U8321 (N_8321,N_3591,N_1271);
nand U8322 (N_8322,N_3600,N_1741);
and U8323 (N_8323,N_1907,N_4254);
and U8324 (N_8324,N_321,N_1812);
and U8325 (N_8325,N_841,N_4951);
nand U8326 (N_8326,N_584,N_924);
nor U8327 (N_8327,N_2176,N_1646);
and U8328 (N_8328,N_3034,N_1203);
nor U8329 (N_8329,N_2397,N_333);
nor U8330 (N_8330,N_112,N_372);
or U8331 (N_8331,N_3096,N_855);
nand U8332 (N_8332,N_3452,N_3974);
or U8333 (N_8333,N_384,N_709);
and U8334 (N_8334,N_4090,N_4804);
nand U8335 (N_8335,N_2412,N_4416);
nor U8336 (N_8336,N_4069,N_2017);
or U8337 (N_8337,N_65,N_788);
nand U8338 (N_8338,N_4214,N_4272);
nand U8339 (N_8339,N_1659,N_4033);
or U8340 (N_8340,N_4007,N_1733);
and U8341 (N_8341,N_1218,N_4022);
nor U8342 (N_8342,N_3185,N_3992);
xor U8343 (N_8343,N_2676,N_1719);
or U8344 (N_8344,N_4005,N_3300);
and U8345 (N_8345,N_92,N_4724);
nor U8346 (N_8346,N_4381,N_1865);
or U8347 (N_8347,N_2757,N_3682);
nor U8348 (N_8348,N_4101,N_182);
nor U8349 (N_8349,N_4790,N_4413);
or U8350 (N_8350,N_3623,N_2215);
or U8351 (N_8351,N_4316,N_3925);
nand U8352 (N_8352,N_2868,N_1913);
nor U8353 (N_8353,N_4253,N_2800);
nor U8354 (N_8354,N_3392,N_2393);
xnor U8355 (N_8355,N_3082,N_3930);
and U8356 (N_8356,N_3680,N_842);
nand U8357 (N_8357,N_2350,N_1743);
and U8358 (N_8358,N_4266,N_3513);
nand U8359 (N_8359,N_425,N_2854);
nor U8360 (N_8360,N_3449,N_2227);
and U8361 (N_8361,N_2720,N_4744);
nor U8362 (N_8362,N_3055,N_4158);
nand U8363 (N_8363,N_4914,N_4378);
nand U8364 (N_8364,N_3964,N_523);
nor U8365 (N_8365,N_2106,N_1187);
nor U8366 (N_8366,N_251,N_967);
or U8367 (N_8367,N_46,N_2960);
nor U8368 (N_8368,N_3873,N_3331);
or U8369 (N_8369,N_3872,N_4521);
nand U8370 (N_8370,N_1645,N_3030);
nor U8371 (N_8371,N_4191,N_1052);
or U8372 (N_8372,N_363,N_4474);
or U8373 (N_8373,N_3051,N_2929);
nand U8374 (N_8374,N_1268,N_4230);
nor U8375 (N_8375,N_1132,N_802);
nand U8376 (N_8376,N_1906,N_2682);
and U8377 (N_8377,N_3192,N_3129);
and U8378 (N_8378,N_4008,N_3286);
or U8379 (N_8379,N_584,N_4308);
nand U8380 (N_8380,N_2136,N_3405);
and U8381 (N_8381,N_2689,N_419);
nor U8382 (N_8382,N_2848,N_302);
nand U8383 (N_8383,N_4463,N_4979);
and U8384 (N_8384,N_2007,N_2469);
and U8385 (N_8385,N_1639,N_2880);
and U8386 (N_8386,N_3324,N_2027);
nand U8387 (N_8387,N_3907,N_725);
nand U8388 (N_8388,N_3933,N_2229);
nand U8389 (N_8389,N_3642,N_379);
nor U8390 (N_8390,N_43,N_854);
and U8391 (N_8391,N_1041,N_3315);
nand U8392 (N_8392,N_3012,N_4108);
xnor U8393 (N_8393,N_4896,N_1588);
and U8394 (N_8394,N_4009,N_103);
nor U8395 (N_8395,N_3980,N_2901);
or U8396 (N_8396,N_3688,N_2566);
and U8397 (N_8397,N_2881,N_1290);
nor U8398 (N_8398,N_1204,N_2605);
or U8399 (N_8399,N_4169,N_3356);
and U8400 (N_8400,N_4330,N_295);
nor U8401 (N_8401,N_1705,N_3405);
nor U8402 (N_8402,N_977,N_3377);
and U8403 (N_8403,N_4728,N_1929);
nand U8404 (N_8404,N_3355,N_4222);
nand U8405 (N_8405,N_2116,N_4042);
and U8406 (N_8406,N_667,N_3934);
nor U8407 (N_8407,N_1553,N_2265);
nand U8408 (N_8408,N_985,N_4811);
or U8409 (N_8409,N_2091,N_497);
and U8410 (N_8410,N_927,N_764);
and U8411 (N_8411,N_4615,N_1335);
nand U8412 (N_8412,N_1082,N_3006);
or U8413 (N_8413,N_4719,N_3132);
and U8414 (N_8414,N_2918,N_1657);
or U8415 (N_8415,N_3341,N_3617);
or U8416 (N_8416,N_1349,N_1295);
xor U8417 (N_8417,N_2841,N_4631);
and U8418 (N_8418,N_821,N_3668);
or U8419 (N_8419,N_4932,N_4014);
and U8420 (N_8420,N_1651,N_1204);
or U8421 (N_8421,N_4402,N_226);
nand U8422 (N_8422,N_1044,N_3624);
nor U8423 (N_8423,N_4724,N_4379);
nand U8424 (N_8424,N_2121,N_4198);
and U8425 (N_8425,N_3868,N_1536);
nor U8426 (N_8426,N_1293,N_3681);
or U8427 (N_8427,N_1917,N_1459);
and U8428 (N_8428,N_1288,N_1491);
or U8429 (N_8429,N_321,N_4712);
nand U8430 (N_8430,N_4470,N_4042);
nand U8431 (N_8431,N_2041,N_187);
nor U8432 (N_8432,N_1064,N_2192);
and U8433 (N_8433,N_2649,N_1567);
and U8434 (N_8434,N_710,N_3336);
and U8435 (N_8435,N_3706,N_4011);
nor U8436 (N_8436,N_4965,N_3463);
and U8437 (N_8437,N_2580,N_2639);
and U8438 (N_8438,N_2110,N_1707);
nand U8439 (N_8439,N_3972,N_3712);
or U8440 (N_8440,N_1079,N_883);
nor U8441 (N_8441,N_4322,N_1252);
nand U8442 (N_8442,N_4145,N_295);
and U8443 (N_8443,N_1892,N_1887);
or U8444 (N_8444,N_3625,N_1296);
or U8445 (N_8445,N_649,N_3409);
or U8446 (N_8446,N_2007,N_3471);
nand U8447 (N_8447,N_1759,N_1237);
or U8448 (N_8448,N_2347,N_1088);
nand U8449 (N_8449,N_2891,N_4453);
or U8450 (N_8450,N_4078,N_3570);
nand U8451 (N_8451,N_3534,N_1076);
nor U8452 (N_8452,N_2369,N_1092);
nor U8453 (N_8453,N_650,N_1893);
and U8454 (N_8454,N_2253,N_351);
nand U8455 (N_8455,N_725,N_44);
nor U8456 (N_8456,N_3923,N_2344);
nand U8457 (N_8457,N_3735,N_332);
or U8458 (N_8458,N_4507,N_2306);
or U8459 (N_8459,N_2179,N_1008);
or U8460 (N_8460,N_983,N_3278);
nand U8461 (N_8461,N_940,N_147);
nand U8462 (N_8462,N_4248,N_1872);
and U8463 (N_8463,N_1239,N_3542);
or U8464 (N_8464,N_4631,N_1207);
nor U8465 (N_8465,N_1682,N_1054);
xnor U8466 (N_8466,N_4864,N_4264);
or U8467 (N_8467,N_979,N_4086);
and U8468 (N_8468,N_3819,N_3370);
nor U8469 (N_8469,N_3760,N_4481);
and U8470 (N_8470,N_3761,N_3835);
nor U8471 (N_8471,N_3282,N_1665);
nand U8472 (N_8472,N_2339,N_524);
nor U8473 (N_8473,N_247,N_1763);
nor U8474 (N_8474,N_4232,N_561);
nand U8475 (N_8475,N_2371,N_1281);
xnor U8476 (N_8476,N_4749,N_4243);
or U8477 (N_8477,N_2552,N_2091);
nor U8478 (N_8478,N_3916,N_1549);
and U8479 (N_8479,N_4428,N_3021);
and U8480 (N_8480,N_4870,N_959);
nor U8481 (N_8481,N_2832,N_575);
or U8482 (N_8482,N_3409,N_293);
or U8483 (N_8483,N_1329,N_1879);
nand U8484 (N_8484,N_143,N_2392);
or U8485 (N_8485,N_3918,N_605);
and U8486 (N_8486,N_4562,N_2509);
nor U8487 (N_8487,N_711,N_3813);
nor U8488 (N_8488,N_737,N_2581);
xor U8489 (N_8489,N_4016,N_3575);
or U8490 (N_8490,N_1663,N_2453);
and U8491 (N_8491,N_523,N_4069);
or U8492 (N_8492,N_570,N_3278);
and U8493 (N_8493,N_2550,N_2690);
nand U8494 (N_8494,N_566,N_3723);
xnor U8495 (N_8495,N_2315,N_4792);
nand U8496 (N_8496,N_2424,N_3046);
nand U8497 (N_8497,N_1946,N_4518);
nor U8498 (N_8498,N_2465,N_2405);
and U8499 (N_8499,N_2635,N_1801);
nor U8500 (N_8500,N_128,N_909);
or U8501 (N_8501,N_3738,N_1825);
nand U8502 (N_8502,N_1202,N_4497);
nand U8503 (N_8503,N_2758,N_4038);
nor U8504 (N_8504,N_3265,N_4459);
nand U8505 (N_8505,N_2498,N_4938);
nor U8506 (N_8506,N_3833,N_3170);
and U8507 (N_8507,N_1759,N_2295);
and U8508 (N_8508,N_3238,N_4336);
nor U8509 (N_8509,N_4607,N_389);
nand U8510 (N_8510,N_643,N_138);
or U8511 (N_8511,N_4826,N_3171);
xor U8512 (N_8512,N_2407,N_761);
nor U8513 (N_8513,N_939,N_4298);
and U8514 (N_8514,N_4585,N_4022);
and U8515 (N_8515,N_1489,N_1516);
nand U8516 (N_8516,N_3939,N_911);
and U8517 (N_8517,N_2950,N_2118);
xor U8518 (N_8518,N_3599,N_305);
nor U8519 (N_8519,N_3635,N_4227);
and U8520 (N_8520,N_3659,N_1814);
nor U8521 (N_8521,N_3458,N_3650);
and U8522 (N_8522,N_4723,N_4644);
nor U8523 (N_8523,N_3962,N_3063);
xnor U8524 (N_8524,N_1550,N_1077);
and U8525 (N_8525,N_360,N_4843);
and U8526 (N_8526,N_3300,N_4709);
and U8527 (N_8527,N_3722,N_4335);
nor U8528 (N_8528,N_2844,N_2657);
nor U8529 (N_8529,N_565,N_1073);
nor U8530 (N_8530,N_2806,N_3809);
nand U8531 (N_8531,N_1250,N_137);
and U8532 (N_8532,N_4726,N_337);
and U8533 (N_8533,N_1759,N_2555);
nor U8534 (N_8534,N_1677,N_4222);
and U8535 (N_8535,N_2230,N_1593);
nand U8536 (N_8536,N_2369,N_4861);
nand U8537 (N_8537,N_4723,N_1891);
or U8538 (N_8538,N_4439,N_2119);
nor U8539 (N_8539,N_2105,N_4657);
and U8540 (N_8540,N_4365,N_2107);
and U8541 (N_8541,N_700,N_2167);
nor U8542 (N_8542,N_1822,N_167);
and U8543 (N_8543,N_1674,N_1589);
or U8544 (N_8544,N_2751,N_1702);
xor U8545 (N_8545,N_1606,N_1437);
nand U8546 (N_8546,N_1161,N_11);
or U8547 (N_8547,N_817,N_1177);
nor U8548 (N_8548,N_4048,N_2558);
and U8549 (N_8549,N_4376,N_3936);
nand U8550 (N_8550,N_1523,N_3975);
and U8551 (N_8551,N_1275,N_3878);
nor U8552 (N_8552,N_4665,N_635);
and U8553 (N_8553,N_1230,N_1010);
nor U8554 (N_8554,N_1613,N_298);
nor U8555 (N_8555,N_1611,N_949);
xnor U8556 (N_8556,N_669,N_2933);
or U8557 (N_8557,N_3931,N_2579);
nor U8558 (N_8558,N_1762,N_4179);
nand U8559 (N_8559,N_2297,N_4016);
or U8560 (N_8560,N_2919,N_4320);
and U8561 (N_8561,N_1399,N_3165);
and U8562 (N_8562,N_141,N_1511);
nand U8563 (N_8563,N_4405,N_396);
xor U8564 (N_8564,N_1591,N_938);
nor U8565 (N_8565,N_3598,N_2934);
and U8566 (N_8566,N_3505,N_3093);
nand U8567 (N_8567,N_3129,N_307);
or U8568 (N_8568,N_806,N_4229);
and U8569 (N_8569,N_1640,N_3037);
or U8570 (N_8570,N_1989,N_594);
nand U8571 (N_8571,N_4393,N_572);
and U8572 (N_8572,N_2564,N_3736);
and U8573 (N_8573,N_4310,N_1126);
or U8574 (N_8574,N_2793,N_1510);
and U8575 (N_8575,N_465,N_2891);
nand U8576 (N_8576,N_1276,N_1813);
and U8577 (N_8577,N_4008,N_2312);
nand U8578 (N_8578,N_24,N_4701);
nand U8579 (N_8579,N_4944,N_4238);
and U8580 (N_8580,N_4957,N_3061);
and U8581 (N_8581,N_1297,N_3001);
nand U8582 (N_8582,N_3496,N_2182);
nor U8583 (N_8583,N_3712,N_4876);
or U8584 (N_8584,N_289,N_4281);
or U8585 (N_8585,N_4685,N_318);
nor U8586 (N_8586,N_1709,N_340);
nor U8587 (N_8587,N_4293,N_1323);
nand U8588 (N_8588,N_3204,N_3093);
and U8589 (N_8589,N_2539,N_4628);
and U8590 (N_8590,N_585,N_1761);
or U8591 (N_8591,N_560,N_373);
or U8592 (N_8592,N_332,N_3256);
or U8593 (N_8593,N_1142,N_1185);
and U8594 (N_8594,N_1429,N_4976);
and U8595 (N_8595,N_1034,N_2911);
nor U8596 (N_8596,N_1003,N_3920);
nor U8597 (N_8597,N_369,N_2696);
nor U8598 (N_8598,N_1475,N_4754);
and U8599 (N_8599,N_4519,N_1515);
and U8600 (N_8600,N_3234,N_1868);
or U8601 (N_8601,N_536,N_3866);
and U8602 (N_8602,N_1090,N_4392);
nand U8603 (N_8603,N_1669,N_258);
and U8604 (N_8604,N_1292,N_1483);
nand U8605 (N_8605,N_457,N_4105);
or U8606 (N_8606,N_3281,N_1947);
nor U8607 (N_8607,N_2241,N_1395);
or U8608 (N_8608,N_4996,N_2602);
nor U8609 (N_8609,N_340,N_3901);
or U8610 (N_8610,N_2528,N_3048);
and U8611 (N_8611,N_2015,N_3281);
and U8612 (N_8612,N_193,N_4534);
nand U8613 (N_8613,N_265,N_237);
or U8614 (N_8614,N_644,N_999);
nor U8615 (N_8615,N_2250,N_1814);
and U8616 (N_8616,N_1340,N_3086);
xnor U8617 (N_8617,N_1530,N_4446);
nand U8618 (N_8618,N_545,N_4641);
and U8619 (N_8619,N_2487,N_1196);
nor U8620 (N_8620,N_4669,N_362);
or U8621 (N_8621,N_2073,N_3326);
nor U8622 (N_8622,N_3706,N_4447);
and U8623 (N_8623,N_547,N_4148);
or U8624 (N_8624,N_4484,N_547);
nor U8625 (N_8625,N_2341,N_3554);
nor U8626 (N_8626,N_966,N_4087);
nand U8627 (N_8627,N_4042,N_4905);
nand U8628 (N_8628,N_37,N_1209);
and U8629 (N_8629,N_3299,N_4409);
nand U8630 (N_8630,N_1934,N_3163);
or U8631 (N_8631,N_1633,N_836);
and U8632 (N_8632,N_606,N_2016);
or U8633 (N_8633,N_1597,N_3902);
or U8634 (N_8634,N_4323,N_2386);
nor U8635 (N_8635,N_865,N_4799);
nand U8636 (N_8636,N_4753,N_3763);
or U8637 (N_8637,N_2823,N_4209);
nand U8638 (N_8638,N_2276,N_3780);
and U8639 (N_8639,N_608,N_634);
nor U8640 (N_8640,N_341,N_1465);
and U8641 (N_8641,N_440,N_1531);
and U8642 (N_8642,N_1350,N_935);
xnor U8643 (N_8643,N_998,N_2606);
nor U8644 (N_8644,N_1110,N_1931);
nor U8645 (N_8645,N_1550,N_825);
nor U8646 (N_8646,N_1423,N_2085);
nor U8647 (N_8647,N_96,N_2889);
or U8648 (N_8648,N_1112,N_4476);
or U8649 (N_8649,N_4414,N_2957);
and U8650 (N_8650,N_3718,N_1388);
nand U8651 (N_8651,N_2918,N_2738);
and U8652 (N_8652,N_3137,N_2367);
or U8653 (N_8653,N_3104,N_4807);
and U8654 (N_8654,N_3266,N_3422);
and U8655 (N_8655,N_2462,N_1234);
nor U8656 (N_8656,N_2753,N_935);
nand U8657 (N_8657,N_1384,N_4771);
xnor U8658 (N_8658,N_4911,N_1484);
and U8659 (N_8659,N_4907,N_2467);
and U8660 (N_8660,N_4946,N_1101);
or U8661 (N_8661,N_1917,N_524);
nor U8662 (N_8662,N_4030,N_2537);
or U8663 (N_8663,N_3263,N_2474);
or U8664 (N_8664,N_4217,N_1683);
nor U8665 (N_8665,N_264,N_166);
and U8666 (N_8666,N_2619,N_2934);
nor U8667 (N_8667,N_823,N_1876);
nor U8668 (N_8668,N_2630,N_2088);
and U8669 (N_8669,N_752,N_304);
and U8670 (N_8670,N_3939,N_4508);
nand U8671 (N_8671,N_4332,N_1329);
or U8672 (N_8672,N_4906,N_4005);
and U8673 (N_8673,N_2491,N_46);
nor U8674 (N_8674,N_3237,N_4713);
nor U8675 (N_8675,N_4800,N_4440);
and U8676 (N_8676,N_205,N_4948);
nand U8677 (N_8677,N_2898,N_2737);
and U8678 (N_8678,N_4929,N_3900);
nor U8679 (N_8679,N_3298,N_3631);
nand U8680 (N_8680,N_356,N_547);
and U8681 (N_8681,N_4659,N_948);
or U8682 (N_8682,N_2336,N_3121);
nor U8683 (N_8683,N_575,N_28);
nor U8684 (N_8684,N_4431,N_4677);
nand U8685 (N_8685,N_4182,N_4996);
or U8686 (N_8686,N_869,N_3861);
nor U8687 (N_8687,N_4440,N_1940);
and U8688 (N_8688,N_4687,N_329);
nand U8689 (N_8689,N_673,N_4118);
nor U8690 (N_8690,N_4610,N_4702);
nor U8691 (N_8691,N_1023,N_4852);
nor U8692 (N_8692,N_1067,N_102);
or U8693 (N_8693,N_3999,N_3240);
or U8694 (N_8694,N_4949,N_817);
nor U8695 (N_8695,N_923,N_4765);
or U8696 (N_8696,N_1279,N_1252);
nand U8697 (N_8697,N_1829,N_1717);
nand U8698 (N_8698,N_4861,N_1451);
and U8699 (N_8699,N_3316,N_2534);
and U8700 (N_8700,N_4072,N_159);
and U8701 (N_8701,N_2837,N_2909);
or U8702 (N_8702,N_4262,N_1391);
or U8703 (N_8703,N_864,N_211);
nor U8704 (N_8704,N_4108,N_2409);
nand U8705 (N_8705,N_797,N_442);
nand U8706 (N_8706,N_108,N_895);
nand U8707 (N_8707,N_2145,N_2152);
or U8708 (N_8708,N_3338,N_2119);
nor U8709 (N_8709,N_4252,N_1920);
nor U8710 (N_8710,N_1345,N_2735);
nor U8711 (N_8711,N_1427,N_4073);
nor U8712 (N_8712,N_1827,N_1723);
or U8713 (N_8713,N_2486,N_2517);
nand U8714 (N_8714,N_1258,N_2238);
and U8715 (N_8715,N_2728,N_3652);
nand U8716 (N_8716,N_2055,N_4160);
nand U8717 (N_8717,N_3675,N_3510);
or U8718 (N_8718,N_4055,N_2578);
and U8719 (N_8719,N_605,N_91);
or U8720 (N_8720,N_3095,N_4636);
nand U8721 (N_8721,N_1557,N_2592);
nand U8722 (N_8722,N_3805,N_432);
or U8723 (N_8723,N_4354,N_555);
nand U8724 (N_8724,N_549,N_321);
nand U8725 (N_8725,N_1537,N_2643);
and U8726 (N_8726,N_1226,N_2415);
nand U8727 (N_8727,N_2470,N_3275);
xnor U8728 (N_8728,N_4126,N_3938);
nor U8729 (N_8729,N_2654,N_3631);
nor U8730 (N_8730,N_4188,N_203);
nor U8731 (N_8731,N_2014,N_4435);
or U8732 (N_8732,N_4681,N_1491);
nor U8733 (N_8733,N_896,N_4820);
nand U8734 (N_8734,N_2171,N_3853);
or U8735 (N_8735,N_3239,N_2357);
or U8736 (N_8736,N_45,N_3034);
nand U8737 (N_8737,N_2312,N_2231);
and U8738 (N_8738,N_4695,N_4352);
and U8739 (N_8739,N_4002,N_102);
nor U8740 (N_8740,N_3292,N_4972);
or U8741 (N_8741,N_3360,N_392);
and U8742 (N_8742,N_3977,N_1271);
xnor U8743 (N_8743,N_429,N_4165);
and U8744 (N_8744,N_4889,N_3259);
or U8745 (N_8745,N_937,N_206);
nand U8746 (N_8746,N_233,N_323);
or U8747 (N_8747,N_436,N_4925);
nor U8748 (N_8748,N_1762,N_1162);
and U8749 (N_8749,N_2926,N_1503);
or U8750 (N_8750,N_3142,N_4728);
nor U8751 (N_8751,N_1351,N_2542);
nor U8752 (N_8752,N_1090,N_3621);
nand U8753 (N_8753,N_1964,N_3492);
or U8754 (N_8754,N_4462,N_382);
and U8755 (N_8755,N_57,N_4236);
nand U8756 (N_8756,N_891,N_1426);
and U8757 (N_8757,N_3883,N_289);
and U8758 (N_8758,N_3229,N_3381);
xor U8759 (N_8759,N_1769,N_432);
xor U8760 (N_8760,N_3882,N_2881);
nor U8761 (N_8761,N_1721,N_2360);
nand U8762 (N_8762,N_1573,N_2923);
nand U8763 (N_8763,N_4940,N_4256);
nor U8764 (N_8764,N_3486,N_2244);
nand U8765 (N_8765,N_3146,N_4280);
and U8766 (N_8766,N_4337,N_4620);
nor U8767 (N_8767,N_1179,N_4617);
nand U8768 (N_8768,N_2075,N_2972);
nand U8769 (N_8769,N_3234,N_3869);
nand U8770 (N_8770,N_2157,N_296);
or U8771 (N_8771,N_436,N_4663);
nor U8772 (N_8772,N_474,N_2552);
nor U8773 (N_8773,N_4628,N_4106);
nand U8774 (N_8774,N_3435,N_1426);
and U8775 (N_8775,N_4590,N_4586);
nor U8776 (N_8776,N_4587,N_859);
nor U8777 (N_8777,N_1308,N_4376);
and U8778 (N_8778,N_2825,N_415);
nor U8779 (N_8779,N_3743,N_3446);
nand U8780 (N_8780,N_1987,N_4479);
or U8781 (N_8781,N_1387,N_730);
nand U8782 (N_8782,N_2838,N_598);
and U8783 (N_8783,N_3140,N_2641);
or U8784 (N_8784,N_4776,N_2886);
nand U8785 (N_8785,N_2105,N_3082);
nand U8786 (N_8786,N_1321,N_2041);
or U8787 (N_8787,N_4445,N_2531);
nor U8788 (N_8788,N_4797,N_2527);
or U8789 (N_8789,N_4889,N_2543);
nor U8790 (N_8790,N_2993,N_2754);
or U8791 (N_8791,N_2703,N_1544);
or U8792 (N_8792,N_3600,N_938);
nand U8793 (N_8793,N_4946,N_2582);
nor U8794 (N_8794,N_3038,N_2337);
and U8795 (N_8795,N_2329,N_759);
nor U8796 (N_8796,N_1822,N_1953);
nand U8797 (N_8797,N_451,N_219);
nand U8798 (N_8798,N_4388,N_677);
or U8799 (N_8799,N_2993,N_1870);
xnor U8800 (N_8800,N_2346,N_4026);
nor U8801 (N_8801,N_2836,N_4440);
and U8802 (N_8802,N_1969,N_2631);
nand U8803 (N_8803,N_1519,N_434);
or U8804 (N_8804,N_4115,N_2309);
nand U8805 (N_8805,N_39,N_3634);
or U8806 (N_8806,N_4935,N_3746);
nor U8807 (N_8807,N_181,N_1728);
nor U8808 (N_8808,N_3952,N_1129);
nor U8809 (N_8809,N_4419,N_2306);
and U8810 (N_8810,N_2088,N_2594);
nor U8811 (N_8811,N_1959,N_1238);
or U8812 (N_8812,N_3848,N_2987);
nand U8813 (N_8813,N_3415,N_905);
nor U8814 (N_8814,N_204,N_2700);
and U8815 (N_8815,N_2407,N_3682);
and U8816 (N_8816,N_2813,N_1607);
nand U8817 (N_8817,N_4156,N_3837);
and U8818 (N_8818,N_3751,N_3482);
nor U8819 (N_8819,N_4167,N_2319);
nor U8820 (N_8820,N_4404,N_932);
nor U8821 (N_8821,N_3841,N_2711);
and U8822 (N_8822,N_2816,N_2102);
and U8823 (N_8823,N_2212,N_4095);
and U8824 (N_8824,N_4523,N_1586);
nand U8825 (N_8825,N_2352,N_4417);
and U8826 (N_8826,N_3325,N_1967);
nor U8827 (N_8827,N_573,N_1530);
and U8828 (N_8828,N_1936,N_2270);
or U8829 (N_8829,N_4023,N_3903);
nor U8830 (N_8830,N_2239,N_3980);
nor U8831 (N_8831,N_712,N_4043);
or U8832 (N_8832,N_3533,N_225);
nand U8833 (N_8833,N_113,N_4002);
nor U8834 (N_8834,N_4746,N_626);
or U8835 (N_8835,N_1172,N_4391);
nand U8836 (N_8836,N_2284,N_1087);
nand U8837 (N_8837,N_3421,N_327);
nand U8838 (N_8838,N_3019,N_3985);
and U8839 (N_8839,N_108,N_1411);
or U8840 (N_8840,N_3401,N_4945);
xor U8841 (N_8841,N_1257,N_2552);
or U8842 (N_8842,N_3303,N_2283);
nand U8843 (N_8843,N_2860,N_1094);
nor U8844 (N_8844,N_4399,N_1481);
nor U8845 (N_8845,N_2221,N_1798);
nand U8846 (N_8846,N_4913,N_2748);
nor U8847 (N_8847,N_3153,N_397);
or U8848 (N_8848,N_2785,N_2686);
and U8849 (N_8849,N_2899,N_1534);
and U8850 (N_8850,N_3183,N_11);
or U8851 (N_8851,N_3042,N_4294);
and U8852 (N_8852,N_1578,N_3693);
or U8853 (N_8853,N_1764,N_3707);
and U8854 (N_8854,N_2436,N_1716);
nand U8855 (N_8855,N_946,N_3175);
or U8856 (N_8856,N_4864,N_484);
nor U8857 (N_8857,N_2019,N_4530);
nand U8858 (N_8858,N_351,N_2163);
and U8859 (N_8859,N_283,N_3632);
or U8860 (N_8860,N_4920,N_4087);
and U8861 (N_8861,N_3952,N_3167);
and U8862 (N_8862,N_2528,N_3271);
nand U8863 (N_8863,N_1408,N_3830);
nor U8864 (N_8864,N_2578,N_2705);
nand U8865 (N_8865,N_1211,N_4760);
and U8866 (N_8866,N_951,N_4743);
nand U8867 (N_8867,N_4935,N_351);
nand U8868 (N_8868,N_4365,N_4759);
nand U8869 (N_8869,N_4234,N_2899);
or U8870 (N_8870,N_2379,N_2060);
or U8871 (N_8871,N_4701,N_428);
or U8872 (N_8872,N_1611,N_831);
nor U8873 (N_8873,N_1396,N_863);
xor U8874 (N_8874,N_4821,N_47);
or U8875 (N_8875,N_545,N_1897);
and U8876 (N_8876,N_1490,N_1009);
or U8877 (N_8877,N_1257,N_1153);
or U8878 (N_8878,N_1924,N_4611);
nor U8879 (N_8879,N_4159,N_4639);
nand U8880 (N_8880,N_4869,N_4407);
and U8881 (N_8881,N_4996,N_1449);
nand U8882 (N_8882,N_3315,N_2289);
and U8883 (N_8883,N_1250,N_3710);
nor U8884 (N_8884,N_4513,N_1136);
nor U8885 (N_8885,N_1020,N_4346);
or U8886 (N_8886,N_3794,N_1837);
and U8887 (N_8887,N_3268,N_1568);
and U8888 (N_8888,N_1133,N_4595);
nor U8889 (N_8889,N_1102,N_178);
nor U8890 (N_8890,N_1446,N_513);
xor U8891 (N_8891,N_341,N_1231);
or U8892 (N_8892,N_2241,N_1121);
xnor U8893 (N_8893,N_2292,N_791);
nor U8894 (N_8894,N_578,N_2580);
or U8895 (N_8895,N_4410,N_2683);
or U8896 (N_8896,N_4290,N_4772);
nor U8897 (N_8897,N_1086,N_2877);
nor U8898 (N_8898,N_359,N_2761);
and U8899 (N_8899,N_514,N_1135);
nor U8900 (N_8900,N_4181,N_4775);
nand U8901 (N_8901,N_3697,N_4203);
nor U8902 (N_8902,N_1793,N_2128);
and U8903 (N_8903,N_3514,N_4025);
nor U8904 (N_8904,N_2647,N_1420);
and U8905 (N_8905,N_3785,N_430);
or U8906 (N_8906,N_3645,N_4349);
nand U8907 (N_8907,N_4201,N_1038);
nor U8908 (N_8908,N_3255,N_4222);
or U8909 (N_8909,N_3134,N_3221);
nor U8910 (N_8910,N_3864,N_3824);
or U8911 (N_8911,N_1778,N_4779);
or U8912 (N_8912,N_4440,N_4026);
and U8913 (N_8913,N_4595,N_3366);
xnor U8914 (N_8914,N_3528,N_1979);
and U8915 (N_8915,N_2514,N_2309);
nor U8916 (N_8916,N_818,N_4801);
or U8917 (N_8917,N_4105,N_855);
nor U8918 (N_8918,N_3714,N_4009);
nand U8919 (N_8919,N_1302,N_4005);
nor U8920 (N_8920,N_2225,N_646);
nor U8921 (N_8921,N_2152,N_3860);
and U8922 (N_8922,N_1592,N_3781);
nor U8923 (N_8923,N_214,N_2884);
or U8924 (N_8924,N_1888,N_1715);
nor U8925 (N_8925,N_2643,N_1000);
nand U8926 (N_8926,N_3773,N_2436);
nand U8927 (N_8927,N_2157,N_3393);
nor U8928 (N_8928,N_1844,N_4388);
and U8929 (N_8929,N_4392,N_797);
or U8930 (N_8930,N_4782,N_1105);
nor U8931 (N_8931,N_4274,N_3326);
and U8932 (N_8932,N_4807,N_2639);
or U8933 (N_8933,N_3053,N_3987);
xor U8934 (N_8934,N_154,N_1529);
nor U8935 (N_8935,N_1616,N_3111);
nor U8936 (N_8936,N_1305,N_109);
and U8937 (N_8937,N_2192,N_2726);
nor U8938 (N_8938,N_1770,N_1487);
nand U8939 (N_8939,N_1574,N_1896);
nor U8940 (N_8940,N_526,N_2511);
nor U8941 (N_8941,N_660,N_1061);
nor U8942 (N_8942,N_3427,N_773);
and U8943 (N_8943,N_3080,N_2239);
xor U8944 (N_8944,N_371,N_3989);
or U8945 (N_8945,N_3854,N_445);
and U8946 (N_8946,N_3824,N_1985);
nand U8947 (N_8947,N_425,N_2119);
nand U8948 (N_8948,N_4373,N_4377);
xnor U8949 (N_8949,N_4617,N_5);
or U8950 (N_8950,N_4847,N_4581);
nand U8951 (N_8951,N_2728,N_4967);
or U8952 (N_8952,N_3505,N_1433);
and U8953 (N_8953,N_996,N_1581);
nor U8954 (N_8954,N_3040,N_4260);
xnor U8955 (N_8955,N_560,N_406);
nand U8956 (N_8956,N_3730,N_1465);
and U8957 (N_8957,N_1520,N_4993);
xor U8958 (N_8958,N_4501,N_3032);
or U8959 (N_8959,N_3235,N_3703);
and U8960 (N_8960,N_1607,N_720);
nor U8961 (N_8961,N_4649,N_905);
nor U8962 (N_8962,N_4919,N_828);
nor U8963 (N_8963,N_2645,N_394);
nor U8964 (N_8964,N_467,N_2575);
and U8965 (N_8965,N_8,N_1999);
and U8966 (N_8966,N_2880,N_4255);
nand U8967 (N_8967,N_2609,N_44);
nand U8968 (N_8968,N_522,N_2476);
nand U8969 (N_8969,N_1413,N_3920);
nand U8970 (N_8970,N_3145,N_3265);
nor U8971 (N_8971,N_1157,N_2212);
nand U8972 (N_8972,N_228,N_2959);
nor U8973 (N_8973,N_980,N_2902);
and U8974 (N_8974,N_3412,N_918);
nand U8975 (N_8975,N_741,N_3650);
nor U8976 (N_8976,N_857,N_4318);
or U8977 (N_8977,N_545,N_3954);
or U8978 (N_8978,N_394,N_2273);
and U8979 (N_8979,N_90,N_2198);
nand U8980 (N_8980,N_3494,N_4878);
and U8981 (N_8981,N_388,N_2149);
or U8982 (N_8982,N_537,N_4287);
or U8983 (N_8983,N_4482,N_3897);
xnor U8984 (N_8984,N_1724,N_1019);
nor U8985 (N_8985,N_2708,N_3755);
and U8986 (N_8986,N_1901,N_2895);
xnor U8987 (N_8987,N_3239,N_470);
nor U8988 (N_8988,N_1296,N_252);
nand U8989 (N_8989,N_79,N_1092);
or U8990 (N_8990,N_4493,N_634);
nand U8991 (N_8991,N_3572,N_1939);
nor U8992 (N_8992,N_3842,N_2632);
nand U8993 (N_8993,N_3084,N_1537);
nand U8994 (N_8994,N_1042,N_1256);
and U8995 (N_8995,N_1522,N_4303);
nand U8996 (N_8996,N_1912,N_4446);
nor U8997 (N_8997,N_3111,N_4516);
nand U8998 (N_8998,N_2860,N_2081);
or U8999 (N_8999,N_2133,N_424);
and U9000 (N_9000,N_4099,N_3693);
nand U9001 (N_9001,N_1876,N_2844);
or U9002 (N_9002,N_162,N_2122);
nand U9003 (N_9003,N_610,N_2968);
and U9004 (N_9004,N_884,N_3970);
or U9005 (N_9005,N_3404,N_2806);
nand U9006 (N_9006,N_1512,N_2391);
or U9007 (N_9007,N_3235,N_1304);
or U9008 (N_9008,N_3601,N_2976);
or U9009 (N_9009,N_3362,N_2019);
and U9010 (N_9010,N_2346,N_2499);
nand U9011 (N_9011,N_995,N_1636);
xnor U9012 (N_9012,N_1895,N_4850);
nand U9013 (N_9013,N_896,N_911);
nand U9014 (N_9014,N_271,N_4105);
and U9015 (N_9015,N_1618,N_3658);
and U9016 (N_9016,N_2420,N_2925);
nor U9017 (N_9017,N_1687,N_1399);
nand U9018 (N_9018,N_3580,N_679);
nor U9019 (N_9019,N_3586,N_4770);
nor U9020 (N_9020,N_2919,N_916);
nand U9021 (N_9021,N_3667,N_4248);
or U9022 (N_9022,N_3653,N_2483);
or U9023 (N_9023,N_1196,N_314);
nand U9024 (N_9024,N_589,N_1754);
and U9025 (N_9025,N_4602,N_2518);
and U9026 (N_9026,N_3121,N_3945);
and U9027 (N_9027,N_1492,N_382);
nor U9028 (N_9028,N_1933,N_4096);
or U9029 (N_9029,N_1350,N_749);
nor U9030 (N_9030,N_594,N_3311);
nor U9031 (N_9031,N_3781,N_4284);
nor U9032 (N_9032,N_1230,N_2534);
nor U9033 (N_9033,N_3548,N_3976);
or U9034 (N_9034,N_1356,N_1678);
nand U9035 (N_9035,N_4040,N_4815);
nor U9036 (N_9036,N_4895,N_1821);
or U9037 (N_9037,N_3461,N_2723);
and U9038 (N_9038,N_1657,N_1468);
or U9039 (N_9039,N_284,N_2280);
or U9040 (N_9040,N_321,N_4977);
or U9041 (N_9041,N_104,N_207);
nand U9042 (N_9042,N_58,N_184);
nand U9043 (N_9043,N_135,N_1077);
and U9044 (N_9044,N_1473,N_1320);
or U9045 (N_9045,N_2651,N_4844);
nand U9046 (N_9046,N_4131,N_4363);
and U9047 (N_9047,N_1236,N_1114);
nor U9048 (N_9048,N_4429,N_2282);
or U9049 (N_9049,N_2826,N_766);
and U9050 (N_9050,N_3992,N_1621);
nand U9051 (N_9051,N_1413,N_1471);
nor U9052 (N_9052,N_541,N_2369);
nand U9053 (N_9053,N_574,N_3400);
nand U9054 (N_9054,N_594,N_3096);
and U9055 (N_9055,N_1439,N_517);
and U9056 (N_9056,N_4761,N_4043);
nand U9057 (N_9057,N_1767,N_677);
or U9058 (N_9058,N_874,N_2590);
nand U9059 (N_9059,N_3000,N_2376);
or U9060 (N_9060,N_222,N_2753);
nand U9061 (N_9061,N_2810,N_3043);
nor U9062 (N_9062,N_3448,N_1439);
or U9063 (N_9063,N_851,N_2231);
and U9064 (N_9064,N_22,N_1445);
nor U9065 (N_9065,N_3867,N_3510);
or U9066 (N_9066,N_1221,N_1593);
nand U9067 (N_9067,N_3654,N_2042);
or U9068 (N_9068,N_1099,N_706);
or U9069 (N_9069,N_544,N_4958);
nand U9070 (N_9070,N_952,N_3167);
nor U9071 (N_9071,N_4826,N_19);
nand U9072 (N_9072,N_2310,N_2605);
or U9073 (N_9073,N_4474,N_3372);
xnor U9074 (N_9074,N_585,N_2630);
nor U9075 (N_9075,N_4364,N_1274);
nor U9076 (N_9076,N_4872,N_4688);
nand U9077 (N_9077,N_2631,N_3415);
nand U9078 (N_9078,N_3753,N_1694);
and U9079 (N_9079,N_1863,N_3460);
nand U9080 (N_9080,N_2702,N_162);
and U9081 (N_9081,N_4414,N_3649);
nand U9082 (N_9082,N_4743,N_2099);
nand U9083 (N_9083,N_2235,N_1282);
nand U9084 (N_9084,N_965,N_4164);
and U9085 (N_9085,N_317,N_1169);
or U9086 (N_9086,N_2465,N_1002);
nor U9087 (N_9087,N_3012,N_1538);
or U9088 (N_9088,N_4974,N_2940);
or U9089 (N_9089,N_401,N_1023);
and U9090 (N_9090,N_2148,N_4580);
or U9091 (N_9091,N_3071,N_4281);
and U9092 (N_9092,N_2990,N_4710);
or U9093 (N_9093,N_424,N_3182);
or U9094 (N_9094,N_4365,N_1690);
nor U9095 (N_9095,N_886,N_2020);
or U9096 (N_9096,N_3809,N_3892);
nand U9097 (N_9097,N_1610,N_2348);
and U9098 (N_9098,N_4156,N_2889);
and U9099 (N_9099,N_4948,N_2717);
nand U9100 (N_9100,N_1977,N_3796);
nor U9101 (N_9101,N_3768,N_1927);
and U9102 (N_9102,N_4798,N_318);
and U9103 (N_9103,N_3004,N_3129);
nand U9104 (N_9104,N_3647,N_1567);
or U9105 (N_9105,N_2664,N_4159);
and U9106 (N_9106,N_3441,N_1580);
and U9107 (N_9107,N_90,N_3039);
nand U9108 (N_9108,N_415,N_85);
and U9109 (N_9109,N_4880,N_4215);
nor U9110 (N_9110,N_4618,N_2075);
nor U9111 (N_9111,N_1976,N_81);
or U9112 (N_9112,N_988,N_676);
nand U9113 (N_9113,N_767,N_1826);
nand U9114 (N_9114,N_1808,N_2869);
nor U9115 (N_9115,N_4446,N_1344);
nor U9116 (N_9116,N_4695,N_1224);
nor U9117 (N_9117,N_4532,N_2898);
and U9118 (N_9118,N_3328,N_2155);
nor U9119 (N_9119,N_1824,N_2503);
nand U9120 (N_9120,N_4115,N_1875);
nand U9121 (N_9121,N_4307,N_888);
and U9122 (N_9122,N_576,N_1661);
nand U9123 (N_9123,N_1648,N_1747);
and U9124 (N_9124,N_1092,N_4371);
nor U9125 (N_9125,N_2045,N_1524);
nand U9126 (N_9126,N_2690,N_1947);
nor U9127 (N_9127,N_4605,N_3372);
and U9128 (N_9128,N_1059,N_1529);
xor U9129 (N_9129,N_383,N_865);
or U9130 (N_9130,N_1323,N_4812);
and U9131 (N_9131,N_4386,N_3221);
nor U9132 (N_9132,N_2462,N_2031);
nor U9133 (N_9133,N_485,N_2850);
nand U9134 (N_9134,N_99,N_286);
and U9135 (N_9135,N_2021,N_519);
nand U9136 (N_9136,N_4045,N_2788);
and U9137 (N_9137,N_4673,N_3645);
or U9138 (N_9138,N_264,N_935);
and U9139 (N_9139,N_3978,N_2102);
nor U9140 (N_9140,N_269,N_3027);
nor U9141 (N_9141,N_175,N_2122);
nand U9142 (N_9142,N_2514,N_4483);
nand U9143 (N_9143,N_1603,N_1262);
nand U9144 (N_9144,N_4021,N_1925);
or U9145 (N_9145,N_1539,N_4177);
nor U9146 (N_9146,N_112,N_873);
or U9147 (N_9147,N_3679,N_2326);
nand U9148 (N_9148,N_632,N_4840);
nand U9149 (N_9149,N_1927,N_4961);
and U9150 (N_9150,N_3408,N_3389);
nand U9151 (N_9151,N_865,N_4332);
nand U9152 (N_9152,N_84,N_650);
or U9153 (N_9153,N_419,N_939);
and U9154 (N_9154,N_2223,N_1342);
nor U9155 (N_9155,N_3433,N_1884);
nor U9156 (N_9156,N_2195,N_782);
and U9157 (N_9157,N_2437,N_1236);
and U9158 (N_9158,N_3487,N_684);
and U9159 (N_9159,N_2756,N_3266);
and U9160 (N_9160,N_2212,N_2633);
nand U9161 (N_9161,N_2536,N_1137);
and U9162 (N_9162,N_4010,N_1271);
nand U9163 (N_9163,N_1071,N_3092);
and U9164 (N_9164,N_2774,N_1039);
and U9165 (N_9165,N_3215,N_2052);
and U9166 (N_9166,N_1092,N_1142);
or U9167 (N_9167,N_72,N_478);
nor U9168 (N_9168,N_3785,N_2757);
or U9169 (N_9169,N_2583,N_3235);
nor U9170 (N_9170,N_3143,N_4884);
and U9171 (N_9171,N_3623,N_2718);
nor U9172 (N_9172,N_1925,N_2722);
and U9173 (N_9173,N_3803,N_1746);
nand U9174 (N_9174,N_4460,N_580);
nand U9175 (N_9175,N_650,N_35);
nand U9176 (N_9176,N_504,N_2589);
nand U9177 (N_9177,N_3287,N_3002);
nand U9178 (N_9178,N_1733,N_1083);
nand U9179 (N_9179,N_3614,N_26);
or U9180 (N_9180,N_4478,N_2542);
and U9181 (N_9181,N_1192,N_4030);
or U9182 (N_9182,N_1855,N_645);
or U9183 (N_9183,N_2344,N_2614);
and U9184 (N_9184,N_4676,N_257);
nor U9185 (N_9185,N_17,N_3785);
nor U9186 (N_9186,N_2142,N_2838);
nor U9187 (N_9187,N_1954,N_3481);
and U9188 (N_9188,N_560,N_1896);
nor U9189 (N_9189,N_1480,N_4504);
nand U9190 (N_9190,N_4228,N_1113);
nor U9191 (N_9191,N_3384,N_349);
nor U9192 (N_9192,N_3058,N_1821);
or U9193 (N_9193,N_1231,N_4697);
and U9194 (N_9194,N_90,N_2847);
or U9195 (N_9195,N_4130,N_345);
nand U9196 (N_9196,N_1690,N_4561);
nor U9197 (N_9197,N_4993,N_3352);
or U9198 (N_9198,N_472,N_3284);
nand U9199 (N_9199,N_2972,N_3557);
or U9200 (N_9200,N_4365,N_1033);
or U9201 (N_9201,N_741,N_1938);
nor U9202 (N_9202,N_4325,N_1114);
nor U9203 (N_9203,N_3822,N_1412);
and U9204 (N_9204,N_2790,N_121);
nor U9205 (N_9205,N_258,N_346);
nand U9206 (N_9206,N_1387,N_4699);
and U9207 (N_9207,N_3887,N_2300);
nor U9208 (N_9208,N_934,N_13);
nand U9209 (N_9209,N_1394,N_2329);
nor U9210 (N_9210,N_1475,N_4043);
nand U9211 (N_9211,N_47,N_3076);
and U9212 (N_9212,N_3828,N_3746);
nand U9213 (N_9213,N_2340,N_3401);
or U9214 (N_9214,N_2317,N_3115);
or U9215 (N_9215,N_4161,N_3173);
or U9216 (N_9216,N_4197,N_17);
or U9217 (N_9217,N_2391,N_4220);
nand U9218 (N_9218,N_4203,N_3048);
or U9219 (N_9219,N_1895,N_4739);
nor U9220 (N_9220,N_4425,N_4510);
nand U9221 (N_9221,N_3617,N_3039);
or U9222 (N_9222,N_466,N_4468);
or U9223 (N_9223,N_1317,N_1831);
nand U9224 (N_9224,N_2560,N_3366);
or U9225 (N_9225,N_3831,N_3447);
nor U9226 (N_9226,N_322,N_4701);
and U9227 (N_9227,N_4976,N_4209);
or U9228 (N_9228,N_1059,N_2631);
and U9229 (N_9229,N_3689,N_4052);
and U9230 (N_9230,N_4225,N_195);
nor U9231 (N_9231,N_4663,N_413);
nor U9232 (N_9232,N_575,N_4681);
nand U9233 (N_9233,N_331,N_712);
or U9234 (N_9234,N_2006,N_2086);
nand U9235 (N_9235,N_4172,N_2343);
nand U9236 (N_9236,N_3004,N_3051);
xnor U9237 (N_9237,N_3643,N_3397);
or U9238 (N_9238,N_537,N_4106);
nor U9239 (N_9239,N_3377,N_3072);
or U9240 (N_9240,N_3797,N_4020);
or U9241 (N_9241,N_2520,N_2792);
and U9242 (N_9242,N_4793,N_81);
and U9243 (N_9243,N_921,N_2349);
or U9244 (N_9244,N_3285,N_3692);
nand U9245 (N_9245,N_3941,N_2053);
or U9246 (N_9246,N_16,N_3014);
nand U9247 (N_9247,N_936,N_2590);
nand U9248 (N_9248,N_4097,N_1853);
and U9249 (N_9249,N_3269,N_2840);
nor U9250 (N_9250,N_4332,N_2196);
nand U9251 (N_9251,N_258,N_312);
nor U9252 (N_9252,N_1850,N_379);
nor U9253 (N_9253,N_583,N_2814);
or U9254 (N_9254,N_3403,N_1972);
or U9255 (N_9255,N_1768,N_825);
nand U9256 (N_9256,N_2453,N_4868);
nand U9257 (N_9257,N_613,N_486);
nand U9258 (N_9258,N_2029,N_1230);
or U9259 (N_9259,N_198,N_3302);
nand U9260 (N_9260,N_3870,N_997);
nor U9261 (N_9261,N_3872,N_715);
nor U9262 (N_9262,N_2282,N_1509);
or U9263 (N_9263,N_3505,N_1345);
or U9264 (N_9264,N_4585,N_3626);
nand U9265 (N_9265,N_4458,N_1322);
or U9266 (N_9266,N_4234,N_4504);
or U9267 (N_9267,N_3933,N_1506);
or U9268 (N_9268,N_1705,N_1687);
nor U9269 (N_9269,N_1650,N_1126);
nand U9270 (N_9270,N_4182,N_1450);
nand U9271 (N_9271,N_2910,N_1890);
xnor U9272 (N_9272,N_901,N_4650);
xor U9273 (N_9273,N_2978,N_3168);
xnor U9274 (N_9274,N_3864,N_375);
and U9275 (N_9275,N_4001,N_206);
and U9276 (N_9276,N_2497,N_2158);
nand U9277 (N_9277,N_3668,N_1621);
or U9278 (N_9278,N_2899,N_1332);
or U9279 (N_9279,N_4650,N_3189);
and U9280 (N_9280,N_600,N_1992);
or U9281 (N_9281,N_2178,N_4102);
nand U9282 (N_9282,N_561,N_1464);
nand U9283 (N_9283,N_2928,N_1739);
nand U9284 (N_9284,N_3744,N_1098);
and U9285 (N_9285,N_3632,N_2842);
and U9286 (N_9286,N_1050,N_4649);
nor U9287 (N_9287,N_2402,N_2285);
and U9288 (N_9288,N_202,N_481);
or U9289 (N_9289,N_3019,N_3415);
nor U9290 (N_9290,N_408,N_1763);
and U9291 (N_9291,N_2778,N_4243);
and U9292 (N_9292,N_2448,N_3572);
nor U9293 (N_9293,N_1706,N_2383);
nand U9294 (N_9294,N_3760,N_2783);
nor U9295 (N_9295,N_2165,N_3060);
and U9296 (N_9296,N_3394,N_4804);
and U9297 (N_9297,N_4327,N_4491);
nor U9298 (N_9298,N_3547,N_3390);
or U9299 (N_9299,N_4498,N_4394);
nor U9300 (N_9300,N_2330,N_1976);
and U9301 (N_9301,N_930,N_4568);
nand U9302 (N_9302,N_996,N_1227);
and U9303 (N_9303,N_794,N_3291);
nand U9304 (N_9304,N_4405,N_4734);
nor U9305 (N_9305,N_4934,N_2871);
and U9306 (N_9306,N_2837,N_124);
or U9307 (N_9307,N_3677,N_1266);
or U9308 (N_9308,N_4376,N_566);
nor U9309 (N_9309,N_2122,N_1849);
nor U9310 (N_9310,N_1211,N_12);
and U9311 (N_9311,N_4594,N_3809);
and U9312 (N_9312,N_1586,N_2766);
xor U9313 (N_9313,N_1655,N_2386);
and U9314 (N_9314,N_1190,N_2157);
and U9315 (N_9315,N_4522,N_3209);
or U9316 (N_9316,N_1792,N_886);
nand U9317 (N_9317,N_4566,N_911);
nand U9318 (N_9318,N_1470,N_1036);
nor U9319 (N_9319,N_4902,N_2865);
or U9320 (N_9320,N_819,N_133);
nand U9321 (N_9321,N_3886,N_279);
nor U9322 (N_9322,N_4856,N_3224);
or U9323 (N_9323,N_3544,N_3589);
or U9324 (N_9324,N_3932,N_3807);
and U9325 (N_9325,N_3337,N_27);
nand U9326 (N_9326,N_849,N_1398);
nand U9327 (N_9327,N_14,N_1820);
nor U9328 (N_9328,N_3884,N_488);
or U9329 (N_9329,N_2424,N_1579);
and U9330 (N_9330,N_4678,N_4065);
and U9331 (N_9331,N_4180,N_3848);
and U9332 (N_9332,N_4386,N_2889);
or U9333 (N_9333,N_4945,N_764);
nor U9334 (N_9334,N_970,N_3851);
and U9335 (N_9335,N_307,N_542);
nor U9336 (N_9336,N_3182,N_1385);
nand U9337 (N_9337,N_1287,N_3191);
nor U9338 (N_9338,N_2670,N_2248);
nand U9339 (N_9339,N_2951,N_1544);
and U9340 (N_9340,N_2054,N_4963);
nand U9341 (N_9341,N_3289,N_3878);
or U9342 (N_9342,N_3009,N_2469);
nor U9343 (N_9343,N_2516,N_1236);
and U9344 (N_9344,N_1845,N_1077);
or U9345 (N_9345,N_219,N_1267);
nor U9346 (N_9346,N_1344,N_1763);
nor U9347 (N_9347,N_2440,N_4025);
or U9348 (N_9348,N_1274,N_2430);
nand U9349 (N_9349,N_3963,N_222);
nor U9350 (N_9350,N_1194,N_1843);
xor U9351 (N_9351,N_4969,N_4708);
nand U9352 (N_9352,N_2628,N_2059);
nand U9353 (N_9353,N_207,N_3705);
and U9354 (N_9354,N_590,N_2937);
nor U9355 (N_9355,N_2335,N_592);
nand U9356 (N_9356,N_2645,N_1816);
xor U9357 (N_9357,N_832,N_3549);
nand U9358 (N_9358,N_1339,N_122);
and U9359 (N_9359,N_3991,N_3729);
nor U9360 (N_9360,N_2940,N_4781);
nor U9361 (N_9361,N_2379,N_1456);
nor U9362 (N_9362,N_3234,N_2879);
or U9363 (N_9363,N_3641,N_2779);
nor U9364 (N_9364,N_1006,N_2642);
nor U9365 (N_9365,N_579,N_3187);
nor U9366 (N_9366,N_11,N_4353);
and U9367 (N_9367,N_3265,N_767);
and U9368 (N_9368,N_2490,N_4247);
and U9369 (N_9369,N_3748,N_4753);
and U9370 (N_9370,N_197,N_2000);
or U9371 (N_9371,N_2124,N_1979);
and U9372 (N_9372,N_1410,N_1974);
and U9373 (N_9373,N_1541,N_1318);
nand U9374 (N_9374,N_1358,N_1321);
nand U9375 (N_9375,N_3319,N_1988);
nand U9376 (N_9376,N_2443,N_4172);
or U9377 (N_9377,N_2187,N_1494);
nand U9378 (N_9378,N_3536,N_1359);
nor U9379 (N_9379,N_513,N_1818);
nor U9380 (N_9380,N_4719,N_42);
nor U9381 (N_9381,N_4707,N_2055);
or U9382 (N_9382,N_1557,N_3640);
nor U9383 (N_9383,N_4037,N_709);
nor U9384 (N_9384,N_320,N_3435);
or U9385 (N_9385,N_743,N_545);
or U9386 (N_9386,N_1068,N_4682);
nand U9387 (N_9387,N_668,N_2609);
nor U9388 (N_9388,N_4337,N_3442);
nand U9389 (N_9389,N_610,N_122);
and U9390 (N_9390,N_1386,N_57);
nand U9391 (N_9391,N_4529,N_931);
nand U9392 (N_9392,N_4690,N_2289);
or U9393 (N_9393,N_3395,N_4116);
nand U9394 (N_9394,N_618,N_4986);
and U9395 (N_9395,N_4094,N_604);
nor U9396 (N_9396,N_4961,N_618);
nand U9397 (N_9397,N_3547,N_1131);
nand U9398 (N_9398,N_332,N_1234);
nor U9399 (N_9399,N_3157,N_1899);
nor U9400 (N_9400,N_729,N_3475);
or U9401 (N_9401,N_4557,N_1316);
and U9402 (N_9402,N_3011,N_912);
and U9403 (N_9403,N_2411,N_4930);
nand U9404 (N_9404,N_3495,N_1951);
nand U9405 (N_9405,N_1040,N_4383);
nand U9406 (N_9406,N_1422,N_2210);
or U9407 (N_9407,N_4558,N_2143);
nand U9408 (N_9408,N_4842,N_2197);
nor U9409 (N_9409,N_1053,N_4581);
nand U9410 (N_9410,N_3936,N_639);
nand U9411 (N_9411,N_1606,N_4548);
nor U9412 (N_9412,N_655,N_2448);
nand U9413 (N_9413,N_2709,N_82);
nand U9414 (N_9414,N_2913,N_2597);
nor U9415 (N_9415,N_4481,N_2592);
or U9416 (N_9416,N_2843,N_2842);
nand U9417 (N_9417,N_4247,N_4743);
or U9418 (N_9418,N_3484,N_3334);
and U9419 (N_9419,N_3939,N_4107);
nor U9420 (N_9420,N_3304,N_3070);
nand U9421 (N_9421,N_4380,N_3821);
or U9422 (N_9422,N_4028,N_681);
nand U9423 (N_9423,N_1875,N_3997);
and U9424 (N_9424,N_4233,N_218);
and U9425 (N_9425,N_1308,N_3551);
and U9426 (N_9426,N_1656,N_1221);
nor U9427 (N_9427,N_1426,N_3110);
nor U9428 (N_9428,N_2853,N_3068);
nand U9429 (N_9429,N_1759,N_4513);
and U9430 (N_9430,N_968,N_3958);
nand U9431 (N_9431,N_3622,N_4145);
nand U9432 (N_9432,N_3407,N_4359);
or U9433 (N_9433,N_852,N_3704);
nor U9434 (N_9434,N_4401,N_1282);
and U9435 (N_9435,N_372,N_180);
or U9436 (N_9436,N_1696,N_2809);
nor U9437 (N_9437,N_2527,N_1251);
nor U9438 (N_9438,N_838,N_3567);
or U9439 (N_9439,N_1163,N_1863);
or U9440 (N_9440,N_515,N_2656);
nand U9441 (N_9441,N_3777,N_4963);
nor U9442 (N_9442,N_4002,N_237);
nand U9443 (N_9443,N_863,N_4885);
or U9444 (N_9444,N_2954,N_1527);
or U9445 (N_9445,N_238,N_3311);
nor U9446 (N_9446,N_1255,N_3681);
nand U9447 (N_9447,N_2895,N_3564);
nor U9448 (N_9448,N_565,N_3474);
nand U9449 (N_9449,N_492,N_4365);
nor U9450 (N_9450,N_4209,N_1907);
or U9451 (N_9451,N_2508,N_2956);
and U9452 (N_9452,N_4525,N_708);
nand U9453 (N_9453,N_3561,N_4644);
and U9454 (N_9454,N_651,N_4835);
nand U9455 (N_9455,N_3460,N_3981);
or U9456 (N_9456,N_1539,N_1771);
nor U9457 (N_9457,N_2673,N_1546);
xnor U9458 (N_9458,N_2829,N_3672);
and U9459 (N_9459,N_4084,N_4427);
nand U9460 (N_9460,N_3283,N_1681);
nand U9461 (N_9461,N_4666,N_3024);
nor U9462 (N_9462,N_4029,N_416);
nor U9463 (N_9463,N_158,N_363);
nand U9464 (N_9464,N_4037,N_4231);
and U9465 (N_9465,N_1380,N_4809);
nor U9466 (N_9466,N_634,N_3848);
nor U9467 (N_9467,N_4251,N_2395);
nor U9468 (N_9468,N_4563,N_4507);
or U9469 (N_9469,N_355,N_2936);
and U9470 (N_9470,N_2686,N_4408);
nor U9471 (N_9471,N_3547,N_1622);
or U9472 (N_9472,N_4815,N_1821);
or U9473 (N_9473,N_4606,N_1170);
nand U9474 (N_9474,N_646,N_2567);
nand U9475 (N_9475,N_2896,N_3548);
nand U9476 (N_9476,N_4973,N_1588);
nor U9477 (N_9477,N_785,N_659);
and U9478 (N_9478,N_3028,N_3367);
nand U9479 (N_9479,N_3045,N_4551);
nand U9480 (N_9480,N_3390,N_1309);
nand U9481 (N_9481,N_3863,N_531);
nor U9482 (N_9482,N_4015,N_1528);
and U9483 (N_9483,N_2783,N_1516);
nand U9484 (N_9484,N_3149,N_3157);
or U9485 (N_9485,N_994,N_3907);
or U9486 (N_9486,N_4899,N_3975);
or U9487 (N_9487,N_432,N_3381);
and U9488 (N_9488,N_4712,N_1200);
nand U9489 (N_9489,N_4295,N_2882);
and U9490 (N_9490,N_504,N_382);
or U9491 (N_9491,N_3303,N_704);
or U9492 (N_9492,N_575,N_2078);
nor U9493 (N_9493,N_2592,N_2780);
and U9494 (N_9494,N_1110,N_545);
or U9495 (N_9495,N_4031,N_2666);
and U9496 (N_9496,N_1755,N_4379);
nand U9497 (N_9497,N_2353,N_3352);
nor U9498 (N_9498,N_1249,N_1467);
and U9499 (N_9499,N_3435,N_3743);
xor U9500 (N_9500,N_3285,N_4744);
nand U9501 (N_9501,N_1117,N_2294);
and U9502 (N_9502,N_4952,N_359);
and U9503 (N_9503,N_4233,N_3201);
or U9504 (N_9504,N_137,N_1712);
or U9505 (N_9505,N_2586,N_1904);
nand U9506 (N_9506,N_3655,N_2593);
nor U9507 (N_9507,N_3989,N_1912);
and U9508 (N_9508,N_345,N_3101);
and U9509 (N_9509,N_2178,N_4200);
nor U9510 (N_9510,N_1146,N_1211);
nand U9511 (N_9511,N_768,N_3891);
or U9512 (N_9512,N_4364,N_1118);
and U9513 (N_9513,N_1009,N_3928);
nor U9514 (N_9514,N_4597,N_3092);
or U9515 (N_9515,N_3079,N_4259);
and U9516 (N_9516,N_1055,N_3602);
and U9517 (N_9517,N_1815,N_324);
and U9518 (N_9518,N_2592,N_4861);
and U9519 (N_9519,N_91,N_322);
and U9520 (N_9520,N_3408,N_3883);
nor U9521 (N_9521,N_3998,N_3108);
and U9522 (N_9522,N_3095,N_4671);
and U9523 (N_9523,N_1620,N_2118);
nor U9524 (N_9524,N_672,N_2994);
or U9525 (N_9525,N_2978,N_4113);
nand U9526 (N_9526,N_1036,N_4574);
nand U9527 (N_9527,N_3955,N_579);
and U9528 (N_9528,N_606,N_2217);
or U9529 (N_9529,N_719,N_917);
and U9530 (N_9530,N_3423,N_3111);
and U9531 (N_9531,N_4564,N_4108);
nand U9532 (N_9532,N_3368,N_277);
nor U9533 (N_9533,N_2986,N_3762);
xnor U9534 (N_9534,N_2852,N_2465);
nand U9535 (N_9535,N_2653,N_4058);
nand U9536 (N_9536,N_1054,N_1546);
nand U9537 (N_9537,N_972,N_2873);
or U9538 (N_9538,N_3101,N_2487);
or U9539 (N_9539,N_3895,N_640);
and U9540 (N_9540,N_85,N_4663);
and U9541 (N_9541,N_3517,N_86);
nor U9542 (N_9542,N_4845,N_4664);
or U9543 (N_9543,N_3046,N_1177);
nor U9544 (N_9544,N_657,N_4902);
nor U9545 (N_9545,N_2512,N_4898);
nand U9546 (N_9546,N_2926,N_4728);
and U9547 (N_9547,N_3387,N_2886);
and U9548 (N_9548,N_4233,N_414);
and U9549 (N_9549,N_3967,N_3948);
nand U9550 (N_9550,N_4623,N_3870);
nor U9551 (N_9551,N_20,N_913);
nor U9552 (N_9552,N_4984,N_3219);
nor U9553 (N_9553,N_926,N_4473);
nand U9554 (N_9554,N_248,N_2095);
and U9555 (N_9555,N_4079,N_4141);
and U9556 (N_9556,N_48,N_2677);
and U9557 (N_9557,N_1386,N_2803);
nor U9558 (N_9558,N_187,N_151);
or U9559 (N_9559,N_3745,N_3197);
or U9560 (N_9560,N_4197,N_873);
nor U9561 (N_9561,N_558,N_4564);
nor U9562 (N_9562,N_3466,N_368);
xor U9563 (N_9563,N_4651,N_1401);
and U9564 (N_9564,N_4751,N_3091);
or U9565 (N_9565,N_518,N_446);
or U9566 (N_9566,N_4226,N_1558);
nand U9567 (N_9567,N_1384,N_2517);
and U9568 (N_9568,N_3444,N_1077);
nand U9569 (N_9569,N_4110,N_2555);
nand U9570 (N_9570,N_3179,N_2645);
and U9571 (N_9571,N_2399,N_1766);
nand U9572 (N_9572,N_1931,N_526);
and U9573 (N_9573,N_2662,N_3571);
and U9574 (N_9574,N_2243,N_4839);
nor U9575 (N_9575,N_4509,N_1371);
or U9576 (N_9576,N_1457,N_1166);
nor U9577 (N_9577,N_824,N_3417);
or U9578 (N_9578,N_1558,N_2357);
nand U9579 (N_9579,N_3162,N_145);
xor U9580 (N_9580,N_3763,N_552);
nand U9581 (N_9581,N_3886,N_4995);
and U9582 (N_9582,N_1030,N_2377);
and U9583 (N_9583,N_470,N_3302);
or U9584 (N_9584,N_194,N_3272);
xor U9585 (N_9585,N_1755,N_2052);
nand U9586 (N_9586,N_181,N_1347);
or U9587 (N_9587,N_3407,N_2251);
nor U9588 (N_9588,N_2501,N_166);
and U9589 (N_9589,N_248,N_2307);
or U9590 (N_9590,N_4994,N_2929);
or U9591 (N_9591,N_1957,N_3326);
and U9592 (N_9592,N_1263,N_2626);
nor U9593 (N_9593,N_1993,N_17);
nand U9594 (N_9594,N_3854,N_776);
or U9595 (N_9595,N_3607,N_1172);
nor U9596 (N_9596,N_3709,N_4431);
nor U9597 (N_9597,N_4091,N_3311);
or U9598 (N_9598,N_4351,N_2864);
or U9599 (N_9599,N_544,N_4093);
and U9600 (N_9600,N_3271,N_3422);
or U9601 (N_9601,N_2014,N_2268);
nand U9602 (N_9602,N_4761,N_2012);
and U9603 (N_9603,N_1065,N_4473);
nand U9604 (N_9604,N_927,N_319);
xnor U9605 (N_9605,N_1571,N_2320);
or U9606 (N_9606,N_2756,N_2962);
or U9607 (N_9607,N_3193,N_4100);
nand U9608 (N_9608,N_2847,N_4335);
nor U9609 (N_9609,N_4482,N_2985);
or U9610 (N_9610,N_2607,N_2506);
nand U9611 (N_9611,N_2561,N_2336);
nor U9612 (N_9612,N_1264,N_323);
or U9613 (N_9613,N_1885,N_2919);
nand U9614 (N_9614,N_4061,N_2924);
nor U9615 (N_9615,N_442,N_4683);
and U9616 (N_9616,N_4642,N_4623);
nand U9617 (N_9617,N_2132,N_2651);
nor U9618 (N_9618,N_4395,N_67);
nor U9619 (N_9619,N_597,N_3858);
or U9620 (N_9620,N_2956,N_904);
and U9621 (N_9621,N_2717,N_359);
nor U9622 (N_9622,N_4853,N_412);
nand U9623 (N_9623,N_588,N_1970);
nor U9624 (N_9624,N_580,N_2467);
or U9625 (N_9625,N_1025,N_97);
or U9626 (N_9626,N_1854,N_3899);
or U9627 (N_9627,N_1830,N_2512);
nor U9628 (N_9628,N_3594,N_1418);
and U9629 (N_9629,N_1911,N_3941);
nor U9630 (N_9630,N_3917,N_3224);
and U9631 (N_9631,N_2541,N_653);
xnor U9632 (N_9632,N_198,N_4040);
or U9633 (N_9633,N_4009,N_69);
nor U9634 (N_9634,N_2602,N_2610);
or U9635 (N_9635,N_3037,N_4278);
and U9636 (N_9636,N_134,N_4950);
nand U9637 (N_9637,N_2773,N_1270);
nand U9638 (N_9638,N_3019,N_1743);
or U9639 (N_9639,N_36,N_2248);
and U9640 (N_9640,N_3687,N_2332);
or U9641 (N_9641,N_1042,N_1478);
nand U9642 (N_9642,N_1541,N_1254);
nand U9643 (N_9643,N_56,N_2736);
nand U9644 (N_9644,N_4762,N_2546);
nor U9645 (N_9645,N_4127,N_4241);
and U9646 (N_9646,N_2753,N_4241);
nand U9647 (N_9647,N_370,N_777);
nand U9648 (N_9648,N_1336,N_2735);
and U9649 (N_9649,N_1333,N_3994);
nand U9650 (N_9650,N_3123,N_393);
or U9651 (N_9651,N_2112,N_4119);
nand U9652 (N_9652,N_4736,N_573);
or U9653 (N_9653,N_1866,N_1129);
or U9654 (N_9654,N_3803,N_4934);
nor U9655 (N_9655,N_980,N_1384);
nand U9656 (N_9656,N_207,N_2283);
nor U9657 (N_9657,N_704,N_1);
and U9658 (N_9658,N_4150,N_1920);
nand U9659 (N_9659,N_4630,N_2974);
and U9660 (N_9660,N_3615,N_1125);
nor U9661 (N_9661,N_4992,N_699);
and U9662 (N_9662,N_3249,N_2722);
nand U9663 (N_9663,N_3734,N_4982);
nor U9664 (N_9664,N_1126,N_1728);
nor U9665 (N_9665,N_2962,N_2520);
or U9666 (N_9666,N_2203,N_3014);
or U9667 (N_9667,N_107,N_2443);
xnor U9668 (N_9668,N_2703,N_2095);
or U9669 (N_9669,N_4106,N_1418);
or U9670 (N_9670,N_3252,N_441);
nor U9671 (N_9671,N_2561,N_4874);
and U9672 (N_9672,N_3376,N_3913);
nand U9673 (N_9673,N_4498,N_4118);
or U9674 (N_9674,N_1053,N_1218);
and U9675 (N_9675,N_2314,N_1705);
nand U9676 (N_9676,N_4478,N_754);
or U9677 (N_9677,N_2223,N_3641);
nand U9678 (N_9678,N_557,N_2472);
and U9679 (N_9679,N_1087,N_4040);
nand U9680 (N_9680,N_2108,N_43);
nor U9681 (N_9681,N_2336,N_3116);
nor U9682 (N_9682,N_4653,N_3915);
or U9683 (N_9683,N_1321,N_661);
nand U9684 (N_9684,N_990,N_329);
nand U9685 (N_9685,N_2626,N_54);
nand U9686 (N_9686,N_3513,N_3227);
nand U9687 (N_9687,N_562,N_3685);
or U9688 (N_9688,N_2225,N_3641);
nor U9689 (N_9689,N_1611,N_4465);
nor U9690 (N_9690,N_1529,N_4763);
or U9691 (N_9691,N_2571,N_4615);
and U9692 (N_9692,N_3282,N_2468);
nor U9693 (N_9693,N_1375,N_1904);
or U9694 (N_9694,N_3687,N_336);
and U9695 (N_9695,N_572,N_2490);
or U9696 (N_9696,N_3198,N_2485);
nand U9697 (N_9697,N_4107,N_4116);
nand U9698 (N_9698,N_2501,N_425);
nor U9699 (N_9699,N_1149,N_2594);
nand U9700 (N_9700,N_4505,N_3550);
nor U9701 (N_9701,N_3460,N_2841);
and U9702 (N_9702,N_3,N_3551);
nor U9703 (N_9703,N_1826,N_4200);
or U9704 (N_9704,N_2598,N_2411);
and U9705 (N_9705,N_2705,N_2523);
and U9706 (N_9706,N_1241,N_3333);
and U9707 (N_9707,N_838,N_2527);
and U9708 (N_9708,N_1867,N_3097);
and U9709 (N_9709,N_590,N_2664);
xor U9710 (N_9710,N_4273,N_786);
and U9711 (N_9711,N_1023,N_4599);
nand U9712 (N_9712,N_3553,N_2576);
or U9713 (N_9713,N_4615,N_4483);
xor U9714 (N_9714,N_2087,N_3673);
nor U9715 (N_9715,N_249,N_3214);
or U9716 (N_9716,N_4575,N_4191);
and U9717 (N_9717,N_4198,N_2098);
or U9718 (N_9718,N_1181,N_3339);
nor U9719 (N_9719,N_3346,N_1146);
nor U9720 (N_9720,N_4952,N_3025);
and U9721 (N_9721,N_1366,N_1885);
nor U9722 (N_9722,N_1102,N_524);
nand U9723 (N_9723,N_3685,N_1610);
and U9724 (N_9724,N_3848,N_2765);
xor U9725 (N_9725,N_3505,N_4753);
or U9726 (N_9726,N_3137,N_4554);
nand U9727 (N_9727,N_385,N_4680);
and U9728 (N_9728,N_2772,N_5);
or U9729 (N_9729,N_199,N_4071);
or U9730 (N_9730,N_547,N_4279);
and U9731 (N_9731,N_1003,N_4663);
and U9732 (N_9732,N_2393,N_2033);
or U9733 (N_9733,N_4517,N_3472);
nand U9734 (N_9734,N_4629,N_363);
and U9735 (N_9735,N_769,N_772);
and U9736 (N_9736,N_1821,N_314);
nor U9737 (N_9737,N_2319,N_4059);
or U9738 (N_9738,N_3226,N_1428);
nand U9739 (N_9739,N_4818,N_4701);
or U9740 (N_9740,N_4317,N_3174);
nor U9741 (N_9741,N_4213,N_3848);
and U9742 (N_9742,N_802,N_4228);
nor U9743 (N_9743,N_1603,N_3059);
nor U9744 (N_9744,N_1662,N_695);
and U9745 (N_9745,N_2309,N_4555);
and U9746 (N_9746,N_3336,N_1440);
nand U9747 (N_9747,N_4921,N_880);
nand U9748 (N_9748,N_2525,N_3171);
and U9749 (N_9749,N_1937,N_1274);
or U9750 (N_9750,N_291,N_3532);
nand U9751 (N_9751,N_1350,N_805);
or U9752 (N_9752,N_1563,N_152);
nor U9753 (N_9753,N_2213,N_1059);
nand U9754 (N_9754,N_1885,N_1074);
nor U9755 (N_9755,N_2564,N_3510);
nand U9756 (N_9756,N_1131,N_3075);
nor U9757 (N_9757,N_2698,N_2764);
nor U9758 (N_9758,N_4634,N_802);
nand U9759 (N_9759,N_1651,N_3563);
nor U9760 (N_9760,N_4685,N_1514);
nor U9761 (N_9761,N_1017,N_3245);
nor U9762 (N_9762,N_304,N_606);
or U9763 (N_9763,N_2181,N_3688);
nand U9764 (N_9764,N_2405,N_3715);
nor U9765 (N_9765,N_198,N_1490);
xnor U9766 (N_9766,N_4312,N_596);
or U9767 (N_9767,N_2626,N_15);
xnor U9768 (N_9768,N_1866,N_1536);
nor U9769 (N_9769,N_1720,N_4952);
and U9770 (N_9770,N_714,N_2146);
or U9771 (N_9771,N_4831,N_1757);
nand U9772 (N_9772,N_1429,N_1765);
nor U9773 (N_9773,N_1012,N_1186);
xor U9774 (N_9774,N_3306,N_4295);
xor U9775 (N_9775,N_1914,N_2976);
nand U9776 (N_9776,N_1271,N_4143);
or U9777 (N_9777,N_2574,N_3474);
or U9778 (N_9778,N_1705,N_1749);
or U9779 (N_9779,N_4525,N_2054);
nand U9780 (N_9780,N_86,N_3420);
nor U9781 (N_9781,N_792,N_615);
and U9782 (N_9782,N_4327,N_2982);
nor U9783 (N_9783,N_1651,N_3475);
nand U9784 (N_9784,N_1950,N_1017);
nand U9785 (N_9785,N_119,N_4507);
nor U9786 (N_9786,N_3630,N_375);
and U9787 (N_9787,N_3600,N_2652);
nand U9788 (N_9788,N_2929,N_3759);
or U9789 (N_9789,N_4611,N_4278);
nor U9790 (N_9790,N_989,N_1962);
or U9791 (N_9791,N_4685,N_2491);
and U9792 (N_9792,N_115,N_4529);
and U9793 (N_9793,N_2419,N_3245);
and U9794 (N_9794,N_4134,N_415);
nor U9795 (N_9795,N_301,N_2270);
nand U9796 (N_9796,N_3493,N_2603);
and U9797 (N_9797,N_1542,N_439);
nor U9798 (N_9798,N_1442,N_3549);
or U9799 (N_9799,N_1094,N_370);
and U9800 (N_9800,N_4824,N_4204);
nor U9801 (N_9801,N_4192,N_4305);
and U9802 (N_9802,N_3692,N_4209);
or U9803 (N_9803,N_586,N_2438);
and U9804 (N_9804,N_4956,N_422);
or U9805 (N_9805,N_4913,N_371);
and U9806 (N_9806,N_799,N_607);
nor U9807 (N_9807,N_4651,N_3751);
nand U9808 (N_9808,N_3068,N_4841);
and U9809 (N_9809,N_575,N_1813);
and U9810 (N_9810,N_2718,N_3109);
nor U9811 (N_9811,N_2135,N_2687);
nand U9812 (N_9812,N_84,N_1226);
nand U9813 (N_9813,N_4107,N_3268);
or U9814 (N_9814,N_605,N_2320);
and U9815 (N_9815,N_4151,N_586);
xor U9816 (N_9816,N_1436,N_2258);
nand U9817 (N_9817,N_4572,N_1781);
nand U9818 (N_9818,N_1175,N_1125);
nand U9819 (N_9819,N_1227,N_130);
or U9820 (N_9820,N_45,N_4680);
nor U9821 (N_9821,N_4065,N_4098);
nor U9822 (N_9822,N_869,N_67);
nand U9823 (N_9823,N_3356,N_1359);
and U9824 (N_9824,N_521,N_4334);
nor U9825 (N_9825,N_1422,N_1324);
nor U9826 (N_9826,N_4094,N_1608);
nand U9827 (N_9827,N_1336,N_937);
nand U9828 (N_9828,N_4821,N_264);
or U9829 (N_9829,N_428,N_317);
or U9830 (N_9830,N_437,N_4195);
xnor U9831 (N_9831,N_3289,N_3352);
nand U9832 (N_9832,N_3135,N_3368);
and U9833 (N_9833,N_3845,N_3029);
or U9834 (N_9834,N_668,N_2558);
nand U9835 (N_9835,N_2218,N_1561);
nand U9836 (N_9836,N_609,N_2025);
and U9837 (N_9837,N_1172,N_4782);
xnor U9838 (N_9838,N_493,N_1656);
and U9839 (N_9839,N_2940,N_752);
nand U9840 (N_9840,N_1365,N_3913);
and U9841 (N_9841,N_950,N_4848);
nor U9842 (N_9842,N_4332,N_2459);
nand U9843 (N_9843,N_4568,N_4955);
nand U9844 (N_9844,N_2140,N_1097);
or U9845 (N_9845,N_2092,N_1576);
nand U9846 (N_9846,N_179,N_337);
nand U9847 (N_9847,N_774,N_4343);
nor U9848 (N_9848,N_692,N_291);
and U9849 (N_9849,N_157,N_2786);
nand U9850 (N_9850,N_2399,N_2917);
nor U9851 (N_9851,N_582,N_3795);
and U9852 (N_9852,N_949,N_883);
or U9853 (N_9853,N_246,N_3771);
nand U9854 (N_9854,N_3646,N_2109);
nor U9855 (N_9855,N_823,N_2454);
nand U9856 (N_9856,N_4968,N_4910);
nand U9857 (N_9857,N_1412,N_3134);
nor U9858 (N_9858,N_1275,N_3886);
nand U9859 (N_9859,N_3038,N_3377);
and U9860 (N_9860,N_3261,N_206);
nor U9861 (N_9861,N_3780,N_2645);
or U9862 (N_9862,N_2237,N_2344);
and U9863 (N_9863,N_1577,N_1963);
or U9864 (N_9864,N_3698,N_101);
nand U9865 (N_9865,N_2553,N_806);
nor U9866 (N_9866,N_4611,N_556);
nand U9867 (N_9867,N_3104,N_3380);
nand U9868 (N_9868,N_2433,N_1964);
nor U9869 (N_9869,N_4921,N_739);
nor U9870 (N_9870,N_2443,N_2944);
nor U9871 (N_9871,N_1361,N_2636);
nor U9872 (N_9872,N_2138,N_2467);
and U9873 (N_9873,N_3814,N_4452);
and U9874 (N_9874,N_58,N_2992);
nand U9875 (N_9875,N_3821,N_91);
nand U9876 (N_9876,N_1476,N_453);
nand U9877 (N_9877,N_173,N_2148);
nand U9878 (N_9878,N_3567,N_2424);
or U9879 (N_9879,N_667,N_1838);
and U9880 (N_9880,N_4078,N_2151);
and U9881 (N_9881,N_795,N_3486);
nor U9882 (N_9882,N_3708,N_1019);
and U9883 (N_9883,N_335,N_482);
and U9884 (N_9884,N_768,N_2641);
or U9885 (N_9885,N_3151,N_2420);
or U9886 (N_9886,N_3501,N_1653);
and U9887 (N_9887,N_361,N_254);
and U9888 (N_9888,N_4036,N_4575);
nand U9889 (N_9889,N_1737,N_746);
nor U9890 (N_9890,N_620,N_3465);
and U9891 (N_9891,N_690,N_3150);
nand U9892 (N_9892,N_1592,N_1576);
or U9893 (N_9893,N_3111,N_4051);
or U9894 (N_9894,N_1262,N_1833);
nand U9895 (N_9895,N_730,N_2385);
nor U9896 (N_9896,N_833,N_3293);
nor U9897 (N_9897,N_4512,N_1746);
nand U9898 (N_9898,N_2867,N_125);
or U9899 (N_9899,N_2816,N_1605);
and U9900 (N_9900,N_4829,N_4608);
nand U9901 (N_9901,N_464,N_2326);
or U9902 (N_9902,N_1541,N_3606);
nand U9903 (N_9903,N_3719,N_3941);
or U9904 (N_9904,N_1291,N_748);
or U9905 (N_9905,N_3405,N_2111);
and U9906 (N_9906,N_2673,N_830);
or U9907 (N_9907,N_1731,N_858);
and U9908 (N_9908,N_4221,N_2561);
and U9909 (N_9909,N_303,N_331);
or U9910 (N_9910,N_2652,N_3351);
nand U9911 (N_9911,N_637,N_2117);
or U9912 (N_9912,N_855,N_2317);
and U9913 (N_9913,N_3087,N_498);
or U9914 (N_9914,N_918,N_4224);
or U9915 (N_9915,N_1957,N_3418);
nor U9916 (N_9916,N_2191,N_4452);
nand U9917 (N_9917,N_4317,N_2724);
or U9918 (N_9918,N_4540,N_1157);
and U9919 (N_9919,N_4472,N_355);
or U9920 (N_9920,N_2818,N_2897);
nor U9921 (N_9921,N_420,N_4510);
nor U9922 (N_9922,N_1310,N_3312);
and U9923 (N_9923,N_3671,N_2668);
and U9924 (N_9924,N_2122,N_4973);
nand U9925 (N_9925,N_2890,N_894);
or U9926 (N_9926,N_36,N_4664);
nand U9927 (N_9927,N_78,N_181);
nand U9928 (N_9928,N_1536,N_801);
nand U9929 (N_9929,N_1216,N_2893);
or U9930 (N_9930,N_4344,N_4761);
nor U9931 (N_9931,N_2128,N_2428);
nand U9932 (N_9932,N_4305,N_4850);
nor U9933 (N_9933,N_4128,N_2418);
and U9934 (N_9934,N_658,N_1720);
nand U9935 (N_9935,N_3693,N_4443);
xnor U9936 (N_9936,N_1006,N_1324);
nor U9937 (N_9937,N_3475,N_4245);
and U9938 (N_9938,N_2284,N_762);
or U9939 (N_9939,N_1955,N_4029);
and U9940 (N_9940,N_3423,N_4554);
nor U9941 (N_9941,N_206,N_3226);
nor U9942 (N_9942,N_3462,N_2452);
xnor U9943 (N_9943,N_779,N_3598);
or U9944 (N_9944,N_2693,N_3383);
nand U9945 (N_9945,N_2877,N_2401);
nand U9946 (N_9946,N_2497,N_805);
and U9947 (N_9947,N_2238,N_3105);
nor U9948 (N_9948,N_2833,N_1506);
nor U9949 (N_9949,N_3639,N_605);
and U9950 (N_9950,N_4345,N_2141);
and U9951 (N_9951,N_895,N_2765);
nand U9952 (N_9952,N_2515,N_2806);
or U9953 (N_9953,N_1473,N_2856);
and U9954 (N_9954,N_2598,N_2926);
or U9955 (N_9955,N_4195,N_3985);
nor U9956 (N_9956,N_2563,N_72);
and U9957 (N_9957,N_3902,N_976);
nand U9958 (N_9958,N_1142,N_87);
nor U9959 (N_9959,N_519,N_2782);
nor U9960 (N_9960,N_797,N_4013);
nand U9961 (N_9961,N_2176,N_1158);
and U9962 (N_9962,N_4942,N_565);
and U9963 (N_9963,N_300,N_847);
xnor U9964 (N_9964,N_2437,N_965);
and U9965 (N_9965,N_66,N_1379);
or U9966 (N_9966,N_1465,N_662);
nand U9967 (N_9967,N_3074,N_3536);
or U9968 (N_9968,N_1811,N_2515);
and U9969 (N_9969,N_1630,N_1196);
nand U9970 (N_9970,N_1762,N_4464);
nor U9971 (N_9971,N_4129,N_1270);
or U9972 (N_9972,N_2927,N_32);
nor U9973 (N_9973,N_1372,N_1091);
and U9974 (N_9974,N_2815,N_4231);
or U9975 (N_9975,N_1493,N_3412);
nor U9976 (N_9976,N_588,N_2530);
nor U9977 (N_9977,N_3388,N_4103);
nor U9978 (N_9978,N_1706,N_2296);
nor U9979 (N_9979,N_1174,N_3392);
or U9980 (N_9980,N_1767,N_1705);
or U9981 (N_9981,N_3656,N_500);
or U9982 (N_9982,N_2657,N_711);
nand U9983 (N_9983,N_2822,N_274);
and U9984 (N_9984,N_2324,N_3515);
nor U9985 (N_9985,N_264,N_3011);
and U9986 (N_9986,N_181,N_4982);
or U9987 (N_9987,N_3815,N_4909);
nand U9988 (N_9988,N_1613,N_1090);
nor U9989 (N_9989,N_304,N_3029);
nand U9990 (N_9990,N_869,N_3921);
and U9991 (N_9991,N_2523,N_700);
and U9992 (N_9992,N_4740,N_2306);
or U9993 (N_9993,N_890,N_1787);
nor U9994 (N_9994,N_3919,N_457);
and U9995 (N_9995,N_1288,N_4187);
nor U9996 (N_9996,N_4322,N_3354);
and U9997 (N_9997,N_371,N_2833);
nand U9998 (N_9998,N_123,N_3631);
nand U9999 (N_9999,N_4503,N_2700);
xnor UO_0 (O_0,N_9348,N_9504);
and UO_1 (O_1,N_5569,N_5725);
and UO_2 (O_2,N_5147,N_9342);
nand UO_3 (O_3,N_6909,N_9589);
and UO_4 (O_4,N_8705,N_5606);
nand UO_5 (O_5,N_5362,N_7755);
nor UO_6 (O_6,N_9784,N_5125);
nand UO_7 (O_7,N_9228,N_8766);
nor UO_8 (O_8,N_7050,N_5932);
or UO_9 (O_9,N_6113,N_8983);
and UO_10 (O_10,N_8260,N_5881);
or UO_11 (O_11,N_8726,N_9237);
nor UO_12 (O_12,N_7799,N_9275);
nand UO_13 (O_13,N_5453,N_7626);
or UO_14 (O_14,N_7087,N_7363);
nand UO_15 (O_15,N_8273,N_7793);
or UO_16 (O_16,N_8321,N_5554);
nand UO_17 (O_17,N_8415,N_7445);
and UO_18 (O_18,N_7441,N_9861);
nand UO_19 (O_19,N_7433,N_7866);
nor UO_20 (O_20,N_6535,N_5162);
and UO_21 (O_21,N_9439,N_5355);
or UO_22 (O_22,N_5027,N_5485);
xor UO_23 (O_23,N_8000,N_5251);
nor UO_24 (O_24,N_7423,N_6196);
and UO_25 (O_25,N_9656,N_5252);
nor UO_26 (O_26,N_6236,N_8394);
nor UO_27 (O_27,N_8457,N_7268);
nor UO_28 (O_28,N_6479,N_9826);
or UO_29 (O_29,N_5006,N_6060);
or UO_30 (O_30,N_7974,N_8424);
nor UO_31 (O_31,N_6262,N_5416);
or UO_32 (O_32,N_8261,N_9605);
and UO_33 (O_33,N_9080,N_6041);
or UO_34 (O_34,N_5180,N_7979);
and UO_35 (O_35,N_5330,N_9007);
xor UO_36 (O_36,N_6175,N_6872);
and UO_37 (O_37,N_9979,N_7951);
nor UO_38 (O_38,N_7372,N_9953);
or UO_39 (O_39,N_5102,N_5175);
nand UO_40 (O_40,N_5492,N_8640);
and UO_41 (O_41,N_7182,N_5702);
nor UO_42 (O_42,N_6255,N_9761);
nand UO_43 (O_43,N_7325,N_8133);
or UO_44 (O_44,N_7887,N_9379);
and UO_45 (O_45,N_8443,N_9010);
nor UO_46 (O_46,N_7537,N_5433);
and UO_47 (O_47,N_8243,N_5685);
nor UO_48 (O_48,N_9577,N_5438);
and UO_49 (O_49,N_5998,N_8530);
nor UO_50 (O_50,N_9217,N_8523);
nand UO_51 (O_51,N_8698,N_5525);
nand UO_52 (O_52,N_7839,N_9367);
nand UO_53 (O_53,N_9611,N_8925);
nand UO_54 (O_54,N_9135,N_7101);
or UO_55 (O_55,N_7547,N_8662);
or UO_56 (O_56,N_6588,N_9083);
nand UO_57 (O_57,N_8054,N_7094);
or UO_58 (O_58,N_9622,N_5807);
and UO_59 (O_59,N_6350,N_6115);
and UO_60 (O_60,N_6348,N_7119);
nand UO_61 (O_61,N_6659,N_8023);
or UO_62 (O_62,N_8211,N_8886);
or UO_63 (O_63,N_8475,N_6982);
nand UO_64 (O_64,N_5971,N_9763);
xor UO_65 (O_65,N_8219,N_9381);
nor UO_66 (O_66,N_7569,N_7779);
nand UO_67 (O_67,N_8645,N_5883);
nand UO_68 (O_68,N_6309,N_9690);
nor UO_69 (O_69,N_8758,N_7987);
and UO_70 (O_70,N_6932,N_8990);
and UO_71 (O_71,N_9998,N_7338);
nor UO_72 (O_72,N_5649,N_5014);
nor UO_73 (O_73,N_7628,N_9549);
or UO_74 (O_74,N_6709,N_9680);
or UO_75 (O_75,N_7237,N_5724);
nor UO_76 (O_76,N_6239,N_5732);
and UO_77 (O_77,N_8388,N_6552);
nor UO_78 (O_78,N_8794,N_7390);
nand UO_79 (O_79,N_9819,N_8269);
nor UO_80 (O_80,N_8467,N_5923);
and UO_81 (O_81,N_8996,N_8188);
nand UO_82 (O_82,N_7361,N_5350);
or UO_83 (O_83,N_6856,N_6871);
or UO_84 (O_84,N_5432,N_8783);
nor UO_85 (O_85,N_9264,N_9664);
nand UO_86 (O_86,N_8717,N_6140);
and UO_87 (O_87,N_8862,N_9357);
and UO_88 (O_88,N_6295,N_8655);
nor UO_89 (O_89,N_5636,N_7303);
or UO_90 (O_90,N_8927,N_7985);
and UO_91 (O_91,N_7369,N_6577);
nand UO_92 (O_92,N_6241,N_6067);
nand UO_93 (O_93,N_8477,N_9049);
nor UO_94 (O_94,N_8421,N_9505);
nand UO_95 (O_95,N_6480,N_8642);
nand UO_96 (O_96,N_7851,N_9644);
nor UO_97 (O_97,N_8406,N_5559);
or UO_98 (O_98,N_8396,N_6341);
and UO_99 (O_99,N_6963,N_9058);
nand UO_100 (O_100,N_6036,N_5710);
nor UO_101 (O_101,N_6234,N_5363);
and UO_102 (O_102,N_5387,N_7199);
and UO_103 (O_103,N_8881,N_5188);
xor UO_104 (O_104,N_9402,N_9646);
nand UO_105 (O_105,N_7929,N_7930);
nor UO_106 (O_106,N_7550,N_7563);
xor UO_107 (O_107,N_6408,N_8974);
and UO_108 (O_108,N_8491,N_9751);
nand UO_109 (O_109,N_9582,N_9478);
nand UO_110 (O_110,N_5228,N_7259);
nor UO_111 (O_111,N_9369,N_5012);
and UO_112 (O_112,N_8091,N_8561);
and UO_113 (O_113,N_6714,N_6939);
nor UO_114 (O_114,N_9684,N_8264);
or UO_115 (O_115,N_7815,N_6985);
nor UO_116 (O_116,N_8108,N_5662);
and UO_117 (O_117,N_5300,N_5641);
nand UO_118 (O_118,N_8663,N_5750);
or UO_119 (O_119,N_6509,N_6565);
nand UO_120 (O_120,N_8131,N_9982);
nand UO_121 (O_121,N_8817,N_5368);
xnor UO_122 (O_122,N_9392,N_7928);
and UO_123 (O_123,N_8044,N_9908);
or UO_124 (O_124,N_6821,N_5161);
and UO_125 (O_125,N_5622,N_7996);
nor UO_126 (O_126,N_9409,N_6655);
and UO_127 (O_127,N_8096,N_8901);
nor UO_128 (O_128,N_6110,N_8757);
or UO_129 (O_129,N_6216,N_6634);
nor UO_130 (O_130,N_9389,N_7680);
nor UO_131 (O_131,N_6089,N_6644);
nor UO_132 (O_132,N_6218,N_9043);
nand UO_133 (O_133,N_6781,N_6306);
or UO_134 (O_134,N_8776,N_8774);
or UO_135 (O_135,N_7570,N_7897);
and UO_136 (O_136,N_7465,N_8356);
nor UO_137 (O_137,N_9932,N_5365);
nor UO_138 (O_138,N_9566,N_6360);
nand UO_139 (O_139,N_8075,N_6725);
and UO_140 (O_140,N_9428,N_7572);
nand UO_141 (O_141,N_8514,N_9978);
and UO_142 (O_142,N_8621,N_6040);
nand UO_143 (O_143,N_7472,N_9195);
or UO_144 (O_144,N_9960,N_6153);
or UO_145 (O_145,N_7451,N_8404);
or UO_146 (O_146,N_8454,N_6305);
nand UO_147 (O_147,N_6590,N_5498);
nand UO_148 (O_148,N_9199,N_7261);
or UO_149 (O_149,N_8770,N_6142);
nor UO_150 (O_150,N_7109,N_6682);
or UO_151 (O_151,N_7927,N_5104);
or UO_152 (O_152,N_9648,N_9300);
nor UO_153 (O_153,N_9554,N_6958);
nor UO_154 (O_154,N_8287,N_5898);
and UO_155 (O_155,N_8105,N_5046);
nor UO_156 (O_156,N_7157,N_7923);
and UO_157 (O_157,N_8857,N_7129);
nor UO_158 (O_158,N_5233,N_9425);
and UO_159 (O_159,N_7986,N_5231);
and UO_160 (O_160,N_8874,N_8239);
nand UO_161 (O_161,N_5292,N_5903);
or UO_162 (O_162,N_6254,N_5527);
nor UO_163 (O_163,N_9820,N_8891);
nand UO_164 (O_164,N_8538,N_7807);
and UO_165 (O_165,N_7753,N_6486);
nand UO_166 (O_166,N_6721,N_6183);
and UO_167 (O_167,N_7694,N_5659);
nor UO_168 (O_168,N_7977,N_9339);
and UO_169 (O_169,N_6191,N_8110);
nor UO_170 (O_170,N_9364,N_7737);
and UO_171 (O_171,N_9437,N_5706);
or UO_172 (O_172,N_8877,N_8749);
nand UO_173 (O_173,N_9781,N_5415);
and UO_174 (O_174,N_5229,N_7952);
nand UO_175 (O_175,N_9806,N_6708);
nor UO_176 (O_176,N_9889,N_7385);
nor UO_177 (O_177,N_7745,N_8437);
nand UO_178 (O_178,N_8816,N_6297);
and UO_179 (O_179,N_6162,N_9140);
or UO_180 (O_180,N_7443,N_5771);
or UO_181 (O_181,N_7350,N_9031);
and UO_182 (O_182,N_6111,N_5537);
nand UO_183 (O_183,N_8658,N_9709);
nor UO_184 (O_184,N_8262,N_5653);
and UO_185 (O_185,N_5604,N_8715);
nand UO_186 (O_186,N_5873,N_9916);
or UO_187 (O_187,N_5047,N_9345);
or UO_188 (O_188,N_8944,N_9874);
or UO_189 (O_189,N_9333,N_6308);
nand UO_190 (O_190,N_7701,N_9666);
nand UO_191 (O_191,N_6393,N_5817);
nand UO_192 (O_192,N_8842,N_5382);
nand UO_193 (O_193,N_8731,N_6505);
nor UO_194 (O_194,N_9662,N_8452);
and UO_195 (O_195,N_8408,N_6704);
nand UO_196 (O_196,N_7598,N_6584);
and UO_197 (O_197,N_9426,N_6056);
or UO_198 (O_198,N_5146,N_7686);
nor UO_199 (O_199,N_6718,N_7111);
nor UO_200 (O_200,N_8524,N_8125);
nor UO_201 (O_201,N_9056,N_9997);
and UO_202 (O_202,N_7647,N_6671);
nand UO_203 (O_203,N_7298,N_9789);
or UO_204 (O_204,N_8307,N_6698);
nor UO_205 (O_205,N_7112,N_5515);
nor UO_206 (O_206,N_9393,N_6520);
and UO_207 (O_207,N_8455,N_9420);
nor UO_208 (O_208,N_7775,N_8200);
and UO_209 (O_209,N_8461,N_9061);
and UO_210 (O_210,N_7912,N_9051);
or UO_211 (O_211,N_6347,N_9655);
or UO_212 (O_212,N_6016,N_9601);
nor UO_213 (O_213,N_5663,N_8166);
xnor UO_214 (O_214,N_9067,N_8340);
or UO_215 (O_215,N_8399,N_9363);
nand UO_216 (O_216,N_7241,N_6276);
and UO_217 (O_217,N_6334,N_9254);
nor UO_218 (O_218,N_9537,N_6460);
nor UO_219 (O_219,N_9187,N_8485);
nand UO_220 (O_220,N_6929,N_5205);
or UO_221 (O_221,N_8285,N_8546);
and UO_222 (O_222,N_9623,N_5192);
nor UO_223 (O_223,N_7789,N_8449);
nor UO_224 (O_224,N_7042,N_6105);
and UO_225 (O_225,N_7797,N_6123);
nand UO_226 (O_226,N_5405,N_8799);
nand UO_227 (O_227,N_8912,N_7613);
nand UO_228 (O_228,N_6788,N_9096);
and UO_229 (O_229,N_6516,N_9054);
and UO_230 (O_230,N_8782,N_8900);
nor UO_231 (O_231,N_6601,N_9474);
nand UO_232 (O_232,N_9436,N_9277);
or UO_233 (O_233,N_7430,N_5909);
or UO_234 (O_234,N_8550,N_6974);
nand UO_235 (O_235,N_9812,N_9695);
and UO_236 (O_236,N_5744,N_6035);
nand UO_237 (O_237,N_8797,N_9640);
nand UO_238 (O_238,N_7475,N_5572);
and UO_239 (O_239,N_8649,N_6228);
nand UO_240 (O_240,N_5912,N_9193);
and UO_241 (O_241,N_9990,N_6453);
and UO_242 (O_242,N_7032,N_6990);
nand UO_243 (O_243,N_7909,N_5581);
nor UO_244 (O_244,N_5099,N_8137);
nor UO_245 (O_245,N_9972,N_9456);
nor UO_246 (O_246,N_6436,N_9471);
or UO_247 (O_247,N_5941,N_5984);
and UO_248 (O_248,N_8892,N_7861);
and UO_249 (O_249,N_8198,N_9580);
nor UO_250 (O_250,N_6832,N_8947);
xnor UO_251 (O_251,N_5978,N_5956);
nor UO_252 (O_252,N_8923,N_8690);
nor UO_253 (O_253,N_7911,N_5183);
nor UO_254 (O_254,N_9071,N_6419);
nand UO_255 (O_255,N_8134,N_8378);
nand UO_256 (O_256,N_8975,N_9029);
nand UO_257 (O_257,N_7968,N_7651);
xnor UO_258 (O_258,N_5331,N_7809);
or UO_259 (O_259,N_7892,N_7343);
or UO_260 (O_260,N_6246,N_9163);
nor UO_261 (O_261,N_8496,N_5277);
or UO_262 (O_262,N_6597,N_9138);
and UO_263 (O_263,N_5810,N_6854);
and UO_264 (O_264,N_7932,N_5566);
or UO_265 (O_265,N_5716,N_8823);
and UO_266 (O_266,N_5308,N_6214);
nor UO_267 (O_267,N_9795,N_9444);
and UO_268 (O_268,N_6518,N_8596);
nand UO_269 (O_269,N_7106,N_9966);
nor UO_270 (O_270,N_6235,N_5507);
xor UO_271 (O_271,N_9980,N_8159);
nand UO_272 (O_272,N_7144,N_5356);
or UO_273 (O_273,N_7047,N_9739);
or UO_274 (O_274,N_9918,N_5217);
nand UO_275 (O_275,N_8368,N_8604);
nand UO_276 (O_276,N_9143,N_5895);
nand UO_277 (O_277,N_8344,N_9541);
and UO_278 (O_278,N_8624,N_5376);
nor UO_279 (O_279,N_5195,N_7484);
or UO_280 (O_280,N_5155,N_9778);
and UO_281 (O_281,N_7405,N_9109);
or UO_282 (O_282,N_5428,N_6225);
nand UO_283 (O_283,N_5271,N_6692);
or UO_284 (O_284,N_7420,N_9876);
and UO_285 (O_285,N_6034,N_6268);
or UO_286 (O_286,N_6193,N_6296);
and UO_287 (O_287,N_8070,N_9074);
or UO_288 (O_288,N_9146,N_6910);
and UO_289 (O_289,N_8410,N_7035);
and UO_290 (O_290,N_6748,N_9190);
and UO_291 (O_291,N_8322,N_9849);
nand UO_292 (O_292,N_9288,N_7057);
nor UO_293 (O_293,N_7041,N_6905);
nor UO_294 (O_294,N_6705,N_9770);
and UO_295 (O_295,N_8025,N_5670);
nor UO_296 (O_296,N_8458,N_8227);
and UO_297 (O_297,N_6512,N_7333);
and UO_298 (O_298,N_6195,N_9914);
and UO_299 (O_299,N_7356,N_5444);
and UO_300 (O_300,N_5799,N_8139);
or UO_301 (O_301,N_7891,N_7786);
and UO_302 (O_302,N_5066,N_7865);
or UO_303 (O_303,N_7473,N_8945);
nor UO_304 (O_304,N_6507,N_5965);
nor UO_305 (O_305,N_7534,N_8627);
and UO_306 (O_306,N_7907,N_5553);
nor UO_307 (O_307,N_7105,N_6904);
and UO_308 (O_308,N_7565,N_7337);
nor UO_309 (O_309,N_7586,N_8436);
nand UO_310 (O_310,N_7762,N_6976);
or UO_311 (O_311,N_9629,N_8522);
nand UO_312 (O_312,N_5281,N_7673);
and UO_313 (O_313,N_9533,N_9606);
nand UO_314 (O_314,N_9085,N_5770);
or UO_315 (O_315,N_6997,N_8807);
nor UO_316 (O_316,N_8329,N_5202);
and UO_317 (O_317,N_6546,N_8024);
nor UO_318 (O_318,N_5057,N_6116);
nor UO_319 (O_319,N_8063,N_9602);
or UO_320 (O_320,N_6828,N_9268);
or UO_321 (O_321,N_9098,N_9529);
and UO_322 (O_322,N_7376,N_5763);
nor UO_323 (O_323,N_6618,N_5509);
and UO_324 (O_324,N_6550,N_6430);
and UO_325 (O_325,N_7611,N_8818);
nand UO_326 (O_326,N_6328,N_6765);
nand UO_327 (O_327,N_9638,N_7699);
nor UO_328 (O_328,N_7198,N_9700);
or UO_329 (O_329,N_5836,N_7277);
nor UO_330 (O_330,N_9122,N_8691);
and UO_331 (O_331,N_6525,N_9612);
or UO_332 (O_332,N_7281,N_9015);
nand UO_333 (O_333,N_9331,N_6540);
and UO_334 (O_334,N_5409,N_5124);
nor UO_335 (O_335,N_5741,N_5263);
nand UO_336 (O_336,N_9343,N_5422);
or UO_337 (O_337,N_7285,N_6126);
nand UO_338 (O_338,N_9139,N_6531);
nand UO_339 (O_339,N_9780,N_7773);
and UO_340 (O_340,N_8360,N_9679);
and UO_341 (O_341,N_6059,N_7317);
and UO_342 (O_342,N_7629,N_5975);
nor UO_343 (O_343,N_5953,N_5671);
or UO_344 (O_344,N_7442,N_8934);
or UO_345 (O_345,N_9000,N_9689);
nand UO_346 (O_346,N_9141,N_8335);
nor UO_347 (O_347,N_5158,N_6727);
and UO_348 (O_348,N_9649,N_7631);
nor UO_349 (O_349,N_7328,N_6485);
and UO_350 (O_350,N_9065,N_9404);
or UO_351 (O_351,N_7409,N_7696);
and UO_352 (O_352,N_5044,N_5561);
and UO_353 (O_353,N_7486,N_5966);
or UO_354 (O_354,N_6771,N_9840);
nor UO_355 (O_355,N_8894,N_8088);
nor UO_356 (O_356,N_5605,N_6421);
nor UO_357 (O_357,N_7406,N_5901);
and UO_358 (O_358,N_5420,N_5088);
and UO_359 (O_359,N_7121,N_7532);
and UO_360 (O_360,N_9654,N_9527);
or UO_361 (O_361,N_9853,N_8354);
nor UO_362 (O_362,N_8614,N_9970);
and UO_363 (O_363,N_7636,N_6962);
nor UO_364 (O_364,N_9711,N_5623);
nand UO_365 (O_365,N_7713,N_8155);
or UO_366 (O_366,N_5549,N_7045);
and UO_367 (O_367,N_9118,N_8895);
nand UO_368 (O_368,N_8634,N_8296);
and UO_369 (O_369,N_5688,N_9848);
or UO_370 (O_370,N_9465,N_9921);
nand UO_371 (O_371,N_7397,N_6957);
nand UO_372 (O_372,N_7082,N_5595);
nor UO_373 (O_373,N_7104,N_8824);
xnor UO_374 (O_374,N_7467,N_6118);
and UO_375 (O_375,N_7068,N_9562);
or UO_376 (O_376,N_9366,N_5040);
or UO_377 (O_377,N_6657,N_7917);
or UO_378 (O_378,N_8221,N_8056);
nor UO_379 (O_379,N_5845,N_8018);
nor UO_380 (O_380,N_5906,N_5403);
nor UO_381 (O_381,N_5291,N_7377);
nand UO_382 (O_382,N_8804,N_7429);
and UO_383 (O_383,N_7899,N_7200);
nor UO_384 (O_384,N_6762,N_6521);
and UO_385 (O_385,N_5787,N_5074);
nand UO_386 (O_386,N_8968,N_8099);
or UO_387 (O_387,N_8949,N_7375);
nand UO_388 (O_388,N_7610,N_5002);
or UO_389 (O_389,N_7846,N_7131);
and UO_390 (O_390,N_7638,N_9941);
nor UO_391 (O_391,N_6425,N_6674);
and UO_392 (O_392,N_5045,N_8199);
or UO_393 (O_393,N_6654,N_5813);
or UO_394 (O_394,N_6282,N_6185);
and UO_395 (O_395,N_9441,N_5338);
nand UO_396 (O_396,N_7955,N_8414);
nor UO_397 (O_397,N_5765,N_7750);
nor UO_398 (O_398,N_8114,N_9131);
xnor UO_399 (O_399,N_8544,N_6023);
nand UO_400 (O_400,N_9121,N_6493);
nor UO_401 (O_401,N_7292,N_9753);
nand UO_402 (O_402,N_9936,N_9240);
nor UO_403 (O_403,N_5950,N_7945);
nand UO_404 (O_404,N_6723,N_6209);
nor UO_405 (O_405,N_8847,N_9150);
nand UO_406 (O_406,N_8147,N_9893);
nand UO_407 (O_407,N_6700,N_5959);
nand UO_408 (O_408,N_7487,N_5607);
or UO_409 (O_409,N_5977,N_7644);
and UO_410 (O_410,N_5550,N_9421);
and UO_411 (O_411,N_5486,N_9183);
nor UO_412 (O_412,N_6605,N_8639);
or UO_413 (O_413,N_6959,N_6906);
and UO_414 (O_414,N_5690,N_5425);
and UO_415 (O_415,N_7953,N_6855);
nand UO_416 (O_416,N_7746,N_6712);
or UO_417 (O_417,N_9295,N_7384);
and UO_418 (O_418,N_7033,N_8019);
and UO_419 (O_419,N_9347,N_5306);
or UO_420 (O_420,N_8681,N_8967);
nor UO_421 (O_421,N_7837,N_8680);
and UO_422 (O_422,N_5853,N_7300);
nand UO_423 (O_423,N_6020,N_7049);
or UO_424 (O_424,N_8599,N_5735);
and UO_425 (O_425,N_6365,N_9106);
and UO_426 (O_426,N_7878,N_9179);
nand UO_427 (O_427,N_8079,N_6984);
nor UO_428 (O_428,N_6028,N_9833);
and UO_429 (O_429,N_8306,N_5426);
or UO_430 (O_430,N_6510,N_5602);
and UO_431 (O_431,N_5065,N_7780);
or UO_432 (O_432,N_5556,N_7253);
nor UO_433 (O_433,N_7118,N_5145);
and UO_434 (O_434,N_9274,N_8622);
and UO_435 (O_435,N_6536,N_6873);
nand UO_436 (O_436,N_7204,N_9231);
nand UO_437 (O_437,N_8637,N_9319);
xor UO_438 (O_438,N_6281,N_7095);
nand UO_439 (O_439,N_5004,N_5258);
and UO_440 (O_440,N_5406,N_9287);
nor UO_441 (O_441,N_5760,N_6138);
nor UO_442 (O_442,N_6455,N_9742);
or UO_443 (O_443,N_6292,N_5773);
xnor UO_444 (O_444,N_5034,N_8153);
and UO_445 (O_445,N_9842,N_7772);
nand UO_446 (O_446,N_7460,N_6833);
nand UO_447 (O_447,N_5962,N_8126);
nor UO_448 (O_448,N_8535,N_6936);
nand UO_449 (O_449,N_6567,N_5051);
nor UO_450 (O_450,N_8802,N_6622);
nand UO_451 (O_451,N_7166,N_8697);
nand UO_452 (O_452,N_9329,N_9276);
nand UO_453 (O_453,N_7291,N_7414);
and UO_454 (O_454,N_9344,N_5746);
nand UO_455 (O_455,N_9519,N_5140);
nor UO_456 (O_456,N_9930,N_7102);
nor UO_457 (O_457,N_6861,N_7785);
or UO_458 (O_458,N_9090,N_7051);
or UO_459 (O_459,N_7189,N_8355);
nand UO_460 (O_460,N_6652,N_5424);
nand UO_461 (O_461,N_6490,N_7079);
or UO_462 (O_462,N_8814,N_8030);
and UO_463 (O_463,N_9208,N_8248);
xor UO_464 (O_464,N_6633,N_9062);
nand UO_465 (O_465,N_8250,N_6903);
nand UO_466 (O_466,N_6613,N_6809);
and UO_467 (O_467,N_9318,N_7224);
or UO_468 (O_468,N_9283,N_9928);
and UO_469 (O_469,N_9373,N_6843);
and UO_470 (O_470,N_9816,N_6775);
nand UO_471 (O_471,N_7058,N_5316);
nand UO_472 (O_472,N_6750,N_6780);
and UO_473 (O_473,N_8745,N_7402);
nor UO_474 (O_474,N_9660,N_6286);
or UO_475 (O_475,N_8065,N_8254);
or UO_476 (O_476,N_9484,N_9515);
nor UO_477 (O_477,N_7860,N_7011);
or UO_478 (O_478,N_7408,N_8113);
nor UO_479 (O_479,N_5132,N_5397);
nand UO_480 (O_480,N_5629,N_7802);
or UO_481 (O_481,N_9467,N_6304);
nand UO_482 (O_482,N_5348,N_5838);
or UO_483 (O_483,N_9744,N_7017);
nor UO_484 (O_484,N_6848,N_7916);
and UO_485 (O_485,N_8298,N_6989);
nand UO_486 (O_486,N_7055,N_5187);
and UO_487 (O_487,N_6791,N_9434);
and UO_488 (O_488,N_6575,N_9093);
nor UO_489 (O_489,N_7918,N_8411);
nand UO_490 (O_490,N_9394,N_6398);
nand UO_491 (O_491,N_9950,N_5824);
nand UO_492 (O_492,N_6739,N_5323);
xor UO_493 (O_493,N_6824,N_6145);
and UO_494 (O_494,N_7961,N_7885);
or UO_495 (O_495,N_5856,N_8428);
or UO_496 (O_496,N_8972,N_7245);
nand UO_497 (O_497,N_8553,N_7876);
or UO_498 (O_498,N_8089,N_6549);
and UO_499 (O_499,N_6889,N_9705);
and UO_500 (O_500,N_7819,N_8186);
or UO_501 (O_501,N_8425,N_8819);
nor UO_502 (O_502,N_5290,N_9002);
xnor UO_503 (O_503,N_5593,N_9783);
and UO_504 (O_504,N_6229,N_7814);
nor UO_505 (O_505,N_5674,N_8775);
nor UO_506 (O_506,N_7393,N_9004);
and UO_507 (O_507,N_7437,N_5893);
nand UO_508 (O_508,N_7542,N_5769);
and UO_509 (O_509,N_9748,N_5875);
and UO_510 (O_510,N_5165,N_7275);
nor UO_511 (O_511,N_9081,N_5859);
nand UO_512 (O_512,N_9963,N_9581);
nor UO_513 (O_513,N_8274,N_8119);
and UO_514 (O_514,N_6072,N_5224);
nand UO_515 (O_515,N_6397,N_9142);
nor UO_516 (O_516,N_7299,N_9845);
or UO_517 (O_517,N_5410,N_9961);
nand UO_518 (O_518,N_5399,N_8441);
and UO_519 (O_519,N_7206,N_8395);
or UO_520 (O_520,N_6586,N_6002);
and UO_521 (O_521,N_6642,N_7736);
nand UO_522 (O_522,N_9880,N_6483);
and UO_523 (O_523,N_8836,N_7886);
or UO_524 (O_524,N_6921,N_7803);
nor UO_525 (O_525,N_7761,N_5111);
or UO_526 (O_526,N_9308,N_9947);
nand UO_527 (O_527,N_6137,N_6606);
nand UO_528 (O_528,N_6491,N_9390);
or UO_529 (O_529,N_6404,N_6171);
and UO_530 (O_530,N_6336,N_5249);
or UO_531 (O_531,N_8174,N_6263);
and UO_532 (O_532,N_6198,N_5620);
nor UO_533 (O_533,N_7392,N_6379);
nand UO_534 (O_534,N_8313,N_8450);
nor UO_535 (O_535,N_7379,N_7302);
nand UO_536 (O_536,N_9865,N_9694);
and UO_537 (O_537,N_7497,N_5178);
nor UO_538 (O_538,N_8080,N_5342);
or UO_539 (O_539,N_8795,N_5131);
or UO_540 (O_540,N_5783,N_5852);
and UO_541 (O_541,N_6969,N_7688);
nand UO_542 (O_542,N_9503,N_6619);
nor UO_543 (O_543,N_5005,N_9238);
and UO_544 (O_544,N_6947,N_7967);
and UO_545 (O_545,N_8659,N_6592);
nand UO_546 (O_546,N_5298,N_7934);
nand UO_547 (O_547,N_7820,N_8201);
and UO_548 (O_548,N_7114,N_6326);
or UO_549 (O_549,N_6805,N_6163);
and UO_550 (O_550,N_8439,N_6437);
nand UO_551 (O_551,N_5384,N_6043);
nand UO_552 (O_552,N_8281,N_8429);
and UO_553 (O_553,N_6445,N_9782);
nand UO_554 (O_554,N_9204,N_6203);
or UO_555 (O_555,N_5644,N_6556);
and UO_556 (O_556,N_6972,N_9745);
and UO_557 (O_557,N_5301,N_5068);
nor UO_558 (O_558,N_5798,N_5170);
and UO_559 (O_559,N_5021,N_5043);
or UO_560 (O_560,N_5321,N_5101);
and UO_561 (O_561,N_5761,N_5567);
or UO_562 (O_562,N_5599,N_6381);
nand UO_563 (O_563,N_8168,N_8087);
and UO_564 (O_564,N_8017,N_7599);
or UO_565 (O_565,N_8385,N_7439);
or UO_566 (O_566,N_6274,N_9946);
nand UO_567 (O_567,N_7187,N_8316);
nand UO_568 (O_568,N_7717,N_8098);
nor UO_569 (O_569,N_6627,N_9985);
nor UO_570 (O_570,N_7346,N_6847);
and UO_571 (O_571,N_7715,N_9650);
and UO_572 (O_572,N_9169,N_6853);
nand UO_573 (O_573,N_6650,N_9633);
nand UO_574 (O_574,N_5815,N_6389);
nand UO_575 (O_575,N_9906,N_6761);
and UO_576 (O_576,N_7107,N_5095);
nand UO_577 (O_577,N_9245,N_5130);
and UO_578 (O_578,N_6769,N_9440);
and UO_579 (O_579,N_6978,N_5834);
xnor UO_580 (O_580,N_6732,N_5577);
nand UO_581 (O_581,N_9321,N_5392);
or UO_582 (O_582,N_9616,N_7209);
nand UO_583 (O_583,N_6164,N_9257);
nand UO_584 (O_584,N_6073,N_6005);
xor UO_585 (O_585,N_5615,N_5097);
or UO_586 (O_586,N_5896,N_9591);
nand UO_587 (O_587,N_8353,N_5031);
or UO_588 (O_588,N_9473,N_6322);
nand UO_589 (O_589,N_6728,N_6071);
nand UO_590 (O_590,N_7760,N_7883);
nand UO_591 (O_591,N_9117,N_8432);
nand UO_592 (O_592,N_7194,N_8754);
nand UO_593 (O_593,N_8128,N_6212);
nand UO_594 (O_594,N_8148,N_7524);
or UO_595 (O_595,N_7791,N_9887);
or UO_596 (O_596,N_7998,N_5528);
nand UO_597 (O_597,N_8061,N_5168);
or UO_598 (O_598,N_6131,N_9647);
and UO_599 (O_599,N_8861,N_9911);
nor UO_600 (O_600,N_9362,N_8100);
or UO_601 (O_601,N_9125,N_8889);
xor UO_602 (O_602,N_5497,N_7152);
nand UO_603 (O_603,N_9064,N_7658);
xnor UO_604 (O_604,N_9101,N_5513);
nand UO_605 (O_605,N_8601,N_6374);
nor UO_606 (O_606,N_9670,N_9877);
and UO_607 (O_607,N_7440,N_5742);
nand UO_608 (O_608,N_6764,N_7858);
and UO_609 (O_609,N_9637,N_5968);
nand UO_610 (O_610,N_6779,N_5656);
nor UO_611 (O_611,N_8879,N_9087);
and UO_612 (O_612,N_8667,N_7481);
nor UO_613 (O_613,N_5112,N_9220);
nand UO_614 (O_614,N_8654,N_5284);
or UO_615 (O_615,N_7595,N_7169);
nand UO_616 (O_616,N_5501,N_8579);
and UO_617 (O_617,N_7562,N_5758);
or UO_618 (O_618,N_6122,N_6944);
nor UO_619 (O_619,N_9634,N_8348);
nor UO_620 (O_620,N_9693,N_5455);
or UO_621 (O_621,N_5558,N_7632);
and UO_622 (O_622,N_6314,N_5126);
nor UO_623 (O_623,N_9814,N_5618);
nand UO_624 (O_624,N_6443,N_7027);
or UO_625 (O_625,N_5207,N_5536);
nand UO_626 (O_626,N_6572,N_6207);
or UO_627 (O_627,N_7190,N_5328);
nor UO_628 (O_628,N_8122,N_7428);
or UO_629 (O_629,N_7924,N_6628);
or UO_630 (O_630,N_6407,N_9181);
and UO_631 (O_631,N_5086,N_9450);
or UO_632 (O_632,N_5121,N_6785);
and UO_633 (O_633,N_8916,N_7536);
nor UO_634 (O_634,N_8665,N_9267);
nor UO_635 (O_635,N_7663,N_5520);
nor UO_636 (O_636,N_7850,N_9852);
nor UO_637 (O_637,N_7578,N_8319);
and UO_638 (O_638,N_9620,N_5668);
xnor UO_639 (O_639,N_6689,N_9777);
nand UO_640 (O_640,N_5056,N_5847);
and UO_641 (O_641,N_8431,N_8366);
and UO_642 (O_642,N_8256,N_6695);
nand UO_643 (O_643,N_6738,N_6677);
and UO_644 (O_644,N_6130,N_9531);
nand UO_645 (O_645,N_7594,N_9712);
or UO_646 (O_646,N_8342,N_7625);
nor UO_647 (O_647,N_7216,N_7588);
or UO_648 (O_648,N_8586,N_5870);
nand UO_649 (O_649,N_5797,N_8118);
nor UO_650 (O_650,N_6083,N_6880);
nand UO_651 (O_651,N_5683,N_9353);
nand UO_652 (O_652,N_8695,N_8844);
nand UO_653 (O_653,N_7516,N_7310);
and UO_654 (O_654,N_5596,N_7271);
or UO_655 (O_655,N_7545,N_6656);
nand UO_656 (O_656,N_6369,N_6461);
and UO_657 (O_657,N_9836,N_6037);
or UO_658 (O_658,N_7052,N_7227);
nor UO_659 (O_659,N_8611,N_8855);
and UO_660 (O_660,N_9256,N_7345);
or UO_661 (O_661,N_8572,N_8865);
and UO_662 (O_662,N_9136,N_6931);
or UO_663 (O_663,N_9273,N_9147);
or UO_664 (O_664,N_5866,N_8067);
and UO_665 (O_665,N_5085,N_9939);
or UO_666 (O_666,N_8291,N_7528);
or UO_667 (O_667,N_5477,N_7777);
nand UO_668 (O_668,N_6635,N_5571);
or UO_669 (O_669,N_6548,N_6951);
nor UO_670 (O_670,N_9675,N_8176);
and UO_671 (O_671,N_9448,N_6842);
nor UO_672 (O_672,N_7692,N_6054);
nor UO_673 (O_673,N_8101,N_5575);
nor UO_674 (O_674,N_9824,N_6703);
nor UO_675 (O_675,N_5214,N_5437);
and UO_676 (O_676,N_8129,N_7220);
nand UO_677 (O_677,N_7168,N_5345);
or UO_678 (O_678,N_5944,N_8510);
nand UO_679 (O_679,N_9202,N_8971);
nor UO_680 (O_680,N_5830,N_6364);
nor UO_681 (O_681,N_5584,N_7763);
or UO_682 (O_682,N_8345,N_6716);
nor UO_683 (O_683,N_8577,N_9999);
nor UO_684 (O_684,N_7005,N_8419);
and UO_685 (O_685,N_7523,N_5723);
nor UO_686 (O_686,N_5992,N_8641);
or UO_687 (O_687,N_5256,N_7267);
and UO_688 (O_688,N_6787,N_8120);
nand UO_689 (O_689,N_6745,N_5667);
nor UO_690 (O_690,N_5227,N_8708);
nor UO_691 (O_691,N_7018,N_9910);
or UO_692 (O_692,N_8066,N_6080);
and UO_693 (O_693,N_7342,N_5583);
nor UO_694 (O_694,N_5935,N_8271);
nor UO_695 (O_695,N_9509,N_8526);
nand UO_696 (O_696,N_7425,N_6498);
nor UO_697 (O_697,N_6807,N_8935);
nor UO_698 (O_698,N_9413,N_8214);
and UO_699 (O_699,N_8037,N_6457);
and UO_700 (O_700,N_9092,N_9243);
and UO_701 (O_701,N_6269,N_9418);
or UO_702 (O_702,N_7926,N_5888);
nand UO_703 (O_703,N_7856,N_7509);
and UO_704 (O_704,N_8253,N_7714);
and UO_705 (O_705,N_9258,N_9959);
nand UO_706 (O_706,N_6047,N_5352);
and UO_707 (O_707,N_9030,N_7874);
nor UO_708 (O_708,N_6722,N_9933);
and UO_709 (O_709,N_8893,N_7995);
and UO_710 (O_710,N_8676,N_9059);
nor UO_711 (O_711,N_5461,N_6260);
nand UO_712 (O_712,N_5351,N_9455);
nand UO_713 (O_713,N_6557,N_7901);
and UO_714 (O_714,N_9535,N_5934);
nor UO_715 (O_715,N_5691,N_6497);
and UO_716 (O_716,N_6270,N_5812);
nor UO_717 (O_717,N_7314,N_9438);
nand UO_718 (O_718,N_7432,N_5924);
nand UO_719 (O_719,N_6038,N_6706);
nand UO_720 (O_720,N_7490,N_5827);
and UO_721 (O_721,N_9557,N_8835);
and UO_722 (O_722,N_8623,N_6760);
or UO_723 (O_723,N_7783,N_8398);
nand UO_724 (O_724,N_8312,N_7412);
or UO_725 (O_725,N_7491,N_8302);
nor UO_726 (O_726,N_9708,N_6166);
nor UO_727 (O_727,N_7023,N_9057);
nand UO_728 (O_728,N_9236,N_7939);
nor UO_729 (O_729,N_9398,N_9801);
and UO_730 (O_730,N_9129,N_5948);
or UO_731 (O_731,N_9798,N_5851);
nor UO_732 (O_732,N_6554,N_8275);
or UO_733 (O_733,N_6839,N_6104);
nand UO_734 (O_734,N_9881,N_8143);
or UO_735 (O_735,N_7958,N_7202);
nand UO_736 (O_736,N_5800,N_5483);
or UO_737 (O_737,N_6204,N_5269);
nor UO_738 (O_738,N_9315,N_5951);
nand UO_739 (O_739,N_6481,N_5110);
nand UO_740 (O_740,N_9304,N_6376);
or UO_741 (O_741,N_5734,N_5117);
and UO_742 (O_742,N_9788,N_7341);
nand UO_743 (O_743,N_9613,N_5164);
and UO_744 (O_744,N_6687,N_5036);
nand UO_745 (O_745,N_8592,N_6349);
nor UO_746 (O_746,N_8969,N_6802);
nand UO_747 (O_747,N_8035,N_8259);
xnor UO_748 (O_748,N_5311,N_6753);
and UO_749 (O_749,N_8460,N_7690);
and UO_750 (O_750,N_7794,N_5222);
or UO_751 (O_751,N_5198,N_6829);
xor UO_752 (O_752,N_6134,N_6955);
and UO_753 (O_753,N_5267,N_6827);
nor UO_754 (O_754,N_8311,N_9429);
nor UO_755 (O_755,N_7744,N_7362);
nand UO_756 (O_756,N_7320,N_5526);
nor UO_757 (O_757,N_7309,N_7037);
nor UO_758 (O_758,N_9735,N_5011);
nand UO_759 (O_759,N_7233,N_5947);
or UO_760 (O_760,N_8277,N_9312);
and UO_761 (O_761,N_6094,N_6585);
xor UO_762 (O_762,N_7682,N_6272);
or UO_763 (O_763,N_9868,N_6450);
nor UO_764 (O_764,N_5022,N_8314);
nand UO_765 (O_765,N_9883,N_7469);
or UO_766 (O_766,N_9749,N_5257);
and UO_767 (O_767,N_9120,N_9452);
and UO_768 (O_768,N_8276,N_9594);
nand UO_769 (O_769,N_6033,N_5774);
and UO_770 (O_770,N_6914,N_6441);
nand UO_771 (O_771,N_6375,N_8341);
nand UO_772 (O_772,N_8762,N_6673);
nand UO_773 (O_773,N_5431,N_6975);
and UO_774 (O_774,N_7074,N_5421);
nand UO_775 (O_775,N_8059,N_7413);
nor UO_776 (O_776,N_9831,N_6323);
or UO_777 (O_777,N_8764,N_8050);
and UO_778 (O_778,N_7581,N_8738);
nor UO_779 (O_779,N_7133,N_7257);
nor UO_780 (O_780,N_5340,N_8498);
and UO_781 (O_781,N_5591,N_5052);
nand UO_782 (O_782,N_6763,N_5303);
and UO_783 (O_783,N_9278,N_6756);
nand UO_784 (O_784,N_6868,N_6517);
or UO_785 (O_785,N_9676,N_6733);
nor UO_786 (O_786,N_5831,N_5522);
or UO_787 (O_787,N_5803,N_9161);
nor UO_788 (O_788,N_6046,N_6093);
nor UO_789 (O_789,N_8377,N_9154);
nor UO_790 (O_790,N_5508,N_7401);
and UO_791 (O_791,N_7810,N_7754);
or UO_792 (O_792,N_5700,N_5479);
or UO_793 (O_793,N_8585,N_8756);
or UO_794 (O_794,N_9153,N_7708);
and UO_795 (O_795,N_7022,N_5199);
or UO_796 (O_796,N_5484,N_7662);
and UO_797 (O_797,N_6730,N_8661);
nand UO_798 (O_798,N_5980,N_5680);
or UO_799 (O_799,N_8556,N_9926);
nor UO_800 (O_800,N_9984,N_5232);
and UO_801 (O_801,N_9506,N_5661);
nor UO_802 (O_802,N_5478,N_5341);
nor UO_803 (O_803,N_5907,N_6128);
or UO_804 (O_804,N_9561,N_8788);
or UO_805 (O_805,N_5137,N_7495);
nor UO_806 (O_806,N_5701,N_6356);
xnor UO_807 (O_807,N_9213,N_6553);
nor UO_808 (O_808,N_9178,N_7221);
nand UO_809 (O_809,N_9326,N_5013);
nand UO_810 (O_810,N_5274,N_5381);
nor UO_811 (O_811,N_8902,N_5445);
or UO_812 (O_812,N_5347,N_9177);
xnor UO_813 (O_813,N_6665,N_8613);
or UO_814 (O_814,N_6666,N_7698);
nor UO_815 (O_815,N_7894,N_6960);
nand UO_816 (O_816,N_5779,N_5465);
or UO_817 (O_817,N_8694,N_9159);
nand UO_818 (O_818,N_8986,N_8675);
nor UO_819 (O_819,N_5580,N_7976);
or UO_820 (O_820,N_7862,N_7305);
nand UO_821 (O_821,N_6890,N_7103);
nand UO_822 (O_822,N_5459,N_6391);
nor UO_823 (O_823,N_7896,N_9078);
or UO_824 (O_824,N_6125,N_9657);
nand UO_825 (O_825,N_8402,N_9011);
and UO_826 (O_826,N_8492,N_9500);
nand UO_827 (O_827,N_9046,N_6996);
nor UO_828 (O_828,N_8742,N_9487);
and UO_829 (O_829,N_9707,N_9469);
or UO_830 (O_830,N_7728,N_9595);
nand UO_831 (O_831,N_6001,N_7009);
xor UO_832 (O_832,N_5185,N_9144);
nand UO_833 (O_833,N_6250,N_7702);
xor UO_834 (O_834,N_7004,N_8123);
nor UO_835 (O_835,N_8625,N_5708);
nor UO_836 (O_836,N_9462,N_8048);
nand UO_837 (O_837,N_7489,N_8845);
and UO_838 (O_838,N_8851,N_8489);
nand UO_839 (O_839,N_7587,N_5684);
and UO_840 (O_840,N_8433,N_9768);
nand UO_841 (O_841,N_7827,N_8950);
nor UO_842 (O_842,N_6992,N_5163);
and UO_843 (O_843,N_5149,N_5926);
or UO_844 (O_844,N_6555,N_9408);
or UO_845 (O_845,N_8741,N_7186);
nand UO_846 (O_846,N_6806,N_5854);
nand UO_847 (O_847,N_9097,N_5386);
and UO_848 (O_848,N_9827,N_9430);
nand UO_849 (O_849,N_8628,N_7734);
nor UO_850 (O_850,N_5472,N_5997);
nor UO_851 (O_851,N_5759,N_7211);
and UO_852 (O_852,N_6908,N_7254);
nor UO_853 (O_853,N_9285,N_7235);
or UO_854 (O_854,N_9102,N_5128);
and UO_855 (O_855,N_7618,N_6574);
and UO_856 (O_856,N_5915,N_8864);
or UO_857 (O_857,N_7243,N_5518);
and UO_858 (O_858,N_7585,N_8136);
nand UO_859 (O_859,N_8317,N_6804);
or UO_860 (O_860,N_8232,N_7164);
or UO_861 (O_861,N_5325,N_8242);
and UO_862 (O_862,N_9976,N_9157);
or UO_863 (O_863,N_9552,N_8482);
nand UO_864 (O_864,N_6146,N_8115);
and UO_865 (O_865,N_7646,N_8980);
and UO_866 (O_866,N_5134,N_8374);
nor UO_867 (O_867,N_5638,N_8124);
and UO_868 (O_868,N_9722,N_8187);
nand UO_869 (O_869,N_5370,N_6070);
nor UO_870 (O_870,N_5621,N_8997);
or UO_871 (O_871,N_9952,N_7691);
or UO_872 (O_872,N_6495,N_8031);
or UO_873 (O_873,N_8206,N_9170);
and UO_874 (O_874,N_7416,N_5648);
or UO_875 (O_875,N_5634,N_5259);
and UO_876 (O_876,N_6658,N_7132);
nand UO_877 (O_877,N_9828,N_9044);
nand UO_878 (O_878,N_8092,N_8897);
nand UO_879 (O_879,N_7643,N_5456);
or UO_880 (O_880,N_5693,N_5703);
and UO_881 (O_881,N_6680,N_8580);
or UO_882 (O_882,N_5651,N_7030);
nand UO_883 (O_883,N_8278,N_5841);
nand UO_884 (O_884,N_8442,N_7177);
and UO_885 (O_885,N_8921,N_8779);
nor UO_886 (O_886,N_8497,N_5820);
nor UO_887 (O_887,N_6870,N_9716);
and UO_888 (O_888,N_7065,N_5268);
or UO_889 (O_889,N_8459,N_7614);
nand UO_890 (O_890,N_8994,N_9039);
and UO_891 (O_891,N_6803,N_8781);
or UO_892 (O_892,N_7048,N_7672);
or UO_893 (O_893,N_5489,N_8069);
nand UO_894 (O_894,N_9235,N_9387);
and UO_895 (O_895,N_7155,N_9167);
and UO_896 (O_896,N_8286,N_9658);
nor UO_897 (O_897,N_8805,N_5967);
and UO_898 (O_898,N_6100,N_8130);
or UO_899 (O_899,N_8843,N_5796);
nor UO_900 (O_900,N_5120,N_8981);
and UO_901 (O_901,N_7373,N_6422);
nor UO_902 (O_902,N_7980,N_5910);
or UO_903 (O_903,N_6427,N_5514);
nand UO_904 (O_904,N_6000,N_9028);
and UO_905 (O_905,N_9507,N_8013);
or UO_906 (O_906,N_6015,N_6109);
nor UO_907 (O_907,N_6696,N_5279);
nand UO_908 (O_908,N_5547,N_6200);
nand UO_909 (O_909,N_9416,N_7738);
nor UO_910 (O_910,N_8058,N_9317);
and UO_911 (O_911,N_6499,N_8872);
and UO_912 (O_912,N_7641,N_8834);
nor UO_913 (O_913,N_9491,N_7539);
or UO_914 (O_914,N_9600,N_8709);
nor UO_915 (O_915,N_9730,N_8064);
or UO_916 (O_916,N_5904,N_7031);
nand UO_917 (O_917,N_7178,N_6576);
nor UO_918 (O_918,N_5070,N_9776);
xor UO_919 (O_919,N_8919,N_5736);
nor UO_920 (O_920,N_9249,N_7989);
and UO_921 (O_921,N_8839,N_8942);
nand UO_922 (O_922,N_5911,N_9247);
or UO_923 (O_923,N_7090,N_5113);
and UO_924 (O_924,N_8739,N_9006);
nor UO_925 (O_925,N_6409,N_5894);
or UO_926 (O_926,N_9289,N_9175);
nor UO_927 (O_927,N_8218,N_9475);
nand UO_928 (O_928,N_5053,N_7485);
and UO_929 (O_929,N_5987,N_9375);
nand UO_930 (O_930,N_5069,N_5512);
and UO_931 (O_931,N_7668,N_5986);
and UO_932 (O_932,N_5529,N_7097);
or UO_933 (O_933,N_9534,N_8860);
nor UO_934 (O_934,N_6173,N_8702);
nand UO_935 (O_935,N_9558,N_6048);
or UO_936 (O_936,N_9350,N_5393);
or UO_937 (O_937,N_8837,N_5876);
nand UO_938 (O_938,N_8699,N_9334);
and UO_939 (O_939,N_6993,N_8765);
and UO_940 (O_940,N_8609,N_6148);
nand UO_941 (O_941,N_9325,N_9564);
nand UO_942 (O_942,N_7368,N_6582);
or UO_943 (O_943,N_6294,N_6983);
nor UO_944 (O_944,N_7527,N_9232);
and UO_945 (O_945,N_7059,N_7434);
nor UO_946 (O_946,N_5100,N_6351);
and UO_947 (O_947,N_6770,N_6607);
or UO_948 (O_948,N_8506,N_6538);
nand UO_949 (O_949,N_9365,N_8631);
and UO_950 (O_950,N_6287,N_9989);
and UO_951 (O_951,N_6653,N_8683);
and UO_952 (O_952,N_8928,N_6999);
nand UO_953 (O_953,N_8652,N_7747);
or UO_954 (O_954,N_5863,N_9715);
or UO_955 (O_955,N_9155,N_9512);
or UO_956 (O_956,N_7036,N_7568);
or UO_957 (O_957,N_6900,N_9296);
or UO_958 (O_958,N_6637,N_7869);
nand UO_959 (O_959,N_7444,N_7792);
or UO_960 (O_960,N_5617,N_5608);
or UO_961 (O_961,N_8693,N_6580);
nor UO_962 (O_962,N_9897,N_9513);
and UO_963 (O_963,N_5999,N_7013);
nor UO_964 (O_964,N_6815,N_5379);
or UO_965 (O_965,N_6529,N_6102);
nand UO_966 (O_966,N_5681,N_5115);
and UO_967 (O_967,N_8752,N_9886);
nor UO_968 (O_968,N_6545,N_5172);
or UO_969 (O_969,N_7705,N_9542);
nor UO_970 (O_970,N_6108,N_5505);
nand UO_971 (O_971,N_9038,N_6991);
or UO_972 (O_972,N_8883,N_5631);
nand UO_973 (O_973,N_5087,N_9821);
or UO_974 (O_974,N_7695,N_7284);
and UO_975 (O_975,N_6691,N_9244);
or UO_976 (O_976,N_5576,N_8140);
nor UO_977 (O_977,N_5105,N_9764);
nand UO_978 (O_978,N_9630,N_9322);
nor UO_979 (O_979,N_9651,N_7366);
nor UO_980 (O_980,N_7171,N_9587);
or UO_981 (O_981,N_7040,N_6994);
nor UO_982 (O_982,N_6987,N_8040);
nor UO_983 (O_983,N_6823,N_5219);
and UO_984 (O_984,N_7642,N_7324);
nor UO_985 (O_985,N_9603,N_5103);
nor UO_986 (O_986,N_9672,N_8416);
xnor UO_987 (O_987,N_8358,N_8772);
nand UO_988 (O_988,N_9119,N_7492);
or UO_989 (O_989,N_5385,N_8409);
nor UO_990 (O_990,N_7326,N_8318);
or UO_991 (O_991,N_8468,N_7670);
and UO_992 (O_992,N_7113,N_6812);
and UO_993 (O_993,N_5719,N_8330);
or UO_994 (O_994,N_9021,N_9686);
or UO_995 (O_995,N_7937,N_8734);
or UO_996 (O_996,N_6135,N_9270);
nor UO_997 (O_997,N_9551,N_5675);
or UO_998 (O_998,N_8995,N_7214);
xor UO_999 (O_999,N_9713,N_9796);
nand UO_1000 (O_1000,N_8768,N_9773);
xnor UO_1001 (O_1001,N_5539,N_5568);
or UO_1002 (O_1002,N_7158,N_7884);
or UO_1003 (O_1003,N_5545,N_8821);
or UO_1004 (O_1004,N_7969,N_7609);
or UO_1005 (O_1005,N_9386,N_6913);
nor UO_1006 (O_1006,N_8052,N_9995);
or UO_1007 (O_1007,N_6513,N_8095);
nand UO_1008 (O_1008,N_5293,N_6599);
or UO_1009 (O_1009,N_6820,N_7844);
or UO_1010 (O_1010,N_7925,N_9024);
and UO_1011 (O_1011,N_7100,N_8517);
nor UO_1012 (O_1012,N_9543,N_7286);
and UO_1013 (O_1013,N_7863,N_7244);
or UO_1014 (O_1014,N_5640,N_5753);
nand UO_1015 (O_1015,N_9019,N_9635);
or UO_1016 (O_1016,N_6473,N_6186);
nand UO_1017 (O_1017,N_6181,N_9866);
nand UO_1018 (O_1018,N_8181,N_5871);
nor UO_1019 (O_1019,N_8719,N_9560);
or UO_1020 (O_1020,N_8241,N_8701);
and UO_1021 (O_1021,N_8325,N_6238);
nand UO_1022 (O_1022,N_6449,N_5366);
or UO_1023 (O_1023,N_5114,N_5067);
or UO_1024 (O_1024,N_9683,N_8202);
and UO_1025 (O_1025,N_6729,N_5673);
and UO_1026 (O_1026,N_8952,N_6981);
and UO_1027 (O_1027,N_5942,N_5862);
nand UO_1028 (O_1028,N_6188,N_8465);
and UO_1029 (O_1029,N_5320,N_7664);
and UO_1030 (O_1030,N_5467,N_7173);
nand UO_1031 (O_1031,N_9328,N_7510);
nor UO_1032 (O_1032,N_8094,N_6261);
nor UO_1033 (O_1033,N_8939,N_7347);
nor UO_1034 (O_1034,N_5464,N_9463);
and UO_1035 (O_1035,N_5407,N_9076);
or UO_1036 (O_1036,N_7418,N_7229);
nor UO_1037 (O_1037,N_9269,N_7821);
nor UO_1038 (O_1038,N_5297,N_5133);
and UO_1039 (O_1039,N_9867,N_8673);
nand UO_1040 (O_1040,N_9123,N_8103);
and UO_1041 (O_1041,N_7711,N_5738);
or UO_1042 (O_1042,N_6099,N_5443);
or UO_1043 (O_1043,N_5929,N_7704);
nor UO_1044 (O_1044,N_6156,N_9501);
and UO_1045 (O_1045,N_9731,N_7448);
nand UO_1046 (O_1046,N_6668,N_7179);
and UO_1047 (O_1047,N_5988,N_8740);
or UO_1048 (O_1048,N_6911,N_5990);
and UO_1049 (O_1049,N_9977,N_6543);
or UO_1050 (O_1050,N_5793,N_6177);
nand UO_1051 (O_1051,N_6335,N_8138);
and UO_1052 (O_1052,N_5928,N_6077);
xor UO_1053 (O_1053,N_7964,N_7576);
or UO_1054 (O_1054,N_8334,N_8251);
and UO_1055 (O_1055,N_7957,N_7999);
nand UO_1056 (O_1056,N_9609,N_5200);
xor UO_1057 (O_1057,N_9338,N_5150);
or UO_1058 (O_1058,N_5108,N_8283);
or UO_1059 (O_1059,N_6624,N_8615);
and UO_1060 (O_1060,N_6616,N_7954);
nand UO_1061 (O_1061,N_8487,N_6266);
nor UO_1062 (O_1062,N_5280,N_9785);
nand UO_1063 (O_1063,N_9294,N_8922);
xnor UO_1064 (O_1064,N_7150,N_6631);
nor UO_1065 (O_1065,N_6500,N_7881);
or UO_1066 (O_1066,N_8004,N_9209);
or UO_1067 (O_1067,N_8029,N_7249);
or UO_1068 (O_1068,N_8830,N_8303);
or UO_1069 (O_1069,N_9197,N_6052);
nor UO_1070 (O_1070,N_6602,N_6547);
nor UO_1071 (O_1071,N_6478,N_8240);
nor UO_1072 (O_1072,N_7589,N_6252);
or UO_1073 (O_1073,N_5020,N_7560);
nor UO_1074 (O_1074,N_9443,N_9830);
nor UO_1075 (O_1075,N_6751,N_7422);
and UO_1076 (O_1076,N_7648,N_9746);
nor UO_1077 (O_1077,N_8381,N_9787);
and UO_1078 (O_1078,N_7436,N_6988);
and UO_1079 (O_1079,N_5972,N_7203);
nand UO_1080 (O_1080,N_6253,N_6256);
and UO_1081 (O_1081,N_8578,N_7683);
and UO_1082 (O_1082,N_8512,N_5654);
nor UO_1083 (O_1083,N_7639,N_6273);
nor UO_1084 (O_1084,N_9316,N_8710);
nand UO_1085 (O_1085,N_5182,N_9598);
nand UO_1086 (O_1086,N_7061,N_6927);
and UO_1087 (O_1087,N_5136,N_7072);
xnor UO_1088 (O_1088,N_6399,N_9599);
nor UO_1089 (O_1089,N_9931,N_7557);
nor UO_1090 (O_1090,N_5946,N_9378);
nor UO_1091 (O_1091,N_7654,N_9489);
nor UO_1092 (O_1092,N_8472,N_8205);
or UO_1093 (O_1093,N_9521,N_8840);
nor UO_1094 (O_1094,N_8555,N_7143);
nor UO_1095 (O_1095,N_8102,N_6053);
or UO_1096 (O_1096,N_6091,N_5696);
nand UO_1097 (O_1097,N_5933,N_5826);
nor UO_1098 (O_1098,N_5495,N_6632);
nor UO_1099 (O_1099,N_9574,N_6302);
nand UO_1100 (O_1100,N_6884,N_9631);
nor UO_1101 (O_1101,N_6226,N_6355);
or UO_1102 (O_1102,N_8154,N_9502);
or UO_1103 (O_1103,N_7684,N_9356);
and UO_1104 (O_1104,N_7219,N_7247);
nand UO_1105 (O_1105,N_5139,N_5963);
nand UO_1106 (O_1106,N_6858,N_8918);
nand UO_1107 (O_1107,N_9632,N_8162);
and UO_1108 (O_1108,N_9018,N_7603);
nand UO_1109 (O_1109,N_7008,N_6675);
nor UO_1110 (O_1110,N_8657,N_9403);
nand UO_1111 (O_1111,N_7265,N_9793);
nand UO_1112 (O_1112,N_5958,N_8076);
nand UO_1113 (O_1113,N_9579,N_5063);
xor UO_1114 (O_1114,N_8090,N_9671);
or UO_1115 (O_1115,N_5383,N_5780);
or UO_1116 (O_1116,N_6862,N_7236);
nand UO_1117 (O_1117,N_7480,N_7938);
and UO_1118 (O_1118,N_5900,N_5869);
nor UO_1119 (O_1119,N_9901,N_6085);
nand UO_1120 (O_1120,N_5860,N_7720);
nand UO_1121 (O_1121,N_7781,N_9496);
and UO_1122 (O_1122,N_7381,N_9040);
nand UO_1123 (O_1123,N_9013,N_9253);
nor UO_1124 (O_1124,N_9674,N_8961);
nand UO_1125 (O_1125,N_8400,N_6475);
nor UO_1126 (O_1126,N_7388,N_9583);
and UO_1127 (O_1127,N_6368,N_5600);
nand UO_1128 (O_1128,N_9862,N_6019);
or UO_1129 (O_1129,N_9458,N_9017);
nand UO_1130 (O_1130,N_6353,N_9808);
or UO_1131 (O_1131,N_7766,N_9003);
or UO_1132 (O_1132,N_6258,N_7893);
and UO_1133 (O_1133,N_7083,N_7184);
and UO_1134 (O_1134,N_7242,N_5969);
and UO_1135 (O_1135,N_5940,N_5313);
nand UO_1136 (O_1136,N_6923,N_8055);
nor UO_1137 (O_1137,N_5805,N_6937);
and UO_1138 (O_1138,N_6042,N_6029);
nand UO_1139 (O_1139,N_9095,N_9703);
nand UO_1140 (O_1140,N_6501,N_9734);
xnor UO_1141 (O_1141,N_6852,N_6032);
and UO_1142 (O_1142,N_7507,N_9835);
nand UO_1143 (O_1143,N_9052,N_9397);
nand UO_1144 (O_1144,N_6819,N_5709);
and UO_1145 (O_1145,N_9508,N_8326);
nand UO_1146 (O_1146,N_5991,N_7450);
nand UO_1147 (O_1147,N_8012,N_8336);
nand UO_1148 (O_1148,N_8046,N_9442);
or UO_1149 (O_1149,N_9720,N_7666);
or UO_1150 (O_1150,N_6794,N_7488);
xor UO_1151 (O_1151,N_9522,N_6817);
or UO_1152 (O_1152,N_6434,N_5666);
nor UO_1153 (O_1153,N_5657,N_5721);
or UO_1154 (O_1154,N_8203,N_6472);
nor UO_1155 (O_1155,N_6710,N_9955);
and UO_1156 (O_1156,N_8712,N_8216);
or UO_1157 (O_1157,N_6248,N_7085);
and UO_1158 (O_1158,N_7751,N_7553);
or UO_1159 (O_1159,N_8798,N_8349);
nor UO_1160 (O_1160,N_5757,N_9307);
and UO_1161 (O_1161,N_6452,N_7296);
or UO_1162 (O_1162,N_7597,N_5287);
or UO_1163 (O_1163,N_9068,N_8646);
and UO_1164 (O_1164,N_7950,N_8562);
and UO_1165 (O_1165,N_5156,N_6917);
and UO_1166 (O_1166,N_9047,N_6811);
nor UO_1167 (O_1167,N_7637,N_6797);
and UO_1168 (O_1168,N_7873,N_5650);
nor UO_1169 (O_1169,N_9909,N_9981);
nor UO_1170 (O_1170,N_9621,N_5949);
and UO_1171 (O_1171,N_5408,N_7240);
and UO_1172 (O_1172,N_6213,N_8265);
nand UO_1173 (O_1173,N_9406,N_9048);
nor UO_1174 (O_1174,N_6388,N_8191);
and UO_1175 (O_1175,N_5333,N_7339);
or UO_1176 (O_1176,N_8190,N_8515);
nor UO_1177 (O_1177,N_5446,N_8963);
and UO_1178 (O_1178,N_5434,N_7567);
or UO_1179 (O_1179,N_9314,N_8587);
nor UO_1180 (O_1180,N_6896,N_7398);
nor UO_1181 (O_1181,N_8707,N_6338);
or UO_1182 (O_1182,N_8479,N_7583);
nor UO_1183 (O_1183,N_8028,N_8252);
or UO_1184 (O_1184,N_7279,N_6405);
and UO_1185 (O_1185,N_6810,N_8998);
and UO_1186 (O_1186,N_5265,N_5642);
nand UO_1187 (O_1187,N_9548,N_5075);
and UO_1188 (O_1188,N_7124,N_5601);
nand UO_1189 (O_1189,N_5633,N_9854);
xnor UO_1190 (O_1190,N_7621,N_8956);
or UO_1191 (O_1191,N_6537,N_8809);
and UO_1192 (O_1192,N_6922,N_5197);
nand UO_1193 (O_1193,N_5974,N_8010);
nand UO_1194 (O_1194,N_8570,N_7407);
nand UO_1195 (O_1195,N_6638,N_7529);
and UO_1196 (O_1196,N_9111,N_5089);
and UO_1197 (O_1197,N_9025,N_8499);
or UO_1198 (O_1198,N_5255,N_6466);
nor UO_1199 (O_1199,N_5748,N_6840);
and UO_1200 (O_1200,N_8820,N_8863);
nand UO_1201 (O_1201,N_6831,N_6082);
and UO_1202 (O_1202,N_9198,N_5902);
nand UO_1203 (O_1203,N_5973,N_6451);
and UO_1204 (O_1204,N_8769,N_8671);
and UO_1205 (O_1205,N_6874,N_9229);
nand UO_1206 (O_1206,N_9559,N_7359);
nand UO_1207 (O_1207,N_7273,N_9221);
xnor UO_1208 (O_1208,N_6358,N_9412);
and UO_1209 (O_1209,N_7571,N_7726);
nand UO_1210 (O_1210,N_6176,N_9807);
nor UO_1211 (O_1211,N_9023,N_9149);
nor UO_1212 (O_1212,N_5107,N_9766);
and UO_1213 (O_1213,N_8263,N_9112);
and UO_1214 (O_1214,N_5936,N_5360);
or UO_1215 (O_1215,N_7419,N_9954);
and UO_1216 (O_1216,N_6428,N_7515);
and UO_1217 (O_1217,N_7687,N_8463);
nand UO_1218 (O_1218,N_5302,N_6058);
or UO_1219 (O_1219,N_5093,N_8859);
nand UO_1220 (O_1220,N_9973,N_6468);
and UO_1221 (O_1221,N_7064,N_9922);
and UO_1222 (O_1222,N_5844,N_8045);
nor UO_1223 (O_1223,N_5658,N_8896);
or UO_1224 (O_1224,N_9988,N_7137);
and UO_1225 (O_1225,N_8670,N_5839);
nor UO_1226 (O_1226,N_5937,N_9900);
and UO_1227 (O_1227,N_7355,N_6774);
and UO_1228 (O_1228,N_7577,N_8144);
and UO_1229 (O_1229,N_8689,N_8744);
or UO_1230 (O_1230,N_7959,N_6101);
or UO_1231 (O_1231,N_6055,N_6026);
and UO_1232 (O_1232,N_9495,N_8146);
or UO_1233 (O_1233,N_9829,N_7331);
nor UO_1234 (O_1234,N_6010,N_9072);
nand UO_1235 (O_1235,N_7871,N_5469);
nand UO_1236 (O_1236,N_5801,N_7016);
or UO_1237 (O_1237,N_6066,N_5010);
nand UO_1238 (O_1238,N_5585,N_8684);
or UO_1239 (O_1239,N_6382,N_9493);
or UO_1240 (O_1240,N_7703,N_6354);
and UO_1241 (O_1241,N_8868,N_9311);
nor UO_1242 (O_1242,N_6792,N_6095);
or UO_1243 (O_1243,N_7922,N_7404);
nor UO_1244 (O_1244,N_8733,N_7870);
nand UO_1245 (O_1245,N_8364,N_6776);
xor UO_1246 (O_1246,N_9461,N_9681);
nor UO_1247 (O_1247,N_6147,N_9352);
nor UO_1248 (O_1248,N_7172,N_9964);
nor UO_1249 (O_1249,N_9625,N_9965);
and UO_1250 (O_1250,N_7387,N_5482);
or UO_1251 (O_1251,N_8500,N_6736);
nor UO_1252 (O_1252,N_7315,N_6158);
and UO_1253 (O_1253,N_9376,N_6841);
nand UO_1254 (O_1254,N_7120,N_8053);
and UO_1255 (O_1255,N_8841,N_9212);
and UO_1256 (O_1256,N_5843,N_9607);
nand UO_1257 (O_1257,N_5614,N_5586);
nand UO_1258 (O_1258,N_7645,N_7110);
nor UO_1259 (O_1259,N_8167,N_8194);
xor UO_1260 (O_1260,N_7543,N_7514);
nor UO_1261 (O_1261,N_9103,N_6219);
nor UO_1262 (O_1262,N_7380,N_8038);
nand UO_1263 (O_1263,N_6966,N_5296);
nand UO_1264 (O_1264,N_8966,N_5955);
or UO_1265 (O_1265,N_8885,N_9271);
nand UO_1266 (O_1266,N_8826,N_7554);
nand UO_1267 (O_1267,N_5349,N_8160);
xnor UO_1268 (O_1268,N_7681,N_5733);
nand UO_1269 (O_1269,N_7769,N_7348);
nand UO_1270 (O_1270,N_7732,N_8906);
nor UO_1271 (O_1271,N_7092,N_5440);
nor UO_1272 (O_1272,N_5867,N_7709);
or UO_1273 (O_1273,N_8688,N_7099);
nor UO_1274 (O_1274,N_9728,N_6747);
and UO_1275 (O_1275,N_8305,N_6247);
nand UO_1276 (O_1276,N_5212,N_8541);
and UO_1277 (O_1277,N_9790,N_6025);
or UO_1278 (O_1278,N_5858,N_8551);
nand UO_1279 (O_1279,N_7556,N_7617);
or UO_1280 (O_1280,N_7879,N_6514);
or UO_1281 (O_1281,N_6313,N_7538);
and UO_1282 (O_1282,N_6332,N_8951);
nand UO_1283 (O_1283,N_5678,N_6620);
nand UO_1284 (O_1284,N_9702,N_6244);
nor UO_1285 (O_1285,N_5535,N_5917);
nand UO_1286 (O_1286,N_8521,N_6883);
and UO_1287 (O_1287,N_8911,N_8727);
and UO_1288 (O_1288,N_9371,N_9476);
nor UO_1289 (O_1289,N_7983,N_8386);
nand UO_1290 (O_1290,N_9395,N_5546);
nor UO_1291 (O_1291,N_8899,N_6645);
and UO_1292 (O_1292,N_8930,N_5081);
and UO_1293 (O_1293,N_9012,N_5982);
nor UO_1294 (O_1294,N_8780,N_9524);
nand UO_1295 (O_1295,N_6724,N_8636);
nand UO_1296 (O_1296,N_8647,N_8870);
or UO_1297 (O_1297,N_6600,N_5436);
or UO_1298 (O_1298,N_7855,N_8525);
and UO_1299 (O_1299,N_6581,N_5952);
and UO_1300 (O_1300,N_6685,N_9624);
or UO_1301 (O_1301,N_9124,N_6251);
nor UO_1302 (O_1302,N_6570,N_7301);
nand UO_1303 (O_1303,N_5414,N_9698);
nor UO_1304 (O_1304,N_9619,N_8767);
nor UO_1305 (O_1305,N_7675,N_7383);
nand UO_1306 (O_1306,N_5698,N_8106);
or UO_1307 (O_1307,N_7946,N_9079);
or UO_1308 (O_1308,N_7205,N_8743);
and UO_1309 (O_1309,N_8268,N_7197);
or UO_1310 (O_1310,N_7805,N_5985);
and UO_1311 (O_1311,N_9692,N_8822);
nand UO_1312 (O_1312,N_6563,N_9354);
nand UO_1313 (O_1313,N_9266,N_7521);
and UO_1314 (O_1314,N_9182,N_7503);
and UO_1315 (O_1315,N_6465,N_7758);
xnor UO_1316 (O_1316,N_7477,N_8244);
and UO_1317 (O_1317,N_6051,N_9578);
or UO_1318 (O_1318,N_6224,N_8389);
nor UO_1319 (O_1319,N_6544,N_7540);
and UO_1320 (O_1320,N_9359,N_5743);
or UO_1321 (O_1321,N_9864,N_6834);
or UO_1322 (O_1322,N_7830,N_8258);
xnor UO_1323 (O_1323,N_7693,N_7824);
nor UO_1324 (O_1324,N_7468,N_9214);
and UO_1325 (O_1325,N_8887,N_5598);
and UO_1326 (O_1326,N_9457,N_8620);
nand UO_1327 (O_1327,N_9663,N_5059);
nor UO_1328 (O_1328,N_8293,N_8478);
and UO_1329 (O_1329,N_8371,N_9729);
and UO_1330 (O_1330,N_6916,N_7591);
or UO_1331 (O_1331,N_9596,N_7630);
and UO_1332 (O_1332,N_5098,N_9724);
or UO_1333 (O_1333,N_6357,N_7274);
and UO_1334 (O_1334,N_8282,N_9050);
nand UO_1335 (O_1335,N_9432,N_7250);
and UO_1336 (O_1336,N_7652,N_8686);
nand UO_1337 (O_1337,N_7825,N_8444);
nand UO_1338 (O_1338,N_5925,N_8737);
or UO_1339 (O_1339,N_5639,N_8786);
and UO_1340 (O_1340,N_7053,N_5814);
nand UO_1341 (O_1341,N_7135,N_6208);
and UO_1342 (O_1342,N_6950,N_9310);
and UO_1343 (O_1343,N_7452,N_6288);
nand UO_1344 (O_1344,N_8829,N_6319);
nand UO_1345 (O_1345,N_9099,N_6320);
nor UO_1346 (O_1346,N_7828,N_7046);
nand UO_1347 (O_1347,N_8309,N_6899);
nand UO_1348 (O_1348,N_5001,N_5369);
nor UO_1349 (O_1349,N_9417,N_5749);
nand UO_1350 (O_1350,N_5475,N_9752);
nor UO_1351 (O_1351,N_7592,N_5712);
xor UO_1352 (O_1352,N_5458,N_8576);
and UO_1353 (O_1353,N_6345,N_6275);
xnor UO_1354 (O_1354,N_6596,N_6965);
nand UO_1355 (O_1355,N_7689,N_5166);
and UO_1356 (O_1356,N_7025,N_6534);
nor UO_1357 (O_1357,N_5534,N_6526);
nor UO_1358 (O_1358,N_9126,N_8107);
nand UO_1359 (O_1359,N_8866,N_7895);
nand UO_1360 (O_1360,N_6964,N_5822);
nor UO_1361 (O_1361,N_7657,N_5468);
xor UO_1362 (O_1362,N_5745,N_5427);
nor UO_1363 (O_1363,N_6078,N_6378);
nand UO_1364 (O_1364,N_5931,N_8047);
nand UO_1365 (O_1365,N_5029,N_6462);
nand UO_1366 (O_1366,N_6464,N_7139);
and UO_1367 (O_1367,N_9818,N_7327);
and UO_1368 (O_1368,N_9422,N_9673);
nor UO_1369 (O_1369,N_9219,N_7191);
nor UO_1370 (O_1370,N_5677,N_9464);
nor UO_1371 (O_1371,N_6569,N_8288);
nor UO_1372 (O_1372,N_6004,N_8170);
and UO_1373 (O_1373,N_9951,N_8790);
nor UO_1374 (O_1374,N_9020,N_7089);
nand UO_1375 (O_1375,N_7787,N_7151);
nor UO_1376 (O_1376,N_5336,N_8266);
and UO_1377 (O_1377,N_6190,N_7518);
nand UO_1378 (O_1378,N_8246,N_9368);
or UO_1379 (O_1379,N_7255,N_5373);
or UO_1380 (O_1380,N_8991,N_9691);
and UO_1381 (O_1381,N_8184,N_5354);
or UO_1382 (O_1382,N_8304,N_7453);
nor UO_1383 (O_1383,N_7988,N_8476);
or UO_1384 (O_1384,N_7811,N_5788);
or UO_1385 (O_1385,N_5396,N_9653);
or UO_1386 (O_1386,N_6169,N_9114);
nand UO_1387 (O_1387,N_8533,N_8204);
or UO_1388 (O_1388,N_6798,N_5009);
nand UO_1389 (O_1389,N_8907,N_9148);
nor UO_1390 (O_1390,N_5727,N_6515);
nand UO_1391 (O_1391,N_5248,N_8626);
nand UO_1392 (O_1392,N_7349,N_7269);
and UO_1393 (O_1393,N_5879,N_5335);
or UO_1394 (O_1394,N_6431,N_8706);
or UO_1395 (O_1395,N_6670,N_7607);
and UO_1396 (O_1396,N_6539,N_9767);
nor UO_1397 (O_1397,N_5122,N_9727);
nor UO_1398 (O_1398,N_6636,N_6943);
or UO_1399 (O_1399,N_9929,N_9239);
nand UO_1400 (O_1400,N_8071,N_9520);
or UO_1401 (O_1401,N_9896,N_8509);
and UO_1402 (O_1402,N_6503,N_6076);
nand UO_1403 (O_1403,N_9041,N_8600);
and UO_1404 (O_1404,N_7888,N_7024);
nor UO_1405 (O_1405,N_8846,N_6290);
nand UO_1406 (O_1406,N_6603,N_8289);
nand UO_1407 (O_1407,N_7602,N_9355);
nor UO_1408 (O_1408,N_7188,N_8890);
or UO_1409 (O_1409,N_8005,N_5030);
nand UO_1410 (O_1410,N_7548,N_6065);
nor UO_1411 (O_1411,N_9572,N_5367);
and UO_1412 (O_1412,N_6285,N_8964);
or UO_1413 (O_1413,N_8962,N_7849);
nor UO_1414 (O_1414,N_5315,N_8593);
or UO_1415 (O_1415,N_5857,N_5939);
nand UO_1416 (O_1416,N_7671,N_9817);
and UO_1417 (O_1417,N_9890,N_9360);
nor UO_1418 (O_1418,N_6877,N_8800);
nand UO_1419 (O_1419,N_9036,N_9399);
nor UO_1420 (O_1420,N_8813,N_8039);
nor UO_1421 (O_1421,N_8973,N_6136);
or UO_1422 (O_1422,N_9483,N_8401);
nand UO_1423 (O_1423,N_8750,N_5169);
or UO_1424 (O_1424,N_7334,N_6096);
xnor UO_1425 (O_1425,N_6742,N_6267);
and UO_1426 (O_1426,N_7470,N_8924);
xnor UO_1427 (O_1427,N_7482,N_7323);
nand UO_1428 (O_1428,N_8573,N_7679);
nand UO_1429 (O_1429,N_7258,N_7248);
nand UO_1430 (O_1430,N_6149,N_7222);
or UO_1431 (O_1431,N_5430,N_7992);
nand UO_1432 (O_1432,N_8753,N_8422);
xor UO_1433 (O_1433,N_9303,N_6283);
nor UO_1434 (O_1434,N_7080,N_8446);
or UO_1435 (O_1435,N_5374,N_5751);
nand UO_1436 (O_1436,N_9636,N_5707);
nand UO_1437 (O_1437,N_6492,N_6595);
nand UO_1438 (O_1438,N_7517,N_6243);
or UO_1439 (O_1439,N_9652,N_6279);
nand UO_1440 (O_1440,N_7336,N_5304);
and UO_1441 (O_1441,N_7790,N_5756);
nand UO_1442 (O_1442,N_9486,N_7462);
or UO_1443 (O_1443,N_6948,N_8036);
or UO_1444 (O_1444,N_9669,N_5389);
and UO_1445 (O_1445,N_6459,N_7635);
and UO_1446 (O_1446,N_8955,N_7378);
nand UO_1447 (O_1447,N_6227,N_5729);
nand UO_1448 (O_1448,N_8728,N_9184);
or UO_1449 (O_1449,N_5388,N_9855);
or UO_1450 (O_1450,N_6968,N_9539);
or UO_1451 (O_1451,N_7604,N_6194);
or UO_1452 (O_1452,N_6865,N_9205);
nand UO_1453 (O_1453,N_7134,N_8173);
or UO_1454 (O_1454,N_7842,N_6420);
nor UO_1455 (O_1455,N_9234,N_5832);
nor UO_1456 (O_1456,N_9639,N_9132);
nor UO_1457 (O_1457,N_9207,N_8189);
nor UO_1458 (O_1458,N_7020,N_5809);
or UO_1459 (O_1459,N_8529,N_9517);
nor UO_1460 (O_1460,N_7330,N_8720);
nor UO_1461 (O_1461,N_5092,N_8026);
or UO_1462 (O_1462,N_7212,N_5339);
nand UO_1463 (O_1463,N_9405,N_7718);
or UO_1464 (O_1464,N_9255,N_7903);
or UO_1465 (O_1465,N_5837,N_7838);
and UO_1466 (O_1466,N_9775,N_9850);
and UO_1467 (O_1467,N_7864,N_5209);
nor UO_1468 (O_1468,N_7908,N_9374);
nand UO_1469 (O_1469,N_5493,N_6998);
or UO_1470 (O_1470,N_8532,N_8960);
or UO_1471 (O_1471,N_5819,N_8618);
or UO_1472 (O_1472,N_7660,N_7415);
and UO_1473 (O_1473,N_5289,N_9176);
or UO_1474 (O_1474,N_7936,N_7627);
or UO_1475 (O_1475,N_7289,N_8332);
and UO_1476 (O_1476,N_9792,N_7531);
and UO_1477 (O_1477,N_6415,N_9320);
and UO_1478 (O_1478,N_7044,N_5007);
nor UO_1479 (O_1479,N_6021,N_5609);
or UO_1480 (O_1480,N_7653,N_7213);
nor UO_1481 (O_1481,N_9222,N_7295);
nand UO_1482 (O_1482,N_7697,N_9759);
or UO_1483 (O_1483,N_7230,N_7234);
nor UO_1484 (O_1484,N_6432,N_9151);
nor UO_1485 (O_1485,N_7836,N_9823);
nand UO_1486 (O_1486,N_6299,N_7685);
and UO_1487 (O_1487,N_7730,N_5842);
or UO_1488 (O_1488,N_6402,N_6433);
nand UO_1489 (O_1489,N_9105,N_5041);
nor UO_1490 (O_1490,N_5884,N_5885);
nor UO_1491 (O_1491,N_8209,N_9497);
and UO_1492 (O_1492,N_8405,N_8785);
nand UO_1493 (O_1493,N_8970,N_8152);
nand UO_1494 (O_1494,N_5877,N_5260);
or UO_1495 (O_1495,N_7843,N_6317);
nor UO_1496 (O_1496,N_5908,N_9536);
xor UO_1497 (O_1497,N_6789,N_8417);
nand UO_1498 (O_1498,N_8878,N_5343);
and UO_1499 (O_1499,N_7181,N_6394);
endmodule