module basic_3000_30000_3500_150_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2592,In_2742);
nor U1 (N_1,In_9,In_109);
and U2 (N_2,In_2893,In_123);
xor U3 (N_3,In_1706,In_1301);
xor U4 (N_4,In_1758,In_2671);
and U5 (N_5,In_1853,In_373);
or U6 (N_6,In_2032,In_736);
nand U7 (N_7,In_2853,In_2276);
nand U8 (N_8,In_1942,In_1736);
or U9 (N_9,In_2808,In_748);
nor U10 (N_10,In_949,In_56);
or U11 (N_11,In_2133,In_1459);
xor U12 (N_12,In_1303,In_1966);
nand U13 (N_13,In_2342,In_2394);
or U14 (N_14,In_1183,In_2116);
or U15 (N_15,In_2249,In_2542);
and U16 (N_16,In_2156,In_2121);
or U17 (N_17,In_1881,In_1198);
xor U18 (N_18,In_103,In_2423);
xor U19 (N_19,In_1211,In_2987);
nand U20 (N_20,In_943,In_1691);
or U21 (N_21,In_1530,In_1813);
nor U22 (N_22,In_2044,In_1484);
or U23 (N_23,In_2840,In_1431);
or U24 (N_24,In_236,In_1118);
xnor U25 (N_25,In_267,In_2502);
and U26 (N_26,In_2930,In_711);
xor U27 (N_27,In_2387,In_356);
or U28 (N_28,In_2645,In_1392);
nand U29 (N_29,In_1564,In_251);
xnor U30 (N_30,In_1039,In_1056);
nor U31 (N_31,In_2662,In_2678);
nor U32 (N_32,In_1250,In_1058);
or U33 (N_33,In_1962,In_810);
nor U34 (N_34,In_2038,In_604);
nor U35 (N_35,In_1831,In_1059);
and U36 (N_36,In_1571,In_746);
nor U37 (N_37,In_211,In_2880);
xor U38 (N_38,In_146,In_2218);
and U39 (N_39,In_309,In_695);
nor U40 (N_40,In_1465,In_1871);
xnor U41 (N_41,In_532,In_1414);
nor U42 (N_42,In_2685,In_634);
nand U43 (N_43,In_2011,In_2246);
nand U44 (N_44,In_2408,In_2475);
and U45 (N_45,In_889,In_322);
xor U46 (N_46,In_1395,In_865);
and U47 (N_47,In_2527,In_1947);
nor U48 (N_48,In_1113,In_2864);
xor U49 (N_49,In_2281,In_2078);
or U50 (N_50,In_2848,In_2779);
nor U51 (N_51,In_1620,In_2457);
or U52 (N_52,In_2179,In_2042);
and U53 (N_53,In_1473,In_199);
or U54 (N_54,In_1950,In_1681);
nor U55 (N_55,In_1151,In_854);
or U56 (N_56,In_830,In_1389);
nor U57 (N_57,In_690,In_1130);
or U58 (N_58,In_1913,In_603);
or U59 (N_59,In_2730,In_1240);
or U60 (N_60,In_2867,In_1196);
xnor U61 (N_61,In_1667,In_1391);
nor U62 (N_62,In_2902,In_2557);
nor U63 (N_63,In_2320,In_2316);
or U64 (N_64,In_589,In_281);
xnor U65 (N_65,In_2154,In_765);
and U66 (N_66,In_105,In_1738);
nor U67 (N_67,In_586,In_2759);
or U68 (N_68,In_659,In_2503);
nor U69 (N_69,In_565,In_122);
or U70 (N_70,In_2396,In_2569);
xnor U71 (N_71,In_2398,In_1908);
and U72 (N_72,In_2973,In_1889);
nor U73 (N_73,In_1293,In_2184);
nand U74 (N_74,In_2755,In_241);
nor U75 (N_75,In_2882,In_1849);
nand U76 (N_76,In_2174,In_2447);
nand U77 (N_77,In_1108,In_1649);
xnor U78 (N_78,In_2980,In_1404);
or U79 (N_79,In_1133,In_1504);
xnor U80 (N_80,In_707,In_2288);
nor U81 (N_81,In_599,In_958);
xnor U82 (N_82,In_1514,In_2574);
nand U83 (N_83,In_2776,In_349);
nand U84 (N_84,In_230,In_2516);
nand U85 (N_85,In_304,In_2014);
xor U86 (N_86,In_519,In_2676);
and U87 (N_87,In_2695,In_272);
nand U88 (N_88,In_2745,In_2054);
and U89 (N_89,In_1223,In_2787);
nor U90 (N_90,In_2362,In_1621);
and U91 (N_91,In_2957,In_1943);
or U92 (N_92,In_2140,In_2245);
or U93 (N_93,In_1317,In_1906);
and U94 (N_94,In_2737,In_1783);
nor U95 (N_95,In_2635,In_2319);
and U96 (N_96,In_1013,In_861);
and U97 (N_97,In_2725,In_1280);
xnor U98 (N_98,In_294,In_588);
and U99 (N_99,In_25,In_214);
nand U100 (N_100,In_1353,In_1606);
nand U101 (N_101,In_1340,In_508);
or U102 (N_102,In_478,In_517);
and U103 (N_103,In_1919,In_273);
and U104 (N_104,In_2169,In_1489);
xnor U105 (N_105,In_1161,In_2188);
xor U106 (N_106,In_2955,In_1442);
nand U107 (N_107,In_2749,In_697);
nand U108 (N_108,In_582,In_2899);
or U109 (N_109,In_310,In_1552);
nor U110 (N_110,In_1413,In_2104);
or U111 (N_111,In_2310,In_2918);
nor U112 (N_112,In_2390,In_142);
nand U113 (N_113,In_511,In_2);
nor U114 (N_114,In_2598,In_60);
and U115 (N_115,In_2177,In_646);
xor U116 (N_116,In_1883,In_1318);
nand U117 (N_117,In_527,In_1337);
and U118 (N_118,In_842,In_999);
xor U119 (N_119,In_1653,In_348);
xor U120 (N_120,In_2572,In_97);
and U121 (N_121,In_2293,In_740);
nand U122 (N_122,In_2139,In_2106);
and U123 (N_123,In_128,In_694);
and U124 (N_124,In_691,In_2798);
nand U125 (N_125,In_846,In_2460);
xor U126 (N_126,In_2380,In_425);
nand U127 (N_127,In_1643,In_483);
nand U128 (N_128,In_203,In_2581);
or U129 (N_129,In_140,In_1580);
and U130 (N_130,In_2356,In_2649);
nor U131 (N_131,In_1440,In_2476);
nand U132 (N_132,In_1265,In_1622);
xor U133 (N_133,In_314,In_29);
or U134 (N_134,In_259,In_2528);
nor U135 (N_135,In_2883,In_1125);
nand U136 (N_136,In_2865,In_1583);
or U137 (N_137,In_709,In_2110);
nor U138 (N_138,In_2182,In_2778);
nand U139 (N_139,In_1312,In_978);
nand U140 (N_140,In_2624,In_876);
nand U141 (N_141,In_1253,In_1602);
or U142 (N_142,In_1278,In_1614);
xor U143 (N_143,In_1061,In_2895);
nand U144 (N_144,In_486,In_1266);
or U145 (N_145,In_817,In_1642);
nor U146 (N_146,In_1714,In_1037);
or U147 (N_147,In_205,In_790);
or U148 (N_148,In_1102,In_474);
and U149 (N_149,In_188,In_2125);
and U150 (N_150,In_57,In_1448);
and U151 (N_151,In_952,In_2782);
nand U152 (N_152,In_13,In_2046);
and U153 (N_153,In_1855,In_1662);
and U154 (N_154,In_1613,In_738);
nand U155 (N_155,In_993,In_473);
xor U156 (N_156,In_1717,In_685);
xor U157 (N_157,In_1210,In_2661);
or U158 (N_158,In_2199,In_643);
nand U159 (N_159,In_2185,In_252);
nand U160 (N_160,In_2146,In_2606);
and U161 (N_161,In_2001,In_1388);
and U162 (N_162,In_117,In_1903);
or U163 (N_163,In_1468,In_1308);
nor U164 (N_164,In_15,In_1986);
and U165 (N_165,In_1399,In_1647);
nand U166 (N_166,In_476,In_641);
nor U167 (N_167,In_1426,In_1296);
or U168 (N_168,In_334,In_648);
and U169 (N_169,In_1619,In_800);
and U170 (N_170,In_149,In_786);
nor U171 (N_171,In_1267,In_916);
nor U172 (N_172,In_2300,In_2709);
or U173 (N_173,In_1336,In_684);
or U174 (N_174,In_2859,In_201);
nor U175 (N_175,In_2385,In_670);
xnor U176 (N_176,In_2171,In_2571);
and U177 (N_177,In_1748,In_372);
nand U178 (N_178,In_2195,In_1115);
or U179 (N_179,In_1684,In_966);
xor U180 (N_180,In_2545,In_2215);
nand U181 (N_181,In_2453,In_1818);
nand U182 (N_182,In_86,In_2752);
xor U183 (N_183,In_111,In_879);
xnor U184 (N_184,In_824,In_701);
or U185 (N_185,In_2167,In_2478);
or U186 (N_186,In_1859,In_1518);
or U187 (N_187,In_1705,In_1633);
xnor U188 (N_188,In_152,In_1900);
or U189 (N_189,In_455,In_2159);
xnor U190 (N_190,In_1026,In_1138);
and U191 (N_191,In_1496,In_615);
and U192 (N_192,In_551,In_387);
nor U193 (N_193,In_852,In_1073);
and U194 (N_194,In_1631,In_1584);
nand U195 (N_195,In_233,In_1599);
xor U196 (N_196,In_1321,In_1260);
xor U197 (N_197,In_1424,In_2541);
nor U198 (N_198,In_2280,In_2242);
nand U199 (N_199,In_1023,In_1241);
xor U200 (N_200,In_2582,In_1628);
nand U201 (N_201,In_189,In_1611);
and U202 (N_202,In_1998,In_1227);
or U203 (N_203,In_2439,In_2713);
and U204 (N_204,In_1741,In_1937);
nand U205 (N_205,In_828,In_1596);
or U206 (N_206,In_2751,In_435);
and U207 (N_207,In_626,In_20);
xor U208 (N_208,In_1866,N_28);
nor U209 (N_209,In_134,In_504);
xor U210 (N_210,In_1995,N_107);
nor U211 (N_211,In_1498,In_2173);
nor U212 (N_212,In_2834,In_540);
nand U213 (N_213,In_625,In_1828);
nor U214 (N_214,In_2481,In_2060);
nor U215 (N_215,In_1992,In_1450);
nor U216 (N_216,In_317,In_992);
nand U217 (N_217,In_1730,In_1712);
and U218 (N_218,In_2471,In_2983);
and U219 (N_219,In_2655,In_156);
and U220 (N_220,In_1066,In_120);
nor U221 (N_221,In_2733,In_627);
xnor U222 (N_222,In_1492,In_1155);
nor U223 (N_223,In_150,N_154);
and U224 (N_224,In_923,In_184);
nor U225 (N_225,In_936,In_413);
or U226 (N_226,N_149,In_737);
nand U227 (N_227,In_2132,In_2648);
and U228 (N_228,In_82,In_1764);
or U229 (N_229,In_1925,In_1352);
nor U230 (N_230,In_1627,In_1439);
and U231 (N_231,In_644,In_1525);
nor U232 (N_232,In_1193,In_2357);
and U233 (N_233,In_138,In_2748);
and U234 (N_234,In_191,In_132);
or U235 (N_235,In_892,In_616);
nor U236 (N_236,In_1742,In_1434);
or U237 (N_237,In_1446,In_312);
nor U238 (N_238,In_2863,In_2731);
nor U239 (N_239,In_1538,In_1832);
and U240 (N_240,In_2877,In_2977);
or U241 (N_241,In_359,In_1261);
nor U242 (N_242,In_2193,In_2768);
or U243 (N_243,In_1005,In_903);
xnor U244 (N_244,In_2535,In_2015);
xor U245 (N_245,N_171,In_580);
or U246 (N_246,In_2846,In_1494);
or U247 (N_247,In_1720,In_1147);
and U248 (N_248,In_2532,In_1382);
and U249 (N_249,In_2227,In_1826);
or U250 (N_250,N_32,In_969);
xor U251 (N_251,In_6,N_131);
nand U252 (N_252,In_100,In_2822);
and U253 (N_253,N_76,In_2697);
and U254 (N_254,In_2732,In_195);
nand U255 (N_255,In_1870,N_40);
nand U256 (N_256,In_2479,In_1170);
and U257 (N_257,In_2463,In_1521);
and U258 (N_258,In_1673,In_238);
nor U259 (N_259,In_2641,In_58);
or U260 (N_260,In_1364,In_2128);
nor U261 (N_261,In_2192,In_2176);
nand U262 (N_262,In_2904,In_1951);
nor U263 (N_263,In_1347,In_1909);
xor U264 (N_264,In_985,In_1032);
and U265 (N_265,In_2148,N_122);
nand U266 (N_266,In_2703,In_1848);
nand U267 (N_267,In_333,In_2888);
xnor U268 (N_268,In_585,In_1641);
nor U269 (N_269,In_2013,In_2927);
or U270 (N_270,N_108,In_2107);
nor U271 (N_271,In_1428,In_1313);
and U272 (N_272,In_2108,In_365);
xor U273 (N_273,In_147,In_2401);
and U274 (N_274,In_133,N_80);
nor U275 (N_275,N_160,In_2313);
and U276 (N_276,In_1990,In_2283);
nor U277 (N_277,In_1954,N_86);
or U278 (N_278,In_1634,In_608);
or U279 (N_279,In_881,In_1356);
or U280 (N_280,In_1245,In_1199);
nand U281 (N_281,In_2739,N_69);
nor U282 (N_282,In_2050,In_1574);
xor U283 (N_283,In_2498,In_656);
xnor U284 (N_284,In_1955,In_1510);
or U285 (N_285,In_2682,In_2360);
nor U286 (N_286,In_2962,In_1542);
nand U287 (N_287,In_401,In_2347);
or U288 (N_288,In_1490,In_470);
xor U289 (N_289,In_1481,In_1761);
nand U290 (N_290,In_206,In_1570);
nor U291 (N_291,In_1996,In_2543);
xnor U292 (N_292,In_2854,In_8);
and U293 (N_293,In_930,In_2909);
nor U294 (N_294,In_2023,N_89);
nor U295 (N_295,In_1784,In_1134);
and U296 (N_296,In_808,In_2756);
or U297 (N_297,In_2698,In_925);
nand U298 (N_298,In_229,In_1650);
nand U299 (N_299,In_2469,In_1884);
nand U300 (N_300,N_10,In_2985);
nand U301 (N_301,In_671,In_2451);
xnor U302 (N_302,N_137,In_1786);
nor U303 (N_303,In_1781,In_2553);
or U304 (N_304,In_2508,In_371);
and U305 (N_305,In_2690,In_61);
nand U306 (N_306,In_12,In_2639);
nand U307 (N_307,In_2949,In_139);
nor U308 (N_308,In_2308,In_2079);
nand U309 (N_309,In_2821,In_2815);
or U310 (N_310,In_1306,In_619);
and U311 (N_311,In_825,In_5);
or U312 (N_312,In_1435,In_2850);
xnor U313 (N_313,In_649,In_1129);
xor U314 (N_314,In_1780,In_2519);
nand U315 (N_315,In_2914,In_2511);
or U316 (N_316,In_255,In_832);
nand U317 (N_317,In_81,N_133);
and U318 (N_318,In_1396,In_716);
nand U319 (N_319,In_1553,In_2129);
nor U320 (N_320,In_1961,In_1987);
nor U321 (N_321,N_175,In_2103);
or U322 (N_322,In_2951,In_98);
nand U323 (N_323,In_323,In_292);
nand U324 (N_324,In_104,In_121);
and U325 (N_325,In_2642,In_2395);
nand U326 (N_326,In_2191,In_980);
and U327 (N_327,In_1390,In_1709);
and U328 (N_328,In_376,N_61);
nor U329 (N_329,In_2879,In_2189);
nand U330 (N_330,In_2063,In_2970);
xnor U331 (N_331,In_979,In_2026);
nand U332 (N_332,In_2548,In_1509);
nor U333 (N_333,N_151,In_340);
and U334 (N_334,In_2225,In_2016);
or U335 (N_335,In_2634,In_1623);
and U336 (N_336,In_621,In_1002);
xnor U337 (N_337,In_1406,In_2209);
or U338 (N_338,In_1558,In_981);
and U339 (N_339,In_946,In_1209);
nand U340 (N_340,N_190,In_1279);
or U341 (N_341,In_2549,In_2204);
nand U342 (N_342,In_1447,In_886);
and U343 (N_343,N_121,In_44);
and U344 (N_344,In_2783,In_332);
and U345 (N_345,In_521,In_1403);
nand U346 (N_346,In_1467,In_1001);
nor U347 (N_347,In_1865,N_45);
xnor U348 (N_348,In_453,In_64);
nor U349 (N_349,In_763,In_1283);
and U350 (N_350,In_2485,In_99);
and U351 (N_351,In_1568,In_2538);
or U352 (N_352,In_2269,In_962);
nor U353 (N_353,In_1541,In_1617);
nand U354 (N_354,In_672,In_2932);
or U355 (N_355,In_183,In_714);
or U356 (N_356,N_172,N_170);
and U357 (N_357,In_2564,In_764);
xnor U358 (N_358,In_2187,In_198);
xor U359 (N_359,In_541,In_1020);
and U360 (N_360,In_90,In_1719);
xor U361 (N_361,In_1018,N_112);
and U362 (N_362,In_548,In_1707);
nor U363 (N_363,In_164,In_2370);
and U364 (N_364,In_2233,In_2435);
nor U365 (N_365,In_2002,In_2770);
and U366 (N_366,In_1915,N_187);
nor U367 (N_367,In_1704,In_460);
nor U368 (N_368,In_2105,In_2540);
nand U369 (N_369,In_577,N_81);
or U370 (N_370,In_1885,In_342);
nand U371 (N_371,In_1487,In_1873);
nand U372 (N_372,In_414,In_2483);
xnor U373 (N_373,N_35,In_938);
nor U374 (N_374,In_750,In_1246);
nand U375 (N_375,In_1640,In_1136);
nand U376 (N_376,In_898,In_27);
and U377 (N_377,In_2414,In_209);
and U378 (N_378,N_183,In_2907);
nor U379 (N_379,In_788,In_136);
and U380 (N_380,In_2386,In_1888);
nor U381 (N_381,In_1454,In_857);
and U382 (N_382,In_1105,In_2762);
or U383 (N_383,In_59,In_596);
xor U384 (N_384,In_1146,N_166);
xor U385 (N_385,In_445,In_1099);
or U386 (N_386,In_1289,In_295);
xnor U387 (N_387,In_1674,In_1263);
xor U388 (N_388,In_344,In_2873);
or U389 (N_389,In_126,In_2450);
and U390 (N_390,In_1247,In_953);
xor U391 (N_391,N_77,In_10);
nor U392 (N_392,In_814,In_1021);
xnor U393 (N_393,In_1632,In_637);
nor U394 (N_394,In_1973,In_2566);
nor U395 (N_395,In_171,In_2136);
or U396 (N_396,In_2750,In_226);
and U397 (N_397,In_112,In_829);
and U398 (N_398,In_2443,In_2102);
nand U399 (N_399,In_2504,In_2743);
or U400 (N_400,In_1302,In_657);
or U401 (N_401,In_1605,In_1204);
and U402 (N_402,In_1305,In_2430);
nand U403 (N_403,In_1676,In_720);
nand U404 (N_404,In_2164,In_2855);
or U405 (N_405,In_22,In_1891);
and U406 (N_406,In_382,In_2994);
and U407 (N_407,In_806,In_2707);
xnor U408 (N_408,In_1491,In_2059);
nor U409 (N_409,In_869,In_2074);
or U410 (N_410,N_164,N_99);
xnor U411 (N_411,In_1346,N_152);
and U412 (N_412,In_2206,In_2432);
nand U413 (N_413,In_1616,In_386);
xnor U414 (N_414,In_991,In_2721);
and U415 (N_415,In_2346,In_1329);
and U416 (N_416,In_787,N_337);
and U417 (N_417,In_1084,In_560);
and U418 (N_418,In_1940,In_2579);
nand U419 (N_419,In_2397,In_1197);
nand U420 (N_420,In_2941,In_1254);
nand U421 (N_421,In_710,N_49);
nor U422 (N_422,In_1095,In_1357);
or U423 (N_423,In_1592,In_668);
or U424 (N_424,In_1524,In_1694);
nand U425 (N_425,In_1791,In_2945);
xnor U426 (N_426,In_1762,N_341);
nand U427 (N_427,In_235,N_224);
and U428 (N_428,In_666,In_160);
nand U429 (N_429,In_579,In_847);
nor U430 (N_430,In_94,In_1180);
and U431 (N_431,In_1922,In_795);
nor U432 (N_432,In_1190,In_1772);
xor U433 (N_433,In_1090,In_1601);
xor U434 (N_434,In_535,In_286);
xnor U435 (N_435,In_931,In_73);
or U436 (N_436,In_1581,In_137);
xnor U437 (N_437,In_821,In_1648);
nor U438 (N_438,In_363,In_2279);
nand U439 (N_439,In_2024,In_963);
or U440 (N_440,In_2706,In_2668);
and U441 (N_441,In_1890,In_2650);
or U442 (N_442,In_1167,In_947);
nand U443 (N_443,In_2622,N_222);
or U444 (N_444,In_2693,In_2349);
and U445 (N_445,N_82,In_1595);
nor U446 (N_446,In_1716,In_747);
nand U447 (N_447,In_1503,In_2391);
and U448 (N_448,In_845,In_2229);
and U449 (N_449,In_1959,In_266);
xor U450 (N_450,In_145,In_2130);
nor U451 (N_451,In_635,In_636);
and U452 (N_452,In_1604,In_1980);
xnor U453 (N_453,In_904,In_509);
nor U454 (N_454,In_2286,In_320);
nand U455 (N_455,In_370,N_85);
xor U456 (N_456,In_1804,In_1964);
and U457 (N_457,In_2522,In_2048);
xor U458 (N_458,In_2900,In_987);
nor U459 (N_459,In_2487,In_2389);
nand U460 (N_460,In_395,In_536);
and U461 (N_461,N_394,In_2406);
and U462 (N_462,In_2222,N_390);
nand U463 (N_463,In_1326,In_2069);
xnor U464 (N_464,N_343,In_92);
nor U465 (N_465,N_130,In_114);
and U466 (N_466,In_2442,In_1098);
nand U467 (N_467,In_2929,In_83);
and U468 (N_468,In_1295,In_223);
nand U469 (N_469,In_813,In_2339);
nand U470 (N_470,In_419,In_2889);
nand U471 (N_471,In_2992,In_2777);
nor U472 (N_472,In_2413,In_1699);
nor U473 (N_473,In_1597,In_618);
xnor U474 (N_474,N_237,In_1006);
nor U475 (N_475,In_1117,In_2067);
nor U476 (N_476,In_935,In_2420);
nand U477 (N_477,N_321,In_1501);
nand U478 (N_478,In_2068,In_1917);
and U479 (N_479,In_1529,In_2312);
nand U480 (N_480,N_239,In_220);
nor U481 (N_481,In_2234,N_138);
nand U482 (N_482,In_253,In_858);
or U483 (N_483,In_1727,In_2012);
nor U484 (N_484,In_1244,In_1923);
xor U485 (N_485,In_2623,N_215);
nor U486 (N_486,N_225,In_833);
nand U487 (N_487,In_1875,N_391);
nand U488 (N_488,In_2144,In_1771);
nand U489 (N_489,In_35,In_2231);
nand U490 (N_490,In_2775,In_1478);
xor U491 (N_491,In_423,In_2021);
and U492 (N_492,N_105,In_2150);
and U493 (N_493,N_288,In_844);
xor U494 (N_494,In_2820,In_642);
and U495 (N_495,In_1578,In_1710);
nor U496 (N_496,In_2066,In_575);
xor U497 (N_497,N_74,N_377);
and U498 (N_498,In_1093,In_2651);
or U499 (N_499,In_875,In_2520);
nand U500 (N_500,In_2325,In_887);
nand U501 (N_501,In_268,N_189);
nor U502 (N_502,In_1270,In_70);
xnor U503 (N_503,In_1217,In_2628);
or U504 (N_504,In_1589,In_2986);
xnor U505 (N_505,In_231,In_1854);
nor U506 (N_506,In_1083,In_2790);
nor U507 (N_507,N_329,In_1825);
xnor U508 (N_508,In_19,In_2753);
nor U509 (N_509,In_1743,In_1754);
and U510 (N_510,In_213,In_1224);
and U511 (N_511,In_1539,In_2175);
nor U512 (N_512,In_2302,N_386);
or U513 (N_513,In_196,N_371);
xor U514 (N_514,In_274,In_1186);
nand U515 (N_515,In_2247,In_2257);
or U516 (N_516,In_920,In_1930);
xor U517 (N_517,In_2824,In_1842);
xor U518 (N_518,In_2112,In_96);
or U519 (N_519,In_1060,N_373);
and U520 (N_520,In_2094,In_1551);
nor U521 (N_521,In_170,In_494);
or U522 (N_522,N_290,In_2480);
and U523 (N_523,In_1255,In_1286);
or U524 (N_524,In_2186,In_1218);
or U525 (N_525,In_1474,In_911);
nand U526 (N_526,N_158,In_495);
nor U527 (N_527,In_1724,In_1091);
xnor U528 (N_528,In_2127,In_1534);
and U529 (N_529,In_1868,N_213);
or U530 (N_530,In_405,In_2747);
and U531 (N_531,In_2332,In_1324);
and U532 (N_532,N_258,N_142);
nor U533 (N_533,In_125,In_1839);
nor U534 (N_534,N_230,In_1896);
nor U535 (N_535,In_2263,In_1798);
nor U536 (N_536,N_381,In_385);
and U537 (N_537,In_2653,In_1577);
and U538 (N_538,In_1561,In_2273);
or U539 (N_539,In_1063,In_2677);
or U540 (N_540,In_477,N_278);
nand U541 (N_541,In_1172,In_2972);
nor U542 (N_542,N_54,In_1753);
nand U543 (N_543,In_1537,In_1252);
nand U544 (N_544,N_156,In_782);
nor U545 (N_545,In_1035,In_102);
nand U546 (N_546,In_2619,In_555);
and U547 (N_547,In_282,In_2604);
and U548 (N_548,In_21,In_2259);
or U549 (N_549,N_376,In_910);
nand U550 (N_550,In_161,In_2612);
and U551 (N_551,In_968,In_341);
nand U552 (N_552,In_2577,N_84);
xor U553 (N_553,In_1898,In_2807);
nand U554 (N_554,In_1608,N_51);
or U555 (N_555,In_970,In_1157);
nand U556 (N_556,In_853,In_2330);
nand U557 (N_557,In_38,In_1081);
nand U558 (N_558,In_1782,In_1097);
and U559 (N_559,In_392,In_2729);
xor U560 (N_560,In_2917,In_1046);
nor U561 (N_561,In_921,In_1100);
nand U562 (N_562,In_2194,In_928);
and U563 (N_563,In_257,In_882);
or U564 (N_564,In_2595,In_1410);
and U565 (N_565,In_1531,In_1835);
nor U566 (N_566,N_226,N_98);
or U567 (N_567,In_1877,In_2704);
xor U568 (N_568,N_362,In_1887);
xnor U569 (N_569,In_1746,In_742);
and U570 (N_570,In_1671,N_236);
xnor U571 (N_571,In_2230,In_2862);
xor U572 (N_572,In_1368,In_998);
nand U573 (N_573,In_2789,In_1455);
and U574 (N_574,In_820,In_544);
or U575 (N_575,In_1402,In_1291);
or U576 (N_576,N_393,In_1007);
xor U577 (N_577,In_2803,In_623);
or U578 (N_578,In_1030,In_1586);
nand U579 (N_579,In_2388,In_510);
xnor U580 (N_580,In_26,In_2800);
nor U581 (N_581,N_319,N_306);
and U582 (N_582,In_2852,In_2568);
nand U583 (N_583,In_75,In_1069);
and U584 (N_584,In_704,In_2780);
and U585 (N_585,In_1814,In_1281);
nor U586 (N_586,In_2984,In_1110);
nand U587 (N_587,In_762,In_1234);
nand U588 (N_588,In_1502,In_700);
nor U589 (N_589,In_2377,N_378);
or U590 (N_590,In_2018,In_2324);
nand U591 (N_591,In_2489,In_2291);
or U592 (N_592,In_590,N_359);
nand U593 (N_593,In_208,In_158);
xor U594 (N_594,In_2382,N_119);
and U595 (N_595,N_96,In_411);
or U596 (N_596,In_542,N_46);
nand U597 (N_597,In_162,In_1166);
and U598 (N_598,In_2901,In_403);
and U599 (N_599,In_1015,In_1335);
and U600 (N_600,In_557,In_352);
and U601 (N_601,In_664,In_1485);
nand U602 (N_602,In_1462,In_1836);
and U603 (N_603,In_217,In_432);
and U604 (N_604,In_1269,In_450);
xor U605 (N_605,In_528,In_2428);
and U606 (N_606,In_1944,In_1016);
nor U607 (N_607,In_2943,N_176);
xor U608 (N_608,In_95,N_566);
nand U609 (N_609,In_1082,N_558);
or U610 (N_610,In_426,N_368);
xnor U611 (N_611,In_1971,In_2817);
nand U612 (N_612,In_2064,In_289);
xor U613 (N_613,In_49,N_355);
xnor U614 (N_614,In_2124,N_211);
xnor U615 (N_615,In_1651,N_526);
nor U616 (N_616,In_1607,N_210);
nand U617 (N_617,In_1958,In_1941);
or U618 (N_618,N_214,In_1600);
xnor U619 (N_619,In_1074,N_395);
nand U620 (N_620,N_300,In_2341);
or U621 (N_621,In_2228,In_2336);
xor U622 (N_622,In_119,In_2052);
or U623 (N_623,In_1797,In_811);
xnor U624 (N_624,In_600,N_38);
and U625 (N_625,In_718,N_2);
and U626 (N_626,In_2866,In_1851);
and U627 (N_627,N_1,In_106);
xnor U628 (N_628,N_481,In_2499);
or U629 (N_629,N_455,In_959);
nand U630 (N_630,In_492,In_567);
xor U631 (N_631,In_93,In_2894);
nor U632 (N_632,In_1918,In_1052);
or U633 (N_633,In_2036,In_1036);
or U634 (N_634,In_630,In_2290);
nor U635 (N_635,In_2358,N_406);
nor U636 (N_636,In_574,In_23);
and U637 (N_637,In_246,In_942);
nand U638 (N_638,N_447,N_414);
nor U639 (N_639,N_97,In_2658);
or U640 (N_640,In_2088,In_2270);
or U641 (N_641,N_220,In_280);
nand U642 (N_642,In_784,In_254);
and U643 (N_643,In_1107,In_870);
or U644 (N_644,In_1794,In_2123);
and U645 (N_645,In_298,In_988);
xor U646 (N_646,In_2361,In_1750);
xnor U647 (N_647,In_1163,N_363);
or U648 (N_648,In_2292,N_413);
nor U649 (N_649,N_459,In_1696);
and U650 (N_650,In_2141,In_873);
xor U651 (N_651,N_298,In_899);
nor U652 (N_652,In_2384,In_1840);
xor U653 (N_653,In_1176,In_2849);
nor U654 (N_654,In_2971,In_2547);
nand U655 (N_655,In_2599,In_498);
nand U656 (N_656,In_2772,N_497);
xnor U657 (N_657,N_400,N_104);
nand U658 (N_658,In_1400,In_760);
or U659 (N_659,In_2404,In_678);
or U660 (N_660,In_669,In_1482);
or U661 (N_661,N_433,In_610);
xor U662 (N_662,In_1886,In_688);
xor U663 (N_663,In_1760,In_2416);
xnor U664 (N_664,In_2376,N_520);
or U665 (N_665,N_423,In_1375);
nor U666 (N_666,N_452,In_1841);
xor U667 (N_667,N_153,In_2567);
and U668 (N_668,N_13,In_2080);
nand U669 (N_669,In_1899,N_126);
nor U670 (N_670,In_2287,N_307);
nand U671 (N_671,In_905,N_150);
xnor U672 (N_672,N_246,In_2626);
nand U673 (N_673,N_93,In_1874);
nor U674 (N_674,In_2411,In_2178);
nand U675 (N_675,In_524,In_1834);
nor U676 (N_676,In_2296,N_280);
nor U677 (N_677,In_1609,In_324);
and U678 (N_678,In_1188,In_816);
nor U679 (N_679,In_1050,In_1732);
nand U680 (N_680,N_62,In_2348);
and U681 (N_681,In_1497,In_393);
xnor U682 (N_682,In_1969,In_2275);
and U683 (N_683,In_658,In_513);
or U684 (N_684,In_62,In_1666);
nor U685 (N_685,In_430,In_2843);
xnor U686 (N_686,N_598,In_2431);
or U687 (N_687,In_2198,In_178);
nand U688 (N_688,N_502,In_2670);
or U689 (N_689,In_2839,In_163);
and U690 (N_690,N_491,N_477);
nor U691 (N_691,In_803,In_2735);
xor U692 (N_692,In_2271,In_431);
nor U693 (N_693,In_2097,In_2326);
or U694 (N_694,In_2486,In_2990);
and U695 (N_695,In_2368,In_1034);
and U696 (N_696,In_2583,In_1790);
and U697 (N_697,In_1569,In_1830);
nand U698 (N_698,N_536,In_338);
nand U699 (N_699,In_202,In_2874);
nand U700 (N_700,In_1031,In_2197);
nand U701 (N_701,N_590,In_155);
nand U702 (N_702,In_2702,In_124);
xnor U703 (N_703,N_486,In_895);
nor U704 (N_704,N_510,N_471);
nand U705 (N_705,N_374,In_2322);
nor U706 (N_706,In_1697,In_919);
and U707 (N_707,In_1562,In_1587);
or U708 (N_708,N_299,In_2514);
or U709 (N_709,In_2205,In_1827);
xnor U710 (N_710,N_456,In_1307);
and U711 (N_711,In_2890,In_468);
or U712 (N_712,In_219,In_285);
nor U713 (N_713,In_1796,In_277);
nand U714 (N_714,In_1397,N_367);
nor U715 (N_715,In_2399,In_632);
xnor U716 (N_716,In_421,In_1309);
or U717 (N_717,N_469,N_454);
nand U718 (N_718,N_181,In_592);
nand U719 (N_719,In_2305,In_1300);
nor U720 (N_720,N_494,In_1976);
nand U721 (N_721,In_729,In_1064);
xnor U722 (N_722,N_268,N_532);
nor U723 (N_723,In_705,N_562);
nor U724 (N_724,N_462,In_1663);
or U725 (N_725,In_559,In_1010);
or U726 (N_726,In_2151,In_2667);
or U727 (N_727,In_726,In_2916);
or U728 (N_728,In_2076,In_194);
or U729 (N_729,N_188,N_241);
nand U730 (N_730,In_2875,In_176);
and U731 (N_731,In_1360,In_1242);
nand U732 (N_732,In_1618,In_2126);
nand U733 (N_733,N_488,In_1603);
nor U734 (N_734,N_569,In_2675);
or U735 (N_735,In_1230,N_223);
nor U736 (N_736,In_190,In_1652);
or U737 (N_737,In_2666,In_2806);
and U738 (N_738,In_2546,In_1041);
xor U739 (N_739,In_1221,In_538);
and U740 (N_740,In_2878,In_288);
nor U741 (N_741,N_506,In_1088);
xor U742 (N_742,In_2095,In_2551);
or U743 (N_743,In_1657,In_730);
and U744 (N_744,In_741,N_490);
nand U745 (N_745,In_2996,In_2022);
or U746 (N_746,N_397,In_2201);
nand U747 (N_747,In_2333,In_2084);
nand U748 (N_748,N_328,N_275);
and U749 (N_749,In_940,In_47);
or U750 (N_750,In_2115,In_1345);
and U751 (N_751,In_2284,In_2311);
xnor U752 (N_752,In_1418,In_712);
nand U753 (N_753,In_2967,In_400);
and U754 (N_754,N_52,In_594);
nand U755 (N_755,In_2881,In_2051);
and U756 (N_756,N_261,In_308);
nand U757 (N_757,In_169,N_479);
xor U758 (N_758,In_1148,In_515);
or U759 (N_759,In_1734,In_1544);
and U760 (N_760,In_1457,In_662);
nor U761 (N_761,In_493,N_578);
or U762 (N_762,In_755,In_751);
nand U763 (N_763,In_1009,In_1332);
nor U764 (N_764,In_1988,In_770);
nand U765 (N_765,N_372,N_492);
nor U766 (N_766,In_441,In_1548);
nand U767 (N_767,In_7,N_221);
or U768 (N_768,In_950,In_2003);
or U769 (N_769,In_1960,In_379);
and U770 (N_770,In_1144,In_1585);
nand U771 (N_771,In_2472,In_1154);
xnor U772 (N_772,N_266,In_838);
nand U773 (N_773,In_1999,N_267);
nor U774 (N_774,N_232,In_2343);
and U775 (N_775,N_272,In_2149);
or U776 (N_776,In_36,In_1268);
nor U777 (N_777,In_1094,In_651);
nand U778 (N_778,N_295,N_444);
nand U779 (N_779,In_539,In_2764);
or U780 (N_780,In_1017,In_1766);
xnor U781 (N_781,In_591,In_2449);
nand U782 (N_782,In_2691,In_1523);
nand U783 (N_783,In_248,In_1808);
nor U784 (N_784,N_14,In_2210);
and U785 (N_785,In_880,N_286);
or U786 (N_786,In_2705,In_1033);
or U787 (N_787,In_14,In_110);
and U788 (N_788,In_2801,N_449);
nor U789 (N_789,In_87,In_1752);
or U790 (N_790,In_1174,N_325);
or U791 (N_791,N_570,In_827);
xor U792 (N_792,In_2353,In_2264);
xnor U793 (N_793,In_2318,In_2953);
or U794 (N_794,N_336,In_2805);
nor U795 (N_795,In_335,In_1860);
or U796 (N_796,N_425,N_495);
and U797 (N_797,In_260,In_449);
or U798 (N_798,In_624,N_442);
nor U799 (N_799,N_583,In_1311);
or U800 (N_800,In_390,In_849);
and U801 (N_801,In_679,In_633);
or U802 (N_802,In_554,In_655);
and U803 (N_803,In_529,In_2905);
nand U804 (N_804,N_587,In_1071);
or U805 (N_805,In_1532,In_1547);
or U806 (N_806,In_576,In_1970);
and U807 (N_807,In_719,In_917);
and U808 (N_808,In_2260,N_7);
or U809 (N_809,In_2620,In_2465);
nor U810 (N_810,In_1594,In_2464);
or U811 (N_811,N_327,N_797);
or U812 (N_812,In_406,In_1806);
nand U813 (N_813,N_549,In_1075);
nand U814 (N_814,N_110,In_2070);
or U815 (N_815,N_707,In_1106);
nand U816 (N_816,In_2219,In_1845);
xor U817 (N_817,In_699,N_301);
xor U818 (N_818,In_1143,In_2689);
nand U819 (N_819,In_1092,In_2767);
xnor U820 (N_820,In_2028,In_76);
nor U821 (N_821,N_780,In_1862);
nand U822 (N_822,N_173,In_2507);
or U823 (N_823,In_350,In_2829);
nor U824 (N_824,In_739,In_1659);
and U825 (N_825,In_2329,N_117);
nand U826 (N_826,N_408,In_2309);
and U827 (N_827,In_1200,In_399);
nand U828 (N_828,In_1872,In_1384);
and U829 (N_829,N_339,In_2584);
xnor U830 (N_830,N_678,N_585);
or U831 (N_831,N_745,In_1864);
xor U832 (N_832,N_658,N_749);
and U833 (N_833,In_2091,In_2183);
and U834 (N_834,In_2744,In_2870);
nor U835 (N_835,N_627,N_572);
and U836 (N_836,In_893,In_2804);
xor U837 (N_837,In_2299,N_205);
xnor U838 (N_838,In_1802,In_1401);
xnor U839 (N_839,In_2638,In_1807);
nor U840 (N_840,N_795,N_23);
and U841 (N_841,In_1453,N_466);
or U842 (N_842,In_1297,In_2093);
xnor U843 (N_843,In_1763,In_1850);
and U844 (N_844,N_784,In_2495);
or U845 (N_845,In_1177,In_1636);
nor U846 (N_846,N_238,In_1054);
nor U847 (N_847,In_1486,In_2160);
nand U848 (N_848,In_501,N_405);
nor U849 (N_849,N_270,N_522);
or U850 (N_850,In_1365,In_1929);
xor U851 (N_851,N_385,In_823);
nor U852 (N_852,In_1892,N_602);
and U853 (N_853,In_2552,In_802);
xor U854 (N_854,N_513,In_1876);
or U855 (N_855,In_1111,In_2392);
nor U856 (N_856,In_1737,In_232);
and U857 (N_857,N_448,In_891);
xnor U858 (N_858,N_686,N_392);
or U859 (N_859,N_732,In_1630);
or U860 (N_860,In_614,In_306);
nor U861 (N_861,In_514,In_573);
nand U862 (N_862,In_182,In_550);
xor U863 (N_863,In_2533,N_198);
or U864 (N_864,In_1298,In_2637);
or U865 (N_865,In_2029,N_437);
and U866 (N_866,N_231,In_1068);
nand U867 (N_867,In_2454,In_2043);
nor U868 (N_868,In_1910,In_1140);
or U869 (N_869,N_264,In_329);
xor U870 (N_870,In_2365,In_88);
nor U871 (N_871,N_793,In_28);
nor U872 (N_872,In_305,In_1319);
and U873 (N_873,In_1989,In_429);
xnor U874 (N_874,In_723,In_2586);
and U875 (N_875,In_2891,In_1282);
or U876 (N_876,In_914,In_2425);
and U877 (N_877,In_1499,In_1735);
and U878 (N_878,In_2618,N_102);
xnor U879 (N_879,N_663,N_725);
or U880 (N_880,N_281,N_694);
and U881 (N_881,In_1612,N_677);
xnor U882 (N_882,N_312,N_623);
or U883 (N_883,In_1358,N_434);
or U884 (N_884,N_601,In_906);
or U885 (N_885,In_2937,N_560);
nor U886 (N_886,In_2172,In_30);
nor U887 (N_887,In_1258,In_2473);
xor U888 (N_888,In_2738,In_291);
nand U889 (N_889,N_634,In_2837);
nand U890 (N_890,N_698,In_264);
xnor U891 (N_891,In_1275,In_2117);
or U892 (N_892,In_638,In_2371);
nor U893 (N_893,In_215,In_945);
nor U894 (N_894,N_750,In_2903);
and U895 (N_895,In_2763,N_755);
xnor U896 (N_896,In_1028,In_2948);
or U897 (N_897,In_2122,In_934);
nor U898 (N_898,In_2625,N_421);
nand U899 (N_899,In_2537,N_689);
nor U900 (N_900,In_1775,In_2988);
and U901 (N_901,N_418,In_2440);
or U902 (N_902,In_1386,N_33);
xor U903 (N_903,In_1731,N_555);
or U904 (N_904,N_88,In_1952);
nor U905 (N_905,In_2403,In_2113);
nand U906 (N_906,In_367,In_2935);
nand U907 (N_907,In_1123,In_503);
and U908 (N_908,In_1328,N_727);
xnor U909 (N_909,In_563,N_661);
nand U910 (N_910,In_1104,N_672);
nor U911 (N_911,In_915,In_300);
or U912 (N_912,In_165,N_726);
xor U913 (N_913,In_135,N_310);
xnor U914 (N_914,In_851,In_446);
nor U915 (N_915,In_2657,In_1011);
nor U916 (N_916,In_2369,In_2912);
and U917 (N_917,N_687,In_63);
nand U918 (N_918,In_2965,N_674);
or U919 (N_919,N_599,N_42);
xnor U920 (N_920,In_2717,N_713);
or U921 (N_921,N_617,In_1185);
and U922 (N_922,N_527,N_507);
and U923 (N_923,In_686,In_1248);
xor U924 (N_924,In_2647,In_212);
xnor U925 (N_925,In_653,In_1451);
and U926 (N_926,In_771,N_139);
nand U927 (N_927,N_467,In_427);
and U928 (N_928,In_113,N_417);
nand U929 (N_929,In_2501,In_2856);
or U930 (N_930,In_313,In_863);
and U931 (N_931,N_465,In_1669);
nor U932 (N_932,In_868,In_1550);
and U933 (N_933,N_641,N_616);
nor U934 (N_934,In_2892,In_2282);
or U935 (N_935,In_1615,In_2448);
and U936 (N_936,N_269,N_387);
and U937 (N_937,In_1495,In_1983);
nand U938 (N_938,N_333,In_2736);
xor U939 (N_939,N_650,N_657);
xnor U940 (N_940,N_608,N_409);
nor U941 (N_941,N_388,In_1087);
or U942 (N_942,In_1264,In_722);
xnor U943 (N_943,N_690,N_518);
and U944 (N_944,N_684,In_1423);
nand U945 (N_945,N_542,N_739);
nand U946 (N_946,In_628,In_327);
nor U947 (N_947,In_2256,In_2086);
and U948 (N_948,In_807,In_2455);
nand U949 (N_949,N_157,In_556);
nand U950 (N_950,In_1795,In_2303);
nor U951 (N_951,N_799,N_370);
nor U952 (N_952,In_1202,In_1935);
or U953 (N_953,N_733,In_1235);
xor U954 (N_954,In_2861,N_401);
or U955 (N_955,N_59,N_411);
and U956 (N_956,In_799,N_769);
xnor U957 (N_957,N_655,N_625);
nor U958 (N_958,In_2165,In_2644);
nor U959 (N_959,N_200,N_375);
nand U960 (N_960,In_346,N_124);
nor U961 (N_961,In_186,In_1408);
xor U962 (N_962,In_568,In_91);
nor U963 (N_963,In_2407,N_197);
or U964 (N_964,In_1048,N_426);
and U965 (N_965,N_283,In_1181);
nand U966 (N_966,In_275,In_885);
nand U967 (N_967,In_2799,N_571);
nand U968 (N_968,N_314,N_346);
or U969 (N_969,In_1978,In_1670);
nor U970 (N_970,In_2047,In_2938);
xnor U971 (N_971,In_2627,In_775);
xnor U972 (N_972,In_2243,N_646);
or U973 (N_973,In_566,In_2700);
nand U974 (N_974,In_484,N_36);
nor U975 (N_975,In_2643,In_2600);
nor U976 (N_976,In_2997,In_791);
xor U977 (N_977,In_1349,In_204);
or U978 (N_978,In_1506,In_1304);
or U979 (N_979,In_1567,In_546);
and U980 (N_980,In_2885,In_108);
nor U981 (N_981,N_619,N_746);
nand U982 (N_982,N_340,N_552);
nand U983 (N_983,In_278,N_609);
nor U984 (N_984,In_2062,In_1685);
nand U985 (N_985,In_663,N_747);
nand U986 (N_986,In_2474,N_292);
xnor U987 (N_987,N_489,In_2119);
nor U988 (N_988,In_673,In_523);
and U989 (N_989,In_1660,In_2409);
nor U990 (N_990,N_643,In_2235);
nor U991 (N_991,In_1675,In_2939);
or U992 (N_992,In_734,In_307);
nand U993 (N_993,In_1938,N_64);
nor U994 (N_994,N_316,In_174);
or U995 (N_995,In_1799,In_2350);
nor U996 (N_996,In_2190,N_415);
or U997 (N_997,In_475,In_442);
nand U998 (N_998,In_2926,In_2004);
nand U999 (N_999,N_547,N_612);
or U1000 (N_1000,In_1626,N_699);
nor U1001 (N_1001,In_418,N_953);
nand U1002 (N_1002,In_1686,N_344);
nor U1003 (N_1003,N_419,In_417);
nor U1004 (N_1004,In_2588,N_39);
nor U1005 (N_1005,In_1132,In_1765);
and U1006 (N_1006,N_703,N_25);
or U1007 (N_1007,In_2826,In_1703);
xnor U1008 (N_1008,N_63,N_174);
or U1009 (N_1009,In_1527,In_297);
or U1010 (N_1010,In_2559,In_1511);
and U1011 (N_1011,In_1273,In_2152);
xnor U1012 (N_1012,In_2512,In_2950);
or U1013 (N_1013,In_1713,N_729);
xnor U1014 (N_1014,N_353,In_1774);
and U1015 (N_1015,In_2629,N_568);
xor U1016 (N_1016,N_987,In_16);
xnor U1017 (N_1017,In_1377,In_1284);
xnor U1018 (N_1018,In_451,N_66);
nor U1019 (N_1019,N_994,N_185);
nor U1020 (N_1020,In_2802,In_1262);
and U1021 (N_1021,N_865,In_2297);
xor U1022 (N_1022,In_2071,In_776);
xnor U1023 (N_1023,In_2575,N_659);
xor U1024 (N_1024,N_323,In_2969);
nor U1025 (N_1025,N_380,In_1993);
xnor U1026 (N_1026,In_1668,In_37);
and U1027 (N_1027,In_2142,N_229);
and U1028 (N_1028,In_1936,N_811);
nand U1029 (N_1029,In_533,In_258);
and U1030 (N_1030,In_835,In_1477);
nor U1031 (N_1031,In_2277,In_2771);
nand U1032 (N_1032,In_1749,N_186);
or U1033 (N_1033,In_2617,N_863);
or U1034 (N_1034,In_864,In_1624);
and U1035 (N_1035,In_2944,In_129);
and U1036 (N_1036,In_1003,In_2010);
nand U1037 (N_1037,In_505,In_681);
xnor U1038 (N_1038,In_639,In_374);
and U1039 (N_1039,N_106,In_1067);
nor U1040 (N_1040,In_2372,In_818);
and U1041 (N_1041,In_2328,N_441);
xor U1042 (N_1042,In_2591,In_1829);
or U1043 (N_1043,In_127,In_2058);
and U1044 (N_1044,N_265,In_489);
and U1045 (N_1045,In_2285,In_2724);
nand U1046 (N_1046,In_227,In_2075);
nor U1047 (N_1047,In_1057,In_1409);
nor U1048 (N_1048,In_1729,In_547);
xnor U1049 (N_1049,In_2838,N_790);
nand U1050 (N_1050,In_2467,N_782);
and U1051 (N_1051,N_600,In_1639);
and U1052 (N_1052,In_2936,N_744);
nand U1053 (N_1053,N_4,In_2687);
nand U1054 (N_1054,In_774,In_1682);
and U1055 (N_1055,N_574,In_1469);
xnor U1056 (N_1056,In_620,In_2422);
or U1057 (N_1057,In_2232,N_924);
xnor U1058 (N_1058,In_481,N_350);
xnor U1059 (N_1059,N_951,In_1449);
xnor U1060 (N_1060,N_928,In_1723);
nand U1061 (N_1061,In_2734,N_514);
nand U1062 (N_1062,N_767,N_629);
nor U1063 (N_1063,In_2827,In_466);
nor U1064 (N_1064,N_358,N_890);
nor U1065 (N_1065,In_708,In_2510);
xnor U1066 (N_1066,In_434,In_116);
xnor U1067 (N_1067,N_632,N_279);
xnor U1068 (N_1068,N_664,N_884);
nor U1069 (N_1069,N_543,In_1153);
nor U1070 (N_1070,N_55,N_311);
or U1071 (N_1071,N_438,In_2886);
nor U1072 (N_1072,N_516,N_958);
and U1073 (N_1073,In_1912,In_1359);
xor U1074 (N_1074,In_34,In_1475);
xnor U1075 (N_1075,N_412,In_2931);
nor U1076 (N_1076,In_290,In_759);
nand U1077 (N_1077,In_2223,N_313);
and U1078 (N_1078,In_2452,N_206);
and U1079 (N_1079,N_883,In_2202);
nand U1080 (N_1080,In_1809,In_1778);
xnor U1081 (N_1081,In_2578,N_476);
xnor U1082 (N_1082,In_1927,N_194);
nand U1083 (N_1083,N_16,N_90);
or U1084 (N_1084,N_906,In_1014);
and U1085 (N_1085,N_683,In_1505);
nor U1086 (N_1086,In_564,In_2111);
nand U1087 (N_1087,N_140,In_1376);
nor U1088 (N_1088,In_680,In_1272);
nor U1089 (N_1089,In_488,In_303);
or U1090 (N_1090,In_2761,In_394);
nor U1091 (N_1091,N_702,In_39);
and U1092 (N_1092,In_2718,In_151);
nand U1093 (N_1093,N_253,In_522);
nand U1094 (N_1094,N_79,In_2692);
nand U1095 (N_1095,In_587,In_1483);
xor U1096 (N_1096,In_843,In_2301);
nor U1097 (N_1097,N_503,N_512);
nor U1098 (N_1098,In_1314,In_850);
xor U1099 (N_1099,N_866,In_1043);
and U1100 (N_1100,In_749,In_561);
or U1101 (N_1101,In_752,N_956);
or U1102 (N_1102,N_293,N_669);
nand U1103 (N_1103,In_2134,In_996);
xnor U1104 (N_1104,N_691,N_615);
nor U1105 (N_1105,In_2602,In_2427);
or U1106 (N_1106,In_1692,In_131);
xor U1107 (N_1107,In_965,In_2468);
xor U1108 (N_1108,N_875,N_606);
nor U1109 (N_1109,In_2252,In_2766);
nand U1110 (N_1110,N_996,In_1931);
xnor U1111 (N_1111,In_676,In_1693);
nand U1112 (N_1112,In_461,In_4);
nor U1113 (N_1113,N_805,In_1285);
or U1114 (N_1114,N_348,N_652);
xor U1115 (N_1115,In_244,N_837);
and U1116 (N_1116,N_15,In_756);
and U1117 (N_1117,In_2554,In_1363);
or U1118 (N_1118,N_808,N_777);
and U1119 (N_1119,N_649,In_983);
xor U1120 (N_1120,In_1967,In_2723);
or U1121 (N_1121,In_293,In_168);
and U1122 (N_1122,In_364,In_490);
or U1123 (N_1123,N_17,In_2217);
nand U1124 (N_1124,In_80,N_891);
and U1125 (N_1125,In_2118,N_993);
and U1126 (N_1126,In_2327,N_428);
xor U1127 (N_1127,In_1792,In_347);
nand U1128 (N_1128,In_1654,In_2842);
nand U1129 (N_1129,N_640,In_1522);
nand U1130 (N_1130,N_87,In_2825);
nand U1131 (N_1131,In_859,N_132);
nor U1132 (N_1132,In_1751,In_2500);
nor U1133 (N_1133,In_2933,N_792);
or U1134 (N_1134,N_320,In_2238);
nand U1135 (N_1135,In_1757,N_988);
and U1136 (N_1136,In_1205,In_971);
nor U1137 (N_1137,In_1556,In_2773);
xor U1138 (N_1138,In_465,In_2462);
xnor U1139 (N_1139,N_435,In_792);
or U1140 (N_1140,In_884,In_758);
and U1141 (N_1141,N_909,In_2792);
xor U1142 (N_1142,In_433,In_1901);
and U1143 (N_1143,In_1801,In_797);
xor U1144 (N_1144,N_475,In_1956);
or U1145 (N_1145,N_895,In_1897);
nor U1146 (N_1146,In_2596,In_2364);
nand U1147 (N_1147,In_471,N_973);
nor U1148 (N_1148,N_18,In_1464);
and U1149 (N_1149,N_159,In_862);
nor U1150 (N_1150,In_396,In_2366);
and U1151 (N_1151,N_743,In_1565);
nor U1152 (N_1152,N_303,In_2402);
and U1153 (N_1153,N_410,In_222);
or U1154 (N_1154,In_51,N_851);
or U1155 (N_1155,In_572,In_1251);
nand U1156 (N_1156,N_929,In_326);
or U1157 (N_1157,N_450,In_2593);
nor U1158 (N_1158,In_262,In_2244);
nand U1159 (N_1159,In_2847,N_27);
xor U1160 (N_1160,In_301,In_1591);
nor U1161 (N_1161,N_111,In_2317);
and U1162 (N_1162,In_2211,In_1114);
xnor U1163 (N_1163,N_219,In_2461);
or U1164 (N_1164,In_2570,In_631);
and U1165 (N_1165,In_1226,In_2758);
nand U1166 (N_1166,N_484,In_997);
and U1167 (N_1167,N_227,In_2030);
or U1168 (N_1168,In_1745,N_881);
nor U1169 (N_1169,In_439,In_185);
xnor U1170 (N_1170,In_2226,In_706);
xor U1171 (N_1171,In_1690,In_1902);
or U1172 (N_1172,In_463,In_2518);
nand U1173 (N_1173,In_54,In_1045);
nor U1174 (N_1174,In_2814,In_1385);
or U1175 (N_1175,In_796,In_2338);
nand U1176 (N_1176,In_944,In_296);
nor U1177 (N_1177,In_497,In_1257);
or U1178 (N_1178,In_777,In_1212);
and U1179 (N_1179,N_668,In_1445);
or U1180 (N_1180,In_1427,N_907);
or U1181 (N_1181,N_334,In_1416);
or U1182 (N_1182,N_908,In_1112);
and U1183 (N_1183,In_302,In_1833);
xnor U1184 (N_1184,In_1500,N_550);
and U1185 (N_1185,In_948,In_1432);
and U1186 (N_1186,In_2872,In_1086);
xnor U1187 (N_1187,In_867,N_975);
nor U1188 (N_1188,In_2565,In_1655);
or U1189 (N_1189,In_1137,N_915);
nor U1190 (N_1190,In_2711,In_2035);
nand U1191 (N_1191,In_926,In_2524);
nor U1192 (N_1192,In_1882,In_687);
and U1193 (N_1193,In_2081,In_299);
xor U1194 (N_1194,In_1638,In_1916);
xor U1195 (N_1195,N_468,In_1290);
nand U1196 (N_1196,In_17,In_696);
nand U1197 (N_1197,In_502,In_2818);
xor U1198 (N_1198,N_700,N_719);
nor U1199 (N_1199,N_342,In_534);
nand U1200 (N_1200,In_1012,N_1112);
nor U1201 (N_1201,In_378,In_1271);
nand U1202 (N_1202,N_919,In_2181);
or U1203 (N_1203,N_1036,N_354);
or U1204 (N_1204,N_1026,N_1042);
xnor U1205 (N_1205,N_1065,In_2754);
xnor U1206 (N_1206,N_825,N_259);
nand U1207 (N_1207,N_758,In_866);
nor U1208 (N_1208,N_129,In_2694);
and U1209 (N_1209,In_2444,In_271);
nor U1210 (N_1210,In_2521,In_976);
xor U1211 (N_1211,In_1062,In_1299);
and U1212 (N_1212,N_1148,N_3);
xor U1213 (N_1213,In_2673,N_815);
and U1214 (N_1214,In_1726,N_534);
nand U1215 (N_1215,N_636,N_116);
xnor U1216 (N_1216,In_2876,N_8);
nand U1217 (N_1217,N_927,N_685);
and U1218 (N_1218,In_2830,In_2794);
nand U1219 (N_1219,In_2509,In_733);
and U1220 (N_1220,N_667,N_19);
xnor U1221 (N_1221,N_1108,In_677);
nand U1222 (N_1222,In_2321,N_240);
nand U1223 (N_1223,N_717,In_984);
or U1224 (N_1224,N_939,In_2746);
and U1225 (N_1225,In_115,In_1077);
or U1226 (N_1226,In_1543,N_1002);
and U1227 (N_1227,N_695,In_420);
xnor U1228 (N_1228,In_467,In_1430);
nand U1229 (N_1229,N_384,In_1040);
nand U1230 (N_1230,N_114,In_1219);
xor U1231 (N_1231,In_2529,N_1005);
nand U1232 (N_1232,In_2180,N_844);
or U1233 (N_1233,In_929,N_666);
xnor U1234 (N_1234,In_1096,N_1160);
nor U1235 (N_1235,In_2608,In_516);
and U1236 (N_1236,In_2214,In_1142);
nand U1237 (N_1237,N_810,N_1139);
and U1238 (N_1238,In_2660,In_2374);
nand U1239 (N_1239,N_846,N_976);
or U1240 (N_1240,N_485,In_593);
and U1241 (N_1241,N_56,In_1816);
nand U1242 (N_1242,In_1343,In_1239);
or U1243 (N_1243,In_2337,In_1008);
or U1244 (N_1244,N_1028,In_1755);
or U1245 (N_1245,In_1162,In_181);
xnor U1246 (N_1246,In_549,In_689);
and U1247 (N_1247,In_2719,N_365);
xnor U1248 (N_1248,In_2961,N_1132);
nor U1249 (N_1249,N_499,In_1563);
xor U1250 (N_1250,N_308,N_1144);
xnor U1251 (N_1251,N_1124,N_622);
nor U1252 (N_1252,In_2956,N_193);
or U1253 (N_1253,N_778,In_443);
or U1254 (N_1254,In_1822,In_2560);
nand U1255 (N_1255,N_1089,N_294);
or U1256 (N_1256,In_1687,In_357);
xor U1257 (N_1257,In_2614,In_1740);
or U1258 (N_1258,In_2359,In_2381);
nor U1259 (N_1259,In_172,N_1187);
nor U1260 (N_1260,N_260,N_1169);
nand U1261 (N_1261,N_1136,N_830);
nand U1262 (N_1262,In_11,In_2942);
xnor U1263 (N_1263,N_981,N_912);
and U1264 (N_1264,In_1287,N_788);
nor U1265 (N_1265,N_624,N_1156);
and U1266 (N_1266,In_2161,In_2610);
xnor U1267 (N_1267,In_1846,N_285);
xor U1268 (N_1268,N_538,In_2470);
nand U1269 (N_1269,N_24,In_2884);
nor U1270 (N_1270,In_531,N_937);
nand U1271 (N_1271,N_880,N_839);
nor U1272 (N_1272,In_1436,In_1869);
and U1273 (N_1273,N_984,In_1805);
xnor U1274 (N_1274,N_347,N_806);
and U1275 (N_1275,In_1744,In_2298);
xor U1276 (N_1276,N_586,In_496);
and U1277 (N_1277,In_46,In_2253);
nand U1278 (N_1278,In_2220,In_856);
or U1279 (N_1279,In_1488,In_2616);
or U1280 (N_1280,N_822,N_943);
nor U1281 (N_1281,N_20,N_244);
xor U1282 (N_1282,In_1471,In_2157);
or U1283 (N_1283,In_456,N_710);
nor U1284 (N_1284,In_2715,In_2680);
xor U1285 (N_1285,N_179,In_2613);
nor U1286 (N_1286,In_197,In_2237);
xor U1287 (N_1287,In_2550,N_605);
nor U1288 (N_1288,In_1844,In_960);
nand U1289 (N_1289,In_2921,N_796);
nand U1290 (N_1290,N_1185,In_1208);
and U1291 (N_1291,N_756,N_948);
nand U1292 (N_1292,In_525,N_487);
nand U1293 (N_1293,In_2250,N_934);
or U1294 (N_1294,N_842,In_2589);
xor U1295 (N_1295,N_961,N_263);
nor U1296 (N_1296,In_328,N_559);
xor U1297 (N_1297,In_2791,In_1629);
and U1298 (N_1298,N_835,N_818);
or U1299 (N_1299,N_1107,N_402);
or U1300 (N_1300,N_73,In_1926);
and U1301 (N_1301,In_912,N_823);
nor U1302 (N_1302,In_1216,N_761);
nand U1303 (N_1303,In_78,In_1220);
and U1304 (N_1304,In_1187,In_1672);
and U1305 (N_1305,In_2785,N_141);
xor U1306 (N_1306,In_1398,N_1093);
and U1307 (N_1307,N_470,In_402);
and U1308 (N_1308,In_2251,N_977);
and U1309 (N_1309,In_2200,N_618);
and U1310 (N_1310,In_424,N_742);
or U1311 (N_1311,N_436,In_1380);
nor U1312 (N_1312,N_1013,In_1429);
nor U1313 (N_1313,N_774,In_2278);
nand U1314 (N_1314,N_47,In_2424);
or U1315 (N_1315,In_2446,In_512);
nor U1316 (N_1316,In_1055,In_179);
and U1317 (N_1317,In_1213,N_965);
nor U1318 (N_1318,In_2809,In_1907);
nor U1319 (N_1319,In_65,In_242);
nand U1320 (N_1320,In_2061,In_1572);
nand U1321 (N_1321,N_809,In_2784);
xnor U1322 (N_1322,In_1546,N_949);
nand U1323 (N_1323,N_296,In_2954);
nand U1324 (N_1324,N_715,N_262);
or U1325 (N_1325,N_271,In_2168);
xor U1326 (N_1326,In_368,N_1033);
nor U1327 (N_1327,N_829,N_581);
xnor U1328 (N_1328,In_1924,N_1130);
nand U1329 (N_1329,N_803,In_785);
xnor U1330 (N_1330,In_2573,In_2998);
xnor U1331 (N_1331,N_1015,In_652);
nand U1332 (N_1332,In_2236,In_2494);
and U1333 (N_1333,In_2421,N_832);
and U1334 (N_1334,In_2354,N_53);
nor U1335 (N_1335,In_2590,In_218);
nand U1336 (N_1336,N_134,In_1369);
xnor U1337 (N_1337,N_445,N_1085);
xor U1338 (N_1338,In_261,N_680);
nand U1339 (N_1339,In_939,In_1150);
and U1340 (N_1340,N_1091,In_1557);
nand U1341 (N_1341,N_802,In_2923);
nand U1342 (N_1342,In_1715,In_1863);
nor U1343 (N_1343,In_1711,N_123);
xnor U1344 (N_1344,In_1070,N_653);
or U1345 (N_1345,N_840,N_1053);
and U1346 (N_1346,N_827,In_1820);
nor U1347 (N_1347,In_311,In_2979);
nand U1348 (N_1348,N_1014,N_850);
nor U1349 (N_1349,In_2858,In_1856);
or U1350 (N_1350,In_1189,In_1770);
nand U1351 (N_1351,In_526,N_1104);
nor U1352 (N_1352,In_1207,N_986);
nor U1353 (N_1353,In_366,In_2515);
or U1354 (N_1354,In_141,In_1517);
or U1355 (N_1355,In_1019,In_1120);
or U1356 (N_1356,In_1047,N_708);
and U1357 (N_1357,In_2090,In_2633);
nand U1358 (N_1358,In_570,In_1512);
nand U1359 (N_1359,In_1461,In_745);
xnor U1360 (N_1360,N_531,In_361);
nand U1361 (N_1361,In_1677,N_736);
nand U1362 (N_1362,In_1991,In_674);
or U1363 (N_1363,In_1688,N_276);
xor U1364 (N_1364,In_2006,N_633);
xor U1365 (N_1365,In_2466,N_431);
and U1366 (N_1366,In_50,In_744);
or U1367 (N_1367,In_175,In_1545);
xnor U1368 (N_1368,In_1420,In_1934);
nand U1369 (N_1369,In_2757,In_545);
and U1370 (N_1370,In_1437,N_1020);
and U1371 (N_1371,In_552,N_1197);
and U1372 (N_1372,N_548,In_571);
nand U1373 (N_1373,N_1078,N_1055);
nand U1374 (N_1374,In_732,In_1858);
and U1375 (N_1375,In_1393,N_1068);
xor U1376 (N_1376,In_2833,N_234);
or U1377 (N_1377,In_1135,In_837);
nor U1378 (N_1378,In_1022,In_2539);
nand U1379 (N_1379,In_1238,N_305);
nor U1380 (N_1380,In_812,N_1047);
nand U1381 (N_1381,N_1058,In_757);
or U1382 (N_1382,In_1076,In_2089);
or U1383 (N_1383,N_955,N_58);
xor U1384 (N_1384,In_315,N_1022);
nor U1385 (N_1385,N_75,N_1097);
nor U1386 (N_1386,In_754,In_2968);
or U1387 (N_1387,N_1048,N_383);
or U1388 (N_1388,N_974,N_1083);
xor U1389 (N_1389,N_789,In_1785);
nor U1390 (N_1390,N_541,In_2482);
nand U1391 (N_1391,In_1101,In_725);
nand U1392 (N_1392,N_770,In_1519);
nand U1393 (N_1393,In_2304,In_1861);
nor U1394 (N_1394,In_2053,N_501);
xor U1395 (N_1395,N_662,N_523);
nor U1396 (N_1396,In_166,In_360);
xnor U1397 (N_1397,In_975,In_3);
nor U1398 (N_1398,N_998,In_900);
nor U1399 (N_1399,N_1072,In_2828);
nand U1400 (N_1400,N_856,N_1358);
or U1401 (N_1401,N_162,In_1109);
nand U1402 (N_1402,In_2055,N_1149);
nand U1403 (N_1403,In_31,In_840);
or U1404 (N_1404,In_650,In_1387);
or U1405 (N_1405,N_1277,In_622);
nor U1406 (N_1406,In_1373,N_216);
or U1407 (N_1407,N_1098,N_1001);
and U1408 (N_1408,In_2663,N_473);
nand U1409 (N_1409,N_968,N_779);
and U1410 (N_1410,N_1182,In_2158);
xnor U1411 (N_1411,In_1237,In_901);
and U1412 (N_1412,N_1246,N_1090);
xnor U1413 (N_1413,N_1252,In_1479);
nand U1414 (N_1414,In_245,N_1087);
or U1415 (N_1415,N_1228,N_184);
nand U1416 (N_1416,In_187,In_167);
xor U1417 (N_1417,N_233,In_2207);
nor U1418 (N_1418,In_1000,N_1269);
or U1419 (N_1419,In_1184,In_1355);
xnor U1420 (N_1420,N_921,In_2536);
and U1421 (N_1421,In_1378,In_74);
nor U1422 (N_1422,In_40,In_1644);
or U1423 (N_1423,In_2632,N_1267);
nor U1424 (N_1424,In_584,N_1140);
or U1425 (N_1425,In_2265,N_1273);
and U1426 (N_1426,In_2417,N_287);
nand U1427 (N_1427,N_1339,N_1045);
xnor U1428 (N_1428,N_349,N_1129);
nand U1429 (N_1429,In_2716,N_1334);
xnor U1430 (N_1430,N_995,N_1133);
xnor U1431 (N_1431,N_714,In_1441);
or U1432 (N_1432,N_1007,In_2506);
or U1433 (N_1433,N_1227,N_1365);
nand U1434 (N_1434,In_1582,N_693);
and U1435 (N_1435,N_277,N_1120);
or U1436 (N_1436,In_1708,N_1352);
nand U1437 (N_1437,N_1123,N_1244);
xnor U1438 (N_1438,N_1302,N_1283);
and U1439 (N_1439,N_168,N_30);
or U1440 (N_1440,N_1336,In_1972);
xnor U1441 (N_1441,N_631,N_1152);
and U1442 (N_1442,In_1232,N_345);
nand U1443 (N_1443,In_1421,N_1122);
and U1444 (N_1444,N_458,N_786);
and U1445 (N_1445,N_403,In_2722);
and U1446 (N_1446,N_356,In_1323);
nor U1447 (N_1447,N_1150,N_228);
nor U1448 (N_1448,N_723,In_972);
xor U1449 (N_1449,N_1194,N_1154);
nor U1450 (N_1450,In_1315,N_1355);
or U1451 (N_1451,N_254,In_986);
nor U1452 (N_1452,In_1381,In_1974);
and U1453 (N_1453,In_1590,In_1963);
or U1454 (N_1454,In_2477,N_100);
or U1455 (N_1455,In_1560,N_505);
xor U1456 (N_1456,N_564,In_793);
xor U1457 (N_1457,In_2911,N_113);
nor U1458 (N_1458,N_1186,In_836);
nor U1459 (N_1459,In_1243,N_1075);
nor U1460 (N_1460,N_478,N_1237);
nor U1461 (N_1461,N_1238,N_1304);
and U1462 (N_1462,N_1209,In_2056);
nor U1463 (N_1463,N_282,In_1419);
xor U1464 (N_1464,N_1296,In_2145);
and U1465 (N_1465,In_2781,N_1370);
nand U1466 (N_1466,N_898,In_1229);
xnor U1467 (N_1467,N_573,N_498);
and U1468 (N_1468,In_239,N_416);
nor U1469 (N_1469,In_2860,In_1516);
nor U1470 (N_1470,In_2728,In_902);
and U1471 (N_1471,In_1195,N_1335);
nor U1472 (N_1472,In_2057,N_711);
nand U1473 (N_1473,N_872,In_1837);
xnor U1474 (N_1474,In_927,In_1773);
xnor U1475 (N_1475,N_1390,In_2334);
or U1476 (N_1476,In_1119,N_740);
and U1477 (N_1477,In_2562,In_937);
and U1478 (N_1478,In_2005,N_597);
nand U1479 (N_1479,N_1016,N_148);
nand U1480 (N_1480,In_1322,N_1290);
xnor U1481 (N_1481,In_1168,In_154);
xnor U1482 (N_1482,In_617,In_2216);
and U1483 (N_1483,N_847,N_1041);
and U1484 (N_1484,In_2993,In_2213);
nor U1485 (N_1485,In_1957,In_1456);
nand U1486 (N_1486,In_377,N_519);
xor U1487 (N_1487,N_217,In_2096);
xnor U1488 (N_1488,N_525,In_369);
nand U1489 (N_1489,In_909,N_807);
or U1490 (N_1490,N_257,In_692);
nor U1491 (N_1491,In_1320,In_2355);
and U1492 (N_1492,N_1183,In_2241);
xor U1493 (N_1493,N_676,N_5);
xor U1494 (N_1494,N_318,In_2007);
nor U1495 (N_1495,N_1147,In_2434);
or U1496 (N_1496,In_860,N_1084);
and U1497 (N_1497,In_1700,N_1177);
xor U1498 (N_1498,In_358,In_2740);
nand U1499 (N_1499,In_1053,N_1366);
xor U1500 (N_1500,In_924,N_879);
and U1501 (N_1501,In_2009,In_2426);
nand U1502 (N_1502,N_1145,N_504);
xor U1503 (N_1503,In_499,In_1933);
or U1504 (N_1504,N_1345,In_743);
and U1505 (N_1505,N_1077,In_316);
or U1506 (N_1506,N_1218,N_1287);
xnor U1507 (N_1507,In_2020,N_567);
xor U1508 (N_1508,In_1089,In_1788);
nor U1509 (N_1509,In_2155,N_1399);
and U1510 (N_1510,N_886,N_155);
and U1511 (N_1511,In_913,In_918);
xnor U1512 (N_1512,N_876,In_2492);
and U1513 (N_1513,N_705,N_1163);
or U1514 (N_1514,In_457,In_2684);
nand U1515 (N_1515,N_1054,N_1000);
nor U1516 (N_1516,In_1787,N_524);
or U1517 (N_1517,N_1205,In_2832);
nor U1518 (N_1518,In_1,N_521);
xnor U1519 (N_1519,In_43,N_1051);
or U1520 (N_1520,In_2656,N_819);
xor U1521 (N_1521,N_493,In_1847);
and U1522 (N_1522,In_1625,N_1243);
nor U1523 (N_1523,In_2975,N_407);
or U1524 (N_1524,In_2898,In_2959);
xnor U1525 (N_1525,In_408,In_974);
nand U1526 (N_1526,In_2810,N_918);
nor U1527 (N_1527,In_1362,N_637);
nand U1528 (N_1528,N_1224,N_630);
nor U1529 (N_1529,N_1357,In_2445);
and U1530 (N_1530,In_2196,N_1106);
nand U1531 (N_1531,In_247,In_1341);
or U1532 (N_1532,N_628,N_335);
or U1533 (N_1533,In_1051,In_1080);
and U1534 (N_1534,N_718,N_787);
and U1535 (N_1535,N_167,In_819);
nor U1536 (N_1536,N_946,In_2240);
and U1537 (N_1537,N_1249,In_1274);
xor U1538 (N_1538,N_1309,N_737);
and U1539 (N_1539,N_885,In_1576);
xor U1540 (N_1540,In_454,N_1378);
xor U1541 (N_1541,N_967,N_1270);
or U1542 (N_1542,N_849,In_728);
nand U1543 (N_1543,In_2306,In_1904);
and U1544 (N_1544,In_1540,In_2897);
or U1545 (N_1545,In_355,In_1169);
nand U1546 (N_1546,In_2615,N_125);
nand U1547 (N_1547,In_537,N_1317);
xnor U1548 (N_1548,N_1211,N_192);
xor U1549 (N_1549,N_37,N_1275);
and U1550 (N_1550,N_1105,In_2331);
nor U1551 (N_1551,N_1159,In_383);
and U1552 (N_1552,In_1575,In_1394);
xnor U1553 (N_1553,In_1610,In_1171);
and U1554 (N_1554,In_640,In_831);
or U1555 (N_1555,In_2654,In_583);
or U1556 (N_1556,N_944,In_2991);
xor U1557 (N_1557,In_1325,In_890);
xor U1558 (N_1558,In_1789,N_854);
nand U1559 (N_1559,N_980,In_2919);
and U1560 (N_1560,In_1513,In_1288);
nand U1561 (N_1561,N_1206,N_992);
nand U1562 (N_1562,N_315,In_562);
or U1563 (N_1563,N_554,In_0);
and U1564 (N_1564,N_1348,In_2400);
or U1565 (N_1565,In_1728,N_529);
or U1566 (N_1566,In_2295,N_763);
xnor U1567 (N_1567,In_2513,N_1288);
nand U1568 (N_1568,In_2120,In_2138);
nor U1569 (N_1569,N_734,In_2981);
nand U1570 (N_1570,N_1095,N_768);
xor U1571 (N_1571,In_606,N_766);
or U1572 (N_1572,In_2488,N_109);
xnor U1573 (N_1573,N_720,N_859);
or U1574 (N_1574,N_1327,N_1307);
or U1575 (N_1575,In_1920,In_2699);
or U1576 (N_1576,N_878,In_1344);
and U1577 (N_1577,N_1173,N_120);
and U1578 (N_1578,N_776,N_255);
and U1579 (N_1579,N_508,N_1008);
or U1580 (N_1580,N_882,In_1024);
xnor U1581 (N_1581,In_177,In_2131);
nand U1582 (N_1582,In_2114,N_563);
and U1583 (N_1583,N_1126,In_249);
nand U1584 (N_1584,In_693,N_1003);
nor U1585 (N_1585,In_1348,In_654);
and U1586 (N_1586,In_834,In_2436);
nand U1587 (N_1587,N_1397,In_613);
nand U1588 (N_1588,In_2101,In_71);
or U1589 (N_1589,In_1549,In_2008);
xor U1590 (N_1590,In_345,In_1277);
xor U1591 (N_1591,N_580,N_893);
nand U1592 (N_1592,N_127,In_437);
xor U1593 (N_1593,N_26,In_1085);
nor U1594 (N_1594,In_2841,N_1245);
or U1595 (N_1595,N_1119,N_163);
nand U1596 (N_1596,N_577,N_1364);
or U1597 (N_1597,In_48,In_1695);
xor U1598 (N_1598,N_1135,In_2576);
nor U1599 (N_1599,N_302,In_2491);
nor U1600 (N_1600,N_874,In_2261);
and U1601 (N_1601,In_2415,N_1221);
or U1602 (N_1602,N_1462,N_1256);
or U1603 (N_1603,N_304,In_153);
nor U1604 (N_1604,N_1526,In_1049);
and U1605 (N_1605,N_161,N_1027);
nand U1606 (N_1606,N_1313,N_551);
and U1607 (N_1607,In_1350,In_1725);
nand U1608 (N_1608,In_1985,In_1555);
nor U1609 (N_1609,N_772,N_1460);
nand U1610 (N_1610,In_2523,N_1536);
nor U1611 (N_1611,N_1017,In_221);
nor U1612 (N_1612,N_1567,In_415);
nand U1613 (N_1613,N_914,In_1372);
xnor U1614 (N_1614,In_1029,In_731);
nor U1615 (N_1615,N_1503,N_1278);
nor U1616 (N_1616,N_1239,N_1247);
nand U1617 (N_1617,In_1817,N_243);
or U1618 (N_1618,In_1164,N_101);
nor U1619 (N_1619,N_730,In_1680);
nor U1620 (N_1620,N_1382,N_1179);
and U1621 (N_1621,N_1408,In_1379);
and U1622 (N_1622,N_1565,N_1234);
xnor U1623 (N_1623,N_1450,N_399);
xor U1624 (N_1624,N_696,In_1131);
and U1625 (N_1625,In_2976,N_1504);
nand U1626 (N_1626,N_420,N_1052);
or U1627 (N_1627,In_2484,In_228);
xnor U1628 (N_1628,N_1299,N_1423);
or U1629 (N_1629,N_191,N_1429);
and U1630 (N_1630,In_1078,In_2989);
nand U1631 (N_1631,In_2274,N_692);
xnor U1632 (N_1632,In_1981,In_2034);
nand U1633 (N_1633,In_809,In_1141);
xor U1634 (N_1634,N_794,N_621);
and U1635 (N_1635,In_2910,N_1146);
nand U1636 (N_1636,N_1088,In_69);
xnor U1637 (N_1637,In_682,N_1235);
nor U1638 (N_1638,N_1471,In_2100);
nand U1639 (N_1639,N_195,In_216);
and U1640 (N_1640,N_1242,N_1061);
nand U1641 (N_1641,N_888,N_1131);
nor U1642 (N_1642,In_1702,N_783);
nand U1643 (N_1643,N_199,In_1405);
nand U1644 (N_1644,N_1557,N_1517);
or U1645 (N_1645,In_1065,N_1591);
or U1646 (N_1646,In_438,N_1321);
nor U1647 (N_1647,In_702,In_1339);
or U1648 (N_1648,In_715,N_364);
or U1649 (N_1649,In_237,N_1279);
nand U1650 (N_1650,N_1447,In_325);
xor U1651 (N_1651,In_487,N_932);
nand U1652 (N_1652,In_200,N_212);
or U1653 (N_1653,N_1251,In_157);
xnor U1654 (N_1654,N_1038,In_2208);
nor U1655 (N_1655,In_595,In_2531);
xnor U1656 (N_1656,N_913,N_1193);
nor U1657 (N_1657,In_2788,N_864);
xnor U1658 (N_1658,N_1455,In_2636);
nor U1659 (N_1659,In_2908,In_2964);
and U1660 (N_1660,N_1480,N_1192);
and U1661 (N_1661,In_1004,N_136);
or U1662 (N_1662,In_2966,N_1377);
and U1663 (N_1663,In_1759,N_1454);
nor U1664 (N_1664,N_1501,N_92);
nand U1665 (N_1665,N_910,In_2934);
nand U1666 (N_1666,In_1664,N_1513);
nand U1667 (N_1667,In_1689,N_1226);
xor U1668 (N_1668,N_1542,N_1232);
xor U1669 (N_1669,In_2072,In_1977);
or U1670 (N_1670,N_1293,N_1486);
or U1671 (N_1671,N_1329,N_1198);
nor U1672 (N_1672,N_1298,N_1342);
nand U1673 (N_1673,N_964,In_1228);
xnor U1674 (N_1674,N_596,N_712);
xnor U1675 (N_1675,In_804,N_889);
or U1676 (N_1676,In_1520,In_2383);
or U1677 (N_1677,In_2258,In_173);
nor U1678 (N_1678,In_2594,N_1376);
and U1679 (N_1679,N_1406,In_2143);
nor U1680 (N_1680,In_1152,N_757);
and U1681 (N_1681,N_50,N_1285);
or U1682 (N_1682,N_1569,N_941);
xor U1683 (N_1683,N_611,N_1258);
and U1684 (N_1684,In_645,In_1159);
or U1685 (N_1685,N_1094,In_2493);
and U1686 (N_1686,N_820,In_1351);
nand U1687 (N_1687,N_607,In_1945);
nor U1688 (N_1688,In_2254,In_2561);
nand U1689 (N_1689,N_78,In_381);
or U1690 (N_1690,N_1525,In_41);
or U1691 (N_1691,N_1322,In_1949);
nand U1692 (N_1692,In_2147,N_1575);
or U1693 (N_1693,N_1442,In_2170);
or U1694 (N_1694,N_1308,In_1968);
xnor U1695 (N_1695,N_1233,N_798);
and U1696 (N_1696,In_2351,N_862);
and U1697 (N_1697,In_1231,In_1236);
or U1698 (N_1698,In_878,N_1519);
nand U1699 (N_1699,In_2544,N_724);
and U1700 (N_1700,In_407,N_1543);
nand U1701 (N_1701,In_780,N_147);
nand U1702 (N_1702,In_1025,N_1257);
and U1703 (N_1703,N_9,In_922);
nand U1704 (N_1704,N_1492,N_1545);
xor U1705 (N_1705,In_256,N_1445);
nor U1706 (N_1706,N_1431,In_321);
xor U1707 (N_1707,In_1559,N_626);
nand U1708 (N_1708,In_391,N_1060);
xor U1709 (N_1709,N_115,N_351);
and U1710 (N_1710,In_1292,N_1594);
xor U1711 (N_1711,N_1403,In_2913);
xor U1712 (N_1712,N_1483,In_2315);
nand U1713 (N_1713,N_1325,In_2611);
nand U1714 (N_1714,N_539,N_660);
nand U1715 (N_1715,In_1444,N_972);
or U1716 (N_1716,N_1300,In_872);
nor U1717 (N_1717,In_422,N_1351);
nor U1718 (N_1718,N_83,N_816);
nand U1719 (N_1719,N_1530,In_721);
xor U1720 (N_1720,N_752,N_1099);
nand U1721 (N_1721,In_2674,N_1214);
or U1722 (N_1722,In_1733,In_2795);
and U1723 (N_1723,N_1380,In_1768);
nand U1724 (N_1724,In_459,In_380);
and U1725 (N_1725,N_1161,N_1059);
and U1726 (N_1726,N_960,In_482);
nor U1727 (N_1727,N_21,N_1074);
nand U1728 (N_1728,N_1113,N_1556);
or U1729 (N_1729,In_234,In_951);
or U1730 (N_1730,N_1369,N_1070);
or U1731 (N_1731,N_145,N_873);
nand U1732 (N_1732,In_908,N_931);
nor U1733 (N_1733,N_1081,In_2664);
or U1734 (N_1734,N_1117,N_1464);
or U1735 (N_1735,In_2835,N_146);
or U1736 (N_1736,In_2819,N_1023);
nand U1737 (N_1737,N_1393,N_1533);
xnor U1738 (N_1738,In_1294,In_1767);
nor U1739 (N_1739,N_453,N_697);
xor U1740 (N_1740,In_2813,In_1333);
xnor U1741 (N_1741,N_1392,N_196);
or U1742 (N_1742,In_192,In_1800);
xnor U1743 (N_1743,N_528,In_1470);
xor U1744 (N_1744,N_1282,N_1151);
xor U1745 (N_1745,In_2153,N_1030);
or U1746 (N_1746,In_1953,In_1823);
xnor U1747 (N_1747,N_962,N_1175);
or U1748 (N_1748,N_1494,N_331);
and U1749 (N_1749,N_1076,In_284);
nor U1750 (N_1750,N_422,N_852);
nor U1751 (N_1751,N_642,N_1465);
xor U1752 (N_1752,N_1435,In_2896);
or U1753 (N_1753,N_1166,N_48);
nor U1754 (N_1754,In_2262,In_1331);
nand U1755 (N_1755,In_1182,In_2221);
nand U1756 (N_1756,N_911,N_638);
nand U1757 (N_1757,N_1268,N_1340);
xnor U1758 (N_1758,N_1432,N_670);
nor U1759 (N_1759,In_761,In_703);
nor U1760 (N_1760,N_457,In_1928);
nor U1761 (N_1761,In_2555,In_409);
xnor U1762 (N_1762,N_203,N_635);
or U1763 (N_1763,N_382,In_55);
xnor U1764 (N_1764,N_1310,N_1383);
and U1765 (N_1765,In_1769,In_2041);
or U1766 (N_1766,N_201,N_1220);
nor U1767 (N_1767,N_1066,N_515);
nand U1768 (N_1768,N_1446,N_870);
and U1769 (N_1769,In_2963,N_1424);
and U1770 (N_1770,N_902,In_130);
and U1771 (N_1771,In_1878,N_1284);
xor U1772 (N_1772,In_491,N_1448);
nand U1773 (N_1773,N_954,In_2135);
or U1774 (N_1774,N_1420,N_1360);
or U1775 (N_1775,In_530,In_2437);
xnor U1776 (N_1776,In_1126,In_2393);
nor U1777 (N_1777,N_352,In_279);
nor U1778 (N_1778,N_1012,In_1249);
nand U1779 (N_1779,In_144,N_11);
and U1780 (N_1780,In_2323,N_979);
and U1781 (N_1781,In_789,In_1880);
nor U1782 (N_1782,In_553,In_1810);
nor U1783 (N_1783,N_369,N_480);
nand U1784 (N_1784,N_309,In_2603);
and U1785 (N_1785,In_2039,N_1395);
nand U1786 (N_1786,N_1453,In_2652);
nand U1787 (N_1787,N_209,In_888);
and U1788 (N_1788,N_1264,In_1330);
xor U1789 (N_1789,N_274,N_1421);
or U1790 (N_1790,N_728,N_565);
nor U1791 (N_1791,N_1597,N_869);
nor U1792 (N_1792,In_973,N_800);
nor U1793 (N_1793,In_148,N_1171);
nor U1794 (N_1794,N_1080,In_2255);
or U1795 (N_1795,N_868,In_1573);
and U1796 (N_1796,In_2679,N_576);
and U1797 (N_1797,In_1433,N_1555);
or U1798 (N_1798,In_1256,N_1153);
and U1799 (N_1799,In_2162,N_511);
xnor U1800 (N_1800,N_1487,N_251);
nor U1801 (N_1801,N_754,In_263);
and U1802 (N_1802,N_1761,In_1122);
nor U1803 (N_1803,N_1172,In_1824);
xnor U1804 (N_1804,In_894,N_595);
or U1805 (N_1805,N_1626,N_1636);
or U1806 (N_1806,N_1289,In_2033);
and U1807 (N_1807,In_1354,N_500);
nand U1808 (N_1808,In_2940,In_1476);
nand U1809 (N_1809,N_1491,N_1674);
nor U1810 (N_1810,In_598,N_679);
nand U1811 (N_1811,In_1683,In_2027);
nand U1812 (N_1812,N_1499,N_1647);
and U1813 (N_1813,In_1124,In_2077);
nor U1814 (N_1814,N_1616,N_218);
nand U1815 (N_1815,In_107,N_579);
and U1816 (N_1816,N_845,N_1384);
nor U1817 (N_1817,In_855,N_1318);
and U1818 (N_1818,In_848,N_860);
xnor U1819 (N_1819,In_507,N_1125);
and U1820 (N_1820,N_1755,N_858);
nand U1821 (N_1821,N_1768,N_1764);
xor U1822 (N_1822,In_1422,N_252);
xor U1823 (N_1823,In_2025,N_1071);
nand U1824 (N_1824,In_2065,N_1461);
nor U1825 (N_1825,N_1697,N_848);
and U1826 (N_1826,In_32,In_1994);
nor U1827 (N_1827,N_950,N_1774);
nor U1828 (N_1828,N_273,N_1564);
xnor U1829 (N_1829,N_836,N_1441);
and U1830 (N_1830,In_2868,N_1143);
nand U1831 (N_1831,N_1797,In_1079);
and U1832 (N_1832,In_53,N_1210);
and U1833 (N_1833,In_932,N_1609);
and U1834 (N_1834,In_410,In_2857);
nand U1835 (N_1835,In_1812,N_1531);
nand U1836 (N_1836,N_1439,In_841);
nand U1837 (N_1837,N_1231,N_366);
xnor U1838 (N_1838,N_1655,In_2497);
nor U1839 (N_1839,N_41,N_1760);
nand U1840 (N_1840,N_12,In_602);
xor U1841 (N_1841,N_1733,In_665);
xnor U1842 (N_1842,In_896,In_2345);
xor U1843 (N_1843,N_1770,N_483);
nor U1844 (N_1844,In_1508,N_1056);
nand U1845 (N_1845,N_317,N_1562);
nand U1846 (N_1846,N_1115,In_1779);
nor U1847 (N_1847,N_70,N_1651);
nor U1848 (N_1848,In_1179,N_1444);
nor U1849 (N_1849,In_2580,N_1748);
nand U1850 (N_1850,In_2073,N_242);
or U1851 (N_1851,N_938,N_1541);
nand U1852 (N_1852,In_1515,N_1769);
or U1853 (N_1853,N_250,In_2367);
nor U1854 (N_1854,In_2496,In_794);
nand U1855 (N_1855,In_331,N_1787);
nand U1856 (N_1856,In_2525,N_1693);
and U1857 (N_1857,N_1359,N_1111);
or U1858 (N_1858,In_1838,N_940);
nor U1859 (N_1859,N_1167,N_801);
nor U1860 (N_1860,In_933,N_952);
and U1861 (N_1861,In_2031,In_977);
nand U1862 (N_1862,N_1632,N_654);
or U1863 (N_1863,In_2109,N_1716);
or U1864 (N_1864,N_1596,N_1333);
xnor U1865 (N_1865,In_2816,N_969);
and U1866 (N_1866,N_1410,N_1758);
nor U1867 (N_1867,N_71,N_1101);
nand U1868 (N_1868,N_1662,In_578);
nor U1869 (N_1869,In_485,In_1438);
nand U1870 (N_1870,N_1488,In_1893);
nand U1871 (N_1871,N_1642,N_1165);
or U1872 (N_1872,N_1698,N_1681);
and U1873 (N_1873,N_1714,N_1763);
and U1874 (N_1874,In_1334,N_1676);
nand U1875 (N_1875,In_24,N_871);
xor U1876 (N_1876,N_1490,In_2558);
or U1877 (N_1877,In_480,N_1722);
xor U1878 (N_1878,In_1206,N_207);
nor U1879 (N_1879,N_1396,N_896);
and U1880 (N_1880,N_297,N_991);
and U1881 (N_1881,In_1665,In_874);
or U1882 (N_1882,N_604,N_396);
or U1883 (N_1883,N_775,N_1178);
or U1884 (N_1884,In_2844,N_648);
nor U1885 (N_1885,In_783,N_899);
and U1886 (N_1886,N_933,N_1326);
nor U1887 (N_1887,N_1103,In_462);
and U1888 (N_1888,In_826,In_2774);
and U1889 (N_1889,N_1598,N_1493);
and U1890 (N_1890,In_1756,In_612);
nand U1891 (N_1891,In_1895,N_1665);
or U1892 (N_1892,N_1731,N_1678);
and U1893 (N_1893,N_204,In_118);
nor U1894 (N_1894,N_1323,In_1843);
or U1895 (N_1895,In_1443,In_2696);
nand U1896 (N_1896,N_95,N_553);
and U1897 (N_1897,N_1643,N_999);
xor U1898 (N_1898,N_1560,N_1043);
nor U1899 (N_1899,N_901,In_2418);
or U1900 (N_1900,N_682,N_1628);
nor U1901 (N_1901,In_458,N_614);
nor U1902 (N_1902,N_1650,N_1682);
xor U1903 (N_1903,N_1417,N_1705);
nor U1904 (N_1904,N_1751,N_1623);
nor U1905 (N_1905,N_1240,N_1157);
nor U1906 (N_1906,In_1701,In_2851);
nor U1907 (N_1907,N_1011,In_1721);
xor U1908 (N_1908,In_1932,N_1202);
xnor U1909 (N_1909,N_561,N_289);
and U1910 (N_1910,N_1527,N_1739);
nand U1911 (N_1911,N_990,In_2166);
nor U1912 (N_1912,In_2248,In_2701);
xor U1913 (N_1913,N_1648,In_2712);
xnor U1914 (N_1914,N_1481,In_1158);
nand U1915 (N_1915,N_1343,N_985);
nor U1916 (N_1916,In_1656,N_169);
and U1917 (N_1917,N_1428,N_1271);
or U1918 (N_1918,N_1563,N_1255);
and U1919 (N_1919,N_540,N_997);
and U1920 (N_1920,N_764,N_1433);
nand U1921 (N_1921,N_1576,N_1398);
or U1922 (N_1922,N_1434,In_2665);
nor U1923 (N_1923,N_603,N_591);
nor U1924 (N_1924,N_1730,N_1466);
nand U1925 (N_1925,N_135,In_1821);
xnor U1926 (N_1926,N_1470,In_1310);
nand U1927 (N_1927,N_1736,In_954);
nand U1928 (N_1928,In_801,N_1702);
nand U1929 (N_1929,N_1387,N_1624);
xor U1930 (N_1930,In_2797,N_1415);
nor U1931 (N_1931,N_360,In_1894);
and U1932 (N_1932,N_509,N_1631);
xor U1933 (N_1933,N_1418,N_673);
nor U1934 (N_1934,N_1677,In_1739);
or U1935 (N_1935,N_1783,N_1586);
nand U1936 (N_1936,N_1427,N_1225);
nor U1937 (N_1937,N_1196,N_897);
nand U1938 (N_1938,In_2019,N_1580);
xor U1939 (N_1939,N_834,In_2378);
nor U1940 (N_1940,N_1506,N_165);
and U1941 (N_1941,In_1480,In_1038);
and U1942 (N_1942,N_1029,In_955);
xnor U1943 (N_1943,N_1469,In_1911);
xnor U1944 (N_1944,N_1645,N_1079);
xor U1945 (N_1945,In_464,N_838);
or U1946 (N_1946,N_389,N_1554);
nor U1947 (N_1947,In_2352,N_182);
nor U1948 (N_1948,In_1975,In_607);
nand U1949 (N_1949,In_42,N_1700);
nor U1950 (N_1950,N_748,N_970);
or U1951 (N_1951,N_1176,N_1771);
nor U1952 (N_1952,N_1049,In_990);
xor U1953 (N_1953,N_935,N_249);
and U1954 (N_1954,N_202,N_43);
xnor U1955 (N_1955,N_332,N_1708);
nand U1956 (N_1956,N_1223,N_1286);
nor U1957 (N_1957,N_1520,In_2340);
xnor U1958 (N_1958,In_724,N_1062);
nand U1959 (N_1959,N_1683,N_1653);
nand U1960 (N_1960,In_2714,N_1622);
and U1961 (N_1961,N_1356,N_1482);
xor U1962 (N_1962,In_2556,N_1757);
xnor U1963 (N_1963,N_1082,N_1727);
and U1964 (N_1964,N_831,N_1127);
xor U1965 (N_1965,N_432,In_336);
and U1966 (N_1966,In_1588,In_543);
and U1967 (N_1967,In_2307,N_1096);
nand U1968 (N_1968,In_1121,N_821);
xnor U1969 (N_1969,N_917,N_68);
or U1970 (N_1970,N_1615,N_1602);
xnor U1971 (N_1971,N_1798,In_772);
or U1972 (N_1972,In_389,N_923);
nand U1973 (N_1973,N_57,In_2831);
nor U1974 (N_1974,In_2092,In_2974);
nor U1975 (N_1975,N_1440,N_1640);
or U1976 (N_1976,N_1346,N_1656);
xnor U1977 (N_1977,In_2314,In_276);
nor U1978 (N_1978,In_1165,N_530);
and U1979 (N_1979,In_1259,N_1735);
xnor U1980 (N_1980,In_1965,N_1500);
and U1981 (N_1981,In_1679,In_2928);
or U1982 (N_1982,N_29,N_1456);
and U1983 (N_1983,In_2659,In_243);
nor U1984 (N_1984,In_67,N_1657);
nor U1985 (N_1985,N_60,In_2605);
xor U1986 (N_1986,N_1759,In_2811);
and U1987 (N_1987,N_1685,In_2958);
and U1988 (N_1988,N_1222,In_2640);
or U1989 (N_1989,In_1718,N_556);
nand U1990 (N_1990,In_2344,In_2906);
or U1991 (N_1991,N_867,N_963);
and U1992 (N_1992,N_1217,N_1375);
xnor U1993 (N_1993,N_1458,N_1672);
nand U1994 (N_1994,N_1568,N_575);
and U1995 (N_1995,In_89,In_1921);
and U1996 (N_1996,In_1225,N_1443);
nand U1997 (N_1997,In_1905,In_2085);
xor U1998 (N_1998,N_1711,In_448);
xnor U1999 (N_1999,In_66,N_651);
or U2000 (N_2000,N_1116,N_1720);
nand U2001 (N_2001,N_1195,N_1886);
nor U2002 (N_2002,In_1367,N_1025);
and U2003 (N_2003,N_1004,In_2272);
and U2004 (N_2004,N_1436,N_1507);
nand U2005 (N_2005,N_430,In_2082);
and U2006 (N_2006,N_1843,N_1031);
xor U2007 (N_2007,N_1834,N_983);
and U2008 (N_2008,N_610,N_1860);
nand U2009 (N_2009,In_1042,In_877);
and U2010 (N_2010,N_1524,In_339);
or U2011 (N_2011,N_841,In_2099);
xnor U2012 (N_2012,N_1841,N_1207);
nor U2013 (N_2013,In_569,N_1809);
nor U2014 (N_2014,N_1590,N_1960);
nor U2015 (N_2015,N_1476,N_1842);
xnor U2016 (N_2016,N_1849,N_361);
nor U2017 (N_2017,N_804,N_256);
or U2018 (N_2018,N_1955,N_1896);
or U2019 (N_2019,N_1895,N_1980);
nor U2020 (N_2020,N_1976,N_1799);
or U2021 (N_2021,N_1824,N_1573);
and U2022 (N_2022,In_2045,In_964);
and U2023 (N_2023,N_1581,N_1523);
and U2024 (N_2024,N_247,In_1661);
and U2025 (N_2025,N_1966,N_1404);
nor U2026 (N_2026,N_1857,N_1999);
nor U2027 (N_2027,N_1851,In_1984);
nor U2028 (N_2028,N_1848,N_904);
or U2029 (N_2029,N_451,In_660);
xnor U2030 (N_2030,In_994,N_1982);
and U2031 (N_2031,In_989,In_68);
and U2032 (N_2032,N_1856,N_1509);
and U2033 (N_2033,N_1930,In_781);
xnor U2034 (N_2034,N_947,In_1463);
and U2035 (N_2035,N_942,In_683);
nor U2036 (N_2036,N_1919,N_1859);
xor U2037 (N_2037,In_2769,N_22);
and U2038 (N_2038,In_1215,N_589);
xor U2039 (N_2039,In_1946,N_1766);
nand U2040 (N_2040,N_1337,N_1362);
xnor U2041 (N_2041,N_1929,In_207);
nor U2042 (N_2042,N_1670,N_1952);
nor U2043 (N_2043,N_1411,N_496);
and U2044 (N_2044,N_1847,In_871);
nor U2045 (N_2045,In_416,N_1889);
and U2046 (N_2046,N_1750,In_2534);
and U2047 (N_2047,N_1922,N_1600);
or U2048 (N_2048,N_1371,N_460);
nor U2049 (N_2049,N_1388,In_85);
or U2050 (N_2050,In_2268,N_1553);
nand U2051 (N_2051,N_1934,N_1475);
xnor U2052 (N_2052,N_1511,In_956);
and U2053 (N_2053,N_1883,N_709);
and U2054 (N_2054,N_982,N_1725);
or U2055 (N_2055,In_2049,N_1971);
nor U2056 (N_2056,N_1838,N_1891);
and U2057 (N_2057,N_1986,N_731);
and U2058 (N_2058,N_1295,N_751);
or U2059 (N_2059,N_1667,In_1815);
nand U2060 (N_2060,N_936,N_1505);
and U2061 (N_2061,N_1821,N_1752);
xnor U2062 (N_2062,In_330,In_269);
and U2063 (N_2063,In_2760,In_779);
or U2064 (N_2064,N_1998,N_1913);
xnor U2065 (N_2065,In_1819,N_1861);
nand U2066 (N_2066,N_1712,In_224);
nand U2067 (N_2067,In_2405,N_1219);
and U2068 (N_2068,N_665,N_1579);
xor U2069 (N_2069,In_2607,In_1103);
xnor U2070 (N_2070,N_1280,In_520);
and U2071 (N_2071,In_753,N_1142);
or U2072 (N_2072,In_1371,In_1201);
nor U2073 (N_2073,In_2441,N_1620);
and U2074 (N_2074,N_1110,N_1729);
and U2075 (N_2075,N_1721,N_1900);
or U2076 (N_2076,N_1818,N_34);
xor U2077 (N_2077,In_2681,N_1669);
nand U2078 (N_2078,N_1710,N_1473);
nor U2079 (N_2079,N_1426,In_1342);
xnor U2080 (N_2080,N_1254,N_833);
xor U2081 (N_2081,In_2289,In_469);
nor U2082 (N_2082,In_2922,N_1361);
nand U2083 (N_2083,In_1458,In_1678);
xor U2084 (N_2084,In_2517,N_1920);
and U2085 (N_2085,In_2017,In_250);
xnor U2086 (N_2086,N_1338,N_1118);
and U2087 (N_2087,N_584,N_1498);
and U2088 (N_2088,N_1102,In_79);
nand U2089 (N_2089,N_557,N_704);
and U2090 (N_2090,N_1539,N_645);
xnor U2091 (N_2091,N_741,N_1741);
nor U2092 (N_2092,In_2621,N_1032);
nor U2093 (N_2093,N_1584,N_1508);
nor U2094 (N_2094,N_1261,N_647);
and U2095 (N_2095,In_287,N_1412);
nand U2096 (N_2096,N_1897,In_1811);
and U2097 (N_2097,N_1121,N_1989);
or U2098 (N_2098,In_1466,N_1561);
nand U2099 (N_2099,In_2587,N_1301);
and U2100 (N_2100,N_1241,N_1819);
nor U2101 (N_2101,N_1635,N_1034);
nand U2102 (N_2102,N_1540,N_1713);
nand U2103 (N_2103,In_1411,N_429);
and U2104 (N_2104,In_2375,N_722);
xnor U2105 (N_2105,N_785,N_1664);
xor U2106 (N_2106,N_1687,In_77);
or U2107 (N_2107,N_1695,N_1825);
and U2108 (N_2108,N_1967,N_1953);
or U2109 (N_2109,N_1495,N_1778);
nor U2110 (N_2110,N_1690,In_159);
or U2111 (N_2111,In_597,N_1806);
and U2112 (N_2112,N_1324,In_839);
nand U2113 (N_2113,In_2823,N_1024);
xor U2114 (N_2114,In_2335,N_1814);
or U2115 (N_2115,N_1888,In_2947);
or U2116 (N_2116,N_1686,N_1840);
nor U2117 (N_2117,N_65,In_2924);
xnor U2118 (N_2118,In_2438,N_957);
xnor U2119 (N_2119,N_1529,N_1582);
xor U2120 (N_2120,N_1935,N_1386);
xor U2121 (N_2121,In_2672,N_404);
nand U2122 (N_2122,In_2087,N_1035);
or U2123 (N_2123,N_1067,N_592);
and U2124 (N_2124,N_1717,N_67);
or U2125 (N_2125,N_1253,N_1855);
or U2126 (N_2126,N_1744,N_814);
nor U2127 (N_2127,N_544,In_2982);
and U2128 (N_2128,N_1201,N_357);
and U2129 (N_2129,N_1274,In_1598);
and U2130 (N_2130,N_1740,N_1184);
or U2131 (N_2131,N_44,N_771);
nor U2132 (N_2132,N_817,N_671);
nand U2133 (N_2133,N_1532,N_1820);
and U2134 (N_2134,N_1850,N_1871);
nand U2135 (N_2135,N_1518,In_18);
or U2136 (N_2136,N_1331,N_1909);
xnor U2137 (N_2137,N_1993,N_1684);
xnor U2138 (N_2138,N_824,N_1835);
nor U2139 (N_2139,In_2459,N_474);
and U2140 (N_2140,N_1601,N_1742);
xnor U2141 (N_2141,N_1407,N_1754);
xnor U2142 (N_2142,N_1899,In_1178);
nand U2143 (N_2143,In_1338,In_1698);
or U2144 (N_2144,N_1605,In_319);
nand U2145 (N_2145,N_877,N_6);
and U2146 (N_2146,N_781,In_2083);
nand U2147 (N_2147,In_1857,N_1793);
nand U2148 (N_2148,In_2683,In_2999);
nor U2149 (N_2149,N_1954,N_1063);
or U2150 (N_2150,N_1964,N_1800);
nand U2151 (N_2151,N_1815,N_1617);
nor U2152 (N_2152,N_1782,N_1230);
xnor U2153 (N_2153,N_1864,N_1260);
and U2154 (N_2154,In_1452,N_461);
or U2155 (N_2155,N_1957,N_1663);
xnor U2156 (N_2156,In_601,In_1276);
xor U2157 (N_2157,N_1879,In_353);
and U2158 (N_2158,N_1773,N_1991);
or U2159 (N_2159,In_240,N_1502);
nand U2160 (N_2160,N_594,N_1633);
or U2161 (N_2161,N_1040,N_1547);
and U2162 (N_2162,N_1463,N_1784);
nand U2163 (N_2163,In_384,In_143);
or U2164 (N_2164,N_1276,N_1625);
xor U2165 (N_2165,In_822,N_1882);
xnor U2166 (N_2166,N_177,N_1923);
and U2167 (N_2167,N_813,In_675);
nor U2168 (N_2168,N_326,N_1158);
nand U2169 (N_2169,N_1887,In_1370);
xnor U2170 (N_2170,N_1621,N_1199);
and U2171 (N_2171,In_388,N_1694);
nand U2172 (N_2172,N_1789,In_2920);
nand U2173 (N_2173,N_721,N_989);
and U2174 (N_2174,N_338,N_1409);
nor U2175 (N_2175,In_265,N_1965);
nor U2176 (N_2176,N_1876,In_1383);
xor U2177 (N_2177,In_2163,N_925);
or U2178 (N_2178,N_1689,N_1983);
xnor U2179 (N_2179,N_1939,In_2224);
or U2180 (N_2180,N_1457,In_1192);
and U2181 (N_2181,N_1707,In_727);
or U2182 (N_2182,In_1175,N_1994);
nand U2183 (N_2183,N_1303,In_1914);
nor U2184 (N_2184,In_2458,N_1660);
xor U2185 (N_2185,N_1981,In_1072);
or U2186 (N_2186,N_1484,N_1973);
nand U2187 (N_2187,In_444,N_681);
or U2188 (N_2188,N_1614,N_1925);
nor U2189 (N_2189,N_1595,N_1827);
and U2190 (N_2190,N_959,N_1385);
nor U2191 (N_2191,N_656,N_1772);
and U2192 (N_2192,N_330,In_1417);
nor U2193 (N_2193,In_2978,N_1259);
or U2194 (N_2194,In_1044,N_1915);
and U2195 (N_2195,In_2646,N_1852);
and U2196 (N_2196,In_1536,In_2946);
and U2197 (N_2197,In_1472,N_1696);
or U2198 (N_2198,N_1802,N_1552);
nand U2199 (N_2199,N_1585,N_1608);
or U2200 (N_2200,N_427,N_1837);
xnor U2201 (N_2201,N_1570,N_2074);
xnor U2202 (N_2202,N_1853,N_1574);
or U2203 (N_2203,N_2045,N_1902);
nor U2204 (N_2204,N_1917,N_379);
nand U2205 (N_2205,In_452,N_1306);
xor U2206 (N_2206,In_1777,In_805);
nand U2207 (N_2207,In_1793,N_1449);
or U2208 (N_2208,N_1354,N_1846);
nor U2209 (N_2209,N_1528,N_2031);
nand U2210 (N_2210,In_1493,N_971);
and U2211 (N_2211,N_2187,In_398);
nand U2212 (N_2212,In_558,N_2182);
nor U2213 (N_2213,In_210,In_2686);
nand U2214 (N_2214,N_2113,N_1641);
and U2215 (N_2215,N_464,In_351);
nand U2216 (N_2216,N_2083,In_1156);
nand U2217 (N_2217,N_1794,N_1918);
nand U2218 (N_2218,N_1777,N_118);
nand U2219 (N_2219,In_1203,N_2073);
nor U2220 (N_2220,N_2119,N_439);
nand U2221 (N_2221,N_1612,N_545);
nand U2222 (N_2222,N_2033,N_2046);
nor U2223 (N_2223,N_716,N_922);
xnor U2224 (N_2224,In_2845,In_2363);
nor U2225 (N_2225,N_2111,N_1330);
xor U2226 (N_2226,In_1803,N_1691);
nand U2227 (N_2227,N_2011,N_2084);
and U2228 (N_2228,N_472,In_1722);
nand U2229 (N_2229,N_2092,N_887);
nor U2230 (N_2230,N_2036,N_2012);
nand U2231 (N_2231,N_2148,N_2002);
or U2232 (N_2232,N_1940,N_1812);
or U2233 (N_2233,N_2000,N_1037);
nand U2234 (N_2234,N_1832,In_2727);
xor U2235 (N_2235,N_1941,N_1137);
nand U2236 (N_2236,N_857,N_1910);
or U2237 (N_2237,N_1350,In_1645);
xnor U2238 (N_2238,N_1968,N_1969);
and U2239 (N_2239,N_2065,N_2149);
nand U2240 (N_2240,N_1884,N_2060);
nand U2241 (N_2241,N_2024,N_675);
and U2242 (N_2242,N_1963,In_270);
and U2243 (N_2243,N_2150,N_443);
nand U2244 (N_2244,N_762,N_1875);
xor U2245 (N_2245,In_1867,N_537);
xor U2246 (N_2246,N_1938,In_2952);
and U2247 (N_2247,N_1367,N_1828);
nor U2248 (N_2248,N_2064,In_436);
or U2249 (N_2249,N_1817,N_1956);
nor U2250 (N_2250,In_1507,N_1639);
or U2251 (N_2251,N_1951,In_2708);
or U2252 (N_2252,In_45,N_1666);
xor U2253 (N_2253,N_1155,N_1497);
nand U2254 (N_2254,N_1961,N_1212);
and U2255 (N_2255,N_2166,In_283);
xnor U2256 (N_2256,In_1535,N_2079);
xor U2257 (N_2257,N_945,N_2070);
or U2258 (N_2258,N_2136,N_324);
nor U2259 (N_2259,In_404,In_2379);
nor U2260 (N_2260,In_773,N_2191);
and U2261 (N_2261,N_2014,N_2030);
and U2262 (N_2262,N_1452,N_2062);
xnor U2263 (N_2263,N_2123,N_2124);
xnor U2264 (N_2264,N_1607,N_208);
or U2265 (N_2265,N_1743,In_412);
or U2266 (N_2266,N_1200,N_1937);
or U2267 (N_2267,In_995,N_1992);
xor U2268 (N_2268,In_354,N_446);
xnor U2269 (N_2269,N_533,N_1534);
and U2270 (N_2270,N_482,N_398);
nor U2271 (N_2271,N_31,N_1363);
and U2272 (N_2272,N_1272,N_1893);
nor U2273 (N_2273,N_1521,In_375);
xnor U2274 (N_2274,N_760,N_1732);
and U2275 (N_2275,N_2087,N_1141);
or U2276 (N_2276,In_1646,N_2165);
or U2277 (N_2277,N_1114,N_2193);
nor U2278 (N_2278,N_1671,N_1320);
or U2279 (N_2279,N_855,N_1381);
nand U2280 (N_2280,In_1160,N_644);
or U2281 (N_2281,N_1215,In_605);
or U2282 (N_2282,N_1312,N_1946);
xnor U2283 (N_2283,N_1745,N_1489);
nor U2284 (N_2284,N_738,N_1803);
and U2285 (N_2285,N_1826,In_2796);
and U2286 (N_2286,N_1905,N_1924);
and U2287 (N_2287,In_1116,In_1128);
xnor U2288 (N_2288,N_2044,N_1109);
nand U2289 (N_2289,N_894,N_1401);
nor U2290 (N_2290,N_2169,N_2180);
nor U2291 (N_2291,N_1629,N_2186);
xor U2292 (N_2292,N_1191,N_1588);
xor U2293 (N_2293,In_1149,N_1990);
xor U2294 (N_2294,N_2027,N_2078);
nor U2295 (N_2295,N_2163,N_1372);
xor U2296 (N_2296,In_397,In_647);
nor U2297 (N_2297,N_2048,N_1638);
or U2298 (N_2298,N_2039,N_2196);
xnor U2299 (N_2299,N_1901,N_2132);
or U2300 (N_2300,N_535,N_1868);
or U2301 (N_2301,N_2199,In_2597);
or U2302 (N_2302,N_1865,N_2109);
nor U2303 (N_2303,N_2181,N_1593);
nor U2304 (N_2304,N_1064,In_2429);
nor U2305 (N_2305,N_2146,N_1311);
nand U2306 (N_2306,N_2049,N_1416);
nand U2307 (N_2307,N_517,N_892);
nand U2308 (N_2308,In_883,N_1373);
xnor U2309 (N_2309,In_2410,N_1894);
xor U2310 (N_2310,N_2029,N_1092);
nor U2311 (N_2311,N_1927,N_2098);
and U2312 (N_2312,N_2157,N_826);
and U2313 (N_2313,N_2104,In_2871);
nor U2314 (N_2314,In_897,N_1767);
nand U2315 (N_2315,N_2183,N_1911);
nand U2316 (N_2316,N_1979,In_629);
nor U2317 (N_2317,N_2054,N_2058);
and U2318 (N_2318,In_2267,N_2001);
nand U2319 (N_2319,N_1180,N_966);
and U2320 (N_2320,N_235,N_1675);
and U2321 (N_2321,N_2171,In_2037);
nand U2322 (N_2322,N_1975,N_1422);
or U2323 (N_2323,In_2688,In_1593);
nand U2324 (N_2324,N_180,N_1906);
and U2325 (N_2325,N_1592,In_2412);
or U2326 (N_2326,N_2016,N_1559);
nand U2327 (N_2327,N_1190,N_1830);
nand U2328 (N_2328,N_2122,N_1822);
nor U2329 (N_2329,N_2097,In_667);
nand U2330 (N_2330,N_2082,N_2094);
nor U2331 (N_2331,N_1057,N_1472);
nor U2332 (N_2332,In_2812,N_2035);
xnor U2333 (N_2333,N_1870,In_2741);
nand U2334 (N_2334,N_1018,N_1451);
nor U2335 (N_2335,N_2134,N_1878);
nor U2336 (N_2336,N_1583,N_1341);
or U2337 (N_2337,N_1188,In_2710);
and U2338 (N_2338,N_1880,N_1549);
xor U2339 (N_2339,In_1979,N_1985);
xor U2340 (N_2340,N_2099,N_2188);
or U2341 (N_2341,N_1213,N_701);
xnor U2342 (N_2342,N_2075,In_1214);
xor U2343 (N_2343,N_1236,N_2009);
nor U2344 (N_2344,N_791,N_1936);
nand U2345 (N_2345,N_2063,N_2189);
xnor U2346 (N_2346,N_1050,N_1810);
nor U2347 (N_2347,In_1407,In_447);
xnor U2348 (N_2348,In_815,In_1776);
nor U2349 (N_2349,N_1972,N_1263);
or U2350 (N_2350,N_2057,N_1419);
nand U2351 (N_2351,N_2155,N_1292);
and U2352 (N_2352,N_1305,N_582);
nor U2353 (N_2353,N_1589,N_2056);
xor U2354 (N_2354,N_978,N_1831);
and U2355 (N_2355,N_2088,N_2017);
and U2356 (N_2356,N_2141,N_1389);
or U2357 (N_2357,N_2138,N_1203);
or U2358 (N_2358,N_1294,N_1546);
or U2359 (N_2359,N_1942,N_1634);
and U2360 (N_2360,N_2178,N_1281);
and U2361 (N_2361,N_1349,N_1808);
or U2362 (N_2362,N_613,N_2096);
nor U2363 (N_2363,N_1478,N_1997);
nor U2364 (N_2364,In_1027,In_609);
or U2365 (N_2365,N_424,N_2071);
nand U2366 (N_2366,N_1266,N_1347);
nor U2367 (N_2367,N_2154,N_1514);
nand U2368 (N_2368,In_2720,N_2089);
xor U2369 (N_2369,N_1715,N_1943);
xor U2370 (N_2370,N_2010,In_1127);
nor U2371 (N_2371,In_2887,N_1932);
nor U2372 (N_2372,N_2105,N_1039);
or U2373 (N_2373,N_2106,N_2137);
xor U2374 (N_2374,N_2179,N_1610);
nand U2375 (N_2375,N_2197,In_1997);
nor U2376 (N_2376,N_1788,N_2061);
or U2377 (N_2377,N_916,N_1316);
xor U2378 (N_2378,N_1984,N_1100);
nand U2379 (N_2379,N_1646,N_2121);
nor U2380 (N_2380,In_982,In_611);
xnor U2381 (N_2381,N_1904,In_2585);
and U2382 (N_2382,N_1661,In_2630);
and U2383 (N_2383,N_2195,N_1988);
nand U2384 (N_2384,N_900,N_2015);
xnor U2385 (N_2385,N_1344,N_2115);
or U2386 (N_2386,N_1587,N_930);
or U2387 (N_2387,N_2172,N_1400);
and U2388 (N_2388,In_500,N_1468);
or U2389 (N_2389,N_2151,In_2609);
or U2390 (N_2390,N_1854,N_2147);
or U2391 (N_2391,In_907,In_337);
nor U2392 (N_2392,N_2130,N_620);
nand U2393 (N_2393,N_1873,N_440);
nand U2394 (N_2394,N_1762,N_2038);
xor U2395 (N_2395,N_2167,N_1673);
xnor U2396 (N_2396,N_1977,N_1069);
nor U2397 (N_2397,N_2023,N_1679);
or U2398 (N_2398,N_2008,In_2631);
nand U2399 (N_2399,In_1316,N_1866);
nor U2400 (N_2400,N_2135,In_766);
nand U2401 (N_2401,N_1829,In_1879);
and U2402 (N_2402,N_2365,In_2793);
or U2403 (N_2403,N_2028,N_1086);
nand U2404 (N_2404,N_2375,N_546);
xnor U2405 (N_2405,N_1044,N_2228);
nand U2406 (N_2406,N_2275,N_2076);
nand U2407 (N_2407,N_2328,N_1379);
nor U2408 (N_2408,N_1391,N_2170);
and U2409 (N_2409,In_84,N_1958);
and U2410 (N_2410,In_1194,N_2072);
nor U2411 (N_2411,N_1823,N_2290);
or U2412 (N_2412,N_2037,N_2203);
nand U2413 (N_2413,N_2093,N_1659);
or U2414 (N_2414,N_2286,N_2140);
and U2415 (N_2415,N_2378,N_2144);
xnor U2416 (N_2416,In_472,N_1944);
or U2417 (N_2417,N_1414,In_713);
nand U2418 (N_2418,N_2370,N_1737);
xor U2419 (N_2419,N_1619,N_2209);
and U2420 (N_2420,N_2204,N_2337);
or U2421 (N_2421,N_735,N_1959);
nor U2422 (N_2422,N_2260,In_1948);
or U2423 (N_2423,N_1749,N_2329);
nand U2424 (N_2424,N_2224,N_2312);
xor U2425 (N_2425,N_1949,In_735);
nor U2426 (N_2426,N_2251,N_2342);
nor U2427 (N_2427,N_1765,In_967);
nand U2428 (N_2428,N_2327,N_1833);
xnor U2429 (N_2429,N_2139,N_1262);
and U2430 (N_2430,N_688,N_2053);
nor U2431 (N_2431,N_2067,N_2091);
and U2432 (N_2432,In_2419,N_2395);
or U2433 (N_2433,N_2040,In_1635);
and U2434 (N_2434,N_1189,N_2086);
xnor U2435 (N_2435,N_2217,N_2116);
nor U2436 (N_2436,N_2102,N_2296);
and U2437 (N_2437,N_94,N_1734);
nor U2438 (N_2438,N_2325,N_2185);
nor U2439 (N_2439,In_1233,N_1869);
nand U2440 (N_2440,N_1724,N_2314);
nor U2441 (N_2441,N_1019,N_1950);
nand U2442 (N_2442,N_2288,N_1692);
nand U2443 (N_2443,N_2214,N_2158);
xnor U2444 (N_2444,N_2285,N_1394);
nor U2445 (N_2445,N_1006,N_2153);
xnor U2446 (N_2446,N_1903,N_2284);
and U2447 (N_2447,N_2164,N_1571);
nand U2448 (N_2448,N_2252,In_957);
and U2449 (N_2449,N_2263,In_428);
or U2450 (N_2450,N_2388,N_2085);
or U2451 (N_2451,N_2095,N_1611);
nand U2452 (N_2452,N_2194,N_1962);
nand U2453 (N_2453,N_2384,N_2225);
or U2454 (N_2454,N_2353,N_2381);
nand U2455 (N_2455,In_1374,N_1947);
xnor U2456 (N_2456,N_1786,N_2277);
nor U2457 (N_2457,N_1738,N_2289);
xor U2458 (N_2458,N_1719,N_2198);
nand U2459 (N_2459,In_1412,N_2025);
nand U2460 (N_2460,N_2059,N_1680);
nor U2461 (N_2461,N_1785,N_2266);
nand U2462 (N_2462,N_2018,N_2250);
and U2463 (N_2463,N_2269,N_1926);
nor U2464 (N_2464,N_1816,N_2175);
or U2465 (N_2465,N_2253,N_2192);
nand U2466 (N_2466,N_1485,N_1668);
nor U2467 (N_2467,N_2320,N_1208);
and U2468 (N_2468,N_2338,N_1603);
xnor U2469 (N_2469,N_2131,N_2077);
xor U2470 (N_2470,N_1987,N_1046);
or U2471 (N_2471,N_1353,N_2377);
nor U2472 (N_2472,In_1939,In_1852);
nand U2473 (N_2473,N_2133,N_2021);
nor U2474 (N_2474,N_861,N_0);
nand U2475 (N_2475,N_2068,N_1867);
nand U2476 (N_2476,N_2243,N_1780);
or U2477 (N_2477,N_2280,N_2223);
and U2478 (N_2478,N_2219,In_1415);
or U2479 (N_2479,N_1402,N_2398);
or U2480 (N_2480,In_1366,N_1438);
nor U2481 (N_2481,N_828,N_1558);
and U2482 (N_2482,In_1173,N_1368);
xnor U2483 (N_2483,N_1858,In_2786);
nand U2484 (N_2484,In_1327,In_1579);
xnor U2485 (N_2485,N_1756,N_1162);
nor U2486 (N_2486,N_2259,In_2098);
nand U2487 (N_2487,N_1995,N_1872);
or U2488 (N_2488,In_52,N_2055);
nor U2489 (N_2489,N_1718,N_1933);
nand U2490 (N_2490,N_2262,N_1477);
xnor U2491 (N_2491,N_2069,In_2456);
nand U2492 (N_2492,N_2202,In_1145);
and U2493 (N_2493,N_128,N_1544);
nand U2494 (N_2494,N_1170,In_767);
and U2495 (N_2495,In_2925,N_2249);
nand U2496 (N_2496,In_2726,N_2354);
xor U2497 (N_2497,N_2293,N_2368);
xor U2498 (N_2498,N_1914,N_2352);
or U2499 (N_2499,N_2316,N_2032);
and U2500 (N_2500,N_2246,N_2235);
xor U2501 (N_2501,N_1836,N_2399);
and U2502 (N_2502,N_1319,In_2239);
or U2503 (N_2503,N_2389,N_2369);
or U2504 (N_2504,In_1139,N_2184);
or U2505 (N_2505,N_1314,N_903);
or U2506 (N_2506,N_2218,In_33);
or U2507 (N_2507,N_2200,N_2173);
nand U2508 (N_2508,N_1928,In_2294);
and U2509 (N_2509,N_1430,N_2367);
xnor U2510 (N_2510,N_2387,N_2274);
or U2511 (N_2511,N_1916,N_1792);
or U2512 (N_2512,N_2222,N_2080);
nor U2513 (N_2513,N_2341,In_2995);
nor U2514 (N_2514,N_1654,N_2310);
nor U2515 (N_2515,N_2291,N_2361);
nor U2516 (N_2516,N_2227,In_1982);
xnor U2517 (N_2517,N_2207,In_1191);
nand U2518 (N_2518,In_2601,N_1813);
and U2519 (N_2519,N_2278,N_2346);
xnor U2520 (N_2520,N_2255,N_2306);
and U2521 (N_2521,N_2240,N_2383);
or U2522 (N_2522,N_1613,N_1021);
or U2523 (N_2523,N_248,In_440);
nor U2524 (N_2524,N_2208,In_2203);
nand U2525 (N_2525,N_2216,N_1658);
nand U2526 (N_2526,N_1474,N_2372);
nand U2527 (N_2527,N_1839,N_588);
nand U2528 (N_2528,N_2343,N_2344);
and U2529 (N_2529,N_1413,In_1361);
nand U2530 (N_2530,N_2373,N_2363);
nand U2531 (N_2531,N_2101,N_2270);
and U2532 (N_2532,N_1801,N_2160);
or U2533 (N_2533,N_1703,N_2351);
or U2534 (N_2534,N_1181,In_2373);
or U2535 (N_2535,N_1578,N_2239);
nor U2536 (N_2536,N_1709,N_245);
xnor U2537 (N_2537,N_2128,N_2386);
nand U2538 (N_2538,N_2005,In_2836);
and U2539 (N_2539,N_1898,N_1845);
nand U2540 (N_2540,N_2234,N_2305);
nor U2541 (N_2541,N_2292,N_2256);
nand U2542 (N_2542,N_2339,N_2265);
or U2543 (N_2543,N_1630,N_2254);
nor U2544 (N_2544,N_2364,N_1577);
nand U2545 (N_2545,N_2242,N_1467);
nand U2546 (N_2546,N_1204,N_1807);
and U2547 (N_2547,In_1533,In_1747);
nor U2548 (N_2548,N_1874,N_2297);
and U2549 (N_2549,N_2392,N_2231);
or U2550 (N_2550,N_1512,N_1315);
xnor U2551 (N_2551,N_2051,N_1881);
nand U2552 (N_2552,N_1974,In_225);
nor U2553 (N_2553,N_2298,N_2307);
nor U2554 (N_2554,N_1877,N_2248);
or U2555 (N_2555,N_1907,N_2385);
nand U2556 (N_2556,N_1496,In_2505);
and U2557 (N_2557,N_2340,N_1291);
and U2558 (N_2558,N_2348,N_759);
nor U2559 (N_2559,N_765,N_2319);
and U2560 (N_2560,N_2350,N_2022);
nor U2561 (N_2561,N_2301,N_2007);
and U2562 (N_2562,In_1222,N_843);
nand U2563 (N_2563,N_91,In_479);
and U2564 (N_2564,N_1796,N_1479);
and U2565 (N_2565,N_463,In_1425);
nor U2566 (N_2566,N_1863,N_322);
and U2567 (N_2567,N_2004,In_661);
and U2568 (N_2568,N_2271,In_180);
or U2569 (N_2569,N_1649,N_2013);
nand U2570 (N_2570,In_343,N_2229);
and U2571 (N_2571,N_2110,N_2283);
xor U2572 (N_2572,N_2322,N_2333);
xnor U2573 (N_2573,N_1890,N_2108);
nand U2574 (N_2574,N_1297,N_1538);
nand U2575 (N_2575,N_2220,In_961);
and U2576 (N_2576,N_1701,In_2530);
or U2577 (N_2577,N_291,N_1652);
and U2578 (N_2578,N_2161,N_2126);
nand U2579 (N_2579,N_2118,N_2230);
nor U2580 (N_2580,N_1515,N_2349);
nor U2581 (N_2581,In_1554,N_1781);
or U2582 (N_2582,N_2331,N_2366);
nor U2583 (N_2583,N_2226,N_2317);
and U2584 (N_2584,N_2213,N_1921);
or U2585 (N_2585,In_2526,N_2332);
or U2586 (N_2586,N_1599,N_2355);
nand U2587 (N_2587,N_2311,N_1128);
and U2588 (N_2588,N_2176,N_2303);
nor U2589 (N_2589,N_2282,N_2168);
nor U2590 (N_2590,N_2391,N_1776);
and U2591 (N_2591,N_1425,N_1138);
nand U2592 (N_2592,N_1537,N_143);
nor U2593 (N_2593,N_1779,N_2026);
and U2594 (N_2594,N_2066,N_1459);
nand U2595 (N_2595,N_1535,N_284);
nor U2596 (N_2596,N_2052,N_1728);
nand U2597 (N_2597,N_2143,N_1704);
and U2598 (N_2598,In_2960,N_2020);
or U2599 (N_2599,N_853,N_1931);
nand U2600 (N_2600,N_2530,N_1010);
nand U2601 (N_2601,N_2512,N_2257);
or U2602 (N_2602,In_778,N_2003);
or U2603 (N_2603,N_2439,N_2447);
xnor U2604 (N_2604,N_2520,N_2465);
nand U2605 (N_2605,N_1548,In_101);
nor U2606 (N_2606,N_2529,N_1885);
and U2607 (N_2607,N_1437,N_1250);
nand U2608 (N_2608,N_2458,N_2413);
or U2609 (N_2609,N_2345,N_2300);
and U2610 (N_2610,N_2485,N_2397);
and U2611 (N_2611,N_2431,N_1948);
nor U2612 (N_2612,N_2238,N_2569);
xnor U2613 (N_2613,N_2390,N_2047);
nand U2614 (N_2614,N_2174,N_1229);
nor U2615 (N_2615,N_2334,N_2568);
xor U2616 (N_2616,N_2446,N_2444);
nor U2617 (N_2617,N_2394,N_1606);
xnor U2618 (N_2618,N_2244,N_2575);
and U2619 (N_2619,N_905,In_2266);
or U2620 (N_2620,In_2915,N_753);
or U2621 (N_2621,N_2587,N_2455);
nand U2622 (N_2622,N_2479,N_2453);
or U2623 (N_2623,N_2117,N_2445);
xnor U2624 (N_2624,N_2464,N_2495);
nor U2625 (N_2625,N_2423,N_2524);
nor U2626 (N_2626,N_2299,N_2090);
or U2627 (N_2627,N_2505,N_2491);
and U2628 (N_2628,N_1970,N_2177);
and U2629 (N_2629,N_2518,N_2599);
xor U2630 (N_2630,N_2376,N_2483);
nand U2631 (N_2631,N_2509,N_2501);
and U2632 (N_2632,N_1073,In_1460);
xor U2633 (N_2633,N_2407,N_2412);
or U2634 (N_2634,N_1637,N_2573);
nand U2635 (N_2635,N_1790,N_2245);
xnor U2636 (N_2636,N_2490,N_1516);
and U2637 (N_2637,In_2137,In_2563);
or U2638 (N_2638,In_362,N_2579);
xnor U2639 (N_2639,N_2578,N_2205);
nor U2640 (N_2640,In_941,N_2409);
and U2641 (N_2641,N_2496,N_2454);
and U2642 (N_2642,N_2503,N_1746);
nand U2643 (N_2643,N_2374,N_920);
and U2644 (N_2644,N_2211,N_2466);
nor U2645 (N_2645,N_2233,N_2410);
xnor U2646 (N_2646,N_2556,N_2210);
and U2647 (N_2647,N_1912,N_2324);
xnor U2648 (N_2648,N_2484,N_2145);
and U2649 (N_2649,N_2081,N_2549);
nor U2650 (N_2650,N_2521,N_1945);
and U2651 (N_2651,N_2156,N_2577);
and U2652 (N_2652,N_2586,N_2557);
nor U2653 (N_2653,N_2534,N_178);
xor U2654 (N_2654,N_2393,N_2330);
and U2655 (N_2655,N_2459,N_144);
or U2656 (N_2656,In_2212,N_2538);
xor U2657 (N_2657,N_2563,N_2335);
nand U2658 (N_2658,N_2507,N_2241);
and U2659 (N_2659,N_2129,N_2437);
nand U2660 (N_2660,In_506,N_2519);
nand U2661 (N_2661,N_2467,N_2434);
xnor U2662 (N_2662,N_2498,N_2585);
or U2663 (N_2663,N_1604,In_1526);
nor U2664 (N_2664,N_2576,N_2565);
nand U2665 (N_2665,N_2588,N_2318);
and U2666 (N_2666,N_2492,N_2500);
nand U2667 (N_2667,N_2589,N_2514);
nand U2668 (N_2668,N_2287,N_1566);
nor U2669 (N_2669,N_2449,N_2405);
and U2670 (N_2670,N_2594,N_2379);
nor U2671 (N_2671,N_2571,N_2120);
nor U2672 (N_2672,In_1566,N_2206);
and U2673 (N_2673,N_2508,N_2424);
nor U2674 (N_2674,N_2542,N_2416);
nand U2675 (N_2675,N_2510,N_2247);
xnor U2676 (N_2676,In_768,N_2050);
nor U2677 (N_2677,N_2477,N_2236);
nor U2678 (N_2678,N_2125,N_2564);
and U2679 (N_2679,N_2162,N_1908);
nand U2680 (N_2680,N_2572,N_2237);
and U2681 (N_2681,N_2598,N_2476);
xor U2682 (N_2682,N_2273,N_2567);
and U2683 (N_2683,N_2313,N_1726);
nand U2684 (N_2684,N_2550,N_1405);
and U2685 (N_2685,N_1510,N_2489);
nand U2686 (N_2686,N_2295,N_2415);
nor U2687 (N_2687,N_2516,N_2480);
and U2688 (N_2688,N_2566,N_2441);
nor U2689 (N_2689,In_1637,N_2482);
or U2690 (N_2690,N_2435,N_773);
nor U2691 (N_2691,N_926,N_2506);
or U2692 (N_2692,N_2593,N_2100);
nand U2693 (N_2693,N_2457,N_2553);
nand U2694 (N_2694,N_2315,In_2433);
nand U2695 (N_2695,N_2570,N_103);
nand U2696 (N_2696,N_2360,N_2422);
nor U2697 (N_2697,N_1328,N_2212);
nor U2698 (N_2698,N_2540,N_2401);
or U2699 (N_2699,N_2411,N_1164);
and U2700 (N_2700,N_2433,N_1551);
and U2701 (N_2701,N_2474,N_2404);
nand U2702 (N_2702,N_1723,N_2536);
and U2703 (N_2703,N_2432,N_2430);
nor U2704 (N_2704,N_2362,N_2418);
xnor U2705 (N_2705,N_1706,N_2408);
and U2706 (N_2706,N_2419,N_2438);
or U2707 (N_2707,N_2561,In_2490);
nor U2708 (N_2708,N_2487,N_1795);
nand U2709 (N_2709,N_1747,N_2400);
and U2710 (N_2710,N_2535,N_2470);
or U2711 (N_2711,N_2543,N_2582);
and U2712 (N_2712,N_2551,In_193);
nand U2713 (N_2713,In_1528,N_2041);
nand U2714 (N_2714,N_1805,N_2190);
xnor U2715 (N_2715,N_2481,N_2347);
nor U2716 (N_2716,In_581,N_2309);
nand U2717 (N_2717,N_2525,N_2426);
or U2718 (N_2718,N_2554,N_1804);
nor U2719 (N_2719,N_1374,N_2471);
nand U2720 (N_2720,N_2473,N_2380);
xor U2721 (N_2721,N_2159,N_2281);
nor U2722 (N_2722,N_2201,N_2595);
xnor U2723 (N_2723,N_2427,N_2522);
nand U2724 (N_2724,N_2531,N_2420);
and U2725 (N_2725,N_2494,N_2451);
and U2726 (N_2726,N_2468,N_2526);
and U2727 (N_2727,N_2359,N_2356);
or U2728 (N_2728,N_639,N_2462);
and U2729 (N_2729,In_72,N_2463);
nand U2730 (N_2730,N_2114,N_2103);
and U2731 (N_2731,N_2429,N_2590);
or U2732 (N_2732,N_2517,N_2596);
xor U2733 (N_2733,N_2502,N_2499);
xnor U2734 (N_2734,N_2460,N_2261);
or U2735 (N_2735,N_812,N_2493);
nor U2736 (N_2736,N_2560,N_2232);
or U2737 (N_2737,N_2539,N_2034);
or U2738 (N_2738,N_2396,N_2469);
and U2739 (N_2739,In_2000,N_1978);
or U2740 (N_2740,N_2436,N_2107);
and U2741 (N_2741,N_2541,N_2545);
and U2742 (N_2742,N_2537,N_2548);
nand U2743 (N_2743,N_2547,N_2440);
and U2744 (N_2744,N_2006,N_2450);
xnor U2745 (N_2745,N_2267,N_1688);
and U2746 (N_2746,N_2357,N_2279);
nand U2747 (N_2747,N_2488,N_2580);
xnor U2748 (N_2748,N_2417,N_1550);
nand U2749 (N_2749,N_2527,N_2528);
xor U2750 (N_2750,N_2574,N_2555);
or U2751 (N_2751,N_1332,N_1791);
xnor U2752 (N_2752,N_1168,N_1248);
xnor U2753 (N_2753,N_1892,N_1811);
xor U2754 (N_2754,N_2448,N_2127);
nor U2755 (N_2755,N_72,N_2276);
xnor U2756 (N_2756,N_2294,In_518);
and U2757 (N_2757,N_1216,In_698);
or U2758 (N_2758,N_2472,N_2583);
xor U2759 (N_2759,N_2532,N_2215);
xnor U2760 (N_2760,N_2597,N_2456);
nand U2761 (N_2761,N_2546,N_1134);
or U2762 (N_2762,N_2584,N_2421);
nor U2763 (N_2763,N_2358,N_2268);
and U2764 (N_2764,N_2533,N_1699);
nor U2765 (N_2765,N_593,N_2414);
xor U2766 (N_2766,N_2478,In_798);
xnor U2767 (N_2767,N_2592,N_2523);
or U2768 (N_2768,N_2042,N_2264);
and U2769 (N_2769,N_2428,N_2308);
and U2770 (N_2770,N_2562,N_2152);
xnor U2771 (N_2771,In_1658,N_2461);
and U2772 (N_2772,N_2591,N_1862);
nand U2773 (N_2773,N_2043,N_2581);
nor U2774 (N_2774,N_1174,In_717);
nor U2775 (N_2775,N_2258,N_1618);
nand U2776 (N_2776,N_2559,N_2552);
or U2777 (N_2777,N_2336,N_2544);
and U2778 (N_2778,N_2019,N_2403);
and U2779 (N_2779,N_2304,N_2504);
or U2780 (N_2780,N_2323,N_1572);
nand U2781 (N_2781,N_1753,N_2326);
nor U2782 (N_2782,N_2272,N_2371);
nor U2783 (N_2783,N_2511,N_2382);
or U2784 (N_2784,In_2040,N_706);
and U2785 (N_2785,N_2443,N_2221);
nand U2786 (N_2786,N_2558,In_2669);
nand U2787 (N_2787,N_2475,N_2402);
and U2788 (N_2788,N_1009,N_2142);
xor U2789 (N_2789,In_318,In_769);
nand U2790 (N_2790,N_1627,N_2321);
nor U2791 (N_2791,N_1644,N_2425);
nand U2792 (N_2792,N_1265,N_2513);
xor U2793 (N_2793,N_1522,N_2452);
and U2794 (N_2794,N_2442,N_2497);
nand U2795 (N_2795,N_2515,N_2486);
nor U2796 (N_2796,In_2869,N_1844);
and U2797 (N_2797,N_1775,N_1996);
or U2798 (N_2798,N_2406,N_2302);
and U2799 (N_2799,In_2765,N_2112);
nor U2800 (N_2800,N_2798,N_2666);
and U2801 (N_2801,N_2772,N_2708);
nand U2802 (N_2802,N_2786,N_2789);
and U2803 (N_2803,N_2717,N_2671);
or U2804 (N_2804,N_2799,N_2796);
or U2805 (N_2805,N_2711,N_2605);
nor U2806 (N_2806,N_2654,N_2655);
and U2807 (N_2807,N_2738,N_2609);
nand U2808 (N_2808,N_2795,N_2653);
nand U2809 (N_2809,N_2704,N_2767);
nand U2810 (N_2810,N_2714,N_2752);
xor U2811 (N_2811,N_2647,N_2601);
nor U2812 (N_2812,N_2707,N_2744);
or U2813 (N_2813,N_2793,N_2614);
xor U2814 (N_2814,N_2762,N_2748);
nor U2815 (N_2815,N_2760,N_2642);
nor U2816 (N_2816,N_2768,N_2742);
nand U2817 (N_2817,N_2718,N_2709);
xor U2818 (N_2818,N_2723,N_2763);
or U2819 (N_2819,N_2741,N_2615);
nor U2820 (N_2820,N_2694,N_2706);
or U2821 (N_2821,N_2715,N_2616);
and U2822 (N_2822,N_2753,N_2667);
and U2823 (N_2823,N_2766,N_2610);
and U2824 (N_2824,N_2620,N_2764);
xor U2825 (N_2825,N_2749,N_2683);
or U2826 (N_2826,N_2630,N_2665);
xnor U2827 (N_2827,N_2774,N_2693);
nand U2828 (N_2828,N_2735,N_2769);
nand U2829 (N_2829,N_2751,N_2644);
xor U2830 (N_2830,N_2690,N_2660);
or U2831 (N_2831,N_2602,N_2780);
nor U2832 (N_2832,N_2739,N_2612);
nand U2833 (N_2833,N_2728,N_2695);
and U2834 (N_2834,N_2737,N_2781);
xor U2835 (N_2835,N_2663,N_2696);
nor U2836 (N_2836,N_2678,N_2726);
xnor U2837 (N_2837,N_2623,N_2758);
or U2838 (N_2838,N_2621,N_2626);
nor U2839 (N_2839,N_2727,N_2681);
nor U2840 (N_2840,N_2661,N_2674);
nor U2841 (N_2841,N_2776,N_2757);
xnor U2842 (N_2842,N_2638,N_2677);
nand U2843 (N_2843,N_2669,N_2622);
xor U2844 (N_2844,N_2759,N_2619);
nor U2845 (N_2845,N_2668,N_2747);
xnor U2846 (N_2846,N_2659,N_2771);
nand U2847 (N_2847,N_2656,N_2794);
nand U2848 (N_2848,N_2785,N_2632);
or U2849 (N_2849,N_2617,N_2697);
xnor U2850 (N_2850,N_2636,N_2713);
nor U2851 (N_2851,N_2652,N_2756);
and U2852 (N_2852,N_2761,N_2724);
nor U2853 (N_2853,N_2603,N_2754);
nand U2854 (N_2854,N_2664,N_2740);
and U2855 (N_2855,N_2604,N_2650);
nand U2856 (N_2856,N_2710,N_2635);
or U2857 (N_2857,N_2645,N_2676);
or U2858 (N_2858,N_2699,N_2733);
or U2859 (N_2859,N_2691,N_2732);
and U2860 (N_2860,N_2779,N_2673);
and U2861 (N_2861,N_2649,N_2631);
or U2862 (N_2862,N_2729,N_2721);
xor U2863 (N_2863,N_2746,N_2606);
xnor U2864 (N_2864,N_2736,N_2790);
nand U2865 (N_2865,N_2687,N_2797);
and U2866 (N_2866,N_2648,N_2702);
or U2867 (N_2867,N_2731,N_2698);
and U2868 (N_2868,N_2705,N_2689);
nand U2869 (N_2869,N_2672,N_2675);
xor U2870 (N_2870,N_2788,N_2703);
and U2871 (N_2871,N_2686,N_2777);
xor U2872 (N_2872,N_2607,N_2716);
nor U2873 (N_2873,N_2633,N_2700);
xor U2874 (N_2874,N_2627,N_2641);
xor U2875 (N_2875,N_2685,N_2624);
or U2876 (N_2876,N_2611,N_2778);
nor U2877 (N_2877,N_2765,N_2670);
nand U2878 (N_2878,N_2782,N_2783);
nand U2879 (N_2879,N_2629,N_2734);
and U2880 (N_2880,N_2634,N_2719);
nand U2881 (N_2881,N_2628,N_2688);
and U2882 (N_2882,N_2684,N_2750);
xor U2883 (N_2883,N_2657,N_2643);
or U2884 (N_2884,N_2600,N_2712);
and U2885 (N_2885,N_2680,N_2787);
nor U2886 (N_2886,N_2792,N_2784);
nand U2887 (N_2887,N_2730,N_2770);
or U2888 (N_2888,N_2618,N_2608);
and U2889 (N_2889,N_2651,N_2646);
nand U2890 (N_2890,N_2692,N_2640);
xor U2891 (N_2891,N_2682,N_2775);
and U2892 (N_2892,N_2720,N_2679);
or U2893 (N_2893,N_2755,N_2613);
nor U2894 (N_2894,N_2722,N_2773);
xnor U2895 (N_2895,N_2701,N_2662);
nand U2896 (N_2896,N_2637,N_2743);
xnor U2897 (N_2897,N_2625,N_2725);
xnor U2898 (N_2898,N_2658,N_2745);
xor U2899 (N_2899,N_2791,N_2639);
or U2900 (N_2900,N_2668,N_2709);
nand U2901 (N_2901,N_2689,N_2674);
nand U2902 (N_2902,N_2799,N_2674);
nor U2903 (N_2903,N_2608,N_2610);
and U2904 (N_2904,N_2677,N_2632);
nor U2905 (N_2905,N_2740,N_2737);
xor U2906 (N_2906,N_2669,N_2730);
or U2907 (N_2907,N_2747,N_2737);
or U2908 (N_2908,N_2706,N_2702);
xor U2909 (N_2909,N_2620,N_2604);
xor U2910 (N_2910,N_2796,N_2732);
nand U2911 (N_2911,N_2645,N_2654);
nor U2912 (N_2912,N_2619,N_2749);
or U2913 (N_2913,N_2678,N_2658);
and U2914 (N_2914,N_2743,N_2620);
and U2915 (N_2915,N_2761,N_2699);
nor U2916 (N_2916,N_2764,N_2610);
xor U2917 (N_2917,N_2614,N_2764);
or U2918 (N_2918,N_2668,N_2682);
or U2919 (N_2919,N_2728,N_2739);
xor U2920 (N_2920,N_2764,N_2704);
or U2921 (N_2921,N_2703,N_2660);
nor U2922 (N_2922,N_2741,N_2705);
xnor U2923 (N_2923,N_2624,N_2663);
and U2924 (N_2924,N_2693,N_2714);
nand U2925 (N_2925,N_2664,N_2658);
or U2926 (N_2926,N_2635,N_2648);
nand U2927 (N_2927,N_2628,N_2611);
xor U2928 (N_2928,N_2658,N_2621);
nand U2929 (N_2929,N_2719,N_2754);
and U2930 (N_2930,N_2632,N_2604);
nor U2931 (N_2931,N_2689,N_2649);
or U2932 (N_2932,N_2684,N_2627);
nor U2933 (N_2933,N_2797,N_2604);
and U2934 (N_2934,N_2622,N_2652);
xnor U2935 (N_2935,N_2744,N_2682);
xor U2936 (N_2936,N_2762,N_2685);
nand U2937 (N_2937,N_2696,N_2760);
nor U2938 (N_2938,N_2761,N_2619);
and U2939 (N_2939,N_2624,N_2748);
and U2940 (N_2940,N_2768,N_2621);
or U2941 (N_2941,N_2635,N_2775);
and U2942 (N_2942,N_2628,N_2793);
nor U2943 (N_2943,N_2610,N_2723);
nand U2944 (N_2944,N_2615,N_2601);
and U2945 (N_2945,N_2736,N_2722);
xor U2946 (N_2946,N_2733,N_2718);
or U2947 (N_2947,N_2669,N_2765);
and U2948 (N_2948,N_2753,N_2631);
and U2949 (N_2949,N_2759,N_2712);
nor U2950 (N_2950,N_2640,N_2610);
nand U2951 (N_2951,N_2643,N_2765);
nor U2952 (N_2952,N_2710,N_2774);
or U2953 (N_2953,N_2699,N_2646);
and U2954 (N_2954,N_2686,N_2606);
xor U2955 (N_2955,N_2679,N_2772);
xnor U2956 (N_2956,N_2647,N_2774);
or U2957 (N_2957,N_2653,N_2658);
or U2958 (N_2958,N_2731,N_2789);
nand U2959 (N_2959,N_2739,N_2614);
and U2960 (N_2960,N_2784,N_2793);
or U2961 (N_2961,N_2773,N_2600);
and U2962 (N_2962,N_2652,N_2612);
nand U2963 (N_2963,N_2660,N_2730);
or U2964 (N_2964,N_2771,N_2742);
and U2965 (N_2965,N_2649,N_2711);
and U2966 (N_2966,N_2677,N_2649);
and U2967 (N_2967,N_2671,N_2723);
nand U2968 (N_2968,N_2735,N_2750);
nand U2969 (N_2969,N_2677,N_2755);
xor U2970 (N_2970,N_2754,N_2721);
xnor U2971 (N_2971,N_2733,N_2777);
or U2972 (N_2972,N_2724,N_2609);
or U2973 (N_2973,N_2671,N_2639);
nor U2974 (N_2974,N_2740,N_2787);
xor U2975 (N_2975,N_2737,N_2694);
xnor U2976 (N_2976,N_2701,N_2624);
and U2977 (N_2977,N_2731,N_2773);
nor U2978 (N_2978,N_2632,N_2612);
or U2979 (N_2979,N_2755,N_2605);
nand U2980 (N_2980,N_2669,N_2799);
xnor U2981 (N_2981,N_2738,N_2791);
nor U2982 (N_2982,N_2755,N_2722);
xor U2983 (N_2983,N_2691,N_2739);
or U2984 (N_2984,N_2674,N_2677);
nand U2985 (N_2985,N_2603,N_2674);
or U2986 (N_2986,N_2714,N_2713);
and U2987 (N_2987,N_2644,N_2787);
nand U2988 (N_2988,N_2640,N_2650);
nand U2989 (N_2989,N_2748,N_2601);
and U2990 (N_2990,N_2774,N_2645);
nand U2991 (N_2991,N_2631,N_2659);
nor U2992 (N_2992,N_2600,N_2721);
nor U2993 (N_2993,N_2652,N_2745);
xor U2994 (N_2994,N_2622,N_2624);
and U2995 (N_2995,N_2616,N_2663);
or U2996 (N_2996,N_2618,N_2708);
nor U2997 (N_2997,N_2653,N_2623);
nand U2998 (N_2998,N_2663,N_2604);
xnor U2999 (N_2999,N_2654,N_2679);
and U3000 (N_3000,N_2806,N_2804);
and U3001 (N_3001,N_2842,N_2987);
or U3002 (N_3002,N_2927,N_2908);
nor U3003 (N_3003,N_2932,N_2925);
nor U3004 (N_3004,N_2862,N_2906);
nand U3005 (N_3005,N_2881,N_2857);
nor U3006 (N_3006,N_2919,N_2817);
nand U3007 (N_3007,N_2922,N_2975);
xor U3008 (N_3008,N_2943,N_2879);
xnor U3009 (N_3009,N_2845,N_2966);
nand U3010 (N_3010,N_2977,N_2989);
or U3011 (N_3011,N_2935,N_2980);
nand U3012 (N_3012,N_2838,N_2848);
nand U3013 (N_3013,N_2897,N_2931);
nand U3014 (N_3014,N_2871,N_2813);
xor U3015 (N_3015,N_2979,N_2946);
nor U3016 (N_3016,N_2913,N_2985);
nor U3017 (N_3017,N_2974,N_2903);
and U3018 (N_3018,N_2971,N_2996);
xnor U3019 (N_3019,N_2866,N_2885);
and U3020 (N_3020,N_2991,N_2942);
nor U3021 (N_3021,N_2868,N_2835);
xor U3022 (N_3022,N_2983,N_2993);
xnor U3023 (N_3023,N_2940,N_2967);
and U3024 (N_3024,N_2962,N_2877);
xnor U3025 (N_3025,N_2970,N_2800);
or U3026 (N_3026,N_2961,N_2957);
nand U3027 (N_3027,N_2861,N_2811);
and U3028 (N_3028,N_2917,N_2854);
nor U3029 (N_3029,N_2909,N_2934);
xor U3030 (N_3030,N_2926,N_2949);
nor U3031 (N_3031,N_2803,N_2812);
or U3032 (N_3032,N_2981,N_2910);
xnor U3033 (N_3033,N_2965,N_2954);
nand U3034 (N_3034,N_2890,N_2828);
xnor U3035 (N_3035,N_2907,N_2850);
xor U3036 (N_3036,N_2911,N_2814);
or U3037 (N_3037,N_2815,N_2825);
nor U3038 (N_3038,N_2976,N_2819);
nand U3039 (N_3039,N_2978,N_2809);
nor U3040 (N_3040,N_2928,N_2923);
xor U3041 (N_3041,N_2872,N_2956);
xnor U3042 (N_3042,N_2924,N_2888);
nand U3043 (N_3043,N_2990,N_2846);
xnor U3044 (N_3044,N_2941,N_2905);
or U3045 (N_3045,N_2858,N_2834);
or U3046 (N_3046,N_2883,N_2859);
or U3047 (N_3047,N_2822,N_2824);
xor U3048 (N_3048,N_2849,N_2829);
xnor U3049 (N_3049,N_2831,N_2856);
nand U3050 (N_3050,N_2999,N_2944);
xnor U3051 (N_3051,N_2843,N_2982);
xnor U3052 (N_3052,N_2865,N_2900);
nand U3053 (N_3053,N_2832,N_2802);
xnor U3054 (N_3054,N_2867,N_2875);
or U3055 (N_3055,N_2847,N_2972);
or U3056 (N_3056,N_2869,N_2807);
nor U3057 (N_3057,N_2860,N_2904);
nand U3058 (N_3058,N_2889,N_2953);
or U3059 (N_3059,N_2986,N_2950);
xor U3060 (N_3060,N_2998,N_2844);
and U3061 (N_3061,N_2892,N_2820);
nand U3062 (N_3062,N_2988,N_2948);
xnor U3063 (N_3063,N_2805,N_2994);
and U3064 (N_3064,N_2836,N_2968);
nand U3065 (N_3065,N_2851,N_2930);
or U3066 (N_3066,N_2898,N_2833);
and U3067 (N_3067,N_2893,N_2837);
nand U3068 (N_3068,N_2826,N_2921);
xor U3069 (N_3069,N_2830,N_2863);
and U3070 (N_3070,N_2918,N_2840);
and U3071 (N_3071,N_2852,N_2959);
xor U3072 (N_3072,N_2945,N_2992);
xor U3073 (N_3073,N_2902,N_2855);
or U3074 (N_3074,N_2969,N_2821);
xnor U3075 (N_3075,N_2929,N_2947);
nand U3076 (N_3076,N_2870,N_2880);
or U3077 (N_3077,N_2997,N_2882);
nor U3078 (N_3078,N_2895,N_2896);
xor U3079 (N_3079,N_2939,N_2958);
nor U3080 (N_3080,N_2920,N_2874);
nor U3081 (N_3081,N_2973,N_2936);
nand U3082 (N_3082,N_2823,N_2876);
nand U3083 (N_3083,N_2886,N_2818);
nor U3084 (N_3084,N_2853,N_2964);
xnor U3085 (N_3085,N_2884,N_2916);
or U3086 (N_3086,N_2960,N_2887);
nand U3087 (N_3087,N_2827,N_2914);
nor U3088 (N_3088,N_2901,N_2995);
nor U3089 (N_3089,N_2937,N_2912);
nor U3090 (N_3090,N_2894,N_2963);
xor U3091 (N_3091,N_2915,N_2873);
and U3092 (N_3092,N_2801,N_2891);
and U3093 (N_3093,N_2878,N_2951);
and U3094 (N_3094,N_2955,N_2839);
nor U3095 (N_3095,N_2808,N_2810);
xor U3096 (N_3096,N_2938,N_2899);
and U3097 (N_3097,N_2841,N_2984);
or U3098 (N_3098,N_2952,N_2864);
nor U3099 (N_3099,N_2933,N_2816);
nor U3100 (N_3100,N_2964,N_2801);
nand U3101 (N_3101,N_2903,N_2981);
nor U3102 (N_3102,N_2957,N_2887);
nor U3103 (N_3103,N_2923,N_2806);
nor U3104 (N_3104,N_2969,N_2961);
nor U3105 (N_3105,N_2896,N_2929);
nand U3106 (N_3106,N_2807,N_2961);
xor U3107 (N_3107,N_2807,N_2931);
nand U3108 (N_3108,N_2859,N_2853);
xnor U3109 (N_3109,N_2855,N_2809);
nand U3110 (N_3110,N_2992,N_2908);
and U3111 (N_3111,N_2934,N_2952);
nor U3112 (N_3112,N_2971,N_2801);
nand U3113 (N_3113,N_2893,N_2930);
or U3114 (N_3114,N_2880,N_2952);
nand U3115 (N_3115,N_2904,N_2838);
or U3116 (N_3116,N_2953,N_2883);
nand U3117 (N_3117,N_2842,N_2961);
xnor U3118 (N_3118,N_2810,N_2906);
nand U3119 (N_3119,N_2828,N_2860);
and U3120 (N_3120,N_2970,N_2840);
xnor U3121 (N_3121,N_2943,N_2864);
and U3122 (N_3122,N_2966,N_2890);
or U3123 (N_3123,N_2983,N_2945);
xor U3124 (N_3124,N_2949,N_2883);
and U3125 (N_3125,N_2872,N_2917);
nand U3126 (N_3126,N_2841,N_2993);
or U3127 (N_3127,N_2873,N_2990);
xnor U3128 (N_3128,N_2927,N_2969);
and U3129 (N_3129,N_2880,N_2878);
nor U3130 (N_3130,N_2821,N_2958);
nand U3131 (N_3131,N_2879,N_2979);
xor U3132 (N_3132,N_2940,N_2875);
nand U3133 (N_3133,N_2931,N_2891);
nand U3134 (N_3134,N_2908,N_2842);
or U3135 (N_3135,N_2852,N_2818);
nor U3136 (N_3136,N_2883,N_2980);
xor U3137 (N_3137,N_2992,N_2852);
or U3138 (N_3138,N_2963,N_2921);
nor U3139 (N_3139,N_2874,N_2923);
xor U3140 (N_3140,N_2897,N_2979);
and U3141 (N_3141,N_2812,N_2876);
nor U3142 (N_3142,N_2833,N_2967);
and U3143 (N_3143,N_2865,N_2898);
nor U3144 (N_3144,N_2968,N_2929);
or U3145 (N_3145,N_2955,N_2989);
xor U3146 (N_3146,N_2921,N_2991);
nand U3147 (N_3147,N_2810,N_2896);
nand U3148 (N_3148,N_2895,N_2857);
xor U3149 (N_3149,N_2938,N_2923);
nand U3150 (N_3150,N_2943,N_2981);
xnor U3151 (N_3151,N_2981,N_2867);
nand U3152 (N_3152,N_2817,N_2905);
nor U3153 (N_3153,N_2824,N_2886);
xor U3154 (N_3154,N_2806,N_2888);
xnor U3155 (N_3155,N_2939,N_2850);
nor U3156 (N_3156,N_2854,N_2828);
and U3157 (N_3157,N_2888,N_2949);
and U3158 (N_3158,N_2854,N_2930);
or U3159 (N_3159,N_2946,N_2988);
nand U3160 (N_3160,N_2874,N_2949);
and U3161 (N_3161,N_2985,N_2937);
xnor U3162 (N_3162,N_2870,N_2877);
nand U3163 (N_3163,N_2913,N_2843);
xnor U3164 (N_3164,N_2897,N_2814);
nor U3165 (N_3165,N_2930,N_2835);
xnor U3166 (N_3166,N_2912,N_2831);
and U3167 (N_3167,N_2867,N_2881);
xnor U3168 (N_3168,N_2985,N_2908);
nand U3169 (N_3169,N_2902,N_2957);
nor U3170 (N_3170,N_2906,N_2871);
or U3171 (N_3171,N_2850,N_2857);
nor U3172 (N_3172,N_2903,N_2946);
nor U3173 (N_3173,N_2950,N_2909);
nor U3174 (N_3174,N_2884,N_2848);
and U3175 (N_3175,N_2947,N_2965);
and U3176 (N_3176,N_2913,N_2941);
xnor U3177 (N_3177,N_2845,N_2994);
nor U3178 (N_3178,N_2961,N_2800);
nand U3179 (N_3179,N_2988,N_2860);
nand U3180 (N_3180,N_2834,N_2977);
nand U3181 (N_3181,N_2989,N_2924);
or U3182 (N_3182,N_2882,N_2852);
and U3183 (N_3183,N_2982,N_2821);
and U3184 (N_3184,N_2940,N_2888);
and U3185 (N_3185,N_2845,N_2935);
nand U3186 (N_3186,N_2815,N_2915);
or U3187 (N_3187,N_2901,N_2812);
nor U3188 (N_3188,N_2998,N_2915);
nor U3189 (N_3189,N_2865,N_2812);
and U3190 (N_3190,N_2867,N_2962);
xnor U3191 (N_3191,N_2850,N_2904);
xnor U3192 (N_3192,N_2897,N_2913);
nand U3193 (N_3193,N_2996,N_2892);
xor U3194 (N_3194,N_2843,N_2880);
or U3195 (N_3195,N_2933,N_2955);
or U3196 (N_3196,N_2958,N_2873);
xnor U3197 (N_3197,N_2889,N_2873);
nand U3198 (N_3198,N_2953,N_2817);
nand U3199 (N_3199,N_2843,N_2860);
xor U3200 (N_3200,N_3003,N_3178);
nand U3201 (N_3201,N_3108,N_3164);
nand U3202 (N_3202,N_3009,N_3105);
nor U3203 (N_3203,N_3194,N_3045);
xnor U3204 (N_3204,N_3093,N_3134);
and U3205 (N_3205,N_3037,N_3118);
or U3206 (N_3206,N_3193,N_3132);
and U3207 (N_3207,N_3044,N_3121);
and U3208 (N_3208,N_3135,N_3199);
or U3209 (N_3209,N_3053,N_3184);
or U3210 (N_3210,N_3196,N_3173);
xor U3211 (N_3211,N_3153,N_3047);
nand U3212 (N_3212,N_3106,N_3162);
nand U3213 (N_3213,N_3185,N_3151);
or U3214 (N_3214,N_3018,N_3086);
nand U3215 (N_3215,N_3058,N_3023);
or U3216 (N_3216,N_3051,N_3049);
and U3217 (N_3217,N_3048,N_3170);
or U3218 (N_3218,N_3103,N_3179);
and U3219 (N_3219,N_3001,N_3136);
and U3220 (N_3220,N_3138,N_3189);
or U3221 (N_3221,N_3091,N_3183);
nand U3222 (N_3222,N_3038,N_3120);
or U3223 (N_3223,N_3078,N_3181);
nand U3224 (N_3224,N_3039,N_3082);
nand U3225 (N_3225,N_3144,N_3169);
and U3226 (N_3226,N_3002,N_3122);
or U3227 (N_3227,N_3195,N_3129);
nand U3228 (N_3228,N_3137,N_3188);
or U3229 (N_3229,N_3064,N_3165);
and U3230 (N_3230,N_3073,N_3031);
nor U3231 (N_3231,N_3042,N_3081);
and U3232 (N_3232,N_3161,N_3066);
nor U3233 (N_3233,N_3030,N_3123);
or U3234 (N_3234,N_3168,N_3124);
nand U3235 (N_3235,N_3085,N_3145);
nand U3236 (N_3236,N_3128,N_3080);
nand U3237 (N_3237,N_3172,N_3154);
or U3238 (N_3238,N_3060,N_3034);
nor U3239 (N_3239,N_3140,N_3107);
or U3240 (N_3240,N_3067,N_3094);
or U3241 (N_3241,N_3027,N_3175);
or U3242 (N_3242,N_3004,N_3159);
nand U3243 (N_3243,N_3177,N_3005);
nor U3244 (N_3244,N_3055,N_3088);
nor U3245 (N_3245,N_3090,N_3156);
or U3246 (N_3246,N_3069,N_3087);
nor U3247 (N_3247,N_3160,N_3021);
nand U3248 (N_3248,N_3111,N_3167);
and U3249 (N_3249,N_3158,N_3074);
nand U3250 (N_3250,N_3041,N_3063);
and U3251 (N_3251,N_3016,N_3100);
or U3252 (N_3252,N_3155,N_3197);
nor U3253 (N_3253,N_3152,N_3065);
nand U3254 (N_3254,N_3119,N_3019);
nor U3255 (N_3255,N_3098,N_3007);
nor U3256 (N_3256,N_3083,N_3110);
xor U3257 (N_3257,N_3157,N_3089);
nor U3258 (N_3258,N_3130,N_3006);
or U3259 (N_3259,N_3149,N_3043);
nand U3260 (N_3260,N_3070,N_3000);
nor U3261 (N_3261,N_3187,N_3036);
xnor U3262 (N_3262,N_3024,N_3015);
or U3263 (N_3263,N_3046,N_3028);
or U3264 (N_3264,N_3020,N_3163);
and U3265 (N_3265,N_3126,N_3014);
xnor U3266 (N_3266,N_3109,N_3099);
nand U3267 (N_3267,N_3142,N_3025);
xor U3268 (N_3268,N_3191,N_3116);
and U3269 (N_3269,N_3139,N_3076);
or U3270 (N_3270,N_3166,N_3012);
or U3271 (N_3271,N_3104,N_3176);
and U3272 (N_3272,N_3054,N_3032);
xnor U3273 (N_3273,N_3117,N_3071);
or U3274 (N_3274,N_3057,N_3131);
and U3275 (N_3275,N_3148,N_3035);
or U3276 (N_3276,N_3033,N_3198);
and U3277 (N_3277,N_3061,N_3125);
xor U3278 (N_3278,N_3072,N_3097);
and U3279 (N_3279,N_3127,N_3174);
xnor U3280 (N_3280,N_3075,N_3052);
xnor U3281 (N_3281,N_3192,N_3133);
nor U3282 (N_3282,N_3147,N_3102);
or U3283 (N_3283,N_3026,N_3114);
nand U3284 (N_3284,N_3077,N_3029);
or U3285 (N_3285,N_3079,N_3186);
nor U3286 (N_3286,N_3143,N_3050);
xnor U3287 (N_3287,N_3056,N_3180);
nor U3288 (N_3288,N_3095,N_3040);
nor U3289 (N_3289,N_3096,N_3146);
or U3290 (N_3290,N_3150,N_3022);
and U3291 (N_3291,N_3059,N_3112);
nor U3292 (N_3292,N_3141,N_3011);
xor U3293 (N_3293,N_3008,N_3115);
or U3294 (N_3294,N_3068,N_3062);
nand U3295 (N_3295,N_3113,N_3190);
nand U3296 (N_3296,N_3101,N_3013);
xnor U3297 (N_3297,N_3010,N_3092);
or U3298 (N_3298,N_3171,N_3182);
and U3299 (N_3299,N_3084,N_3017);
nand U3300 (N_3300,N_3095,N_3054);
nor U3301 (N_3301,N_3094,N_3106);
and U3302 (N_3302,N_3106,N_3197);
xnor U3303 (N_3303,N_3013,N_3019);
and U3304 (N_3304,N_3131,N_3078);
and U3305 (N_3305,N_3009,N_3164);
nand U3306 (N_3306,N_3033,N_3015);
and U3307 (N_3307,N_3116,N_3136);
or U3308 (N_3308,N_3121,N_3150);
nor U3309 (N_3309,N_3030,N_3035);
nor U3310 (N_3310,N_3107,N_3113);
xor U3311 (N_3311,N_3083,N_3172);
xor U3312 (N_3312,N_3155,N_3165);
or U3313 (N_3313,N_3054,N_3171);
or U3314 (N_3314,N_3137,N_3182);
xnor U3315 (N_3315,N_3132,N_3098);
nand U3316 (N_3316,N_3157,N_3010);
and U3317 (N_3317,N_3073,N_3076);
and U3318 (N_3318,N_3174,N_3075);
and U3319 (N_3319,N_3034,N_3068);
nor U3320 (N_3320,N_3163,N_3151);
and U3321 (N_3321,N_3062,N_3084);
or U3322 (N_3322,N_3093,N_3145);
nand U3323 (N_3323,N_3151,N_3114);
and U3324 (N_3324,N_3138,N_3015);
and U3325 (N_3325,N_3078,N_3186);
and U3326 (N_3326,N_3146,N_3190);
and U3327 (N_3327,N_3047,N_3070);
and U3328 (N_3328,N_3060,N_3177);
xnor U3329 (N_3329,N_3164,N_3116);
nand U3330 (N_3330,N_3162,N_3177);
xor U3331 (N_3331,N_3112,N_3077);
nor U3332 (N_3332,N_3195,N_3150);
nand U3333 (N_3333,N_3018,N_3186);
or U3334 (N_3334,N_3149,N_3162);
nor U3335 (N_3335,N_3058,N_3053);
and U3336 (N_3336,N_3157,N_3027);
or U3337 (N_3337,N_3029,N_3031);
or U3338 (N_3338,N_3196,N_3138);
or U3339 (N_3339,N_3076,N_3054);
nor U3340 (N_3340,N_3114,N_3120);
or U3341 (N_3341,N_3102,N_3198);
or U3342 (N_3342,N_3007,N_3023);
xor U3343 (N_3343,N_3194,N_3161);
nand U3344 (N_3344,N_3127,N_3066);
or U3345 (N_3345,N_3114,N_3186);
nor U3346 (N_3346,N_3085,N_3053);
nor U3347 (N_3347,N_3019,N_3063);
or U3348 (N_3348,N_3152,N_3193);
and U3349 (N_3349,N_3132,N_3042);
nand U3350 (N_3350,N_3038,N_3009);
nor U3351 (N_3351,N_3095,N_3069);
and U3352 (N_3352,N_3107,N_3136);
xnor U3353 (N_3353,N_3023,N_3151);
and U3354 (N_3354,N_3142,N_3161);
nor U3355 (N_3355,N_3058,N_3143);
nand U3356 (N_3356,N_3033,N_3102);
nand U3357 (N_3357,N_3061,N_3019);
nor U3358 (N_3358,N_3192,N_3116);
nor U3359 (N_3359,N_3037,N_3029);
nand U3360 (N_3360,N_3110,N_3011);
xor U3361 (N_3361,N_3192,N_3079);
nor U3362 (N_3362,N_3031,N_3196);
xor U3363 (N_3363,N_3035,N_3196);
nand U3364 (N_3364,N_3119,N_3069);
nand U3365 (N_3365,N_3007,N_3197);
and U3366 (N_3366,N_3138,N_3004);
and U3367 (N_3367,N_3078,N_3018);
nor U3368 (N_3368,N_3077,N_3086);
xor U3369 (N_3369,N_3036,N_3193);
or U3370 (N_3370,N_3172,N_3110);
nor U3371 (N_3371,N_3069,N_3015);
and U3372 (N_3372,N_3159,N_3178);
xor U3373 (N_3373,N_3027,N_3188);
nor U3374 (N_3374,N_3017,N_3135);
and U3375 (N_3375,N_3041,N_3032);
and U3376 (N_3376,N_3130,N_3166);
and U3377 (N_3377,N_3079,N_3092);
and U3378 (N_3378,N_3096,N_3081);
nor U3379 (N_3379,N_3008,N_3134);
or U3380 (N_3380,N_3121,N_3083);
and U3381 (N_3381,N_3119,N_3135);
nor U3382 (N_3382,N_3114,N_3116);
or U3383 (N_3383,N_3003,N_3022);
xnor U3384 (N_3384,N_3189,N_3016);
nor U3385 (N_3385,N_3126,N_3048);
and U3386 (N_3386,N_3196,N_3199);
or U3387 (N_3387,N_3188,N_3037);
xor U3388 (N_3388,N_3078,N_3061);
or U3389 (N_3389,N_3153,N_3193);
nor U3390 (N_3390,N_3137,N_3117);
nand U3391 (N_3391,N_3134,N_3060);
xor U3392 (N_3392,N_3131,N_3136);
and U3393 (N_3393,N_3024,N_3095);
and U3394 (N_3394,N_3134,N_3020);
nand U3395 (N_3395,N_3128,N_3123);
nand U3396 (N_3396,N_3158,N_3076);
nand U3397 (N_3397,N_3075,N_3051);
and U3398 (N_3398,N_3006,N_3062);
nand U3399 (N_3399,N_3139,N_3038);
nand U3400 (N_3400,N_3274,N_3263);
or U3401 (N_3401,N_3376,N_3244);
and U3402 (N_3402,N_3314,N_3207);
and U3403 (N_3403,N_3239,N_3371);
or U3404 (N_3404,N_3321,N_3227);
nand U3405 (N_3405,N_3323,N_3238);
xnor U3406 (N_3406,N_3335,N_3330);
and U3407 (N_3407,N_3324,N_3295);
and U3408 (N_3408,N_3357,N_3273);
and U3409 (N_3409,N_3206,N_3232);
and U3410 (N_3410,N_3287,N_3364);
and U3411 (N_3411,N_3299,N_3278);
and U3412 (N_3412,N_3215,N_3396);
nand U3413 (N_3413,N_3200,N_3248);
and U3414 (N_3414,N_3212,N_3270);
or U3415 (N_3415,N_3265,N_3208);
nand U3416 (N_3416,N_3289,N_3288);
or U3417 (N_3417,N_3285,N_3202);
xnor U3418 (N_3418,N_3241,N_3332);
nor U3419 (N_3419,N_3333,N_3219);
nand U3420 (N_3420,N_3290,N_3392);
and U3421 (N_3421,N_3268,N_3217);
nor U3422 (N_3422,N_3224,N_3379);
nor U3423 (N_3423,N_3228,N_3283);
nor U3424 (N_3424,N_3384,N_3251);
nor U3425 (N_3425,N_3372,N_3351);
and U3426 (N_3426,N_3308,N_3218);
nand U3427 (N_3427,N_3209,N_3349);
nor U3428 (N_3428,N_3210,N_3368);
xnor U3429 (N_3429,N_3306,N_3353);
xor U3430 (N_3430,N_3380,N_3394);
xnor U3431 (N_3431,N_3229,N_3373);
and U3432 (N_3432,N_3375,N_3214);
xor U3433 (N_3433,N_3340,N_3231);
and U3434 (N_3434,N_3301,N_3267);
nor U3435 (N_3435,N_3261,N_3316);
xnor U3436 (N_3436,N_3362,N_3203);
and U3437 (N_3437,N_3284,N_3225);
xnor U3438 (N_3438,N_3370,N_3281);
and U3439 (N_3439,N_3211,N_3243);
or U3440 (N_3440,N_3302,N_3319);
xor U3441 (N_3441,N_3226,N_3264);
or U3442 (N_3442,N_3390,N_3360);
or U3443 (N_3443,N_3275,N_3240);
or U3444 (N_3444,N_3237,N_3358);
or U3445 (N_3445,N_3297,N_3234);
xnor U3446 (N_3446,N_3338,N_3369);
and U3447 (N_3447,N_3205,N_3236);
and U3448 (N_3448,N_3391,N_3255);
and U3449 (N_3449,N_3242,N_3397);
or U3450 (N_3450,N_3307,N_3359);
nand U3451 (N_3451,N_3387,N_3339);
and U3452 (N_3452,N_3266,N_3317);
xor U3453 (N_3453,N_3367,N_3309);
xor U3454 (N_3454,N_3343,N_3253);
nand U3455 (N_3455,N_3250,N_3336);
and U3456 (N_3456,N_3366,N_3328);
nor U3457 (N_3457,N_3318,N_3213);
xnor U3458 (N_3458,N_3262,N_3386);
nand U3459 (N_3459,N_3320,N_3277);
and U3460 (N_3460,N_3310,N_3259);
and U3461 (N_3461,N_3395,N_3389);
xnor U3462 (N_3462,N_3279,N_3216);
nand U3463 (N_3463,N_3235,N_3280);
xor U3464 (N_3464,N_3325,N_3381);
nor U3465 (N_3465,N_3315,N_3254);
xnor U3466 (N_3466,N_3383,N_3233);
nand U3467 (N_3467,N_3377,N_3399);
nor U3468 (N_3468,N_3345,N_3342);
nor U3469 (N_3469,N_3303,N_3245);
xor U3470 (N_3470,N_3247,N_3293);
or U3471 (N_3471,N_3271,N_3322);
xor U3472 (N_3472,N_3292,N_3252);
xor U3473 (N_3473,N_3344,N_3346);
nor U3474 (N_3474,N_3222,N_3249);
nand U3475 (N_3475,N_3347,N_3365);
nand U3476 (N_3476,N_3223,N_3276);
and U3477 (N_3477,N_3327,N_3334);
nor U3478 (N_3478,N_3350,N_3286);
nand U3479 (N_3479,N_3313,N_3296);
or U3480 (N_3480,N_3221,N_3282);
or U3481 (N_3481,N_3388,N_3300);
and U3482 (N_3482,N_3348,N_3294);
and U3483 (N_3483,N_3374,N_3257);
xor U3484 (N_3484,N_3272,N_3291);
and U3485 (N_3485,N_3311,N_3260);
nor U3486 (N_3486,N_3378,N_3354);
or U3487 (N_3487,N_3312,N_3385);
or U3488 (N_3488,N_3355,N_3204);
xnor U3489 (N_3489,N_3398,N_3305);
or U3490 (N_3490,N_3352,N_3269);
and U3491 (N_3491,N_3382,N_3298);
and U3492 (N_3492,N_3361,N_3363);
xor U3493 (N_3493,N_3341,N_3326);
and U3494 (N_3494,N_3331,N_3220);
and U3495 (N_3495,N_3356,N_3258);
nor U3496 (N_3496,N_3304,N_3337);
nand U3497 (N_3497,N_3201,N_3230);
nor U3498 (N_3498,N_3393,N_3256);
nand U3499 (N_3499,N_3246,N_3329);
or U3500 (N_3500,N_3322,N_3224);
xnor U3501 (N_3501,N_3388,N_3326);
and U3502 (N_3502,N_3344,N_3236);
or U3503 (N_3503,N_3316,N_3326);
nand U3504 (N_3504,N_3212,N_3302);
nand U3505 (N_3505,N_3286,N_3357);
nand U3506 (N_3506,N_3216,N_3371);
xnor U3507 (N_3507,N_3235,N_3224);
nor U3508 (N_3508,N_3246,N_3273);
nor U3509 (N_3509,N_3380,N_3316);
or U3510 (N_3510,N_3370,N_3317);
xnor U3511 (N_3511,N_3278,N_3388);
or U3512 (N_3512,N_3344,N_3322);
and U3513 (N_3513,N_3369,N_3392);
or U3514 (N_3514,N_3250,N_3300);
nor U3515 (N_3515,N_3311,N_3375);
nand U3516 (N_3516,N_3394,N_3233);
nand U3517 (N_3517,N_3210,N_3209);
nand U3518 (N_3518,N_3238,N_3308);
xor U3519 (N_3519,N_3331,N_3390);
and U3520 (N_3520,N_3321,N_3271);
nor U3521 (N_3521,N_3392,N_3206);
and U3522 (N_3522,N_3380,N_3227);
and U3523 (N_3523,N_3336,N_3295);
nor U3524 (N_3524,N_3232,N_3356);
nand U3525 (N_3525,N_3392,N_3399);
nor U3526 (N_3526,N_3261,N_3395);
xor U3527 (N_3527,N_3287,N_3376);
or U3528 (N_3528,N_3375,N_3219);
or U3529 (N_3529,N_3378,N_3396);
nand U3530 (N_3530,N_3355,N_3337);
xor U3531 (N_3531,N_3388,N_3358);
nand U3532 (N_3532,N_3268,N_3319);
xnor U3533 (N_3533,N_3273,N_3209);
and U3534 (N_3534,N_3270,N_3289);
or U3535 (N_3535,N_3282,N_3242);
xnor U3536 (N_3536,N_3288,N_3331);
nand U3537 (N_3537,N_3257,N_3355);
and U3538 (N_3538,N_3241,N_3207);
xor U3539 (N_3539,N_3215,N_3245);
or U3540 (N_3540,N_3290,N_3309);
or U3541 (N_3541,N_3364,N_3301);
nor U3542 (N_3542,N_3219,N_3364);
nand U3543 (N_3543,N_3252,N_3336);
xor U3544 (N_3544,N_3344,N_3359);
nor U3545 (N_3545,N_3280,N_3312);
xnor U3546 (N_3546,N_3259,N_3372);
or U3547 (N_3547,N_3305,N_3211);
nand U3548 (N_3548,N_3271,N_3295);
and U3549 (N_3549,N_3335,N_3202);
nor U3550 (N_3550,N_3256,N_3218);
and U3551 (N_3551,N_3354,N_3219);
nand U3552 (N_3552,N_3256,N_3293);
or U3553 (N_3553,N_3258,N_3242);
or U3554 (N_3554,N_3396,N_3327);
and U3555 (N_3555,N_3358,N_3214);
nand U3556 (N_3556,N_3395,N_3258);
nor U3557 (N_3557,N_3235,N_3249);
and U3558 (N_3558,N_3373,N_3318);
nand U3559 (N_3559,N_3280,N_3291);
nand U3560 (N_3560,N_3317,N_3250);
and U3561 (N_3561,N_3366,N_3354);
or U3562 (N_3562,N_3246,N_3356);
and U3563 (N_3563,N_3313,N_3255);
and U3564 (N_3564,N_3236,N_3308);
and U3565 (N_3565,N_3329,N_3342);
nand U3566 (N_3566,N_3348,N_3303);
or U3567 (N_3567,N_3326,N_3343);
nor U3568 (N_3568,N_3305,N_3243);
nor U3569 (N_3569,N_3208,N_3259);
nand U3570 (N_3570,N_3272,N_3203);
or U3571 (N_3571,N_3230,N_3329);
nor U3572 (N_3572,N_3381,N_3289);
nand U3573 (N_3573,N_3392,N_3242);
nor U3574 (N_3574,N_3275,N_3229);
nand U3575 (N_3575,N_3389,N_3367);
or U3576 (N_3576,N_3248,N_3357);
and U3577 (N_3577,N_3253,N_3226);
xor U3578 (N_3578,N_3272,N_3221);
xnor U3579 (N_3579,N_3329,N_3275);
nor U3580 (N_3580,N_3329,N_3220);
and U3581 (N_3581,N_3334,N_3383);
or U3582 (N_3582,N_3315,N_3277);
nor U3583 (N_3583,N_3256,N_3274);
and U3584 (N_3584,N_3399,N_3366);
and U3585 (N_3585,N_3285,N_3234);
xnor U3586 (N_3586,N_3288,N_3306);
nor U3587 (N_3587,N_3348,N_3364);
and U3588 (N_3588,N_3205,N_3266);
nor U3589 (N_3589,N_3216,N_3229);
nand U3590 (N_3590,N_3210,N_3337);
and U3591 (N_3591,N_3384,N_3296);
and U3592 (N_3592,N_3228,N_3399);
or U3593 (N_3593,N_3316,N_3343);
and U3594 (N_3594,N_3282,N_3210);
or U3595 (N_3595,N_3288,N_3360);
or U3596 (N_3596,N_3288,N_3247);
xnor U3597 (N_3597,N_3205,N_3256);
xnor U3598 (N_3598,N_3243,N_3387);
and U3599 (N_3599,N_3247,N_3336);
nor U3600 (N_3600,N_3407,N_3509);
or U3601 (N_3601,N_3544,N_3537);
nand U3602 (N_3602,N_3543,N_3538);
or U3603 (N_3603,N_3476,N_3501);
nor U3604 (N_3604,N_3595,N_3448);
nor U3605 (N_3605,N_3415,N_3529);
xor U3606 (N_3606,N_3459,N_3508);
xnor U3607 (N_3607,N_3436,N_3488);
or U3608 (N_3608,N_3457,N_3539);
or U3609 (N_3609,N_3556,N_3572);
nor U3610 (N_3610,N_3551,N_3548);
or U3611 (N_3611,N_3433,N_3525);
and U3612 (N_3612,N_3587,N_3568);
or U3613 (N_3613,N_3541,N_3571);
xor U3614 (N_3614,N_3413,N_3427);
and U3615 (N_3615,N_3560,N_3493);
and U3616 (N_3616,N_3513,N_3514);
and U3617 (N_3617,N_3434,N_3507);
xnor U3618 (N_3618,N_3497,N_3517);
or U3619 (N_3619,N_3582,N_3515);
or U3620 (N_3620,N_3406,N_3449);
xor U3621 (N_3621,N_3502,N_3404);
nor U3622 (N_3622,N_3504,N_3467);
nand U3623 (N_3623,N_3416,N_3536);
nand U3624 (N_3624,N_3482,N_3461);
nand U3625 (N_3625,N_3424,N_3518);
nand U3626 (N_3626,N_3534,N_3565);
or U3627 (N_3627,N_3439,N_3462);
xnor U3628 (N_3628,N_3589,N_3567);
and U3629 (N_3629,N_3522,N_3435);
nor U3630 (N_3630,N_3426,N_3599);
nand U3631 (N_3631,N_3473,N_3574);
or U3632 (N_3632,N_3447,N_3440);
nor U3633 (N_3633,N_3466,N_3414);
xor U3634 (N_3634,N_3546,N_3532);
nor U3635 (N_3635,N_3499,N_3437);
and U3636 (N_3636,N_3512,N_3429);
or U3637 (N_3637,N_3455,N_3550);
nor U3638 (N_3638,N_3533,N_3422);
nand U3639 (N_3639,N_3510,N_3495);
or U3640 (N_3640,N_3483,N_3490);
nand U3641 (N_3641,N_3446,N_3477);
and U3642 (N_3642,N_3552,N_3549);
nand U3643 (N_3643,N_3594,N_3472);
or U3644 (N_3644,N_3484,N_3478);
and U3645 (N_3645,N_3516,N_3580);
and U3646 (N_3646,N_3593,N_3419);
xor U3647 (N_3647,N_3405,N_3445);
nor U3648 (N_3648,N_3475,N_3485);
nand U3649 (N_3649,N_3469,N_3425);
nor U3650 (N_3650,N_3530,N_3468);
nor U3651 (N_3651,N_3470,N_3418);
xor U3652 (N_3652,N_3591,N_3566);
nand U3653 (N_3653,N_3463,N_3590);
or U3654 (N_3654,N_3500,N_3431);
and U3655 (N_3655,N_3442,N_3526);
or U3656 (N_3656,N_3401,N_3527);
nor U3657 (N_3657,N_3400,N_3519);
nor U3658 (N_3658,N_3402,N_3581);
xnor U3659 (N_3659,N_3464,N_3570);
or U3660 (N_3660,N_3487,N_3553);
or U3661 (N_3661,N_3411,N_3576);
and U3662 (N_3662,N_3573,N_3443);
and U3663 (N_3663,N_3496,N_3597);
and U3664 (N_3664,N_3535,N_3506);
or U3665 (N_3665,N_3524,N_3410);
and U3666 (N_3666,N_3521,N_3554);
and U3667 (N_3667,N_3489,N_3454);
xor U3668 (N_3668,N_3491,N_3555);
xor U3669 (N_3669,N_3444,N_3585);
nand U3670 (N_3670,N_3481,N_3430);
xnor U3671 (N_3671,N_3438,N_3465);
xor U3672 (N_3672,N_3421,N_3575);
or U3673 (N_3673,N_3562,N_3456);
or U3674 (N_3674,N_3417,N_3586);
xnor U3675 (N_3675,N_3460,N_3531);
or U3676 (N_3676,N_3540,N_3561);
or U3677 (N_3677,N_3583,N_3494);
or U3678 (N_3678,N_3584,N_3598);
or U3679 (N_3679,N_3432,N_3428);
or U3680 (N_3680,N_3420,N_3503);
and U3681 (N_3681,N_3505,N_3403);
and U3682 (N_3682,N_3545,N_3579);
nor U3683 (N_3683,N_3588,N_3577);
or U3684 (N_3684,N_3450,N_3523);
nand U3685 (N_3685,N_3486,N_3451);
and U3686 (N_3686,N_3596,N_3564);
nor U3687 (N_3687,N_3458,N_3441);
nor U3688 (N_3688,N_3511,N_3592);
or U3689 (N_3689,N_3409,N_3412);
or U3690 (N_3690,N_3558,N_3408);
xnor U3691 (N_3691,N_3578,N_3542);
or U3692 (N_3692,N_3520,N_3569);
nand U3693 (N_3693,N_3480,N_3547);
and U3694 (N_3694,N_3453,N_3498);
nand U3695 (N_3695,N_3452,N_3479);
nand U3696 (N_3696,N_3528,N_3563);
nand U3697 (N_3697,N_3474,N_3423);
xor U3698 (N_3698,N_3559,N_3557);
nand U3699 (N_3699,N_3492,N_3471);
nand U3700 (N_3700,N_3591,N_3581);
or U3701 (N_3701,N_3502,N_3580);
and U3702 (N_3702,N_3417,N_3505);
and U3703 (N_3703,N_3412,N_3594);
xor U3704 (N_3704,N_3562,N_3512);
xor U3705 (N_3705,N_3402,N_3468);
nor U3706 (N_3706,N_3555,N_3594);
xnor U3707 (N_3707,N_3538,N_3422);
nand U3708 (N_3708,N_3473,N_3550);
nand U3709 (N_3709,N_3506,N_3561);
and U3710 (N_3710,N_3502,N_3457);
xnor U3711 (N_3711,N_3577,N_3531);
nor U3712 (N_3712,N_3530,N_3439);
nor U3713 (N_3713,N_3410,N_3500);
xor U3714 (N_3714,N_3512,N_3568);
nand U3715 (N_3715,N_3520,N_3460);
or U3716 (N_3716,N_3427,N_3486);
nor U3717 (N_3717,N_3561,N_3441);
and U3718 (N_3718,N_3598,N_3519);
or U3719 (N_3719,N_3465,N_3522);
or U3720 (N_3720,N_3599,N_3455);
and U3721 (N_3721,N_3539,N_3597);
nand U3722 (N_3722,N_3549,N_3499);
and U3723 (N_3723,N_3569,N_3414);
or U3724 (N_3724,N_3400,N_3564);
nor U3725 (N_3725,N_3518,N_3469);
nand U3726 (N_3726,N_3416,N_3401);
nand U3727 (N_3727,N_3501,N_3432);
and U3728 (N_3728,N_3594,N_3480);
xnor U3729 (N_3729,N_3543,N_3530);
nand U3730 (N_3730,N_3495,N_3577);
nand U3731 (N_3731,N_3498,N_3597);
xor U3732 (N_3732,N_3567,N_3565);
and U3733 (N_3733,N_3479,N_3465);
nor U3734 (N_3734,N_3558,N_3564);
xor U3735 (N_3735,N_3570,N_3449);
and U3736 (N_3736,N_3487,N_3409);
nand U3737 (N_3737,N_3558,N_3436);
xor U3738 (N_3738,N_3494,N_3501);
xor U3739 (N_3739,N_3437,N_3544);
nand U3740 (N_3740,N_3418,N_3431);
and U3741 (N_3741,N_3402,N_3575);
nor U3742 (N_3742,N_3521,N_3450);
nand U3743 (N_3743,N_3409,N_3456);
xor U3744 (N_3744,N_3505,N_3466);
nor U3745 (N_3745,N_3412,N_3593);
nor U3746 (N_3746,N_3469,N_3411);
or U3747 (N_3747,N_3588,N_3407);
or U3748 (N_3748,N_3561,N_3452);
or U3749 (N_3749,N_3481,N_3505);
nand U3750 (N_3750,N_3531,N_3526);
nor U3751 (N_3751,N_3527,N_3515);
and U3752 (N_3752,N_3406,N_3490);
nor U3753 (N_3753,N_3486,N_3433);
or U3754 (N_3754,N_3484,N_3526);
nor U3755 (N_3755,N_3575,N_3471);
or U3756 (N_3756,N_3458,N_3560);
nand U3757 (N_3757,N_3496,N_3538);
xor U3758 (N_3758,N_3424,N_3458);
nand U3759 (N_3759,N_3496,N_3553);
and U3760 (N_3760,N_3411,N_3539);
nor U3761 (N_3761,N_3544,N_3454);
nand U3762 (N_3762,N_3531,N_3521);
nand U3763 (N_3763,N_3405,N_3429);
and U3764 (N_3764,N_3434,N_3492);
or U3765 (N_3765,N_3535,N_3456);
and U3766 (N_3766,N_3520,N_3512);
xnor U3767 (N_3767,N_3506,N_3510);
nor U3768 (N_3768,N_3429,N_3511);
nand U3769 (N_3769,N_3577,N_3500);
nand U3770 (N_3770,N_3510,N_3431);
nor U3771 (N_3771,N_3565,N_3429);
and U3772 (N_3772,N_3475,N_3564);
xnor U3773 (N_3773,N_3404,N_3428);
nand U3774 (N_3774,N_3589,N_3524);
nand U3775 (N_3775,N_3556,N_3597);
nand U3776 (N_3776,N_3413,N_3524);
nand U3777 (N_3777,N_3479,N_3493);
nand U3778 (N_3778,N_3406,N_3443);
and U3779 (N_3779,N_3574,N_3483);
or U3780 (N_3780,N_3590,N_3428);
xnor U3781 (N_3781,N_3474,N_3462);
and U3782 (N_3782,N_3525,N_3409);
nand U3783 (N_3783,N_3426,N_3536);
or U3784 (N_3784,N_3527,N_3526);
nor U3785 (N_3785,N_3498,N_3584);
nor U3786 (N_3786,N_3521,N_3401);
or U3787 (N_3787,N_3475,N_3546);
nand U3788 (N_3788,N_3529,N_3515);
or U3789 (N_3789,N_3458,N_3535);
or U3790 (N_3790,N_3407,N_3508);
nor U3791 (N_3791,N_3574,N_3443);
or U3792 (N_3792,N_3507,N_3427);
nor U3793 (N_3793,N_3441,N_3588);
xnor U3794 (N_3794,N_3497,N_3475);
and U3795 (N_3795,N_3519,N_3548);
nand U3796 (N_3796,N_3505,N_3452);
nand U3797 (N_3797,N_3406,N_3558);
xor U3798 (N_3798,N_3469,N_3439);
nand U3799 (N_3799,N_3534,N_3539);
or U3800 (N_3800,N_3656,N_3634);
xor U3801 (N_3801,N_3689,N_3643);
nand U3802 (N_3802,N_3792,N_3706);
and U3803 (N_3803,N_3758,N_3767);
xnor U3804 (N_3804,N_3737,N_3623);
xnor U3805 (N_3805,N_3764,N_3785);
and U3806 (N_3806,N_3672,N_3644);
and U3807 (N_3807,N_3715,N_3621);
and U3808 (N_3808,N_3647,N_3695);
nand U3809 (N_3809,N_3771,N_3744);
xor U3810 (N_3810,N_3603,N_3633);
and U3811 (N_3811,N_3654,N_3752);
nand U3812 (N_3812,N_3684,N_3775);
and U3813 (N_3813,N_3607,N_3657);
nor U3814 (N_3814,N_3671,N_3754);
xor U3815 (N_3815,N_3739,N_3734);
or U3816 (N_3816,N_3681,N_3743);
xnor U3817 (N_3817,N_3702,N_3719);
xnor U3818 (N_3818,N_3777,N_3664);
or U3819 (N_3819,N_3655,N_3738);
xor U3820 (N_3820,N_3641,N_3658);
and U3821 (N_3821,N_3604,N_3600);
nand U3822 (N_3822,N_3776,N_3690);
or U3823 (N_3823,N_3778,N_3617);
xnor U3824 (N_3824,N_3700,N_3760);
nand U3825 (N_3825,N_3781,N_3619);
nor U3826 (N_3826,N_3769,N_3653);
and U3827 (N_3827,N_3756,N_3768);
and U3828 (N_3828,N_3707,N_3665);
and U3829 (N_3829,N_3708,N_3786);
xor U3830 (N_3830,N_3753,N_3787);
nor U3831 (N_3831,N_3799,N_3703);
nand U3832 (N_3832,N_3635,N_3774);
or U3833 (N_3833,N_3659,N_3608);
or U3834 (N_3834,N_3729,N_3639);
nand U3835 (N_3835,N_3615,N_3627);
nand U3836 (N_3836,N_3782,N_3742);
and U3837 (N_3837,N_3735,N_3755);
nand U3838 (N_3838,N_3685,N_3745);
nor U3839 (N_3839,N_3788,N_3796);
xnor U3840 (N_3840,N_3687,N_3676);
and U3841 (N_3841,N_3646,N_3736);
xor U3842 (N_3842,N_3610,N_3730);
and U3843 (N_3843,N_3698,N_3747);
xnor U3844 (N_3844,N_3688,N_3605);
nand U3845 (N_3845,N_3749,N_3670);
nand U3846 (N_3846,N_3650,N_3773);
or U3847 (N_3847,N_3631,N_3795);
xnor U3848 (N_3848,N_3667,N_3616);
nor U3849 (N_3849,N_3678,N_3725);
and U3850 (N_3850,N_3682,N_3630);
xor U3851 (N_3851,N_3668,N_3618);
or U3852 (N_3852,N_3704,N_3772);
nand U3853 (N_3853,N_3728,N_3640);
nand U3854 (N_3854,N_3709,N_3762);
nand U3855 (N_3855,N_3716,N_3660);
nand U3856 (N_3856,N_3666,N_3691);
or U3857 (N_3857,N_3696,N_3675);
nor U3858 (N_3858,N_3770,N_3727);
and U3859 (N_3859,N_3751,N_3759);
nand U3860 (N_3860,N_3711,N_3601);
nor U3861 (N_3861,N_3705,N_3726);
xor U3862 (N_3862,N_3680,N_3780);
nand U3863 (N_3863,N_3732,N_3779);
xnor U3864 (N_3864,N_3740,N_3720);
nand U3865 (N_3865,N_3645,N_3602);
nand U3866 (N_3866,N_3789,N_3798);
nor U3867 (N_3867,N_3710,N_3750);
nand U3868 (N_3868,N_3648,N_3636);
nor U3869 (N_3869,N_3613,N_3614);
nor U3870 (N_3870,N_3761,N_3797);
nand U3871 (N_3871,N_3637,N_3626);
or U3872 (N_3872,N_3638,N_3692);
nand U3873 (N_3873,N_3733,N_3784);
nand U3874 (N_3874,N_3662,N_3790);
nor U3875 (N_3875,N_3632,N_3679);
xnor U3876 (N_3876,N_3628,N_3699);
nand U3877 (N_3877,N_3629,N_3746);
or U3878 (N_3878,N_3765,N_3712);
xor U3879 (N_3879,N_3794,N_3713);
nor U3880 (N_3880,N_3741,N_3693);
nor U3881 (N_3881,N_3661,N_3694);
nor U3882 (N_3882,N_3717,N_3731);
nand U3883 (N_3883,N_3674,N_3757);
xnor U3884 (N_3884,N_3609,N_3651);
and U3885 (N_3885,N_3721,N_3763);
nor U3886 (N_3886,N_3697,N_3783);
nor U3887 (N_3887,N_3611,N_3723);
and U3888 (N_3888,N_3724,N_3625);
and U3889 (N_3889,N_3606,N_3701);
or U3890 (N_3890,N_3683,N_3722);
and U3891 (N_3891,N_3649,N_3620);
xor U3892 (N_3892,N_3686,N_3677);
and U3893 (N_3893,N_3624,N_3718);
and U3894 (N_3894,N_3673,N_3793);
nand U3895 (N_3895,N_3612,N_3766);
or U3896 (N_3896,N_3642,N_3652);
or U3897 (N_3897,N_3791,N_3714);
and U3898 (N_3898,N_3622,N_3663);
nor U3899 (N_3899,N_3748,N_3669);
xnor U3900 (N_3900,N_3690,N_3689);
and U3901 (N_3901,N_3726,N_3715);
or U3902 (N_3902,N_3734,N_3748);
nor U3903 (N_3903,N_3612,N_3736);
and U3904 (N_3904,N_3701,N_3667);
nor U3905 (N_3905,N_3687,N_3764);
and U3906 (N_3906,N_3759,N_3654);
or U3907 (N_3907,N_3787,N_3635);
and U3908 (N_3908,N_3689,N_3744);
xnor U3909 (N_3909,N_3653,N_3622);
nor U3910 (N_3910,N_3718,N_3724);
nor U3911 (N_3911,N_3786,N_3718);
or U3912 (N_3912,N_3796,N_3608);
nor U3913 (N_3913,N_3770,N_3762);
nand U3914 (N_3914,N_3748,N_3690);
nand U3915 (N_3915,N_3679,N_3688);
or U3916 (N_3916,N_3652,N_3723);
nand U3917 (N_3917,N_3791,N_3663);
and U3918 (N_3918,N_3779,N_3640);
and U3919 (N_3919,N_3643,N_3735);
or U3920 (N_3920,N_3743,N_3688);
nor U3921 (N_3921,N_3668,N_3692);
nor U3922 (N_3922,N_3763,N_3638);
nor U3923 (N_3923,N_3766,N_3675);
or U3924 (N_3924,N_3693,N_3672);
nand U3925 (N_3925,N_3620,N_3739);
nand U3926 (N_3926,N_3797,N_3772);
xnor U3927 (N_3927,N_3603,N_3743);
or U3928 (N_3928,N_3716,N_3659);
nand U3929 (N_3929,N_3741,N_3770);
nand U3930 (N_3930,N_3700,N_3666);
nand U3931 (N_3931,N_3797,N_3686);
xnor U3932 (N_3932,N_3641,N_3711);
nand U3933 (N_3933,N_3693,N_3774);
or U3934 (N_3934,N_3775,N_3761);
xnor U3935 (N_3935,N_3756,N_3662);
xor U3936 (N_3936,N_3672,N_3665);
nand U3937 (N_3937,N_3764,N_3732);
nor U3938 (N_3938,N_3678,N_3787);
or U3939 (N_3939,N_3791,N_3679);
and U3940 (N_3940,N_3660,N_3620);
or U3941 (N_3941,N_3776,N_3682);
nor U3942 (N_3942,N_3616,N_3780);
nand U3943 (N_3943,N_3675,N_3719);
nand U3944 (N_3944,N_3713,N_3654);
and U3945 (N_3945,N_3687,N_3717);
or U3946 (N_3946,N_3607,N_3616);
and U3947 (N_3947,N_3695,N_3702);
xor U3948 (N_3948,N_3799,N_3626);
or U3949 (N_3949,N_3710,N_3672);
xor U3950 (N_3950,N_3703,N_3732);
or U3951 (N_3951,N_3712,N_3689);
or U3952 (N_3952,N_3711,N_3666);
nand U3953 (N_3953,N_3746,N_3741);
or U3954 (N_3954,N_3675,N_3736);
nor U3955 (N_3955,N_3716,N_3617);
nor U3956 (N_3956,N_3696,N_3615);
xnor U3957 (N_3957,N_3634,N_3780);
and U3958 (N_3958,N_3782,N_3696);
and U3959 (N_3959,N_3791,N_3731);
and U3960 (N_3960,N_3775,N_3694);
nor U3961 (N_3961,N_3604,N_3696);
or U3962 (N_3962,N_3767,N_3618);
nor U3963 (N_3963,N_3796,N_3721);
or U3964 (N_3964,N_3693,N_3637);
nand U3965 (N_3965,N_3705,N_3617);
or U3966 (N_3966,N_3696,N_3673);
nor U3967 (N_3967,N_3747,N_3767);
and U3968 (N_3968,N_3642,N_3760);
xor U3969 (N_3969,N_3641,N_3746);
or U3970 (N_3970,N_3662,N_3744);
nor U3971 (N_3971,N_3795,N_3661);
nor U3972 (N_3972,N_3710,N_3689);
xor U3973 (N_3973,N_3791,N_3684);
and U3974 (N_3974,N_3797,N_3709);
or U3975 (N_3975,N_3743,N_3748);
nand U3976 (N_3976,N_3696,N_3662);
and U3977 (N_3977,N_3764,N_3714);
nand U3978 (N_3978,N_3600,N_3702);
nand U3979 (N_3979,N_3657,N_3755);
or U3980 (N_3980,N_3668,N_3746);
and U3981 (N_3981,N_3627,N_3600);
and U3982 (N_3982,N_3625,N_3623);
or U3983 (N_3983,N_3765,N_3721);
nand U3984 (N_3984,N_3670,N_3726);
or U3985 (N_3985,N_3606,N_3627);
and U3986 (N_3986,N_3778,N_3793);
nor U3987 (N_3987,N_3697,N_3636);
or U3988 (N_3988,N_3793,N_3776);
nand U3989 (N_3989,N_3649,N_3799);
and U3990 (N_3990,N_3750,N_3766);
and U3991 (N_3991,N_3603,N_3788);
and U3992 (N_3992,N_3742,N_3656);
xnor U3993 (N_3993,N_3670,N_3648);
nor U3994 (N_3994,N_3667,N_3753);
or U3995 (N_3995,N_3753,N_3642);
xor U3996 (N_3996,N_3777,N_3659);
xor U3997 (N_3997,N_3630,N_3608);
nor U3998 (N_3998,N_3600,N_3773);
and U3999 (N_3999,N_3646,N_3744);
xor U4000 (N_4000,N_3804,N_3916);
nor U4001 (N_4001,N_3933,N_3929);
xnor U4002 (N_4002,N_3802,N_3858);
and U4003 (N_4003,N_3866,N_3835);
or U4004 (N_4004,N_3880,N_3811);
or U4005 (N_4005,N_3831,N_3986);
nor U4006 (N_4006,N_3870,N_3926);
xnor U4007 (N_4007,N_3989,N_3907);
nand U4008 (N_4008,N_3894,N_3867);
nor U4009 (N_4009,N_3936,N_3879);
nor U4010 (N_4010,N_3853,N_3959);
and U4011 (N_4011,N_3851,N_3854);
nor U4012 (N_4012,N_3843,N_3940);
nor U4013 (N_4013,N_3817,N_3924);
or U4014 (N_4014,N_3998,N_3984);
nand U4015 (N_4015,N_3850,N_3948);
and U4016 (N_4016,N_3969,N_3946);
or U4017 (N_4017,N_3859,N_3912);
nor U4018 (N_4018,N_3938,N_3947);
and U4019 (N_4019,N_3857,N_3905);
xnor U4020 (N_4020,N_3820,N_3801);
or U4021 (N_4021,N_3836,N_3856);
xor U4022 (N_4022,N_3983,N_3960);
xnor U4023 (N_4023,N_3891,N_3895);
and U4024 (N_4024,N_3819,N_3808);
xor U4025 (N_4025,N_3980,N_3968);
nor U4026 (N_4026,N_3997,N_3963);
xnor U4027 (N_4027,N_3825,N_3848);
nor U4028 (N_4028,N_3944,N_3822);
xor U4029 (N_4029,N_3985,N_3945);
nor U4030 (N_4030,N_3846,N_3878);
nor U4031 (N_4031,N_3976,N_3821);
or U4032 (N_4032,N_3937,N_3809);
or U4033 (N_4033,N_3893,N_3996);
nor U4034 (N_4034,N_3807,N_3881);
nor U4035 (N_4035,N_3800,N_3877);
xor U4036 (N_4036,N_3885,N_3844);
and U4037 (N_4037,N_3932,N_3845);
or U4038 (N_4038,N_3823,N_3862);
nand U4039 (N_4039,N_3861,N_3864);
and U4040 (N_4040,N_3806,N_3826);
xor U4041 (N_4041,N_3832,N_3900);
nor U4042 (N_4042,N_3909,N_3955);
or U4043 (N_4043,N_3868,N_3952);
nor U4044 (N_4044,N_3888,N_3884);
and U4045 (N_4045,N_3896,N_3901);
nor U4046 (N_4046,N_3908,N_3911);
xnor U4047 (N_4047,N_3987,N_3816);
and U4048 (N_4048,N_3914,N_3965);
and U4049 (N_4049,N_3897,N_3957);
or U4050 (N_4050,N_3849,N_3935);
and U4051 (N_4051,N_3803,N_3824);
or U4052 (N_4052,N_3966,N_3991);
xnor U4053 (N_4053,N_3982,N_3814);
xnor U4054 (N_4054,N_3863,N_3918);
nand U4055 (N_4055,N_3889,N_3904);
nor U4056 (N_4056,N_3964,N_3978);
nand U4057 (N_4057,N_3913,N_3981);
and U4058 (N_4058,N_3842,N_3827);
nand U4059 (N_4059,N_3873,N_3812);
xor U4060 (N_4060,N_3830,N_3934);
xor U4061 (N_4061,N_3838,N_3869);
and U4062 (N_4062,N_3818,N_3833);
or U4063 (N_4063,N_3805,N_3990);
nor U4064 (N_4064,N_3974,N_3992);
and U4065 (N_4065,N_3883,N_3890);
or U4066 (N_4066,N_3910,N_3875);
or U4067 (N_4067,N_3923,N_3828);
xnor U4068 (N_4068,N_3829,N_3925);
or U4069 (N_4069,N_3915,N_3865);
nor U4070 (N_4070,N_3815,N_3951);
xnor U4071 (N_4071,N_3906,N_3837);
nand U4072 (N_4072,N_3872,N_3993);
nand U4073 (N_4073,N_3971,N_3973);
xnor U4074 (N_4074,N_3962,N_3942);
or U4075 (N_4075,N_3855,N_3961);
and U4076 (N_4076,N_3898,N_3922);
nand U4077 (N_4077,N_3921,N_3919);
nand U4078 (N_4078,N_3876,N_3954);
xnor U4079 (N_4079,N_3994,N_3852);
xor U4080 (N_4080,N_3886,N_3927);
and U4081 (N_4081,N_3917,N_3902);
and U4082 (N_4082,N_3999,N_3892);
xnor U4083 (N_4083,N_3958,N_3970);
xnor U4084 (N_4084,N_3871,N_3943);
xnor U4085 (N_4085,N_3956,N_3887);
nand U4086 (N_4086,N_3813,N_3928);
and U4087 (N_4087,N_3899,N_3841);
or U4088 (N_4088,N_3903,N_3874);
or U4089 (N_4089,N_3988,N_3975);
nor U4090 (N_4090,N_3840,N_3847);
nor U4091 (N_4091,N_3967,N_3930);
xnor U4092 (N_4092,N_3977,N_3972);
or U4093 (N_4093,N_3810,N_3941);
xnor U4094 (N_4094,N_3949,N_3979);
nor U4095 (N_4095,N_3839,N_3939);
or U4096 (N_4096,N_3953,N_3920);
xnor U4097 (N_4097,N_3995,N_3931);
nor U4098 (N_4098,N_3860,N_3882);
xnor U4099 (N_4099,N_3950,N_3834);
or U4100 (N_4100,N_3901,N_3839);
nor U4101 (N_4101,N_3889,N_3888);
and U4102 (N_4102,N_3801,N_3804);
xor U4103 (N_4103,N_3849,N_3827);
nor U4104 (N_4104,N_3956,N_3890);
nand U4105 (N_4105,N_3824,N_3841);
or U4106 (N_4106,N_3963,N_3882);
xnor U4107 (N_4107,N_3977,N_3853);
and U4108 (N_4108,N_3944,N_3810);
xnor U4109 (N_4109,N_3940,N_3870);
and U4110 (N_4110,N_3924,N_3894);
and U4111 (N_4111,N_3881,N_3941);
nor U4112 (N_4112,N_3874,N_3891);
nand U4113 (N_4113,N_3847,N_3809);
nor U4114 (N_4114,N_3951,N_3986);
xnor U4115 (N_4115,N_3981,N_3946);
nand U4116 (N_4116,N_3855,N_3978);
nand U4117 (N_4117,N_3851,N_3987);
or U4118 (N_4118,N_3908,N_3951);
and U4119 (N_4119,N_3988,N_3902);
nand U4120 (N_4120,N_3815,N_3945);
nand U4121 (N_4121,N_3905,N_3989);
nand U4122 (N_4122,N_3899,N_3829);
xnor U4123 (N_4123,N_3838,N_3820);
nor U4124 (N_4124,N_3939,N_3965);
nor U4125 (N_4125,N_3887,N_3833);
nor U4126 (N_4126,N_3851,N_3894);
xor U4127 (N_4127,N_3885,N_3895);
and U4128 (N_4128,N_3881,N_3954);
nor U4129 (N_4129,N_3860,N_3872);
or U4130 (N_4130,N_3802,N_3994);
nand U4131 (N_4131,N_3939,N_3914);
or U4132 (N_4132,N_3830,N_3839);
xnor U4133 (N_4133,N_3918,N_3964);
or U4134 (N_4134,N_3875,N_3839);
and U4135 (N_4135,N_3821,N_3823);
nor U4136 (N_4136,N_3816,N_3899);
xnor U4137 (N_4137,N_3863,N_3905);
nor U4138 (N_4138,N_3935,N_3889);
and U4139 (N_4139,N_3854,N_3874);
nand U4140 (N_4140,N_3932,N_3818);
or U4141 (N_4141,N_3895,N_3919);
nor U4142 (N_4142,N_3824,N_3933);
xnor U4143 (N_4143,N_3929,N_3808);
nand U4144 (N_4144,N_3890,N_3806);
xor U4145 (N_4145,N_3969,N_3859);
or U4146 (N_4146,N_3963,N_3976);
xor U4147 (N_4147,N_3923,N_3811);
xor U4148 (N_4148,N_3996,N_3942);
nor U4149 (N_4149,N_3982,N_3959);
and U4150 (N_4150,N_3894,N_3957);
nor U4151 (N_4151,N_3973,N_3837);
and U4152 (N_4152,N_3918,N_3853);
nand U4153 (N_4153,N_3861,N_3897);
nor U4154 (N_4154,N_3827,N_3847);
and U4155 (N_4155,N_3867,N_3821);
xor U4156 (N_4156,N_3889,N_3877);
xnor U4157 (N_4157,N_3965,N_3978);
or U4158 (N_4158,N_3891,N_3805);
nand U4159 (N_4159,N_3954,N_3978);
nand U4160 (N_4160,N_3922,N_3860);
and U4161 (N_4161,N_3886,N_3843);
nor U4162 (N_4162,N_3869,N_3991);
and U4163 (N_4163,N_3822,N_3974);
and U4164 (N_4164,N_3828,N_3846);
or U4165 (N_4165,N_3862,N_3987);
and U4166 (N_4166,N_3813,N_3916);
nand U4167 (N_4167,N_3815,N_3935);
xor U4168 (N_4168,N_3879,N_3811);
or U4169 (N_4169,N_3835,N_3904);
and U4170 (N_4170,N_3895,N_3813);
nor U4171 (N_4171,N_3882,N_3902);
and U4172 (N_4172,N_3801,N_3868);
or U4173 (N_4173,N_3898,N_3808);
nor U4174 (N_4174,N_3994,N_3833);
xor U4175 (N_4175,N_3876,N_3953);
nor U4176 (N_4176,N_3893,N_3970);
or U4177 (N_4177,N_3942,N_3886);
and U4178 (N_4178,N_3975,N_3848);
xnor U4179 (N_4179,N_3909,N_3959);
nor U4180 (N_4180,N_3895,N_3862);
and U4181 (N_4181,N_3928,N_3965);
or U4182 (N_4182,N_3917,N_3916);
and U4183 (N_4183,N_3994,N_3832);
xnor U4184 (N_4184,N_3999,N_3996);
xor U4185 (N_4185,N_3876,N_3830);
xor U4186 (N_4186,N_3965,N_3900);
xnor U4187 (N_4187,N_3977,N_3933);
and U4188 (N_4188,N_3975,N_3984);
xnor U4189 (N_4189,N_3829,N_3838);
or U4190 (N_4190,N_3846,N_3879);
nor U4191 (N_4191,N_3941,N_3908);
nor U4192 (N_4192,N_3949,N_3837);
xnor U4193 (N_4193,N_3939,N_3807);
nand U4194 (N_4194,N_3993,N_3855);
nor U4195 (N_4195,N_3953,N_3870);
nor U4196 (N_4196,N_3825,N_3865);
and U4197 (N_4197,N_3950,N_3880);
xor U4198 (N_4198,N_3979,N_3919);
xor U4199 (N_4199,N_3880,N_3878);
and U4200 (N_4200,N_4096,N_4030);
xnor U4201 (N_4201,N_4121,N_4001);
nand U4202 (N_4202,N_4159,N_4113);
and U4203 (N_4203,N_4125,N_4179);
and U4204 (N_4204,N_4077,N_4199);
nor U4205 (N_4205,N_4083,N_4136);
and U4206 (N_4206,N_4072,N_4186);
nor U4207 (N_4207,N_4092,N_4052);
or U4208 (N_4208,N_4173,N_4112);
and U4209 (N_4209,N_4016,N_4074);
or U4210 (N_4210,N_4032,N_4148);
and U4211 (N_4211,N_4114,N_4105);
or U4212 (N_4212,N_4007,N_4138);
xnor U4213 (N_4213,N_4165,N_4188);
xnor U4214 (N_4214,N_4005,N_4012);
or U4215 (N_4215,N_4055,N_4141);
and U4216 (N_4216,N_4118,N_4163);
and U4217 (N_4217,N_4107,N_4010);
xnor U4218 (N_4218,N_4004,N_4053);
nor U4219 (N_4219,N_4094,N_4154);
or U4220 (N_4220,N_4137,N_4026);
and U4221 (N_4221,N_4117,N_4189);
or U4222 (N_4222,N_4041,N_4031);
nor U4223 (N_4223,N_4106,N_4021);
xor U4224 (N_4224,N_4057,N_4102);
and U4225 (N_4225,N_4014,N_4069);
and U4226 (N_4226,N_4011,N_4143);
and U4227 (N_4227,N_4175,N_4192);
or U4228 (N_4228,N_4104,N_4139);
nor U4229 (N_4229,N_4101,N_4128);
nand U4230 (N_4230,N_4071,N_4049);
or U4231 (N_4231,N_4115,N_4028);
nand U4232 (N_4232,N_4065,N_4070);
or U4233 (N_4233,N_4079,N_4038);
or U4234 (N_4234,N_4171,N_4194);
or U4235 (N_4235,N_4034,N_4110);
and U4236 (N_4236,N_4044,N_4190);
and U4237 (N_4237,N_4039,N_4153);
nor U4238 (N_4238,N_4051,N_4178);
or U4239 (N_4239,N_4066,N_4095);
nand U4240 (N_4240,N_4149,N_4158);
nor U4241 (N_4241,N_4120,N_4098);
nand U4242 (N_4242,N_4081,N_4062);
xor U4243 (N_4243,N_4046,N_4119);
nor U4244 (N_4244,N_4111,N_4015);
nand U4245 (N_4245,N_4076,N_4078);
and U4246 (N_4246,N_4027,N_4135);
and U4247 (N_4247,N_4147,N_4142);
nand U4248 (N_4248,N_4090,N_4036);
nand U4249 (N_4249,N_4024,N_4129);
or U4250 (N_4250,N_4146,N_4187);
xor U4251 (N_4251,N_4182,N_4164);
or U4252 (N_4252,N_4020,N_4172);
nor U4253 (N_4253,N_4108,N_4093);
nor U4254 (N_4254,N_4048,N_4050);
nor U4255 (N_4255,N_4160,N_4167);
nor U4256 (N_4256,N_4124,N_4185);
or U4257 (N_4257,N_4029,N_4018);
and U4258 (N_4258,N_4183,N_4145);
nand U4259 (N_4259,N_4162,N_4045);
nand U4260 (N_4260,N_4195,N_4064);
xnor U4261 (N_4261,N_4009,N_4060);
xor U4262 (N_4262,N_4073,N_4123);
and U4263 (N_4263,N_4131,N_4127);
or U4264 (N_4264,N_4176,N_4130);
xor U4265 (N_4265,N_4084,N_4089);
and U4266 (N_4266,N_4035,N_4085);
nand U4267 (N_4267,N_4174,N_4099);
and U4268 (N_4268,N_4140,N_4097);
nor U4269 (N_4269,N_4109,N_4132);
nor U4270 (N_4270,N_4116,N_4122);
nand U4271 (N_4271,N_4144,N_4006);
and U4272 (N_4272,N_4042,N_4061);
nand U4273 (N_4273,N_4087,N_4100);
and U4274 (N_4274,N_4196,N_4040);
nand U4275 (N_4275,N_4082,N_4017);
or U4276 (N_4276,N_4067,N_4166);
nor U4277 (N_4277,N_4091,N_4181);
xor U4278 (N_4278,N_4059,N_4133);
or U4279 (N_4279,N_4033,N_4054);
xor U4280 (N_4280,N_4088,N_4169);
and U4281 (N_4281,N_4170,N_4086);
xnor U4282 (N_4282,N_4157,N_4156);
and U4283 (N_4283,N_4193,N_4063);
or U4284 (N_4284,N_4025,N_4013);
nor U4285 (N_4285,N_4019,N_4150);
or U4286 (N_4286,N_4056,N_4177);
and U4287 (N_4287,N_4184,N_4155);
xor U4288 (N_4288,N_4180,N_4080);
nor U4289 (N_4289,N_4152,N_4000);
xor U4290 (N_4290,N_4198,N_4008);
nand U4291 (N_4291,N_4068,N_4022);
and U4292 (N_4292,N_4191,N_4075);
nor U4293 (N_4293,N_4003,N_4126);
and U4294 (N_4294,N_4023,N_4058);
nor U4295 (N_4295,N_4037,N_4002);
nand U4296 (N_4296,N_4161,N_4043);
nand U4297 (N_4297,N_4103,N_4197);
and U4298 (N_4298,N_4047,N_4168);
nor U4299 (N_4299,N_4134,N_4151);
nor U4300 (N_4300,N_4060,N_4094);
nor U4301 (N_4301,N_4029,N_4151);
nand U4302 (N_4302,N_4169,N_4017);
xnor U4303 (N_4303,N_4092,N_4063);
xor U4304 (N_4304,N_4012,N_4146);
or U4305 (N_4305,N_4083,N_4138);
nor U4306 (N_4306,N_4190,N_4125);
or U4307 (N_4307,N_4086,N_4025);
nand U4308 (N_4308,N_4053,N_4060);
or U4309 (N_4309,N_4192,N_4120);
xnor U4310 (N_4310,N_4147,N_4031);
or U4311 (N_4311,N_4044,N_4110);
nand U4312 (N_4312,N_4099,N_4086);
xor U4313 (N_4313,N_4123,N_4011);
nor U4314 (N_4314,N_4161,N_4002);
nor U4315 (N_4315,N_4123,N_4100);
nor U4316 (N_4316,N_4184,N_4078);
nand U4317 (N_4317,N_4151,N_4020);
xnor U4318 (N_4318,N_4196,N_4170);
or U4319 (N_4319,N_4128,N_4172);
and U4320 (N_4320,N_4172,N_4131);
nand U4321 (N_4321,N_4178,N_4166);
xnor U4322 (N_4322,N_4066,N_4118);
xnor U4323 (N_4323,N_4188,N_4179);
nand U4324 (N_4324,N_4120,N_4024);
or U4325 (N_4325,N_4110,N_4188);
nor U4326 (N_4326,N_4160,N_4020);
nand U4327 (N_4327,N_4158,N_4045);
or U4328 (N_4328,N_4007,N_4024);
or U4329 (N_4329,N_4010,N_4109);
or U4330 (N_4330,N_4032,N_4142);
or U4331 (N_4331,N_4065,N_4066);
nand U4332 (N_4332,N_4196,N_4032);
nand U4333 (N_4333,N_4025,N_4134);
or U4334 (N_4334,N_4004,N_4142);
or U4335 (N_4335,N_4186,N_4122);
nor U4336 (N_4336,N_4172,N_4065);
nand U4337 (N_4337,N_4175,N_4190);
nand U4338 (N_4338,N_4036,N_4095);
and U4339 (N_4339,N_4051,N_4164);
or U4340 (N_4340,N_4014,N_4146);
nor U4341 (N_4341,N_4035,N_4173);
xnor U4342 (N_4342,N_4091,N_4094);
or U4343 (N_4343,N_4188,N_4017);
and U4344 (N_4344,N_4166,N_4103);
and U4345 (N_4345,N_4001,N_4175);
nand U4346 (N_4346,N_4035,N_4193);
and U4347 (N_4347,N_4040,N_4065);
and U4348 (N_4348,N_4140,N_4102);
xnor U4349 (N_4349,N_4056,N_4049);
nand U4350 (N_4350,N_4170,N_4030);
and U4351 (N_4351,N_4030,N_4135);
xnor U4352 (N_4352,N_4168,N_4071);
and U4353 (N_4353,N_4052,N_4018);
xnor U4354 (N_4354,N_4097,N_4191);
or U4355 (N_4355,N_4143,N_4167);
and U4356 (N_4356,N_4136,N_4198);
and U4357 (N_4357,N_4128,N_4091);
xnor U4358 (N_4358,N_4189,N_4139);
or U4359 (N_4359,N_4069,N_4090);
and U4360 (N_4360,N_4009,N_4143);
or U4361 (N_4361,N_4136,N_4172);
nand U4362 (N_4362,N_4051,N_4131);
xor U4363 (N_4363,N_4065,N_4121);
xnor U4364 (N_4364,N_4053,N_4129);
nor U4365 (N_4365,N_4127,N_4143);
and U4366 (N_4366,N_4157,N_4074);
nand U4367 (N_4367,N_4074,N_4104);
and U4368 (N_4368,N_4039,N_4085);
or U4369 (N_4369,N_4125,N_4063);
nand U4370 (N_4370,N_4172,N_4156);
nand U4371 (N_4371,N_4091,N_4025);
and U4372 (N_4372,N_4029,N_4062);
and U4373 (N_4373,N_4065,N_4123);
or U4374 (N_4374,N_4084,N_4188);
or U4375 (N_4375,N_4098,N_4009);
nor U4376 (N_4376,N_4037,N_4117);
xnor U4377 (N_4377,N_4132,N_4037);
nand U4378 (N_4378,N_4097,N_4037);
and U4379 (N_4379,N_4192,N_4064);
and U4380 (N_4380,N_4113,N_4111);
nor U4381 (N_4381,N_4157,N_4022);
or U4382 (N_4382,N_4193,N_4186);
and U4383 (N_4383,N_4194,N_4080);
nor U4384 (N_4384,N_4102,N_4059);
nor U4385 (N_4385,N_4167,N_4177);
nand U4386 (N_4386,N_4033,N_4082);
and U4387 (N_4387,N_4079,N_4034);
nor U4388 (N_4388,N_4092,N_4171);
and U4389 (N_4389,N_4182,N_4020);
xnor U4390 (N_4390,N_4029,N_4092);
nand U4391 (N_4391,N_4055,N_4044);
nand U4392 (N_4392,N_4162,N_4194);
xor U4393 (N_4393,N_4050,N_4068);
or U4394 (N_4394,N_4077,N_4010);
nor U4395 (N_4395,N_4083,N_4040);
and U4396 (N_4396,N_4190,N_4055);
xor U4397 (N_4397,N_4002,N_4009);
xor U4398 (N_4398,N_4082,N_4130);
or U4399 (N_4399,N_4004,N_4165);
nor U4400 (N_4400,N_4325,N_4327);
xor U4401 (N_4401,N_4243,N_4361);
nand U4402 (N_4402,N_4352,N_4349);
and U4403 (N_4403,N_4363,N_4256);
xor U4404 (N_4404,N_4278,N_4294);
nor U4405 (N_4405,N_4268,N_4380);
and U4406 (N_4406,N_4215,N_4379);
nor U4407 (N_4407,N_4290,N_4205);
or U4408 (N_4408,N_4329,N_4229);
xnor U4409 (N_4409,N_4200,N_4344);
and U4410 (N_4410,N_4399,N_4387);
or U4411 (N_4411,N_4252,N_4386);
nor U4412 (N_4412,N_4242,N_4259);
nand U4413 (N_4413,N_4223,N_4266);
xnor U4414 (N_4414,N_4355,N_4263);
nor U4415 (N_4415,N_4335,N_4336);
nand U4416 (N_4416,N_4322,N_4382);
or U4417 (N_4417,N_4241,N_4312);
or U4418 (N_4418,N_4232,N_4314);
xor U4419 (N_4419,N_4346,N_4244);
xor U4420 (N_4420,N_4230,N_4318);
and U4421 (N_4421,N_4393,N_4293);
nand U4422 (N_4422,N_4367,N_4370);
nand U4423 (N_4423,N_4378,N_4328);
nor U4424 (N_4424,N_4350,N_4313);
or U4425 (N_4425,N_4358,N_4300);
and U4426 (N_4426,N_4385,N_4257);
and U4427 (N_4427,N_4341,N_4359);
nor U4428 (N_4428,N_4283,N_4234);
xor U4429 (N_4429,N_4236,N_4245);
nor U4430 (N_4430,N_4331,N_4345);
and U4431 (N_4431,N_4303,N_4334);
xor U4432 (N_4432,N_4306,N_4265);
xnor U4433 (N_4433,N_4307,N_4337);
or U4434 (N_4434,N_4301,N_4332);
nor U4435 (N_4435,N_4231,N_4396);
nand U4436 (N_4436,N_4248,N_4319);
xnor U4437 (N_4437,N_4289,N_4302);
xnor U4438 (N_4438,N_4207,N_4233);
nor U4439 (N_4439,N_4254,N_4282);
and U4440 (N_4440,N_4255,N_4240);
and U4441 (N_4441,N_4383,N_4376);
and U4442 (N_4442,N_4368,N_4262);
and U4443 (N_4443,N_4261,N_4281);
and U4444 (N_4444,N_4384,N_4227);
and U4445 (N_4445,N_4398,N_4343);
nand U4446 (N_4446,N_4213,N_4237);
nand U4447 (N_4447,N_4274,N_4296);
xor U4448 (N_4448,N_4204,N_4298);
xor U4449 (N_4449,N_4320,N_4270);
or U4450 (N_4450,N_4291,N_4218);
nor U4451 (N_4451,N_4389,N_4315);
or U4452 (N_4452,N_4264,N_4220);
xnor U4453 (N_4453,N_4238,N_4308);
nor U4454 (N_4454,N_4221,N_4375);
and U4455 (N_4455,N_4228,N_4285);
xnor U4456 (N_4456,N_4208,N_4397);
xor U4457 (N_4457,N_4395,N_4369);
nor U4458 (N_4458,N_4347,N_4326);
nand U4459 (N_4459,N_4216,N_4366);
xnor U4460 (N_4460,N_4280,N_4351);
nand U4461 (N_4461,N_4304,N_4250);
xnor U4462 (N_4462,N_4235,N_4212);
or U4463 (N_4463,N_4356,N_4284);
nor U4464 (N_4464,N_4371,N_4279);
xnor U4465 (N_4465,N_4305,N_4364);
or U4466 (N_4466,N_4211,N_4288);
and U4467 (N_4467,N_4339,N_4394);
nand U4468 (N_4468,N_4286,N_4239);
and U4469 (N_4469,N_4357,N_4247);
or U4470 (N_4470,N_4373,N_4365);
nor U4471 (N_4471,N_4354,N_4330);
nand U4472 (N_4472,N_4273,N_4340);
xor U4473 (N_4473,N_4260,N_4209);
and U4474 (N_4474,N_4321,N_4377);
xnor U4475 (N_4475,N_4297,N_4277);
xnor U4476 (N_4476,N_4251,N_4202);
xnor U4477 (N_4477,N_4224,N_4258);
xnor U4478 (N_4478,N_4348,N_4323);
nor U4479 (N_4479,N_4206,N_4210);
and U4480 (N_4480,N_4267,N_4362);
nor U4481 (N_4481,N_4253,N_4392);
nand U4482 (N_4482,N_4226,N_4214);
nand U4483 (N_4483,N_4353,N_4292);
nor U4484 (N_4484,N_4317,N_4316);
nand U4485 (N_4485,N_4309,N_4391);
xor U4486 (N_4486,N_4287,N_4246);
nor U4487 (N_4487,N_4271,N_4276);
nand U4488 (N_4488,N_4390,N_4311);
nand U4489 (N_4489,N_4342,N_4372);
nand U4490 (N_4490,N_4269,N_4249);
nand U4491 (N_4491,N_4203,N_4272);
and U4492 (N_4492,N_4299,N_4388);
nand U4493 (N_4493,N_4225,N_4219);
nor U4494 (N_4494,N_4275,N_4222);
and U4495 (N_4495,N_4333,N_4338);
xor U4496 (N_4496,N_4381,N_4201);
nor U4497 (N_4497,N_4324,N_4374);
nor U4498 (N_4498,N_4310,N_4295);
or U4499 (N_4499,N_4360,N_4217);
or U4500 (N_4500,N_4322,N_4319);
nor U4501 (N_4501,N_4365,N_4261);
nor U4502 (N_4502,N_4349,N_4201);
nand U4503 (N_4503,N_4377,N_4263);
nand U4504 (N_4504,N_4351,N_4258);
or U4505 (N_4505,N_4366,N_4231);
xnor U4506 (N_4506,N_4264,N_4381);
and U4507 (N_4507,N_4237,N_4392);
xnor U4508 (N_4508,N_4330,N_4312);
nor U4509 (N_4509,N_4279,N_4235);
nand U4510 (N_4510,N_4259,N_4331);
and U4511 (N_4511,N_4306,N_4312);
nor U4512 (N_4512,N_4246,N_4290);
xnor U4513 (N_4513,N_4256,N_4211);
or U4514 (N_4514,N_4292,N_4337);
or U4515 (N_4515,N_4239,N_4248);
nor U4516 (N_4516,N_4204,N_4351);
nor U4517 (N_4517,N_4315,N_4309);
and U4518 (N_4518,N_4261,N_4241);
xor U4519 (N_4519,N_4208,N_4252);
nand U4520 (N_4520,N_4381,N_4213);
xnor U4521 (N_4521,N_4276,N_4388);
nand U4522 (N_4522,N_4278,N_4237);
nand U4523 (N_4523,N_4318,N_4378);
nor U4524 (N_4524,N_4256,N_4384);
nand U4525 (N_4525,N_4245,N_4279);
nand U4526 (N_4526,N_4322,N_4278);
or U4527 (N_4527,N_4254,N_4326);
xnor U4528 (N_4528,N_4231,N_4376);
or U4529 (N_4529,N_4322,N_4256);
nor U4530 (N_4530,N_4360,N_4305);
nand U4531 (N_4531,N_4286,N_4228);
nor U4532 (N_4532,N_4304,N_4392);
and U4533 (N_4533,N_4389,N_4234);
xor U4534 (N_4534,N_4294,N_4203);
or U4535 (N_4535,N_4347,N_4356);
nand U4536 (N_4536,N_4305,N_4228);
nand U4537 (N_4537,N_4286,N_4272);
or U4538 (N_4538,N_4297,N_4228);
nand U4539 (N_4539,N_4342,N_4360);
nor U4540 (N_4540,N_4281,N_4231);
xnor U4541 (N_4541,N_4280,N_4347);
nor U4542 (N_4542,N_4394,N_4376);
or U4543 (N_4543,N_4319,N_4211);
nand U4544 (N_4544,N_4383,N_4240);
nand U4545 (N_4545,N_4254,N_4242);
and U4546 (N_4546,N_4391,N_4250);
xnor U4547 (N_4547,N_4313,N_4318);
and U4548 (N_4548,N_4222,N_4399);
or U4549 (N_4549,N_4341,N_4246);
or U4550 (N_4550,N_4334,N_4244);
or U4551 (N_4551,N_4342,N_4296);
nand U4552 (N_4552,N_4264,N_4252);
nand U4553 (N_4553,N_4344,N_4266);
nand U4554 (N_4554,N_4322,N_4341);
or U4555 (N_4555,N_4218,N_4389);
nand U4556 (N_4556,N_4229,N_4295);
xnor U4557 (N_4557,N_4381,N_4395);
xor U4558 (N_4558,N_4348,N_4265);
or U4559 (N_4559,N_4393,N_4290);
xnor U4560 (N_4560,N_4297,N_4226);
xnor U4561 (N_4561,N_4320,N_4393);
and U4562 (N_4562,N_4343,N_4238);
or U4563 (N_4563,N_4216,N_4251);
nand U4564 (N_4564,N_4280,N_4241);
nor U4565 (N_4565,N_4304,N_4390);
and U4566 (N_4566,N_4230,N_4277);
xor U4567 (N_4567,N_4266,N_4297);
or U4568 (N_4568,N_4313,N_4242);
nand U4569 (N_4569,N_4287,N_4389);
xor U4570 (N_4570,N_4245,N_4324);
nand U4571 (N_4571,N_4357,N_4241);
nand U4572 (N_4572,N_4229,N_4314);
or U4573 (N_4573,N_4368,N_4297);
xor U4574 (N_4574,N_4320,N_4306);
and U4575 (N_4575,N_4330,N_4277);
nand U4576 (N_4576,N_4270,N_4397);
xnor U4577 (N_4577,N_4277,N_4237);
nor U4578 (N_4578,N_4399,N_4216);
or U4579 (N_4579,N_4331,N_4290);
and U4580 (N_4580,N_4264,N_4364);
nand U4581 (N_4581,N_4260,N_4365);
and U4582 (N_4582,N_4297,N_4256);
or U4583 (N_4583,N_4299,N_4320);
and U4584 (N_4584,N_4303,N_4257);
nor U4585 (N_4585,N_4359,N_4354);
xor U4586 (N_4586,N_4366,N_4219);
xor U4587 (N_4587,N_4394,N_4269);
xor U4588 (N_4588,N_4339,N_4206);
or U4589 (N_4589,N_4357,N_4343);
and U4590 (N_4590,N_4269,N_4349);
and U4591 (N_4591,N_4374,N_4298);
and U4592 (N_4592,N_4385,N_4287);
xnor U4593 (N_4593,N_4282,N_4200);
or U4594 (N_4594,N_4233,N_4212);
and U4595 (N_4595,N_4209,N_4347);
or U4596 (N_4596,N_4243,N_4389);
and U4597 (N_4597,N_4338,N_4335);
or U4598 (N_4598,N_4262,N_4363);
or U4599 (N_4599,N_4380,N_4288);
or U4600 (N_4600,N_4457,N_4482);
and U4601 (N_4601,N_4499,N_4418);
and U4602 (N_4602,N_4444,N_4401);
or U4603 (N_4603,N_4589,N_4424);
and U4604 (N_4604,N_4497,N_4493);
nand U4605 (N_4605,N_4408,N_4478);
or U4606 (N_4606,N_4475,N_4443);
and U4607 (N_4607,N_4577,N_4413);
xnor U4608 (N_4608,N_4464,N_4470);
nand U4609 (N_4609,N_4542,N_4400);
nor U4610 (N_4610,N_4459,N_4540);
xor U4611 (N_4611,N_4455,N_4407);
nor U4612 (N_4612,N_4436,N_4437);
nand U4613 (N_4613,N_4513,N_4501);
or U4614 (N_4614,N_4532,N_4485);
or U4615 (N_4615,N_4557,N_4515);
xor U4616 (N_4616,N_4503,N_4519);
nor U4617 (N_4617,N_4525,N_4427);
and U4618 (N_4618,N_4546,N_4432);
nor U4619 (N_4619,N_4586,N_4495);
nor U4620 (N_4620,N_4576,N_4410);
or U4621 (N_4621,N_4544,N_4466);
nor U4622 (N_4622,N_4581,N_4488);
nand U4623 (N_4623,N_4504,N_4453);
and U4624 (N_4624,N_4403,N_4523);
nand U4625 (N_4625,N_4450,N_4541);
or U4626 (N_4626,N_4554,N_4484);
nor U4627 (N_4627,N_4426,N_4578);
or U4628 (N_4628,N_4406,N_4440);
or U4629 (N_4629,N_4476,N_4555);
nand U4630 (N_4630,N_4414,N_4489);
and U4631 (N_4631,N_4536,N_4458);
or U4632 (N_4632,N_4508,N_4526);
nor U4633 (N_4633,N_4452,N_4569);
or U4634 (N_4634,N_4518,N_4582);
and U4635 (N_4635,N_4528,N_4421);
or U4636 (N_4636,N_4556,N_4454);
or U4637 (N_4637,N_4509,N_4471);
nor U4638 (N_4638,N_4593,N_4469);
nor U4639 (N_4639,N_4533,N_4516);
xnor U4640 (N_4640,N_4438,N_4575);
or U4641 (N_4641,N_4531,N_4417);
and U4642 (N_4642,N_4598,N_4415);
nand U4643 (N_4643,N_4545,N_4416);
xor U4644 (N_4644,N_4590,N_4448);
or U4645 (N_4645,N_4588,N_4461);
xor U4646 (N_4646,N_4429,N_4490);
or U4647 (N_4647,N_4583,N_4492);
nor U4648 (N_4648,N_4404,N_4563);
and U4649 (N_4649,N_4442,N_4562);
nand U4650 (N_4650,N_4551,N_4434);
nand U4651 (N_4651,N_4433,N_4511);
nand U4652 (N_4652,N_4505,N_4502);
nand U4653 (N_4653,N_4498,N_4439);
xnor U4654 (N_4654,N_4566,N_4570);
nor U4655 (N_4655,N_4468,N_4594);
nor U4656 (N_4656,N_4596,N_4521);
nor U4657 (N_4657,N_4580,N_4462);
or U4658 (N_4658,N_4574,N_4483);
nor U4659 (N_4659,N_4571,N_4481);
or U4660 (N_4660,N_4445,N_4547);
and U4661 (N_4661,N_4573,N_4549);
or U4662 (N_4662,N_4599,N_4524);
xnor U4663 (N_4663,N_4435,N_4467);
xor U4664 (N_4664,N_4535,N_4465);
nor U4665 (N_4665,N_4587,N_4585);
nand U4666 (N_4666,N_4409,N_4486);
xnor U4667 (N_4667,N_4520,N_4510);
and U4668 (N_4668,N_4572,N_4534);
nor U4669 (N_4669,N_4474,N_4514);
and U4670 (N_4670,N_4412,N_4477);
or U4671 (N_4671,N_4480,N_4451);
and U4672 (N_4672,N_4422,N_4479);
nor U4673 (N_4673,N_4506,N_4472);
nand U4674 (N_4674,N_4496,N_4552);
and U4675 (N_4675,N_4405,N_4463);
nor U4676 (N_4676,N_4512,N_4446);
and U4677 (N_4677,N_4560,N_4584);
or U4678 (N_4678,N_4564,N_4411);
xor U4679 (N_4679,N_4568,N_4529);
nor U4680 (N_4680,N_4567,N_4420);
nor U4681 (N_4681,N_4430,N_4507);
or U4682 (N_4682,N_4419,N_4565);
nand U4683 (N_4683,N_4431,N_4494);
and U4684 (N_4684,N_4423,N_4538);
and U4685 (N_4685,N_4500,N_4539);
nand U4686 (N_4686,N_4553,N_4428);
or U4687 (N_4687,N_4517,N_4473);
nand U4688 (N_4688,N_4561,N_4447);
nand U4689 (N_4689,N_4592,N_4530);
xnor U4690 (N_4690,N_4550,N_4548);
and U4691 (N_4691,N_4491,N_4522);
nand U4692 (N_4692,N_4456,N_4595);
and U4693 (N_4693,N_4441,N_4487);
nor U4694 (N_4694,N_4591,N_4537);
xor U4695 (N_4695,N_4425,N_4597);
xnor U4696 (N_4696,N_4559,N_4543);
and U4697 (N_4697,N_4527,N_4460);
nor U4698 (N_4698,N_4402,N_4558);
xnor U4699 (N_4699,N_4449,N_4579);
nor U4700 (N_4700,N_4431,N_4471);
nor U4701 (N_4701,N_4434,N_4427);
xor U4702 (N_4702,N_4542,N_4492);
or U4703 (N_4703,N_4475,N_4582);
nor U4704 (N_4704,N_4478,N_4409);
nor U4705 (N_4705,N_4501,N_4480);
nor U4706 (N_4706,N_4599,N_4480);
and U4707 (N_4707,N_4530,N_4544);
and U4708 (N_4708,N_4584,N_4476);
and U4709 (N_4709,N_4516,N_4424);
or U4710 (N_4710,N_4490,N_4550);
or U4711 (N_4711,N_4474,N_4552);
xnor U4712 (N_4712,N_4572,N_4428);
nor U4713 (N_4713,N_4511,N_4510);
xor U4714 (N_4714,N_4553,N_4418);
nor U4715 (N_4715,N_4413,N_4578);
nor U4716 (N_4716,N_4477,N_4506);
or U4717 (N_4717,N_4483,N_4583);
and U4718 (N_4718,N_4437,N_4467);
or U4719 (N_4719,N_4419,N_4524);
and U4720 (N_4720,N_4531,N_4569);
and U4721 (N_4721,N_4532,N_4481);
and U4722 (N_4722,N_4597,N_4440);
and U4723 (N_4723,N_4470,N_4438);
and U4724 (N_4724,N_4535,N_4474);
nor U4725 (N_4725,N_4522,N_4519);
nand U4726 (N_4726,N_4521,N_4440);
nor U4727 (N_4727,N_4409,N_4570);
nor U4728 (N_4728,N_4501,N_4430);
nand U4729 (N_4729,N_4518,N_4402);
nand U4730 (N_4730,N_4423,N_4553);
or U4731 (N_4731,N_4583,N_4527);
and U4732 (N_4732,N_4495,N_4494);
xnor U4733 (N_4733,N_4444,N_4575);
xor U4734 (N_4734,N_4472,N_4539);
nor U4735 (N_4735,N_4445,N_4538);
nor U4736 (N_4736,N_4593,N_4507);
and U4737 (N_4737,N_4455,N_4566);
xnor U4738 (N_4738,N_4547,N_4517);
or U4739 (N_4739,N_4444,N_4464);
xor U4740 (N_4740,N_4559,N_4566);
or U4741 (N_4741,N_4596,N_4463);
or U4742 (N_4742,N_4471,N_4465);
nor U4743 (N_4743,N_4462,N_4599);
nor U4744 (N_4744,N_4556,N_4479);
nand U4745 (N_4745,N_4487,N_4535);
nor U4746 (N_4746,N_4555,N_4561);
nor U4747 (N_4747,N_4419,N_4416);
or U4748 (N_4748,N_4495,N_4535);
xnor U4749 (N_4749,N_4599,N_4499);
nor U4750 (N_4750,N_4461,N_4557);
and U4751 (N_4751,N_4501,N_4434);
or U4752 (N_4752,N_4429,N_4441);
xnor U4753 (N_4753,N_4465,N_4420);
or U4754 (N_4754,N_4403,N_4558);
and U4755 (N_4755,N_4488,N_4449);
xnor U4756 (N_4756,N_4485,N_4492);
xnor U4757 (N_4757,N_4592,N_4457);
or U4758 (N_4758,N_4437,N_4422);
xor U4759 (N_4759,N_4582,N_4453);
nand U4760 (N_4760,N_4475,N_4470);
or U4761 (N_4761,N_4524,N_4435);
xor U4762 (N_4762,N_4480,N_4458);
and U4763 (N_4763,N_4463,N_4409);
or U4764 (N_4764,N_4536,N_4572);
nor U4765 (N_4765,N_4549,N_4443);
nand U4766 (N_4766,N_4525,N_4491);
nor U4767 (N_4767,N_4586,N_4496);
and U4768 (N_4768,N_4450,N_4443);
or U4769 (N_4769,N_4571,N_4512);
nor U4770 (N_4770,N_4486,N_4408);
and U4771 (N_4771,N_4579,N_4429);
or U4772 (N_4772,N_4566,N_4424);
and U4773 (N_4773,N_4577,N_4422);
or U4774 (N_4774,N_4416,N_4442);
or U4775 (N_4775,N_4421,N_4593);
and U4776 (N_4776,N_4525,N_4526);
xnor U4777 (N_4777,N_4513,N_4519);
and U4778 (N_4778,N_4597,N_4543);
xnor U4779 (N_4779,N_4512,N_4449);
or U4780 (N_4780,N_4418,N_4433);
and U4781 (N_4781,N_4484,N_4479);
or U4782 (N_4782,N_4467,N_4488);
xor U4783 (N_4783,N_4580,N_4514);
nor U4784 (N_4784,N_4557,N_4564);
xnor U4785 (N_4785,N_4469,N_4530);
nand U4786 (N_4786,N_4457,N_4540);
nor U4787 (N_4787,N_4555,N_4433);
xnor U4788 (N_4788,N_4414,N_4412);
and U4789 (N_4789,N_4484,N_4500);
nand U4790 (N_4790,N_4437,N_4546);
or U4791 (N_4791,N_4549,N_4546);
nand U4792 (N_4792,N_4431,N_4403);
nand U4793 (N_4793,N_4549,N_4404);
and U4794 (N_4794,N_4506,N_4493);
xor U4795 (N_4795,N_4484,N_4556);
xnor U4796 (N_4796,N_4472,N_4423);
nor U4797 (N_4797,N_4555,N_4582);
xnor U4798 (N_4798,N_4452,N_4572);
nor U4799 (N_4799,N_4497,N_4549);
or U4800 (N_4800,N_4703,N_4719);
xnor U4801 (N_4801,N_4665,N_4658);
xor U4802 (N_4802,N_4761,N_4708);
and U4803 (N_4803,N_4768,N_4734);
xor U4804 (N_4804,N_4695,N_4773);
or U4805 (N_4805,N_4652,N_4687);
nand U4806 (N_4806,N_4739,N_4779);
xnor U4807 (N_4807,N_4644,N_4740);
and U4808 (N_4808,N_4758,N_4612);
or U4809 (N_4809,N_4711,N_4627);
nor U4810 (N_4810,N_4678,N_4682);
xor U4811 (N_4811,N_4771,N_4737);
or U4812 (N_4812,N_4704,N_4726);
or U4813 (N_4813,N_4759,N_4750);
or U4814 (N_4814,N_4661,N_4632);
and U4815 (N_4815,N_4664,N_4693);
nor U4816 (N_4816,N_4622,N_4662);
nor U4817 (N_4817,N_4784,N_4718);
nand U4818 (N_4818,N_4756,N_4694);
xor U4819 (N_4819,N_4769,N_4600);
or U4820 (N_4820,N_4729,N_4616);
or U4821 (N_4821,N_4651,N_4723);
xor U4822 (N_4822,N_4765,N_4645);
or U4823 (N_4823,N_4762,N_4710);
xnor U4824 (N_4824,N_4775,N_4684);
xor U4825 (N_4825,N_4618,N_4639);
nor U4826 (N_4826,N_4626,N_4787);
nor U4827 (N_4827,N_4748,N_4667);
nand U4828 (N_4828,N_4701,N_4780);
nor U4829 (N_4829,N_4716,N_4713);
or U4830 (N_4830,N_4741,N_4605);
or U4831 (N_4831,N_4625,N_4659);
xor U4832 (N_4832,N_4673,N_4637);
xor U4833 (N_4833,N_4619,N_4776);
or U4834 (N_4834,N_4725,N_4670);
or U4835 (N_4835,N_4689,N_4757);
nand U4836 (N_4836,N_4636,N_4717);
nor U4837 (N_4837,N_4763,N_4743);
nor U4838 (N_4838,N_4609,N_4677);
nand U4839 (N_4839,N_4793,N_4614);
or U4840 (N_4840,N_4751,N_4706);
xnor U4841 (N_4841,N_4755,N_4714);
and U4842 (N_4842,N_4640,N_4753);
or U4843 (N_4843,N_4727,N_4754);
or U4844 (N_4844,N_4642,N_4786);
and U4845 (N_4845,N_4766,N_4728);
or U4846 (N_4846,N_4767,N_4646);
xor U4847 (N_4847,N_4730,N_4715);
and U4848 (N_4848,N_4702,N_4615);
nand U4849 (N_4849,N_4660,N_4772);
or U4850 (N_4850,N_4795,N_4641);
and U4851 (N_4851,N_4604,N_4613);
xor U4852 (N_4852,N_4672,N_4668);
nor U4853 (N_4853,N_4746,N_4606);
nand U4854 (N_4854,N_4623,N_4679);
or U4855 (N_4855,N_4690,N_4676);
nor U4856 (N_4856,N_4634,N_4601);
nor U4857 (N_4857,N_4620,N_4791);
and U4858 (N_4858,N_4731,N_4778);
xnor U4859 (N_4859,N_4752,N_4732);
or U4860 (N_4860,N_4745,N_4610);
nor U4861 (N_4861,N_4736,N_4788);
xnor U4862 (N_4862,N_4783,N_4671);
nor U4863 (N_4863,N_4770,N_4656);
or U4864 (N_4864,N_4697,N_4712);
nand U4865 (N_4865,N_4698,N_4735);
and U4866 (N_4866,N_4692,N_4685);
and U4867 (N_4867,N_4603,N_4624);
nand U4868 (N_4868,N_4633,N_4655);
nor U4869 (N_4869,N_4797,N_4647);
or U4870 (N_4870,N_4629,N_4781);
xnor U4871 (N_4871,N_4691,N_4738);
nor U4872 (N_4872,N_4631,N_4749);
nor U4873 (N_4873,N_4721,N_4635);
and U4874 (N_4874,N_4675,N_4621);
nor U4875 (N_4875,N_4798,N_4777);
and U4876 (N_4876,N_4617,N_4669);
xor U4877 (N_4877,N_4648,N_4782);
xor U4878 (N_4878,N_4747,N_4796);
nor U4879 (N_4879,N_4680,N_4683);
xor U4880 (N_4880,N_4709,N_4602);
nand U4881 (N_4881,N_4744,N_4774);
xor U4882 (N_4882,N_4760,N_4607);
and U4883 (N_4883,N_4643,N_4666);
nand U4884 (N_4884,N_4653,N_4794);
or U4885 (N_4885,N_4705,N_4654);
nand U4886 (N_4886,N_4707,N_4688);
nor U4887 (N_4887,N_4663,N_4681);
and U4888 (N_4888,N_4611,N_4724);
nand U4889 (N_4889,N_4649,N_4789);
nor U4890 (N_4890,N_4790,N_4742);
nand U4891 (N_4891,N_4764,N_4792);
or U4892 (N_4892,N_4696,N_4628);
xor U4893 (N_4893,N_4638,N_4733);
nand U4894 (N_4894,N_4700,N_4799);
nor U4895 (N_4895,N_4686,N_4785);
nor U4896 (N_4896,N_4630,N_4699);
xnor U4897 (N_4897,N_4722,N_4608);
nor U4898 (N_4898,N_4657,N_4674);
nand U4899 (N_4899,N_4650,N_4720);
nand U4900 (N_4900,N_4738,N_4776);
xnor U4901 (N_4901,N_4793,N_4674);
or U4902 (N_4902,N_4786,N_4643);
or U4903 (N_4903,N_4634,N_4717);
nand U4904 (N_4904,N_4714,N_4682);
nand U4905 (N_4905,N_4679,N_4682);
or U4906 (N_4906,N_4745,N_4657);
and U4907 (N_4907,N_4779,N_4685);
xor U4908 (N_4908,N_4666,N_4693);
xnor U4909 (N_4909,N_4781,N_4720);
or U4910 (N_4910,N_4694,N_4619);
and U4911 (N_4911,N_4734,N_4659);
xnor U4912 (N_4912,N_4726,N_4723);
xor U4913 (N_4913,N_4610,N_4788);
and U4914 (N_4914,N_4752,N_4618);
xor U4915 (N_4915,N_4778,N_4661);
nor U4916 (N_4916,N_4723,N_4661);
xnor U4917 (N_4917,N_4672,N_4771);
xor U4918 (N_4918,N_4654,N_4656);
or U4919 (N_4919,N_4737,N_4635);
or U4920 (N_4920,N_4770,N_4695);
or U4921 (N_4921,N_4694,N_4700);
nand U4922 (N_4922,N_4649,N_4792);
or U4923 (N_4923,N_4752,N_4711);
nor U4924 (N_4924,N_4649,N_4796);
nor U4925 (N_4925,N_4791,N_4729);
or U4926 (N_4926,N_4686,N_4667);
nand U4927 (N_4927,N_4690,N_4648);
nand U4928 (N_4928,N_4667,N_4764);
xnor U4929 (N_4929,N_4689,N_4722);
or U4930 (N_4930,N_4696,N_4751);
nand U4931 (N_4931,N_4693,N_4752);
nor U4932 (N_4932,N_4653,N_4708);
and U4933 (N_4933,N_4736,N_4749);
nand U4934 (N_4934,N_4740,N_4627);
nor U4935 (N_4935,N_4693,N_4710);
and U4936 (N_4936,N_4698,N_4670);
nor U4937 (N_4937,N_4755,N_4615);
nand U4938 (N_4938,N_4649,N_4690);
or U4939 (N_4939,N_4601,N_4635);
xnor U4940 (N_4940,N_4699,N_4650);
xnor U4941 (N_4941,N_4795,N_4698);
and U4942 (N_4942,N_4791,N_4799);
nand U4943 (N_4943,N_4668,N_4727);
and U4944 (N_4944,N_4762,N_4651);
nor U4945 (N_4945,N_4788,N_4692);
nor U4946 (N_4946,N_4601,N_4722);
nor U4947 (N_4947,N_4743,N_4731);
nor U4948 (N_4948,N_4771,N_4656);
nand U4949 (N_4949,N_4636,N_4700);
nand U4950 (N_4950,N_4674,N_4621);
nor U4951 (N_4951,N_4778,N_4768);
nor U4952 (N_4952,N_4620,N_4767);
and U4953 (N_4953,N_4794,N_4792);
xnor U4954 (N_4954,N_4623,N_4682);
nor U4955 (N_4955,N_4721,N_4777);
nor U4956 (N_4956,N_4716,N_4752);
nor U4957 (N_4957,N_4769,N_4734);
xnor U4958 (N_4958,N_4712,N_4626);
or U4959 (N_4959,N_4620,N_4759);
nand U4960 (N_4960,N_4659,N_4796);
xnor U4961 (N_4961,N_4735,N_4754);
or U4962 (N_4962,N_4704,N_4724);
nor U4963 (N_4963,N_4636,N_4650);
nand U4964 (N_4964,N_4726,N_4624);
or U4965 (N_4965,N_4777,N_4637);
and U4966 (N_4966,N_4757,N_4769);
or U4967 (N_4967,N_4746,N_4762);
xor U4968 (N_4968,N_4687,N_4792);
nor U4969 (N_4969,N_4643,N_4727);
and U4970 (N_4970,N_4608,N_4782);
nor U4971 (N_4971,N_4695,N_4658);
xor U4972 (N_4972,N_4696,N_4680);
nor U4973 (N_4973,N_4648,N_4640);
nor U4974 (N_4974,N_4769,N_4749);
nand U4975 (N_4975,N_4693,N_4679);
or U4976 (N_4976,N_4674,N_4788);
and U4977 (N_4977,N_4707,N_4741);
or U4978 (N_4978,N_4716,N_4678);
nor U4979 (N_4979,N_4738,N_4775);
and U4980 (N_4980,N_4653,N_4689);
nand U4981 (N_4981,N_4779,N_4677);
xnor U4982 (N_4982,N_4678,N_4740);
and U4983 (N_4983,N_4638,N_4788);
nor U4984 (N_4984,N_4722,N_4681);
nand U4985 (N_4985,N_4632,N_4774);
nor U4986 (N_4986,N_4723,N_4708);
and U4987 (N_4987,N_4755,N_4768);
or U4988 (N_4988,N_4607,N_4669);
or U4989 (N_4989,N_4751,N_4615);
xnor U4990 (N_4990,N_4760,N_4779);
xor U4991 (N_4991,N_4614,N_4797);
nand U4992 (N_4992,N_4753,N_4642);
and U4993 (N_4993,N_4602,N_4743);
and U4994 (N_4994,N_4768,N_4706);
or U4995 (N_4995,N_4674,N_4772);
xnor U4996 (N_4996,N_4653,N_4603);
nor U4997 (N_4997,N_4741,N_4774);
and U4998 (N_4998,N_4602,N_4717);
nor U4999 (N_4999,N_4601,N_4746);
or U5000 (N_5000,N_4816,N_4822);
and U5001 (N_5001,N_4872,N_4910);
xor U5002 (N_5002,N_4940,N_4946);
and U5003 (N_5003,N_4800,N_4879);
xor U5004 (N_5004,N_4884,N_4936);
or U5005 (N_5005,N_4804,N_4916);
xnor U5006 (N_5006,N_4904,N_4999);
nand U5007 (N_5007,N_4896,N_4856);
nor U5008 (N_5008,N_4829,N_4931);
and U5009 (N_5009,N_4906,N_4923);
nor U5010 (N_5010,N_4888,N_4960);
and U5011 (N_5011,N_4813,N_4998);
or U5012 (N_5012,N_4964,N_4847);
nor U5013 (N_5013,N_4803,N_4994);
nand U5014 (N_5014,N_4870,N_4966);
or U5015 (N_5015,N_4893,N_4915);
nand U5016 (N_5016,N_4945,N_4920);
and U5017 (N_5017,N_4868,N_4877);
nor U5018 (N_5018,N_4836,N_4984);
nand U5019 (N_5019,N_4842,N_4841);
nor U5020 (N_5020,N_4883,N_4860);
nor U5021 (N_5021,N_4832,N_4809);
nor U5022 (N_5022,N_4972,N_4821);
or U5023 (N_5023,N_4963,N_4948);
nand U5024 (N_5024,N_4876,N_4957);
and U5025 (N_5025,N_4887,N_4970);
or U5026 (N_5026,N_4983,N_4834);
xor U5027 (N_5027,N_4875,N_4878);
nor U5028 (N_5028,N_4808,N_4993);
nor U5029 (N_5029,N_4955,N_4965);
nor U5030 (N_5030,N_4918,N_4973);
or U5031 (N_5031,N_4978,N_4996);
and U5032 (N_5032,N_4845,N_4944);
nor U5033 (N_5033,N_4864,N_4928);
or U5034 (N_5034,N_4982,N_4979);
nand U5035 (N_5035,N_4851,N_4871);
nand U5036 (N_5036,N_4837,N_4953);
nand U5037 (N_5037,N_4924,N_4812);
nand U5038 (N_5038,N_4988,N_4891);
nor U5039 (N_5039,N_4853,N_4905);
xor U5040 (N_5040,N_4838,N_4956);
xor U5041 (N_5041,N_4861,N_4850);
or U5042 (N_5042,N_4977,N_4814);
or U5043 (N_5043,N_4943,N_4952);
or U5044 (N_5044,N_4818,N_4810);
xor U5045 (N_5045,N_4912,N_4911);
and U5046 (N_5046,N_4846,N_4852);
and U5047 (N_5047,N_4902,N_4898);
nor U5048 (N_5048,N_4863,N_4951);
xnor U5049 (N_5049,N_4947,N_4806);
xnor U5050 (N_5050,N_4865,N_4817);
nand U5051 (N_5051,N_4941,N_4843);
or U5052 (N_5052,N_4828,N_4919);
xor U5053 (N_5053,N_4981,N_4913);
or U5054 (N_5054,N_4932,N_4985);
xor U5055 (N_5055,N_4989,N_4938);
nor U5056 (N_5056,N_4901,N_4921);
and U5057 (N_5057,N_4844,N_4987);
or U5058 (N_5058,N_4926,N_4908);
or U5059 (N_5059,N_4967,N_4899);
and U5060 (N_5060,N_4820,N_4885);
nor U5061 (N_5061,N_4805,N_4819);
and U5062 (N_5062,N_4975,N_4854);
or U5063 (N_5063,N_4831,N_4857);
xnor U5064 (N_5064,N_4897,N_4825);
xor U5065 (N_5065,N_4930,N_4866);
and U5066 (N_5066,N_4824,N_4811);
nor U5067 (N_5067,N_4874,N_4990);
nor U5068 (N_5068,N_4886,N_4802);
and U5069 (N_5069,N_4937,N_4942);
nand U5070 (N_5070,N_4917,N_4929);
or U5071 (N_5071,N_4949,N_4889);
or U5072 (N_5072,N_4968,N_4992);
xnor U5073 (N_5073,N_4950,N_4873);
nor U5074 (N_5074,N_4986,N_4991);
or U5075 (N_5075,N_4858,N_4974);
or U5076 (N_5076,N_4959,N_4823);
nand U5077 (N_5077,N_4976,N_4934);
and U5078 (N_5078,N_4835,N_4840);
nor U5079 (N_5079,N_4848,N_4907);
or U5080 (N_5080,N_4859,N_4958);
nand U5081 (N_5081,N_4839,N_4890);
and U5082 (N_5082,N_4939,N_4880);
nand U5083 (N_5083,N_4922,N_4869);
xnor U5084 (N_5084,N_4815,N_4995);
xor U5085 (N_5085,N_4881,N_4980);
nor U5086 (N_5086,N_4807,N_4833);
nand U5087 (N_5087,N_4954,N_4971);
nand U5088 (N_5088,N_4909,N_4855);
xor U5089 (N_5089,N_4892,N_4826);
xor U5090 (N_5090,N_4961,N_4969);
and U5091 (N_5091,N_4925,N_4914);
nor U5092 (N_5092,N_4933,N_4882);
nor U5093 (N_5093,N_4935,N_4827);
xnor U5094 (N_5094,N_4997,N_4862);
and U5095 (N_5095,N_4900,N_4903);
or U5096 (N_5096,N_4927,N_4895);
and U5097 (N_5097,N_4801,N_4849);
nand U5098 (N_5098,N_4894,N_4830);
nor U5099 (N_5099,N_4867,N_4962);
xnor U5100 (N_5100,N_4919,N_4971);
nand U5101 (N_5101,N_4945,N_4977);
and U5102 (N_5102,N_4828,N_4890);
or U5103 (N_5103,N_4875,N_4915);
xor U5104 (N_5104,N_4967,N_4989);
or U5105 (N_5105,N_4933,N_4980);
or U5106 (N_5106,N_4847,N_4830);
and U5107 (N_5107,N_4827,N_4841);
and U5108 (N_5108,N_4830,N_4886);
xnor U5109 (N_5109,N_4824,N_4996);
and U5110 (N_5110,N_4907,N_4958);
nand U5111 (N_5111,N_4825,N_4821);
xor U5112 (N_5112,N_4940,N_4871);
and U5113 (N_5113,N_4924,N_4942);
xnor U5114 (N_5114,N_4946,N_4986);
xnor U5115 (N_5115,N_4890,N_4886);
nand U5116 (N_5116,N_4956,N_4831);
xnor U5117 (N_5117,N_4902,N_4981);
nand U5118 (N_5118,N_4933,N_4869);
nand U5119 (N_5119,N_4887,N_4972);
and U5120 (N_5120,N_4823,N_4837);
xor U5121 (N_5121,N_4904,N_4814);
and U5122 (N_5122,N_4904,N_4883);
nor U5123 (N_5123,N_4898,N_4818);
xor U5124 (N_5124,N_4896,N_4956);
nor U5125 (N_5125,N_4858,N_4827);
and U5126 (N_5126,N_4988,N_4896);
and U5127 (N_5127,N_4977,N_4928);
nand U5128 (N_5128,N_4875,N_4849);
nand U5129 (N_5129,N_4900,N_4858);
xor U5130 (N_5130,N_4807,N_4980);
nand U5131 (N_5131,N_4926,N_4988);
nor U5132 (N_5132,N_4995,N_4862);
nand U5133 (N_5133,N_4848,N_4807);
nand U5134 (N_5134,N_4888,N_4928);
nand U5135 (N_5135,N_4954,N_4910);
xnor U5136 (N_5136,N_4818,N_4901);
xor U5137 (N_5137,N_4856,N_4845);
xor U5138 (N_5138,N_4847,N_4931);
xor U5139 (N_5139,N_4878,N_4845);
xnor U5140 (N_5140,N_4821,N_4948);
nor U5141 (N_5141,N_4961,N_4940);
and U5142 (N_5142,N_4961,N_4933);
nor U5143 (N_5143,N_4825,N_4894);
nor U5144 (N_5144,N_4876,N_4976);
nand U5145 (N_5145,N_4877,N_4909);
or U5146 (N_5146,N_4914,N_4865);
or U5147 (N_5147,N_4829,N_4952);
nand U5148 (N_5148,N_4975,N_4963);
nor U5149 (N_5149,N_4924,N_4977);
nor U5150 (N_5150,N_4987,N_4927);
xnor U5151 (N_5151,N_4934,N_4948);
or U5152 (N_5152,N_4885,N_4874);
nand U5153 (N_5153,N_4969,N_4883);
and U5154 (N_5154,N_4904,N_4816);
or U5155 (N_5155,N_4862,N_4956);
and U5156 (N_5156,N_4811,N_4924);
nand U5157 (N_5157,N_4990,N_4916);
or U5158 (N_5158,N_4944,N_4839);
xor U5159 (N_5159,N_4889,N_4877);
and U5160 (N_5160,N_4811,N_4967);
and U5161 (N_5161,N_4968,N_4935);
or U5162 (N_5162,N_4934,N_4807);
nor U5163 (N_5163,N_4905,N_4919);
and U5164 (N_5164,N_4934,N_4997);
xor U5165 (N_5165,N_4898,N_4863);
or U5166 (N_5166,N_4820,N_4873);
xnor U5167 (N_5167,N_4846,N_4911);
and U5168 (N_5168,N_4806,N_4820);
and U5169 (N_5169,N_4917,N_4954);
and U5170 (N_5170,N_4848,N_4999);
and U5171 (N_5171,N_4910,N_4957);
xor U5172 (N_5172,N_4860,N_4811);
xnor U5173 (N_5173,N_4809,N_4970);
nand U5174 (N_5174,N_4824,N_4983);
or U5175 (N_5175,N_4901,N_4953);
nand U5176 (N_5176,N_4943,N_4924);
and U5177 (N_5177,N_4868,N_4992);
xor U5178 (N_5178,N_4987,N_4869);
or U5179 (N_5179,N_4905,N_4894);
or U5180 (N_5180,N_4945,N_4823);
nand U5181 (N_5181,N_4959,N_4995);
and U5182 (N_5182,N_4841,N_4860);
xor U5183 (N_5183,N_4941,N_4989);
nor U5184 (N_5184,N_4900,N_4848);
nand U5185 (N_5185,N_4903,N_4996);
and U5186 (N_5186,N_4889,N_4934);
and U5187 (N_5187,N_4818,N_4850);
nand U5188 (N_5188,N_4823,N_4936);
or U5189 (N_5189,N_4821,N_4927);
nand U5190 (N_5190,N_4864,N_4873);
xor U5191 (N_5191,N_4911,N_4948);
xnor U5192 (N_5192,N_4949,N_4818);
nand U5193 (N_5193,N_4868,N_4964);
nor U5194 (N_5194,N_4942,N_4821);
and U5195 (N_5195,N_4862,N_4922);
xor U5196 (N_5196,N_4982,N_4948);
xnor U5197 (N_5197,N_4819,N_4859);
nand U5198 (N_5198,N_4835,N_4881);
nand U5199 (N_5199,N_4831,N_4931);
or U5200 (N_5200,N_5174,N_5181);
and U5201 (N_5201,N_5173,N_5039);
xor U5202 (N_5202,N_5031,N_5194);
nor U5203 (N_5203,N_5095,N_5193);
or U5204 (N_5204,N_5102,N_5028);
nand U5205 (N_5205,N_5166,N_5001);
nand U5206 (N_5206,N_5184,N_5033);
or U5207 (N_5207,N_5189,N_5070);
and U5208 (N_5208,N_5148,N_5195);
nor U5209 (N_5209,N_5065,N_5067);
and U5210 (N_5210,N_5085,N_5069);
or U5211 (N_5211,N_5025,N_5160);
or U5212 (N_5212,N_5097,N_5197);
xnor U5213 (N_5213,N_5192,N_5199);
nand U5214 (N_5214,N_5037,N_5086);
or U5215 (N_5215,N_5052,N_5021);
and U5216 (N_5216,N_5058,N_5168);
or U5217 (N_5217,N_5083,N_5124);
nand U5218 (N_5218,N_5146,N_5182);
or U5219 (N_5219,N_5010,N_5096);
nor U5220 (N_5220,N_5051,N_5081);
nand U5221 (N_5221,N_5163,N_5005);
and U5222 (N_5222,N_5153,N_5015);
nor U5223 (N_5223,N_5161,N_5141);
or U5224 (N_5224,N_5105,N_5123);
or U5225 (N_5225,N_5013,N_5130);
and U5226 (N_5226,N_5167,N_5026);
nor U5227 (N_5227,N_5009,N_5027);
or U5228 (N_5228,N_5063,N_5186);
nand U5229 (N_5229,N_5034,N_5149);
or U5230 (N_5230,N_5073,N_5147);
or U5231 (N_5231,N_5156,N_5041);
and U5232 (N_5232,N_5094,N_5103);
or U5233 (N_5233,N_5177,N_5183);
or U5234 (N_5234,N_5162,N_5171);
or U5235 (N_5235,N_5113,N_5008);
xnor U5236 (N_5236,N_5061,N_5158);
or U5237 (N_5237,N_5165,N_5022);
xnor U5238 (N_5238,N_5169,N_5134);
nor U5239 (N_5239,N_5032,N_5084);
xnor U5240 (N_5240,N_5191,N_5030);
nand U5241 (N_5241,N_5108,N_5078);
nor U5242 (N_5242,N_5040,N_5072);
xor U5243 (N_5243,N_5057,N_5104);
xor U5244 (N_5244,N_5132,N_5012);
and U5245 (N_5245,N_5143,N_5109);
nand U5246 (N_5246,N_5098,N_5029);
or U5247 (N_5247,N_5106,N_5110);
and U5248 (N_5248,N_5131,N_5055);
nor U5249 (N_5249,N_5068,N_5119);
nor U5250 (N_5250,N_5175,N_5107);
xor U5251 (N_5251,N_5079,N_5135);
nor U5252 (N_5252,N_5101,N_5114);
xnor U5253 (N_5253,N_5053,N_5198);
nor U5254 (N_5254,N_5017,N_5154);
nand U5255 (N_5255,N_5064,N_5118);
nand U5256 (N_5256,N_5044,N_5170);
and U5257 (N_5257,N_5150,N_5122);
nor U5258 (N_5258,N_5112,N_5002);
or U5259 (N_5259,N_5187,N_5020);
or U5260 (N_5260,N_5144,N_5159);
nand U5261 (N_5261,N_5140,N_5116);
nor U5262 (N_5262,N_5076,N_5023);
nand U5263 (N_5263,N_5011,N_5007);
nor U5264 (N_5264,N_5090,N_5120);
xnor U5265 (N_5265,N_5050,N_5045);
and U5266 (N_5266,N_5136,N_5049);
and U5267 (N_5267,N_5059,N_5093);
nand U5268 (N_5268,N_5151,N_5185);
xor U5269 (N_5269,N_5074,N_5139);
and U5270 (N_5270,N_5180,N_5099);
and U5271 (N_5271,N_5176,N_5054);
xnor U5272 (N_5272,N_5047,N_5121);
or U5273 (N_5273,N_5137,N_5035);
or U5274 (N_5274,N_5000,N_5129);
xor U5275 (N_5275,N_5127,N_5066);
or U5276 (N_5276,N_5077,N_5080);
xnor U5277 (N_5277,N_5016,N_5196);
nor U5278 (N_5278,N_5133,N_5060);
nor U5279 (N_5279,N_5089,N_5138);
nand U5280 (N_5280,N_5046,N_5125);
xor U5281 (N_5281,N_5024,N_5164);
nor U5282 (N_5282,N_5004,N_5014);
or U5283 (N_5283,N_5006,N_5038);
xnor U5284 (N_5284,N_5117,N_5100);
xnor U5285 (N_5285,N_5178,N_5092);
xnor U5286 (N_5286,N_5082,N_5075);
xor U5287 (N_5287,N_5111,N_5190);
or U5288 (N_5288,N_5003,N_5126);
nor U5289 (N_5289,N_5179,N_5152);
or U5290 (N_5290,N_5071,N_5188);
and U5291 (N_5291,N_5157,N_5048);
xnor U5292 (N_5292,N_5172,N_5062);
and U5293 (N_5293,N_5128,N_5088);
xnor U5294 (N_5294,N_5036,N_5142);
nor U5295 (N_5295,N_5043,N_5145);
nand U5296 (N_5296,N_5042,N_5056);
and U5297 (N_5297,N_5019,N_5091);
or U5298 (N_5298,N_5115,N_5087);
nand U5299 (N_5299,N_5155,N_5018);
and U5300 (N_5300,N_5148,N_5180);
nand U5301 (N_5301,N_5112,N_5060);
xor U5302 (N_5302,N_5066,N_5069);
xnor U5303 (N_5303,N_5134,N_5130);
or U5304 (N_5304,N_5163,N_5000);
or U5305 (N_5305,N_5030,N_5061);
nor U5306 (N_5306,N_5179,N_5049);
nor U5307 (N_5307,N_5138,N_5121);
or U5308 (N_5308,N_5080,N_5007);
nor U5309 (N_5309,N_5103,N_5085);
xnor U5310 (N_5310,N_5047,N_5089);
xor U5311 (N_5311,N_5048,N_5133);
nand U5312 (N_5312,N_5056,N_5152);
xor U5313 (N_5313,N_5071,N_5195);
or U5314 (N_5314,N_5097,N_5148);
xnor U5315 (N_5315,N_5055,N_5112);
and U5316 (N_5316,N_5191,N_5098);
xor U5317 (N_5317,N_5178,N_5063);
nor U5318 (N_5318,N_5041,N_5153);
xnor U5319 (N_5319,N_5139,N_5115);
xnor U5320 (N_5320,N_5096,N_5015);
or U5321 (N_5321,N_5192,N_5166);
nand U5322 (N_5322,N_5135,N_5113);
nor U5323 (N_5323,N_5150,N_5184);
xnor U5324 (N_5324,N_5052,N_5059);
and U5325 (N_5325,N_5192,N_5023);
or U5326 (N_5326,N_5115,N_5062);
xor U5327 (N_5327,N_5018,N_5024);
nor U5328 (N_5328,N_5082,N_5017);
or U5329 (N_5329,N_5157,N_5150);
nor U5330 (N_5330,N_5154,N_5111);
and U5331 (N_5331,N_5095,N_5120);
and U5332 (N_5332,N_5127,N_5022);
nand U5333 (N_5333,N_5199,N_5019);
nor U5334 (N_5334,N_5084,N_5069);
and U5335 (N_5335,N_5031,N_5148);
or U5336 (N_5336,N_5057,N_5109);
nand U5337 (N_5337,N_5090,N_5129);
and U5338 (N_5338,N_5097,N_5124);
or U5339 (N_5339,N_5059,N_5028);
nor U5340 (N_5340,N_5148,N_5019);
nand U5341 (N_5341,N_5076,N_5143);
or U5342 (N_5342,N_5194,N_5026);
xnor U5343 (N_5343,N_5027,N_5064);
xor U5344 (N_5344,N_5005,N_5043);
and U5345 (N_5345,N_5180,N_5005);
or U5346 (N_5346,N_5003,N_5170);
nor U5347 (N_5347,N_5016,N_5134);
and U5348 (N_5348,N_5189,N_5102);
and U5349 (N_5349,N_5081,N_5147);
nand U5350 (N_5350,N_5152,N_5012);
nand U5351 (N_5351,N_5108,N_5166);
nand U5352 (N_5352,N_5099,N_5109);
and U5353 (N_5353,N_5011,N_5129);
and U5354 (N_5354,N_5073,N_5154);
and U5355 (N_5355,N_5082,N_5186);
and U5356 (N_5356,N_5046,N_5098);
nand U5357 (N_5357,N_5139,N_5192);
and U5358 (N_5358,N_5064,N_5158);
and U5359 (N_5359,N_5015,N_5184);
nor U5360 (N_5360,N_5009,N_5048);
or U5361 (N_5361,N_5082,N_5080);
or U5362 (N_5362,N_5050,N_5115);
nor U5363 (N_5363,N_5008,N_5062);
xor U5364 (N_5364,N_5022,N_5191);
xnor U5365 (N_5365,N_5111,N_5043);
nand U5366 (N_5366,N_5015,N_5188);
and U5367 (N_5367,N_5114,N_5006);
xnor U5368 (N_5368,N_5003,N_5041);
or U5369 (N_5369,N_5174,N_5080);
xnor U5370 (N_5370,N_5094,N_5122);
and U5371 (N_5371,N_5055,N_5114);
and U5372 (N_5372,N_5025,N_5145);
or U5373 (N_5373,N_5034,N_5093);
or U5374 (N_5374,N_5158,N_5144);
and U5375 (N_5375,N_5108,N_5042);
and U5376 (N_5376,N_5046,N_5021);
and U5377 (N_5377,N_5190,N_5185);
nor U5378 (N_5378,N_5057,N_5024);
nand U5379 (N_5379,N_5181,N_5159);
nor U5380 (N_5380,N_5113,N_5144);
xnor U5381 (N_5381,N_5027,N_5160);
and U5382 (N_5382,N_5061,N_5100);
nor U5383 (N_5383,N_5131,N_5151);
xnor U5384 (N_5384,N_5026,N_5127);
nor U5385 (N_5385,N_5069,N_5096);
xor U5386 (N_5386,N_5125,N_5059);
nor U5387 (N_5387,N_5190,N_5177);
nor U5388 (N_5388,N_5152,N_5133);
and U5389 (N_5389,N_5068,N_5088);
nor U5390 (N_5390,N_5106,N_5061);
or U5391 (N_5391,N_5187,N_5183);
and U5392 (N_5392,N_5069,N_5009);
xor U5393 (N_5393,N_5048,N_5051);
xor U5394 (N_5394,N_5133,N_5164);
or U5395 (N_5395,N_5135,N_5140);
nand U5396 (N_5396,N_5093,N_5169);
nand U5397 (N_5397,N_5185,N_5120);
xnor U5398 (N_5398,N_5045,N_5099);
nand U5399 (N_5399,N_5049,N_5059);
or U5400 (N_5400,N_5204,N_5270);
and U5401 (N_5401,N_5207,N_5316);
nor U5402 (N_5402,N_5216,N_5311);
or U5403 (N_5403,N_5217,N_5236);
xor U5404 (N_5404,N_5266,N_5338);
and U5405 (N_5405,N_5239,N_5278);
and U5406 (N_5406,N_5276,N_5214);
xnor U5407 (N_5407,N_5227,N_5347);
nor U5408 (N_5408,N_5326,N_5357);
nand U5409 (N_5409,N_5301,N_5255);
or U5410 (N_5410,N_5244,N_5298);
nor U5411 (N_5411,N_5283,N_5291);
xor U5412 (N_5412,N_5224,N_5238);
or U5413 (N_5413,N_5257,N_5287);
xnor U5414 (N_5414,N_5372,N_5215);
xnor U5415 (N_5415,N_5218,N_5213);
xnor U5416 (N_5416,N_5233,N_5340);
nor U5417 (N_5417,N_5376,N_5303);
nand U5418 (N_5418,N_5265,N_5329);
nor U5419 (N_5419,N_5264,N_5379);
or U5420 (N_5420,N_5263,N_5286);
or U5421 (N_5421,N_5354,N_5353);
or U5422 (N_5422,N_5267,N_5350);
nor U5423 (N_5423,N_5281,N_5334);
and U5424 (N_5424,N_5200,N_5261);
or U5425 (N_5425,N_5229,N_5295);
nor U5426 (N_5426,N_5302,N_5325);
nor U5427 (N_5427,N_5314,N_5285);
nor U5428 (N_5428,N_5332,N_5210);
nand U5429 (N_5429,N_5304,N_5247);
nor U5430 (N_5430,N_5253,N_5331);
or U5431 (N_5431,N_5346,N_5256);
and U5432 (N_5432,N_5203,N_5367);
and U5433 (N_5433,N_5380,N_5361);
xor U5434 (N_5434,N_5237,N_5232);
nor U5435 (N_5435,N_5387,N_5313);
xor U5436 (N_5436,N_5292,N_5308);
nand U5437 (N_5437,N_5339,N_5275);
nor U5438 (N_5438,N_5363,N_5274);
xor U5439 (N_5439,N_5359,N_5319);
or U5440 (N_5440,N_5254,N_5374);
xnor U5441 (N_5441,N_5317,N_5235);
nor U5442 (N_5442,N_5320,N_5395);
nand U5443 (N_5443,N_5370,N_5230);
nor U5444 (N_5444,N_5343,N_5392);
xor U5445 (N_5445,N_5335,N_5234);
or U5446 (N_5446,N_5269,N_5352);
or U5447 (N_5447,N_5279,N_5397);
or U5448 (N_5448,N_5362,N_5322);
nand U5449 (N_5449,N_5251,N_5226);
nor U5450 (N_5450,N_5321,N_5383);
nand U5451 (N_5451,N_5222,N_5345);
nand U5452 (N_5452,N_5356,N_5299);
nor U5453 (N_5453,N_5318,N_5341);
xor U5454 (N_5454,N_5300,N_5373);
or U5455 (N_5455,N_5242,N_5305);
or U5456 (N_5456,N_5202,N_5271);
and U5457 (N_5457,N_5310,N_5307);
nor U5458 (N_5458,N_5240,N_5272);
nor U5459 (N_5459,N_5327,N_5360);
and U5460 (N_5460,N_5220,N_5288);
or U5461 (N_5461,N_5246,N_5228);
and U5462 (N_5462,N_5368,N_5315);
nand U5463 (N_5463,N_5280,N_5208);
nand U5464 (N_5464,N_5337,N_5297);
and U5465 (N_5465,N_5394,N_5223);
nand U5466 (N_5466,N_5324,N_5323);
or U5467 (N_5467,N_5366,N_5348);
nand U5468 (N_5468,N_5277,N_5262);
xnor U5469 (N_5469,N_5282,N_5349);
nor U5470 (N_5470,N_5309,N_5389);
and U5471 (N_5471,N_5396,N_5289);
and U5472 (N_5472,N_5211,N_5273);
and U5473 (N_5473,N_5393,N_5312);
xor U5474 (N_5474,N_5260,N_5342);
xnor U5475 (N_5475,N_5250,N_5293);
or U5476 (N_5476,N_5371,N_5290);
or U5477 (N_5477,N_5245,N_5209);
and U5478 (N_5478,N_5221,N_5384);
or U5479 (N_5479,N_5385,N_5399);
xnor U5480 (N_5480,N_5248,N_5294);
and U5481 (N_5481,N_5382,N_5398);
and U5482 (N_5482,N_5268,N_5377);
nand U5483 (N_5483,N_5391,N_5375);
xor U5484 (N_5484,N_5201,N_5296);
or U5485 (N_5485,N_5206,N_5358);
and U5486 (N_5486,N_5369,N_5306);
xor U5487 (N_5487,N_5205,N_5212);
or U5488 (N_5488,N_5330,N_5344);
nand U5489 (N_5489,N_5388,N_5333);
and U5490 (N_5490,N_5364,N_5258);
nor U5491 (N_5491,N_5351,N_5386);
nor U5492 (N_5492,N_5252,N_5243);
or U5493 (N_5493,N_5231,N_5355);
nor U5494 (N_5494,N_5328,N_5336);
xor U5495 (N_5495,N_5365,N_5378);
or U5496 (N_5496,N_5219,N_5259);
xnor U5497 (N_5497,N_5249,N_5241);
and U5498 (N_5498,N_5390,N_5381);
xor U5499 (N_5499,N_5225,N_5284);
nand U5500 (N_5500,N_5227,N_5248);
or U5501 (N_5501,N_5317,N_5212);
xor U5502 (N_5502,N_5221,N_5245);
and U5503 (N_5503,N_5258,N_5375);
nand U5504 (N_5504,N_5308,N_5335);
nor U5505 (N_5505,N_5203,N_5250);
and U5506 (N_5506,N_5291,N_5242);
nor U5507 (N_5507,N_5228,N_5338);
xnor U5508 (N_5508,N_5259,N_5310);
and U5509 (N_5509,N_5205,N_5306);
xnor U5510 (N_5510,N_5266,N_5337);
and U5511 (N_5511,N_5366,N_5206);
or U5512 (N_5512,N_5304,N_5376);
or U5513 (N_5513,N_5381,N_5391);
or U5514 (N_5514,N_5283,N_5321);
or U5515 (N_5515,N_5354,N_5341);
or U5516 (N_5516,N_5202,N_5326);
nor U5517 (N_5517,N_5370,N_5304);
nor U5518 (N_5518,N_5371,N_5340);
nand U5519 (N_5519,N_5369,N_5288);
or U5520 (N_5520,N_5228,N_5256);
nand U5521 (N_5521,N_5361,N_5232);
nand U5522 (N_5522,N_5315,N_5286);
and U5523 (N_5523,N_5215,N_5345);
xnor U5524 (N_5524,N_5272,N_5317);
nor U5525 (N_5525,N_5278,N_5255);
xnor U5526 (N_5526,N_5337,N_5366);
nor U5527 (N_5527,N_5218,N_5360);
nor U5528 (N_5528,N_5399,N_5282);
nor U5529 (N_5529,N_5263,N_5289);
xor U5530 (N_5530,N_5268,N_5254);
nand U5531 (N_5531,N_5235,N_5205);
xor U5532 (N_5532,N_5320,N_5267);
nand U5533 (N_5533,N_5209,N_5248);
nand U5534 (N_5534,N_5265,N_5368);
xor U5535 (N_5535,N_5349,N_5231);
or U5536 (N_5536,N_5219,N_5342);
xnor U5537 (N_5537,N_5369,N_5200);
and U5538 (N_5538,N_5219,N_5377);
or U5539 (N_5539,N_5304,N_5299);
nand U5540 (N_5540,N_5261,N_5385);
or U5541 (N_5541,N_5370,N_5325);
or U5542 (N_5542,N_5275,N_5364);
nor U5543 (N_5543,N_5380,N_5354);
nand U5544 (N_5544,N_5223,N_5329);
nand U5545 (N_5545,N_5380,N_5322);
nor U5546 (N_5546,N_5353,N_5367);
and U5547 (N_5547,N_5387,N_5368);
or U5548 (N_5548,N_5308,N_5399);
xnor U5549 (N_5549,N_5323,N_5268);
xor U5550 (N_5550,N_5246,N_5269);
nor U5551 (N_5551,N_5318,N_5387);
and U5552 (N_5552,N_5393,N_5379);
or U5553 (N_5553,N_5340,N_5319);
xor U5554 (N_5554,N_5226,N_5349);
nand U5555 (N_5555,N_5248,N_5226);
nand U5556 (N_5556,N_5269,N_5334);
and U5557 (N_5557,N_5211,N_5221);
nor U5558 (N_5558,N_5269,N_5204);
nand U5559 (N_5559,N_5313,N_5251);
or U5560 (N_5560,N_5219,N_5333);
or U5561 (N_5561,N_5359,N_5393);
or U5562 (N_5562,N_5311,N_5364);
nor U5563 (N_5563,N_5342,N_5237);
nand U5564 (N_5564,N_5340,N_5290);
or U5565 (N_5565,N_5385,N_5299);
nor U5566 (N_5566,N_5271,N_5299);
nand U5567 (N_5567,N_5385,N_5223);
or U5568 (N_5568,N_5369,N_5379);
nand U5569 (N_5569,N_5399,N_5303);
nand U5570 (N_5570,N_5393,N_5295);
or U5571 (N_5571,N_5240,N_5336);
xor U5572 (N_5572,N_5391,N_5350);
nor U5573 (N_5573,N_5201,N_5358);
or U5574 (N_5574,N_5287,N_5288);
xnor U5575 (N_5575,N_5363,N_5307);
and U5576 (N_5576,N_5239,N_5373);
and U5577 (N_5577,N_5380,N_5284);
and U5578 (N_5578,N_5399,N_5365);
nand U5579 (N_5579,N_5324,N_5294);
and U5580 (N_5580,N_5241,N_5393);
xnor U5581 (N_5581,N_5260,N_5314);
and U5582 (N_5582,N_5280,N_5343);
or U5583 (N_5583,N_5306,N_5257);
nand U5584 (N_5584,N_5284,N_5252);
or U5585 (N_5585,N_5292,N_5350);
and U5586 (N_5586,N_5267,N_5274);
or U5587 (N_5587,N_5329,N_5383);
or U5588 (N_5588,N_5254,N_5206);
nand U5589 (N_5589,N_5230,N_5318);
or U5590 (N_5590,N_5284,N_5204);
and U5591 (N_5591,N_5383,N_5399);
nand U5592 (N_5592,N_5269,N_5369);
and U5593 (N_5593,N_5253,N_5351);
and U5594 (N_5594,N_5296,N_5388);
nand U5595 (N_5595,N_5350,N_5242);
xor U5596 (N_5596,N_5255,N_5235);
nand U5597 (N_5597,N_5294,N_5359);
nor U5598 (N_5598,N_5370,N_5208);
or U5599 (N_5599,N_5340,N_5200);
nor U5600 (N_5600,N_5544,N_5509);
or U5601 (N_5601,N_5554,N_5446);
or U5602 (N_5602,N_5481,N_5433);
and U5603 (N_5603,N_5489,N_5470);
nor U5604 (N_5604,N_5583,N_5573);
xor U5605 (N_5605,N_5469,N_5448);
nor U5606 (N_5606,N_5514,N_5474);
xor U5607 (N_5607,N_5464,N_5598);
nand U5608 (N_5608,N_5457,N_5571);
nand U5609 (N_5609,N_5528,N_5415);
and U5610 (N_5610,N_5599,N_5406);
or U5611 (N_5611,N_5404,N_5475);
nor U5612 (N_5612,N_5540,N_5531);
nand U5613 (N_5613,N_5451,N_5543);
and U5614 (N_5614,N_5494,N_5483);
nor U5615 (N_5615,N_5575,N_5566);
and U5616 (N_5616,N_5576,N_5513);
nand U5617 (N_5617,N_5527,N_5518);
and U5618 (N_5618,N_5577,N_5491);
nand U5619 (N_5619,N_5591,N_5560);
nor U5620 (N_5620,N_5520,N_5553);
nor U5621 (N_5621,N_5568,N_5542);
xnor U5622 (N_5622,N_5432,N_5449);
and U5623 (N_5623,N_5421,N_5480);
or U5624 (N_5624,N_5570,N_5442);
or U5625 (N_5625,N_5535,N_5594);
xor U5626 (N_5626,N_5502,N_5521);
nor U5627 (N_5627,N_5505,N_5403);
and U5628 (N_5628,N_5431,N_5556);
xnor U5629 (N_5629,N_5425,N_5596);
xnor U5630 (N_5630,N_5511,N_5471);
and U5631 (N_5631,N_5485,N_5492);
nand U5632 (N_5632,N_5487,N_5562);
nand U5633 (N_5633,N_5418,N_5557);
xnor U5634 (N_5634,N_5588,N_5525);
xor U5635 (N_5635,N_5472,N_5524);
or U5636 (N_5636,N_5538,N_5584);
and U5637 (N_5637,N_5461,N_5529);
xnor U5638 (N_5638,N_5532,N_5405);
xor U5639 (N_5639,N_5581,N_5586);
or U5640 (N_5640,N_5440,N_5417);
or U5641 (N_5641,N_5565,N_5507);
xnor U5642 (N_5642,N_5445,N_5547);
xnor U5643 (N_5643,N_5447,N_5597);
xnor U5644 (N_5644,N_5455,N_5467);
nand U5645 (N_5645,N_5443,N_5436);
nand U5646 (N_5646,N_5490,N_5468);
nand U5647 (N_5647,N_5437,N_5515);
or U5648 (N_5648,N_5408,N_5530);
nand U5649 (N_5649,N_5498,N_5508);
xnor U5650 (N_5650,N_5402,N_5574);
and U5651 (N_5651,N_5477,N_5559);
xnor U5652 (N_5652,N_5593,N_5587);
or U5653 (N_5653,N_5476,N_5595);
nand U5654 (N_5654,N_5579,N_5409);
xnor U5655 (N_5655,N_5541,N_5499);
nor U5656 (N_5656,N_5493,N_5428);
nand U5657 (N_5657,N_5567,N_5510);
or U5658 (N_5658,N_5504,N_5563);
and U5659 (N_5659,N_5426,N_5572);
or U5660 (N_5660,N_5463,N_5558);
nand U5661 (N_5661,N_5484,N_5454);
nor U5662 (N_5662,N_5512,N_5410);
nor U5663 (N_5663,N_5545,N_5400);
nand U5664 (N_5664,N_5533,N_5548);
xnor U5665 (N_5665,N_5439,N_5549);
nand U5666 (N_5666,N_5500,N_5479);
and U5667 (N_5667,N_5456,N_5424);
or U5668 (N_5668,N_5478,N_5427);
and U5669 (N_5669,N_5561,N_5430);
nand U5670 (N_5670,N_5420,N_5495);
nand U5671 (N_5671,N_5452,N_5522);
and U5672 (N_5672,N_5585,N_5552);
and U5673 (N_5673,N_5569,N_5555);
and U5674 (N_5674,N_5401,N_5429);
nand U5675 (N_5675,N_5416,N_5482);
and U5676 (N_5676,N_5496,N_5458);
and U5677 (N_5677,N_5501,N_5413);
and U5678 (N_5678,N_5460,N_5497);
or U5679 (N_5679,N_5592,N_5407);
or U5680 (N_5680,N_5590,N_5412);
xor U5681 (N_5681,N_5589,N_5434);
nor U5682 (N_5682,N_5546,N_5551);
or U5683 (N_5683,N_5486,N_5414);
and U5684 (N_5684,N_5450,N_5459);
nand U5685 (N_5685,N_5422,N_5488);
nand U5686 (N_5686,N_5419,N_5550);
or U5687 (N_5687,N_5539,N_5441);
and U5688 (N_5688,N_5444,N_5582);
or U5689 (N_5689,N_5465,N_5534);
or U5690 (N_5690,N_5503,N_5580);
or U5691 (N_5691,N_5578,N_5438);
nor U5692 (N_5692,N_5466,N_5523);
nand U5693 (N_5693,N_5526,N_5517);
nor U5694 (N_5694,N_5564,N_5506);
nor U5695 (N_5695,N_5516,N_5519);
nand U5696 (N_5696,N_5435,N_5537);
nor U5697 (N_5697,N_5453,N_5423);
and U5698 (N_5698,N_5473,N_5411);
nand U5699 (N_5699,N_5462,N_5536);
nand U5700 (N_5700,N_5407,N_5516);
or U5701 (N_5701,N_5511,N_5412);
xnor U5702 (N_5702,N_5467,N_5446);
and U5703 (N_5703,N_5466,N_5599);
xor U5704 (N_5704,N_5410,N_5459);
or U5705 (N_5705,N_5567,N_5591);
or U5706 (N_5706,N_5556,N_5529);
or U5707 (N_5707,N_5450,N_5412);
xor U5708 (N_5708,N_5435,N_5451);
and U5709 (N_5709,N_5480,N_5546);
nor U5710 (N_5710,N_5509,N_5576);
nand U5711 (N_5711,N_5453,N_5455);
xor U5712 (N_5712,N_5477,N_5452);
nor U5713 (N_5713,N_5462,N_5498);
nand U5714 (N_5714,N_5488,N_5423);
nand U5715 (N_5715,N_5451,N_5478);
nand U5716 (N_5716,N_5469,N_5582);
and U5717 (N_5717,N_5445,N_5564);
or U5718 (N_5718,N_5556,N_5485);
and U5719 (N_5719,N_5479,N_5507);
xor U5720 (N_5720,N_5583,N_5472);
or U5721 (N_5721,N_5509,N_5499);
or U5722 (N_5722,N_5512,N_5503);
nand U5723 (N_5723,N_5436,N_5508);
nor U5724 (N_5724,N_5581,N_5462);
xnor U5725 (N_5725,N_5454,N_5561);
xor U5726 (N_5726,N_5578,N_5473);
and U5727 (N_5727,N_5569,N_5453);
nand U5728 (N_5728,N_5522,N_5474);
nor U5729 (N_5729,N_5571,N_5545);
or U5730 (N_5730,N_5413,N_5499);
nor U5731 (N_5731,N_5482,N_5578);
xnor U5732 (N_5732,N_5491,N_5494);
and U5733 (N_5733,N_5534,N_5469);
and U5734 (N_5734,N_5481,N_5469);
or U5735 (N_5735,N_5586,N_5408);
nor U5736 (N_5736,N_5564,N_5565);
nand U5737 (N_5737,N_5449,N_5409);
nand U5738 (N_5738,N_5556,N_5543);
nand U5739 (N_5739,N_5528,N_5477);
xor U5740 (N_5740,N_5537,N_5409);
nor U5741 (N_5741,N_5598,N_5448);
nand U5742 (N_5742,N_5592,N_5564);
xor U5743 (N_5743,N_5466,N_5472);
nand U5744 (N_5744,N_5433,N_5558);
and U5745 (N_5745,N_5494,N_5473);
nor U5746 (N_5746,N_5447,N_5446);
and U5747 (N_5747,N_5560,N_5586);
nand U5748 (N_5748,N_5408,N_5546);
and U5749 (N_5749,N_5460,N_5421);
nor U5750 (N_5750,N_5592,N_5400);
xnor U5751 (N_5751,N_5458,N_5482);
nor U5752 (N_5752,N_5534,N_5585);
and U5753 (N_5753,N_5456,N_5563);
xnor U5754 (N_5754,N_5591,N_5436);
xor U5755 (N_5755,N_5427,N_5552);
xnor U5756 (N_5756,N_5493,N_5400);
xnor U5757 (N_5757,N_5541,N_5457);
nor U5758 (N_5758,N_5440,N_5563);
xor U5759 (N_5759,N_5511,N_5557);
nand U5760 (N_5760,N_5548,N_5519);
nor U5761 (N_5761,N_5501,N_5538);
and U5762 (N_5762,N_5436,N_5538);
nand U5763 (N_5763,N_5550,N_5570);
or U5764 (N_5764,N_5481,N_5547);
and U5765 (N_5765,N_5545,N_5526);
or U5766 (N_5766,N_5558,N_5513);
and U5767 (N_5767,N_5535,N_5579);
nand U5768 (N_5768,N_5585,N_5449);
xnor U5769 (N_5769,N_5501,N_5543);
nor U5770 (N_5770,N_5578,N_5531);
nand U5771 (N_5771,N_5447,N_5486);
xnor U5772 (N_5772,N_5434,N_5534);
nand U5773 (N_5773,N_5512,N_5588);
nand U5774 (N_5774,N_5424,N_5573);
or U5775 (N_5775,N_5546,N_5507);
nand U5776 (N_5776,N_5434,N_5484);
or U5777 (N_5777,N_5589,N_5429);
and U5778 (N_5778,N_5470,N_5501);
nor U5779 (N_5779,N_5530,N_5492);
nor U5780 (N_5780,N_5498,N_5554);
or U5781 (N_5781,N_5402,N_5428);
xor U5782 (N_5782,N_5589,N_5564);
xor U5783 (N_5783,N_5559,N_5439);
xor U5784 (N_5784,N_5418,N_5541);
and U5785 (N_5785,N_5565,N_5555);
and U5786 (N_5786,N_5401,N_5494);
nand U5787 (N_5787,N_5423,N_5536);
nor U5788 (N_5788,N_5472,N_5597);
xnor U5789 (N_5789,N_5486,N_5506);
nor U5790 (N_5790,N_5472,N_5422);
and U5791 (N_5791,N_5563,N_5579);
or U5792 (N_5792,N_5400,N_5578);
nand U5793 (N_5793,N_5491,N_5458);
nand U5794 (N_5794,N_5461,N_5499);
nand U5795 (N_5795,N_5498,N_5540);
or U5796 (N_5796,N_5597,N_5579);
nor U5797 (N_5797,N_5556,N_5434);
xor U5798 (N_5798,N_5454,N_5429);
xnor U5799 (N_5799,N_5486,N_5485);
or U5800 (N_5800,N_5744,N_5653);
nand U5801 (N_5801,N_5772,N_5778);
and U5802 (N_5802,N_5708,N_5659);
and U5803 (N_5803,N_5682,N_5685);
xor U5804 (N_5804,N_5738,N_5788);
xnor U5805 (N_5805,N_5748,N_5719);
or U5806 (N_5806,N_5775,N_5779);
and U5807 (N_5807,N_5794,N_5705);
nor U5808 (N_5808,N_5601,N_5619);
or U5809 (N_5809,N_5656,N_5605);
nand U5810 (N_5810,N_5782,N_5667);
nand U5811 (N_5811,N_5798,N_5650);
and U5812 (N_5812,N_5799,N_5690);
nor U5813 (N_5813,N_5683,N_5641);
nand U5814 (N_5814,N_5736,N_5628);
nand U5815 (N_5815,N_5696,N_5695);
nor U5816 (N_5816,N_5774,N_5612);
xnor U5817 (N_5817,N_5725,N_5675);
nand U5818 (N_5818,N_5634,N_5637);
or U5819 (N_5819,N_5604,N_5661);
xor U5820 (N_5820,N_5746,N_5686);
xor U5821 (N_5821,N_5723,N_5678);
xnor U5822 (N_5822,N_5743,N_5733);
or U5823 (N_5823,N_5711,N_5609);
nor U5824 (N_5824,N_5718,N_5726);
and U5825 (N_5825,N_5737,N_5669);
and U5826 (N_5826,N_5663,N_5734);
xnor U5827 (N_5827,N_5643,N_5728);
or U5828 (N_5828,N_5611,N_5654);
xnor U5829 (N_5829,N_5727,N_5707);
and U5830 (N_5830,N_5679,N_5632);
and U5831 (N_5831,N_5674,N_5765);
nor U5832 (N_5832,N_5739,N_5760);
and U5833 (N_5833,N_5730,N_5790);
nand U5834 (N_5834,N_5660,N_5614);
or U5835 (N_5835,N_5786,N_5729);
nand U5836 (N_5836,N_5664,N_5710);
xnor U5837 (N_5837,N_5703,N_5791);
nand U5838 (N_5838,N_5645,N_5780);
nor U5839 (N_5839,N_5768,N_5607);
xor U5840 (N_5840,N_5709,N_5750);
or U5841 (N_5841,N_5694,N_5714);
and U5842 (N_5842,N_5613,N_5668);
xnor U5843 (N_5843,N_5691,N_5702);
and U5844 (N_5844,N_5624,N_5783);
nor U5845 (N_5845,N_5745,N_5606);
xnor U5846 (N_5846,N_5716,N_5698);
or U5847 (N_5847,N_5647,N_5764);
or U5848 (N_5848,N_5701,N_5626);
and U5849 (N_5849,N_5700,N_5741);
nor U5850 (N_5850,N_5673,N_5642);
and U5851 (N_5851,N_5635,N_5681);
xnor U5852 (N_5852,N_5692,N_5740);
or U5853 (N_5853,N_5757,N_5697);
and U5854 (N_5854,N_5776,N_5610);
or U5855 (N_5855,N_5721,N_5680);
and U5856 (N_5856,N_5600,N_5639);
and U5857 (N_5857,N_5769,N_5758);
and U5858 (N_5858,N_5706,N_5704);
and U5859 (N_5859,N_5652,N_5648);
or U5860 (N_5860,N_5784,N_5658);
xnor U5861 (N_5861,N_5712,N_5785);
nand U5862 (N_5862,N_5753,N_5684);
and U5863 (N_5863,N_5602,N_5713);
xor U5864 (N_5864,N_5620,N_5603);
nor U5865 (N_5865,N_5636,N_5759);
and U5866 (N_5866,N_5781,N_5756);
xor U5867 (N_5867,N_5793,N_5724);
xor U5868 (N_5868,N_5671,N_5735);
xnor U5869 (N_5869,N_5665,N_5676);
nor U5870 (N_5870,N_5621,N_5762);
and U5871 (N_5871,N_5644,N_5770);
nor U5872 (N_5872,N_5715,N_5751);
or U5873 (N_5873,N_5731,N_5651);
and U5874 (N_5874,N_5689,N_5761);
and U5875 (N_5875,N_5655,N_5789);
nor U5876 (N_5876,N_5649,N_5638);
xnor U5877 (N_5877,N_5687,N_5699);
and U5878 (N_5878,N_5752,N_5693);
xor U5879 (N_5879,N_5795,N_5657);
xnor U5880 (N_5880,N_5732,N_5672);
and U5881 (N_5881,N_5742,N_5630);
nor U5882 (N_5882,N_5631,N_5767);
xnor U5883 (N_5883,N_5662,N_5771);
nand U5884 (N_5884,N_5777,N_5627);
or U5885 (N_5885,N_5720,N_5646);
nor U5886 (N_5886,N_5618,N_5677);
nand U5887 (N_5887,N_5670,N_5796);
xnor U5888 (N_5888,N_5787,N_5747);
nor U5889 (N_5889,N_5616,N_5623);
nor U5890 (N_5890,N_5722,N_5797);
xnor U5891 (N_5891,N_5608,N_5792);
or U5892 (N_5892,N_5625,N_5754);
and U5893 (N_5893,N_5666,N_5633);
xnor U5894 (N_5894,N_5615,N_5640);
xor U5895 (N_5895,N_5755,N_5688);
xor U5896 (N_5896,N_5629,N_5763);
or U5897 (N_5897,N_5773,N_5717);
nand U5898 (N_5898,N_5766,N_5622);
nand U5899 (N_5899,N_5617,N_5749);
or U5900 (N_5900,N_5709,N_5722);
and U5901 (N_5901,N_5756,N_5712);
and U5902 (N_5902,N_5663,N_5766);
xor U5903 (N_5903,N_5620,N_5792);
xnor U5904 (N_5904,N_5735,N_5631);
or U5905 (N_5905,N_5711,N_5748);
nand U5906 (N_5906,N_5637,N_5798);
nor U5907 (N_5907,N_5686,N_5784);
xor U5908 (N_5908,N_5614,N_5659);
nand U5909 (N_5909,N_5607,N_5619);
xor U5910 (N_5910,N_5673,N_5721);
nand U5911 (N_5911,N_5686,N_5612);
or U5912 (N_5912,N_5701,N_5681);
or U5913 (N_5913,N_5779,N_5788);
xor U5914 (N_5914,N_5618,N_5756);
xnor U5915 (N_5915,N_5750,N_5774);
and U5916 (N_5916,N_5742,N_5755);
nor U5917 (N_5917,N_5619,N_5655);
nor U5918 (N_5918,N_5672,N_5795);
xor U5919 (N_5919,N_5774,N_5745);
xor U5920 (N_5920,N_5687,N_5655);
xor U5921 (N_5921,N_5735,N_5721);
nand U5922 (N_5922,N_5645,N_5660);
nor U5923 (N_5923,N_5751,N_5669);
xor U5924 (N_5924,N_5769,N_5630);
and U5925 (N_5925,N_5654,N_5724);
xnor U5926 (N_5926,N_5717,N_5726);
nand U5927 (N_5927,N_5698,N_5618);
xor U5928 (N_5928,N_5621,N_5631);
and U5929 (N_5929,N_5624,N_5763);
nor U5930 (N_5930,N_5602,N_5785);
nor U5931 (N_5931,N_5694,N_5796);
nor U5932 (N_5932,N_5633,N_5745);
and U5933 (N_5933,N_5769,N_5783);
or U5934 (N_5934,N_5762,N_5695);
or U5935 (N_5935,N_5757,N_5705);
nand U5936 (N_5936,N_5765,N_5630);
and U5937 (N_5937,N_5791,N_5614);
or U5938 (N_5938,N_5690,N_5619);
xor U5939 (N_5939,N_5632,N_5684);
nand U5940 (N_5940,N_5763,N_5703);
and U5941 (N_5941,N_5663,N_5758);
nand U5942 (N_5942,N_5699,N_5605);
or U5943 (N_5943,N_5771,N_5609);
xnor U5944 (N_5944,N_5713,N_5629);
and U5945 (N_5945,N_5775,N_5613);
or U5946 (N_5946,N_5628,N_5767);
or U5947 (N_5947,N_5679,N_5647);
nand U5948 (N_5948,N_5613,N_5735);
and U5949 (N_5949,N_5654,N_5727);
or U5950 (N_5950,N_5754,N_5784);
or U5951 (N_5951,N_5636,N_5614);
xnor U5952 (N_5952,N_5648,N_5721);
and U5953 (N_5953,N_5796,N_5625);
or U5954 (N_5954,N_5660,N_5699);
xor U5955 (N_5955,N_5625,N_5779);
or U5956 (N_5956,N_5639,N_5740);
xor U5957 (N_5957,N_5779,N_5769);
and U5958 (N_5958,N_5784,N_5609);
xor U5959 (N_5959,N_5701,N_5779);
or U5960 (N_5960,N_5741,N_5709);
nand U5961 (N_5961,N_5771,N_5698);
or U5962 (N_5962,N_5613,N_5649);
xor U5963 (N_5963,N_5623,N_5685);
and U5964 (N_5964,N_5697,N_5767);
and U5965 (N_5965,N_5758,N_5797);
nand U5966 (N_5966,N_5730,N_5658);
or U5967 (N_5967,N_5761,N_5620);
or U5968 (N_5968,N_5633,N_5629);
or U5969 (N_5969,N_5707,N_5691);
nor U5970 (N_5970,N_5636,N_5768);
nand U5971 (N_5971,N_5691,N_5607);
or U5972 (N_5972,N_5718,N_5765);
xor U5973 (N_5973,N_5663,N_5732);
or U5974 (N_5974,N_5628,N_5787);
nor U5975 (N_5975,N_5699,N_5763);
and U5976 (N_5976,N_5789,N_5712);
or U5977 (N_5977,N_5601,N_5628);
and U5978 (N_5978,N_5634,N_5728);
nand U5979 (N_5979,N_5794,N_5648);
xor U5980 (N_5980,N_5652,N_5692);
xor U5981 (N_5981,N_5620,N_5772);
or U5982 (N_5982,N_5704,N_5792);
or U5983 (N_5983,N_5778,N_5635);
nor U5984 (N_5984,N_5693,N_5785);
nand U5985 (N_5985,N_5745,N_5746);
nand U5986 (N_5986,N_5682,N_5749);
or U5987 (N_5987,N_5720,N_5617);
and U5988 (N_5988,N_5731,N_5639);
xor U5989 (N_5989,N_5600,N_5652);
or U5990 (N_5990,N_5666,N_5629);
xnor U5991 (N_5991,N_5774,N_5708);
and U5992 (N_5992,N_5782,N_5776);
nand U5993 (N_5993,N_5735,N_5703);
nor U5994 (N_5994,N_5759,N_5796);
or U5995 (N_5995,N_5742,N_5617);
xnor U5996 (N_5996,N_5703,N_5779);
nor U5997 (N_5997,N_5627,N_5723);
xor U5998 (N_5998,N_5754,N_5761);
or U5999 (N_5999,N_5795,N_5768);
and U6000 (N_6000,N_5866,N_5925);
and U6001 (N_6001,N_5966,N_5935);
xor U6002 (N_6002,N_5850,N_5950);
nand U6003 (N_6003,N_5881,N_5937);
xnor U6004 (N_6004,N_5807,N_5914);
nor U6005 (N_6005,N_5823,N_5969);
nand U6006 (N_6006,N_5913,N_5974);
nor U6007 (N_6007,N_5855,N_5803);
nand U6008 (N_6008,N_5890,N_5951);
xor U6009 (N_6009,N_5865,N_5957);
xnor U6010 (N_6010,N_5814,N_5897);
nor U6011 (N_6011,N_5856,N_5845);
nor U6012 (N_6012,N_5980,N_5987);
xor U6013 (N_6013,N_5992,N_5903);
and U6014 (N_6014,N_5922,N_5862);
xor U6015 (N_6015,N_5820,N_5843);
nand U6016 (N_6016,N_5811,N_5996);
xor U6017 (N_6017,N_5822,N_5800);
nor U6018 (N_6018,N_5841,N_5930);
nor U6019 (N_6019,N_5839,N_5967);
nand U6020 (N_6020,N_5977,N_5805);
and U6021 (N_6021,N_5812,N_5932);
xor U6022 (N_6022,N_5829,N_5946);
nand U6023 (N_6023,N_5864,N_5892);
nand U6024 (N_6024,N_5896,N_5886);
nand U6025 (N_6025,N_5982,N_5885);
nand U6026 (N_6026,N_5947,N_5934);
nor U6027 (N_6027,N_5875,N_5810);
xnor U6028 (N_6028,N_5817,N_5834);
and U6029 (N_6029,N_5975,N_5943);
xnor U6030 (N_6030,N_5861,N_5906);
nand U6031 (N_6031,N_5952,N_5835);
or U6032 (N_6032,N_5883,N_5920);
nor U6033 (N_6033,N_5824,N_5859);
or U6034 (N_6034,N_5877,N_5899);
nor U6035 (N_6035,N_5876,N_5954);
nand U6036 (N_6036,N_5942,N_5918);
nor U6037 (N_6037,N_5962,N_5851);
nand U6038 (N_6038,N_5905,N_5979);
nor U6039 (N_6039,N_5915,N_5888);
xor U6040 (N_6040,N_5832,N_5878);
and U6041 (N_6041,N_5898,N_5808);
xnor U6042 (N_6042,N_5928,N_5959);
xor U6043 (N_6043,N_5840,N_5821);
nor U6044 (N_6044,N_5926,N_5860);
nor U6045 (N_6045,N_5804,N_5911);
and U6046 (N_6046,N_5801,N_5872);
xor U6047 (N_6047,N_5924,N_5844);
nor U6048 (N_6048,N_5940,N_5816);
and U6049 (N_6049,N_5830,N_5931);
or U6050 (N_6050,N_5993,N_5893);
and U6051 (N_6051,N_5884,N_5880);
and U6052 (N_6052,N_5868,N_5994);
nor U6053 (N_6053,N_5904,N_5852);
and U6054 (N_6054,N_5981,N_5846);
and U6055 (N_6055,N_5964,N_5983);
nand U6056 (N_6056,N_5939,N_5976);
xnor U6057 (N_6057,N_5825,N_5986);
or U6058 (N_6058,N_5857,N_5978);
and U6059 (N_6059,N_5900,N_5916);
nand U6060 (N_6060,N_5960,N_5863);
nand U6061 (N_6061,N_5972,N_5889);
nor U6062 (N_6062,N_5827,N_5985);
or U6063 (N_6063,N_5813,N_5910);
xor U6064 (N_6064,N_5945,N_5956);
or U6065 (N_6065,N_5988,N_5984);
xor U6066 (N_6066,N_5815,N_5948);
nor U6067 (N_6067,N_5887,N_5891);
nor U6068 (N_6068,N_5873,N_5949);
and U6069 (N_6069,N_5895,N_5867);
nand U6070 (N_6070,N_5936,N_5995);
xnor U6071 (N_6071,N_5858,N_5991);
and U6072 (N_6072,N_5836,N_5809);
or U6073 (N_6073,N_5842,N_5837);
or U6074 (N_6074,N_5963,N_5912);
nor U6075 (N_6075,N_5938,N_5879);
and U6076 (N_6076,N_5849,N_5802);
nand U6077 (N_6077,N_5908,N_5848);
nand U6078 (N_6078,N_5944,N_5970);
nand U6079 (N_6079,N_5933,N_5869);
nand U6080 (N_6080,N_5941,N_5917);
xor U6081 (N_6081,N_5958,N_5971);
or U6082 (N_6082,N_5882,N_5965);
and U6083 (N_6083,N_5894,N_5997);
and U6084 (N_6084,N_5874,N_5989);
nand U6085 (N_6085,N_5973,N_5831);
nor U6086 (N_6086,N_5909,N_5919);
nand U6087 (N_6087,N_5907,N_5923);
or U6088 (N_6088,N_5833,N_5853);
and U6089 (N_6089,N_5838,N_5901);
and U6090 (N_6090,N_5921,N_5854);
and U6091 (N_6091,N_5929,N_5998);
xnor U6092 (N_6092,N_5902,N_5847);
xnor U6093 (N_6093,N_5999,N_5818);
and U6094 (N_6094,N_5968,N_5927);
nand U6095 (N_6095,N_5961,N_5828);
or U6096 (N_6096,N_5871,N_5870);
nor U6097 (N_6097,N_5806,N_5819);
nand U6098 (N_6098,N_5826,N_5953);
nand U6099 (N_6099,N_5990,N_5955);
nand U6100 (N_6100,N_5816,N_5829);
xnor U6101 (N_6101,N_5875,N_5863);
nor U6102 (N_6102,N_5844,N_5809);
and U6103 (N_6103,N_5854,N_5823);
and U6104 (N_6104,N_5917,N_5998);
xor U6105 (N_6105,N_5909,N_5817);
nor U6106 (N_6106,N_5905,N_5947);
nor U6107 (N_6107,N_5921,N_5897);
or U6108 (N_6108,N_5865,N_5999);
or U6109 (N_6109,N_5855,N_5889);
or U6110 (N_6110,N_5938,N_5952);
or U6111 (N_6111,N_5852,N_5840);
nor U6112 (N_6112,N_5926,N_5952);
xor U6113 (N_6113,N_5821,N_5816);
and U6114 (N_6114,N_5834,N_5854);
nor U6115 (N_6115,N_5817,N_5866);
or U6116 (N_6116,N_5829,N_5896);
nand U6117 (N_6117,N_5872,N_5922);
nand U6118 (N_6118,N_5965,N_5826);
nand U6119 (N_6119,N_5941,N_5973);
xnor U6120 (N_6120,N_5980,N_5854);
nand U6121 (N_6121,N_5987,N_5958);
nor U6122 (N_6122,N_5953,N_5906);
xnor U6123 (N_6123,N_5998,N_5944);
and U6124 (N_6124,N_5829,N_5952);
nand U6125 (N_6125,N_5821,N_5893);
xor U6126 (N_6126,N_5980,N_5992);
and U6127 (N_6127,N_5825,N_5823);
and U6128 (N_6128,N_5927,N_5813);
and U6129 (N_6129,N_5894,N_5972);
nor U6130 (N_6130,N_5870,N_5876);
nor U6131 (N_6131,N_5904,N_5894);
nor U6132 (N_6132,N_5904,N_5859);
xnor U6133 (N_6133,N_5819,N_5896);
nand U6134 (N_6134,N_5836,N_5973);
nand U6135 (N_6135,N_5963,N_5942);
nor U6136 (N_6136,N_5936,N_5961);
and U6137 (N_6137,N_5912,N_5910);
and U6138 (N_6138,N_5907,N_5862);
and U6139 (N_6139,N_5874,N_5985);
or U6140 (N_6140,N_5849,N_5928);
xor U6141 (N_6141,N_5812,N_5925);
nor U6142 (N_6142,N_5870,N_5923);
xnor U6143 (N_6143,N_5917,N_5950);
nor U6144 (N_6144,N_5804,N_5887);
nand U6145 (N_6145,N_5841,N_5864);
and U6146 (N_6146,N_5801,N_5933);
nand U6147 (N_6147,N_5976,N_5913);
nor U6148 (N_6148,N_5973,N_5875);
nand U6149 (N_6149,N_5891,N_5859);
nand U6150 (N_6150,N_5993,N_5859);
nand U6151 (N_6151,N_5895,N_5953);
xnor U6152 (N_6152,N_5803,N_5952);
or U6153 (N_6153,N_5857,N_5947);
nor U6154 (N_6154,N_5966,N_5849);
and U6155 (N_6155,N_5944,N_5839);
nor U6156 (N_6156,N_5834,N_5966);
and U6157 (N_6157,N_5851,N_5965);
nor U6158 (N_6158,N_5867,N_5868);
and U6159 (N_6159,N_5907,N_5885);
nor U6160 (N_6160,N_5912,N_5823);
and U6161 (N_6161,N_5961,N_5935);
or U6162 (N_6162,N_5931,N_5966);
nor U6163 (N_6163,N_5930,N_5924);
xor U6164 (N_6164,N_5911,N_5891);
xnor U6165 (N_6165,N_5818,N_5833);
xnor U6166 (N_6166,N_5820,N_5921);
nand U6167 (N_6167,N_5827,N_5971);
or U6168 (N_6168,N_5917,N_5967);
and U6169 (N_6169,N_5821,N_5972);
nand U6170 (N_6170,N_5934,N_5836);
nor U6171 (N_6171,N_5973,N_5835);
xor U6172 (N_6172,N_5844,N_5855);
nand U6173 (N_6173,N_5831,N_5828);
xor U6174 (N_6174,N_5952,N_5985);
xor U6175 (N_6175,N_5955,N_5860);
nand U6176 (N_6176,N_5963,N_5924);
or U6177 (N_6177,N_5918,N_5978);
xnor U6178 (N_6178,N_5841,N_5803);
nor U6179 (N_6179,N_5991,N_5826);
nor U6180 (N_6180,N_5969,N_5942);
xor U6181 (N_6181,N_5981,N_5908);
nor U6182 (N_6182,N_5872,N_5995);
nand U6183 (N_6183,N_5930,N_5949);
nor U6184 (N_6184,N_5936,N_5902);
nor U6185 (N_6185,N_5965,N_5801);
and U6186 (N_6186,N_5850,N_5817);
xor U6187 (N_6187,N_5937,N_5853);
nor U6188 (N_6188,N_5907,N_5846);
xor U6189 (N_6189,N_5966,N_5840);
and U6190 (N_6190,N_5898,N_5935);
nor U6191 (N_6191,N_5812,N_5857);
nor U6192 (N_6192,N_5874,N_5926);
nor U6193 (N_6193,N_5829,N_5944);
nor U6194 (N_6194,N_5969,N_5848);
nor U6195 (N_6195,N_5954,N_5902);
nor U6196 (N_6196,N_5865,N_5843);
xnor U6197 (N_6197,N_5843,N_5841);
or U6198 (N_6198,N_5961,N_5844);
and U6199 (N_6199,N_5905,N_5836);
or U6200 (N_6200,N_6181,N_6087);
nand U6201 (N_6201,N_6066,N_6047);
nand U6202 (N_6202,N_6184,N_6013);
xnor U6203 (N_6203,N_6045,N_6086);
xor U6204 (N_6204,N_6142,N_6058);
nand U6205 (N_6205,N_6146,N_6077);
or U6206 (N_6206,N_6057,N_6010);
nand U6207 (N_6207,N_6129,N_6117);
xnor U6208 (N_6208,N_6056,N_6133);
or U6209 (N_6209,N_6051,N_6131);
nand U6210 (N_6210,N_6007,N_6093);
nor U6211 (N_6211,N_6016,N_6062);
nand U6212 (N_6212,N_6178,N_6120);
nor U6213 (N_6213,N_6179,N_6116);
nand U6214 (N_6214,N_6174,N_6011);
xor U6215 (N_6215,N_6065,N_6055);
or U6216 (N_6216,N_6031,N_6143);
and U6217 (N_6217,N_6180,N_6199);
and U6218 (N_6218,N_6027,N_6028);
xnor U6219 (N_6219,N_6072,N_6134);
xor U6220 (N_6220,N_6194,N_6132);
nor U6221 (N_6221,N_6170,N_6046);
nor U6222 (N_6222,N_6126,N_6138);
xor U6223 (N_6223,N_6118,N_6036);
nand U6224 (N_6224,N_6030,N_6003);
or U6225 (N_6225,N_6006,N_6145);
or U6226 (N_6226,N_6149,N_6019);
or U6227 (N_6227,N_6157,N_6043);
nor U6228 (N_6228,N_6033,N_6196);
xor U6229 (N_6229,N_6122,N_6192);
nor U6230 (N_6230,N_6035,N_6082);
xor U6231 (N_6231,N_6139,N_6026);
or U6232 (N_6232,N_6037,N_6067);
nor U6233 (N_6233,N_6048,N_6171);
or U6234 (N_6234,N_6154,N_6012);
nand U6235 (N_6235,N_6063,N_6130);
or U6236 (N_6236,N_6023,N_6156);
and U6237 (N_6237,N_6081,N_6024);
nor U6238 (N_6238,N_6085,N_6075);
nor U6239 (N_6239,N_6014,N_6177);
and U6240 (N_6240,N_6095,N_6176);
or U6241 (N_6241,N_6042,N_6106);
nor U6242 (N_6242,N_6197,N_6161);
nand U6243 (N_6243,N_6071,N_6061);
xor U6244 (N_6244,N_6034,N_6185);
and U6245 (N_6245,N_6108,N_6152);
or U6246 (N_6246,N_6115,N_6096);
or U6247 (N_6247,N_6005,N_6104);
nand U6248 (N_6248,N_6070,N_6092);
xnor U6249 (N_6249,N_6148,N_6008);
and U6250 (N_6250,N_6069,N_6080);
or U6251 (N_6251,N_6160,N_6105);
or U6252 (N_6252,N_6136,N_6128);
nor U6253 (N_6253,N_6172,N_6187);
or U6254 (N_6254,N_6103,N_6173);
nor U6255 (N_6255,N_6074,N_6041);
xor U6256 (N_6256,N_6083,N_6021);
and U6257 (N_6257,N_6137,N_6091);
and U6258 (N_6258,N_6064,N_6110);
xnor U6259 (N_6259,N_6119,N_6114);
nand U6260 (N_6260,N_6165,N_6166);
nand U6261 (N_6261,N_6112,N_6127);
xnor U6262 (N_6262,N_6076,N_6052);
xnor U6263 (N_6263,N_6102,N_6191);
xor U6264 (N_6264,N_6100,N_6125);
and U6265 (N_6265,N_6101,N_6000);
and U6266 (N_6266,N_6195,N_6001);
nand U6267 (N_6267,N_6140,N_6169);
or U6268 (N_6268,N_6113,N_6162);
nor U6269 (N_6269,N_6094,N_6060);
and U6270 (N_6270,N_6109,N_6153);
xnor U6271 (N_6271,N_6098,N_6078);
or U6272 (N_6272,N_6032,N_6059);
or U6273 (N_6273,N_6039,N_6015);
and U6274 (N_6274,N_6099,N_6189);
xor U6275 (N_6275,N_6004,N_6159);
or U6276 (N_6276,N_6017,N_6188);
or U6277 (N_6277,N_6135,N_6124);
nand U6278 (N_6278,N_6089,N_6123);
nor U6279 (N_6279,N_6022,N_6088);
and U6280 (N_6280,N_6147,N_6155);
nand U6281 (N_6281,N_6025,N_6038);
or U6282 (N_6282,N_6029,N_6164);
or U6283 (N_6283,N_6018,N_6198);
nor U6284 (N_6284,N_6054,N_6193);
or U6285 (N_6285,N_6097,N_6111);
nor U6286 (N_6286,N_6079,N_6158);
nor U6287 (N_6287,N_6163,N_6053);
nor U6288 (N_6288,N_6020,N_6141);
xnor U6289 (N_6289,N_6167,N_6049);
and U6290 (N_6290,N_6182,N_6190);
or U6291 (N_6291,N_6150,N_6183);
nand U6292 (N_6292,N_6168,N_6151);
and U6293 (N_6293,N_6121,N_6073);
nand U6294 (N_6294,N_6040,N_6107);
or U6295 (N_6295,N_6068,N_6144);
xor U6296 (N_6296,N_6084,N_6090);
nand U6297 (N_6297,N_6002,N_6050);
nand U6298 (N_6298,N_6009,N_6175);
or U6299 (N_6299,N_6044,N_6186);
and U6300 (N_6300,N_6009,N_6092);
nor U6301 (N_6301,N_6190,N_6026);
nand U6302 (N_6302,N_6092,N_6121);
or U6303 (N_6303,N_6052,N_6015);
nand U6304 (N_6304,N_6070,N_6029);
nand U6305 (N_6305,N_6155,N_6003);
nor U6306 (N_6306,N_6133,N_6071);
nor U6307 (N_6307,N_6108,N_6076);
xnor U6308 (N_6308,N_6000,N_6056);
or U6309 (N_6309,N_6057,N_6168);
xnor U6310 (N_6310,N_6041,N_6114);
nor U6311 (N_6311,N_6140,N_6015);
nor U6312 (N_6312,N_6093,N_6006);
xor U6313 (N_6313,N_6170,N_6086);
nor U6314 (N_6314,N_6014,N_6149);
or U6315 (N_6315,N_6024,N_6183);
and U6316 (N_6316,N_6077,N_6117);
nor U6317 (N_6317,N_6047,N_6081);
or U6318 (N_6318,N_6043,N_6122);
or U6319 (N_6319,N_6160,N_6087);
xor U6320 (N_6320,N_6002,N_6018);
nand U6321 (N_6321,N_6119,N_6194);
xnor U6322 (N_6322,N_6170,N_6045);
nor U6323 (N_6323,N_6011,N_6117);
nor U6324 (N_6324,N_6050,N_6156);
nand U6325 (N_6325,N_6029,N_6156);
and U6326 (N_6326,N_6095,N_6138);
xor U6327 (N_6327,N_6087,N_6089);
xor U6328 (N_6328,N_6136,N_6096);
nand U6329 (N_6329,N_6064,N_6057);
nor U6330 (N_6330,N_6196,N_6041);
nand U6331 (N_6331,N_6018,N_6042);
nand U6332 (N_6332,N_6033,N_6015);
and U6333 (N_6333,N_6030,N_6117);
or U6334 (N_6334,N_6103,N_6016);
xor U6335 (N_6335,N_6132,N_6054);
or U6336 (N_6336,N_6124,N_6012);
or U6337 (N_6337,N_6024,N_6006);
nor U6338 (N_6338,N_6111,N_6126);
nor U6339 (N_6339,N_6011,N_6032);
nor U6340 (N_6340,N_6168,N_6136);
xor U6341 (N_6341,N_6132,N_6020);
and U6342 (N_6342,N_6051,N_6163);
or U6343 (N_6343,N_6085,N_6058);
xnor U6344 (N_6344,N_6075,N_6035);
xor U6345 (N_6345,N_6124,N_6142);
nor U6346 (N_6346,N_6044,N_6154);
and U6347 (N_6347,N_6083,N_6188);
nand U6348 (N_6348,N_6186,N_6185);
xor U6349 (N_6349,N_6071,N_6005);
and U6350 (N_6350,N_6070,N_6050);
xor U6351 (N_6351,N_6059,N_6016);
xor U6352 (N_6352,N_6011,N_6183);
xnor U6353 (N_6353,N_6188,N_6180);
nor U6354 (N_6354,N_6124,N_6033);
and U6355 (N_6355,N_6004,N_6165);
or U6356 (N_6356,N_6101,N_6159);
and U6357 (N_6357,N_6127,N_6189);
nand U6358 (N_6358,N_6008,N_6108);
nand U6359 (N_6359,N_6189,N_6148);
nand U6360 (N_6360,N_6129,N_6199);
xnor U6361 (N_6361,N_6039,N_6043);
or U6362 (N_6362,N_6072,N_6148);
nor U6363 (N_6363,N_6046,N_6145);
nor U6364 (N_6364,N_6089,N_6171);
nor U6365 (N_6365,N_6150,N_6090);
nand U6366 (N_6366,N_6154,N_6069);
and U6367 (N_6367,N_6103,N_6124);
or U6368 (N_6368,N_6168,N_6144);
nor U6369 (N_6369,N_6112,N_6077);
nand U6370 (N_6370,N_6106,N_6086);
xnor U6371 (N_6371,N_6169,N_6173);
or U6372 (N_6372,N_6144,N_6119);
xor U6373 (N_6373,N_6035,N_6051);
nor U6374 (N_6374,N_6173,N_6123);
or U6375 (N_6375,N_6002,N_6081);
or U6376 (N_6376,N_6020,N_6187);
nor U6377 (N_6377,N_6121,N_6094);
xor U6378 (N_6378,N_6175,N_6013);
nor U6379 (N_6379,N_6005,N_6073);
nor U6380 (N_6380,N_6183,N_6081);
and U6381 (N_6381,N_6090,N_6028);
nand U6382 (N_6382,N_6197,N_6048);
or U6383 (N_6383,N_6036,N_6032);
and U6384 (N_6384,N_6044,N_6189);
nand U6385 (N_6385,N_6075,N_6007);
xnor U6386 (N_6386,N_6131,N_6070);
or U6387 (N_6387,N_6020,N_6180);
or U6388 (N_6388,N_6172,N_6100);
and U6389 (N_6389,N_6191,N_6080);
xnor U6390 (N_6390,N_6004,N_6132);
nor U6391 (N_6391,N_6032,N_6126);
xnor U6392 (N_6392,N_6183,N_6192);
or U6393 (N_6393,N_6031,N_6026);
xor U6394 (N_6394,N_6147,N_6126);
and U6395 (N_6395,N_6174,N_6018);
xnor U6396 (N_6396,N_6082,N_6023);
and U6397 (N_6397,N_6049,N_6138);
or U6398 (N_6398,N_6169,N_6048);
nor U6399 (N_6399,N_6034,N_6138);
nor U6400 (N_6400,N_6220,N_6347);
nor U6401 (N_6401,N_6263,N_6283);
xnor U6402 (N_6402,N_6341,N_6296);
nand U6403 (N_6403,N_6392,N_6289);
and U6404 (N_6404,N_6333,N_6364);
nor U6405 (N_6405,N_6367,N_6250);
xnor U6406 (N_6406,N_6264,N_6348);
nand U6407 (N_6407,N_6397,N_6211);
xnor U6408 (N_6408,N_6226,N_6320);
and U6409 (N_6409,N_6329,N_6368);
xnor U6410 (N_6410,N_6342,N_6370);
or U6411 (N_6411,N_6282,N_6291);
and U6412 (N_6412,N_6277,N_6349);
and U6413 (N_6413,N_6233,N_6378);
or U6414 (N_6414,N_6396,N_6390);
xnor U6415 (N_6415,N_6243,N_6350);
or U6416 (N_6416,N_6253,N_6212);
xor U6417 (N_6417,N_6269,N_6223);
and U6418 (N_6418,N_6302,N_6251);
nand U6419 (N_6419,N_6351,N_6389);
nand U6420 (N_6420,N_6280,N_6312);
xor U6421 (N_6421,N_6391,N_6340);
or U6422 (N_6422,N_6356,N_6395);
xnor U6423 (N_6423,N_6319,N_6361);
and U6424 (N_6424,N_6228,N_6377);
xor U6425 (N_6425,N_6240,N_6380);
xor U6426 (N_6426,N_6295,N_6248);
nand U6427 (N_6427,N_6242,N_6239);
and U6428 (N_6428,N_6245,N_6262);
nor U6429 (N_6429,N_6306,N_6357);
xnor U6430 (N_6430,N_6308,N_6343);
and U6431 (N_6431,N_6304,N_6209);
or U6432 (N_6432,N_6215,N_6275);
nor U6433 (N_6433,N_6241,N_6274);
nor U6434 (N_6434,N_6288,N_6205);
and U6435 (N_6435,N_6388,N_6322);
xnor U6436 (N_6436,N_6303,N_6297);
or U6437 (N_6437,N_6221,N_6258);
or U6438 (N_6438,N_6214,N_6399);
nor U6439 (N_6439,N_6252,N_6309);
or U6440 (N_6440,N_6246,N_6284);
xor U6441 (N_6441,N_6267,N_6244);
nor U6442 (N_6442,N_6344,N_6373);
nor U6443 (N_6443,N_6227,N_6363);
xor U6444 (N_6444,N_6270,N_6318);
nand U6445 (N_6445,N_6316,N_6383);
and U6446 (N_6446,N_6210,N_6225);
nor U6447 (N_6447,N_6379,N_6256);
xor U6448 (N_6448,N_6324,N_6305);
xnor U6449 (N_6449,N_6265,N_6235);
xor U6450 (N_6450,N_6268,N_6247);
xnor U6451 (N_6451,N_6224,N_6230);
or U6452 (N_6452,N_6332,N_6217);
xnor U6453 (N_6453,N_6384,N_6328);
and U6454 (N_6454,N_6371,N_6381);
nand U6455 (N_6455,N_6337,N_6293);
and U6456 (N_6456,N_6259,N_6339);
and U6457 (N_6457,N_6327,N_6234);
xnor U6458 (N_6458,N_6208,N_6229);
xor U6459 (N_6459,N_6354,N_6294);
nor U6460 (N_6460,N_6300,N_6352);
nand U6461 (N_6461,N_6206,N_6260);
and U6462 (N_6462,N_6355,N_6375);
nor U6463 (N_6463,N_6201,N_6372);
nor U6464 (N_6464,N_6310,N_6271);
nor U6465 (N_6465,N_6386,N_6307);
nand U6466 (N_6466,N_6299,N_6231);
nor U6467 (N_6467,N_6353,N_6285);
xnor U6468 (N_6468,N_6362,N_6338);
nand U6469 (N_6469,N_6336,N_6279);
nor U6470 (N_6470,N_6382,N_6222);
xnor U6471 (N_6471,N_6236,N_6330);
xor U6472 (N_6472,N_6281,N_6323);
xor U6473 (N_6473,N_6276,N_6387);
and U6474 (N_6474,N_6237,N_6232);
or U6475 (N_6475,N_6272,N_6257);
nand U6476 (N_6476,N_6207,N_6202);
or U6477 (N_6477,N_6331,N_6358);
or U6478 (N_6478,N_6334,N_6314);
xor U6479 (N_6479,N_6266,N_6286);
and U6480 (N_6480,N_6398,N_6326);
nand U6481 (N_6481,N_6345,N_6366);
nand U6482 (N_6482,N_6219,N_6360);
nand U6483 (N_6483,N_6321,N_6385);
or U6484 (N_6484,N_6216,N_6273);
and U6485 (N_6485,N_6255,N_6369);
and U6486 (N_6486,N_6204,N_6365);
nand U6487 (N_6487,N_6317,N_6249);
or U6488 (N_6488,N_6301,N_6374);
nand U6489 (N_6489,N_6203,N_6292);
and U6490 (N_6490,N_6238,N_6287);
xor U6491 (N_6491,N_6254,N_6313);
xnor U6492 (N_6492,N_6376,N_6200);
or U6493 (N_6493,N_6335,N_6290);
or U6494 (N_6494,N_6325,N_6298);
xnor U6495 (N_6495,N_6213,N_6315);
xnor U6496 (N_6496,N_6311,N_6218);
or U6497 (N_6497,N_6394,N_6346);
xor U6498 (N_6498,N_6393,N_6278);
xor U6499 (N_6499,N_6261,N_6359);
nand U6500 (N_6500,N_6281,N_6239);
nor U6501 (N_6501,N_6247,N_6287);
xor U6502 (N_6502,N_6322,N_6239);
nand U6503 (N_6503,N_6324,N_6212);
nand U6504 (N_6504,N_6344,N_6294);
nand U6505 (N_6505,N_6243,N_6349);
nand U6506 (N_6506,N_6257,N_6219);
nand U6507 (N_6507,N_6208,N_6246);
and U6508 (N_6508,N_6343,N_6277);
xnor U6509 (N_6509,N_6363,N_6221);
and U6510 (N_6510,N_6300,N_6345);
nor U6511 (N_6511,N_6217,N_6297);
or U6512 (N_6512,N_6300,N_6368);
and U6513 (N_6513,N_6295,N_6353);
or U6514 (N_6514,N_6242,N_6311);
nor U6515 (N_6515,N_6364,N_6273);
nand U6516 (N_6516,N_6235,N_6346);
nor U6517 (N_6517,N_6351,N_6356);
and U6518 (N_6518,N_6344,N_6253);
xor U6519 (N_6519,N_6282,N_6200);
nand U6520 (N_6520,N_6226,N_6259);
and U6521 (N_6521,N_6295,N_6370);
nor U6522 (N_6522,N_6378,N_6392);
nor U6523 (N_6523,N_6287,N_6362);
nand U6524 (N_6524,N_6326,N_6272);
and U6525 (N_6525,N_6346,N_6203);
xor U6526 (N_6526,N_6378,N_6298);
or U6527 (N_6527,N_6370,N_6364);
nand U6528 (N_6528,N_6310,N_6344);
xnor U6529 (N_6529,N_6292,N_6209);
nor U6530 (N_6530,N_6333,N_6358);
or U6531 (N_6531,N_6386,N_6290);
xnor U6532 (N_6532,N_6234,N_6233);
nor U6533 (N_6533,N_6283,N_6233);
nand U6534 (N_6534,N_6278,N_6334);
nor U6535 (N_6535,N_6232,N_6286);
xnor U6536 (N_6536,N_6370,N_6222);
and U6537 (N_6537,N_6377,N_6309);
nand U6538 (N_6538,N_6387,N_6229);
xor U6539 (N_6539,N_6335,N_6377);
xor U6540 (N_6540,N_6303,N_6219);
xnor U6541 (N_6541,N_6242,N_6258);
nand U6542 (N_6542,N_6235,N_6224);
or U6543 (N_6543,N_6337,N_6360);
nor U6544 (N_6544,N_6333,N_6276);
nand U6545 (N_6545,N_6213,N_6365);
nand U6546 (N_6546,N_6315,N_6306);
xnor U6547 (N_6547,N_6256,N_6305);
and U6548 (N_6548,N_6253,N_6269);
and U6549 (N_6549,N_6237,N_6358);
or U6550 (N_6550,N_6346,N_6338);
and U6551 (N_6551,N_6364,N_6298);
xor U6552 (N_6552,N_6303,N_6213);
nor U6553 (N_6553,N_6344,N_6356);
nor U6554 (N_6554,N_6218,N_6233);
and U6555 (N_6555,N_6335,N_6256);
and U6556 (N_6556,N_6201,N_6304);
or U6557 (N_6557,N_6277,N_6352);
or U6558 (N_6558,N_6360,N_6287);
xnor U6559 (N_6559,N_6352,N_6227);
and U6560 (N_6560,N_6223,N_6300);
nand U6561 (N_6561,N_6249,N_6224);
nand U6562 (N_6562,N_6297,N_6347);
and U6563 (N_6563,N_6288,N_6255);
and U6564 (N_6564,N_6267,N_6305);
or U6565 (N_6565,N_6235,N_6276);
nor U6566 (N_6566,N_6277,N_6212);
nand U6567 (N_6567,N_6237,N_6254);
or U6568 (N_6568,N_6215,N_6290);
and U6569 (N_6569,N_6244,N_6211);
or U6570 (N_6570,N_6358,N_6284);
nor U6571 (N_6571,N_6307,N_6244);
or U6572 (N_6572,N_6290,N_6316);
nand U6573 (N_6573,N_6332,N_6286);
nor U6574 (N_6574,N_6283,N_6385);
and U6575 (N_6575,N_6293,N_6332);
and U6576 (N_6576,N_6245,N_6296);
or U6577 (N_6577,N_6306,N_6390);
xnor U6578 (N_6578,N_6217,N_6325);
nor U6579 (N_6579,N_6265,N_6294);
nand U6580 (N_6580,N_6271,N_6327);
nor U6581 (N_6581,N_6247,N_6386);
nor U6582 (N_6582,N_6289,N_6280);
or U6583 (N_6583,N_6217,N_6223);
nand U6584 (N_6584,N_6306,N_6260);
nor U6585 (N_6585,N_6271,N_6247);
or U6586 (N_6586,N_6378,N_6265);
nor U6587 (N_6587,N_6368,N_6226);
and U6588 (N_6588,N_6204,N_6266);
nor U6589 (N_6589,N_6390,N_6265);
or U6590 (N_6590,N_6200,N_6342);
nor U6591 (N_6591,N_6221,N_6209);
and U6592 (N_6592,N_6246,N_6392);
nand U6593 (N_6593,N_6276,N_6299);
nor U6594 (N_6594,N_6240,N_6363);
xnor U6595 (N_6595,N_6269,N_6277);
nor U6596 (N_6596,N_6244,N_6288);
xnor U6597 (N_6597,N_6282,N_6218);
xor U6598 (N_6598,N_6369,N_6399);
and U6599 (N_6599,N_6353,N_6373);
nand U6600 (N_6600,N_6585,N_6405);
nand U6601 (N_6601,N_6534,N_6520);
and U6602 (N_6602,N_6506,N_6452);
or U6603 (N_6603,N_6578,N_6433);
or U6604 (N_6604,N_6503,N_6402);
or U6605 (N_6605,N_6422,N_6404);
nand U6606 (N_6606,N_6507,N_6525);
xor U6607 (N_6607,N_6544,N_6476);
or U6608 (N_6608,N_6494,N_6439);
and U6609 (N_6609,N_6593,N_6523);
xor U6610 (N_6610,N_6545,N_6467);
nand U6611 (N_6611,N_6474,N_6565);
nand U6612 (N_6612,N_6418,N_6429);
or U6613 (N_6613,N_6481,N_6460);
nand U6614 (N_6614,N_6519,N_6497);
or U6615 (N_6615,N_6504,N_6448);
nand U6616 (N_6616,N_6482,N_6438);
nor U6617 (N_6617,N_6532,N_6556);
nand U6618 (N_6618,N_6581,N_6595);
and U6619 (N_6619,N_6562,N_6498);
and U6620 (N_6620,N_6459,N_6462);
and U6621 (N_6621,N_6457,N_6566);
nor U6622 (N_6622,N_6555,N_6415);
nand U6623 (N_6623,N_6445,N_6543);
or U6624 (N_6624,N_6434,N_6490);
xnor U6625 (N_6625,N_6473,N_6586);
or U6626 (N_6626,N_6496,N_6466);
or U6627 (N_6627,N_6589,N_6569);
nor U6628 (N_6628,N_6561,N_6584);
or U6629 (N_6629,N_6553,N_6444);
and U6630 (N_6630,N_6518,N_6488);
or U6631 (N_6631,N_6538,N_6411);
nand U6632 (N_6632,N_6501,N_6407);
and U6633 (N_6633,N_6436,N_6582);
xnor U6634 (N_6634,N_6500,N_6597);
and U6635 (N_6635,N_6419,N_6430);
nand U6636 (N_6636,N_6548,N_6567);
or U6637 (N_6637,N_6594,N_6468);
xnor U6638 (N_6638,N_6531,N_6479);
xnor U6639 (N_6639,N_6447,N_6401);
nor U6640 (N_6640,N_6557,N_6486);
nor U6641 (N_6641,N_6435,N_6575);
and U6642 (N_6642,N_6514,N_6588);
and U6643 (N_6643,N_6477,N_6550);
nor U6644 (N_6644,N_6591,N_6546);
and U6645 (N_6645,N_6484,N_6472);
and U6646 (N_6646,N_6470,N_6527);
nand U6647 (N_6647,N_6492,N_6446);
and U6648 (N_6648,N_6571,N_6540);
nor U6649 (N_6649,N_6590,N_6464);
or U6650 (N_6650,N_6536,N_6513);
and U6651 (N_6651,N_6420,N_6437);
or U6652 (N_6652,N_6552,N_6412);
or U6653 (N_6653,N_6592,N_6549);
nand U6654 (N_6654,N_6539,N_6480);
nand U6655 (N_6655,N_6400,N_6576);
or U6656 (N_6656,N_6414,N_6441);
xor U6657 (N_6657,N_6432,N_6443);
and U6658 (N_6658,N_6572,N_6522);
nand U6659 (N_6659,N_6568,N_6587);
nor U6660 (N_6660,N_6421,N_6461);
and U6661 (N_6661,N_6426,N_6424);
or U6662 (N_6662,N_6508,N_6509);
nand U6663 (N_6663,N_6502,N_6563);
and U6664 (N_6664,N_6528,N_6583);
nor U6665 (N_6665,N_6469,N_6535);
and U6666 (N_6666,N_6450,N_6558);
xor U6667 (N_6667,N_6451,N_6579);
or U6668 (N_6668,N_6521,N_6403);
and U6669 (N_6669,N_6431,N_6599);
xnor U6670 (N_6670,N_6570,N_6408);
and U6671 (N_6671,N_6596,N_6453);
xnor U6672 (N_6672,N_6560,N_6577);
or U6673 (N_6673,N_6442,N_6489);
nand U6674 (N_6674,N_6416,N_6487);
xnor U6675 (N_6675,N_6471,N_6598);
and U6676 (N_6676,N_6530,N_6491);
xor U6677 (N_6677,N_6574,N_6463);
nor U6678 (N_6678,N_6505,N_6427);
or U6679 (N_6679,N_6515,N_6413);
and U6680 (N_6680,N_6478,N_6495);
nand U6681 (N_6681,N_6458,N_6533);
and U6682 (N_6682,N_6485,N_6512);
nand U6683 (N_6683,N_6524,N_6559);
nor U6684 (N_6684,N_6564,N_6529);
nor U6685 (N_6685,N_6526,N_6541);
nand U6686 (N_6686,N_6537,N_6428);
or U6687 (N_6687,N_6475,N_6417);
nand U6688 (N_6688,N_6554,N_6410);
or U6689 (N_6689,N_6440,N_6551);
and U6690 (N_6690,N_6510,N_6483);
xor U6691 (N_6691,N_6455,N_6454);
nor U6692 (N_6692,N_6406,N_6499);
xor U6693 (N_6693,N_6493,N_6580);
nor U6694 (N_6694,N_6423,N_6456);
xnor U6695 (N_6695,N_6425,N_6449);
or U6696 (N_6696,N_6511,N_6465);
nand U6697 (N_6697,N_6516,N_6409);
nor U6698 (N_6698,N_6547,N_6517);
or U6699 (N_6699,N_6573,N_6542);
nand U6700 (N_6700,N_6542,N_6416);
and U6701 (N_6701,N_6430,N_6520);
xor U6702 (N_6702,N_6465,N_6567);
nand U6703 (N_6703,N_6442,N_6453);
nand U6704 (N_6704,N_6404,N_6553);
and U6705 (N_6705,N_6555,N_6551);
xor U6706 (N_6706,N_6451,N_6597);
or U6707 (N_6707,N_6532,N_6409);
xor U6708 (N_6708,N_6471,N_6412);
nand U6709 (N_6709,N_6515,N_6554);
or U6710 (N_6710,N_6582,N_6578);
xnor U6711 (N_6711,N_6466,N_6511);
nor U6712 (N_6712,N_6580,N_6576);
nand U6713 (N_6713,N_6559,N_6563);
xnor U6714 (N_6714,N_6432,N_6567);
or U6715 (N_6715,N_6461,N_6565);
xnor U6716 (N_6716,N_6502,N_6478);
nand U6717 (N_6717,N_6551,N_6446);
nor U6718 (N_6718,N_6489,N_6540);
nand U6719 (N_6719,N_6530,N_6430);
or U6720 (N_6720,N_6461,N_6438);
nand U6721 (N_6721,N_6501,N_6548);
nand U6722 (N_6722,N_6472,N_6536);
or U6723 (N_6723,N_6530,N_6487);
xnor U6724 (N_6724,N_6455,N_6548);
and U6725 (N_6725,N_6590,N_6402);
nand U6726 (N_6726,N_6461,N_6511);
or U6727 (N_6727,N_6427,N_6524);
nor U6728 (N_6728,N_6596,N_6545);
nand U6729 (N_6729,N_6554,N_6529);
or U6730 (N_6730,N_6548,N_6487);
nand U6731 (N_6731,N_6484,N_6421);
and U6732 (N_6732,N_6420,N_6529);
nor U6733 (N_6733,N_6531,N_6527);
or U6734 (N_6734,N_6530,N_6532);
or U6735 (N_6735,N_6492,N_6451);
nor U6736 (N_6736,N_6544,N_6502);
xnor U6737 (N_6737,N_6417,N_6412);
and U6738 (N_6738,N_6534,N_6453);
and U6739 (N_6739,N_6452,N_6487);
nor U6740 (N_6740,N_6554,N_6540);
xor U6741 (N_6741,N_6470,N_6476);
and U6742 (N_6742,N_6487,N_6414);
nor U6743 (N_6743,N_6581,N_6405);
xor U6744 (N_6744,N_6503,N_6457);
and U6745 (N_6745,N_6562,N_6412);
nor U6746 (N_6746,N_6432,N_6484);
nor U6747 (N_6747,N_6513,N_6520);
or U6748 (N_6748,N_6571,N_6513);
nor U6749 (N_6749,N_6412,N_6528);
nand U6750 (N_6750,N_6572,N_6484);
nor U6751 (N_6751,N_6592,N_6510);
nor U6752 (N_6752,N_6533,N_6462);
and U6753 (N_6753,N_6579,N_6588);
nand U6754 (N_6754,N_6497,N_6407);
and U6755 (N_6755,N_6536,N_6533);
and U6756 (N_6756,N_6420,N_6564);
nor U6757 (N_6757,N_6437,N_6537);
or U6758 (N_6758,N_6429,N_6493);
nor U6759 (N_6759,N_6586,N_6513);
or U6760 (N_6760,N_6597,N_6470);
nand U6761 (N_6761,N_6447,N_6468);
nor U6762 (N_6762,N_6403,N_6453);
xor U6763 (N_6763,N_6483,N_6491);
nand U6764 (N_6764,N_6454,N_6583);
nand U6765 (N_6765,N_6447,N_6591);
or U6766 (N_6766,N_6565,N_6505);
nand U6767 (N_6767,N_6440,N_6502);
and U6768 (N_6768,N_6549,N_6575);
nand U6769 (N_6769,N_6566,N_6595);
nand U6770 (N_6770,N_6505,N_6461);
or U6771 (N_6771,N_6561,N_6415);
or U6772 (N_6772,N_6403,N_6547);
nand U6773 (N_6773,N_6513,N_6421);
nor U6774 (N_6774,N_6471,N_6505);
or U6775 (N_6775,N_6461,N_6587);
xnor U6776 (N_6776,N_6562,N_6500);
xor U6777 (N_6777,N_6584,N_6437);
xor U6778 (N_6778,N_6489,N_6405);
nand U6779 (N_6779,N_6478,N_6479);
and U6780 (N_6780,N_6556,N_6401);
nand U6781 (N_6781,N_6439,N_6420);
and U6782 (N_6782,N_6470,N_6461);
or U6783 (N_6783,N_6534,N_6458);
nand U6784 (N_6784,N_6592,N_6413);
nor U6785 (N_6785,N_6540,N_6561);
nand U6786 (N_6786,N_6582,N_6555);
nand U6787 (N_6787,N_6423,N_6512);
xor U6788 (N_6788,N_6572,N_6428);
nor U6789 (N_6789,N_6473,N_6574);
or U6790 (N_6790,N_6404,N_6416);
and U6791 (N_6791,N_6585,N_6501);
nor U6792 (N_6792,N_6487,N_6540);
or U6793 (N_6793,N_6429,N_6402);
and U6794 (N_6794,N_6412,N_6485);
xnor U6795 (N_6795,N_6474,N_6469);
nor U6796 (N_6796,N_6474,N_6404);
nand U6797 (N_6797,N_6434,N_6529);
xor U6798 (N_6798,N_6481,N_6480);
or U6799 (N_6799,N_6459,N_6530);
nand U6800 (N_6800,N_6637,N_6745);
and U6801 (N_6801,N_6699,N_6754);
and U6802 (N_6802,N_6786,N_6622);
xnor U6803 (N_6803,N_6767,N_6661);
nor U6804 (N_6804,N_6755,N_6607);
and U6805 (N_6805,N_6645,N_6610);
xnor U6806 (N_6806,N_6707,N_6706);
or U6807 (N_6807,N_6605,N_6652);
and U6808 (N_6808,N_6611,N_6759);
nand U6809 (N_6809,N_6757,N_6743);
nand U6810 (N_6810,N_6783,N_6647);
nor U6811 (N_6811,N_6679,N_6692);
or U6812 (N_6812,N_6667,N_6775);
xnor U6813 (N_6813,N_6697,N_6792);
or U6814 (N_6814,N_6771,N_6604);
xor U6815 (N_6815,N_6772,N_6705);
nor U6816 (N_6816,N_6734,N_6644);
nand U6817 (N_6817,N_6632,N_6753);
nor U6818 (N_6818,N_6684,N_6781);
nand U6819 (N_6819,N_6694,N_6634);
nor U6820 (N_6820,N_6638,N_6768);
xnor U6821 (N_6821,N_6640,N_6613);
or U6822 (N_6822,N_6776,N_6618);
or U6823 (N_6823,N_6646,N_6691);
xnor U6824 (N_6824,N_6765,N_6678);
xor U6825 (N_6825,N_6628,N_6633);
and U6826 (N_6826,N_6724,N_6780);
xnor U6827 (N_6827,N_6749,N_6601);
or U6828 (N_6828,N_6614,N_6666);
nand U6829 (N_6829,N_6671,N_6630);
nand U6830 (N_6830,N_6631,N_6760);
nand U6831 (N_6831,N_6761,N_6681);
or U6832 (N_6832,N_6766,N_6793);
nand U6833 (N_6833,N_6711,N_6627);
nor U6834 (N_6834,N_6663,N_6798);
or U6835 (N_6835,N_6777,N_6785);
nor U6836 (N_6836,N_6725,N_6680);
nand U6837 (N_6837,N_6769,N_6696);
nand U6838 (N_6838,N_6704,N_6695);
xnor U6839 (N_6839,N_6670,N_6729);
or U6840 (N_6840,N_6625,N_6762);
and U6841 (N_6841,N_6741,N_6700);
xor U6842 (N_6842,N_6799,N_6612);
nor U6843 (N_6843,N_6600,N_6672);
and U6844 (N_6844,N_6702,N_6656);
nand U6845 (N_6845,N_6617,N_6752);
or U6846 (N_6846,N_6779,N_6626);
or U6847 (N_6847,N_6728,N_6606);
nand U6848 (N_6848,N_6687,N_6674);
xor U6849 (N_6849,N_6782,N_6732);
nor U6850 (N_6850,N_6701,N_6698);
or U6851 (N_6851,N_6688,N_6709);
and U6852 (N_6852,N_6721,N_6658);
xnor U6853 (N_6853,N_6778,N_6677);
xnor U6854 (N_6854,N_6756,N_6736);
and U6855 (N_6855,N_6673,N_6620);
nor U6856 (N_6856,N_6748,N_6693);
xnor U6857 (N_6857,N_6720,N_6722);
nor U6858 (N_6858,N_6682,N_6794);
xor U6859 (N_6859,N_6648,N_6730);
and U6860 (N_6860,N_6787,N_6657);
nor U6861 (N_6861,N_6738,N_6665);
nor U6862 (N_6862,N_6791,N_6784);
nor U6863 (N_6863,N_6710,N_6712);
or U6864 (N_6864,N_6764,N_6795);
xnor U6865 (N_6865,N_6735,N_6788);
and U6866 (N_6866,N_6763,N_6750);
nor U6867 (N_6867,N_6723,N_6608);
nand U6868 (N_6868,N_6603,N_6742);
nand U6869 (N_6869,N_6650,N_6770);
xnor U6870 (N_6870,N_6651,N_6718);
and U6871 (N_6871,N_6727,N_6602);
nor U6872 (N_6872,N_6797,N_6683);
and U6873 (N_6873,N_6773,N_6636);
or U6874 (N_6874,N_6653,N_6642);
and U6875 (N_6875,N_6668,N_6616);
and U6876 (N_6876,N_6719,N_6703);
xor U6877 (N_6877,N_6639,N_6740);
and U6878 (N_6878,N_6686,N_6747);
nor U6879 (N_6879,N_6731,N_6737);
nor U6880 (N_6880,N_6629,N_6758);
nand U6881 (N_6881,N_6654,N_6649);
xor U6882 (N_6882,N_6609,N_6746);
or U6883 (N_6883,N_6774,N_6664);
nor U6884 (N_6884,N_6690,N_6635);
nor U6885 (N_6885,N_6669,N_6708);
nand U6886 (N_6886,N_6789,N_6621);
nand U6887 (N_6887,N_6623,N_6641);
or U6888 (N_6888,N_6659,N_6662);
nand U6889 (N_6889,N_6717,N_6655);
or U6890 (N_6890,N_6660,N_6751);
nand U6891 (N_6891,N_6739,N_6714);
xor U6892 (N_6892,N_6643,N_6790);
xnor U6893 (N_6893,N_6615,N_6675);
xor U6894 (N_6894,N_6676,N_6689);
nand U6895 (N_6895,N_6726,N_6713);
nor U6896 (N_6896,N_6716,N_6744);
xor U6897 (N_6897,N_6685,N_6715);
or U6898 (N_6898,N_6733,N_6619);
nand U6899 (N_6899,N_6796,N_6624);
or U6900 (N_6900,N_6724,N_6660);
or U6901 (N_6901,N_6738,N_6637);
nor U6902 (N_6902,N_6752,N_6667);
nor U6903 (N_6903,N_6703,N_6677);
xor U6904 (N_6904,N_6741,N_6679);
nor U6905 (N_6905,N_6765,N_6747);
or U6906 (N_6906,N_6673,N_6775);
nand U6907 (N_6907,N_6703,N_6702);
or U6908 (N_6908,N_6664,N_6710);
and U6909 (N_6909,N_6791,N_6793);
nand U6910 (N_6910,N_6674,N_6711);
xnor U6911 (N_6911,N_6659,N_6763);
and U6912 (N_6912,N_6638,N_6795);
nand U6913 (N_6913,N_6696,N_6759);
or U6914 (N_6914,N_6751,N_6766);
and U6915 (N_6915,N_6740,N_6672);
nor U6916 (N_6916,N_6718,N_6690);
or U6917 (N_6917,N_6723,N_6795);
or U6918 (N_6918,N_6742,N_6623);
nor U6919 (N_6919,N_6658,N_6769);
nand U6920 (N_6920,N_6674,N_6699);
nand U6921 (N_6921,N_6609,N_6635);
nand U6922 (N_6922,N_6771,N_6629);
nand U6923 (N_6923,N_6746,N_6781);
or U6924 (N_6924,N_6743,N_6677);
nand U6925 (N_6925,N_6798,N_6633);
or U6926 (N_6926,N_6709,N_6760);
or U6927 (N_6927,N_6749,N_6640);
xor U6928 (N_6928,N_6777,N_6602);
nor U6929 (N_6929,N_6616,N_6617);
nor U6930 (N_6930,N_6629,N_6793);
and U6931 (N_6931,N_6769,N_6618);
xor U6932 (N_6932,N_6735,N_6615);
xnor U6933 (N_6933,N_6735,N_6616);
and U6934 (N_6934,N_6684,N_6713);
nand U6935 (N_6935,N_6792,N_6666);
or U6936 (N_6936,N_6652,N_6724);
nand U6937 (N_6937,N_6785,N_6600);
or U6938 (N_6938,N_6751,N_6724);
nor U6939 (N_6939,N_6613,N_6757);
nand U6940 (N_6940,N_6725,N_6678);
and U6941 (N_6941,N_6609,N_6692);
nand U6942 (N_6942,N_6722,N_6798);
and U6943 (N_6943,N_6776,N_6652);
and U6944 (N_6944,N_6658,N_6719);
or U6945 (N_6945,N_6635,N_6723);
xor U6946 (N_6946,N_6625,N_6737);
nor U6947 (N_6947,N_6705,N_6794);
and U6948 (N_6948,N_6621,N_6773);
and U6949 (N_6949,N_6633,N_6618);
or U6950 (N_6950,N_6657,N_6625);
and U6951 (N_6951,N_6621,N_6610);
or U6952 (N_6952,N_6736,N_6699);
xor U6953 (N_6953,N_6636,N_6761);
nor U6954 (N_6954,N_6789,N_6690);
xor U6955 (N_6955,N_6745,N_6700);
nand U6956 (N_6956,N_6725,N_6698);
and U6957 (N_6957,N_6666,N_6673);
xor U6958 (N_6958,N_6655,N_6770);
or U6959 (N_6959,N_6629,N_6792);
nand U6960 (N_6960,N_6716,N_6795);
xor U6961 (N_6961,N_6733,N_6749);
nor U6962 (N_6962,N_6770,N_6696);
nor U6963 (N_6963,N_6612,N_6697);
xnor U6964 (N_6964,N_6732,N_6711);
xnor U6965 (N_6965,N_6715,N_6604);
or U6966 (N_6966,N_6742,N_6629);
and U6967 (N_6967,N_6632,N_6723);
or U6968 (N_6968,N_6646,N_6775);
nand U6969 (N_6969,N_6603,N_6607);
xor U6970 (N_6970,N_6731,N_6732);
or U6971 (N_6971,N_6723,N_6758);
or U6972 (N_6972,N_6627,N_6609);
and U6973 (N_6973,N_6699,N_6654);
nand U6974 (N_6974,N_6649,N_6699);
or U6975 (N_6975,N_6764,N_6653);
nand U6976 (N_6976,N_6690,N_6759);
or U6977 (N_6977,N_6712,N_6718);
nor U6978 (N_6978,N_6761,N_6758);
and U6979 (N_6979,N_6730,N_6773);
xnor U6980 (N_6980,N_6641,N_6788);
and U6981 (N_6981,N_6730,N_6619);
nand U6982 (N_6982,N_6706,N_6746);
and U6983 (N_6983,N_6627,N_6742);
or U6984 (N_6984,N_6743,N_6763);
nand U6985 (N_6985,N_6760,N_6661);
and U6986 (N_6986,N_6672,N_6762);
or U6987 (N_6987,N_6706,N_6623);
or U6988 (N_6988,N_6603,N_6609);
nand U6989 (N_6989,N_6728,N_6693);
and U6990 (N_6990,N_6739,N_6675);
or U6991 (N_6991,N_6653,N_6691);
xnor U6992 (N_6992,N_6678,N_6755);
or U6993 (N_6993,N_6719,N_6710);
nand U6994 (N_6994,N_6783,N_6765);
and U6995 (N_6995,N_6733,N_6784);
xnor U6996 (N_6996,N_6718,N_6641);
or U6997 (N_6997,N_6754,N_6788);
and U6998 (N_6998,N_6685,N_6628);
nand U6999 (N_6999,N_6686,N_6795);
or U7000 (N_7000,N_6850,N_6828);
nor U7001 (N_7001,N_6812,N_6922);
xnor U7002 (N_7002,N_6880,N_6911);
or U7003 (N_7003,N_6969,N_6981);
xor U7004 (N_7004,N_6886,N_6957);
nor U7005 (N_7005,N_6825,N_6913);
xnor U7006 (N_7006,N_6811,N_6876);
nor U7007 (N_7007,N_6838,N_6910);
xor U7008 (N_7008,N_6961,N_6968);
nor U7009 (N_7009,N_6834,N_6996);
and U7010 (N_7010,N_6835,N_6832);
nor U7011 (N_7011,N_6921,N_6955);
or U7012 (N_7012,N_6837,N_6898);
nor U7013 (N_7013,N_6973,N_6925);
nand U7014 (N_7014,N_6950,N_6853);
or U7015 (N_7015,N_6836,N_6967);
nor U7016 (N_7016,N_6875,N_6942);
and U7017 (N_7017,N_6872,N_6936);
and U7018 (N_7018,N_6993,N_6866);
nor U7019 (N_7019,N_6982,N_6839);
nor U7020 (N_7020,N_6804,N_6907);
nor U7021 (N_7021,N_6935,N_6851);
and U7022 (N_7022,N_6818,N_6855);
and U7023 (N_7023,N_6823,N_6831);
nor U7024 (N_7024,N_6975,N_6966);
nor U7025 (N_7025,N_6939,N_6879);
nand U7026 (N_7026,N_6802,N_6934);
nand U7027 (N_7027,N_6927,N_6801);
and U7028 (N_7028,N_6900,N_6958);
and U7029 (N_7029,N_6928,N_6926);
nor U7030 (N_7030,N_6809,N_6891);
nor U7031 (N_7031,N_6972,N_6862);
nand U7032 (N_7032,N_6941,N_6960);
nor U7033 (N_7033,N_6882,N_6817);
or U7034 (N_7034,N_6870,N_6971);
xor U7035 (N_7035,N_6937,N_6991);
nand U7036 (N_7036,N_6978,N_6874);
and U7037 (N_7037,N_6884,N_6877);
and U7038 (N_7038,N_6888,N_6814);
and U7039 (N_7039,N_6918,N_6956);
nor U7040 (N_7040,N_6945,N_6822);
or U7041 (N_7041,N_6871,N_6923);
xnor U7042 (N_7042,N_6819,N_6917);
nand U7043 (N_7043,N_6827,N_6830);
or U7044 (N_7044,N_6906,N_6965);
and U7045 (N_7045,N_6909,N_6845);
xnor U7046 (N_7046,N_6805,N_6897);
or U7047 (N_7047,N_6854,N_6990);
or U7048 (N_7048,N_6873,N_6901);
and U7049 (N_7049,N_6985,N_6896);
and U7050 (N_7050,N_6868,N_6826);
xnor U7051 (N_7051,N_6930,N_6994);
nand U7052 (N_7052,N_6915,N_6849);
nor U7053 (N_7053,N_6895,N_6887);
nor U7054 (N_7054,N_6952,N_6892);
nand U7055 (N_7055,N_6998,N_6905);
or U7056 (N_7056,N_6829,N_6964);
or U7057 (N_7057,N_6869,N_6806);
nand U7058 (N_7058,N_6940,N_6903);
xnor U7059 (N_7059,N_6933,N_6867);
nor U7060 (N_7060,N_6943,N_6963);
xnor U7061 (N_7061,N_6983,N_6919);
nand U7062 (N_7062,N_6904,N_6995);
nand U7063 (N_7063,N_6916,N_6987);
and U7064 (N_7064,N_6989,N_6999);
and U7065 (N_7065,N_6899,N_6890);
nor U7066 (N_7066,N_6848,N_6979);
nand U7067 (N_7067,N_6949,N_6931);
nand U7068 (N_7068,N_6807,N_6912);
xor U7069 (N_7069,N_6800,N_6840);
or U7070 (N_7070,N_6929,N_6988);
nor U7071 (N_7071,N_6951,N_6980);
xor U7072 (N_7072,N_6997,N_6986);
nor U7073 (N_7073,N_6842,N_6932);
and U7074 (N_7074,N_6908,N_6865);
and U7075 (N_7075,N_6803,N_6847);
nand U7076 (N_7076,N_6813,N_6858);
and U7077 (N_7077,N_6824,N_6893);
nand U7078 (N_7078,N_6902,N_6959);
nand U7079 (N_7079,N_6859,N_6841);
and U7080 (N_7080,N_6810,N_6970);
xor U7081 (N_7081,N_6962,N_6863);
or U7082 (N_7082,N_6860,N_6976);
nor U7083 (N_7083,N_6914,N_6881);
or U7084 (N_7084,N_6864,N_6857);
and U7085 (N_7085,N_6852,N_6953);
and U7086 (N_7086,N_6889,N_6816);
xnor U7087 (N_7087,N_6885,N_6883);
nand U7088 (N_7088,N_6948,N_6833);
and U7089 (N_7089,N_6846,N_6808);
and U7090 (N_7090,N_6878,N_6974);
xor U7091 (N_7091,N_6843,N_6954);
and U7092 (N_7092,N_6894,N_6944);
nor U7093 (N_7093,N_6984,N_6861);
nor U7094 (N_7094,N_6992,N_6820);
nor U7095 (N_7095,N_6844,N_6815);
xnor U7096 (N_7096,N_6947,N_6977);
xnor U7097 (N_7097,N_6821,N_6924);
and U7098 (N_7098,N_6938,N_6920);
xor U7099 (N_7099,N_6856,N_6946);
or U7100 (N_7100,N_6897,N_6949);
and U7101 (N_7101,N_6834,N_6919);
xor U7102 (N_7102,N_6878,N_6880);
nor U7103 (N_7103,N_6898,N_6957);
nand U7104 (N_7104,N_6974,N_6958);
or U7105 (N_7105,N_6985,N_6920);
nand U7106 (N_7106,N_6837,N_6881);
or U7107 (N_7107,N_6957,N_6861);
nor U7108 (N_7108,N_6908,N_6834);
xor U7109 (N_7109,N_6930,N_6929);
and U7110 (N_7110,N_6840,N_6887);
and U7111 (N_7111,N_6814,N_6937);
xor U7112 (N_7112,N_6949,N_6814);
nor U7113 (N_7113,N_6906,N_6917);
and U7114 (N_7114,N_6907,N_6995);
or U7115 (N_7115,N_6835,N_6834);
nand U7116 (N_7116,N_6987,N_6982);
or U7117 (N_7117,N_6958,N_6908);
nor U7118 (N_7118,N_6819,N_6818);
xor U7119 (N_7119,N_6865,N_6880);
or U7120 (N_7120,N_6898,N_6871);
and U7121 (N_7121,N_6885,N_6977);
xor U7122 (N_7122,N_6908,N_6809);
and U7123 (N_7123,N_6905,N_6951);
or U7124 (N_7124,N_6958,N_6972);
or U7125 (N_7125,N_6955,N_6931);
nor U7126 (N_7126,N_6919,N_6877);
or U7127 (N_7127,N_6868,N_6839);
nor U7128 (N_7128,N_6806,N_6974);
xnor U7129 (N_7129,N_6817,N_6902);
nand U7130 (N_7130,N_6851,N_6958);
xnor U7131 (N_7131,N_6846,N_6822);
nor U7132 (N_7132,N_6881,N_6953);
or U7133 (N_7133,N_6809,N_6800);
nand U7134 (N_7134,N_6813,N_6897);
and U7135 (N_7135,N_6888,N_6896);
or U7136 (N_7136,N_6919,N_6959);
and U7137 (N_7137,N_6805,N_6935);
nand U7138 (N_7138,N_6961,N_6912);
nand U7139 (N_7139,N_6973,N_6883);
and U7140 (N_7140,N_6998,N_6848);
or U7141 (N_7141,N_6906,N_6884);
or U7142 (N_7142,N_6985,N_6902);
xor U7143 (N_7143,N_6994,N_6884);
xor U7144 (N_7144,N_6863,N_6954);
and U7145 (N_7145,N_6981,N_6918);
xnor U7146 (N_7146,N_6861,N_6891);
and U7147 (N_7147,N_6989,N_6993);
nor U7148 (N_7148,N_6861,N_6898);
nand U7149 (N_7149,N_6998,N_6908);
nor U7150 (N_7150,N_6946,N_6801);
nor U7151 (N_7151,N_6822,N_6930);
and U7152 (N_7152,N_6889,N_6901);
xor U7153 (N_7153,N_6899,N_6859);
or U7154 (N_7154,N_6846,N_6976);
or U7155 (N_7155,N_6976,N_6867);
nand U7156 (N_7156,N_6968,N_6970);
or U7157 (N_7157,N_6862,N_6974);
nor U7158 (N_7158,N_6948,N_6861);
xnor U7159 (N_7159,N_6965,N_6973);
nand U7160 (N_7160,N_6815,N_6965);
nand U7161 (N_7161,N_6965,N_6998);
nor U7162 (N_7162,N_6997,N_6925);
or U7163 (N_7163,N_6852,N_6912);
or U7164 (N_7164,N_6903,N_6824);
or U7165 (N_7165,N_6973,N_6861);
xor U7166 (N_7166,N_6950,N_6829);
nor U7167 (N_7167,N_6907,N_6993);
and U7168 (N_7168,N_6880,N_6841);
xor U7169 (N_7169,N_6860,N_6913);
or U7170 (N_7170,N_6936,N_6920);
or U7171 (N_7171,N_6902,N_6972);
or U7172 (N_7172,N_6802,N_6943);
and U7173 (N_7173,N_6944,N_6859);
nand U7174 (N_7174,N_6901,N_6932);
and U7175 (N_7175,N_6904,N_6837);
or U7176 (N_7176,N_6923,N_6849);
or U7177 (N_7177,N_6963,N_6983);
nor U7178 (N_7178,N_6822,N_6839);
and U7179 (N_7179,N_6916,N_6985);
and U7180 (N_7180,N_6813,N_6823);
and U7181 (N_7181,N_6828,N_6995);
xor U7182 (N_7182,N_6800,N_6944);
or U7183 (N_7183,N_6818,N_6856);
xor U7184 (N_7184,N_6959,N_6925);
xor U7185 (N_7185,N_6958,N_6876);
or U7186 (N_7186,N_6993,N_6807);
nand U7187 (N_7187,N_6922,N_6806);
nand U7188 (N_7188,N_6876,N_6836);
nor U7189 (N_7189,N_6925,N_6804);
nor U7190 (N_7190,N_6968,N_6847);
xnor U7191 (N_7191,N_6871,N_6910);
nand U7192 (N_7192,N_6964,N_6939);
nor U7193 (N_7193,N_6833,N_6953);
nand U7194 (N_7194,N_6944,N_6856);
nand U7195 (N_7195,N_6824,N_6846);
nand U7196 (N_7196,N_6992,N_6874);
or U7197 (N_7197,N_6978,N_6943);
nand U7198 (N_7198,N_6898,N_6911);
nor U7199 (N_7199,N_6855,N_6895);
or U7200 (N_7200,N_7055,N_7049);
nor U7201 (N_7201,N_7066,N_7071);
or U7202 (N_7202,N_7112,N_7152);
nand U7203 (N_7203,N_7180,N_7107);
or U7204 (N_7204,N_7185,N_7114);
nor U7205 (N_7205,N_7094,N_7189);
or U7206 (N_7206,N_7103,N_7104);
xnor U7207 (N_7207,N_7096,N_7053);
xnor U7208 (N_7208,N_7051,N_7172);
nor U7209 (N_7209,N_7080,N_7087);
nor U7210 (N_7210,N_7121,N_7048);
xor U7211 (N_7211,N_7007,N_7128);
and U7212 (N_7212,N_7068,N_7110);
xnor U7213 (N_7213,N_7034,N_7070);
nand U7214 (N_7214,N_7092,N_7173);
or U7215 (N_7215,N_7024,N_7109);
or U7216 (N_7216,N_7134,N_7009);
nand U7217 (N_7217,N_7117,N_7129);
xor U7218 (N_7218,N_7085,N_7165);
or U7219 (N_7219,N_7041,N_7072);
xor U7220 (N_7220,N_7136,N_7157);
and U7221 (N_7221,N_7101,N_7016);
nand U7222 (N_7222,N_7124,N_7175);
or U7223 (N_7223,N_7042,N_7018);
nor U7224 (N_7224,N_7057,N_7137);
xnor U7225 (N_7225,N_7133,N_7073);
nor U7226 (N_7226,N_7091,N_7111);
or U7227 (N_7227,N_7154,N_7193);
and U7228 (N_7228,N_7196,N_7043);
nand U7229 (N_7229,N_7075,N_7145);
and U7230 (N_7230,N_7195,N_7008);
xnor U7231 (N_7231,N_7064,N_7184);
and U7232 (N_7232,N_7026,N_7058);
nor U7233 (N_7233,N_7187,N_7151);
nand U7234 (N_7234,N_7159,N_7001);
xor U7235 (N_7235,N_7106,N_7002);
nand U7236 (N_7236,N_7127,N_7030);
nor U7237 (N_7237,N_7181,N_7105);
nor U7238 (N_7238,N_7141,N_7168);
or U7239 (N_7239,N_7156,N_7097);
nor U7240 (N_7240,N_7183,N_7131);
and U7241 (N_7241,N_7093,N_7033);
and U7242 (N_7242,N_7010,N_7149);
xnor U7243 (N_7243,N_7054,N_7169);
nor U7244 (N_7244,N_7084,N_7166);
or U7245 (N_7245,N_7147,N_7120);
and U7246 (N_7246,N_7179,N_7148);
nor U7247 (N_7247,N_7046,N_7031);
and U7248 (N_7248,N_7047,N_7176);
or U7249 (N_7249,N_7090,N_7142);
xnor U7250 (N_7250,N_7078,N_7050);
nand U7251 (N_7251,N_7089,N_7059);
or U7252 (N_7252,N_7029,N_7186);
nand U7253 (N_7253,N_7170,N_7188);
nand U7254 (N_7254,N_7130,N_7045);
nand U7255 (N_7255,N_7155,N_7062);
nand U7256 (N_7256,N_7038,N_7119);
nand U7257 (N_7257,N_7012,N_7199);
or U7258 (N_7258,N_7003,N_7140);
or U7259 (N_7259,N_7076,N_7113);
nor U7260 (N_7260,N_7023,N_7138);
and U7261 (N_7261,N_7011,N_7100);
nand U7262 (N_7262,N_7162,N_7126);
nand U7263 (N_7263,N_7164,N_7074);
and U7264 (N_7264,N_7146,N_7099);
nand U7265 (N_7265,N_7019,N_7088);
or U7266 (N_7266,N_7178,N_7021);
nand U7267 (N_7267,N_7095,N_7198);
nand U7268 (N_7268,N_7061,N_7060);
nand U7269 (N_7269,N_7108,N_7160);
xor U7270 (N_7270,N_7102,N_7115);
and U7271 (N_7271,N_7067,N_7077);
and U7272 (N_7272,N_7167,N_7005);
xor U7273 (N_7273,N_7150,N_7079);
xor U7274 (N_7274,N_7144,N_7020);
and U7275 (N_7275,N_7035,N_7083);
xor U7276 (N_7276,N_7177,N_7065);
nor U7277 (N_7277,N_7039,N_7081);
or U7278 (N_7278,N_7158,N_7118);
and U7279 (N_7279,N_7153,N_7000);
nor U7280 (N_7280,N_7191,N_7069);
nor U7281 (N_7281,N_7052,N_7132);
nor U7282 (N_7282,N_7116,N_7163);
or U7283 (N_7283,N_7125,N_7135);
nand U7284 (N_7284,N_7197,N_7098);
xnor U7285 (N_7285,N_7028,N_7082);
and U7286 (N_7286,N_7192,N_7022);
and U7287 (N_7287,N_7006,N_7013);
and U7288 (N_7288,N_7139,N_7086);
xnor U7289 (N_7289,N_7171,N_7015);
and U7290 (N_7290,N_7025,N_7040);
nand U7291 (N_7291,N_7063,N_7174);
or U7292 (N_7292,N_7014,N_7032);
nand U7293 (N_7293,N_7044,N_7161);
xnor U7294 (N_7294,N_7122,N_7004);
nand U7295 (N_7295,N_7123,N_7194);
nand U7296 (N_7296,N_7027,N_7190);
xor U7297 (N_7297,N_7036,N_7143);
nand U7298 (N_7298,N_7182,N_7017);
or U7299 (N_7299,N_7037,N_7056);
or U7300 (N_7300,N_7149,N_7057);
or U7301 (N_7301,N_7021,N_7183);
xor U7302 (N_7302,N_7114,N_7099);
and U7303 (N_7303,N_7084,N_7031);
and U7304 (N_7304,N_7058,N_7169);
nor U7305 (N_7305,N_7046,N_7154);
nand U7306 (N_7306,N_7070,N_7140);
and U7307 (N_7307,N_7022,N_7105);
or U7308 (N_7308,N_7092,N_7116);
or U7309 (N_7309,N_7067,N_7022);
or U7310 (N_7310,N_7197,N_7117);
nand U7311 (N_7311,N_7046,N_7185);
and U7312 (N_7312,N_7144,N_7036);
nor U7313 (N_7313,N_7196,N_7036);
and U7314 (N_7314,N_7072,N_7143);
or U7315 (N_7315,N_7148,N_7177);
or U7316 (N_7316,N_7154,N_7162);
or U7317 (N_7317,N_7064,N_7120);
or U7318 (N_7318,N_7123,N_7175);
nand U7319 (N_7319,N_7161,N_7065);
nor U7320 (N_7320,N_7072,N_7076);
or U7321 (N_7321,N_7132,N_7126);
or U7322 (N_7322,N_7168,N_7187);
nand U7323 (N_7323,N_7090,N_7176);
or U7324 (N_7324,N_7054,N_7082);
nand U7325 (N_7325,N_7152,N_7199);
nor U7326 (N_7326,N_7028,N_7097);
and U7327 (N_7327,N_7075,N_7061);
nor U7328 (N_7328,N_7067,N_7034);
or U7329 (N_7329,N_7098,N_7187);
nand U7330 (N_7330,N_7050,N_7088);
xor U7331 (N_7331,N_7155,N_7031);
or U7332 (N_7332,N_7050,N_7037);
xnor U7333 (N_7333,N_7033,N_7010);
or U7334 (N_7334,N_7045,N_7108);
nand U7335 (N_7335,N_7008,N_7018);
nor U7336 (N_7336,N_7060,N_7050);
or U7337 (N_7337,N_7012,N_7021);
or U7338 (N_7338,N_7193,N_7094);
xor U7339 (N_7339,N_7044,N_7073);
nor U7340 (N_7340,N_7166,N_7006);
xor U7341 (N_7341,N_7012,N_7029);
xor U7342 (N_7342,N_7046,N_7047);
and U7343 (N_7343,N_7194,N_7063);
xor U7344 (N_7344,N_7119,N_7089);
nor U7345 (N_7345,N_7142,N_7000);
nor U7346 (N_7346,N_7085,N_7162);
and U7347 (N_7347,N_7137,N_7035);
nand U7348 (N_7348,N_7023,N_7025);
or U7349 (N_7349,N_7056,N_7035);
xor U7350 (N_7350,N_7122,N_7055);
and U7351 (N_7351,N_7133,N_7130);
nand U7352 (N_7352,N_7072,N_7199);
nand U7353 (N_7353,N_7084,N_7098);
and U7354 (N_7354,N_7005,N_7004);
nand U7355 (N_7355,N_7020,N_7008);
nand U7356 (N_7356,N_7065,N_7195);
nand U7357 (N_7357,N_7060,N_7118);
nand U7358 (N_7358,N_7185,N_7126);
nor U7359 (N_7359,N_7099,N_7177);
and U7360 (N_7360,N_7187,N_7107);
xor U7361 (N_7361,N_7003,N_7107);
nand U7362 (N_7362,N_7011,N_7176);
or U7363 (N_7363,N_7012,N_7180);
and U7364 (N_7364,N_7120,N_7171);
nor U7365 (N_7365,N_7045,N_7067);
xor U7366 (N_7366,N_7097,N_7058);
nor U7367 (N_7367,N_7165,N_7019);
and U7368 (N_7368,N_7110,N_7125);
nor U7369 (N_7369,N_7149,N_7015);
nor U7370 (N_7370,N_7020,N_7192);
or U7371 (N_7371,N_7070,N_7194);
or U7372 (N_7372,N_7045,N_7159);
nand U7373 (N_7373,N_7156,N_7013);
or U7374 (N_7374,N_7030,N_7052);
and U7375 (N_7375,N_7160,N_7068);
xor U7376 (N_7376,N_7136,N_7021);
and U7377 (N_7377,N_7159,N_7100);
and U7378 (N_7378,N_7124,N_7168);
nand U7379 (N_7379,N_7143,N_7110);
nand U7380 (N_7380,N_7040,N_7145);
nor U7381 (N_7381,N_7154,N_7073);
xnor U7382 (N_7382,N_7047,N_7179);
and U7383 (N_7383,N_7024,N_7017);
xor U7384 (N_7384,N_7058,N_7027);
nor U7385 (N_7385,N_7132,N_7196);
and U7386 (N_7386,N_7072,N_7164);
nand U7387 (N_7387,N_7178,N_7189);
nand U7388 (N_7388,N_7064,N_7111);
nor U7389 (N_7389,N_7172,N_7184);
or U7390 (N_7390,N_7006,N_7099);
or U7391 (N_7391,N_7167,N_7126);
nor U7392 (N_7392,N_7192,N_7071);
nand U7393 (N_7393,N_7106,N_7020);
nand U7394 (N_7394,N_7142,N_7158);
nor U7395 (N_7395,N_7102,N_7186);
xnor U7396 (N_7396,N_7118,N_7062);
nor U7397 (N_7397,N_7155,N_7141);
and U7398 (N_7398,N_7104,N_7049);
or U7399 (N_7399,N_7022,N_7056);
nor U7400 (N_7400,N_7313,N_7205);
xor U7401 (N_7401,N_7229,N_7364);
and U7402 (N_7402,N_7376,N_7253);
xor U7403 (N_7403,N_7237,N_7339);
nand U7404 (N_7404,N_7280,N_7201);
or U7405 (N_7405,N_7221,N_7219);
or U7406 (N_7406,N_7378,N_7325);
nand U7407 (N_7407,N_7356,N_7332);
and U7408 (N_7408,N_7210,N_7289);
and U7409 (N_7409,N_7244,N_7296);
and U7410 (N_7410,N_7304,N_7264);
or U7411 (N_7411,N_7366,N_7348);
xnor U7412 (N_7412,N_7246,N_7389);
and U7413 (N_7413,N_7248,N_7225);
and U7414 (N_7414,N_7334,N_7355);
or U7415 (N_7415,N_7218,N_7267);
and U7416 (N_7416,N_7252,N_7240);
and U7417 (N_7417,N_7336,N_7395);
xnor U7418 (N_7418,N_7272,N_7343);
nand U7419 (N_7419,N_7266,N_7394);
and U7420 (N_7420,N_7274,N_7352);
and U7421 (N_7421,N_7242,N_7231);
xnor U7422 (N_7422,N_7263,N_7373);
or U7423 (N_7423,N_7206,N_7305);
or U7424 (N_7424,N_7350,N_7234);
and U7425 (N_7425,N_7388,N_7261);
or U7426 (N_7426,N_7207,N_7391);
and U7427 (N_7427,N_7213,N_7357);
and U7428 (N_7428,N_7281,N_7317);
nor U7429 (N_7429,N_7249,N_7200);
nand U7430 (N_7430,N_7291,N_7299);
or U7431 (N_7431,N_7380,N_7258);
or U7432 (N_7432,N_7302,N_7337);
nor U7433 (N_7433,N_7294,N_7370);
xor U7434 (N_7434,N_7278,N_7368);
and U7435 (N_7435,N_7220,N_7393);
or U7436 (N_7436,N_7275,N_7297);
nor U7437 (N_7437,N_7271,N_7345);
or U7438 (N_7438,N_7341,N_7212);
or U7439 (N_7439,N_7236,N_7360);
or U7440 (N_7440,N_7224,N_7367);
or U7441 (N_7441,N_7318,N_7331);
nor U7442 (N_7442,N_7319,N_7362);
xnor U7443 (N_7443,N_7397,N_7365);
nand U7444 (N_7444,N_7354,N_7239);
and U7445 (N_7445,N_7342,N_7273);
or U7446 (N_7446,N_7384,N_7335);
xor U7447 (N_7447,N_7311,N_7320);
and U7448 (N_7448,N_7288,N_7321);
nand U7449 (N_7449,N_7260,N_7340);
nand U7450 (N_7450,N_7309,N_7347);
nor U7451 (N_7451,N_7303,N_7270);
nor U7452 (N_7452,N_7315,N_7215);
or U7453 (N_7453,N_7371,N_7359);
or U7454 (N_7454,N_7312,N_7290);
or U7455 (N_7455,N_7282,N_7287);
and U7456 (N_7456,N_7308,N_7284);
and U7457 (N_7457,N_7310,N_7227);
nand U7458 (N_7458,N_7247,N_7230);
and U7459 (N_7459,N_7265,N_7292);
nand U7460 (N_7460,N_7392,N_7387);
nor U7461 (N_7461,N_7202,N_7324);
or U7462 (N_7462,N_7301,N_7208);
and U7463 (N_7463,N_7369,N_7251);
and U7464 (N_7464,N_7353,N_7222);
and U7465 (N_7465,N_7344,N_7255);
xnor U7466 (N_7466,N_7358,N_7214);
nor U7467 (N_7467,N_7257,N_7295);
and U7468 (N_7468,N_7346,N_7361);
nand U7469 (N_7469,N_7241,N_7306);
nand U7470 (N_7470,N_7398,N_7211);
and U7471 (N_7471,N_7277,N_7327);
xor U7472 (N_7472,N_7245,N_7233);
nand U7473 (N_7473,N_7283,N_7243);
xnor U7474 (N_7474,N_7250,N_7279);
nor U7475 (N_7475,N_7381,N_7385);
nand U7476 (N_7476,N_7363,N_7322);
nand U7477 (N_7477,N_7383,N_7226);
xor U7478 (N_7478,N_7382,N_7307);
nor U7479 (N_7479,N_7323,N_7262);
or U7480 (N_7480,N_7349,N_7209);
and U7481 (N_7481,N_7399,N_7390);
nand U7482 (N_7482,N_7386,N_7228);
nand U7483 (N_7483,N_7293,N_7269);
xnor U7484 (N_7484,N_7256,N_7276);
nand U7485 (N_7485,N_7217,N_7238);
nor U7486 (N_7486,N_7223,N_7351);
nand U7487 (N_7487,N_7286,N_7328);
xor U7488 (N_7488,N_7377,N_7316);
or U7489 (N_7489,N_7314,N_7232);
nor U7490 (N_7490,N_7338,N_7259);
or U7491 (N_7491,N_7298,N_7330);
and U7492 (N_7492,N_7300,N_7329);
nor U7493 (N_7493,N_7379,N_7203);
or U7494 (N_7494,N_7235,N_7372);
nand U7495 (N_7495,N_7375,N_7204);
nand U7496 (N_7496,N_7268,N_7396);
nand U7497 (N_7497,N_7333,N_7254);
or U7498 (N_7498,N_7374,N_7285);
or U7499 (N_7499,N_7326,N_7216);
nand U7500 (N_7500,N_7259,N_7382);
nand U7501 (N_7501,N_7399,N_7262);
or U7502 (N_7502,N_7300,N_7373);
xnor U7503 (N_7503,N_7212,N_7244);
and U7504 (N_7504,N_7306,N_7257);
nor U7505 (N_7505,N_7363,N_7229);
and U7506 (N_7506,N_7281,N_7387);
nand U7507 (N_7507,N_7314,N_7305);
nand U7508 (N_7508,N_7368,N_7386);
or U7509 (N_7509,N_7254,N_7373);
xor U7510 (N_7510,N_7363,N_7289);
xnor U7511 (N_7511,N_7325,N_7294);
and U7512 (N_7512,N_7220,N_7331);
or U7513 (N_7513,N_7352,N_7252);
and U7514 (N_7514,N_7282,N_7387);
and U7515 (N_7515,N_7384,N_7360);
nand U7516 (N_7516,N_7375,N_7338);
nor U7517 (N_7517,N_7222,N_7259);
and U7518 (N_7518,N_7275,N_7324);
xnor U7519 (N_7519,N_7293,N_7263);
and U7520 (N_7520,N_7370,N_7215);
nor U7521 (N_7521,N_7234,N_7236);
xor U7522 (N_7522,N_7329,N_7380);
and U7523 (N_7523,N_7387,N_7228);
or U7524 (N_7524,N_7380,N_7327);
or U7525 (N_7525,N_7291,N_7395);
nor U7526 (N_7526,N_7326,N_7328);
and U7527 (N_7527,N_7389,N_7338);
or U7528 (N_7528,N_7289,N_7351);
nand U7529 (N_7529,N_7263,N_7383);
or U7530 (N_7530,N_7297,N_7229);
or U7531 (N_7531,N_7366,N_7259);
or U7532 (N_7532,N_7260,N_7310);
and U7533 (N_7533,N_7208,N_7392);
or U7534 (N_7534,N_7261,N_7387);
and U7535 (N_7535,N_7237,N_7376);
or U7536 (N_7536,N_7368,N_7305);
nor U7537 (N_7537,N_7293,N_7262);
nand U7538 (N_7538,N_7317,N_7236);
xor U7539 (N_7539,N_7233,N_7230);
xnor U7540 (N_7540,N_7316,N_7227);
nand U7541 (N_7541,N_7314,N_7249);
and U7542 (N_7542,N_7287,N_7247);
or U7543 (N_7543,N_7376,N_7396);
nor U7544 (N_7544,N_7258,N_7359);
and U7545 (N_7545,N_7215,N_7364);
and U7546 (N_7546,N_7322,N_7213);
xor U7547 (N_7547,N_7393,N_7275);
nand U7548 (N_7548,N_7340,N_7368);
nor U7549 (N_7549,N_7240,N_7370);
nand U7550 (N_7550,N_7324,N_7306);
or U7551 (N_7551,N_7212,N_7387);
nand U7552 (N_7552,N_7204,N_7394);
and U7553 (N_7553,N_7393,N_7232);
nand U7554 (N_7554,N_7374,N_7210);
xor U7555 (N_7555,N_7215,N_7320);
nand U7556 (N_7556,N_7362,N_7329);
and U7557 (N_7557,N_7253,N_7382);
or U7558 (N_7558,N_7218,N_7311);
nor U7559 (N_7559,N_7308,N_7298);
nor U7560 (N_7560,N_7297,N_7288);
or U7561 (N_7561,N_7315,N_7311);
nor U7562 (N_7562,N_7288,N_7245);
or U7563 (N_7563,N_7336,N_7362);
nand U7564 (N_7564,N_7230,N_7393);
nor U7565 (N_7565,N_7297,N_7328);
nand U7566 (N_7566,N_7269,N_7275);
xor U7567 (N_7567,N_7325,N_7349);
nand U7568 (N_7568,N_7307,N_7265);
xnor U7569 (N_7569,N_7380,N_7275);
and U7570 (N_7570,N_7387,N_7286);
xnor U7571 (N_7571,N_7230,N_7213);
or U7572 (N_7572,N_7241,N_7323);
and U7573 (N_7573,N_7368,N_7356);
and U7574 (N_7574,N_7307,N_7313);
and U7575 (N_7575,N_7244,N_7375);
or U7576 (N_7576,N_7364,N_7208);
and U7577 (N_7577,N_7342,N_7295);
and U7578 (N_7578,N_7306,N_7242);
and U7579 (N_7579,N_7330,N_7231);
nor U7580 (N_7580,N_7295,N_7392);
or U7581 (N_7581,N_7296,N_7392);
and U7582 (N_7582,N_7320,N_7374);
xor U7583 (N_7583,N_7242,N_7350);
nand U7584 (N_7584,N_7292,N_7334);
nor U7585 (N_7585,N_7298,N_7396);
and U7586 (N_7586,N_7357,N_7321);
xnor U7587 (N_7587,N_7212,N_7261);
and U7588 (N_7588,N_7396,N_7321);
nor U7589 (N_7589,N_7381,N_7380);
xor U7590 (N_7590,N_7380,N_7370);
or U7591 (N_7591,N_7215,N_7250);
and U7592 (N_7592,N_7245,N_7260);
and U7593 (N_7593,N_7215,N_7204);
and U7594 (N_7594,N_7220,N_7353);
xor U7595 (N_7595,N_7216,N_7319);
or U7596 (N_7596,N_7212,N_7287);
xor U7597 (N_7597,N_7310,N_7284);
and U7598 (N_7598,N_7348,N_7329);
xor U7599 (N_7599,N_7304,N_7221);
nand U7600 (N_7600,N_7578,N_7436);
and U7601 (N_7601,N_7585,N_7408);
and U7602 (N_7602,N_7583,N_7596);
nand U7603 (N_7603,N_7444,N_7594);
xnor U7604 (N_7604,N_7454,N_7524);
nand U7605 (N_7605,N_7491,N_7402);
nor U7606 (N_7606,N_7564,N_7477);
xnor U7607 (N_7607,N_7409,N_7472);
or U7608 (N_7608,N_7542,N_7465);
xor U7609 (N_7609,N_7495,N_7514);
or U7610 (N_7610,N_7410,N_7414);
xnor U7611 (N_7611,N_7516,N_7582);
nand U7612 (N_7612,N_7430,N_7561);
and U7613 (N_7613,N_7401,N_7577);
nand U7614 (N_7614,N_7486,N_7494);
xnor U7615 (N_7615,N_7441,N_7425);
nand U7616 (N_7616,N_7534,N_7433);
and U7617 (N_7617,N_7499,N_7469);
nor U7618 (N_7618,N_7558,N_7566);
xor U7619 (N_7619,N_7569,N_7550);
or U7620 (N_7620,N_7413,N_7576);
nand U7621 (N_7621,N_7515,N_7573);
nand U7622 (N_7622,N_7503,N_7468);
or U7623 (N_7623,N_7467,N_7497);
xnor U7624 (N_7624,N_7431,N_7562);
nand U7625 (N_7625,N_7405,N_7533);
or U7626 (N_7626,N_7547,N_7443);
nor U7627 (N_7627,N_7590,N_7529);
xnor U7628 (N_7628,N_7537,N_7543);
or U7629 (N_7629,N_7531,N_7521);
or U7630 (N_7630,N_7442,N_7449);
and U7631 (N_7631,N_7571,N_7451);
and U7632 (N_7632,N_7522,N_7539);
or U7633 (N_7633,N_7427,N_7555);
nor U7634 (N_7634,N_7510,N_7496);
and U7635 (N_7635,N_7591,N_7584);
nor U7636 (N_7636,N_7593,N_7538);
and U7637 (N_7637,N_7567,N_7581);
nor U7638 (N_7638,N_7570,N_7453);
xor U7639 (N_7639,N_7508,N_7504);
and U7640 (N_7640,N_7525,N_7492);
nor U7641 (N_7641,N_7455,N_7528);
xor U7642 (N_7642,N_7426,N_7520);
xnor U7643 (N_7643,N_7461,N_7517);
nand U7644 (N_7644,N_7511,N_7456);
or U7645 (N_7645,N_7588,N_7490);
or U7646 (N_7646,N_7415,N_7400);
nor U7647 (N_7647,N_7519,N_7450);
nand U7648 (N_7648,N_7458,N_7485);
nor U7649 (N_7649,N_7432,N_7404);
or U7650 (N_7650,N_7505,N_7556);
or U7651 (N_7651,N_7423,N_7471);
and U7652 (N_7652,N_7575,N_7587);
and U7653 (N_7653,N_7563,N_7478);
nor U7654 (N_7654,N_7448,N_7476);
or U7655 (N_7655,N_7435,N_7483);
and U7656 (N_7656,N_7509,N_7438);
nor U7657 (N_7657,N_7502,N_7464);
nand U7658 (N_7658,N_7463,N_7560);
or U7659 (N_7659,N_7473,N_7457);
nor U7660 (N_7660,N_7545,N_7437);
and U7661 (N_7661,N_7549,N_7552);
nand U7662 (N_7662,N_7507,N_7527);
and U7663 (N_7663,N_7480,N_7479);
or U7664 (N_7664,N_7407,N_7532);
and U7665 (N_7665,N_7523,N_7541);
nand U7666 (N_7666,N_7406,N_7422);
xor U7667 (N_7667,N_7459,N_7416);
and U7668 (N_7668,N_7548,N_7429);
or U7669 (N_7669,N_7421,N_7540);
xor U7670 (N_7670,N_7482,N_7474);
nand U7671 (N_7671,N_7452,N_7513);
and U7672 (N_7672,N_7554,N_7418);
or U7673 (N_7673,N_7411,N_7498);
nor U7674 (N_7674,N_7428,N_7530);
nor U7675 (N_7675,N_7544,N_7470);
nand U7676 (N_7676,N_7481,N_7501);
or U7677 (N_7677,N_7493,N_7417);
nand U7678 (N_7678,N_7518,N_7589);
xnor U7679 (N_7679,N_7599,N_7489);
nor U7680 (N_7680,N_7551,N_7598);
xnor U7681 (N_7681,N_7572,N_7500);
xnor U7682 (N_7682,N_7412,N_7559);
and U7683 (N_7683,N_7488,N_7475);
xnor U7684 (N_7684,N_7565,N_7595);
nor U7685 (N_7685,N_7446,N_7466);
and U7686 (N_7686,N_7440,N_7424);
or U7687 (N_7687,N_7592,N_7546);
nor U7688 (N_7688,N_7447,N_7574);
or U7689 (N_7689,N_7553,N_7484);
and U7690 (N_7690,N_7568,N_7420);
or U7691 (N_7691,N_7536,N_7445);
or U7692 (N_7692,N_7535,N_7434);
and U7693 (N_7693,N_7419,N_7462);
xor U7694 (N_7694,N_7597,N_7586);
nand U7695 (N_7695,N_7506,N_7403);
nor U7696 (N_7696,N_7512,N_7487);
and U7697 (N_7697,N_7526,N_7460);
and U7698 (N_7698,N_7557,N_7579);
or U7699 (N_7699,N_7439,N_7580);
nor U7700 (N_7700,N_7426,N_7552);
nand U7701 (N_7701,N_7499,N_7444);
nand U7702 (N_7702,N_7484,N_7528);
xor U7703 (N_7703,N_7588,N_7545);
or U7704 (N_7704,N_7556,N_7598);
or U7705 (N_7705,N_7568,N_7505);
and U7706 (N_7706,N_7425,N_7533);
nor U7707 (N_7707,N_7517,N_7498);
xor U7708 (N_7708,N_7594,N_7544);
xor U7709 (N_7709,N_7422,N_7578);
or U7710 (N_7710,N_7431,N_7591);
or U7711 (N_7711,N_7402,N_7443);
nor U7712 (N_7712,N_7511,N_7589);
xnor U7713 (N_7713,N_7571,N_7540);
xnor U7714 (N_7714,N_7531,N_7551);
and U7715 (N_7715,N_7567,N_7481);
nor U7716 (N_7716,N_7452,N_7587);
nand U7717 (N_7717,N_7547,N_7407);
or U7718 (N_7718,N_7595,N_7509);
xor U7719 (N_7719,N_7426,N_7401);
or U7720 (N_7720,N_7410,N_7456);
and U7721 (N_7721,N_7468,N_7477);
and U7722 (N_7722,N_7467,N_7585);
or U7723 (N_7723,N_7480,N_7477);
nor U7724 (N_7724,N_7420,N_7560);
nor U7725 (N_7725,N_7501,N_7454);
nor U7726 (N_7726,N_7482,N_7505);
nand U7727 (N_7727,N_7546,N_7480);
nand U7728 (N_7728,N_7444,N_7410);
nor U7729 (N_7729,N_7556,N_7440);
nand U7730 (N_7730,N_7513,N_7557);
or U7731 (N_7731,N_7569,N_7449);
xor U7732 (N_7732,N_7408,N_7489);
xor U7733 (N_7733,N_7573,N_7504);
xor U7734 (N_7734,N_7526,N_7502);
and U7735 (N_7735,N_7421,N_7417);
nand U7736 (N_7736,N_7407,N_7461);
nor U7737 (N_7737,N_7549,N_7598);
nor U7738 (N_7738,N_7550,N_7590);
and U7739 (N_7739,N_7566,N_7563);
nor U7740 (N_7740,N_7528,N_7576);
or U7741 (N_7741,N_7410,N_7475);
or U7742 (N_7742,N_7556,N_7483);
nand U7743 (N_7743,N_7418,N_7577);
nor U7744 (N_7744,N_7465,N_7552);
or U7745 (N_7745,N_7455,N_7520);
nand U7746 (N_7746,N_7411,N_7471);
nand U7747 (N_7747,N_7439,N_7411);
and U7748 (N_7748,N_7463,N_7449);
xnor U7749 (N_7749,N_7428,N_7450);
or U7750 (N_7750,N_7506,N_7407);
nand U7751 (N_7751,N_7521,N_7508);
or U7752 (N_7752,N_7475,N_7480);
xor U7753 (N_7753,N_7410,N_7543);
and U7754 (N_7754,N_7423,N_7489);
xor U7755 (N_7755,N_7497,N_7413);
or U7756 (N_7756,N_7564,N_7503);
and U7757 (N_7757,N_7493,N_7483);
nor U7758 (N_7758,N_7529,N_7592);
nor U7759 (N_7759,N_7433,N_7532);
nor U7760 (N_7760,N_7523,N_7558);
or U7761 (N_7761,N_7503,N_7551);
nor U7762 (N_7762,N_7461,N_7441);
nor U7763 (N_7763,N_7569,N_7492);
xnor U7764 (N_7764,N_7460,N_7515);
nor U7765 (N_7765,N_7430,N_7475);
or U7766 (N_7766,N_7486,N_7441);
nand U7767 (N_7767,N_7582,N_7517);
nor U7768 (N_7768,N_7408,N_7574);
xnor U7769 (N_7769,N_7406,N_7441);
xor U7770 (N_7770,N_7488,N_7577);
and U7771 (N_7771,N_7598,N_7543);
nor U7772 (N_7772,N_7529,N_7472);
or U7773 (N_7773,N_7472,N_7451);
or U7774 (N_7774,N_7587,N_7442);
and U7775 (N_7775,N_7514,N_7581);
and U7776 (N_7776,N_7554,N_7439);
or U7777 (N_7777,N_7593,N_7535);
nand U7778 (N_7778,N_7406,N_7469);
and U7779 (N_7779,N_7564,N_7412);
nor U7780 (N_7780,N_7450,N_7462);
nand U7781 (N_7781,N_7579,N_7422);
and U7782 (N_7782,N_7575,N_7558);
and U7783 (N_7783,N_7520,N_7414);
xor U7784 (N_7784,N_7455,N_7587);
xnor U7785 (N_7785,N_7549,N_7479);
and U7786 (N_7786,N_7582,N_7462);
or U7787 (N_7787,N_7549,N_7451);
xor U7788 (N_7788,N_7424,N_7462);
xnor U7789 (N_7789,N_7522,N_7489);
nand U7790 (N_7790,N_7481,N_7432);
and U7791 (N_7791,N_7453,N_7415);
nand U7792 (N_7792,N_7404,N_7421);
and U7793 (N_7793,N_7560,N_7430);
and U7794 (N_7794,N_7453,N_7593);
or U7795 (N_7795,N_7542,N_7489);
nand U7796 (N_7796,N_7585,N_7509);
nand U7797 (N_7797,N_7439,N_7538);
or U7798 (N_7798,N_7497,N_7484);
or U7799 (N_7799,N_7405,N_7584);
and U7800 (N_7800,N_7635,N_7763);
xnor U7801 (N_7801,N_7717,N_7722);
or U7802 (N_7802,N_7666,N_7652);
nand U7803 (N_7803,N_7795,N_7607);
nand U7804 (N_7804,N_7703,N_7742);
nor U7805 (N_7805,N_7725,N_7641);
and U7806 (N_7806,N_7656,N_7748);
nand U7807 (N_7807,N_7674,N_7749);
or U7808 (N_7808,N_7788,N_7659);
xor U7809 (N_7809,N_7636,N_7649);
xnor U7810 (N_7810,N_7610,N_7690);
nor U7811 (N_7811,N_7713,N_7790);
nand U7812 (N_7812,N_7664,N_7798);
nor U7813 (N_7813,N_7732,N_7768);
nor U7814 (N_7814,N_7718,N_7716);
xnor U7815 (N_7815,N_7601,N_7612);
nand U7816 (N_7816,N_7743,N_7619);
and U7817 (N_7817,N_7632,N_7724);
or U7818 (N_7818,N_7694,N_7657);
nor U7819 (N_7819,N_7786,N_7627);
nand U7820 (N_7820,N_7726,N_7730);
nor U7821 (N_7821,N_7762,N_7735);
nor U7822 (N_7822,N_7665,N_7617);
or U7823 (N_7823,N_7746,N_7775);
xnor U7824 (N_7824,N_7611,N_7728);
nand U7825 (N_7825,N_7797,N_7731);
and U7826 (N_7826,N_7643,N_7661);
xnor U7827 (N_7827,N_7751,N_7624);
or U7828 (N_7828,N_7729,N_7692);
or U7829 (N_7829,N_7700,N_7626);
xnor U7830 (N_7830,N_7616,N_7648);
nand U7831 (N_7831,N_7785,N_7638);
nor U7832 (N_7832,N_7630,N_7660);
xnor U7833 (N_7833,N_7633,N_7782);
xor U7834 (N_7834,N_7758,N_7625);
xnor U7835 (N_7835,N_7734,N_7608);
nand U7836 (N_7836,N_7675,N_7738);
or U7837 (N_7837,N_7655,N_7774);
nor U7838 (N_7838,N_7688,N_7764);
nand U7839 (N_7839,N_7777,N_7760);
xnor U7840 (N_7840,N_7752,N_7676);
nand U7841 (N_7841,N_7693,N_7642);
and U7842 (N_7842,N_7698,N_7712);
nand U7843 (N_7843,N_7702,N_7677);
nand U7844 (N_7844,N_7714,N_7631);
and U7845 (N_7845,N_7680,N_7793);
nand U7846 (N_7846,N_7791,N_7723);
nand U7847 (N_7847,N_7720,N_7622);
nor U7848 (N_7848,N_7685,N_7678);
nor U7849 (N_7849,N_7697,N_7747);
nor U7850 (N_7850,N_7600,N_7647);
nor U7851 (N_7851,N_7603,N_7629);
nor U7852 (N_7852,N_7606,N_7668);
nor U7853 (N_7853,N_7789,N_7778);
nand U7854 (N_7854,N_7662,N_7766);
and U7855 (N_7855,N_7770,N_7645);
xor U7856 (N_7856,N_7640,N_7695);
xor U7857 (N_7857,N_7715,N_7709);
xnor U7858 (N_7858,N_7672,N_7745);
nor U7859 (N_7859,N_7651,N_7609);
nor U7860 (N_7860,N_7759,N_7799);
xnor U7861 (N_7861,N_7781,N_7621);
nand U7862 (N_7862,N_7605,N_7771);
nor U7863 (N_7863,N_7634,N_7744);
xnor U7864 (N_7864,N_7684,N_7754);
nor U7865 (N_7865,N_7761,N_7604);
nor U7866 (N_7866,N_7701,N_7773);
nand U7867 (N_7867,N_7721,N_7740);
xnor U7868 (N_7868,N_7658,N_7699);
nor U7869 (N_7869,N_7787,N_7769);
and U7870 (N_7870,N_7739,N_7757);
or U7871 (N_7871,N_7708,N_7727);
xnor U7872 (N_7872,N_7615,N_7620);
nand U7873 (N_7873,N_7671,N_7669);
or U7874 (N_7874,N_7779,N_7602);
nand U7875 (N_7875,N_7696,N_7719);
nand U7876 (N_7876,N_7737,N_7767);
or U7877 (N_7877,N_7654,N_7673);
or U7878 (N_7878,N_7689,N_7772);
nor U7879 (N_7879,N_7613,N_7683);
and U7880 (N_7880,N_7637,N_7670);
nand U7881 (N_7881,N_7796,N_7750);
or U7882 (N_7882,N_7618,N_7780);
xor U7883 (N_7883,N_7794,N_7755);
nand U7884 (N_7884,N_7765,N_7733);
and U7885 (N_7885,N_7628,N_7736);
or U7886 (N_7886,N_7711,N_7682);
and U7887 (N_7887,N_7784,N_7667);
nand U7888 (N_7888,N_7639,N_7686);
nor U7889 (N_7889,N_7783,N_7704);
nand U7890 (N_7890,N_7691,N_7653);
nand U7891 (N_7891,N_7644,N_7705);
nand U7892 (N_7892,N_7776,N_7646);
nor U7893 (N_7893,N_7663,N_7741);
or U7894 (N_7894,N_7710,N_7681);
nor U7895 (N_7895,N_7753,N_7623);
nand U7896 (N_7896,N_7707,N_7679);
nand U7897 (N_7897,N_7706,N_7792);
or U7898 (N_7898,N_7756,N_7614);
xor U7899 (N_7899,N_7650,N_7687);
nand U7900 (N_7900,N_7724,N_7764);
and U7901 (N_7901,N_7720,N_7626);
nand U7902 (N_7902,N_7798,N_7734);
xor U7903 (N_7903,N_7727,N_7776);
xor U7904 (N_7904,N_7786,N_7750);
and U7905 (N_7905,N_7701,N_7722);
and U7906 (N_7906,N_7689,N_7765);
xnor U7907 (N_7907,N_7788,N_7653);
xnor U7908 (N_7908,N_7695,N_7766);
xor U7909 (N_7909,N_7633,N_7620);
nand U7910 (N_7910,N_7778,N_7758);
xor U7911 (N_7911,N_7669,N_7785);
nor U7912 (N_7912,N_7690,N_7784);
xor U7913 (N_7913,N_7689,N_7735);
xor U7914 (N_7914,N_7692,N_7753);
nor U7915 (N_7915,N_7642,N_7703);
and U7916 (N_7916,N_7795,N_7721);
and U7917 (N_7917,N_7749,N_7773);
xor U7918 (N_7918,N_7695,N_7646);
and U7919 (N_7919,N_7640,N_7633);
xor U7920 (N_7920,N_7776,N_7640);
and U7921 (N_7921,N_7739,N_7667);
nor U7922 (N_7922,N_7656,N_7631);
xor U7923 (N_7923,N_7737,N_7747);
and U7924 (N_7924,N_7622,N_7787);
nor U7925 (N_7925,N_7740,N_7774);
nor U7926 (N_7926,N_7647,N_7683);
nor U7927 (N_7927,N_7729,N_7784);
xnor U7928 (N_7928,N_7627,N_7666);
nand U7929 (N_7929,N_7697,N_7726);
xnor U7930 (N_7930,N_7639,N_7795);
and U7931 (N_7931,N_7674,N_7646);
xor U7932 (N_7932,N_7619,N_7740);
and U7933 (N_7933,N_7778,N_7647);
nand U7934 (N_7934,N_7767,N_7617);
nand U7935 (N_7935,N_7671,N_7729);
nor U7936 (N_7936,N_7726,N_7660);
xor U7937 (N_7937,N_7625,N_7612);
nand U7938 (N_7938,N_7664,N_7720);
nand U7939 (N_7939,N_7792,N_7757);
or U7940 (N_7940,N_7655,N_7661);
and U7941 (N_7941,N_7636,N_7655);
xnor U7942 (N_7942,N_7763,N_7739);
xor U7943 (N_7943,N_7642,N_7696);
nor U7944 (N_7944,N_7657,N_7791);
and U7945 (N_7945,N_7798,N_7695);
and U7946 (N_7946,N_7631,N_7712);
nand U7947 (N_7947,N_7710,N_7670);
nor U7948 (N_7948,N_7674,N_7642);
and U7949 (N_7949,N_7623,N_7788);
nor U7950 (N_7950,N_7753,N_7729);
nor U7951 (N_7951,N_7794,N_7735);
or U7952 (N_7952,N_7611,N_7751);
and U7953 (N_7953,N_7761,N_7628);
and U7954 (N_7954,N_7647,N_7689);
or U7955 (N_7955,N_7668,N_7762);
nor U7956 (N_7956,N_7601,N_7653);
nand U7957 (N_7957,N_7627,N_7642);
and U7958 (N_7958,N_7609,N_7719);
or U7959 (N_7959,N_7633,N_7662);
xor U7960 (N_7960,N_7725,N_7683);
nand U7961 (N_7961,N_7702,N_7681);
or U7962 (N_7962,N_7640,N_7611);
xnor U7963 (N_7963,N_7780,N_7670);
xor U7964 (N_7964,N_7640,N_7798);
and U7965 (N_7965,N_7683,N_7787);
xnor U7966 (N_7966,N_7706,N_7680);
and U7967 (N_7967,N_7795,N_7789);
xor U7968 (N_7968,N_7663,N_7772);
nand U7969 (N_7969,N_7751,N_7650);
and U7970 (N_7970,N_7682,N_7693);
nand U7971 (N_7971,N_7776,N_7736);
and U7972 (N_7972,N_7604,N_7610);
nand U7973 (N_7973,N_7718,N_7633);
and U7974 (N_7974,N_7716,N_7687);
nand U7975 (N_7975,N_7611,N_7726);
nand U7976 (N_7976,N_7748,N_7666);
or U7977 (N_7977,N_7735,N_7684);
or U7978 (N_7978,N_7690,N_7780);
nand U7979 (N_7979,N_7685,N_7627);
or U7980 (N_7980,N_7669,N_7759);
and U7981 (N_7981,N_7789,N_7702);
nor U7982 (N_7982,N_7643,N_7736);
xor U7983 (N_7983,N_7628,N_7617);
and U7984 (N_7984,N_7665,N_7608);
nand U7985 (N_7985,N_7619,N_7771);
or U7986 (N_7986,N_7717,N_7740);
nor U7987 (N_7987,N_7643,N_7658);
xor U7988 (N_7988,N_7729,N_7764);
xnor U7989 (N_7989,N_7657,N_7640);
nand U7990 (N_7990,N_7683,N_7722);
nand U7991 (N_7991,N_7774,N_7713);
xor U7992 (N_7992,N_7717,N_7688);
and U7993 (N_7993,N_7765,N_7636);
and U7994 (N_7994,N_7626,N_7674);
and U7995 (N_7995,N_7753,N_7612);
and U7996 (N_7996,N_7742,N_7631);
or U7997 (N_7997,N_7693,N_7652);
nand U7998 (N_7998,N_7765,N_7741);
nand U7999 (N_7999,N_7743,N_7621);
and U8000 (N_8000,N_7854,N_7935);
and U8001 (N_8001,N_7818,N_7861);
nor U8002 (N_8002,N_7834,N_7871);
or U8003 (N_8003,N_7940,N_7931);
nor U8004 (N_8004,N_7884,N_7881);
and U8005 (N_8005,N_7900,N_7866);
xor U8006 (N_8006,N_7849,N_7902);
nand U8007 (N_8007,N_7862,N_7949);
or U8008 (N_8008,N_7801,N_7972);
xor U8009 (N_8009,N_7987,N_7872);
nand U8010 (N_8010,N_7805,N_7970);
or U8011 (N_8011,N_7980,N_7858);
xor U8012 (N_8012,N_7901,N_7812);
xor U8013 (N_8013,N_7981,N_7955);
nor U8014 (N_8014,N_7961,N_7994);
nor U8015 (N_8015,N_7963,N_7856);
nor U8016 (N_8016,N_7897,N_7843);
or U8017 (N_8017,N_7847,N_7817);
nor U8018 (N_8018,N_7997,N_7825);
and U8019 (N_8019,N_7879,N_7996);
nand U8020 (N_8020,N_7964,N_7841);
xnor U8021 (N_8021,N_7833,N_7907);
nand U8022 (N_8022,N_7969,N_7877);
or U8023 (N_8023,N_7917,N_7930);
and U8024 (N_8024,N_7808,N_7839);
xor U8025 (N_8025,N_7889,N_7912);
xor U8026 (N_8026,N_7982,N_7903);
and U8027 (N_8027,N_7810,N_7948);
nor U8028 (N_8028,N_7892,N_7971);
and U8029 (N_8029,N_7827,N_7937);
and U8030 (N_8030,N_7814,N_7836);
or U8031 (N_8031,N_7929,N_7837);
nor U8032 (N_8032,N_7842,N_7959);
nor U8033 (N_8033,N_7840,N_7813);
nor U8034 (N_8034,N_7911,N_7956);
xor U8035 (N_8035,N_7922,N_7886);
and U8036 (N_8036,N_7891,N_7983);
xor U8037 (N_8037,N_7976,N_7977);
or U8038 (N_8038,N_7864,N_7893);
xor U8039 (N_8039,N_7979,N_7826);
xnor U8040 (N_8040,N_7890,N_7823);
nor U8041 (N_8041,N_7899,N_7945);
or U8042 (N_8042,N_7925,N_7832);
or U8043 (N_8043,N_7873,N_7906);
nor U8044 (N_8044,N_7820,N_7985);
nor U8045 (N_8045,N_7916,N_7845);
nand U8046 (N_8046,N_7888,N_7848);
and U8047 (N_8047,N_7802,N_7953);
xnor U8048 (N_8048,N_7965,N_7855);
or U8049 (N_8049,N_7860,N_7991);
xor U8050 (N_8050,N_7896,N_7933);
nand U8051 (N_8051,N_7943,N_7992);
nand U8052 (N_8052,N_7821,N_7934);
or U8053 (N_8053,N_7914,N_7824);
xnor U8054 (N_8054,N_7838,N_7904);
nand U8055 (N_8055,N_7830,N_7958);
nand U8056 (N_8056,N_7829,N_7957);
or U8057 (N_8057,N_7804,N_7844);
or U8058 (N_8058,N_7816,N_7942);
nand U8059 (N_8059,N_7898,N_7876);
or U8060 (N_8060,N_7887,N_7946);
or U8061 (N_8061,N_7921,N_7883);
and U8062 (N_8062,N_7993,N_7950);
nor U8063 (N_8063,N_7857,N_7800);
nand U8064 (N_8064,N_7952,N_7869);
xor U8065 (N_8065,N_7870,N_7919);
nor U8066 (N_8066,N_7913,N_7852);
xnor U8067 (N_8067,N_7960,N_7932);
nor U8068 (N_8068,N_7962,N_7999);
nand U8069 (N_8069,N_7998,N_7909);
and U8070 (N_8070,N_7905,N_7924);
nor U8071 (N_8071,N_7809,N_7926);
or U8072 (N_8072,N_7974,N_7910);
and U8073 (N_8073,N_7859,N_7895);
nor U8074 (N_8074,N_7915,N_7851);
nor U8075 (N_8075,N_7967,N_7865);
nand U8076 (N_8076,N_7988,N_7989);
nand U8077 (N_8077,N_7885,N_7975);
nor U8078 (N_8078,N_7863,N_7894);
nor U8079 (N_8079,N_7966,N_7986);
xnor U8080 (N_8080,N_7846,N_7868);
xnor U8081 (N_8081,N_7828,N_7938);
and U8082 (N_8082,N_7878,N_7923);
nand U8083 (N_8083,N_7968,N_7927);
nand U8084 (N_8084,N_7875,N_7954);
nand U8085 (N_8085,N_7984,N_7867);
nand U8086 (N_8086,N_7880,N_7908);
or U8087 (N_8087,N_7806,N_7815);
xor U8088 (N_8088,N_7990,N_7947);
xnor U8089 (N_8089,N_7803,N_7995);
and U8090 (N_8090,N_7882,N_7928);
or U8091 (N_8091,N_7874,N_7951);
or U8092 (N_8092,N_7918,N_7936);
or U8093 (N_8093,N_7939,N_7973);
nor U8094 (N_8094,N_7831,N_7920);
xor U8095 (N_8095,N_7978,N_7850);
nand U8096 (N_8096,N_7853,N_7944);
xor U8097 (N_8097,N_7807,N_7819);
xor U8098 (N_8098,N_7941,N_7835);
nor U8099 (N_8099,N_7811,N_7822);
or U8100 (N_8100,N_7981,N_7954);
nand U8101 (N_8101,N_7922,N_7906);
nand U8102 (N_8102,N_7806,N_7826);
or U8103 (N_8103,N_7828,N_7851);
and U8104 (N_8104,N_7956,N_7915);
and U8105 (N_8105,N_7872,N_7910);
nand U8106 (N_8106,N_7862,N_7838);
xnor U8107 (N_8107,N_7882,N_7902);
nor U8108 (N_8108,N_7801,N_7983);
xnor U8109 (N_8109,N_7839,N_7820);
nand U8110 (N_8110,N_7945,N_7908);
or U8111 (N_8111,N_7810,N_7942);
xnor U8112 (N_8112,N_7839,N_7960);
nand U8113 (N_8113,N_7897,N_7976);
xor U8114 (N_8114,N_7869,N_7841);
xor U8115 (N_8115,N_7812,N_7905);
or U8116 (N_8116,N_7813,N_7906);
and U8117 (N_8117,N_7974,N_7972);
or U8118 (N_8118,N_7861,N_7800);
xnor U8119 (N_8119,N_7824,N_7816);
or U8120 (N_8120,N_7969,N_7910);
and U8121 (N_8121,N_7966,N_7948);
or U8122 (N_8122,N_7834,N_7917);
nand U8123 (N_8123,N_7948,N_7951);
and U8124 (N_8124,N_7816,N_7863);
or U8125 (N_8125,N_7909,N_7866);
and U8126 (N_8126,N_7868,N_7879);
and U8127 (N_8127,N_7810,N_7867);
xnor U8128 (N_8128,N_7912,N_7923);
nand U8129 (N_8129,N_7924,N_7823);
nor U8130 (N_8130,N_7929,N_7828);
and U8131 (N_8131,N_7823,N_7944);
and U8132 (N_8132,N_7956,N_7932);
xor U8133 (N_8133,N_7926,N_7965);
and U8134 (N_8134,N_7968,N_7811);
nand U8135 (N_8135,N_7836,N_7930);
xor U8136 (N_8136,N_7863,N_7866);
nand U8137 (N_8137,N_7910,N_7916);
nand U8138 (N_8138,N_7808,N_7821);
and U8139 (N_8139,N_7816,N_7904);
or U8140 (N_8140,N_7886,N_7952);
nor U8141 (N_8141,N_7962,N_7869);
xor U8142 (N_8142,N_7932,N_7831);
xnor U8143 (N_8143,N_7901,N_7954);
nor U8144 (N_8144,N_7855,N_7974);
nor U8145 (N_8145,N_7893,N_7999);
and U8146 (N_8146,N_7894,N_7856);
nor U8147 (N_8147,N_7886,N_7925);
and U8148 (N_8148,N_7939,N_7952);
and U8149 (N_8149,N_7885,N_7862);
nand U8150 (N_8150,N_7945,N_7915);
xnor U8151 (N_8151,N_7894,N_7845);
and U8152 (N_8152,N_7801,N_7892);
nand U8153 (N_8153,N_7901,N_7933);
or U8154 (N_8154,N_7902,N_7924);
nor U8155 (N_8155,N_7867,N_7958);
or U8156 (N_8156,N_7906,N_7981);
nand U8157 (N_8157,N_7806,N_7822);
xnor U8158 (N_8158,N_7880,N_7877);
or U8159 (N_8159,N_7998,N_7898);
and U8160 (N_8160,N_7877,N_7821);
nand U8161 (N_8161,N_7924,N_7860);
nand U8162 (N_8162,N_7933,N_7978);
nor U8163 (N_8163,N_7830,N_7966);
nor U8164 (N_8164,N_7967,N_7992);
and U8165 (N_8165,N_7978,N_7973);
and U8166 (N_8166,N_7839,N_7895);
or U8167 (N_8167,N_7925,N_7819);
xor U8168 (N_8168,N_7999,N_7978);
xnor U8169 (N_8169,N_7804,N_7903);
xor U8170 (N_8170,N_7808,N_7836);
nand U8171 (N_8171,N_7941,N_7999);
and U8172 (N_8172,N_7957,N_7907);
or U8173 (N_8173,N_7976,N_7962);
and U8174 (N_8174,N_7804,N_7967);
nand U8175 (N_8175,N_7876,N_7991);
nand U8176 (N_8176,N_7810,N_7959);
nand U8177 (N_8177,N_7916,N_7920);
and U8178 (N_8178,N_7970,N_7816);
and U8179 (N_8179,N_7925,N_7908);
and U8180 (N_8180,N_7941,N_7833);
nand U8181 (N_8181,N_7814,N_7891);
and U8182 (N_8182,N_7833,N_7911);
and U8183 (N_8183,N_7939,N_7948);
nand U8184 (N_8184,N_7807,N_7997);
nand U8185 (N_8185,N_7970,N_7971);
or U8186 (N_8186,N_7991,N_7937);
and U8187 (N_8187,N_7928,N_7935);
or U8188 (N_8188,N_7919,N_7854);
nand U8189 (N_8189,N_7916,N_7931);
nor U8190 (N_8190,N_7884,N_7893);
or U8191 (N_8191,N_7903,N_7809);
or U8192 (N_8192,N_7827,N_7899);
nand U8193 (N_8193,N_7963,N_7860);
or U8194 (N_8194,N_7886,N_7803);
nand U8195 (N_8195,N_7996,N_7928);
or U8196 (N_8196,N_7809,N_7855);
xnor U8197 (N_8197,N_7942,N_7979);
and U8198 (N_8198,N_7837,N_7980);
xor U8199 (N_8199,N_7892,N_7937);
nand U8200 (N_8200,N_8140,N_8120);
or U8201 (N_8201,N_8131,N_8130);
nand U8202 (N_8202,N_8137,N_8191);
xnor U8203 (N_8203,N_8157,N_8171);
xor U8204 (N_8204,N_8155,N_8142);
nor U8205 (N_8205,N_8153,N_8156);
and U8206 (N_8206,N_8098,N_8065);
or U8207 (N_8207,N_8049,N_8112);
xnor U8208 (N_8208,N_8020,N_8177);
xor U8209 (N_8209,N_8044,N_8113);
and U8210 (N_8210,N_8135,N_8041);
nand U8211 (N_8211,N_8022,N_8192);
xnor U8212 (N_8212,N_8062,N_8176);
nor U8213 (N_8213,N_8015,N_8076);
xnor U8214 (N_8214,N_8073,N_8045);
and U8215 (N_8215,N_8111,N_8057);
and U8216 (N_8216,N_8084,N_8165);
nand U8217 (N_8217,N_8000,N_8081);
xnor U8218 (N_8218,N_8121,N_8188);
nand U8219 (N_8219,N_8037,N_8096);
or U8220 (N_8220,N_8043,N_8028);
or U8221 (N_8221,N_8152,N_8128);
or U8222 (N_8222,N_8054,N_8150);
nor U8223 (N_8223,N_8019,N_8039);
xnor U8224 (N_8224,N_8197,N_8116);
nor U8225 (N_8225,N_8129,N_8125);
nand U8226 (N_8226,N_8115,N_8136);
nor U8227 (N_8227,N_8173,N_8048);
or U8228 (N_8228,N_8161,N_8051);
nand U8229 (N_8229,N_8091,N_8080);
xnor U8230 (N_8230,N_8029,N_8069);
nand U8231 (N_8231,N_8074,N_8196);
xnor U8232 (N_8232,N_8053,N_8033);
nor U8233 (N_8233,N_8127,N_8148);
xor U8234 (N_8234,N_8035,N_8059);
or U8235 (N_8235,N_8169,N_8175);
or U8236 (N_8236,N_8042,N_8182);
nor U8237 (N_8237,N_8187,N_8193);
nor U8238 (N_8238,N_8031,N_8003);
nor U8239 (N_8239,N_8070,N_8164);
nor U8240 (N_8240,N_8174,N_8160);
nand U8241 (N_8241,N_8021,N_8077);
and U8242 (N_8242,N_8198,N_8141);
or U8243 (N_8243,N_8145,N_8009);
nand U8244 (N_8244,N_8027,N_8016);
and U8245 (N_8245,N_8154,N_8168);
xor U8246 (N_8246,N_8109,N_8058);
xor U8247 (N_8247,N_8002,N_8184);
nor U8248 (N_8248,N_8122,N_8163);
nor U8249 (N_8249,N_8133,N_8101);
nor U8250 (N_8250,N_8063,N_8170);
nor U8251 (N_8251,N_8099,N_8088);
and U8252 (N_8252,N_8146,N_8186);
or U8253 (N_8253,N_8066,N_8167);
and U8254 (N_8254,N_8090,N_8159);
and U8255 (N_8255,N_8071,N_8026);
nand U8256 (N_8256,N_8106,N_8083);
and U8257 (N_8257,N_8036,N_8014);
and U8258 (N_8258,N_8194,N_8006);
or U8259 (N_8259,N_8107,N_8189);
nand U8260 (N_8260,N_8185,N_8134);
nor U8261 (N_8261,N_8199,N_8147);
nor U8262 (N_8262,N_8007,N_8190);
nand U8263 (N_8263,N_8183,N_8105);
nor U8264 (N_8264,N_8038,N_8005);
xnor U8265 (N_8265,N_8060,N_8004);
or U8266 (N_8266,N_8102,N_8072);
nand U8267 (N_8267,N_8013,N_8166);
nand U8268 (N_8268,N_8126,N_8047);
or U8269 (N_8269,N_8138,N_8158);
and U8270 (N_8270,N_8162,N_8095);
nor U8271 (N_8271,N_8100,N_8144);
nand U8272 (N_8272,N_8087,N_8024);
or U8273 (N_8273,N_8011,N_8079);
or U8274 (N_8274,N_8075,N_8017);
nand U8275 (N_8275,N_8108,N_8119);
nor U8276 (N_8276,N_8117,N_8180);
and U8277 (N_8277,N_8132,N_8181);
nor U8278 (N_8278,N_8118,N_8068);
nand U8279 (N_8279,N_8178,N_8110);
nand U8280 (N_8280,N_8052,N_8114);
nand U8281 (N_8281,N_8061,N_8018);
nand U8282 (N_8282,N_8012,N_8008);
nor U8283 (N_8283,N_8195,N_8032);
and U8284 (N_8284,N_8034,N_8025);
xor U8285 (N_8285,N_8123,N_8104);
nand U8286 (N_8286,N_8086,N_8124);
nand U8287 (N_8287,N_8064,N_8092);
nand U8288 (N_8288,N_8078,N_8093);
nand U8289 (N_8289,N_8094,N_8055);
nand U8290 (N_8290,N_8040,N_8172);
or U8291 (N_8291,N_8089,N_8097);
nor U8292 (N_8292,N_8010,N_8085);
nand U8293 (N_8293,N_8046,N_8030);
and U8294 (N_8294,N_8151,N_8067);
or U8295 (N_8295,N_8023,N_8149);
xor U8296 (N_8296,N_8050,N_8143);
xnor U8297 (N_8297,N_8056,N_8082);
or U8298 (N_8298,N_8139,N_8103);
nor U8299 (N_8299,N_8001,N_8179);
nand U8300 (N_8300,N_8074,N_8147);
xor U8301 (N_8301,N_8112,N_8044);
nand U8302 (N_8302,N_8074,N_8014);
nor U8303 (N_8303,N_8047,N_8004);
nand U8304 (N_8304,N_8174,N_8080);
or U8305 (N_8305,N_8152,N_8055);
xnor U8306 (N_8306,N_8154,N_8128);
xor U8307 (N_8307,N_8171,N_8019);
nor U8308 (N_8308,N_8149,N_8178);
and U8309 (N_8309,N_8197,N_8018);
and U8310 (N_8310,N_8055,N_8124);
xnor U8311 (N_8311,N_8150,N_8049);
nor U8312 (N_8312,N_8161,N_8000);
xor U8313 (N_8313,N_8150,N_8153);
nand U8314 (N_8314,N_8033,N_8030);
xor U8315 (N_8315,N_8092,N_8054);
nor U8316 (N_8316,N_8039,N_8080);
nand U8317 (N_8317,N_8037,N_8196);
nand U8318 (N_8318,N_8043,N_8134);
nor U8319 (N_8319,N_8127,N_8149);
nand U8320 (N_8320,N_8101,N_8068);
nor U8321 (N_8321,N_8099,N_8066);
or U8322 (N_8322,N_8130,N_8177);
and U8323 (N_8323,N_8084,N_8006);
nor U8324 (N_8324,N_8156,N_8101);
or U8325 (N_8325,N_8046,N_8117);
and U8326 (N_8326,N_8131,N_8021);
nand U8327 (N_8327,N_8009,N_8104);
or U8328 (N_8328,N_8199,N_8127);
and U8329 (N_8329,N_8016,N_8078);
xnor U8330 (N_8330,N_8188,N_8028);
nand U8331 (N_8331,N_8126,N_8104);
or U8332 (N_8332,N_8046,N_8193);
and U8333 (N_8333,N_8077,N_8157);
or U8334 (N_8334,N_8006,N_8019);
xor U8335 (N_8335,N_8135,N_8174);
or U8336 (N_8336,N_8146,N_8102);
nand U8337 (N_8337,N_8187,N_8046);
nand U8338 (N_8338,N_8094,N_8052);
and U8339 (N_8339,N_8054,N_8146);
or U8340 (N_8340,N_8091,N_8113);
and U8341 (N_8341,N_8134,N_8198);
nor U8342 (N_8342,N_8124,N_8182);
nor U8343 (N_8343,N_8031,N_8115);
nor U8344 (N_8344,N_8157,N_8101);
xnor U8345 (N_8345,N_8167,N_8084);
nand U8346 (N_8346,N_8098,N_8192);
nor U8347 (N_8347,N_8058,N_8067);
nor U8348 (N_8348,N_8103,N_8149);
or U8349 (N_8349,N_8017,N_8079);
or U8350 (N_8350,N_8090,N_8018);
nor U8351 (N_8351,N_8031,N_8128);
nor U8352 (N_8352,N_8121,N_8047);
xnor U8353 (N_8353,N_8164,N_8009);
nand U8354 (N_8354,N_8124,N_8198);
and U8355 (N_8355,N_8179,N_8199);
nor U8356 (N_8356,N_8175,N_8071);
or U8357 (N_8357,N_8000,N_8051);
nand U8358 (N_8358,N_8149,N_8119);
nand U8359 (N_8359,N_8142,N_8168);
nor U8360 (N_8360,N_8061,N_8053);
nand U8361 (N_8361,N_8103,N_8110);
or U8362 (N_8362,N_8155,N_8177);
or U8363 (N_8363,N_8037,N_8023);
nor U8364 (N_8364,N_8144,N_8032);
and U8365 (N_8365,N_8072,N_8113);
nand U8366 (N_8366,N_8009,N_8092);
or U8367 (N_8367,N_8157,N_8177);
xnor U8368 (N_8368,N_8079,N_8062);
nand U8369 (N_8369,N_8014,N_8162);
and U8370 (N_8370,N_8108,N_8166);
nand U8371 (N_8371,N_8079,N_8139);
nor U8372 (N_8372,N_8094,N_8123);
xor U8373 (N_8373,N_8147,N_8032);
and U8374 (N_8374,N_8083,N_8187);
or U8375 (N_8375,N_8139,N_8071);
nor U8376 (N_8376,N_8043,N_8131);
and U8377 (N_8377,N_8032,N_8070);
or U8378 (N_8378,N_8086,N_8025);
or U8379 (N_8379,N_8019,N_8067);
and U8380 (N_8380,N_8008,N_8079);
xnor U8381 (N_8381,N_8146,N_8007);
xor U8382 (N_8382,N_8022,N_8064);
nand U8383 (N_8383,N_8028,N_8027);
or U8384 (N_8384,N_8034,N_8183);
or U8385 (N_8385,N_8106,N_8012);
and U8386 (N_8386,N_8185,N_8111);
nor U8387 (N_8387,N_8101,N_8013);
nor U8388 (N_8388,N_8081,N_8054);
and U8389 (N_8389,N_8118,N_8087);
xor U8390 (N_8390,N_8043,N_8011);
xnor U8391 (N_8391,N_8174,N_8073);
or U8392 (N_8392,N_8115,N_8005);
or U8393 (N_8393,N_8078,N_8092);
and U8394 (N_8394,N_8154,N_8111);
nor U8395 (N_8395,N_8034,N_8137);
nor U8396 (N_8396,N_8125,N_8036);
nor U8397 (N_8397,N_8027,N_8090);
nand U8398 (N_8398,N_8057,N_8081);
or U8399 (N_8399,N_8034,N_8152);
and U8400 (N_8400,N_8359,N_8210);
nand U8401 (N_8401,N_8254,N_8315);
or U8402 (N_8402,N_8341,N_8287);
or U8403 (N_8403,N_8202,N_8355);
or U8404 (N_8404,N_8395,N_8328);
nand U8405 (N_8405,N_8369,N_8284);
and U8406 (N_8406,N_8267,N_8245);
or U8407 (N_8407,N_8326,N_8277);
xnor U8408 (N_8408,N_8374,N_8244);
nand U8409 (N_8409,N_8218,N_8236);
nand U8410 (N_8410,N_8251,N_8338);
nand U8411 (N_8411,N_8261,N_8331);
xor U8412 (N_8412,N_8292,N_8235);
nor U8413 (N_8413,N_8353,N_8356);
nand U8414 (N_8414,N_8246,N_8376);
or U8415 (N_8415,N_8368,N_8209);
xor U8416 (N_8416,N_8379,N_8345);
nor U8417 (N_8417,N_8213,N_8311);
and U8418 (N_8418,N_8329,N_8257);
or U8419 (N_8419,N_8312,N_8327);
xor U8420 (N_8420,N_8384,N_8208);
nand U8421 (N_8421,N_8296,N_8268);
nand U8422 (N_8422,N_8373,N_8299);
nor U8423 (N_8423,N_8212,N_8260);
xnor U8424 (N_8424,N_8207,N_8222);
xnor U8425 (N_8425,N_8305,N_8200);
and U8426 (N_8426,N_8201,N_8203);
and U8427 (N_8427,N_8351,N_8352);
or U8428 (N_8428,N_8288,N_8383);
nand U8429 (N_8429,N_8286,N_8386);
xnor U8430 (N_8430,N_8274,N_8233);
and U8431 (N_8431,N_8360,N_8364);
and U8432 (N_8432,N_8275,N_8318);
and U8433 (N_8433,N_8221,N_8295);
nor U8434 (N_8434,N_8340,N_8300);
nor U8435 (N_8435,N_8216,N_8324);
nand U8436 (N_8436,N_8332,N_8393);
xnor U8437 (N_8437,N_8371,N_8271);
xnor U8438 (N_8438,N_8224,N_8242);
and U8439 (N_8439,N_8396,N_8265);
nand U8440 (N_8440,N_8323,N_8223);
nor U8441 (N_8441,N_8380,N_8249);
or U8442 (N_8442,N_8301,N_8256);
or U8443 (N_8443,N_8333,N_8297);
xnor U8444 (N_8444,N_8347,N_8298);
and U8445 (N_8445,N_8307,N_8270);
or U8446 (N_8446,N_8308,N_8334);
or U8447 (N_8447,N_8392,N_8217);
nand U8448 (N_8448,N_8316,N_8262);
or U8449 (N_8449,N_8336,N_8399);
xnor U8450 (N_8450,N_8227,N_8349);
nor U8451 (N_8451,N_8258,N_8237);
nand U8452 (N_8452,N_8238,N_8255);
xnor U8453 (N_8453,N_8241,N_8252);
nor U8454 (N_8454,N_8330,N_8240);
or U8455 (N_8455,N_8220,N_8391);
or U8456 (N_8456,N_8322,N_8319);
and U8457 (N_8457,N_8266,N_8219);
nand U8458 (N_8458,N_8234,N_8283);
or U8459 (N_8459,N_8278,N_8304);
or U8460 (N_8460,N_8272,N_8377);
or U8461 (N_8461,N_8358,N_8243);
xor U8462 (N_8462,N_8293,N_8205);
nor U8463 (N_8463,N_8367,N_8206);
or U8464 (N_8464,N_8214,N_8248);
xnor U8465 (N_8465,N_8398,N_8390);
nor U8466 (N_8466,N_8342,N_8344);
or U8467 (N_8467,N_8228,N_8211);
and U8468 (N_8468,N_8276,N_8337);
nand U8469 (N_8469,N_8397,N_8321);
or U8470 (N_8470,N_8361,N_8215);
or U8471 (N_8471,N_8372,N_8282);
nand U8472 (N_8472,N_8230,N_8247);
nor U8473 (N_8473,N_8354,N_8273);
and U8474 (N_8474,N_8285,N_8302);
or U8475 (N_8475,N_8310,N_8314);
and U8476 (N_8476,N_8229,N_8280);
nor U8477 (N_8477,N_8339,N_8350);
or U8478 (N_8478,N_8250,N_8370);
xor U8479 (N_8479,N_8264,N_8313);
nor U8480 (N_8480,N_8263,N_8362);
and U8481 (N_8481,N_8309,N_8290);
or U8482 (N_8482,N_8269,N_8232);
or U8483 (N_8483,N_8385,N_8357);
nor U8484 (N_8484,N_8231,N_8289);
xor U8485 (N_8485,N_8320,N_8363);
xnor U8486 (N_8486,N_8303,N_8306);
or U8487 (N_8487,N_8382,N_8365);
xor U8488 (N_8488,N_8226,N_8291);
xnor U8489 (N_8489,N_8378,N_8366);
nand U8490 (N_8490,N_8348,N_8259);
and U8491 (N_8491,N_8394,N_8387);
nand U8492 (N_8492,N_8346,N_8388);
and U8493 (N_8493,N_8335,N_8389);
nor U8494 (N_8494,N_8317,N_8294);
nor U8495 (N_8495,N_8204,N_8239);
and U8496 (N_8496,N_8325,N_8253);
xor U8497 (N_8497,N_8375,N_8279);
xnor U8498 (N_8498,N_8225,N_8343);
or U8499 (N_8499,N_8281,N_8381);
nand U8500 (N_8500,N_8262,N_8319);
xor U8501 (N_8501,N_8312,N_8230);
nor U8502 (N_8502,N_8311,N_8269);
and U8503 (N_8503,N_8380,N_8255);
and U8504 (N_8504,N_8389,N_8307);
or U8505 (N_8505,N_8312,N_8275);
and U8506 (N_8506,N_8254,N_8370);
nor U8507 (N_8507,N_8200,N_8319);
nand U8508 (N_8508,N_8238,N_8211);
xnor U8509 (N_8509,N_8382,N_8301);
nor U8510 (N_8510,N_8282,N_8313);
nor U8511 (N_8511,N_8371,N_8396);
and U8512 (N_8512,N_8271,N_8341);
nor U8513 (N_8513,N_8395,N_8396);
xor U8514 (N_8514,N_8230,N_8298);
and U8515 (N_8515,N_8243,N_8389);
or U8516 (N_8516,N_8223,N_8287);
or U8517 (N_8517,N_8232,N_8336);
nand U8518 (N_8518,N_8331,N_8324);
or U8519 (N_8519,N_8224,N_8298);
or U8520 (N_8520,N_8238,N_8314);
nor U8521 (N_8521,N_8306,N_8305);
and U8522 (N_8522,N_8206,N_8280);
or U8523 (N_8523,N_8398,N_8370);
and U8524 (N_8524,N_8314,N_8258);
and U8525 (N_8525,N_8202,N_8266);
and U8526 (N_8526,N_8366,N_8384);
and U8527 (N_8527,N_8273,N_8342);
and U8528 (N_8528,N_8337,N_8309);
nand U8529 (N_8529,N_8329,N_8382);
xnor U8530 (N_8530,N_8366,N_8201);
nor U8531 (N_8531,N_8386,N_8246);
nor U8532 (N_8532,N_8212,N_8354);
xor U8533 (N_8533,N_8387,N_8364);
nand U8534 (N_8534,N_8381,N_8288);
nand U8535 (N_8535,N_8292,N_8375);
and U8536 (N_8536,N_8270,N_8268);
nor U8537 (N_8537,N_8277,N_8349);
or U8538 (N_8538,N_8210,N_8242);
nand U8539 (N_8539,N_8233,N_8220);
xnor U8540 (N_8540,N_8218,N_8388);
nor U8541 (N_8541,N_8305,N_8235);
nor U8542 (N_8542,N_8393,N_8216);
nor U8543 (N_8543,N_8269,N_8320);
nor U8544 (N_8544,N_8315,N_8309);
nor U8545 (N_8545,N_8297,N_8387);
xor U8546 (N_8546,N_8250,N_8304);
and U8547 (N_8547,N_8227,N_8245);
xor U8548 (N_8548,N_8257,N_8336);
nor U8549 (N_8549,N_8335,N_8360);
nor U8550 (N_8550,N_8349,N_8325);
nand U8551 (N_8551,N_8304,N_8233);
or U8552 (N_8552,N_8365,N_8275);
and U8553 (N_8553,N_8264,N_8265);
nor U8554 (N_8554,N_8356,N_8287);
or U8555 (N_8555,N_8362,N_8244);
or U8556 (N_8556,N_8222,N_8273);
or U8557 (N_8557,N_8275,N_8279);
or U8558 (N_8558,N_8376,N_8215);
nand U8559 (N_8559,N_8344,N_8325);
and U8560 (N_8560,N_8245,N_8328);
xor U8561 (N_8561,N_8342,N_8260);
or U8562 (N_8562,N_8353,N_8364);
and U8563 (N_8563,N_8318,N_8202);
or U8564 (N_8564,N_8371,N_8274);
nor U8565 (N_8565,N_8258,N_8300);
nor U8566 (N_8566,N_8251,N_8223);
xnor U8567 (N_8567,N_8392,N_8386);
nand U8568 (N_8568,N_8307,N_8212);
xor U8569 (N_8569,N_8204,N_8263);
nand U8570 (N_8570,N_8220,N_8305);
xnor U8571 (N_8571,N_8245,N_8213);
or U8572 (N_8572,N_8370,N_8368);
and U8573 (N_8573,N_8311,N_8233);
or U8574 (N_8574,N_8394,N_8211);
and U8575 (N_8575,N_8207,N_8213);
xnor U8576 (N_8576,N_8326,N_8324);
nand U8577 (N_8577,N_8264,N_8372);
nor U8578 (N_8578,N_8378,N_8372);
xnor U8579 (N_8579,N_8360,N_8260);
xor U8580 (N_8580,N_8230,N_8296);
xnor U8581 (N_8581,N_8314,N_8322);
nand U8582 (N_8582,N_8340,N_8272);
or U8583 (N_8583,N_8218,N_8387);
nor U8584 (N_8584,N_8220,N_8354);
and U8585 (N_8585,N_8274,N_8275);
nor U8586 (N_8586,N_8249,N_8292);
and U8587 (N_8587,N_8225,N_8336);
nand U8588 (N_8588,N_8388,N_8200);
nand U8589 (N_8589,N_8352,N_8305);
xnor U8590 (N_8590,N_8229,N_8302);
and U8591 (N_8591,N_8288,N_8268);
and U8592 (N_8592,N_8395,N_8211);
nand U8593 (N_8593,N_8326,N_8313);
nor U8594 (N_8594,N_8378,N_8214);
nand U8595 (N_8595,N_8248,N_8296);
nor U8596 (N_8596,N_8220,N_8275);
xor U8597 (N_8597,N_8319,N_8321);
nor U8598 (N_8598,N_8399,N_8384);
and U8599 (N_8599,N_8265,N_8383);
nor U8600 (N_8600,N_8458,N_8402);
nor U8601 (N_8601,N_8503,N_8464);
or U8602 (N_8602,N_8528,N_8538);
xor U8603 (N_8603,N_8545,N_8448);
nor U8604 (N_8604,N_8466,N_8469);
nand U8605 (N_8605,N_8584,N_8472);
nor U8606 (N_8606,N_8430,N_8429);
or U8607 (N_8607,N_8487,N_8517);
nand U8608 (N_8608,N_8587,N_8546);
xor U8609 (N_8609,N_8568,N_8533);
xnor U8610 (N_8610,N_8462,N_8415);
nand U8611 (N_8611,N_8510,N_8486);
nor U8612 (N_8612,N_8582,N_8502);
and U8613 (N_8613,N_8467,N_8427);
and U8614 (N_8614,N_8581,N_8432);
xor U8615 (N_8615,N_8509,N_8483);
nand U8616 (N_8616,N_8514,N_8445);
or U8617 (N_8617,N_8406,N_8409);
or U8618 (N_8618,N_8554,N_8426);
or U8619 (N_8619,N_8489,N_8594);
nand U8620 (N_8620,N_8562,N_8526);
and U8621 (N_8621,N_8515,N_8527);
xnor U8622 (N_8622,N_8563,N_8590);
nor U8623 (N_8623,N_8475,N_8410);
nor U8624 (N_8624,N_8488,N_8566);
and U8625 (N_8625,N_8598,N_8529);
nor U8626 (N_8626,N_8485,N_8508);
and U8627 (N_8627,N_8520,N_8542);
or U8628 (N_8628,N_8534,N_8403);
nand U8629 (N_8629,N_8492,N_8419);
xnor U8630 (N_8630,N_8400,N_8440);
nor U8631 (N_8631,N_8457,N_8512);
xor U8632 (N_8632,N_8552,N_8519);
and U8633 (N_8633,N_8453,N_8575);
nor U8634 (N_8634,N_8535,N_8561);
nand U8635 (N_8635,N_8468,N_8567);
or U8636 (N_8636,N_8585,N_8549);
and U8637 (N_8637,N_8441,N_8404);
or U8638 (N_8638,N_8418,N_8421);
or U8639 (N_8639,N_8556,N_8592);
xor U8640 (N_8640,N_8470,N_8442);
nand U8641 (N_8641,N_8536,N_8551);
and U8642 (N_8642,N_8439,N_8417);
and U8643 (N_8643,N_8449,N_8569);
or U8644 (N_8644,N_8484,N_8411);
nand U8645 (N_8645,N_8577,N_8495);
or U8646 (N_8646,N_8401,N_8463);
nor U8647 (N_8647,N_8559,N_8422);
xor U8648 (N_8648,N_8452,N_8565);
and U8649 (N_8649,N_8586,N_8540);
xnor U8650 (N_8650,N_8460,N_8532);
nand U8651 (N_8651,N_8479,N_8576);
nand U8652 (N_8652,N_8412,N_8591);
nand U8653 (N_8653,N_8446,N_8423);
or U8654 (N_8654,N_8588,N_8571);
nor U8655 (N_8655,N_8456,N_8560);
and U8656 (N_8656,N_8522,N_8553);
nand U8657 (N_8657,N_8433,N_8541);
and U8658 (N_8658,N_8498,N_8513);
xor U8659 (N_8659,N_8505,N_8405);
nor U8660 (N_8660,N_8420,N_8416);
and U8661 (N_8661,N_8504,N_8493);
or U8662 (N_8662,N_8497,N_8428);
nor U8663 (N_8663,N_8511,N_8523);
and U8664 (N_8664,N_8524,N_8574);
nor U8665 (N_8665,N_8471,N_8555);
or U8666 (N_8666,N_8506,N_8438);
or U8667 (N_8667,N_8455,N_8572);
and U8668 (N_8668,N_8482,N_8435);
xnor U8669 (N_8669,N_8459,N_8477);
nand U8670 (N_8670,N_8461,N_8499);
and U8671 (N_8671,N_8408,N_8516);
nor U8672 (N_8672,N_8573,N_8521);
and U8673 (N_8673,N_8531,N_8491);
or U8674 (N_8674,N_8437,N_8413);
nor U8675 (N_8675,N_8593,N_8490);
and U8676 (N_8676,N_8507,N_8578);
or U8677 (N_8677,N_8454,N_8580);
nor U8678 (N_8678,N_8599,N_8450);
xor U8679 (N_8679,N_8496,N_8530);
xnor U8680 (N_8680,N_8518,N_8407);
nor U8681 (N_8681,N_8597,N_8525);
xnor U8682 (N_8682,N_8595,N_8596);
or U8683 (N_8683,N_8500,N_8431);
or U8684 (N_8684,N_8539,N_8547);
nand U8685 (N_8685,N_8579,N_8473);
xnor U8686 (N_8686,N_8583,N_8414);
or U8687 (N_8687,N_8474,N_8589);
xor U8688 (N_8688,N_8465,N_8480);
nand U8689 (N_8689,N_8443,N_8501);
xor U8690 (N_8690,N_8436,N_8537);
nand U8691 (N_8691,N_8564,N_8444);
xor U8692 (N_8692,N_8494,N_8557);
nand U8693 (N_8693,N_8434,N_8543);
nor U8694 (N_8694,N_8548,N_8550);
nor U8695 (N_8695,N_8451,N_8425);
nand U8696 (N_8696,N_8544,N_8424);
xnor U8697 (N_8697,N_8476,N_8481);
xnor U8698 (N_8698,N_8558,N_8570);
and U8699 (N_8699,N_8447,N_8478);
xnor U8700 (N_8700,N_8415,N_8531);
xnor U8701 (N_8701,N_8506,N_8493);
and U8702 (N_8702,N_8544,N_8410);
and U8703 (N_8703,N_8596,N_8550);
and U8704 (N_8704,N_8415,N_8409);
nor U8705 (N_8705,N_8456,N_8433);
nand U8706 (N_8706,N_8404,N_8409);
or U8707 (N_8707,N_8491,N_8539);
and U8708 (N_8708,N_8481,N_8561);
xor U8709 (N_8709,N_8472,N_8438);
xor U8710 (N_8710,N_8553,N_8533);
xnor U8711 (N_8711,N_8546,N_8553);
or U8712 (N_8712,N_8567,N_8437);
xnor U8713 (N_8713,N_8521,N_8429);
and U8714 (N_8714,N_8585,N_8577);
nand U8715 (N_8715,N_8548,N_8510);
and U8716 (N_8716,N_8561,N_8573);
or U8717 (N_8717,N_8524,N_8562);
nand U8718 (N_8718,N_8417,N_8401);
xor U8719 (N_8719,N_8490,N_8506);
and U8720 (N_8720,N_8593,N_8481);
and U8721 (N_8721,N_8426,N_8409);
or U8722 (N_8722,N_8593,N_8407);
xor U8723 (N_8723,N_8496,N_8466);
and U8724 (N_8724,N_8565,N_8530);
nand U8725 (N_8725,N_8575,N_8491);
nor U8726 (N_8726,N_8424,N_8515);
nand U8727 (N_8727,N_8574,N_8492);
nand U8728 (N_8728,N_8475,N_8597);
and U8729 (N_8729,N_8530,N_8520);
nor U8730 (N_8730,N_8579,N_8414);
xor U8731 (N_8731,N_8539,N_8434);
and U8732 (N_8732,N_8468,N_8549);
xnor U8733 (N_8733,N_8513,N_8468);
nand U8734 (N_8734,N_8474,N_8464);
and U8735 (N_8735,N_8500,N_8493);
nor U8736 (N_8736,N_8588,N_8469);
or U8737 (N_8737,N_8597,N_8444);
and U8738 (N_8738,N_8401,N_8549);
nor U8739 (N_8739,N_8477,N_8587);
or U8740 (N_8740,N_8590,N_8573);
and U8741 (N_8741,N_8468,N_8404);
or U8742 (N_8742,N_8490,N_8477);
nand U8743 (N_8743,N_8416,N_8545);
or U8744 (N_8744,N_8488,N_8540);
and U8745 (N_8745,N_8482,N_8417);
nor U8746 (N_8746,N_8407,N_8461);
and U8747 (N_8747,N_8491,N_8410);
xnor U8748 (N_8748,N_8587,N_8545);
nor U8749 (N_8749,N_8543,N_8588);
or U8750 (N_8750,N_8479,N_8453);
xor U8751 (N_8751,N_8578,N_8419);
and U8752 (N_8752,N_8523,N_8486);
nor U8753 (N_8753,N_8411,N_8508);
nor U8754 (N_8754,N_8532,N_8441);
nand U8755 (N_8755,N_8564,N_8464);
or U8756 (N_8756,N_8441,N_8425);
xnor U8757 (N_8757,N_8595,N_8556);
nor U8758 (N_8758,N_8429,N_8406);
and U8759 (N_8759,N_8519,N_8543);
nor U8760 (N_8760,N_8506,N_8442);
nor U8761 (N_8761,N_8592,N_8538);
nor U8762 (N_8762,N_8429,N_8450);
xor U8763 (N_8763,N_8423,N_8482);
and U8764 (N_8764,N_8478,N_8520);
nand U8765 (N_8765,N_8581,N_8464);
and U8766 (N_8766,N_8501,N_8436);
xnor U8767 (N_8767,N_8416,N_8494);
nand U8768 (N_8768,N_8459,N_8575);
and U8769 (N_8769,N_8584,N_8561);
nor U8770 (N_8770,N_8536,N_8519);
xor U8771 (N_8771,N_8536,N_8515);
and U8772 (N_8772,N_8421,N_8467);
and U8773 (N_8773,N_8525,N_8599);
nand U8774 (N_8774,N_8407,N_8508);
nand U8775 (N_8775,N_8422,N_8489);
or U8776 (N_8776,N_8514,N_8525);
nor U8777 (N_8777,N_8566,N_8565);
and U8778 (N_8778,N_8548,N_8533);
or U8779 (N_8779,N_8565,N_8436);
and U8780 (N_8780,N_8469,N_8405);
and U8781 (N_8781,N_8477,N_8468);
or U8782 (N_8782,N_8499,N_8588);
nor U8783 (N_8783,N_8469,N_8549);
and U8784 (N_8784,N_8496,N_8525);
nor U8785 (N_8785,N_8572,N_8478);
xnor U8786 (N_8786,N_8524,N_8421);
and U8787 (N_8787,N_8598,N_8450);
xnor U8788 (N_8788,N_8534,N_8438);
xnor U8789 (N_8789,N_8557,N_8480);
xnor U8790 (N_8790,N_8556,N_8489);
or U8791 (N_8791,N_8574,N_8582);
nand U8792 (N_8792,N_8516,N_8456);
or U8793 (N_8793,N_8405,N_8570);
xnor U8794 (N_8794,N_8472,N_8452);
or U8795 (N_8795,N_8549,N_8577);
or U8796 (N_8796,N_8529,N_8517);
nor U8797 (N_8797,N_8427,N_8414);
and U8798 (N_8798,N_8413,N_8431);
and U8799 (N_8799,N_8454,N_8520);
xor U8800 (N_8800,N_8645,N_8767);
xor U8801 (N_8801,N_8606,N_8637);
and U8802 (N_8802,N_8786,N_8757);
and U8803 (N_8803,N_8613,N_8628);
nor U8804 (N_8804,N_8698,N_8760);
xor U8805 (N_8805,N_8795,N_8788);
nor U8806 (N_8806,N_8758,N_8662);
nor U8807 (N_8807,N_8658,N_8718);
or U8808 (N_8808,N_8629,N_8648);
or U8809 (N_8809,N_8784,N_8665);
xnor U8810 (N_8810,N_8787,N_8731);
and U8811 (N_8811,N_8791,N_8689);
and U8812 (N_8812,N_8745,N_8635);
nand U8813 (N_8813,N_8724,N_8756);
and U8814 (N_8814,N_8730,N_8746);
xor U8815 (N_8815,N_8609,N_8602);
nand U8816 (N_8816,N_8691,N_8650);
or U8817 (N_8817,N_8616,N_8687);
or U8818 (N_8818,N_8772,N_8793);
nand U8819 (N_8819,N_8721,N_8727);
nand U8820 (N_8820,N_8726,N_8610);
and U8821 (N_8821,N_8693,N_8782);
xor U8822 (N_8822,N_8776,N_8652);
xnor U8823 (N_8823,N_8608,N_8747);
xor U8824 (N_8824,N_8759,N_8622);
nand U8825 (N_8825,N_8711,N_8749);
or U8826 (N_8826,N_8625,N_8636);
nand U8827 (N_8827,N_8642,N_8684);
nand U8828 (N_8828,N_8792,N_8669);
nand U8829 (N_8829,N_8785,N_8603);
nand U8830 (N_8830,N_8748,N_8742);
xor U8831 (N_8831,N_8601,N_8769);
nor U8832 (N_8832,N_8663,N_8670);
nor U8833 (N_8833,N_8640,N_8704);
nand U8834 (N_8834,N_8619,N_8755);
nand U8835 (N_8835,N_8764,N_8634);
and U8836 (N_8836,N_8761,N_8725);
xnor U8837 (N_8837,N_8656,N_8617);
xnor U8838 (N_8838,N_8678,N_8728);
and U8839 (N_8839,N_8799,N_8743);
xnor U8840 (N_8840,N_8703,N_8719);
xor U8841 (N_8841,N_8796,N_8778);
xnor U8842 (N_8842,N_8690,N_8614);
and U8843 (N_8843,N_8646,N_8686);
xor U8844 (N_8844,N_8692,N_8660);
nand U8845 (N_8845,N_8683,N_8671);
nand U8846 (N_8846,N_8604,N_8774);
xnor U8847 (N_8847,N_8685,N_8702);
xor U8848 (N_8848,N_8667,N_8618);
and U8849 (N_8849,N_8639,N_8713);
and U8850 (N_8850,N_8661,N_8717);
nand U8851 (N_8851,N_8754,N_8666);
or U8852 (N_8852,N_8798,N_8664);
xor U8853 (N_8853,N_8680,N_8688);
and U8854 (N_8854,N_8779,N_8773);
nor U8855 (N_8855,N_8643,N_8737);
and U8856 (N_8856,N_8600,N_8710);
and U8857 (N_8857,N_8729,N_8674);
and U8858 (N_8858,N_8783,N_8715);
xor U8859 (N_8859,N_8720,N_8716);
or U8860 (N_8860,N_8709,N_8615);
nor U8861 (N_8861,N_8797,N_8722);
xnor U8862 (N_8862,N_8647,N_8620);
nor U8863 (N_8863,N_8705,N_8752);
or U8864 (N_8864,N_8697,N_8775);
or U8865 (N_8865,N_8699,N_8630);
nor U8866 (N_8866,N_8633,N_8790);
xnor U8867 (N_8867,N_8627,N_8765);
xor U8868 (N_8868,N_8657,N_8741);
xor U8869 (N_8869,N_8644,N_8682);
nor U8870 (N_8870,N_8654,N_8621);
xnor U8871 (N_8871,N_8623,N_8734);
nor U8872 (N_8872,N_8675,N_8751);
xor U8873 (N_8873,N_8712,N_8771);
nor U8874 (N_8874,N_8612,N_8739);
nor U8875 (N_8875,N_8641,N_8676);
xor U8876 (N_8876,N_8651,N_8794);
or U8877 (N_8877,N_8673,N_8780);
xor U8878 (N_8878,N_8753,N_8694);
and U8879 (N_8879,N_8624,N_8738);
or U8880 (N_8880,N_8649,N_8732);
or U8881 (N_8881,N_8777,N_8632);
or U8882 (N_8882,N_8679,N_8681);
or U8883 (N_8883,N_8750,N_8626);
nand U8884 (N_8884,N_8605,N_8607);
xor U8885 (N_8885,N_8735,N_8707);
nand U8886 (N_8886,N_8701,N_8763);
xnor U8887 (N_8887,N_8638,N_8762);
xnor U8888 (N_8888,N_8696,N_8770);
nand U8889 (N_8889,N_8695,N_8744);
and U8890 (N_8890,N_8706,N_8659);
and U8891 (N_8891,N_8700,N_8611);
and U8892 (N_8892,N_8733,N_8714);
nor U8893 (N_8893,N_8740,N_8723);
or U8894 (N_8894,N_8766,N_8736);
nand U8895 (N_8895,N_8768,N_8789);
or U8896 (N_8896,N_8677,N_8655);
xor U8897 (N_8897,N_8653,N_8668);
nand U8898 (N_8898,N_8672,N_8708);
xor U8899 (N_8899,N_8631,N_8781);
nor U8900 (N_8900,N_8615,N_8618);
nor U8901 (N_8901,N_8773,N_8654);
xnor U8902 (N_8902,N_8671,N_8657);
or U8903 (N_8903,N_8657,N_8612);
xnor U8904 (N_8904,N_8742,N_8774);
or U8905 (N_8905,N_8782,N_8731);
nor U8906 (N_8906,N_8686,N_8789);
xor U8907 (N_8907,N_8748,N_8733);
or U8908 (N_8908,N_8755,N_8691);
or U8909 (N_8909,N_8781,N_8686);
or U8910 (N_8910,N_8706,N_8773);
xor U8911 (N_8911,N_8669,N_8619);
or U8912 (N_8912,N_8713,N_8759);
and U8913 (N_8913,N_8657,N_8799);
xnor U8914 (N_8914,N_8760,N_8649);
nand U8915 (N_8915,N_8678,N_8772);
or U8916 (N_8916,N_8612,N_8798);
nand U8917 (N_8917,N_8659,N_8783);
and U8918 (N_8918,N_8679,N_8638);
and U8919 (N_8919,N_8780,N_8645);
nand U8920 (N_8920,N_8625,N_8710);
nor U8921 (N_8921,N_8776,N_8785);
or U8922 (N_8922,N_8605,N_8702);
nand U8923 (N_8923,N_8770,N_8666);
xnor U8924 (N_8924,N_8757,N_8701);
or U8925 (N_8925,N_8655,N_8693);
or U8926 (N_8926,N_8741,N_8647);
xnor U8927 (N_8927,N_8612,N_8655);
xnor U8928 (N_8928,N_8796,N_8723);
nand U8929 (N_8929,N_8784,N_8650);
nand U8930 (N_8930,N_8730,N_8602);
or U8931 (N_8931,N_8696,N_8727);
nand U8932 (N_8932,N_8749,N_8601);
nor U8933 (N_8933,N_8624,N_8614);
and U8934 (N_8934,N_8664,N_8678);
and U8935 (N_8935,N_8658,N_8728);
or U8936 (N_8936,N_8701,N_8654);
nor U8937 (N_8937,N_8698,N_8684);
nor U8938 (N_8938,N_8778,N_8791);
nand U8939 (N_8939,N_8771,N_8629);
and U8940 (N_8940,N_8710,N_8761);
and U8941 (N_8941,N_8669,N_8729);
nor U8942 (N_8942,N_8786,N_8707);
or U8943 (N_8943,N_8618,N_8651);
nand U8944 (N_8944,N_8765,N_8750);
nor U8945 (N_8945,N_8748,N_8775);
nor U8946 (N_8946,N_8748,N_8702);
or U8947 (N_8947,N_8642,N_8746);
nor U8948 (N_8948,N_8720,N_8767);
nor U8949 (N_8949,N_8709,N_8725);
xnor U8950 (N_8950,N_8656,N_8689);
xor U8951 (N_8951,N_8712,N_8692);
or U8952 (N_8952,N_8794,N_8633);
and U8953 (N_8953,N_8658,N_8782);
and U8954 (N_8954,N_8650,N_8775);
xor U8955 (N_8955,N_8720,N_8748);
and U8956 (N_8956,N_8691,N_8664);
and U8957 (N_8957,N_8755,N_8696);
nand U8958 (N_8958,N_8675,N_8693);
nor U8959 (N_8959,N_8653,N_8781);
xnor U8960 (N_8960,N_8747,N_8666);
nor U8961 (N_8961,N_8691,N_8776);
nand U8962 (N_8962,N_8681,N_8767);
and U8963 (N_8963,N_8656,N_8622);
nor U8964 (N_8964,N_8755,N_8673);
xnor U8965 (N_8965,N_8695,N_8781);
xor U8966 (N_8966,N_8684,N_8657);
and U8967 (N_8967,N_8790,N_8632);
nand U8968 (N_8968,N_8749,N_8761);
or U8969 (N_8969,N_8757,N_8660);
nand U8970 (N_8970,N_8769,N_8687);
or U8971 (N_8971,N_8752,N_8720);
xor U8972 (N_8972,N_8794,N_8632);
xor U8973 (N_8973,N_8765,N_8649);
and U8974 (N_8974,N_8717,N_8697);
or U8975 (N_8975,N_8765,N_8656);
or U8976 (N_8976,N_8775,N_8624);
nor U8977 (N_8977,N_8723,N_8666);
nand U8978 (N_8978,N_8654,N_8611);
or U8979 (N_8979,N_8726,N_8649);
xnor U8980 (N_8980,N_8621,N_8746);
and U8981 (N_8981,N_8642,N_8682);
and U8982 (N_8982,N_8756,N_8687);
nand U8983 (N_8983,N_8606,N_8779);
and U8984 (N_8984,N_8787,N_8793);
and U8985 (N_8985,N_8725,N_8608);
nor U8986 (N_8986,N_8758,N_8611);
or U8987 (N_8987,N_8756,N_8680);
and U8988 (N_8988,N_8657,N_8610);
nor U8989 (N_8989,N_8665,N_8601);
and U8990 (N_8990,N_8769,N_8668);
nand U8991 (N_8991,N_8664,N_8698);
or U8992 (N_8992,N_8771,N_8730);
xor U8993 (N_8993,N_8724,N_8637);
nand U8994 (N_8994,N_8641,N_8704);
nand U8995 (N_8995,N_8683,N_8688);
and U8996 (N_8996,N_8755,N_8626);
nor U8997 (N_8997,N_8763,N_8765);
or U8998 (N_8998,N_8730,N_8705);
nand U8999 (N_8999,N_8611,N_8625);
xnor U9000 (N_9000,N_8888,N_8913);
nand U9001 (N_9001,N_8801,N_8925);
or U9002 (N_9002,N_8997,N_8963);
and U9003 (N_9003,N_8854,N_8969);
nor U9004 (N_9004,N_8885,N_8852);
xnor U9005 (N_9005,N_8965,N_8961);
and U9006 (N_9006,N_8826,N_8919);
nand U9007 (N_9007,N_8865,N_8896);
and U9008 (N_9008,N_8816,N_8900);
nand U9009 (N_9009,N_8908,N_8891);
nor U9010 (N_9010,N_8892,N_8993);
or U9011 (N_9011,N_8860,N_8846);
nand U9012 (N_9012,N_8867,N_8808);
nor U9013 (N_9013,N_8861,N_8809);
xor U9014 (N_9014,N_8928,N_8890);
or U9015 (N_9015,N_8986,N_8933);
and U9016 (N_9016,N_8876,N_8817);
and U9017 (N_9017,N_8921,N_8847);
and U9018 (N_9018,N_8995,N_8974);
nand U9019 (N_9019,N_8818,N_8953);
xnor U9020 (N_9020,N_8806,N_8882);
nand U9021 (N_9021,N_8981,N_8853);
and U9022 (N_9022,N_8996,N_8980);
xnor U9023 (N_9023,N_8887,N_8884);
nand U9024 (N_9024,N_8813,N_8845);
xnor U9025 (N_9025,N_8917,N_8841);
or U9026 (N_9026,N_8889,N_8807);
nor U9027 (N_9027,N_8849,N_8869);
xnor U9028 (N_9028,N_8901,N_8832);
nand U9029 (N_9029,N_8934,N_8920);
nand U9030 (N_9030,N_8989,N_8870);
and U9031 (N_9031,N_8827,N_8964);
xnor U9032 (N_9032,N_8883,N_8930);
xor U9033 (N_9033,N_8825,N_8911);
nor U9034 (N_9034,N_8830,N_8987);
nor U9035 (N_9035,N_8983,N_8822);
xor U9036 (N_9036,N_8951,N_8923);
xnor U9037 (N_9037,N_8863,N_8984);
nand U9038 (N_9038,N_8897,N_8916);
xor U9039 (N_9039,N_8828,N_8834);
and U9040 (N_9040,N_8850,N_8856);
xnor U9041 (N_9041,N_8910,N_8970);
or U9042 (N_9042,N_8945,N_8950);
and U9043 (N_9043,N_8851,N_8968);
nor U9044 (N_9044,N_8804,N_8924);
or U9045 (N_9045,N_8873,N_8904);
xnor U9046 (N_9046,N_8999,N_8994);
xor U9047 (N_9047,N_8927,N_8814);
and U9048 (N_9048,N_8812,N_8922);
xor U9049 (N_9049,N_8948,N_8903);
or U9050 (N_9050,N_8898,N_8819);
or U9051 (N_9051,N_8975,N_8952);
and U9052 (N_9052,N_8811,N_8829);
nand U9053 (N_9053,N_8862,N_8905);
nor U9054 (N_9054,N_8979,N_8843);
and U9055 (N_9055,N_8886,N_8929);
or U9056 (N_9056,N_8824,N_8820);
or U9057 (N_9057,N_8875,N_8982);
nor U9058 (N_9058,N_8977,N_8914);
and U9059 (N_9059,N_8857,N_8958);
or U9060 (N_9060,N_8985,N_8895);
xnor U9061 (N_9061,N_8973,N_8837);
nand U9062 (N_9062,N_8967,N_8972);
or U9063 (N_9063,N_8855,N_8976);
xor U9064 (N_9064,N_8918,N_8840);
nor U9065 (N_9065,N_8858,N_8844);
nor U9066 (N_9066,N_8879,N_8915);
nor U9067 (N_9067,N_8956,N_8954);
nand U9068 (N_9068,N_8866,N_8836);
xor U9069 (N_9069,N_8815,N_8874);
or U9070 (N_9070,N_8909,N_8971);
and U9071 (N_9071,N_8937,N_8939);
or U9072 (N_9072,N_8962,N_8803);
or U9073 (N_9073,N_8931,N_8823);
nor U9074 (N_9074,N_8881,N_8912);
xor U9075 (N_9075,N_8998,N_8944);
or U9076 (N_9076,N_8926,N_8880);
nor U9077 (N_9077,N_8894,N_8848);
nor U9078 (N_9078,N_8988,N_8864);
nand U9079 (N_9079,N_8899,N_8842);
or U9080 (N_9080,N_8932,N_8838);
or U9081 (N_9081,N_8941,N_8991);
and U9082 (N_9082,N_8802,N_8871);
nor U9083 (N_9083,N_8906,N_8805);
nand U9084 (N_9084,N_8957,N_8960);
xor U9085 (N_9085,N_8966,N_8940);
or U9086 (N_9086,N_8833,N_8949);
or U9087 (N_9087,N_8835,N_8868);
and U9088 (N_9088,N_8821,N_8810);
xor U9089 (N_9089,N_8893,N_8946);
nor U9090 (N_9090,N_8992,N_8955);
nand U9091 (N_9091,N_8907,N_8859);
nor U9092 (N_9092,N_8839,N_8877);
nor U9093 (N_9093,N_8935,N_8902);
nor U9094 (N_9094,N_8990,N_8878);
and U9095 (N_9095,N_8943,N_8947);
nor U9096 (N_9096,N_8831,N_8959);
nor U9097 (N_9097,N_8800,N_8938);
or U9098 (N_9098,N_8936,N_8942);
and U9099 (N_9099,N_8978,N_8872);
nor U9100 (N_9100,N_8884,N_8986);
xor U9101 (N_9101,N_8901,N_8820);
and U9102 (N_9102,N_8908,N_8893);
xor U9103 (N_9103,N_8972,N_8989);
xor U9104 (N_9104,N_8948,N_8964);
xor U9105 (N_9105,N_8855,N_8806);
nand U9106 (N_9106,N_8828,N_8921);
or U9107 (N_9107,N_8827,N_8841);
and U9108 (N_9108,N_8856,N_8981);
nor U9109 (N_9109,N_8818,N_8898);
nand U9110 (N_9110,N_8951,N_8905);
xnor U9111 (N_9111,N_8909,N_8876);
xnor U9112 (N_9112,N_8814,N_8995);
or U9113 (N_9113,N_8800,N_8897);
nor U9114 (N_9114,N_8877,N_8809);
nand U9115 (N_9115,N_8976,N_8891);
xor U9116 (N_9116,N_8933,N_8947);
or U9117 (N_9117,N_8887,N_8982);
nor U9118 (N_9118,N_8830,N_8940);
nor U9119 (N_9119,N_8802,N_8801);
nand U9120 (N_9120,N_8983,N_8920);
xor U9121 (N_9121,N_8825,N_8831);
nor U9122 (N_9122,N_8893,N_8802);
nor U9123 (N_9123,N_8886,N_8956);
xnor U9124 (N_9124,N_8974,N_8973);
nor U9125 (N_9125,N_8820,N_8941);
nand U9126 (N_9126,N_8928,N_8862);
xor U9127 (N_9127,N_8817,N_8900);
and U9128 (N_9128,N_8893,N_8870);
and U9129 (N_9129,N_8914,N_8958);
or U9130 (N_9130,N_8988,N_8838);
and U9131 (N_9131,N_8927,N_8863);
or U9132 (N_9132,N_8826,N_8973);
nor U9133 (N_9133,N_8865,N_8937);
or U9134 (N_9134,N_8867,N_8989);
or U9135 (N_9135,N_8970,N_8987);
xnor U9136 (N_9136,N_8900,N_8978);
xor U9137 (N_9137,N_8859,N_8872);
and U9138 (N_9138,N_8954,N_8964);
xnor U9139 (N_9139,N_8820,N_8936);
nand U9140 (N_9140,N_8825,N_8998);
or U9141 (N_9141,N_8917,N_8838);
or U9142 (N_9142,N_8984,N_8857);
or U9143 (N_9143,N_8844,N_8902);
or U9144 (N_9144,N_8889,N_8982);
nand U9145 (N_9145,N_8913,N_8898);
or U9146 (N_9146,N_8897,N_8960);
xnor U9147 (N_9147,N_8822,N_8845);
nand U9148 (N_9148,N_8805,N_8803);
and U9149 (N_9149,N_8872,N_8925);
nor U9150 (N_9150,N_8995,N_8850);
xnor U9151 (N_9151,N_8873,N_8805);
nor U9152 (N_9152,N_8853,N_8918);
and U9153 (N_9153,N_8815,N_8816);
nor U9154 (N_9154,N_8986,N_8889);
xnor U9155 (N_9155,N_8884,N_8905);
nand U9156 (N_9156,N_8854,N_8914);
nor U9157 (N_9157,N_8870,N_8841);
or U9158 (N_9158,N_8809,N_8889);
xor U9159 (N_9159,N_8809,N_8890);
nor U9160 (N_9160,N_8937,N_8804);
nor U9161 (N_9161,N_8959,N_8919);
nor U9162 (N_9162,N_8993,N_8814);
xnor U9163 (N_9163,N_8807,N_8998);
and U9164 (N_9164,N_8882,N_8953);
and U9165 (N_9165,N_8855,N_8899);
nand U9166 (N_9166,N_8844,N_8815);
or U9167 (N_9167,N_8839,N_8957);
xnor U9168 (N_9168,N_8856,N_8984);
or U9169 (N_9169,N_8803,N_8923);
xnor U9170 (N_9170,N_8827,N_8940);
or U9171 (N_9171,N_8991,N_8997);
and U9172 (N_9172,N_8921,N_8949);
and U9173 (N_9173,N_8879,N_8896);
xor U9174 (N_9174,N_8956,N_8981);
xnor U9175 (N_9175,N_8978,N_8869);
xor U9176 (N_9176,N_8832,N_8828);
or U9177 (N_9177,N_8870,N_8938);
or U9178 (N_9178,N_8819,N_8956);
xor U9179 (N_9179,N_8925,N_8990);
xnor U9180 (N_9180,N_8975,N_8819);
and U9181 (N_9181,N_8856,N_8827);
nand U9182 (N_9182,N_8814,N_8802);
xor U9183 (N_9183,N_8874,N_8953);
xor U9184 (N_9184,N_8821,N_8902);
xnor U9185 (N_9185,N_8810,N_8891);
and U9186 (N_9186,N_8964,N_8847);
xnor U9187 (N_9187,N_8888,N_8863);
or U9188 (N_9188,N_8985,N_8915);
xnor U9189 (N_9189,N_8857,N_8872);
nand U9190 (N_9190,N_8976,N_8926);
xnor U9191 (N_9191,N_8825,N_8816);
xor U9192 (N_9192,N_8948,N_8838);
nor U9193 (N_9193,N_8927,N_8895);
or U9194 (N_9194,N_8971,N_8994);
nor U9195 (N_9195,N_8927,N_8867);
nand U9196 (N_9196,N_8951,N_8985);
nor U9197 (N_9197,N_8945,N_8896);
nor U9198 (N_9198,N_8920,N_8847);
nor U9199 (N_9199,N_8853,N_8838);
nand U9200 (N_9200,N_9159,N_9142);
and U9201 (N_9201,N_9173,N_9128);
xnor U9202 (N_9202,N_9119,N_9080);
xnor U9203 (N_9203,N_9070,N_9189);
or U9204 (N_9204,N_9065,N_9112);
and U9205 (N_9205,N_9054,N_9038);
nand U9206 (N_9206,N_9008,N_9176);
or U9207 (N_9207,N_9178,N_9023);
nor U9208 (N_9208,N_9103,N_9073);
and U9209 (N_9209,N_9022,N_9061);
and U9210 (N_9210,N_9107,N_9168);
or U9211 (N_9211,N_9147,N_9110);
xor U9212 (N_9212,N_9018,N_9174);
xor U9213 (N_9213,N_9184,N_9089);
or U9214 (N_9214,N_9124,N_9043);
nand U9215 (N_9215,N_9028,N_9033);
xnor U9216 (N_9216,N_9118,N_9076);
or U9217 (N_9217,N_9031,N_9049);
xor U9218 (N_9218,N_9003,N_9177);
nor U9219 (N_9219,N_9036,N_9091);
and U9220 (N_9220,N_9152,N_9059);
xor U9221 (N_9221,N_9143,N_9111);
nand U9222 (N_9222,N_9006,N_9130);
and U9223 (N_9223,N_9074,N_9007);
nor U9224 (N_9224,N_9196,N_9083);
or U9225 (N_9225,N_9120,N_9027);
nand U9226 (N_9226,N_9109,N_9092);
nor U9227 (N_9227,N_9063,N_9187);
nand U9228 (N_9228,N_9005,N_9077);
nand U9229 (N_9229,N_9134,N_9058);
nand U9230 (N_9230,N_9141,N_9150);
nor U9231 (N_9231,N_9047,N_9072);
nand U9232 (N_9232,N_9144,N_9052);
nor U9233 (N_9233,N_9132,N_9001);
and U9234 (N_9234,N_9166,N_9138);
and U9235 (N_9235,N_9048,N_9123);
and U9236 (N_9236,N_9115,N_9160);
nor U9237 (N_9237,N_9067,N_9095);
and U9238 (N_9238,N_9026,N_9066);
nand U9239 (N_9239,N_9002,N_9040);
or U9240 (N_9240,N_9094,N_9163);
nor U9241 (N_9241,N_9183,N_9011);
nand U9242 (N_9242,N_9030,N_9009);
nand U9243 (N_9243,N_9169,N_9190);
nand U9244 (N_9244,N_9034,N_9131);
xnor U9245 (N_9245,N_9105,N_9055);
nor U9246 (N_9246,N_9153,N_9188);
and U9247 (N_9247,N_9068,N_9162);
and U9248 (N_9248,N_9167,N_9180);
xor U9249 (N_9249,N_9161,N_9149);
nand U9250 (N_9250,N_9041,N_9129);
and U9251 (N_9251,N_9020,N_9039);
xor U9252 (N_9252,N_9079,N_9133);
xnor U9253 (N_9253,N_9137,N_9093);
nor U9254 (N_9254,N_9148,N_9019);
nor U9255 (N_9255,N_9081,N_9108);
nor U9256 (N_9256,N_9125,N_9098);
xnor U9257 (N_9257,N_9114,N_9010);
or U9258 (N_9258,N_9170,N_9017);
nand U9259 (N_9259,N_9145,N_9172);
nor U9260 (N_9260,N_9165,N_9175);
nor U9261 (N_9261,N_9127,N_9014);
xnor U9262 (N_9262,N_9194,N_9000);
nand U9263 (N_9263,N_9082,N_9084);
nand U9264 (N_9264,N_9154,N_9064);
xnor U9265 (N_9265,N_9102,N_9053);
and U9266 (N_9266,N_9140,N_9100);
or U9267 (N_9267,N_9191,N_9056);
nor U9268 (N_9268,N_9035,N_9139);
nor U9269 (N_9269,N_9051,N_9069);
nor U9270 (N_9270,N_9121,N_9078);
xnor U9271 (N_9271,N_9117,N_9136);
nor U9272 (N_9272,N_9057,N_9164);
nor U9273 (N_9273,N_9186,N_9016);
xor U9274 (N_9274,N_9013,N_9193);
and U9275 (N_9275,N_9060,N_9096);
nor U9276 (N_9276,N_9044,N_9012);
nand U9277 (N_9277,N_9029,N_9195);
and U9278 (N_9278,N_9126,N_9199);
xnor U9279 (N_9279,N_9197,N_9046);
nor U9280 (N_9280,N_9045,N_9024);
or U9281 (N_9281,N_9071,N_9085);
nor U9282 (N_9282,N_9104,N_9015);
or U9283 (N_9283,N_9158,N_9090);
and U9284 (N_9284,N_9025,N_9086);
or U9285 (N_9285,N_9099,N_9156);
xnor U9286 (N_9286,N_9062,N_9181);
nor U9287 (N_9287,N_9004,N_9042);
or U9288 (N_9288,N_9146,N_9135);
xor U9289 (N_9289,N_9151,N_9050);
and U9290 (N_9290,N_9113,N_9155);
nand U9291 (N_9291,N_9088,N_9171);
and U9292 (N_9292,N_9032,N_9106);
and U9293 (N_9293,N_9087,N_9037);
xnor U9294 (N_9294,N_9182,N_9075);
xnor U9295 (N_9295,N_9198,N_9021);
and U9296 (N_9296,N_9179,N_9122);
nand U9297 (N_9297,N_9116,N_9157);
or U9298 (N_9298,N_9192,N_9097);
nand U9299 (N_9299,N_9101,N_9185);
and U9300 (N_9300,N_9046,N_9144);
or U9301 (N_9301,N_9173,N_9148);
or U9302 (N_9302,N_9140,N_9020);
xnor U9303 (N_9303,N_9197,N_9151);
and U9304 (N_9304,N_9077,N_9097);
or U9305 (N_9305,N_9045,N_9064);
and U9306 (N_9306,N_9068,N_9080);
xnor U9307 (N_9307,N_9034,N_9190);
xnor U9308 (N_9308,N_9132,N_9048);
or U9309 (N_9309,N_9094,N_9158);
nor U9310 (N_9310,N_9105,N_9100);
or U9311 (N_9311,N_9057,N_9014);
and U9312 (N_9312,N_9013,N_9094);
nand U9313 (N_9313,N_9091,N_9097);
nor U9314 (N_9314,N_9098,N_9151);
or U9315 (N_9315,N_9129,N_9046);
or U9316 (N_9316,N_9124,N_9002);
or U9317 (N_9317,N_9192,N_9123);
xnor U9318 (N_9318,N_9057,N_9172);
or U9319 (N_9319,N_9078,N_9153);
xor U9320 (N_9320,N_9102,N_9076);
nor U9321 (N_9321,N_9082,N_9043);
nand U9322 (N_9322,N_9130,N_9067);
xnor U9323 (N_9323,N_9107,N_9132);
nand U9324 (N_9324,N_9047,N_9053);
and U9325 (N_9325,N_9039,N_9048);
nor U9326 (N_9326,N_9144,N_9030);
and U9327 (N_9327,N_9057,N_9145);
nor U9328 (N_9328,N_9139,N_9008);
or U9329 (N_9329,N_9028,N_9118);
or U9330 (N_9330,N_9162,N_9074);
and U9331 (N_9331,N_9049,N_9023);
nand U9332 (N_9332,N_9101,N_9007);
and U9333 (N_9333,N_9051,N_9197);
nand U9334 (N_9334,N_9044,N_9127);
nand U9335 (N_9335,N_9010,N_9099);
nor U9336 (N_9336,N_9148,N_9125);
xor U9337 (N_9337,N_9031,N_9132);
and U9338 (N_9338,N_9195,N_9130);
xnor U9339 (N_9339,N_9197,N_9007);
xor U9340 (N_9340,N_9194,N_9105);
and U9341 (N_9341,N_9198,N_9003);
and U9342 (N_9342,N_9093,N_9040);
or U9343 (N_9343,N_9024,N_9035);
and U9344 (N_9344,N_9121,N_9171);
or U9345 (N_9345,N_9165,N_9004);
nand U9346 (N_9346,N_9198,N_9112);
xor U9347 (N_9347,N_9092,N_9065);
nand U9348 (N_9348,N_9151,N_9008);
or U9349 (N_9349,N_9065,N_9023);
nor U9350 (N_9350,N_9025,N_9125);
nand U9351 (N_9351,N_9060,N_9195);
xnor U9352 (N_9352,N_9073,N_9014);
nand U9353 (N_9353,N_9149,N_9018);
xnor U9354 (N_9354,N_9167,N_9063);
and U9355 (N_9355,N_9050,N_9053);
xnor U9356 (N_9356,N_9070,N_9023);
xor U9357 (N_9357,N_9090,N_9156);
and U9358 (N_9358,N_9088,N_9065);
xnor U9359 (N_9359,N_9060,N_9156);
or U9360 (N_9360,N_9129,N_9169);
or U9361 (N_9361,N_9177,N_9031);
nand U9362 (N_9362,N_9178,N_9125);
or U9363 (N_9363,N_9168,N_9128);
xor U9364 (N_9364,N_9121,N_9007);
or U9365 (N_9365,N_9006,N_9047);
nor U9366 (N_9366,N_9070,N_9069);
nor U9367 (N_9367,N_9014,N_9015);
or U9368 (N_9368,N_9120,N_9051);
nor U9369 (N_9369,N_9035,N_9192);
nand U9370 (N_9370,N_9074,N_9172);
or U9371 (N_9371,N_9057,N_9042);
and U9372 (N_9372,N_9118,N_9105);
or U9373 (N_9373,N_9188,N_9039);
and U9374 (N_9374,N_9000,N_9154);
and U9375 (N_9375,N_9060,N_9130);
and U9376 (N_9376,N_9040,N_9175);
nor U9377 (N_9377,N_9182,N_9098);
xnor U9378 (N_9378,N_9091,N_9191);
nand U9379 (N_9379,N_9174,N_9027);
or U9380 (N_9380,N_9127,N_9005);
xnor U9381 (N_9381,N_9044,N_9195);
xor U9382 (N_9382,N_9042,N_9196);
nor U9383 (N_9383,N_9075,N_9029);
nand U9384 (N_9384,N_9005,N_9109);
and U9385 (N_9385,N_9151,N_9187);
nor U9386 (N_9386,N_9017,N_9193);
xnor U9387 (N_9387,N_9152,N_9114);
or U9388 (N_9388,N_9189,N_9135);
xor U9389 (N_9389,N_9061,N_9057);
nand U9390 (N_9390,N_9154,N_9146);
nand U9391 (N_9391,N_9014,N_9124);
nor U9392 (N_9392,N_9088,N_9143);
and U9393 (N_9393,N_9144,N_9127);
nand U9394 (N_9394,N_9169,N_9069);
xor U9395 (N_9395,N_9132,N_9195);
xor U9396 (N_9396,N_9188,N_9175);
nor U9397 (N_9397,N_9154,N_9028);
and U9398 (N_9398,N_9092,N_9195);
and U9399 (N_9399,N_9027,N_9147);
and U9400 (N_9400,N_9327,N_9238);
nor U9401 (N_9401,N_9208,N_9353);
and U9402 (N_9402,N_9319,N_9224);
nor U9403 (N_9403,N_9226,N_9249);
nor U9404 (N_9404,N_9252,N_9376);
nand U9405 (N_9405,N_9324,N_9269);
or U9406 (N_9406,N_9370,N_9299);
and U9407 (N_9407,N_9356,N_9213);
or U9408 (N_9408,N_9383,N_9337);
and U9409 (N_9409,N_9245,N_9315);
or U9410 (N_9410,N_9289,N_9292);
nand U9411 (N_9411,N_9264,N_9281);
or U9412 (N_9412,N_9367,N_9207);
and U9413 (N_9413,N_9274,N_9293);
or U9414 (N_9414,N_9246,N_9374);
nor U9415 (N_9415,N_9270,N_9278);
nand U9416 (N_9416,N_9240,N_9254);
nand U9417 (N_9417,N_9256,N_9312);
nor U9418 (N_9418,N_9314,N_9237);
and U9419 (N_9419,N_9379,N_9355);
or U9420 (N_9420,N_9211,N_9334);
xnor U9421 (N_9421,N_9345,N_9307);
and U9422 (N_9422,N_9287,N_9310);
or U9423 (N_9423,N_9272,N_9375);
and U9424 (N_9424,N_9248,N_9318);
nor U9425 (N_9425,N_9372,N_9255);
or U9426 (N_9426,N_9222,N_9275);
or U9427 (N_9427,N_9390,N_9369);
nor U9428 (N_9428,N_9219,N_9215);
nor U9429 (N_9429,N_9386,N_9244);
xnor U9430 (N_9430,N_9282,N_9262);
nor U9431 (N_9431,N_9392,N_9331);
xor U9432 (N_9432,N_9216,N_9266);
and U9433 (N_9433,N_9247,N_9394);
and U9434 (N_9434,N_9399,N_9251);
or U9435 (N_9435,N_9243,N_9389);
xnor U9436 (N_9436,N_9218,N_9357);
and U9437 (N_9437,N_9286,N_9348);
or U9438 (N_9438,N_9214,N_9384);
xor U9439 (N_9439,N_9298,N_9295);
and U9440 (N_9440,N_9230,N_9202);
or U9441 (N_9441,N_9349,N_9229);
nand U9442 (N_9442,N_9223,N_9225);
or U9443 (N_9443,N_9209,N_9291);
nor U9444 (N_9444,N_9380,N_9210);
or U9445 (N_9445,N_9311,N_9313);
or U9446 (N_9446,N_9276,N_9288);
and U9447 (N_9447,N_9341,N_9263);
xnor U9448 (N_9448,N_9290,N_9306);
or U9449 (N_9449,N_9339,N_9396);
nor U9450 (N_9450,N_9338,N_9340);
or U9451 (N_9451,N_9297,N_9371);
nand U9452 (N_9452,N_9351,N_9265);
or U9453 (N_9453,N_9258,N_9301);
xnor U9454 (N_9454,N_9232,N_9316);
or U9455 (N_9455,N_9382,N_9362);
and U9456 (N_9456,N_9304,N_9280);
nor U9457 (N_9457,N_9271,N_9317);
xor U9458 (N_9458,N_9234,N_9268);
nand U9459 (N_9459,N_9359,N_9373);
and U9460 (N_9460,N_9328,N_9397);
and U9461 (N_9461,N_9201,N_9279);
or U9462 (N_9462,N_9242,N_9308);
and U9463 (N_9463,N_9342,N_9361);
xnor U9464 (N_9464,N_9366,N_9320);
xnor U9465 (N_9465,N_9294,N_9335);
xor U9466 (N_9466,N_9388,N_9360);
or U9467 (N_9467,N_9231,N_9323);
and U9468 (N_9468,N_9393,N_9391);
nand U9469 (N_9469,N_9239,N_9220);
xor U9470 (N_9470,N_9343,N_9259);
nor U9471 (N_9471,N_9277,N_9363);
and U9472 (N_9472,N_9336,N_9253);
or U9473 (N_9473,N_9296,N_9364);
nor U9474 (N_9474,N_9395,N_9200);
nand U9475 (N_9475,N_9233,N_9354);
nand U9476 (N_9476,N_9352,N_9321);
nor U9477 (N_9477,N_9385,N_9300);
xnor U9478 (N_9478,N_9261,N_9267);
xor U9479 (N_9479,N_9309,N_9241);
or U9480 (N_9480,N_9305,N_9283);
or U9481 (N_9481,N_9346,N_9204);
or U9482 (N_9482,N_9227,N_9250);
nand U9483 (N_9483,N_9332,N_9381);
and U9484 (N_9484,N_9358,N_9284);
or U9485 (N_9485,N_9333,N_9221);
xnor U9486 (N_9486,N_9257,N_9205);
nor U9487 (N_9487,N_9347,N_9377);
nand U9488 (N_9488,N_9273,N_9325);
and U9489 (N_9489,N_9260,N_9236);
and U9490 (N_9490,N_9235,N_9303);
and U9491 (N_9491,N_9330,N_9344);
nand U9492 (N_9492,N_9322,N_9329);
nand U9493 (N_9493,N_9285,N_9212);
and U9494 (N_9494,N_9228,N_9217);
and U9495 (N_9495,N_9378,N_9350);
or U9496 (N_9496,N_9326,N_9206);
nor U9497 (N_9497,N_9398,N_9302);
and U9498 (N_9498,N_9387,N_9365);
and U9499 (N_9499,N_9368,N_9203);
nor U9500 (N_9500,N_9283,N_9377);
or U9501 (N_9501,N_9365,N_9223);
nor U9502 (N_9502,N_9356,N_9231);
and U9503 (N_9503,N_9365,N_9271);
and U9504 (N_9504,N_9218,N_9374);
xnor U9505 (N_9505,N_9230,N_9337);
nand U9506 (N_9506,N_9284,N_9367);
and U9507 (N_9507,N_9292,N_9315);
and U9508 (N_9508,N_9287,N_9247);
nor U9509 (N_9509,N_9231,N_9278);
or U9510 (N_9510,N_9288,N_9227);
and U9511 (N_9511,N_9399,N_9363);
nor U9512 (N_9512,N_9334,N_9360);
xnor U9513 (N_9513,N_9363,N_9338);
nand U9514 (N_9514,N_9335,N_9250);
and U9515 (N_9515,N_9239,N_9241);
xor U9516 (N_9516,N_9225,N_9384);
nand U9517 (N_9517,N_9324,N_9396);
nand U9518 (N_9518,N_9214,N_9379);
nor U9519 (N_9519,N_9398,N_9361);
xnor U9520 (N_9520,N_9384,N_9236);
or U9521 (N_9521,N_9219,N_9262);
nand U9522 (N_9522,N_9348,N_9352);
or U9523 (N_9523,N_9251,N_9389);
or U9524 (N_9524,N_9236,N_9307);
or U9525 (N_9525,N_9284,N_9312);
nor U9526 (N_9526,N_9305,N_9206);
or U9527 (N_9527,N_9391,N_9256);
and U9528 (N_9528,N_9336,N_9327);
nor U9529 (N_9529,N_9286,N_9307);
nand U9530 (N_9530,N_9224,N_9311);
or U9531 (N_9531,N_9300,N_9279);
or U9532 (N_9532,N_9348,N_9364);
or U9533 (N_9533,N_9335,N_9305);
or U9534 (N_9534,N_9306,N_9299);
and U9535 (N_9535,N_9270,N_9291);
nor U9536 (N_9536,N_9389,N_9351);
nor U9537 (N_9537,N_9205,N_9293);
nand U9538 (N_9538,N_9315,N_9380);
or U9539 (N_9539,N_9358,N_9212);
nand U9540 (N_9540,N_9378,N_9382);
xnor U9541 (N_9541,N_9302,N_9399);
and U9542 (N_9542,N_9202,N_9310);
nand U9543 (N_9543,N_9370,N_9241);
nor U9544 (N_9544,N_9376,N_9374);
and U9545 (N_9545,N_9360,N_9348);
or U9546 (N_9546,N_9279,N_9210);
or U9547 (N_9547,N_9325,N_9285);
nand U9548 (N_9548,N_9362,N_9230);
and U9549 (N_9549,N_9300,N_9340);
nor U9550 (N_9550,N_9361,N_9351);
and U9551 (N_9551,N_9295,N_9306);
or U9552 (N_9552,N_9218,N_9384);
xnor U9553 (N_9553,N_9372,N_9282);
and U9554 (N_9554,N_9221,N_9265);
and U9555 (N_9555,N_9279,N_9397);
nor U9556 (N_9556,N_9225,N_9220);
nand U9557 (N_9557,N_9292,N_9303);
nor U9558 (N_9558,N_9333,N_9275);
nor U9559 (N_9559,N_9224,N_9316);
xor U9560 (N_9560,N_9312,N_9204);
nand U9561 (N_9561,N_9301,N_9272);
or U9562 (N_9562,N_9297,N_9200);
xnor U9563 (N_9563,N_9262,N_9280);
nor U9564 (N_9564,N_9336,N_9291);
nor U9565 (N_9565,N_9235,N_9370);
and U9566 (N_9566,N_9285,N_9294);
nor U9567 (N_9567,N_9270,N_9321);
or U9568 (N_9568,N_9275,N_9369);
nand U9569 (N_9569,N_9383,N_9390);
xnor U9570 (N_9570,N_9269,N_9367);
xor U9571 (N_9571,N_9251,N_9280);
nor U9572 (N_9572,N_9252,N_9316);
and U9573 (N_9573,N_9219,N_9283);
nand U9574 (N_9574,N_9366,N_9391);
or U9575 (N_9575,N_9381,N_9337);
and U9576 (N_9576,N_9279,N_9324);
or U9577 (N_9577,N_9348,N_9398);
or U9578 (N_9578,N_9330,N_9283);
nor U9579 (N_9579,N_9224,N_9332);
nor U9580 (N_9580,N_9288,N_9211);
nand U9581 (N_9581,N_9213,N_9245);
and U9582 (N_9582,N_9311,N_9281);
or U9583 (N_9583,N_9210,N_9289);
or U9584 (N_9584,N_9285,N_9235);
or U9585 (N_9585,N_9231,N_9205);
or U9586 (N_9586,N_9385,N_9309);
xor U9587 (N_9587,N_9214,N_9202);
or U9588 (N_9588,N_9271,N_9319);
nor U9589 (N_9589,N_9219,N_9263);
or U9590 (N_9590,N_9318,N_9226);
or U9591 (N_9591,N_9353,N_9393);
nand U9592 (N_9592,N_9315,N_9368);
nor U9593 (N_9593,N_9227,N_9358);
nor U9594 (N_9594,N_9389,N_9200);
xor U9595 (N_9595,N_9230,N_9283);
xnor U9596 (N_9596,N_9218,N_9256);
and U9597 (N_9597,N_9237,N_9371);
nand U9598 (N_9598,N_9305,N_9334);
and U9599 (N_9599,N_9274,N_9285);
nor U9600 (N_9600,N_9403,N_9544);
xnor U9601 (N_9601,N_9588,N_9454);
and U9602 (N_9602,N_9582,N_9580);
xor U9603 (N_9603,N_9466,N_9423);
nor U9604 (N_9604,N_9409,N_9504);
nor U9605 (N_9605,N_9431,N_9439);
and U9606 (N_9606,N_9595,N_9484);
nor U9607 (N_9607,N_9450,N_9438);
or U9608 (N_9608,N_9523,N_9591);
xnor U9609 (N_9609,N_9428,N_9496);
nand U9610 (N_9610,N_9557,N_9568);
or U9611 (N_9611,N_9491,N_9579);
nand U9612 (N_9612,N_9503,N_9546);
or U9613 (N_9613,N_9573,N_9448);
or U9614 (N_9614,N_9402,N_9463);
and U9615 (N_9615,N_9447,N_9485);
and U9616 (N_9616,N_9585,N_9514);
xor U9617 (N_9617,N_9455,N_9538);
and U9618 (N_9618,N_9480,N_9525);
nand U9619 (N_9619,N_9469,N_9540);
nor U9620 (N_9620,N_9482,N_9511);
and U9621 (N_9621,N_9476,N_9596);
or U9622 (N_9622,N_9433,N_9550);
nor U9623 (N_9623,N_9571,N_9471);
nand U9624 (N_9624,N_9589,N_9444);
or U9625 (N_9625,N_9489,N_9461);
nor U9626 (N_9626,N_9554,N_9578);
nand U9627 (N_9627,N_9558,N_9533);
nor U9628 (N_9628,N_9531,N_9417);
xor U9629 (N_9629,N_9590,N_9408);
or U9630 (N_9630,N_9572,N_9567);
and U9631 (N_9631,N_9518,N_9553);
and U9632 (N_9632,N_9472,N_9440);
or U9633 (N_9633,N_9495,N_9425);
nor U9634 (N_9634,N_9412,N_9537);
or U9635 (N_9635,N_9494,N_9416);
and U9636 (N_9636,N_9468,N_9493);
and U9637 (N_9637,N_9552,N_9526);
or U9638 (N_9638,N_9593,N_9509);
and U9639 (N_9639,N_9517,N_9457);
nor U9640 (N_9640,N_9551,N_9479);
nor U9641 (N_9641,N_9497,N_9547);
nand U9642 (N_9642,N_9432,N_9442);
and U9643 (N_9643,N_9422,N_9532);
and U9644 (N_9644,N_9421,N_9401);
nor U9645 (N_9645,N_9555,N_9420);
nand U9646 (N_9646,N_9445,N_9426);
nor U9647 (N_9647,N_9586,N_9404);
and U9648 (N_9648,N_9464,N_9446);
nand U9649 (N_9649,N_9477,N_9449);
or U9650 (N_9650,N_9598,N_9451);
xor U9651 (N_9651,N_9516,N_9441);
or U9652 (N_9652,N_9467,N_9599);
and U9653 (N_9653,N_9475,N_9478);
and U9654 (N_9654,N_9499,N_9597);
nand U9655 (N_9655,N_9520,N_9414);
and U9656 (N_9656,N_9453,N_9443);
xor U9657 (N_9657,N_9459,N_9508);
or U9658 (N_9658,N_9576,N_9530);
or U9659 (N_9659,N_9515,N_9456);
nand U9660 (N_9660,N_9594,N_9470);
or U9661 (N_9661,N_9498,N_9535);
nand U9662 (N_9662,N_9430,N_9566);
xor U9663 (N_9663,N_9536,N_9510);
or U9664 (N_9664,N_9565,N_9562);
nand U9665 (N_9665,N_9501,N_9587);
xnor U9666 (N_9666,N_9556,N_9542);
nor U9667 (N_9667,N_9539,N_9474);
or U9668 (N_9668,N_9505,N_9502);
nor U9669 (N_9669,N_9500,N_9490);
nand U9670 (N_9670,N_9427,N_9410);
nor U9671 (N_9671,N_9434,N_9400);
or U9672 (N_9672,N_9569,N_9481);
or U9673 (N_9673,N_9488,N_9458);
and U9674 (N_9674,N_9583,N_9521);
nor U9675 (N_9675,N_9534,N_9436);
nor U9676 (N_9676,N_9581,N_9460);
nand U9677 (N_9677,N_9524,N_9574);
xnor U9678 (N_9678,N_9473,N_9418);
and U9679 (N_9679,N_9492,N_9527);
xor U9680 (N_9680,N_9584,N_9577);
nor U9681 (N_9681,N_9413,N_9415);
or U9682 (N_9682,N_9560,N_9541);
or U9683 (N_9683,N_9545,N_9435);
and U9684 (N_9684,N_9528,N_9486);
nor U9685 (N_9685,N_9437,N_9483);
xor U9686 (N_9686,N_9592,N_9462);
xor U9687 (N_9687,N_9564,N_9419);
nor U9688 (N_9688,N_9519,N_9506);
xor U9689 (N_9689,N_9570,N_9563);
or U9690 (N_9690,N_9407,N_9548);
and U9691 (N_9691,N_9513,N_9405);
nor U9692 (N_9692,N_9512,N_9411);
or U9693 (N_9693,N_9529,N_9406);
nor U9694 (N_9694,N_9424,N_9522);
xnor U9695 (N_9695,N_9549,N_9429);
xnor U9696 (N_9696,N_9487,N_9559);
xor U9697 (N_9697,N_9507,N_9561);
and U9698 (N_9698,N_9575,N_9543);
or U9699 (N_9699,N_9452,N_9465);
or U9700 (N_9700,N_9452,N_9403);
xnor U9701 (N_9701,N_9502,N_9571);
nand U9702 (N_9702,N_9593,N_9466);
nor U9703 (N_9703,N_9519,N_9572);
or U9704 (N_9704,N_9419,N_9562);
and U9705 (N_9705,N_9501,N_9486);
nor U9706 (N_9706,N_9472,N_9538);
or U9707 (N_9707,N_9534,N_9415);
nor U9708 (N_9708,N_9553,N_9468);
nand U9709 (N_9709,N_9548,N_9444);
or U9710 (N_9710,N_9417,N_9464);
nand U9711 (N_9711,N_9554,N_9420);
nand U9712 (N_9712,N_9439,N_9404);
and U9713 (N_9713,N_9591,N_9407);
nor U9714 (N_9714,N_9570,N_9504);
nand U9715 (N_9715,N_9579,N_9460);
or U9716 (N_9716,N_9416,N_9481);
nand U9717 (N_9717,N_9597,N_9561);
nand U9718 (N_9718,N_9429,N_9452);
nor U9719 (N_9719,N_9434,N_9475);
and U9720 (N_9720,N_9538,N_9593);
or U9721 (N_9721,N_9592,N_9409);
nand U9722 (N_9722,N_9576,N_9498);
xor U9723 (N_9723,N_9450,N_9591);
and U9724 (N_9724,N_9417,N_9410);
and U9725 (N_9725,N_9498,N_9570);
or U9726 (N_9726,N_9518,N_9508);
nand U9727 (N_9727,N_9444,N_9465);
nand U9728 (N_9728,N_9489,N_9551);
xor U9729 (N_9729,N_9517,N_9502);
or U9730 (N_9730,N_9565,N_9486);
and U9731 (N_9731,N_9475,N_9413);
xnor U9732 (N_9732,N_9559,N_9567);
nor U9733 (N_9733,N_9532,N_9409);
and U9734 (N_9734,N_9432,N_9571);
nor U9735 (N_9735,N_9420,N_9516);
xnor U9736 (N_9736,N_9456,N_9572);
xor U9737 (N_9737,N_9523,N_9467);
xnor U9738 (N_9738,N_9505,N_9473);
and U9739 (N_9739,N_9542,N_9534);
nor U9740 (N_9740,N_9426,N_9548);
and U9741 (N_9741,N_9483,N_9581);
nand U9742 (N_9742,N_9528,N_9563);
or U9743 (N_9743,N_9589,N_9594);
nor U9744 (N_9744,N_9596,N_9570);
or U9745 (N_9745,N_9543,N_9558);
nand U9746 (N_9746,N_9402,N_9459);
and U9747 (N_9747,N_9419,N_9581);
nand U9748 (N_9748,N_9453,N_9559);
nor U9749 (N_9749,N_9482,N_9595);
xor U9750 (N_9750,N_9436,N_9492);
and U9751 (N_9751,N_9543,N_9495);
xor U9752 (N_9752,N_9541,N_9591);
xor U9753 (N_9753,N_9466,N_9543);
and U9754 (N_9754,N_9552,N_9429);
or U9755 (N_9755,N_9555,N_9445);
nor U9756 (N_9756,N_9482,N_9548);
xor U9757 (N_9757,N_9542,N_9503);
xor U9758 (N_9758,N_9488,N_9439);
xnor U9759 (N_9759,N_9458,N_9486);
and U9760 (N_9760,N_9539,N_9438);
xor U9761 (N_9761,N_9409,N_9480);
xnor U9762 (N_9762,N_9415,N_9542);
xor U9763 (N_9763,N_9410,N_9489);
nand U9764 (N_9764,N_9554,N_9489);
and U9765 (N_9765,N_9526,N_9489);
or U9766 (N_9766,N_9566,N_9496);
and U9767 (N_9767,N_9554,N_9433);
nand U9768 (N_9768,N_9439,N_9496);
nor U9769 (N_9769,N_9528,N_9451);
nor U9770 (N_9770,N_9558,N_9587);
nor U9771 (N_9771,N_9475,N_9449);
or U9772 (N_9772,N_9557,N_9551);
nand U9773 (N_9773,N_9536,N_9425);
or U9774 (N_9774,N_9482,N_9557);
and U9775 (N_9775,N_9494,N_9551);
nor U9776 (N_9776,N_9484,N_9555);
xnor U9777 (N_9777,N_9460,N_9437);
nand U9778 (N_9778,N_9574,N_9473);
or U9779 (N_9779,N_9473,N_9462);
xnor U9780 (N_9780,N_9596,N_9423);
and U9781 (N_9781,N_9405,N_9435);
xor U9782 (N_9782,N_9411,N_9410);
nand U9783 (N_9783,N_9415,N_9406);
and U9784 (N_9784,N_9527,N_9453);
nand U9785 (N_9785,N_9591,N_9461);
and U9786 (N_9786,N_9418,N_9421);
nand U9787 (N_9787,N_9458,N_9574);
and U9788 (N_9788,N_9547,N_9593);
or U9789 (N_9789,N_9596,N_9513);
and U9790 (N_9790,N_9432,N_9462);
and U9791 (N_9791,N_9498,N_9548);
nand U9792 (N_9792,N_9558,N_9555);
nor U9793 (N_9793,N_9518,N_9421);
xnor U9794 (N_9794,N_9400,N_9403);
and U9795 (N_9795,N_9581,N_9509);
nand U9796 (N_9796,N_9575,N_9556);
nand U9797 (N_9797,N_9404,N_9536);
nand U9798 (N_9798,N_9451,N_9573);
and U9799 (N_9799,N_9440,N_9530);
xor U9800 (N_9800,N_9792,N_9732);
nor U9801 (N_9801,N_9717,N_9692);
or U9802 (N_9802,N_9740,N_9691);
xor U9803 (N_9803,N_9693,N_9775);
xnor U9804 (N_9804,N_9615,N_9795);
or U9805 (N_9805,N_9751,N_9741);
nor U9806 (N_9806,N_9648,N_9799);
nor U9807 (N_9807,N_9722,N_9632);
nor U9808 (N_9808,N_9603,N_9619);
or U9809 (N_9809,N_9781,N_9748);
xnor U9810 (N_9810,N_9716,N_9734);
nor U9811 (N_9811,N_9678,N_9672);
nand U9812 (N_9812,N_9778,N_9773);
xnor U9813 (N_9813,N_9701,N_9765);
xnor U9814 (N_9814,N_9736,N_9770);
and U9815 (N_9815,N_9608,N_9735);
nand U9816 (N_9816,N_9629,N_9784);
nand U9817 (N_9817,N_9779,N_9798);
or U9818 (N_9818,N_9675,N_9746);
and U9819 (N_9819,N_9652,N_9647);
and U9820 (N_9820,N_9663,N_9626);
or U9821 (N_9821,N_9636,N_9610);
nor U9822 (N_9822,N_9657,N_9646);
nand U9823 (N_9823,N_9762,N_9714);
nand U9824 (N_9824,N_9669,N_9712);
nor U9825 (N_9825,N_9612,N_9682);
and U9826 (N_9826,N_9627,N_9709);
nand U9827 (N_9827,N_9640,N_9763);
and U9828 (N_9828,N_9679,N_9630);
xor U9829 (N_9829,N_9644,N_9606);
or U9830 (N_9830,N_9694,N_9670);
or U9831 (N_9831,N_9638,N_9757);
or U9832 (N_9832,N_9768,N_9696);
xor U9833 (N_9833,N_9700,N_9789);
and U9834 (N_9834,N_9786,N_9634);
or U9835 (N_9835,N_9726,N_9689);
nand U9836 (N_9836,N_9643,N_9797);
nand U9837 (N_9837,N_9738,N_9686);
nand U9838 (N_9838,N_9720,N_9767);
xnor U9839 (N_9839,N_9725,N_9739);
and U9840 (N_9840,N_9618,N_9713);
xor U9841 (N_9841,N_9637,N_9649);
or U9842 (N_9842,N_9698,N_9769);
nor U9843 (N_9843,N_9614,N_9774);
or U9844 (N_9844,N_9661,N_9704);
xor U9845 (N_9845,N_9695,N_9705);
or U9846 (N_9846,N_9656,N_9707);
nand U9847 (N_9847,N_9699,N_9772);
nand U9848 (N_9848,N_9756,N_9723);
and U9849 (N_9849,N_9783,N_9605);
nor U9850 (N_9850,N_9766,N_9787);
xnor U9851 (N_9851,N_9688,N_9750);
nand U9852 (N_9852,N_9613,N_9651);
xnor U9853 (N_9853,N_9602,N_9758);
or U9854 (N_9854,N_9666,N_9664);
or U9855 (N_9855,N_9743,N_9650);
nor U9856 (N_9856,N_9607,N_9753);
and U9857 (N_9857,N_9780,N_9761);
nor U9858 (N_9858,N_9622,N_9633);
and U9859 (N_9859,N_9760,N_9715);
xnor U9860 (N_9860,N_9794,N_9628);
nor U9861 (N_9861,N_9641,N_9600);
or U9862 (N_9862,N_9677,N_9673);
and U9863 (N_9863,N_9729,N_9796);
and U9864 (N_9864,N_9771,N_9625);
nand U9865 (N_9865,N_9690,N_9676);
xor U9866 (N_9866,N_9730,N_9721);
nor U9867 (N_9867,N_9711,N_9731);
xor U9868 (N_9868,N_9737,N_9621);
or U9869 (N_9869,N_9755,N_9684);
xor U9870 (N_9870,N_9665,N_9604);
or U9871 (N_9871,N_9645,N_9710);
and U9872 (N_9872,N_9759,N_9655);
xor U9873 (N_9873,N_9687,N_9790);
nand U9874 (N_9874,N_9706,N_9616);
nand U9875 (N_9875,N_9718,N_9658);
nor U9876 (N_9876,N_9788,N_9754);
or U9877 (N_9877,N_9642,N_9683);
xor U9878 (N_9878,N_9660,N_9659);
or U9879 (N_9879,N_9703,N_9620);
nand U9880 (N_9880,N_9785,N_9601);
and U9881 (N_9881,N_9609,N_9776);
and U9882 (N_9882,N_9719,N_9728);
and U9883 (N_9883,N_9733,N_9662);
xnor U9884 (N_9884,N_9671,N_9653);
or U9885 (N_9885,N_9680,N_9611);
nor U9886 (N_9886,N_9702,N_9749);
nor U9887 (N_9887,N_9617,N_9668);
or U9888 (N_9888,N_9744,N_9745);
or U9889 (N_9889,N_9747,N_9635);
xor U9890 (N_9890,N_9697,N_9681);
xnor U9891 (N_9891,N_9782,N_9724);
nor U9892 (N_9892,N_9752,N_9654);
nor U9893 (N_9893,N_9674,N_9623);
and U9894 (N_9894,N_9791,N_9624);
nand U9895 (N_9895,N_9727,N_9631);
or U9896 (N_9896,N_9742,N_9777);
and U9897 (N_9897,N_9685,N_9793);
nor U9898 (N_9898,N_9764,N_9639);
nand U9899 (N_9899,N_9708,N_9667);
and U9900 (N_9900,N_9666,N_9685);
nor U9901 (N_9901,N_9674,N_9677);
nor U9902 (N_9902,N_9704,N_9799);
xor U9903 (N_9903,N_9757,N_9654);
nand U9904 (N_9904,N_9775,N_9691);
nor U9905 (N_9905,N_9788,N_9645);
nor U9906 (N_9906,N_9697,N_9623);
nor U9907 (N_9907,N_9633,N_9722);
nor U9908 (N_9908,N_9641,N_9674);
nor U9909 (N_9909,N_9625,N_9665);
and U9910 (N_9910,N_9609,N_9714);
or U9911 (N_9911,N_9765,N_9633);
or U9912 (N_9912,N_9674,N_9654);
xnor U9913 (N_9913,N_9611,N_9722);
and U9914 (N_9914,N_9677,N_9755);
nor U9915 (N_9915,N_9785,N_9602);
xnor U9916 (N_9916,N_9687,N_9635);
nand U9917 (N_9917,N_9661,N_9639);
nor U9918 (N_9918,N_9740,N_9786);
xnor U9919 (N_9919,N_9705,N_9772);
xnor U9920 (N_9920,N_9771,N_9742);
nor U9921 (N_9921,N_9688,N_9762);
or U9922 (N_9922,N_9692,N_9796);
nand U9923 (N_9923,N_9723,N_9747);
nand U9924 (N_9924,N_9643,N_9612);
or U9925 (N_9925,N_9666,N_9756);
xor U9926 (N_9926,N_9787,N_9658);
xor U9927 (N_9927,N_9611,N_9795);
nand U9928 (N_9928,N_9742,N_9715);
and U9929 (N_9929,N_9783,N_9671);
or U9930 (N_9930,N_9720,N_9743);
and U9931 (N_9931,N_9687,N_9664);
nand U9932 (N_9932,N_9738,N_9718);
and U9933 (N_9933,N_9622,N_9757);
xnor U9934 (N_9934,N_9728,N_9696);
or U9935 (N_9935,N_9699,N_9724);
nor U9936 (N_9936,N_9785,N_9711);
or U9937 (N_9937,N_9659,N_9752);
and U9938 (N_9938,N_9673,N_9772);
nand U9939 (N_9939,N_9695,N_9625);
and U9940 (N_9940,N_9768,N_9638);
nand U9941 (N_9941,N_9669,N_9762);
xnor U9942 (N_9942,N_9643,N_9783);
xor U9943 (N_9943,N_9792,N_9691);
nor U9944 (N_9944,N_9759,N_9753);
and U9945 (N_9945,N_9675,N_9631);
nor U9946 (N_9946,N_9652,N_9780);
nor U9947 (N_9947,N_9602,N_9737);
nand U9948 (N_9948,N_9712,N_9699);
nor U9949 (N_9949,N_9772,N_9613);
nor U9950 (N_9950,N_9628,N_9629);
xor U9951 (N_9951,N_9717,N_9699);
nor U9952 (N_9952,N_9789,N_9726);
nor U9953 (N_9953,N_9641,N_9643);
xor U9954 (N_9954,N_9683,N_9659);
nor U9955 (N_9955,N_9717,N_9759);
and U9956 (N_9956,N_9729,N_9679);
or U9957 (N_9957,N_9796,N_9633);
nor U9958 (N_9958,N_9638,N_9616);
nand U9959 (N_9959,N_9756,N_9783);
xor U9960 (N_9960,N_9780,N_9731);
xor U9961 (N_9961,N_9719,N_9761);
xor U9962 (N_9962,N_9612,N_9683);
or U9963 (N_9963,N_9652,N_9749);
xnor U9964 (N_9964,N_9652,N_9798);
nand U9965 (N_9965,N_9719,N_9792);
xnor U9966 (N_9966,N_9711,N_9727);
or U9967 (N_9967,N_9639,N_9772);
and U9968 (N_9968,N_9660,N_9651);
and U9969 (N_9969,N_9619,N_9627);
and U9970 (N_9970,N_9601,N_9758);
nand U9971 (N_9971,N_9614,N_9627);
nand U9972 (N_9972,N_9759,N_9764);
nand U9973 (N_9973,N_9648,N_9634);
nand U9974 (N_9974,N_9775,N_9610);
nor U9975 (N_9975,N_9732,N_9666);
nor U9976 (N_9976,N_9682,N_9746);
and U9977 (N_9977,N_9603,N_9680);
or U9978 (N_9978,N_9663,N_9634);
nand U9979 (N_9979,N_9725,N_9638);
or U9980 (N_9980,N_9749,N_9690);
nor U9981 (N_9981,N_9611,N_9767);
nor U9982 (N_9982,N_9706,N_9702);
or U9983 (N_9983,N_9649,N_9790);
and U9984 (N_9984,N_9730,N_9636);
or U9985 (N_9985,N_9687,N_9763);
nand U9986 (N_9986,N_9707,N_9651);
nand U9987 (N_9987,N_9779,N_9602);
xnor U9988 (N_9988,N_9652,N_9727);
nor U9989 (N_9989,N_9747,N_9780);
or U9990 (N_9990,N_9760,N_9774);
nand U9991 (N_9991,N_9735,N_9666);
nor U9992 (N_9992,N_9764,N_9690);
nand U9993 (N_9993,N_9790,N_9673);
xnor U9994 (N_9994,N_9634,N_9754);
or U9995 (N_9995,N_9729,N_9622);
or U9996 (N_9996,N_9690,N_9645);
nor U9997 (N_9997,N_9741,N_9708);
xor U9998 (N_9998,N_9712,N_9770);
nor U9999 (N_9999,N_9653,N_9677);
xnor U10000 (N_10000,N_9826,N_9803);
or U10001 (N_10001,N_9890,N_9867);
nor U10002 (N_10002,N_9897,N_9889);
nor U10003 (N_10003,N_9933,N_9992);
nand U10004 (N_10004,N_9962,N_9991);
or U10005 (N_10005,N_9809,N_9912);
and U10006 (N_10006,N_9902,N_9996);
nand U10007 (N_10007,N_9925,N_9972);
and U10008 (N_10008,N_9917,N_9949);
nand U10009 (N_10009,N_9885,N_9987);
or U10010 (N_10010,N_9907,N_9979);
and U10011 (N_10011,N_9805,N_9873);
nand U10012 (N_10012,N_9845,N_9927);
nor U10013 (N_10013,N_9994,N_9843);
nor U10014 (N_10014,N_9888,N_9801);
nand U10015 (N_10015,N_9938,N_9945);
nand U10016 (N_10016,N_9922,N_9831);
or U10017 (N_10017,N_9971,N_9862);
or U10018 (N_10018,N_9977,N_9984);
nor U10019 (N_10019,N_9882,N_9837);
nand U10020 (N_10020,N_9856,N_9956);
nor U10021 (N_10021,N_9995,N_9986);
and U10022 (N_10022,N_9869,N_9930);
and U10023 (N_10023,N_9921,N_9865);
xor U10024 (N_10024,N_9828,N_9924);
or U10025 (N_10025,N_9963,N_9827);
and U10026 (N_10026,N_9881,N_9957);
and U10027 (N_10027,N_9834,N_9931);
nand U10028 (N_10028,N_9838,N_9948);
nand U10029 (N_10029,N_9969,N_9974);
nand U10030 (N_10030,N_9981,N_9893);
nor U10031 (N_10031,N_9959,N_9887);
or U10032 (N_10032,N_9989,N_9965);
or U10033 (N_10033,N_9941,N_9944);
nor U10034 (N_10034,N_9901,N_9868);
nand U10035 (N_10035,N_9980,N_9810);
nor U10036 (N_10036,N_9999,N_9990);
xor U10037 (N_10037,N_9906,N_9832);
and U10038 (N_10038,N_9821,N_9952);
or U10039 (N_10039,N_9839,N_9954);
or U10040 (N_10040,N_9823,N_9947);
nor U10041 (N_10041,N_9825,N_9848);
or U10042 (N_10042,N_9892,N_9814);
or U10043 (N_10043,N_9966,N_9960);
nor U10044 (N_10044,N_9951,N_9953);
nand U10045 (N_10045,N_9985,N_9864);
nand U10046 (N_10046,N_9935,N_9998);
xor U10047 (N_10047,N_9928,N_9855);
nand U10048 (N_10048,N_9886,N_9860);
xor U10049 (N_10049,N_9923,N_9807);
nand U10050 (N_10050,N_9911,N_9894);
and U10051 (N_10051,N_9820,N_9849);
nor U10052 (N_10052,N_9877,N_9905);
and U10053 (N_10053,N_9942,N_9940);
and U10054 (N_10054,N_9878,N_9866);
nand U10055 (N_10055,N_9920,N_9851);
nor U10056 (N_10056,N_9936,N_9909);
and U10057 (N_10057,N_9943,N_9958);
nand U10058 (N_10058,N_9816,N_9926);
nor U10059 (N_10059,N_9910,N_9833);
nor U10060 (N_10060,N_9968,N_9871);
or U10061 (N_10061,N_9817,N_9844);
nor U10062 (N_10062,N_9880,N_9808);
or U10063 (N_10063,N_9861,N_9883);
and U10064 (N_10064,N_9993,N_9847);
xnor U10065 (N_10065,N_9819,N_9876);
nand U10066 (N_10066,N_9852,N_9811);
and U10067 (N_10067,N_9982,N_9891);
or U10068 (N_10068,N_9997,N_9896);
or U10069 (N_10069,N_9824,N_9854);
nand U10070 (N_10070,N_9950,N_9908);
xnor U10071 (N_10071,N_9964,N_9970);
xor U10072 (N_10072,N_9858,N_9975);
and U10073 (N_10073,N_9872,N_9903);
and U10074 (N_10074,N_9988,N_9812);
xnor U10075 (N_10075,N_9874,N_9946);
nor U10076 (N_10076,N_9967,N_9904);
xor U10077 (N_10077,N_9863,N_9850);
or U10078 (N_10078,N_9914,N_9840);
or U10079 (N_10079,N_9802,N_9934);
and U10080 (N_10080,N_9815,N_9879);
xnor U10081 (N_10081,N_9929,N_9898);
or U10082 (N_10082,N_9961,N_9853);
and U10083 (N_10083,N_9916,N_9813);
or U10084 (N_10084,N_9842,N_9915);
nor U10085 (N_10085,N_9875,N_9841);
and U10086 (N_10086,N_9804,N_9937);
and U10087 (N_10087,N_9913,N_9870);
nor U10088 (N_10088,N_9835,N_9806);
xor U10089 (N_10089,N_9932,N_9857);
and U10090 (N_10090,N_9884,N_9830);
nand U10091 (N_10091,N_9895,N_9822);
or U10092 (N_10092,N_9846,N_9976);
and U10093 (N_10093,N_9919,N_9983);
xor U10094 (N_10094,N_9955,N_9818);
xor U10095 (N_10095,N_9900,N_9829);
nand U10096 (N_10096,N_9939,N_9859);
nand U10097 (N_10097,N_9973,N_9918);
nor U10098 (N_10098,N_9836,N_9899);
nor U10099 (N_10099,N_9978,N_9800);
nand U10100 (N_10100,N_9813,N_9849);
nand U10101 (N_10101,N_9984,N_9846);
and U10102 (N_10102,N_9838,N_9908);
or U10103 (N_10103,N_9806,N_9923);
nand U10104 (N_10104,N_9859,N_9877);
nor U10105 (N_10105,N_9985,N_9906);
nand U10106 (N_10106,N_9848,N_9988);
or U10107 (N_10107,N_9831,N_9850);
nand U10108 (N_10108,N_9813,N_9914);
xnor U10109 (N_10109,N_9920,N_9909);
and U10110 (N_10110,N_9810,N_9965);
nor U10111 (N_10111,N_9909,N_9956);
nor U10112 (N_10112,N_9907,N_9936);
or U10113 (N_10113,N_9884,N_9912);
nand U10114 (N_10114,N_9915,N_9955);
and U10115 (N_10115,N_9834,N_9807);
nand U10116 (N_10116,N_9911,N_9974);
nand U10117 (N_10117,N_9995,N_9855);
nand U10118 (N_10118,N_9976,N_9927);
nand U10119 (N_10119,N_9909,N_9892);
xnor U10120 (N_10120,N_9970,N_9885);
or U10121 (N_10121,N_9912,N_9808);
nand U10122 (N_10122,N_9924,N_9947);
nand U10123 (N_10123,N_9977,N_9880);
nand U10124 (N_10124,N_9908,N_9882);
nor U10125 (N_10125,N_9805,N_9838);
nand U10126 (N_10126,N_9824,N_9929);
nand U10127 (N_10127,N_9971,N_9898);
nor U10128 (N_10128,N_9955,N_9896);
xnor U10129 (N_10129,N_9802,N_9844);
and U10130 (N_10130,N_9817,N_9935);
nand U10131 (N_10131,N_9869,N_9919);
or U10132 (N_10132,N_9954,N_9858);
or U10133 (N_10133,N_9908,N_9987);
nand U10134 (N_10134,N_9881,N_9883);
nand U10135 (N_10135,N_9906,N_9975);
xnor U10136 (N_10136,N_9912,N_9872);
or U10137 (N_10137,N_9922,N_9879);
nand U10138 (N_10138,N_9962,N_9846);
nor U10139 (N_10139,N_9908,N_9862);
and U10140 (N_10140,N_9992,N_9944);
nand U10141 (N_10141,N_9839,N_9882);
nor U10142 (N_10142,N_9830,N_9846);
nand U10143 (N_10143,N_9908,N_9819);
and U10144 (N_10144,N_9967,N_9932);
nand U10145 (N_10145,N_9989,N_9898);
and U10146 (N_10146,N_9867,N_9985);
or U10147 (N_10147,N_9957,N_9981);
nor U10148 (N_10148,N_9926,N_9881);
xor U10149 (N_10149,N_9840,N_9843);
and U10150 (N_10150,N_9837,N_9938);
and U10151 (N_10151,N_9917,N_9948);
nor U10152 (N_10152,N_9836,N_9824);
nor U10153 (N_10153,N_9811,N_9938);
and U10154 (N_10154,N_9947,N_9920);
nor U10155 (N_10155,N_9816,N_9989);
nand U10156 (N_10156,N_9946,N_9835);
and U10157 (N_10157,N_9871,N_9822);
or U10158 (N_10158,N_9811,N_9930);
and U10159 (N_10159,N_9888,N_9964);
xor U10160 (N_10160,N_9893,N_9898);
and U10161 (N_10161,N_9998,N_9804);
nand U10162 (N_10162,N_9979,N_9816);
xor U10163 (N_10163,N_9942,N_9939);
nor U10164 (N_10164,N_9969,N_9922);
and U10165 (N_10165,N_9949,N_9827);
or U10166 (N_10166,N_9824,N_9935);
and U10167 (N_10167,N_9854,N_9846);
xor U10168 (N_10168,N_9993,N_9880);
nand U10169 (N_10169,N_9902,N_9994);
or U10170 (N_10170,N_9923,N_9867);
xnor U10171 (N_10171,N_9866,N_9857);
or U10172 (N_10172,N_9927,N_9803);
xnor U10173 (N_10173,N_9932,N_9971);
nor U10174 (N_10174,N_9931,N_9830);
nor U10175 (N_10175,N_9831,N_9857);
xnor U10176 (N_10176,N_9874,N_9806);
nand U10177 (N_10177,N_9955,N_9879);
nand U10178 (N_10178,N_9973,N_9924);
nor U10179 (N_10179,N_9913,N_9915);
nor U10180 (N_10180,N_9898,N_9814);
and U10181 (N_10181,N_9864,N_9989);
xnor U10182 (N_10182,N_9845,N_9982);
nor U10183 (N_10183,N_9938,N_9956);
and U10184 (N_10184,N_9807,N_9830);
or U10185 (N_10185,N_9980,N_9910);
nor U10186 (N_10186,N_9917,N_9936);
xnor U10187 (N_10187,N_9856,N_9822);
or U10188 (N_10188,N_9852,N_9815);
or U10189 (N_10189,N_9908,N_9832);
nand U10190 (N_10190,N_9896,N_9969);
xnor U10191 (N_10191,N_9808,N_9889);
xnor U10192 (N_10192,N_9866,N_9917);
nor U10193 (N_10193,N_9984,N_9854);
xnor U10194 (N_10194,N_9869,N_9971);
nor U10195 (N_10195,N_9916,N_9962);
xnor U10196 (N_10196,N_9958,N_9911);
xnor U10197 (N_10197,N_9817,N_9920);
or U10198 (N_10198,N_9870,N_9985);
or U10199 (N_10199,N_9949,N_9975);
nand U10200 (N_10200,N_10046,N_10196);
nor U10201 (N_10201,N_10000,N_10020);
nand U10202 (N_10202,N_10002,N_10098);
and U10203 (N_10203,N_10092,N_10106);
xnor U10204 (N_10204,N_10141,N_10067);
and U10205 (N_10205,N_10198,N_10191);
and U10206 (N_10206,N_10073,N_10057);
nand U10207 (N_10207,N_10039,N_10111);
and U10208 (N_10208,N_10012,N_10147);
nor U10209 (N_10209,N_10010,N_10154);
nand U10210 (N_10210,N_10116,N_10108);
and U10211 (N_10211,N_10014,N_10053);
and U10212 (N_10212,N_10072,N_10150);
xnor U10213 (N_10213,N_10120,N_10084);
or U10214 (N_10214,N_10097,N_10100);
nand U10215 (N_10215,N_10135,N_10071);
xnor U10216 (N_10216,N_10048,N_10146);
nor U10217 (N_10217,N_10035,N_10037);
nor U10218 (N_10218,N_10021,N_10158);
xor U10219 (N_10219,N_10043,N_10132);
or U10220 (N_10220,N_10065,N_10041);
xnor U10221 (N_10221,N_10190,N_10159);
and U10222 (N_10222,N_10110,N_10181);
and U10223 (N_10223,N_10164,N_10183);
or U10224 (N_10224,N_10082,N_10155);
or U10225 (N_10225,N_10042,N_10031);
and U10226 (N_10226,N_10079,N_10160);
and U10227 (N_10227,N_10173,N_10148);
nor U10228 (N_10228,N_10194,N_10033);
nor U10229 (N_10229,N_10130,N_10161);
nor U10230 (N_10230,N_10124,N_10142);
and U10231 (N_10231,N_10143,N_10023);
or U10232 (N_10232,N_10001,N_10015);
xor U10233 (N_10233,N_10123,N_10151);
and U10234 (N_10234,N_10188,N_10032);
nor U10235 (N_10235,N_10118,N_10126);
and U10236 (N_10236,N_10077,N_10176);
nor U10237 (N_10237,N_10127,N_10112);
xnor U10238 (N_10238,N_10027,N_10099);
nor U10239 (N_10239,N_10066,N_10051);
nor U10240 (N_10240,N_10102,N_10007);
nand U10241 (N_10241,N_10004,N_10081);
or U10242 (N_10242,N_10018,N_10045);
or U10243 (N_10243,N_10166,N_10179);
or U10244 (N_10244,N_10157,N_10115);
nand U10245 (N_10245,N_10145,N_10090);
nand U10246 (N_10246,N_10061,N_10131);
and U10247 (N_10247,N_10133,N_10156);
nor U10248 (N_10248,N_10059,N_10063);
and U10249 (N_10249,N_10034,N_10017);
xnor U10250 (N_10250,N_10186,N_10170);
nand U10251 (N_10251,N_10008,N_10144);
nor U10252 (N_10252,N_10050,N_10013);
xnor U10253 (N_10253,N_10049,N_10128);
or U10254 (N_10254,N_10189,N_10094);
nand U10255 (N_10255,N_10006,N_10058);
or U10256 (N_10256,N_10182,N_10119);
nor U10257 (N_10257,N_10138,N_10104);
and U10258 (N_10258,N_10140,N_10083);
nor U10259 (N_10259,N_10174,N_10184);
nor U10260 (N_10260,N_10019,N_10047);
nor U10261 (N_10261,N_10187,N_10080);
nand U10262 (N_10262,N_10022,N_10134);
and U10263 (N_10263,N_10056,N_10030);
or U10264 (N_10264,N_10093,N_10052);
or U10265 (N_10265,N_10162,N_10011);
xor U10266 (N_10266,N_10152,N_10070);
nor U10267 (N_10267,N_10180,N_10168);
or U10268 (N_10268,N_10025,N_10029);
xor U10269 (N_10269,N_10105,N_10064);
nand U10270 (N_10270,N_10129,N_10171);
or U10271 (N_10271,N_10195,N_10177);
xnor U10272 (N_10272,N_10044,N_10193);
or U10273 (N_10273,N_10103,N_10062);
and U10274 (N_10274,N_10026,N_10109);
and U10275 (N_10275,N_10096,N_10085);
or U10276 (N_10276,N_10121,N_10016);
xor U10277 (N_10277,N_10076,N_10172);
or U10278 (N_10278,N_10038,N_10192);
nor U10279 (N_10279,N_10122,N_10087);
nand U10280 (N_10280,N_10054,N_10153);
or U10281 (N_10281,N_10089,N_10101);
and U10282 (N_10282,N_10024,N_10003);
and U10283 (N_10283,N_10197,N_10068);
xnor U10284 (N_10284,N_10175,N_10091);
or U10285 (N_10285,N_10149,N_10117);
and U10286 (N_10286,N_10163,N_10036);
nand U10287 (N_10287,N_10167,N_10075);
nor U10288 (N_10288,N_10199,N_10107);
nand U10289 (N_10289,N_10040,N_10055);
and U10290 (N_10290,N_10113,N_10028);
xnor U10291 (N_10291,N_10078,N_10069);
and U10292 (N_10292,N_10136,N_10005);
or U10293 (N_10293,N_10074,N_10114);
nor U10294 (N_10294,N_10185,N_10169);
nor U10295 (N_10295,N_10060,N_10178);
or U10296 (N_10296,N_10125,N_10009);
and U10297 (N_10297,N_10086,N_10139);
nor U10298 (N_10298,N_10095,N_10088);
and U10299 (N_10299,N_10165,N_10137);
nor U10300 (N_10300,N_10070,N_10099);
nor U10301 (N_10301,N_10020,N_10178);
or U10302 (N_10302,N_10175,N_10066);
nand U10303 (N_10303,N_10171,N_10091);
xor U10304 (N_10304,N_10003,N_10127);
nor U10305 (N_10305,N_10156,N_10194);
or U10306 (N_10306,N_10084,N_10022);
or U10307 (N_10307,N_10023,N_10108);
and U10308 (N_10308,N_10063,N_10162);
or U10309 (N_10309,N_10017,N_10126);
or U10310 (N_10310,N_10120,N_10086);
xor U10311 (N_10311,N_10179,N_10128);
or U10312 (N_10312,N_10016,N_10066);
xnor U10313 (N_10313,N_10115,N_10006);
and U10314 (N_10314,N_10069,N_10079);
nand U10315 (N_10315,N_10008,N_10096);
and U10316 (N_10316,N_10139,N_10013);
and U10317 (N_10317,N_10102,N_10171);
nand U10318 (N_10318,N_10173,N_10163);
and U10319 (N_10319,N_10002,N_10179);
or U10320 (N_10320,N_10024,N_10076);
or U10321 (N_10321,N_10146,N_10151);
xor U10322 (N_10322,N_10102,N_10049);
nand U10323 (N_10323,N_10167,N_10089);
or U10324 (N_10324,N_10040,N_10140);
or U10325 (N_10325,N_10098,N_10058);
or U10326 (N_10326,N_10083,N_10161);
nand U10327 (N_10327,N_10155,N_10163);
or U10328 (N_10328,N_10119,N_10048);
xnor U10329 (N_10329,N_10047,N_10055);
xor U10330 (N_10330,N_10175,N_10070);
xor U10331 (N_10331,N_10089,N_10132);
xnor U10332 (N_10332,N_10108,N_10028);
nor U10333 (N_10333,N_10020,N_10050);
or U10334 (N_10334,N_10096,N_10083);
nand U10335 (N_10335,N_10105,N_10194);
or U10336 (N_10336,N_10019,N_10135);
nand U10337 (N_10337,N_10153,N_10118);
or U10338 (N_10338,N_10031,N_10199);
nand U10339 (N_10339,N_10029,N_10003);
or U10340 (N_10340,N_10147,N_10011);
and U10341 (N_10341,N_10139,N_10006);
nand U10342 (N_10342,N_10015,N_10197);
nand U10343 (N_10343,N_10005,N_10056);
and U10344 (N_10344,N_10107,N_10169);
and U10345 (N_10345,N_10155,N_10021);
nor U10346 (N_10346,N_10127,N_10194);
and U10347 (N_10347,N_10091,N_10086);
xor U10348 (N_10348,N_10078,N_10145);
and U10349 (N_10349,N_10145,N_10077);
nand U10350 (N_10350,N_10006,N_10104);
or U10351 (N_10351,N_10148,N_10104);
nor U10352 (N_10352,N_10161,N_10120);
and U10353 (N_10353,N_10039,N_10031);
and U10354 (N_10354,N_10105,N_10011);
nand U10355 (N_10355,N_10103,N_10001);
nor U10356 (N_10356,N_10133,N_10072);
or U10357 (N_10357,N_10164,N_10113);
and U10358 (N_10358,N_10069,N_10083);
or U10359 (N_10359,N_10018,N_10060);
or U10360 (N_10360,N_10197,N_10142);
nor U10361 (N_10361,N_10036,N_10141);
xor U10362 (N_10362,N_10093,N_10080);
nor U10363 (N_10363,N_10079,N_10169);
and U10364 (N_10364,N_10198,N_10112);
nand U10365 (N_10365,N_10086,N_10020);
or U10366 (N_10366,N_10000,N_10022);
nand U10367 (N_10367,N_10094,N_10180);
or U10368 (N_10368,N_10117,N_10018);
or U10369 (N_10369,N_10134,N_10173);
nand U10370 (N_10370,N_10010,N_10182);
xor U10371 (N_10371,N_10016,N_10026);
nor U10372 (N_10372,N_10184,N_10164);
nand U10373 (N_10373,N_10022,N_10035);
or U10374 (N_10374,N_10177,N_10154);
xnor U10375 (N_10375,N_10096,N_10077);
nand U10376 (N_10376,N_10057,N_10098);
nand U10377 (N_10377,N_10056,N_10115);
nand U10378 (N_10378,N_10040,N_10132);
nor U10379 (N_10379,N_10044,N_10005);
and U10380 (N_10380,N_10014,N_10025);
and U10381 (N_10381,N_10187,N_10188);
xor U10382 (N_10382,N_10021,N_10034);
nand U10383 (N_10383,N_10187,N_10140);
xor U10384 (N_10384,N_10026,N_10092);
nand U10385 (N_10385,N_10068,N_10027);
or U10386 (N_10386,N_10014,N_10129);
or U10387 (N_10387,N_10021,N_10127);
xor U10388 (N_10388,N_10152,N_10125);
nand U10389 (N_10389,N_10080,N_10180);
xnor U10390 (N_10390,N_10150,N_10160);
nor U10391 (N_10391,N_10045,N_10032);
or U10392 (N_10392,N_10194,N_10120);
xnor U10393 (N_10393,N_10008,N_10169);
nand U10394 (N_10394,N_10016,N_10148);
and U10395 (N_10395,N_10110,N_10006);
xor U10396 (N_10396,N_10021,N_10105);
and U10397 (N_10397,N_10173,N_10029);
xor U10398 (N_10398,N_10078,N_10156);
or U10399 (N_10399,N_10018,N_10056);
nand U10400 (N_10400,N_10268,N_10296);
nand U10401 (N_10401,N_10346,N_10228);
or U10402 (N_10402,N_10306,N_10290);
xnor U10403 (N_10403,N_10374,N_10235);
nor U10404 (N_10404,N_10365,N_10261);
nor U10405 (N_10405,N_10209,N_10264);
and U10406 (N_10406,N_10387,N_10210);
nor U10407 (N_10407,N_10372,N_10240);
xor U10408 (N_10408,N_10398,N_10300);
and U10409 (N_10409,N_10325,N_10265);
nand U10410 (N_10410,N_10285,N_10271);
xor U10411 (N_10411,N_10330,N_10313);
and U10412 (N_10412,N_10348,N_10280);
xor U10413 (N_10413,N_10308,N_10212);
or U10414 (N_10414,N_10328,N_10294);
nand U10415 (N_10415,N_10373,N_10215);
nand U10416 (N_10416,N_10226,N_10258);
nand U10417 (N_10417,N_10288,N_10303);
xor U10418 (N_10418,N_10218,N_10270);
nand U10419 (N_10419,N_10231,N_10362);
or U10420 (N_10420,N_10309,N_10329);
nor U10421 (N_10421,N_10252,N_10291);
nor U10422 (N_10422,N_10301,N_10394);
xnor U10423 (N_10423,N_10223,N_10342);
and U10424 (N_10424,N_10333,N_10253);
xnor U10425 (N_10425,N_10241,N_10356);
nor U10426 (N_10426,N_10319,N_10393);
and U10427 (N_10427,N_10287,N_10345);
or U10428 (N_10428,N_10299,N_10322);
nand U10429 (N_10429,N_10315,N_10278);
nor U10430 (N_10430,N_10321,N_10395);
and U10431 (N_10431,N_10366,N_10376);
xnor U10432 (N_10432,N_10351,N_10332);
xnor U10433 (N_10433,N_10380,N_10255);
nor U10434 (N_10434,N_10205,N_10281);
and U10435 (N_10435,N_10324,N_10219);
or U10436 (N_10436,N_10353,N_10227);
nor U10437 (N_10437,N_10314,N_10260);
nand U10438 (N_10438,N_10208,N_10368);
nand U10439 (N_10439,N_10317,N_10282);
nor U10440 (N_10440,N_10310,N_10347);
nand U10441 (N_10441,N_10383,N_10279);
or U10442 (N_10442,N_10236,N_10349);
nor U10443 (N_10443,N_10254,N_10316);
xor U10444 (N_10444,N_10269,N_10247);
or U10445 (N_10445,N_10386,N_10369);
nand U10446 (N_10446,N_10272,N_10354);
nor U10447 (N_10447,N_10297,N_10232);
xor U10448 (N_10448,N_10357,N_10293);
or U10449 (N_10449,N_10256,N_10338);
nand U10450 (N_10450,N_10382,N_10298);
nand U10451 (N_10451,N_10263,N_10305);
nor U10452 (N_10452,N_10370,N_10273);
nand U10453 (N_10453,N_10233,N_10267);
nand U10454 (N_10454,N_10204,N_10385);
xor U10455 (N_10455,N_10350,N_10363);
or U10456 (N_10456,N_10331,N_10304);
and U10457 (N_10457,N_10239,N_10248);
xnor U10458 (N_10458,N_10379,N_10202);
nand U10459 (N_10459,N_10375,N_10245);
nand U10460 (N_10460,N_10203,N_10359);
and U10461 (N_10461,N_10334,N_10339);
xor U10462 (N_10462,N_10399,N_10220);
or U10463 (N_10463,N_10207,N_10200);
or U10464 (N_10464,N_10237,N_10388);
and U10465 (N_10465,N_10230,N_10266);
and U10466 (N_10466,N_10243,N_10367);
xnor U10467 (N_10467,N_10286,N_10327);
xor U10468 (N_10468,N_10323,N_10214);
and U10469 (N_10469,N_10246,N_10312);
nor U10470 (N_10470,N_10336,N_10335);
xor U10471 (N_10471,N_10352,N_10397);
or U10472 (N_10472,N_10392,N_10384);
nor U10473 (N_10473,N_10201,N_10274);
or U10474 (N_10474,N_10242,N_10225);
or U10475 (N_10475,N_10326,N_10216);
and U10476 (N_10476,N_10259,N_10343);
nand U10477 (N_10477,N_10361,N_10371);
and U10478 (N_10478,N_10378,N_10307);
nor U10479 (N_10479,N_10337,N_10234);
and U10480 (N_10480,N_10360,N_10340);
nor U10481 (N_10481,N_10244,N_10390);
xnor U10482 (N_10482,N_10276,N_10222);
nand U10483 (N_10483,N_10275,N_10295);
or U10484 (N_10484,N_10389,N_10320);
or U10485 (N_10485,N_10396,N_10238);
nor U10486 (N_10486,N_10249,N_10213);
and U10487 (N_10487,N_10229,N_10221);
nand U10488 (N_10488,N_10358,N_10217);
xor U10489 (N_10489,N_10250,N_10377);
nor U10490 (N_10490,N_10318,N_10341);
xnor U10491 (N_10491,N_10311,N_10283);
xor U10492 (N_10492,N_10364,N_10381);
or U10493 (N_10493,N_10292,N_10206);
xor U10494 (N_10494,N_10302,N_10262);
nand U10495 (N_10495,N_10257,N_10391);
xor U10496 (N_10496,N_10355,N_10344);
or U10497 (N_10497,N_10289,N_10251);
nand U10498 (N_10498,N_10211,N_10284);
and U10499 (N_10499,N_10224,N_10277);
xor U10500 (N_10500,N_10365,N_10278);
nand U10501 (N_10501,N_10374,N_10247);
nor U10502 (N_10502,N_10368,N_10273);
or U10503 (N_10503,N_10210,N_10315);
nor U10504 (N_10504,N_10209,N_10281);
nand U10505 (N_10505,N_10353,N_10256);
nor U10506 (N_10506,N_10290,N_10216);
and U10507 (N_10507,N_10355,N_10330);
nor U10508 (N_10508,N_10234,N_10235);
nor U10509 (N_10509,N_10372,N_10293);
and U10510 (N_10510,N_10200,N_10283);
or U10511 (N_10511,N_10397,N_10241);
and U10512 (N_10512,N_10381,N_10395);
nor U10513 (N_10513,N_10274,N_10279);
nor U10514 (N_10514,N_10228,N_10363);
or U10515 (N_10515,N_10260,N_10268);
nand U10516 (N_10516,N_10256,N_10369);
and U10517 (N_10517,N_10208,N_10333);
nand U10518 (N_10518,N_10256,N_10313);
nand U10519 (N_10519,N_10230,N_10202);
and U10520 (N_10520,N_10231,N_10370);
xor U10521 (N_10521,N_10387,N_10337);
xor U10522 (N_10522,N_10223,N_10372);
xnor U10523 (N_10523,N_10331,N_10283);
nor U10524 (N_10524,N_10296,N_10232);
nor U10525 (N_10525,N_10268,N_10317);
xnor U10526 (N_10526,N_10285,N_10260);
nor U10527 (N_10527,N_10378,N_10239);
or U10528 (N_10528,N_10321,N_10283);
xor U10529 (N_10529,N_10209,N_10348);
nor U10530 (N_10530,N_10324,N_10375);
nand U10531 (N_10531,N_10267,N_10344);
nand U10532 (N_10532,N_10293,N_10316);
and U10533 (N_10533,N_10255,N_10261);
xor U10534 (N_10534,N_10347,N_10306);
xnor U10535 (N_10535,N_10215,N_10286);
nand U10536 (N_10536,N_10368,N_10205);
nor U10537 (N_10537,N_10204,N_10314);
or U10538 (N_10538,N_10350,N_10301);
xor U10539 (N_10539,N_10367,N_10332);
xor U10540 (N_10540,N_10214,N_10316);
nor U10541 (N_10541,N_10242,N_10319);
nor U10542 (N_10542,N_10227,N_10378);
and U10543 (N_10543,N_10320,N_10350);
and U10544 (N_10544,N_10359,N_10321);
or U10545 (N_10545,N_10341,N_10362);
or U10546 (N_10546,N_10238,N_10333);
or U10547 (N_10547,N_10297,N_10341);
xor U10548 (N_10548,N_10337,N_10248);
and U10549 (N_10549,N_10329,N_10262);
and U10550 (N_10550,N_10325,N_10224);
xor U10551 (N_10551,N_10239,N_10260);
or U10552 (N_10552,N_10349,N_10290);
and U10553 (N_10553,N_10367,N_10249);
nand U10554 (N_10554,N_10381,N_10282);
nor U10555 (N_10555,N_10310,N_10228);
or U10556 (N_10556,N_10205,N_10350);
nor U10557 (N_10557,N_10385,N_10304);
nand U10558 (N_10558,N_10213,N_10323);
nor U10559 (N_10559,N_10352,N_10363);
nand U10560 (N_10560,N_10206,N_10337);
and U10561 (N_10561,N_10288,N_10254);
nor U10562 (N_10562,N_10310,N_10359);
nand U10563 (N_10563,N_10223,N_10247);
nand U10564 (N_10564,N_10289,N_10308);
and U10565 (N_10565,N_10271,N_10280);
nor U10566 (N_10566,N_10234,N_10205);
nor U10567 (N_10567,N_10388,N_10371);
or U10568 (N_10568,N_10262,N_10226);
or U10569 (N_10569,N_10340,N_10363);
or U10570 (N_10570,N_10254,N_10318);
or U10571 (N_10571,N_10336,N_10229);
xnor U10572 (N_10572,N_10244,N_10296);
nand U10573 (N_10573,N_10296,N_10241);
nor U10574 (N_10574,N_10263,N_10313);
nor U10575 (N_10575,N_10317,N_10374);
and U10576 (N_10576,N_10322,N_10256);
xnor U10577 (N_10577,N_10290,N_10321);
nor U10578 (N_10578,N_10381,N_10342);
nor U10579 (N_10579,N_10298,N_10387);
or U10580 (N_10580,N_10233,N_10248);
xnor U10581 (N_10581,N_10248,N_10245);
and U10582 (N_10582,N_10279,N_10241);
and U10583 (N_10583,N_10352,N_10222);
and U10584 (N_10584,N_10212,N_10221);
and U10585 (N_10585,N_10319,N_10320);
and U10586 (N_10586,N_10331,N_10397);
nor U10587 (N_10587,N_10349,N_10281);
or U10588 (N_10588,N_10376,N_10289);
or U10589 (N_10589,N_10351,N_10366);
nand U10590 (N_10590,N_10308,N_10225);
or U10591 (N_10591,N_10244,N_10222);
xor U10592 (N_10592,N_10298,N_10345);
nand U10593 (N_10593,N_10364,N_10304);
xor U10594 (N_10594,N_10333,N_10392);
nor U10595 (N_10595,N_10292,N_10397);
and U10596 (N_10596,N_10231,N_10318);
nor U10597 (N_10597,N_10332,N_10323);
nand U10598 (N_10598,N_10288,N_10236);
nand U10599 (N_10599,N_10314,N_10254);
and U10600 (N_10600,N_10437,N_10436);
xor U10601 (N_10601,N_10550,N_10571);
or U10602 (N_10602,N_10466,N_10499);
nand U10603 (N_10603,N_10524,N_10450);
nand U10604 (N_10604,N_10575,N_10409);
or U10605 (N_10605,N_10465,N_10449);
nor U10606 (N_10606,N_10498,N_10541);
nand U10607 (N_10607,N_10504,N_10461);
nand U10608 (N_10608,N_10472,N_10442);
xnor U10609 (N_10609,N_10425,N_10464);
nand U10610 (N_10610,N_10573,N_10458);
or U10611 (N_10611,N_10510,N_10496);
or U10612 (N_10612,N_10563,N_10518);
xnor U10613 (N_10613,N_10569,N_10444);
xor U10614 (N_10614,N_10511,N_10561);
xor U10615 (N_10615,N_10583,N_10572);
xnor U10616 (N_10616,N_10567,N_10579);
and U10617 (N_10617,N_10570,N_10537);
nor U10618 (N_10618,N_10426,N_10580);
or U10619 (N_10619,N_10482,N_10456);
nor U10620 (N_10620,N_10495,N_10405);
xnor U10621 (N_10621,N_10556,N_10497);
nand U10622 (N_10622,N_10417,N_10544);
nor U10623 (N_10623,N_10508,N_10485);
nand U10624 (N_10624,N_10493,N_10592);
xnor U10625 (N_10625,N_10515,N_10586);
or U10626 (N_10626,N_10527,N_10433);
and U10627 (N_10627,N_10401,N_10462);
nor U10628 (N_10628,N_10529,N_10574);
and U10629 (N_10629,N_10588,N_10419);
nand U10630 (N_10630,N_10438,N_10542);
nand U10631 (N_10631,N_10422,N_10451);
nand U10632 (N_10632,N_10516,N_10483);
nor U10633 (N_10633,N_10589,N_10519);
or U10634 (N_10634,N_10528,N_10596);
xor U10635 (N_10635,N_10407,N_10531);
or U10636 (N_10636,N_10530,N_10502);
nand U10637 (N_10637,N_10512,N_10494);
nand U10638 (N_10638,N_10533,N_10559);
xor U10639 (N_10639,N_10427,N_10525);
and U10640 (N_10640,N_10474,N_10584);
nand U10641 (N_10641,N_10565,N_10413);
nand U10642 (N_10642,N_10539,N_10412);
xnor U10643 (N_10643,N_10546,N_10553);
or U10644 (N_10644,N_10489,N_10507);
nand U10645 (N_10645,N_10501,N_10500);
or U10646 (N_10646,N_10514,N_10414);
nor U10647 (N_10647,N_10562,N_10408);
or U10648 (N_10648,N_10487,N_10471);
nor U10649 (N_10649,N_10446,N_10459);
xor U10650 (N_10650,N_10517,N_10439);
or U10651 (N_10651,N_10420,N_10540);
and U10652 (N_10652,N_10503,N_10490);
and U10653 (N_10653,N_10587,N_10476);
or U10654 (N_10654,N_10416,N_10473);
and U10655 (N_10655,N_10534,N_10448);
nor U10656 (N_10656,N_10453,N_10447);
xnor U10657 (N_10657,N_10430,N_10429);
nor U10658 (N_10658,N_10479,N_10481);
or U10659 (N_10659,N_10566,N_10468);
or U10660 (N_10660,N_10411,N_10576);
and U10661 (N_10661,N_10526,N_10492);
nand U10662 (N_10662,N_10421,N_10467);
nand U10663 (N_10663,N_10591,N_10547);
nand U10664 (N_10664,N_10597,N_10478);
and U10665 (N_10665,N_10470,N_10406);
nor U10666 (N_10666,N_10554,N_10548);
nand U10667 (N_10667,N_10577,N_10509);
xnor U10668 (N_10668,N_10488,N_10404);
or U10669 (N_10669,N_10545,N_10480);
and U10670 (N_10670,N_10506,N_10555);
and U10671 (N_10671,N_10560,N_10428);
and U10672 (N_10672,N_10423,N_10536);
nor U10673 (N_10673,N_10403,N_10424);
or U10674 (N_10674,N_10477,N_10558);
nor U10675 (N_10675,N_10418,N_10469);
nand U10676 (N_10676,N_10457,N_10486);
nand U10677 (N_10677,N_10475,N_10452);
xnor U10678 (N_10678,N_10593,N_10443);
or U10679 (N_10679,N_10400,N_10538);
xor U10680 (N_10680,N_10460,N_10505);
xnor U10681 (N_10681,N_10513,N_10582);
xnor U10682 (N_10682,N_10521,N_10595);
nor U10683 (N_10683,N_10520,N_10578);
xnor U10684 (N_10684,N_10549,N_10410);
or U10685 (N_10685,N_10491,N_10434);
or U10686 (N_10686,N_10440,N_10598);
or U10687 (N_10687,N_10535,N_10532);
and U10688 (N_10688,N_10435,N_10543);
or U10689 (N_10689,N_10402,N_10581);
nor U10690 (N_10690,N_10523,N_10568);
xnor U10691 (N_10691,N_10415,N_10454);
nor U10692 (N_10692,N_10431,N_10594);
or U10693 (N_10693,N_10590,N_10484);
nand U10694 (N_10694,N_10463,N_10522);
xor U10695 (N_10695,N_10564,N_10455);
or U10696 (N_10696,N_10551,N_10432);
nand U10697 (N_10697,N_10441,N_10445);
xnor U10698 (N_10698,N_10557,N_10552);
or U10699 (N_10699,N_10585,N_10599);
and U10700 (N_10700,N_10477,N_10567);
xor U10701 (N_10701,N_10432,N_10526);
xnor U10702 (N_10702,N_10454,N_10579);
nor U10703 (N_10703,N_10410,N_10401);
or U10704 (N_10704,N_10405,N_10433);
nand U10705 (N_10705,N_10489,N_10460);
or U10706 (N_10706,N_10593,N_10407);
or U10707 (N_10707,N_10483,N_10436);
xnor U10708 (N_10708,N_10408,N_10527);
nor U10709 (N_10709,N_10487,N_10429);
xnor U10710 (N_10710,N_10555,N_10574);
and U10711 (N_10711,N_10499,N_10425);
or U10712 (N_10712,N_10580,N_10531);
and U10713 (N_10713,N_10439,N_10549);
and U10714 (N_10714,N_10513,N_10480);
xnor U10715 (N_10715,N_10520,N_10510);
or U10716 (N_10716,N_10486,N_10410);
and U10717 (N_10717,N_10533,N_10405);
or U10718 (N_10718,N_10504,N_10580);
or U10719 (N_10719,N_10464,N_10548);
xnor U10720 (N_10720,N_10437,N_10468);
nor U10721 (N_10721,N_10577,N_10540);
or U10722 (N_10722,N_10599,N_10528);
nand U10723 (N_10723,N_10577,N_10534);
xor U10724 (N_10724,N_10567,N_10544);
and U10725 (N_10725,N_10518,N_10469);
nor U10726 (N_10726,N_10485,N_10446);
xnor U10727 (N_10727,N_10465,N_10488);
and U10728 (N_10728,N_10556,N_10486);
and U10729 (N_10729,N_10467,N_10506);
nand U10730 (N_10730,N_10543,N_10571);
nor U10731 (N_10731,N_10524,N_10506);
nor U10732 (N_10732,N_10425,N_10543);
and U10733 (N_10733,N_10427,N_10532);
nor U10734 (N_10734,N_10580,N_10539);
nand U10735 (N_10735,N_10580,N_10485);
or U10736 (N_10736,N_10566,N_10537);
nand U10737 (N_10737,N_10594,N_10406);
and U10738 (N_10738,N_10541,N_10474);
nor U10739 (N_10739,N_10588,N_10488);
nor U10740 (N_10740,N_10557,N_10520);
and U10741 (N_10741,N_10453,N_10555);
xor U10742 (N_10742,N_10577,N_10532);
and U10743 (N_10743,N_10429,N_10563);
or U10744 (N_10744,N_10461,N_10489);
nand U10745 (N_10745,N_10598,N_10560);
nand U10746 (N_10746,N_10444,N_10475);
nand U10747 (N_10747,N_10568,N_10541);
nor U10748 (N_10748,N_10563,N_10473);
and U10749 (N_10749,N_10433,N_10457);
xnor U10750 (N_10750,N_10422,N_10454);
and U10751 (N_10751,N_10491,N_10480);
nand U10752 (N_10752,N_10420,N_10533);
nor U10753 (N_10753,N_10578,N_10558);
nand U10754 (N_10754,N_10437,N_10464);
and U10755 (N_10755,N_10521,N_10423);
nor U10756 (N_10756,N_10475,N_10514);
xor U10757 (N_10757,N_10520,N_10508);
or U10758 (N_10758,N_10418,N_10494);
xor U10759 (N_10759,N_10460,N_10529);
nand U10760 (N_10760,N_10475,N_10563);
or U10761 (N_10761,N_10550,N_10489);
or U10762 (N_10762,N_10526,N_10487);
and U10763 (N_10763,N_10529,N_10415);
and U10764 (N_10764,N_10463,N_10555);
or U10765 (N_10765,N_10478,N_10411);
nor U10766 (N_10766,N_10463,N_10565);
xnor U10767 (N_10767,N_10527,N_10466);
nand U10768 (N_10768,N_10566,N_10575);
or U10769 (N_10769,N_10437,N_10500);
and U10770 (N_10770,N_10530,N_10565);
nor U10771 (N_10771,N_10455,N_10523);
and U10772 (N_10772,N_10580,N_10560);
nand U10773 (N_10773,N_10586,N_10476);
nor U10774 (N_10774,N_10587,N_10538);
nor U10775 (N_10775,N_10436,N_10448);
nand U10776 (N_10776,N_10500,N_10516);
and U10777 (N_10777,N_10505,N_10587);
xnor U10778 (N_10778,N_10416,N_10483);
xnor U10779 (N_10779,N_10496,N_10482);
or U10780 (N_10780,N_10523,N_10520);
nand U10781 (N_10781,N_10433,N_10458);
xnor U10782 (N_10782,N_10450,N_10597);
nand U10783 (N_10783,N_10448,N_10407);
or U10784 (N_10784,N_10513,N_10552);
nand U10785 (N_10785,N_10433,N_10475);
or U10786 (N_10786,N_10477,N_10416);
xnor U10787 (N_10787,N_10440,N_10509);
xnor U10788 (N_10788,N_10559,N_10567);
and U10789 (N_10789,N_10544,N_10515);
nand U10790 (N_10790,N_10410,N_10474);
or U10791 (N_10791,N_10488,N_10494);
or U10792 (N_10792,N_10473,N_10515);
nand U10793 (N_10793,N_10508,N_10424);
or U10794 (N_10794,N_10473,N_10495);
nand U10795 (N_10795,N_10591,N_10555);
or U10796 (N_10796,N_10563,N_10446);
and U10797 (N_10797,N_10574,N_10548);
nand U10798 (N_10798,N_10502,N_10477);
and U10799 (N_10799,N_10482,N_10410);
or U10800 (N_10800,N_10634,N_10641);
or U10801 (N_10801,N_10704,N_10678);
nand U10802 (N_10802,N_10688,N_10728);
xnor U10803 (N_10803,N_10789,N_10772);
nor U10804 (N_10804,N_10647,N_10787);
nand U10805 (N_10805,N_10726,N_10783);
xor U10806 (N_10806,N_10636,N_10627);
nand U10807 (N_10807,N_10645,N_10701);
nor U10808 (N_10808,N_10680,N_10664);
nand U10809 (N_10809,N_10775,N_10697);
nand U10810 (N_10810,N_10747,N_10796);
nor U10811 (N_10811,N_10718,N_10719);
nor U10812 (N_10812,N_10721,N_10785);
nor U10813 (N_10813,N_10668,N_10742);
xnor U10814 (N_10814,N_10629,N_10607);
nor U10815 (N_10815,N_10705,N_10687);
nor U10816 (N_10816,N_10694,N_10649);
or U10817 (N_10817,N_10610,N_10652);
nand U10818 (N_10818,N_10755,N_10600);
or U10819 (N_10819,N_10765,N_10767);
nand U10820 (N_10820,N_10630,N_10727);
xor U10821 (N_10821,N_10637,N_10738);
and U10822 (N_10822,N_10653,N_10656);
nand U10823 (N_10823,N_10773,N_10735);
nor U10824 (N_10824,N_10703,N_10615);
nor U10825 (N_10825,N_10609,N_10716);
xnor U10826 (N_10826,N_10679,N_10768);
xor U10827 (N_10827,N_10715,N_10675);
nor U10828 (N_10828,N_10608,N_10628);
nor U10829 (N_10829,N_10640,N_10739);
nor U10830 (N_10830,N_10794,N_10695);
nor U10831 (N_10831,N_10717,N_10760);
and U10832 (N_10832,N_10706,N_10691);
nor U10833 (N_10833,N_10696,N_10766);
xor U10834 (N_10834,N_10731,N_10776);
nor U10835 (N_10835,N_10677,N_10603);
or U10836 (N_10836,N_10606,N_10746);
nor U10837 (N_10837,N_10780,N_10611);
or U10838 (N_10838,N_10722,N_10799);
and U10839 (N_10839,N_10622,N_10661);
or U10840 (N_10840,N_10782,N_10779);
nand U10841 (N_10841,N_10674,N_10660);
and U10842 (N_10842,N_10756,N_10659);
nor U10843 (N_10843,N_10620,N_10777);
nand U10844 (N_10844,N_10693,N_10672);
xor U10845 (N_10845,N_10748,N_10751);
nand U10846 (N_10846,N_10792,N_10788);
nor U10847 (N_10847,N_10708,N_10725);
nand U10848 (N_10848,N_10761,N_10650);
xnor U10849 (N_10849,N_10778,N_10663);
or U10850 (N_10850,N_10790,N_10713);
nand U10851 (N_10851,N_10774,N_10723);
xnor U10852 (N_10852,N_10605,N_10654);
nand U10853 (N_10853,N_10784,N_10741);
and U10854 (N_10854,N_10681,N_10651);
nand U10855 (N_10855,N_10632,N_10714);
xnor U10856 (N_10856,N_10740,N_10724);
xor U10857 (N_10857,N_10631,N_10757);
nor U10858 (N_10858,N_10643,N_10657);
xor U10859 (N_10859,N_10710,N_10683);
nor U10860 (N_10860,N_10754,N_10621);
or U10861 (N_10861,N_10662,N_10689);
and U10862 (N_10862,N_10639,N_10638);
nor U10863 (N_10863,N_10749,N_10769);
xor U10864 (N_10864,N_10646,N_10730);
xor U10865 (N_10865,N_10682,N_10762);
or U10866 (N_10866,N_10644,N_10711);
and U10867 (N_10867,N_10658,N_10625);
or U10868 (N_10868,N_10617,N_10759);
or U10869 (N_10869,N_10729,N_10752);
nor U10870 (N_10870,N_10795,N_10737);
or U10871 (N_10871,N_10763,N_10791);
xor U10872 (N_10872,N_10684,N_10770);
and U10873 (N_10873,N_10758,N_10793);
xor U10874 (N_10874,N_10702,N_10619);
nand U10875 (N_10875,N_10601,N_10750);
and U10876 (N_10876,N_10602,N_10786);
nand U10877 (N_10877,N_10753,N_10736);
and U10878 (N_10878,N_10616,N_10642);
or U10879 (N_10879,N_10692,N_10699);
xor U10880 (N_10880,N_10734,N_10670);
or U10881 (N_10881,N_10612,N_10667);
nand U10882 (N_10882,N_10733,N_10732);
or U10883 (N_10883,N_10624,N_10676);
xor U10884 (N_10884,N_10709,N_10613);
nand U10885 (N_10885,N_10781,N_10686);
and U10886 (N_10886,N_10614,N_10626);
and U10887 (N_10887,N_10744,N_10764);
nand U10888 (N_10888,N_10623,N_10633);
nor U10889 (N_10889,N_10666,N_10685);
or U10890 (N_10890,N_10798,N_10771);
xnor U10891 (N_10891,N_10707,N_10669);
and U10892 (N_10892,N_10720,N_10690);
nand U10893 (N_10893,N_10655,N_10673);
nor U10894 (N_10894,N_10665,N_10671);
nand U10895 (N_10895,N_10797,N_10743);
nor U10896 (N_10896,N_10618,N_10604);
nand U10897 (N_10897,N_10712,N_10700);
xor U10898 (N_10898,N_10745,N_10698);
and U10899 (N_10899,N_10635,N_10648);
nand U10900 (N_10900,N_10714,N_10621);
or U10901 (N_10901,N_10664,N_10765);
and U10902 (N_10902,N_10689,N_10604);
nor U10903 (N_10903,N_10701,N_10654);
xor U10904 (N_10904,N_10699,N_10729);
nand U10905 (N_10905,N_10777,N_10639);
xor U10906 (N_10906,N_10628,N_10784);
nand U10907 (N_10907,N_10771,N_10698);
nor U10908 (N_10908,N_10643,N_10616);
nor U10909 (N_10909,N_10618,N_10799);
and U10910 (N_10910,N_10758,N_10662);
or U10911 (N_10911,N_10670,N_10716);
and U10912 (N_10912,N_10606,N_10644);
nor U10913 (N_10913,N_10762,N_10658);
xor U10914 (N_10914,N_10750,N_10611);
and U10915 (N_10915,N_10688,N_10742);
nand U10916 (N_10916,N_10636,N_10616);
xor U10917 (N_10917,N_10644,N_10742);
xnor U10918 (N_10918,N_10684,N_10652);
or U10919 (N_10919,N_10673,N_10638);
or U10920 (N_10920,N_10682,N_10701);
xnor U10921 (N_10921,N_10718,N_10775);
xor U10922 (N_10922,N_10612,N_10732);
nand U10923 (N_10923,N_10672,N_10600);
nor U10924 (N_10924,N_10642,N_10617);
nand U10925 (N_10925,N_10756,N_10762);
nor U10926 (N_10926,N_10606,N_10610);
or U10927 (N_10927,N_10709,N_10668);
nand U10928 (N_10928,N_10605,N_10602);
and U10929 (N_10929,N_10668,N_10616);
xnor U10930 (N_10930,N_10721,N_10681);
nand U10931 (N_10931,N_10623,N_10651);
xor U10932 (N_10932,N_10706,N_10747);
nand U10933 (N_10933,N_10690,N_10714);
xor U10934 (N_10934,N_10646,N_10700);
nor U10935 (N_10935,N_10605,N_10747);
or U10936 (N_10936,N_10795,N_10716);
or U10937 (N_10937,N_10714,N_10654);
and U10938 (N_10938,N_10765,N_10747);
nor U10939 (N_10939,N_10728,N_10709);
and U10940 (N_10940,N_10616,N_10681);
nand U10941 (N_10941,N_10698,N_10657);
nor U10942 (N_10942,N_10714,N_10694);
or U10943 (N_10943,N_10689,N_10618);
and U10944 (N_10944,N_10640,N_10747);
nand U10945 (N_10945,N_10789,N_10788);
nor U10946 (N_10946,N_10609,N_10746);
and U10947 (N_10947,N_10747,N_10733);
nor U10948 (N_10948,N_10634,N_10785);
xor U10949 (N_10949,N_10774,N_10737);
nand U10950 (N_10950,N_10617,N_10644);
and U10951 (N_10951,N_10722,N_10691);
and U10952 (N_10952,N_10694,N_10782);
xor U10953 (N_10953,N_10794,N_10633);
and U10954 (N_10954,N_10734,N_10773);
nand U10955 (N_10955,N_10602,N_10641);
nor U10956 (N_10956,N_10699,N_10784);
and U10957 (N_10957,N_10637,N_10645);
or U10958 (N_10958,N_10670,N_10691);
xor U10959 (N_10959,N_10671,N_10786);
nor U10960 (N_10960,N_10704,N_10657);
nor U10961 (N_10961,N_10694,N_10686);
or U10962 (N_10962,N_10761,N_10769);
nand U10963 (N_10963,N_10636,N_10767);
and U10964 (N_10964,N_10668,N_10630);
xnor U10965 (N_10965,N_10674,N_10646);
or U10966 (N_10966,N_10700,N_10709);
or U10967 (N_10967,N_10715,N_10669);
xor U10968 (N_10968,N_10730,N_10765);
xor U10969 (N_10969,N_10684,N_10610);
xnor U10970 (N_10970,N_10638,N_10681);
or U10971 (N_10971,N_10600,N_10703);
or U10972 (N_10972,N_10795,N_10609);
nor U10973 (N_10973,N_10693,N_10641);
nor U10974 (N_10974,N_10759,N_10692);
and U10975 (N_10975,N_10682,N_10725);
nor U10976 (N_10976,N_10761,N_10731);
nor U10977 (N_10977,N_10742,N_10672);
or U10978 (N_10978,N_10669,N_10639);
nor U10979 (N_10979,N_10716,N_10686);
and U10980 (N_10980,N_10702,N_10792);
and U10981 (N_10981,N_10701,N_10737);
or U10982 (N_10982,N_10716,N_10705);
xnor U10983 (N_10983,N_10602,N_10644);
or U10984 (N_10984,N_10792,N_10766);
nor U10985 (N_10985,N_10788,N_10746);
nor U10986 (N_10986,N_10623,N_10698);
or U10987 (N_10987,N_10708,N_10659);
nor U10988 (N_10988,N_10678,N_10710);
nor U10989 (N_10989,N_10686,N_10641);
and U10990 (N_10990,N_10635,N_10616);
and U10991 (N_10991,N_10617,N_10755);
nand U10992 (N_10992,N_10643,N_10788);
xor U10993 (N_10993,N_10630,N_10676);
nor U10994 (N_10994,N_10751,N_10757);
or U10995 (N_10995,N_10675,N_10724);
nand U10996 (N_10996,N_10793,N_10691);
and U10997 (N_10997,N_10714,N_10727);
nand U10998 (N_10998,N_10684,N_10741);
nand U10999 (N_10999,N_10631,N_10660);
nand U11000 (N_11000,N_10862,N_10835);
nand U11001 (N_11001,N_10806,N_10879);
xor U11002 (N_11002,N_10824,N_10864);
xor U11003 (N_11003,N_10929,N_10966);
or U11004 (N_11004,N_10845,N_10922);
nand U11005 (N_11005,N_10906,N_10938);
xor U11006 (N_11006,N_10855,N_10858);
and U11007 (N_11007,N_10836,N_10869);
nand U11008 (N_11008,N_10890,N_10829);
or U11009 (N_11009,N_10988,N_10943);
or U11010 (N_11010,N_10942,N_10956);
and U11011 (N_11011,N_10838,N_10860);
nand U11012 (N_11012,N_10971,N_10908);
and U11013 (N_11013,N_10953,N_10861);
xor U11014 (N_11014,N_10833,N_10877);
xor U11015 (N_11015,N_10904,N_10818);
nand U11016 (N_11016,N_10882,N_10949);
and U11017 (N_11017,N_10808,N_10989);
or U11018 (N_11018,N_10910,N_10962);
nand U11019 (N_11019,N_10987,N_10873);
nand U11020 (N_11020,N_10940,N_10967);
nand U11021 (N_11021,N_10853,N_10802);
nor U11022 (N_11022,N_10895,N_10856);
and U11023 (N_11023,N_10918,N_10871);
or U11024 (N_11024,N_10839,N_10897);
nand U11025 (N_11025,N_10933,N_10841);
nor U11026 (N_11026,N_10800,N_10955);
and U11027 (N_11027,N_10954,N_10983);
and U11028 (N_11028,N_10960,N_10843);
nor U11029 (N_11029,N_10851,N_10916);
nand U11030 (N_11030,N_10848,N_10857);
nor U11031 (N_11031,N_10973,N_10867);
nand U11032 (N_11032,N_10982,N_10849);
nand U11033 (N_11033,N_10951,N_10801);
or U11034 (N_11034,N_10868,N_10875);
nand U11035 (N_11035,N_10957,N_10844);
nand U11036 (N_11036,N_10821,N_10985);
nor U11037 (N_11037,N_10899,N_10902);
nand U11038 (N_11038,N_10930,N_10993);
and U11039 (N_11039,N_10823,N_10827);
and U11040 (N_11040,N_10850,N_10837);
and U11041 (N_11041,N_10925,N_10874);
nor U11042 (N_11042,N_10979,N_10996);
xnor U11043 (N_11043,N_10932,N_10820);
xnor U11044 (N_11044,N_10923,N_10921);
nor U11045 (N_11045,N_10950,N_10936);
xor U11046 (N_11046,N_10815,N_10990);
and U11047 (N_11047,N_10900,N_10822);
and U11048 (N_11048,N_10984,N_10852);
xnor U11049 (N_11049,N_10881,N_10944);
or U11050 (N_11050,N_10927,N_10919);
or U11051 (N_11051,N_10961,N_10937);
and U11052 (N_11052,N_10924,N_10969);
and U11053 (N_11053,N_10978,N_10813);
xnor U11054 (N_11054,N_10870,N_10888);
nand U11055 (N_11055,N_10935,N_10998);
and U11056 (N_11056,N_10830,N_10828);
nor U11057 (N_11057,N_10886,N_10941);
nor U11058 (N_11058,N_10804,N_10959);
and U11059 (N_11059,N_10885,N_10872);
xnor U11060 (N_11060,N_10903,N_10958);
nand U11061 (N_11061,N_10816,N_10894);
and U11062 (N_11062,N_10840,N_10939);
nor U11063 (N_11063,N_10970,N_10934);
nor U11064 (N_11064,N_10901,N_10952);
xnor U11065 (N_11065,N_10847,N_10999);
xor U11066 (N_11066,N_10814,N_10909);
or U11067 (N_11067,N_10963,N_10965);
xor U11068 (N_11068,N_10883,N_10807);
xor U11069 (N_11069,N_10891,N_10994);
xor U11070 (N_11070,N_10896,N_10878);
nand U11071 (N_11071,N_10810,N_10995);
nor U11072 (N_11072,N_10831,N_10905);
xor U11073 (N_11073,N_10948,N_10842);
or U11074 (N_11074,N_10884,N_10915);
xor U11075 (N_11075,N_10825,N_10803);
nor U11076 (N_11076,N_10859,N_10834);
and U11077 (N_11077,N_10887,N_10972);
nand U11078 (N_11078,N_10968,N_10991);
xor U11079 (N_11079,N_10880,N_10892);
nand U11080 (N_11080,N_10876,N_10974);
nand U11081 (N_11081,N_10912,N_10889);
nand U11082 (N_11082,N_10866,N_10946);
nand U11083 (N_11083,N_10914,N_10964);
nand U11084 (N_11084,N_10854,N_10812);
nand U11085 (N_11085,N_10931,N_10917);
nand U11086 (N_11086,N_10826,N_10846);
and U11087 (N_11087,N_10832,N_10986);
nor U11088 (N_11088,N_10819,N_10947);
nor U11089 (N_11089,N_10913,N_10976);
and U11090 (N_11090,N_10975,N_10863);
nor U11091 (N_11091,N_10980,N_10865);
or U11092 (N_11092,N_10928,N_10809);
nand U11093 (N_11093,N_10997,N_10805);
and U11094 (N_11094,N_10977,N_10911);
or U11095 (N_11095,N_10893,N_10981);
nor U11096 (N_11096,N_10811,N_10920);
xnor U11097 (N_11097,N_10898,N_10907);
nand U11098 (N_11098,N_10926,N_10992);
or U11099 (N_11099,N_10817,N_10945);
xnor U11100 (N_11100,N_10987,N_10816);
nor U11101 (N_11101,N_10868,N_10998);
nand U11102 (N_11102,N_10916,N_10850);
or U11103 (N_11103,N_10889,N_10994);
nand U11104 (N_11104,N_10841,N_10897);
and U11105 (N_11105,N_10991,N_10945);
nand U11106 (N_11106,N_10954,N_10933);
xor U11107 (N_11107,N_10870,N_10967);
xnor U11108 (N_11108,N_10887,N_10843);
nand U11109 (N_11109,N_10890,N_10816);
or U11110 (N_11110,N_10873,N_10812);
xor U11111 (N_11111,N_10876,N_10951);
nand U11112 (N_11112,N_10860,N_10870);
nand U11113 (N_11113,N_10808,N_10926);
nand U11114 (N_11114,N_10984,N_10816);
nand U11115 (N_11115,N_10843,N_10813);
xnor U11116 (N_11116,N_10867,N_10958);
or U11117 (N_11117,N_10815,N_10963);
nand U11118 (N_11118,N_10878,N_10904);
xnor U11119 (N_11119,N_10923,N_10895);
nor U11120 (N_11120,N_10960,N_10982);
or U11121 (N_11121,N_10968,N_10949);
and U11122 (N_11122,N_10899,N_10805);
xnor U11123 (N_11123,N_10982,N_10892);
xnor U11124 (N_11124,N_10904,N_10955);
nand U11125 (N_11125,N_10934,N_10965);
nand U11126 (N_11126,N_10808,N_10896);
xor U11127 (N_11127,N_10973,N_10950);
and U11128 (N_11128,N_10998,N_10833);
nor U11129 (N_11129,N_10869,N_10984);
nor U11130 (N_11130,N_10854,N_10906);
or U11131 (N_11131,N_10814,N_10806);
xor U11132 (N_11132,N_10984,N_10886);
xor U11133 (N_11133,N_10890,N_10878);
nand U11134 (N_11134,N_10871,N_10973);
nor U11135 (N_11135,N_10848,N_10804);
nand U11136 (N_11136,N_10910,N_10860);
xor U11137 (N_11137,N_10852,N_10822);
or U11138 (N_11138,N_10869,N_10982);
xnor U11139 (N_11139,N_10938,N_10883);
nor U11140 (N_11140,N_10872,N_10947);
nand U11141 (N_11141,N_10922,N_10909);
nand U11142 (N_11142,N_10808,N_10890);
or U11143 (N_11143,N_10861,N_10814);
xor U11144 (N_11144,N_10826,N_10894);
and U11145 (N_11145,N_10914,N_10845);
and U11146 (N_11146,N_10880,N_10903);
xor U11147 (N_11147,N_10841,N_10871);
and U11148 (N_11148,N_10854,N_10867);
nor U11149 (N_11149,N_10998,N_10829);
nor U11150 (N_11150,N_10817,N_10935);
nor U11151 (N_11151,N_10957,N_10885);
and U11152 (N_11152,N_10961,N_10909);
and U11153 (N_11153,N_10891,N_10829);
xnor U11154 (N_11154,N_10924,N_10917);
or U11155 (N_11155,N_10858,N_10947);
and U11156 (N_11156,N_10896,N_10850);
xnor U11157 (N_11157,N_10897,N_10935);
xor U11158 (N_11158,N_10892,N_10861);
nand U11159 (N_11159,N_10965,N_10808);
nand U11160 (N_11160,N_10999,N_10980);
nand U11161 (N_11161,N_10892,N_10857);
or U11162 (N_11162,N_10815,N_10950);
and U11163 (N_11163,N_10989,N_10838);
xor U11164 (N_11164,N_10975,N_10895);
nand U11165 (N_11165,N_10882,N_10893);
nand U11166 (N_11166,N_10856,N_10965);
xor U11167 (N_11167,N_10953,N_10844);
and U11168 (N_11168,N_10949,N_10950);
nor U11169 (N_11169,N_10996,N_10806);
nand U11170 (N_11170,N_10817,N_10882);
xor U11171 (N_11171,N_10873,N_10932);
nand U11172 (N_11172,N_10826,N_10963);
or U11173 (N_11173,N_10938,N_10956);
or U11174 (N_11174,N_10817,N_10913);
nor U11175 (N_11175,N_10957,N_10894);
and U11176 (N_11176,N_10870,N_10975);
nand U11177 (N_11177,N_10815,N_10885);
nor U11178 (N_11178,N_10843,N_10953);
or U11179 (N_11179,N_10859,N_10943);
nor U11180 (N_11180,N_10949,N_10985);
or U11181 (N_11181,N_10856,N_10867);
xnor U11182 (N_11182,N_10956,N_10989);
xor U11183 (N_11183,N_10813,N_10873);
xor U11184 (N_11184,N_10947,N_10994);
and U11185 (N_11185,N_10859,N_10914);
or U11186 (N_11186,N_10824,N_10812);
and U11187 (N_11187,N_10948,N_10916);
xor U11188 (N_11188,N_10966,N_10829);
and U11189 (N_11189,N_10812,N_10850);
nor U11190 (N_11190,N_10946,N_10889);
and U11191 (N_11191,N_10850,N_10929);
or U11192 (N_11192,N_10824,N_10894);
or U11193 (N_11193,N_10873,N_10887);
xnor U11194 (N_11194,N_10847,N_10929);
and U11195 (N_11195,N_10967,N_10864);
nand U11196 (N_11196,N_10931,N_10830);
xnor U11197 (N_11197,N_10824,N_10907);
nand U11198 (N_11198,N_10894,N_10906);
nand U11199 (N_11199,N_10843,N_10982);
nor U11200 (N_11200,N_11180,N_11075);
or U11201 (N_11201,N_11020,N_11029);
nor U11202 (N_11202,N_11090,N_11087);
or U11203 (N_11203,N_11153,N_11164);
nor U11204 (N_11204,N_11152,N_11141);
or U11205 (N_11205,N_11139,N_11154);
nor U11206 (N_11206,N_11144,N_11148);
or U11207 (N_11207,N_11138,N_11042);
and U11208 (N_11208,N_11110,N_11074);
nor U11209 (N_11209,N_11078,N_11050);
and U11210 (N_11210,N_11175,N_11051);
and U11211 (N_11211,N_11168,N_11098);
and U11212 (N_11212,N_11105,N_11004);
and U11213 (N_11213,N_11072,N_11140);
xnor U11214 (N_11214,N_11032,N_11162);
and U11215 (N_11215,N_11066,N_11116);
nor U11216 (N_11216,N_11089,N_11189);
nand U11217 (N_11217,N_11000,N_11045);
nor U11218 (N_11218,N_11161,N_11080);
xnor U11219 (N_11219,N_11177,N_11195);
and U11220 (N_11220,N_11060,N_11117);
nand U11221 (N_11221,N_11064,N_11120);
nand U11222 (N_11222,N_11037,N_11002);
nor U11223 (N_11223,N_11113,N_11132);
nor U11224 (N_11224,N_11021,N_11068);
and U11225 (N_11225,N_11142,N_11058);
nand U11226 (N_11226,N_11143,N_11077);
or U11227 (N_11227,N_11149,N_11019);
nor U11228 (N_11228,N_11088,N_11026);
nand U11229 (N_11229,N_11010,N_11119);
nor U11230 (N_11230,N_11191,N_11056);
nand U11231 (N_11231,N_11016,N_11012);
and U11232 (N_11232,N_11003,N_11197);
nor U11233 (N_11233,N_11055,N_11150);
or U11234 (N_11234,N_11025,N_11147);
nand U11235 (N_11235,N_11178,N_11100);
and U11236 (N_11236,N_11085,N_11052);
xor U11237 (N_11237,N_11107,N_11157);
and U11238 (N_11238,N_11190,N_11108);
nor U11239 (N_11239,N_11038,N_11170);
and U11240 (N_11240,N_11165,N_11093);
or U11241 (N_11241,N_11167,N_11023);
or U11242 (N_11242,N_11122,N_11131);
and U11243 (N_11243,N_11008,N_11070);
xor U11244 (N_11244,N_11181,N_11047);
or U11245 (N_11245,N_11159,N_11151);
nand U11246 (N_11246,N_11076,N_11194);
or U11247 (N_11247,N_11043,N_11035);
xnor U11248 (N_11248,N_11104,N_11171);
xor U11249 (N_11249,N_11134,N_11028);
or U11250 (N_11250,N_11083,N_11185);
nor U11251 (N_11251,N_11014,N_11015);
xor U11252 (N_11252,N_11095,N_11166);
or U11253 (N_11253,N_11124,N_11099);
xnor U11254 (N_11254,N_11086,N_11091);
and U11255 (N_11255,N_11173,N_11183);
nand U11256 (N_11256,N_11174,N_11033);
nand U11257 (N_11257,N_11053,N_11102);
xor U11258 (N_11258,N_11188,N_11041);
xnor U11259 (N_11259,N_11094,N_11017);
nand U11260 (N_11260,N_11186,N_11057);
xnor U11261 (N_11261,N_11160,N_11184);
nor U11262 (N_11262,N_11063,N_11169);
nor U11263 (N_11263,N_11081,N_11109);
or U11264 (N_11264,N_11062,N_11069);
nor U11265 (N_11265,N_11011,N_11048);
nand U11266 (N_11266,N_11137,N_11193);
and U11267 (N_11267,N_11106,N_11018);
and U11268 (N_11268,N_11061,N_11133);
or U11269 (N_11269,N_11067,N_11046);
or U11270 (N_11270,N_11158,N_11125);
and U11271 (N_11271,N_11082,N_11036);
and U11272 (N_11272,N_11027,N_11049);
nor U11273 (N_11273,N_11129,N_11155);
and U11274 (N_11274,N_11039,N_11044);
nor U11275 (N_11275,N_11092,N_11146);
or U11276 (N_11276,N_11040,N_11007);
xnor U11277 (N_11277,N_11054,N_11006);
nand U11278 (N_11278,N_11121,N_11156);
or U11279 (N_11279,N_11084,N_11071);
nand U11280 (N_11280,N_11198,N_11172);
nor U11281 (N_11281,N_11013,N_11024);
xor U11282 (N_11282,N_11127,N_11136);
xnor U11283 (N_11283,N_11079,N_11135);
or U11284 (N_11284,N_11128,N_11065);
and U11285 (N_11285,N_11114,N_11130);
nor U11286 (N_11286,N_11022,N_11176);
or U11287 (N_11287,N_11103,N_11192);
or U11288 (N_11288,N_11030,N_11115);
or U11289 (N_11289,N_11145,N_11199);
or U11290 (N_11290,N_11112,N_11126);
xnor U11291 (N_11291,N_11163,N_11059);
and U11292 (N_11292,N_11123,N_11196);
nor U11293 (N_11293,N_11111,N_11031);
and U11294 (N_11294,N_11187,N_11001);
and U11295 (N_11295,N_11118,N_11096);
xnor U11296 (N_11296,N_11073,N_11179);
and U11297 (N_11297,N_11005,N_11034);
nor U11298 (N_11298,N_11097,N_11182);
nor U11299 (N_11299,N_11101,N_11009);
xnor U11300 (N_11300,N_11160,N_11070);
nor U11301 (N_11301,N_11085,N_11194);
xnor U11302 (N_11302,N_11062,N_11162);
and U11303 (N_11303,N_11177,N_11164);
xor U11304 (N_11304,N_11083,N_11072);
nor U11305 (N_11305,N_11088,N_11131);
or U11306 (N_11306,N_11039,N_11049);
nand U11307 (N_11307,N_11021,N_11023);
nor U11308 (N_11308,N_11003,N_11085);
or U11309 (N_11309,N_11161,N_11064);
and U11310 (N_11310,N_11105,N_11112);
nand U11311 (N_11311,N_11127,N_11199);
or U11312 (N_11312,N_11077,N_11046);
or U11313 (N_11313,N_11010,N_11075);
and U11314 (N_11314,N_11012,N_11116);
nor U11315 (N_11315,N_11102,N_11172);
nor U11316 (N_11316,N_11032,N_11078);
or U11317 (N_11317,N_11138,N_11081);
nor U11318 (N_11318,N_11043,N_11105);
and U11319 (N_11319,N_11111,N_11008);
and U11320 (N_11320,N_11076,N_11135);
xnor U11321 (N_11321,N_11097,N_11173);
nand U11322 (N_11322,N_11087,N_11065);
or U11323 (N_11323,N_11111,N_11011);
and U11324 (N_11324,N_11004,N_11051);
and U11325 (N_11325,N_11133,N_11125);
xnor U11326 (N_11326,N_11134,N_11075);
nand U11327 (N_11327,N_11063,N_11155);
or U11328 (N_11328,N_11038,N_11082);
or U11329 (N_11329,N_11013,N_11186);
nor U11330 (N_11330,N_11171,N_11110);
nor U11331 (N_11331,N_11083,N_11170);
or U11332 (N_11332,N_11135,N_11095);
xor U11333 (N_11333,N_11078,N_11052);
xor U11334 (N_11334,N_11026,N_11073);
and U11335 (N_11335,N_11159,N_11105);
nand U11336 (N_11336,N_11178,N_11035);
nand U11337 (N_11337,N_11109,N_11052);
and U11338 (N_11338,N_11099,N_11046);
and U11339 (N_11339,N_11180,N_11102);
or U11340 (N_11340,N_11110,N_11163);
nor U11341 (N_11341,N_11012,N_11079);
nor U11342 (N_11342,N_11177,N_11031);
and U11343 (N_11343,N_11068,N_11169);
or U11344 (N_11344,N_11075,N_11163);
nor U11345 (N_11345,N_11101,N_11015);
nor U11346 (N_11346,N_11187,N_11018);
xnor U11347 (N_11347,N_11170,N_11104);
xor U11348 (N_11348,N_11196,N_11063);
or U11349 (N_11349,N_11073,N_11012);
xor U11350 (N_11350,N_11093,N_11009);
nor U11351 (N_11351,N_11061,N_11041);
nor U11352 (N_11352,N_11088,N_11152);
or U11353 (N_11353,N_11040,N_11145);
xor U11354 (N_11354,N_11130,N_11010);
nand U11355 (N_11355,N_11186,N_11122);
nand U11356 (N_11356,N_11185,N_11058);
xnor U11357 (N_11357,N_11140,N_11155);
nand U11358 (N_11358,N_11112,N_11195);
or U11359 (N_11359,N_11189,N_11032);
and U11360 (N_11360,N_11195,N_11165);
nand U11361 (N_11361,N_11178,N_11084);
nand U11362 (N_11362,N_11011,N_11091);
and U11363 (N_11363,N_11115,N_11136);
xnor U11364 (N_11364,N_11065,N_11186);
xor U11365 (N_11365,N_11103,N_11076);
xnor U11366 (N_11366,N_11045,N_11082);
xnor U11367 (N_11367,N_11092,N_11061);
xnor U11368 (N_11368,N_11156,N_11054);
or U11369 (N_11369,N_11045,N_11105);
nand U11370 (N_11370,N_11117,N_11068);
and U11371 (N_11371,N_11084,N_11046);
and U11372 (N_11372,N_11091,N_11125);
or U11373 (N_11373,N_11157,N_11170);
or U11374 (N_11374,N_11158,N_11008);
xnor U11375 (N_11375,N_11176,N_11191);
and U11376 (N_11376,N_11064,N_11184);
nor U11377 (N_11377,N_11035,N_11118);
and U11378 (N_11378,N_11015,N_11122);
or U11379 (N_11379,N_11010,N_11140);
or U11380 (N_11380,N_11063,N_11014);
nor U11381 (N_11381,N_11101,N_11166);
or U11382 (N_11382,N_11059,N_11062);
nand U11383 (N_11383,N_11020,N_11037);
and U11384 (N_11384,N_11118,N_11170);
nand U11385 (N_11385,N_11173,N_11127);
or U11386 (N_11386,N_11051,N_11123);
xor U11387 (N_11387,N_11079,N_11033);
nand U11388 (N_11388,N_11121,N_11181);
xor U11389 (N_11389,N_11166,N_11020);
nand U11390 (N_11390,N_11011,N_11112);
and U11391 (N_11391,N_11146,N_11018);
xor U11392 (N_11392,N_11091,N_11015);
nor U11393 (N_11393,N_11125,N_11094);
or U11394 (N_11394,N_11023,N_11155);
xnor U11395 (N_11395,N_11188,N_11072);
nand U11396 (N_11396,N_11104,N_11036);
nor U11397 (N_11397,N_11064,N_11167);
and U11398 (N_11398,N_11091,N_11030);
xor U11399 (N_11399,N_11128,N_11016);
and U11400 (N_11400,N_11273,N_11281);
or U11401 (N_11401,N_11307,N_11371);
and U11402 (N_11402,N_11296,N_11324);
nor U11403 (N_11403,N_11318,N_11383);
xor U11404 (N_11404,N_11344,N_11381);
nand U11405 (N_11405,N_11304,N_11360);
nor U11406 (N_11406,N_11239,N_11361);
nor U11407 (N_11407,N_11250,N_11300);
and U11408 (N_11408,N_11372,N_11235);
xnor U11409 (N_11409,N_11395,N_11275);
or U11410 (N_11410,N_11214,N_11282);
nor U11411 (N_11411,N_11325,N_11340);
or U11412 (N_11412,N_11306,N_11370);
or U11413 (N_11413,N_11295,N_11261);
nand U11414 (N_11414,N_11397,N_11299);
and U11415 (N_11415,N_11277,N_11346);
nor U11416 (N_11416,N_11331,N_11270);
and U11417 (N_11417,N_11268,N_11216);
and U11418 (N_11418,N_11218,N_11319);
xnor U11419 (N_11419,N_11394,N_11366);
or U11420 (N_11420,N_11212,N_11352);
or U11421 (N_11421,N_11380,N_11351);
and U11422 (N_11422,N_11386,N_11206);
or U11423 (N_11423,N_11271,N_11338);
xor U11424 (N_11424,N_11312,N_11356);
and U11425 (N_11425,N_11263,N_11251);
or U11426 (N_11426,N_11339,N_11285);
or U11427 (N_11427,N_11327,N_11228);
and U11428 (N_11428,N_11389,N_11208);
or U11429 (N_11429,N_11237,N_11376);
xnor U11430 (N_11430,N_11258,N_11230);
or U11431 (N_11431,N_11238,N_11269);
nand U11432 (N_11432,N_11278,N_11320);
nor U11433 (N_11433,N_11355,N_11232);
and U11434 (N_11434,N_11233,N_11336);
nor U11435 (N_11435,N_11375,N_11350);
or U11436 (N_11436,N_11315,N_11220);
xor U11437 (N_11437,N_11219,N_11321);
nand U11438 (N_11438,N_11367,N_11288);
and U11439 (N_11439,N_11293,N_11294);
or U11440 (N_11440,N_11290,N_11333);
nand U11441 (N_11441,N_11378,N_11347);
or U11442 (N_11442,N_11283,N_11213);
and U11443 (N_11443,N_11255,N_11203);
xor U11444 (N_11444,N_11259,N_11326);
or U11445 (N_11445,N_11354,N_11246);
or U11446 (N_11446,N_11279,N_11374);
nor U11447 (N_11447,N_11314,N_11210);
or U11448 (N_11448,N_11265,N_11217);
and U11449 (N_11449,N_11398,N_11317);
or U11450 (N_11450,N_11349,N_11335);
xor U11451 (N_11451,N_11254,N_11382);
nor U11452 (N_11452,N_11393,N_11241);
xnor U11453 (N_11453,N_11345,N_11364);
nor U11454 (N_11454,N_11363,N_11262);
nand U11455 (N_11455,N_11234,N_11209);
xor U11456 (N_11456,N_11253,N_11342);
nand U11457 (N_11457,N_11266,N_11298);
nor U11458 (N_11458,N_11256,N_11245);
nor U11459 (N_11459,N_11303,N_11353);
or U11460 (N_11460,N_11276,N_11286);
or U11461 (N_11461,N_11343,N_11201);
or U11462 (N_11462,N_11316,N_11249);
nand U11463 (N_11463,N_11247,N_11248);
or U11464 (N_11464,N_11231,N_11387);
xor U11465 (N_11465,N_11292,N_11243);
nor U11466 (N_11466,N_11240,N_11384);
and U11467 (N_11467,N_11310,N_11396);
nor U11468 (N_11468,N_11392,N_11297);
nor U11469 (N_11469,N_11244,N_11272);
xnor U11470 (N_11470,N_11313,N_11267);
and U11471 (N_11471,N_11221,N_11202);
nor U11472 (N_11472,N_11229,N_11260);
nor U11473 (N_11473,N_11385,N_11274);
and U11474 (N_11474,N_11204,N_11226);
and U11475 (N_11475,N_11284,N_11330);
nor U11476 (N_11476,N_11391,N_11358);
and U11477 (N_11477,N_11379,N_11301);
or U11478 (N_11478,N_11287,N_11236);
xnor U11479 (N_11479,N_11215,N_11264);
xor U11480 (N_11480,N_11329,N_11311);
or U11481 (N_11481,N_11305,N_11308);
nand U11482 (N_11482,N_11390,N_11224);
nand U11483 (N_11483,N_11337,N_11377);
nand U11484 (N_11484,N_11280,N_11323);
and U11485 (N_11485,N_11205,N_11362);
xor U11486 (N_11486,N_11348,N_11365);
and U11487 (N_11487,N_11200,N_11399);
or U11488 (N_11488,N_11341,N_11211);
xor U11489 (N_11489,N_11242,N_11289);
nand U11490 (N_11490,N_11291,N_11332);
or U11491 (N_11491,N_11359,N_11223);
xor U11492 (N_11492,N_11388,N_11369);
xor U11493 (N_11493,N_11322,N_11222);
xor U11494 (N_11494,N_11257,N_11373);
nand U11495 (N_11495,N_11309,N_11334);
or U11496 (N_11496,N_11207,N_11252);
and U11497 (N_11497,N_11227,N_11357);
xor U11498 (N_11498,N_11225,N_11368);
xnor U11499 (N_11499,N_11302,N_11328);
nor U11500 (N_11500,N_11249,N_11340);
xor U11501 (N_11501,N_11327,N_11287);
or U11502 (N_11502,N_11264,N_11334);
nand U11503 (N_11503,N_11308,N_11298);
nor U11504 (N_11504,N_11253,N_11336);
xor U11505 (N_11505,N_11310,N_11305);
nor U11506 (N_11506,N_11379,N_11370);
or U11507 (N_11507,N_11318,N_11235);
nor U11508 (N_11508,N_11201,N_11360);
xnor U11509 (N_11509,N_11296,N_11242);
nand U11510 (N_11510,N_11311,N_11246);
nand U11511 (N_11511,N_11363,N_11240);
nor U11512 (N_11512,N_11374,N_11300);
and U11513 (N_11513,N_11259,N_11269);
nand U11514 (N_11514,N_11382,N_11243);
or U11515 (N_11515,N_11248,N_11343);
or U11516 (N_11516,N_11214,N_11344);
or U11517 (N_11517,N_11380,N_11224);
nand U11518 (N_11518,N_11368,N_11241);
or U11519 (N_11519,N_11252,N_11399);
or U11520 (N_11520,N_11219,N_11218);
xnor U11521 (N_11521,N_11349,N_11324);
xor U11522 (N_11522,N_11310,N_11211);
nand U11523 (N_11523,N_11236,N_11372);
and U11524 (N_11524,N_11369,N_11234);
nor U11525 (N_11525,N_11339,N_11316);
and U11526 (N_11526,N_11351,N_11236);
or U11527 (N_11527,N_11362,N_11239);
xnor U11528 (N_11528,N_11386,N_11239);
nor U11529 (N_11529,N_11363,N_11324);
nor U11530 (N_11530,N_11352,N_11293);
nand U11531 (N_11531,N_11297,N_11364);
nand U11532 (N_11532,N_11231,N_11319);
nand U11533 (N_11533,N_11379,N_11239);
nor U11534 (N_11534,N_11233,N_11304);
and U11535 (N_11535,N_11325,N_11377);
xor U11536 (N_11536,N_11277,N_11254);
or U11537 (N_11537,N_11365,N_11223);
nand U11538 (N_11538,N_11204,N_11253);
and U11539 (N_11539,N_11272,N_11254);
nand U11540 (N_11540,N_11364,N_11225);
and U11541 (N_11541,N_11248,N_11203);
xnor U11542 (N_11542,N_11368,N_11342);
or U11543 (N_11543,N_11215,N_11363);
and U11544 (N_11544,N_11360,N_11349);
or U11545 (N_11545,N_11262,N_11274);
nor U11546 (N_11546,N_11239,N_11228);
nor U11547 (N_11547,N_11271,N_11215);
nor U11548 (N_11548,N_11368,N_11239);
xnor U11549 (N_11549,N_11363,N_11294);
or U11550 (N_11550,N_11344,N_11231);
or U11551 (N_11551,N_11220,N_11249);
nand U11552 (N_11552,N_11344,N_11308);
nand U11553 (N_11553,N_11349,N_11333);
or U11554 (N_11554,N_11389,N_11317);
and U11555 (N_11555,N_11360,N_11328);
and U11556 (N_11556,N_11346,N_11236);
and U11557 (N_11557,N_11273,N_11254);
nand U11558 (N_11558,N_11211,N_11201);
xor U11559 (N_11559,N_11260,N_11227);
xor U11560 (N_11560,N_11226,N_11398);
or U11561 (N_11561,N_11317,N_11335);
and U11562 (N_11562,N_11312,N_11255);
nand U11563 (N_11563,N_11320,N_11287);
or U11564 (N_11564,N_11261,N_11364);
nor U11565 (N_11565,N_11236,N_11349);
nand U11566 (N_11566,N_11215,N_11337);
or U11567 (N_11567,N_11285,N_11220);
or U11568 (N_11568,N_11215,N_11388);
nand U11569 (N_11569,N_11258,N_11231);
or U11570 (N_11570,N_11393,N_11212);
and U11571 (N_11571,N_11226,N_11307);
nand U11572 (N_11572,N_11249,N_11234);
and U11573 (N_11573,N_11357,N_11281);
or U11574 (N_11574,N_11344,N_11293);
nor U11575 (N_11575,N_11365,N_11278);
nor U11576 (N_11576,N_11372,N_11399);
nor U11577 (N_11577,N_11224,N_11266);
nor U11578 (N_11578,N_11268,N_11326);
nand U11579 (N_11579,N_11366,N_11208);
or U11580 (N_11580,N_11258,N_11302);
nand U11581 (N_11581,N_11332,N_11296);
and U11582 (N_11582,N_11239,N_11277);
nor U11583 (N_11583,N_11260,N_11206);
xnor U11584 (N_11584,N_11217,N_11367);
and U11585 (N_11585,N_11394,N_11343);
xnor U11586 (N_11586,N_11362,N_11204);
nor U11587 (N_11587,N_11259,N_11201);
nand U11588 (N_11588,N_11255,N_11384);
nor U11589 (N_11589,N_11386,N_11302);
nand U11590 (N_11590,N_11290,N_11365);
nor U11591 (N_11591,N_11247,N_11398);
nor U11592 (N_11592,N_11205,N_11309);
nand U11593 (N_11593,N_11246,N_11368);
xor U11594 (N_11594,N_11222,N_11203);
and U11595 (N_11595,N_11219,N_11331);
xnor U11596 (N_11596,N_11370,N_11285);
xor U11597 (N_11597,N_11254,N_11263);
and U11598 (N_11598,N_11268,N_11286);
nor U11599 (N_11599,N_11264,N_11306);
or U11600 (N_11600,N_11550,N_11529);
xnor U11601 (N_11601,N_11538,N_11598);
xnor U11602 (N_11602,N_11522,N_11430);
xnor U11603 (N_11603,N_11542,N_11473);
and U11604 (N_11604,N_11541,N_11585);
nor U11605 (N_11605,N_11444,N_11419);
xnor U11606 (N_11606,N_11545,N_11517);
xor U11607 (N_11607,N_11401,N_11425);
and U11608 (N_11608,N_11488,N_11532);
nand U11609 (N_11609,N_11597,N_11526);
and U11610 (N_11610,N_11505,N_11451);
and U11611 (N_11611,N_11596,N_11470);
and U11612 (N_11612,N_11589,N_11495);
nand U11613 (N_11613,N_11429,N_11551);
nand U11614 (N_11614,N_11439,N_11588);
nand U11615 (N_11615,N_11516,N_11530);
nor U11616 (N_11616,N_11410,N_11485);
and U11617 (N_11617,N_11533,N_11564);
and U11618 (N_11618,N_11497,N_11464);
nand U11619 (N_11619,N_11524,N_11463);
and U11620 (N_11620,N_11574,N_11513);
and U11621 (N_11621,N_11456,N_11504);
xnor U11622 (N_11622,N_11440,N_11527);
nor U11623 (N_11623,N_11549,N_11432);
xor U11624 (N_11624,N_11474,N_11537);
or U11625 (N_11625,N_11431,N_11577);
nand U11626 (N_11626,N_11466,N_11400);
or U11627 (N_11627,N_11565,N_11515);
and U11628 (N_11628,N_11482,N_11540);
xnor U11629 (N_11629,N_11594,N_11519);
xor U11630 (N_11630,N_11479,N_11567);
nand U11631 (N_11631,N_11460,N_11490);
nor U11632 (N_11632,N_11592,N_11560);
and U11633 (N_11633,N_11536,N_11579);
or U11634 (N_11634,N_11489,N_11581);
or U11635 (N_11635,N_11418,N_11499);
nand U11636 (N_11636,N_11465,N_11544);
nand U11637 (N_11637,N_11476,N_11468);
nor U11638 (N_11638,N_11571,N_11539);
or U11639 (N_11639,N_11423,N_11576);
and U11640 (N_11640,N_11434,N_11555);
and U11641 (N_11641,N_11484,N_11518);
and U11642 (N_11642,N_11500,N_11573);
or U11643 (N_11643,N_11587,N_11453);
and U11644 (N_11644,N_11559,N_11591);
and U11645 (N_11645,N_11520,N_11417);
or U11646 (N_11646,N_11409,N_11510);
nor U11647 (N_11647,N_11575,N_11424);
xor U11648 (N_11648,N_11547,N_11411);
xor U11649 (N_11649,N_11442,N_11584);
xnor U11650 (N_11650,N_11512,N_11452);
and U11651 (N_11651,N_11438,N_11523);
nand U11652 (N_11652,N_11507,N_11494);
nand U11653 (N_11653,N_11435,N_11552);
nor U11654 (N_11654,N_11449,N_11459);
nor U11655 (N_11655,N_11590,N_11531);
xnor U11656 (N_11656,N_11480,N_11428);
nor U11657 (N_11657,N_11582,N_11487);
xor U11658 (N_11658,N_11471,N_11416);
nand U11659 (N_11659,N_11501,N_11553);
nand U11660 (N_11660,N_11441,N_11483);
xor U11661 (N_11661,N_11569,N_11508);
or U11662 (N_11662,N_11427,N_11593);
xnor U11663 (N_11663,N_11445,N_11437);
nand U11664 (N_11664,N_11448,N_11525);
xnor U11665 (N_11665,N_11422,N_11511);
nand U11666 (N_11666,N_11405,N_11583);
xnor U11667 (N_11667,N_11469,N_11412);
nand U11668 (N_11668,N_11570,N_11514);
or U11669 (N_11669,N_11415,N_11458);
or U11670 (N_11670,N_11481,N_11454);
or U11671 (N_11671,N_11478,N_11420);
and U11672 (N_11672,N_11436,N_11580);
nor U11673 (N_11673,N_11599,N_11509);
and U11674 (N_11674,N_11462,N_11486);
or U11675 (N_11675,N_11556,N_11461);
nand U11676 (N_11676,N_11595,N_11457);
or U11677 (N_11677,N_11414,N_11433);
and U11678 (N_11678,N_11491,N_11402);
nor U11679 (N_11679,N_11421,N_11408);
or U11680 (N_11680,N_11563,N_11443);
and U11681 (N_11681,N_11546,N_11455);
nor U11682 (N_11682,N_11450,N_11406);
and U11683 (N_11683,N_11426,N_11534);
or U11684 (N_11684,N_11543,N_11561);
or U11685 (N_11685,N_11535,N_11578);
nand U11686 (N_11686,N_11528,N_11493);
nor U11687 (N_11687,N_11562,N_11566);
and U11688 (N_11688,N_11572,N_11404);
nand U11689 (N_11689,N_11496,N_11413);
xnor U11690 (N_11690,N_11502,N_11467);
nand U11691 (N_11691,N_11554,N_11506);
xnor U11692 (N_11692,N_11477,N_11447);
nand U11693 (N_11693,N_11503,N_11568);
and U11694 (N_11694,N_11407,N_11446);
and U11695 (N_11695,N_11475,N_11558);
nor U11696 (N_11696,N_11472,N_11586);
nor U11697 (N_11697,N_11498,N_11557);
and U11698 (N_11698,N_11492,N_11521);
nand U11699 (N_11699,N_11548,N_11403);
nand U11700 (N_11700,N_11598,N_11579);
nand U11701 (N_11701,N_11486,N_11593);
xor U11702 (N_11702,N_11575,N_11580);
or U11703 (N_11703,N_11478,N_11411);
or U11704 (N_11704,N_11560,N_11446);
or U11705 (N_11705,N_11503,N_11484);
nand U11706 (N_11706,N_11559,N_11545);
nand U11707 (N_11707,N_11480,N_11445);
nand U11708 (N_11708,N_11404,N_11411);
and U11709 (N_11709,N_11595,N_11463);
nor U11710 (N_11710,N_11434,N_11499);
or U11711 (N_11711,N_11477,N_11571);
and U11712 (N_11712,N_11427,N_11472);
or U11713 (N_11713,N_11465,N_11586);
or U11714 (N_11714,N_11497,N_11544);
or U11715 (N_11715,N_11432,N_11402);
xnor U11716 (N_11716,N_11529,N_11598);
xor U11717 (N_11717,N_11483,N_11583);
nand U11718 (N_11718,N_11598,N_11499);
xnor U11719 (N_11719,N_11400,N_11582);
and U11720 (N_11720,N_11482,N_11433);
and U11721 (N_11721,N_11511,N_11587);
nand U11722 (N_11722,N_11539,N_11457);
or U11723 (N_11723,N_11580,N_11432);
nor U11724 (N_11724,N_11548,N_11444);
nand U11725 (N_11725,N_11597,N_11416);
nand U11726 (N_11726,N_11410,N_11522);
or U11727 (N_11727,N_11421,N_11560);
and U11728 (N_11728,N_11591,N_11529);
or U11729 (N_11729,N_11438,N_11428);
nor U11730 (N_11730,N_11432,N_11527);
and U11731 (N_11731,N_11516,N_11579);
or U11732 (N_11732,N_11441,N_11571);
nand U11733 (N_11733,N_11410,N_11470);
and U11734 (N_11734,N_11411,N_11586);
and U11735 (N_11735,N_11550,N_11501);
nand U11736 (N_11736,N_11548,N_11472);
and U11737 (N_11737,N_11460,N_11469);
and U11738 (N_11738,N_11489,N_11427);
xor U11739 (N_11739,N_11470,N_11477);
or U11740 (N_11740,N_11409,N_11414);
xnor U11741 (N_11741,N_11526,N_11517);
and U11742 (N_11742,N_11550,N_11413);
nand U11743 (N_11743,N_11569,N_11401);
xor U11744 (N_11744,N_11515,N_11541);
and U11745 (N_11745,N_11494,N_11584);
nor U11746 (N_11746,N_11581,N_11496);
or U11747 (N_11747,N_11503,N_11562);
xor U11748 (N_11748,N_11488,N_11510);
or U11749 (N_11749,N_11457,N_11551);
nand U11750 (N_11750,N_11505,N_11532);
xnor U11751 (N_11751,N_11546,N_11483);
nand U11752 (N_11752,N_11401,N_11465);
nor U11753 (N_11753,N_11547,N_11552);
nand U11754 (N_11754,N_11484,N_11487);
and U11755 (N_11755,N_11529,N_11506);
nand U11756 (N_11756,N_11576,N_11479);
or U11757 (N_11757,N_11467,N_11464);
nor U11758 (N_11758,N_11538,N_11570);
nand U11759 (N_11759,N_11529,N_11492);
or U11760 (N_11760,N_11593,N_11491);
nand U11761 (N_11761,N_11443,N_11571);
nand U11762 (N_11762,N_11562,N_11556);
nand U11763 (N_11763,N_11501,N_11522);
nor U11764 (N_11764,N_11453,N_11416);
xor U11765 (N_11765,N_11503,N_11402);
xnor U11766 (N_11766,N_11579,N_11566);
nand U11767 (N_11767,N_11501,N_11470);
and U11768 (N_11768,N_11552,N_11561);
nor U11769 (N_11769,N_11577,N_11422);
nand U11770 (N_11770,N_11585,N_11415);
nand U11771 (N_11771,N_11560,N_11451);
and U11772 (N_11772,N_11546,N_11573);
nand U11773 (N_11773,N_11439,N_11403);
nor U11774 (N_11774,N_11507,N_11500);
xnor U11775 (N_11775,N_11565,N_11418);
or U11776 (N_11776,N_11436,N_11561);
or U11777 (N_11777,N_11502,N_11535);
and U11778 (N_11778,N_11503,N_11468);
or U11779 (N_11779,N_11501,N_11554);
or U11780 (N_11780,N_11554,N_11482);
nand U11781 (N_11781,N_11415,N_11420);
nand U11782 (N_11782,N_11470,N_11534);
and U11783 (N_11783,N_11562,N_11404);
xor U11784 (N_11784,N_11576,N_11447);
or U11785 (N_11785,N_11468,N_11422);
and U11786 (N_11786,N_11460,N_11474);
xnor U11787 (N_11787,N_11547,N_11579);
nand U11788 (N_11788,N_11543,N_11491);
nand U11789 (N_11789,N_11505,N_11581);
xnor U11790 (N_11790,N_11475,N_11416);
and U11791 (N_11791,N_11484,N_11430);
and U11792 (N_11792,N_11574,N_11442);
and U11793 (N_11793,N_11429,N_11435);
nor U11794 (N_11794,N_11454,N_11491);
nand U11795 (N_11795,N_11512,N_11460);
nor U11796 (N_11796,N_11412,N_11571);
and U11797 (N_11797,N_11459,N_11479);
nor U11798 (N_11798,N_11547,N_11436);
xnor U11799 (N_11799,N_11425,N_11459);
xnor U11800 (N_11800,N_11628,N_11738);
nor U11801 (N_11801,N_11656,N_11630);
nand U11802 (N_11802,N_11649,N_11781);
or U11803 (N_11803,N_11728,N_11724);
nand U11804 (N_11804,N_11777,N_11689);
nand U11805 (N_11805,N_11690,N_11679);
nand U11806 (N_11806,N_11662,N_11796);
or U11807 (N_11807,N_11652,N_11703);
nor U11808 (N_11808,N_11665,N_11647);
or U11809 (N_11809,N_11697,N_11623);
and U11810 (N_11810,N_11775,N_11766);
nor U11811 (N_11811,N_11734,N_11650);
xnor U11812 (N_11812,N_11735,N_11745);
nand U11813 (N_11813,N_11671,N_11711);
nand U11814 (N_11814,N_11789,N_11718);
xnor U11815 (N_11815,N_11691,N_11622);
nand U11816 (N_11816,N_11799,N_11765);
and U11817 (N_11817,N_11706,N_11715);
or U11818 (N_11818,N_11739,N_11700);
and U11819 (N_11819,N_11615,N_11772);
nor U11820 (N_11820,N_11756,N_11627);
nand U11821 (N_11821,N_11654,N_11644);
nor U11822 (N_11822,N_11680,N_11741);
and U11823 (N_11823,N_11790,N_11674);
xor U11824 (N_11824,N_11714,N_11784);
or U11825 (N_11825,N_11685,N_11768);
nor U11826 (N_11826,N_11707,N_11661);
xor U11827 (N_11827,N_11698,N_11636);
xor U11828 (N_11828,N_11776,N_11732);
nor U11829 (N_11829,N_11709,N_11641);
nand U11830 (N_11830,N_11786,N_11648);
and U11831 (N_11831,N_11607,N_11693);
nor U11832 (N_11832,N_11792,N_11663);
nand U11833 (N_11833,N_11687,N_11755);
or U11834 (N_11834,N_11631,N_11740);
xor U11835 (N_11835,N_11730,N_11651);
and U11836 (N_11836,N_11609,N_11645);
or U11837 (N_11837,N_11702,N_11721);
or U11838 (N_11838,N_11795,N_11722);
nand U11839 (N_11839,N_11770,N_11646);
nand U11840 (N_11840,N_11759,N_11643);
xnor U11841 (N_11841,N_11794,N_11601);
nand U11842 (N_11842,N_11664,N_11639);
nand U11843 (N_11843,N_11783,N_11633);
nor U11844 (N_11844,N_11752,N_11604);
and U11845 (N_11845,N_11637,N_11798);
nor U11846 (N_11846,N_11769,N_11780);
nor U11847 (N_11847,N_11611,N_11600);
nand U11848 (N_11848,N_11712,N_11653);
nand U11849 (N_11849,N_11655,N_11625);
nand U11850 (N_11850,N_11729,N_11632);
xnor U11851 (N_11851,N_11678,N_11761);
nor U11852 (N_11852,N_11793,N_11713);
xor U11853 (N_11853,N_11725,N_11668);
xnor U11854 (N_11854,N_11701,N_11767);
or U11855 (N_11855,N_11719,N_11788);
nor U11856 (N_11856,N_11708,N_11749);
and U11857 (N_11857,N_11757,N_11660);
and U11858 (N_11858,N_11629,N_11603);
and U11859 (N_11859,N_11602,N_11751);
or U11860 (N_11860,N_11797,N_11620);
and U11861 (N_11861,N_11605,N_11758);
or U11862 (N_11862,N_11624,N_11753);
nand U11863 (N_11863,N_11720,N_11778);
or U11864 (N_11864,N_11677,N_11747);
xnor U11865 (N_11865,N_11705,N_11688);
and U11866 (N_11866,N_11617,N_11676);
xor U11867 (N_11867,N_11785,N_11670);
xnor U11868 (N_11868,N_11726,N_11658);
and U11869 (N_11869,N_11657,N_11616);
nor U11870 (N_11870,N_11686,N_11672);
and U11871 (N_11871,N_11774,N_11748);
nor U11872 (N_11872,N_11710,N_11659);
and U11873 (N_11873,N_11779,N_11736);
nand U11874 (N_11874,N_11760,N_11764);
nand U11875 (N_11875,N_11744,N_11762);
and U11876 (N_11876,N_11723,N_11699);
xnor U11877 (N_11877,N_11737,N_11684);
nand U11878 (N_11878,N_11666,N_11704);
nor U11879 (N_11879,N_11773,N_11621);
and U11880 (N_11880,N_11743,N_11669);
or U11881 (N_11881,N_11608,N_11675);
nand U11882 (N_11882,N_11750,N_11613);
nor U11883 (N_11883,N_11754,N_11618);
and U11884 (N_11884,N_11695,N_11727);
nand U11885 (N_11885,N_11746,N_11642);
xor U11886 (N_11886,N_11731,N_11638);
and U11887 (N_11887,N_11667,N_11640);
or U11888 (N_11888,N_11763,N_11610);
and U11889 (N_11889,N_11782,N_11635);
nor U11890 (N_11890,N_11626,N_11681);
or U11891 (N_11891,N_11614,N_11673);
and U11892 (N_11892,N_11742,N_11696);
and U11893 (N_11893,N_11717,N_11733);
nand U11894 (N_11894,N_11682,N_11771);
or U11895 (N_11895,N_11612,N_11692);
nand U11896 (N_11896,N_11791,N_11683);
nor U11897 (N_11897,N_11716,N_11619);
nor U11898 (N_11898,N_11787,N_11694);
nor U11899 (N_11899,N_11634,N_11606);
or U11900 (N_11900,N_11647,N_11747);
xor U11901 (N_11901,N_11716,N_11767);
nand U11902 (N_11902,N_11621,N_11639);
or U11903 (N_11903,N_11689,N_11660);
or U11904 (N_11904,N_11715,N_11739);
xnor U11905 (N_11905,N_11696,N_11744);
xnor U11906 (N_11906,N_11794,N_11793);
or U11907 (N_11907,N_11776,N_11708);
nor U11908 (N_11908,N_11768,N_11793);
and U11909 (N_11909,N_11707,N_11772);
and U11910 (N_11910,N_11604,N_11749);
and U11911 (N_11911,N_11691,N_11696);
nand U11912 (N_11912,N_11603,N_11661);
nand U11913 (N_11913,N_11721,N_11688);
nand U11914 (N_11914,N_11636,N_11612);
and U11915 (N_11915,N_11771,N_11784);
xor U11916 (N_11916,N_11715,N_11609);
and U11917 (N_11917,N_11768,N_11672);
xor U11918 (N_11918,N_11773,N_11767);
and U11919 (N_11919,N_11677,N_11716);
and U11920 (N_11920,N_11638,N_11673);
and U11921 (N_11921,N_11661,N_11692);
nand U11922 (N_11922,N_11694,N_11617);
nand U11923 (N_11923,N_11645,N_11734);
or U11924 (N_11924,N_11606,N_11761);
xnor U11925 (N_11925,N_11670,N_11677);
nand U11926 (N_11926,N_11703,N_11684);
and U11927 (N_11927,N_11736,N_11788);
or U11928 (N_11928,N_11776,N_11661);
xor U11929 (N_11929,N_11688,N_11712);
nor U11930 (N_11930,N_11716,N_11785);
or U11931 (N_11931,N_11742,N_11656);
or U11932 (N_11932,N_11762,N_11699);
xnor U11933 (N_11933,N_11703,N_11620);
nand U11934 (N_11934,N_11709,N_11788);
and U11935 (N_11935,N_11756,N_11691);
xnor U11936 (N_11936,N_11753,N_11745);
and U11937 (N_11937,N_11788,N_11742);
or U11938 (N_11938,N_11765,N_11719);
nor U11939 (N_11939,N_11684,N_11655);
and U11940 (N_11940,N_11723,N_11652);
nor U11941 (N_11941,N_11679,N_11789);
xnor U11942 (N_11942,N_11782,N_11601);
nor U11943 (N_11943,N_11695,N_11736);
xor U11944 (N_11944,N_11644,N_11759);
or U11945 (N_11945,N_11647,N_11689);
nand U11946 (N_11946,N_11656,N_11644);
nor U11947 (N_11947,N_11773,N_11783);
xnor U11948 (N_11948,N_11711,N_11767);
and U11949 (N_11949,N_11620,N_11659);
nand U11950 (N_11950,N_11617,N_11625);
nand U11951 (N_11951,N_11744,N_11659);
nor U11952 (N_11952,N_11691,N_11752);
nor U11953 (N_11953,N_11605,N_11699);
nand U11954 (N_11954,N_11778,N_11775);
or U11955 (N_11955,N_11741,N_11654);
nand U11956 (N_11956,N_11752,N_11746);
xnor U11957 (N_11957,N_11770,N_11608);
xnor U11958 (N_11958,N_11717,N_11725);
nor U11959 (N_11959,N_11782,N_11600);
xor U11960 (N_11960,N_11715,N_11724);
xor U11961 (N_11961,N_11785,N_11795);
xnor U11962 (N_11962,N_11609,N_11746);
or U11963 (N_11963,N_11688,N_11738);
nand U11964 (N_11964,N_11720,N_11603);
or U11965 (N_11965,N_11721,N_11686);
or U11966 (N_11966,N_11734,N_11765);
nor U11967 (N_11967,N_11768,N_11606);
nand U11968 (N_11968,N_11685,N_11673);
or U11969 (N_11969,N_11745,N_11787);
nor U11970 (N_11970,N_11752,N_11780);
nor U11971 (N_11971,N_11600,N_11765);
nand U11972 (N_11972,N_11785,N_11701);
xor U11973 (N_11973,N_11708,N_11735);
xor U11974 (N_11974,N_11740,N_11798);
nor U11975 (N_11975,N_11733,N_11625);
nor U11976 (N_11976,N_11611,N_11692);
xor U11977 (N_11977,N_11743,N_11733);
and U11978 (N_11978,N_11741,N_11759);
nand U11979 (N_11979,N_11622,N_11774);
xor U11980 (N_11980,N_11696,N_11705);
or U11981 (N_11981,N_11798,N_11705);
and U11982 (N_11982,N_11706,N_11625);
xor U11983 (N_11983,N_11782,N_11665);
nor U11984 (N_11984,N_11654,N_11680);
nand U11985 (N_11985,N_11786,N_11626);
nand U11986 (N_11986,N_11709,N_11765);
nor U11987 (N_11987,N_11790,N_11614);
nand U11988 (N_11988,N_11770,N_11794);
xor U11989 (N_11989,N_11767,N_11655);
or U11990 (N_11990,N_11692,N_11788);
and U11991 (N_11991,N_11697,N_11610);
nor U11992 (N_11992,N_11703,N_11649);
and U11993 (N_11993,N_11685,N_11666);
and U11994 (N_11994,N_11643,N_11629);
and U11995 (N_11995,N_11689,N_11616);
and U11996 (N_11996,N_11714,N_11708);
nor U11997 (N_11997,N_11609,N_11632);
nor U11998 (N_11998,N_11641,N_11648);
nor U11999 (N_11999,N_11701,N_11739);
and U12000 (N_12000,N_11958,N_11904);
xnor U12001 (N_12001,N_11963,N_11872);
xnor U12002 (N_12002,N_11964,N_11892);
and U12003 (N_12003,N_11837,N_11985);
nor U12004 (N_12004,N_11979,N_11959);
nor U12005 (N_12005,N_11899,N_11801);
or U12006 (N_12006,N_11867,N_11877);
or U12007 (N_12007,N_11853,N_11978);
xor U12008 (N_12008,N_11950,N_11934);
nand U12009 (N_12009,N_11905,N_11921);
or U12010 (N_12010,N_11819,N_11893);
xnor U12011 (N_12011,N_11957,N_11891);
nand U12012 (N_12012,N_11831,N_11902);
xor U12013 (N_12013,N_11937,N_11940);
and U12014 (N_12014,N_11879,N_11823);
nor U12015 (N_12015,N_11929,N_11960);
xnor U12016 (N_12016,N_11806,N_11884);
and U12017 (N_12017,N_11843,N_11896);
or U12018 (N_12018,N_11862,N_11961);
or U12019 (N_12019,N_11920,N_11817);
nand U12020 (N_12020,N_11822,N_11995);
or U12021 (N_12021,N_11821,N_11873);
or U12022 (N_12022,N_11974,N_11878);
or U12023 (N_12023,N_11887,N_11973);
nand U12024 (N_12024,N_11888,N_11859);
or U12025 (N_12025,N_11871,N_11881);
nand U12026 (N_12026,N_11952,N_11983);
xor U12027 (N_12027,N_11971,N_11953);
or U12028 (N_12028,N_11918,N_11816);
and U12029 (N_12029,N_11970,N_11815);
xor U12030 (N_12030,N_11908,N_11809);
xor U12031 (N_12031,N_11839,N_11863);
or U12032 (N_12032,N_11860,N_11939);
and U12033 (N_12033,N_11840,N_11868);
nand U12034 (N_12034,N_11900,N_11930);
and U12035 (N_12035,N_11852,N_11814);
nand U12036 (N_12036,N_11906,N_11987);
or U12037 (N_12037,N_11890,N_11850);
and U12038 (N_12038,N_11870,N_11812);
or U12039 (N_12039,N_11803,N_11975);
nor U12040 (N_12040,N_11966,N_11886);
xor U12041 (N_12041,N_11914,N_11829);
and U12042 (N_12042,N_11866,N_11986);
nand U12043 (N_12043,N_11810,N_11869);
nor U12044 (N_12044,N_11947,N_11933);
nor U12045 (N_12045,N_11999,N_11827);
and U12046 (N_12046,N_11844,N_11845);
xor U12047 (N_12047,N_11944,N_11976);
nand U12048 (N_12048,N_11898,N_11993);
nand U12049 (N_12049,N_11931,N_11805);
or U12050 (N_12050,N_11855,N_11991);
nand U12051 (N_12051,N_11980,N_11928);
or U12052 (N_12052,N_11962,N_11897);
nor U12053 (N_12053,N_11820,N_11932);
nand U12054 (N_12054,N_11936,N_11923);
nor U12055 (N_12055,N_11834,N_11955);
or U12056 (N_12056,N_11903,N_11941);
xor U12057 (N_12057,N_11846,N_11917);
nand U12058 (N_12058,N_11996,N_11984);
xor U12059 (N_12059,N_11838,N_11948);
nor U12060 (N_12060,N_11800,N_11938);
nor U12061 (N_12061,N_11942,N_11924);
nor U12062 (N_12062,N_11885,N_11949);
xor U12063 (N_12063,N_11992,N_11981);
and U12064 (N_12064,N_11998,N_11828);
and U12065 (N_12065,N_11858,N_11830);
nor U12066 (N_12066,N_11874,N_11851);
xor U12067 (N_12067,N_11802,N_11915);
nor U12068 (N_12068,N_11876,N_11836);
nand U12069 (N_12069,N_11927,N_11907);
xor U12070 (N_12070,N_11926,N_11824);
nor U12071 (N_12071,N_11841,N_11875);
or U12072 (N_12072,N_11857,N_11894);
and U12073 (N_12073,N_11968,N_11982);
nand U12074 (N_12074,N_11910,N_11832);
nand U12075 (N_12075,N_11901,N_11882);
xnor U12076 (N_12076,N_11811,N_11861);
nand U12077 (N_12077,N_11818,N_11977);
nand U12078 (N_12078,N_11916,N_11895);
nor U12079 (N_12079,N_11842,N_11804);
nor U12080 (N_12080,N_11833,N_11965);
and U12081 (N_12081,N_11972,N_11854);
and U12082 (N_12082,N_11951,N_11909);
nor U12083 (N_12083,N_11922,N_11847);
xor U12084 (N_12084,N_11826,N_11925);
and U12085 (N_12085,N_11807,N_11813);
nand U12086 (N_12086,N_11994,N_11883);
nor U12087 (N_12087,N_11989,N_11864);
xor U12088 (N_12088,N_11956,N_11889);
or U12089 (N_12089,N_11913,N_11919);
or U12090 (N_12090,N_11835,N_11954);
nor U12091 (N_12091,N_11911,N_11856);
or U12092 (N_12092,N_11865,N_11990);
nand U12093 (N_12093,N_11880,N_11988);
xnor U12094 (N_12094,N_11945,N_11912);
nand U12095 (N_12095,N_11997,N_11946);
or U12096 (N_12096,N_11825,N_11849);
xor U12097 (N_12097,N_11969,N_11943);
nor U12098 (N_12098,N_11808,N_11935);
nor U12099 (N_12099,N_11967,N_11848);
and U12100 (N_12100,N_11808,N_11946);
or U12101 (N_12101,N_11960,N_11992);
and U12102 (N_12102,N_11869,N_11855);
nor U12103 (N_12103,N_11980,N_11956);
nor U12104 (N_12104,N_11849,N_11835);
and U12105 (N_12105,N_11892,N_11980);
or U12106 (N_12106,N_11959,N_11800);
nand U12107 (N_12107,N_11956,N_11906);
or U12108 (N_12108,N_11806,N_11972);
nand U12109 (N_12109,N_11945,N_11854);
xnor U12110 (N_12110,N_11849,N_11988);
nor U12111 (N_12111,N_11918,N_11959);
nor U12112 (N_12112,N_11908,N_11862);
and U12113 (N_12113,N_11808,N_11942);
nand U12114 (N_12114,N_11860,N_11945);
nor U12115 (N_12115,N_11923,N_11917);
nand U12116 (N_12116,N_11822,N_11854);
nand U12117 (N_12117,N_11910,N_11874);
or U12118 (N_12118,N_11931,N_11866);
or U12119 (N_12119,N_11818,N_11814);
nand U12120 (N_12120,N_11962,N_11909);
nand U12121 (N_12121,N_11819,N_11925);
and U12122 (N_12122,N_11922,N_11842);
or U12123 (N_12123,N_11940,N_11984);
xnor U12124 (N_12124,N_11925,N_11864);
nor U12125 (N_12125,N_11821,N_11846);
and U12126 (N_12126,N_11915,N_11934);
nor U12127 (N_12127,N_11834,N_11835);
nand U12128 (N_12128,N_11964,N_11898);
nor U12129 (N_12129,N_11814,N_11802);
xor U12130 (N_12130,N_11956,N_11800);
or U12131 (N_12131,N_11838,N_11935);
nor U12132 (N_12132,N_11800,N_11953);
or U12133 (N_12133,N_11825,N_11873);
xnor U12134 (N_12134,N_11823,N_11854);
nand U12135 (N_12135,N_11851,N_11803);
and U12136 (N_12136,N_11801,N_11893);
xnor U12137 (N_12137,N_11871,N_11964);
nor U12138 (N_12138,N_11860,N_11999);
nor U12139 (N_12139,N_11950,N_11866);
nor U12140 (N_12140,N_11802,N_11866);
nor U12141 (N_12141,N_11962,N_11852);
nand U12142 (N_12142,N_11911,N_11813);
nand U12143 (N_12143,N_11904,N_11880);
nand U12144 (N_12144,N_11844,N_11812);
xnor U12145 (N_12145,N_11893,N_11860);
and U12146 (N_12146,N_11937,N_11992);
nor U12147 (N_12147,N_11970,N_11850);
nor U12148 (N_12148,N_11834,N_11979);
nor U12149 (N_12149,N_11835,N_11897);
xor U12150 (N_12150,N_11886,N_11834);
and U12151 (N_12151,N_11820,N_11949);
nor U12152 (N_12152,N_11899,N_11802);
nor U12153 (N_12153,N_11931,N_11979);
and U12154 (N_12154,N_11827,N_11967);
xor U12155 (N_12155,N_11916,N_11911);
nor U12156 (N_12156,N_11888,N_11863);
xnor U12157 (N_12157,N_11832,N_11846);
xnor U12158 (N_12158,N_11961,N_11845);
and U12159 (N_12159,N_11891,N_11848);
or U12160 (N_12160,N_11896,N_11889);
nor U12161 (N_12161,N_11849,N_11928);
or U12162 (N_12162,N_11804,N_11820);
xor U12163 (N_12163,N_11954,N_11900);
or U12164 (N_12164,N_11824,N_11921);
or U12165 (N_12165,N_11877,N_11955);
or U12166 (N_12166,N_11957,N_11963);
nor U12167 (N_12167,N_11892,N_11868);
nand U12168 (N_12168,N_11941,N_11816);
nand U12169 (N_12169,N_11831,N_11823);
nor U12170 (N_12170,N_11850,N_11936);
or U12171 (N_12171,N_11812,N_11926);
xor U12172 (N_12172,N_11903,N_11872);
nand U12173 (N_12173,N_11933,N_11851);
and U12174 (N_12174,N_11912,N_11903);
and U12175 (N_12175,N_11947,N_11941);
nand U12176 (N_12176,N_11896,N_11918);
nor U12177 (N_12177,N_11877,N_11907);
xor U12178 (N_12178,N_11866,N_11837);
xnor U12179 (N_12179,N_11922,N_11846);
nor U12180 (N_12180,N_11927,N_11887);
nand U12181 (N_12181,N_11954,N_11857);
and U12182 (N_12182,N_11980,N_11989);
or U12183 (N_12183,N_11953,N_11915);
xor U12184 (N_12184,N_11851,N_11804);
and U12185 (N_12185,N_11987,N_11891);
nor U12186 (N_12186,N_11912,N_11839);
nor U12187 (N_12187,N_11911,N_11995);
nor U12188 (N_12188,N_11906,N_11912);
and U12189 (N_12189,N_11932,N_11956);
or U12190 (N_12190,N_11962,N_11817);
nor U12191 (N_12191,N_11947,N_11810);
xnor U12192 (N_12192,N_11866,N_11864);
or U12193 (N_12193,N_11973,N_11929);
xnor U12194 (N_12194,N_11820,N_11840);
and U12195 (N_12195,N_11841,N_11845);
and U12196 (N_12196,N_11922,N_11924);
nor U12197 (N_12197,N_11868,N_11887);
xor U12198 (N_12198,N_11876,N_11806);
xor U12199 (N_12199,N_11832,N_11874);
xor U12200 (N_12200,N_12124,N_12197);
nor U12201 (N_12201,N_12161,N_12152);
and U12202 (N_12202,N_12041,N_12067);
xor U12203 (N_12203,N_12131,N_12142);
nor U12204 (N_12204,N_12149,N_12045);
and U12205 (N_12205,N_12155,N_12125);
nor U12206 (N_12206,N_12174,N_12099);
or U12207 (N_12207,N_12009,N_12052);
or U12208 (N_12208,N_12051,N_12071);
nand U12209 (N_12209,N_12141,N_12169);
nor U12210 (N_12210,N_12111,N_12048);
nor U12211 (N_12211,N_12016,N_12158);
xnor U12212 (N_12212,N_12094,N_12096);
nand U12213 (N_12213,N_12066,N_12098);
xor U12214 (N_12214,N_12157,N_12178);
nand U12215 (N_12215,N_12011,N_12177);
nor U12216 (N_12216,N_12053,N_12187);
nor U12217 (N_12217,N_12018,N_12032);
nor U12218 (N_12218,N_12105,N_12074);
nor U12219 (N_12219,N_12077,N_12181);
nand U12220 (N_12220,N_12024,N_12143);
nand U12221 (N_12221,N_12198,N_12191);
nor U12222 (N_12222,N_12122,N_12021);
or U12223 (N_12223,N_12026,N_12055);
xnor U12224 (N_12224,N_12019,N_12084);
or U12225 (N_12225,N_12138,N_12069);
nand U12226 (N_12226,N_12081,N_12092);
and U12227 (N_12227,N_12164,N_12091);
nor U12228 (N_12228,N_12027,N_12188);
and U12229 (N_12229,N_12190,N_12126);
xor U12230 (N_12230,N_12132,N_12006);
xor U12231 (N_12231,N_12043,N_12054);
or U12232 (N_12232,N_12014,N_12113);
or U12233 (N_12233,N_12022,N_12145);
and U12234 (N_12234,N_12107,N_12037);
nand U12235 (N_12235,N_12086,N_12097);
and U12236 (N_12236,N_12088,N_12015);
and U12237 (N_12237,N_12115,N_12118);
nand U12238 (N_12238,N_12038,N_12108);
nand U12239 (N_12239,N_12001,N_12109);
nor U12240 (N_12240,N_12196,N_12146);
or U12241 (N_12241,N_12072,N_12062);
xnor U12242 (N_12242,N_12139,N_12183);
xnor U12243 (N_12243,N_12112,N_12172);
or U12244 (N_12244,N_12044,N_12080);
nand U12245 (N_12245,N_12083,N_12195);
nor U12246 (N_12246,N_12023,N_12117);
xnor U12247 (N_12247,N_12154,N_12165);
nand U12248 (N_12248,N_12007,N_12156);
or U12249 (N_12249,N_12005,N_12136);
nand U12250 (N_12250,N_12189,N_12159);
or U12251 (N_12251,N_12121,N_12160);
xor U12252 (N_12252,N_12192,N_12153);
and U12253 (N_12253,N_12110,N_12058);
xor U12254 (N_12254,N_12163,N_12076);
or U12255 (N_12255,N_12061,N_12000);
nand U12256 (N_12256,N_12013,N_12025);
xor U12257 (N_12257,N_12167,N_12144);
xnor U12258 (N_12258,N_12137,N_12184);
xor U12259 (N_12259,N_12040,N_12134);
xor U12260 (N_12260,N_12186,N_12150);
nor U12261 (N_12261,N_12180,N_12147);
xnor U12262 (N_12262,N_12176,N_12140);
and U12263 (N_12263,N_12114,N_12070);
xnor U12264 (N_12264,N_12033,N_12085);
nor U12265 (N_12265,N_12101,N_12042);
nor U12266 (N_12266,N_12179,N_12068);
xnor U12267 (N_12267,N_12004,N_12129);
nor U12268 (N_12268,N_12012,N_12028);
or U12269 (N_12269,N_12127,N_12079);
nand U12270 (N_12270,N_12093,N_12103);
nand U12271 (N_12271,N_12166,N_12130);
nand U12272 (N_12272,N_12020,N_12078);
and U12273 (N_12273,N_12135,N_12104);
or U12274 (N_12274,N_12162,N_12119);
and U12275 (N_12275,N_12095,N_12031);
nor U12276 (N_12276,N_12120,N_12010);
nor U12277 (N_12277,N_12123,N_12035);
nor U12278 (N_12278,N_12039,N_12128);
nor U12279 (N_12279,N_12065,N_12170);
nor U12280 (N_12280,N_12182,N_12193);
xor U12281 (N_12281,N_12175,N_12017);
and U12282 (N_12282,N_12056,N_12049);
nand U12283 (N_12283,N_12075,N_12171);
nor U12284 (N_12284,N_12057,N_12064);
or U12285 (N_12285,N_12102,N_12002);
nand U12286 (N_12286,N_12046,N_12030);
and U12287 (N_12287,N_12036,N_12059);
and U12288 (N_12288,N_12090,N_12100);
or U12289 (N_12289,N_12060,N_12047);
nand U12290 (N_12290,N_12133,N_12173);
or U12291 (N_12291,N_12008,N_12087);
nand U12292 (N_12292,N_12106,N_12168);
nand U12293 (N_12293,N_12194,N_12063);
nor U12294 (N_12294,N_12034,N_12082);
and U12295 (N_12295,N_12029,N_12003);
xor U12296 (N_12296,N_12089,N_12148);
nor U12297 (N_12297,N_12185,N_12199);
and U12298 (N_12298,N_12151,N_12073);
nand U12299 (N_12299,N_12050,N_12116);
nor U12300 (N_12300,N_12093,N_12062);
xnor U12301 (N_12301,N_12143,N_12170);
nand U12302 (N_12302,N_12123,N_12006);
nand U12303 (N_12303,N_12010,N_12047);
and U12304 (N_12304,N_12057,N_12178);
xor U12305 (N_12305,N_12168,N_12062);
or U12306 (N_12306,N_12059,N_12046);
nor U12307 (N_12307,N_12025,N_12007);
or U12308 (N_12308,N_12181,N_12197);
xnor U12309 (N_12309,N_12118,N_12059);
or U12310 (N_12310,N_12180,N_12082);
nand U12311 (N_12311,N_12187,N_12086);
xor U12312 (N_12312,N_12007,N_12033);
xnor U12313 (N_12313,N_12081,N_12006);
xor U12314 (N_12314,N_12011,N_12055);
xor U12315 (N_12315,N_12071,N_12138);
nand U12316 (N_12316,N_12033,N_12101);
and U12317 (N_12317,N_12130,N_12039);
xor U12318 (N_12318,N_12043,N_12156);
and U12319 (N_12319,N_12076,N_12169);
nand U12320 (N_12320,N_12089,N_12077);
or U12321 (N_12321,N_12017,N_12159);
xor U12322 (N_12322,N_12133,N_12186);
xnor U12323 (N_12323,N_12098,N_12030);
nor U12324 (N_12324,N_12061,N_12087);
or U12325 (N_12325,N_12099,N_12006);
nand U12326 (N_12326,N_12031,N_12109);
nor U12327 (N_12327,N_12075,N_12162);
xnor U12328 (N_12328,N_12133,N_12128);
nor U12329 (N_12329,N_12163,N_12156);
and U12330 (N_12330,N_12009,N_12182);
nand U12331 (N_12331,N_12021,N_12127);
and U12332 (N_12332,N_12117,N_12173);
xor U12333 (N_12333,N_12039,N_12162);
xnor U12334 (N_12334,N_12099,N_12129);
nand U12335 (N_12335,N_12155,N_12009);
nor U12336 (N_12336,N_12194,N_12031);
nor U12337 (N_12337,N_12026,N_12037);
or U12338 (N_12338,N_12013,N_12130);
and U12339 (N_12339,N_12143,N_12102);
or U12340 (N_12340,N_12170,N_12097);
and U12341 (N_12341,N_12032,N_12190);
xor U12342 (N_12342,N_12019,N_12016);
xor U12343 (N_12343,N_12021,N_12171);
xnor U12344 (N_12344,N_12040,N_12100);
or U12345 (N_12345,N_12125,N_12152);
or U12346 (N_12346,N_12192,N_12118);
and U12347 (N_12347,N_12039,N_12097);
xnor U12348 (N_12348,N_12073,N_12098);
or U12349 (N_12349,N_12189,N_12090);
xnor U12350 (N_12350,N_12034,N_12022);
xnor U12351 (N_12351,N_12137,N_12064);
and U12352 (N_12352,N_12023,N_12112);
or U12353 (N_12353,N_12191,N_12017);
nand U12354 (N_12354,N_12010,N_12035);
and U12355 (N_12355,N_12084,N_12044);
xnor U12356 (N_12356,N_12065,N_12000);
nor U12357 (N_12357,N_12042,N_12029);
xnor U12358 (N_12358,N_12117,N_12009);
and U12359 (N_12359,N_12097,N_12053);
nor U12360 (N_12360,N_12158,N_12166);
nand U12361 (N_12361,N_12086,N_12107);
and U12362 (N_12362,N_12076,N_12111);
xnor U12363 (N_12363,N_12171,N_12066);
nor U12364 (N_12364,N_12178,N_12027);
nor U12365 (N_12365,N_12041,N_12068);
or U12366 (N_12366,N_12085,N_12064);
and U12367 (N_12367,N_12117,N_12129);
and U12368 (N_12368,N_12180,N_12126);
nand U12369 (N_12369,N_12187,N_12074);
nand U12370 (N_12370,N_12182,N_12021);
xor U12371 (N_12371,N_12036,N_12077);
and U12372 (N_12372,N_12189,N_12061);
nand U12373 (N_12373,N_12129,N_12105);
xor U12374 (N_12374,N_12044,N_12112);
or U12375 (N_12375,N_12167,N_12084);
xor U12376 (N_12376,N_12015,N_12151);
or U12377 (N_12377,N_12078,N_12126);
and U12378 (N_12378,N_12088,N_12086);
xnor U12379 (N_12379,N_12160,N_12104);
nor U12380 (N_12380,N_12093,N_12127);
nand U12381 (N_12381,N_12181,N_12107);
nand U12382 (N_12382,N_12111,N_12023);
and U12383 (N_12383,N_12081,N_12047);
nor U12384 (N_12384,N_12049,N_12062);
or U12385 (N_12385,N_12069,N_12159);
or U12386 (N_12386,N_12170,N_12072);
and U12387 (N_12387,N_12166,N_12046);
nand U12388 (N_12388,N_12127,N_12124);
and U12389 (N_12389,N_12156,N_12033);
nand U12390 (N_12390,N_12172,N_12187);
xnor U12391 (N_12391,N_12191,N_12149);
or U12392 (N_12392,N_12145,N_12081);
or U12393 (N_12393,N_12106,N_12007);
nand U12394 (N_12394,N_12181,N_12073);
nor U12395 (N_12395,N_12178,N_12153);
nand U12396 (N_12396,N_12108,N_12182);
and U12397 (N_12397,N_12189,N_12166);
nand U12398 (N_12398,N_12172,N_12175);
nor U12399 (N_12399,N_12193,N_12102);
nor U12400 (N_12400,N_12354,N_12272);
nand U12401 (N_12401,N_12204,N_12359);
or U12402 (N_12402,N_12238,N_12301);
nor U12403 (N_12403,N_12207,N_12235);
or U12404 (N_12404,N_12266,N_12399);
and U12405 (N_12405,N_12335,N_12268);
xor U12406 (N_12406,N_12377,N_12270);
nor U12407 (N_12407,N_12275,N_12228);
or U12408 (N_12408,N_12362,N_12345);
xnor U12409 (N_12409,N_12251,N_12325);
or U12410 (N_12410,N_12358,N_12216);
nor U12411 (N_12411,N_12302,N_12245);
nor U12412 (N_12412,N_12203,N_12348);
nand U12413 (N_12413,N_12291,N_12289);
xnor U12414 (N_12414,N_12384,N_12338);
xnor U12415 (N_12415,N_12392,N_12208);
nor U12416 (N_12416,N_12264,N_12282);
nor U12417 (N_12417,N_12363,N_12274);
nand U12418 (N_12418,N_12393,N_12379);
nor U12419 (N_12419,N_12336,N_12319);
nand U12420 (N_12420,N_12278,N_12202);
nand U12421 (N_12421,N_12323,N_12372);
nor U12422 (N_12422,N_12322,N_12257);
xnor U12423 (N_12423,N_12394,N_12220);
or U12424 (N_12424,N_12351,N_12263);
xor U12425 (N_12425,N_12217,N_12284);
xor U12426 (N_12426,N_12373,N_12305);
nand U12427 (N_12427,N_12380,N_12389);
nand U12428 (N_12428,N_12261,N_12339);
nand U12429 (N_12429,N_12365,N_12306);
or U12430 (N_12430,N_12360,N_12246);
nand U12431 (N_12431,N_12293,N_12382);
and U12432 (N_12432,N_12213,N_12340);
xnor U12433 (N_12433,N_12386,N_12314);
nor U12434 (N_12434,N_12313,N_12371);
and U12435 (N_12435,N_12288,N_12375);
nand U12436 (N_12436,N_12299,N_12308);
nand U12437 (N_12437,N_12317,N_12328);
or U12438 (N_12438,N_12397,N_12256);
xor U12439 (N_12439,N_12396,N_12254);
nor U12440 (N_12440,N_12296,N_12349);
nand U12441 (N_12441,N_12240,N_12234);
and U12442 (N_12442,N_12242,N_12295);
xnor U12443 (N_12443,N_12347,N_12364);
nor U12444 (N_12444,N_12330,N_12241);
nor U12445 (N_12445,N_12267,N_12233);
nand U12446 (N_12446,N_12292,N_12294);
nor U12447 (N_12447,N_12329,N_12285);
and U12448 (N_12448,N_12260,N_12366);
or U12449 (N_12449,N_12258,N_12269);
nand U12450 (N_12450,N_12237,N_12200);
or U12451 (N_12451,N_12212,N_12318);
nor U12452 (N_12452,N_12381,N_12350);
xor U12453 (N_12453,N_12370,N_12279);
nor U12454 (N_12454,N_12385,N_12290);
nand U12455 (N_12455,N_12367,N_12355);
and U12456 (N_12456,N_12337,N_12315);
nor U12457 (N_12457,N_12300,N_12250);
or U12458 (N_12458,N_12346,N_12222);
and U12459 (N_12459,N_12230,N_12227);
or U12460 (N_12460,N_12221,N_12206);
and U12461 (N_12461,N_12320,N_12297);
xnor U12462 (N_12462,N_12368,N_12312);
nor U12463 (N_12463,N_12215,N_12333);
nor U12464 (N_12464,N_12210,N_12259);
xor U12465 (N_12465,N_12225,N_12253);
nor U12466 (N_12466,N_12304,N_12209);
xnor U12467 (N_12467,N_12342,N_12214);
nor U12468 (N_12468,N_12310,N_12262);
or U12469 (N_12469,N_12249,N_12369);
and U12470 (N_12470,N_12353,N_12356);
and U12471 (N_12471,N_12218,N_12280);
nor U12472 (N_12472,N_12224,N_12316);
and U12473 (N_12473,N_12307,N_12229);
nand U12474 (N_12474,N_12331,N_12239);
nand U12475 (N_12475,N_12391,N_12276);
nor U12476 (N_12476,N_12281,N_12376);
and U12477 (N_12477,N_12341,N_12243);
or U12478 (N_12478,N_12326,N_12309);
xnor U12479 (N_12479,N_12286,N_12223);
or U12480 (N_12480,N_12357,N_12219);
xnor U12481 (N_12481,N_12378,N_12387);
or U12482 (N_12482,N_12374,N_12205);
xnor U12483 (N_12483,N_12324,N_12252);
xor U12484 (N_12484,N_12332,N_12248);
nor U12485 (N_12485,N_12273,N_12287);
and U12486 (N_12486,N_12231,N_12352);
and U12487 (N_12487,N_12236,N_12211);
xor U12488 (N_12488,N_12247,N_12361);
nor U12489 (N_12489,N_12383,N_12298);
nor U12490 (N_12490,N_12334,N_12321);
and U12491 (N_12491,N_12390,N_12277);
and U12492 (N_12492,N_12344,N_12244);
nand U12493 (N_12493,N_12255,N_12388);
nor U12494 (N_12494,N_12265,N_12395);
or U12495 (N_12495,N_12327,N_12226);
xor U12496 (N_12496,N_12311,N_12232);
and U12497 (N_12497,N_12343,N_12271);
or U12498 (N_12498,N_12303,N_12398);
nand U12499 (N_12499,N_12201,N_12283);
xnor U12500 (N_12500,N_12382,N_12383);
or U12501 (N_12501,N_12225,N_12245);
nand U12502 (N_12502,N_12221,N_12327);
or U12503 (N_12503,N_12383,N_12341);
nor U12504 (N_12504,N_12300,N_12253);
nand U12505 (N_12505,N_12306,N_12282);
or U12506 (N_12506,N_12328,N_12308);
or U12507 (N_12507,N_12394,N_12358);
nor U12508 (N_12508,N_12365,N_12252);
xor U12509 (N_12509,N_12396,N_12397);
and U12510 (N_12510,N_12206,N_12375);
nand U12511 (N_12511,N_12336,N_12280);
nand U12512 (N_12512,N_12293,N_12330);
nor U12513 (N_12513,N_12207,N_12301);
or U12514 (N_12514,N_12372,N_12302);
or U12515 (N_12515,N_12224,N_12308);
or U12516 (N_12516,N_12274,N_12207);
nor U12517 (N_12517,N_12392,N_12399);
and U12518 (N_12518,N_12386,N_12344);
nor U12519 (N_12519,N_12360,N_12272);
or U12520 (N_12520,N_12229,N_12258);
nor U12521 (N_12521,N_12364,N_12235);
nor U12522 (N_12522,N_12378,N_12291);
and U12523 (N_12523,N_12386,N_12371);
nand U12524 (N_12524,N_12230,N_12317);
nand U12525 (N_12525,N_12259,N_12204);
xnor U12526 (N_12526,N_12270,N_12325);
or U12527 (N_12527,N_12253,N_12335);
nand U12528 (N_12528,N_12228,N_12255);
or U12529 (N_12529,N_12320,N_12200);
and U12530 (N_12530,N_12326,N_12358);
nor U12531 (N_12531,N_12379,N_12367);
xor U12532 (N_12532,N_12221,N_12227);
nor U12533 (N_12533,N_12308,N_12234);
nor U12534 (N_12534,N_12289,N_12230);
nand U12535 (N_12535,N_12355,N_12390);
xor U12536 (N_12536,N_12338,N_12368);
or U12537 (N_12537,N_12398,N_12352);
xnor U12538 (N_12538,N_12340,N_12216);
and U12539 (N_12539,N_12323,N_12222);
or U12540 (N_12540,N_12291,N_12318);
xnor U12541 (N_12541,N_12269,N_12321);
and U12542 (N_12542,N_12291,N_12205);
nor U12543 (N_12543,N_12211,N_12362);
and U12544 (N_12544,N_12354,N_12303);
nor U12545 (N_12545,N_12301,N_12259);
xor U12546 (N_12546,N_12323,N_12213);
and U12547 (N_12547,N_12300,N_12230);
xor U12548 (N_12548,N_12279,N_12360);
nand U12549 (N_12549,N_12203,N_12367);
and U12550 (N_12550,N_12309,N_12263);
or U12551 (N_12551,N_12288,N_12280);
or U12552 (N_12552,N_12205,N_12222);
nand U12553 (N_12553,N_12314,N_12216);
nor U12554 (N_12554,N_12316,N_12382);
and U12555 (N_12555,N_12302,N_12398);
or U12556 (N_12556,N_12236,N_12207);
and U12557 (N_12557,N_12218,N_12361);
nand U12558 (N_12558,N_12371,N_12253);
xor U12559 (N_12559,N_12349,N_12267);
or U12560 (N_12560,N_12327,N_12262);
or U12561 (N_12561,N_12296,N_12258);
and U12562 (N_12562,N_12230,N_12314);
or U12563 (N_12563,N_12339,N_12381);
xnor U12564 (N_12564,N_12358,N_12364);
or U12565 (N_12565,N_12208,N_12329);
xnor U12566 (N_12566,N_12330,N_12215);
nand U12567 (N_12567,N_12356,N_12262);
nand U12568 (N_12568,N_12306,N_12317);
nor U12569 (N_12569,N_12384,N_12254);
xor U12570 (N_12570,N_12314,N_12347);
nand U12571 (N_12571,N_12204,N_12334);
and U12572 (N_12572,N_12288,N_12385);
xnor U12573 (N_12573,N_12226,N_12261);
and U12574 (N_12574,N_12355,N_12308);
nor U12575 (N_12575,N_12341,N_12302);
nand U12576 (N_12576,N_12366,N_12262);
nand U12577 (N_12577,N_12262,N_12344);
nor U12578 (N_12578,N_12302,N_12390);
or U12579 (N_12579,N_12321,N_12387);
xor U12580 (N_12580,N_12203,N_12379);
xnor U12581 (N_12581,N_12390,N_12213);
nand U12582 (N_12582,N_12322,N_12369);
nor U12583 (N_12583,N_12260,N_12213);
xnor U12584 (N_12584,N_12266,N_12346);
and U12585 (N_12585,N_12232,N_12397);
and U12586 (N_12586,N_12390,N_12397);
or U12587 (N_12587,N_12296,N_12206);
nand U12588 (N_12588,N_12354,N_12301);
nor U12589 (N_12589,N_12243,N_12393);
and U12590 (N_12590,N_12307,N_12357);
or U12591 (N_12591,N_12358,N_12275);
or U12592 (N_12592,N_12352,N_12228);
and U12593 (N_12593,N_12255,N_12270);
and U12594 (N_12594,N_12332,N_12301);
or U12595 (N_12595,N_12241,N_12309);
xnor U12596 (N_12596,N_12203,N_12374);
and U12597 (N_12597,N_12342,N_12298);
and U12598 (N_12598,N_12301,N_12348);
or U12599 (N_12599,N_12384,N_12223);
nor U12600 (N_12600,N_12562,N_12410);
nand U12601 (N_12601,N_12574,N_12435);
nor U12602 (N_12602,N_12498,N_12587);
or U12603 (N_12603,N_12465,N_12523);
or U12604 (N_12604,N_12489,N_12490);
nor U12605 (N_12605,N_12597,N_12566);
xnor U12606 (N_12606,N_12484,N_12516);
nor U12607 (N_12607,N_12553,N_12423);
or U12608 (N_12608,N_12470,N_12416);
xnor U12609 (N_12609,N_12459,N_12411);
or U12610 (N_12610,N_12431,N_12573);
xnor U12611 (N_12611,N_12437,N_12598);
and U12612 (N_12612,N_12544,N_12430);
xnor U12613 (N_12613,N_12527,N_12590);
or U12614 (N_12614,N_12591,N_12549);
nand U12615 (N_12615,N_12578,N_12452);
or U12616 (N_12616,N_12589,N_12506);
xor U12617 (N_12617,N_12412,N_12570);
or U12618 (N_12618,N_12497,N_12482);
and U12619 (N_12619,N_12480,N_12584);
nor U12620 (N_12620,N_12466,N_12560);
xnor U12621 (N_12621,N_12415,N_12406);
and U12622 (N_12622,N_12467,N_12426);
or U12623 (N_12623,N_12534,N_12531);
nand U12624 (N_12624,N_12402,N_12515);
and U12625 (N_12625,N_12505,N_12583);
and U12626 (N_12626,N_12520,N_12502);
nand U12627 (N_12627,N_12407,N_12433);
nand U12628 (N_12628,N_12593,N_12456);
nand U12629 (N_12629,N_12447,N_12414);
nand U12630 (N_12630,N_12567,N_12448);
or U12631 (N_12631,N_12585,N_12472);
xor U12632 (N_12632,N_12454,N_12540);
xnor U12633 (N_12633,N_12577,N_12417);
or U12634 (N_12634,N_12438,N_12599);
nand U12635 (N_12635,N_12401,N_12537);
nand U12636 (N_12636,N_12538,N_12439);
xor U12637 (N_12637,N_12461,N_12477);
nor U12638 (N_12638,N_12425,N_12463);
nand U12639 (N_12639,N_12525,N_12441);
and U12640 (N_12640,N_12428,N_12487);
and U12641 (N_12641,N_12494,N_12404);
or U12642 (N_12642,N_12582,N_12485);
and U12643 (N_12643,N_12403,N_12413);
and U12644 (N_12644,N_12408,N_12517);
or U12645 (N_12645,N_12548,N_12444);
and U12646 (N_12646,N_12491,N_12405);
or U12647 (N_12647,N_12521,N_12501);
nand U12648 (N_12648,N_12530,N_12507);
xor U12649 (N_12649,N_12453,N_12471);
xor U12650 (N_12650,N_12564,N_12421);
xor U12651 (N_12651,N_12592,N_12440);
nand U12652 (N_12652,N_12568,N_12518);
or U12653 (N_12653,N_12478,N_12561);
nand U12654 (N_12654,N_12541,N_12446);
nand U12655 (N_12655,N_12569,N_12565);
nor U12656 (N_12656,N_12576,N_12547);
and U12657 (N_12657,N_12422,N_12535);
nand U12658 (N_12658,N_12594,N_12432);
or U12659 (N_12659,N_12409,N_12500);
and U12660 (N_12660,N_12575,N_12419);
nor U12661 (N_12661,N_12512,N_12558);
nor U12662 (N_12662,N_12526,N_12563);
and U12663 (N_12663,N_12481,N_12418);
and U12664 (N_12664,N_12474,N_12479);
nor U12665 (N_12665,N_12503,N_12588);
nand U12666 (N_12666,N_12464,N_12468);
or U12667 (N_12667,N_12429,N_12495);
and U12668 (N_12668,N_12460,N_12522);
and U12669 (N_12669,N_12473,N_12427);
xor U12670 (N_12670,N_12509,N_12551);
and U12671 (N_12671,N_12499,N_12571);
nand U12672 (N_12672,N_12436,N_12488);
nor U12673 (N_12673,N_12508,N_12443);
nor U12674 (N_12674,N_12524,N_12442);
nand U12675 (N_12675,N_12559,N_12476);
nand U12676 (N_12676,N_12533,N_12511);
nand U12677 (N_12677,N_12586,N_12581);
xnor U12678 (N_12678,N_12492,N_12557);
nand U12679 (N_12679,N_12539,N_12545);
nand U12680 (N_12680,N_12457,N_12543);
nand U12681 (N_12681,N_12572,N_12554);
xor U12682 (N_12682,N_12552,N_12400);
nor U12683 (N_12683,N_12536,N_12510);
or U12684 (N_12684,N_12424,N_12434);
xor U12685 (N_12685,N_12596,N_12580);
and U12686 (N_12686,N_12519,N_12532);
and U12687 (N_12687,N_12451,N_12462);
nand U12688 (N_12688,N_12542,N_12496);
xor U12689 (N_12689,N_12513,N_12555);
and U12690 (N_12690,N_12475,N_12550);
or U12691 (N_12691,N_12579,N_12420);
or U12692 (N_12692,N_12450,N_12469);
nand U12693 (N_12693,N_12445,N_12528);
xnor U12694 (N_12694,N_12483,N_12529);
nand U12695 (N_12695,N_12458,N_12449);
or U12696 (N_12696,N_12504,N_12455);
and U12697 (N_12697,N_12595,N_12486);
or U12698 (N_12698,N_12546,N_12514);
nor U12699 (N_12699,N_12556,N_12493);
nand U12700 (N_12700,N_12558,N_12509);
nor U12701 (N_12701,N_12419,N_12544);
xor U12702 (N_12702,N_12459,N_12574);
and U12703 (N_12703,N_12501,N_12484);
and U12704 (N_12704,N_12505,N_12542);
xnor U12705 (N_12705,N_12583,N_12551);
nor U12706 (N_12706,N_12582,N_12461);
and U12707 (N_12707,N_12557,N_12501);
or U12708 (N_12708,N_12539,N_12468);
and U12709 (N_12709,N_12434,N_12406);
nand U12710 (N_12710,N_12570,N_12400);
xor U12711 (N_12711,N_12561,N_12557);
or U12712 (N_12712,N_12587,N_12516);
xnor U12713 (N_12713,N_12427,N_12413);
nor U12714 (N_12714,N_12513,N_12563);
nor U12715 (N_12715,N_12423,N_12566);
nand U12716 (N_12716,N_12485,N_12415);
or U12717 (N_12717,N_12430,N_12509);
or U12718 (N_12718,N_12594,N_12458);
or U12719 (N_12719,N_12569,N_12548);
and U12720 (N_12720,N_12583,N_12578);
and U12721 (N_12721,N_12537,N_12400);
and U12722 (N_12722,N_12446,N_12512);
nor U12723 (N_12723,N_12443,N_12528);
and U12724 (N_12724,N_12580,N_12552);
or U12725 (N_12725,N_12556,N_12462);
or U12726 (N_12726,N_12520,N_12403);
xor U12727 (N_12727,N_12440,N_12468);
or U12728 (N_12728,N_12426,N_12499);
and U12729 (N_12729,N_12572,N_12579);
nand U12730 (N_12730,N_12504,N_12588);
or U12731 (N_12731,N_12418,N_12431);
nor U12732 (N_12732,N_12553,N_12532);
nand U12733 (N_12733,N_12551,N_12580);
and U12734 (N_12734,N_12505,N_12489);
nand U12735 (N_12735,N_12521,N_12495);
nor U12736 (N_12736,N_12483,N_12513);
or U12737 (N_12737,N_12432,N_12546);
nand U12738 (N_12738,N_12524,N_12525);
and U12739 (N_12739,N_12495,N_12415);
xnor U12740 (N_12740,N_12426,N_12561);
xnor U12741 (N_12741,N_12491,N_12555);
and U12742 (N_12742,N_12528,N_12420);
nor U12743 (N_12743,N_12516,N_12439);
nor U12744 (N_12744,N_12525,N_12545);
nor U12745 (N_12745,N_12496,N_12441);
and U12746 (N_12746,N_12522,N_12484);
nor U12747 (N_12747,N_12424,N_12557);
or U12748 (N_12748,N_12592,N_12464);
and U12749 (N_12749,N_12548,N_12563);
or U12750 (N_12750,N_12465,N_12405);
nor U12751 (N_12751,N_12480,N_12540);
and U12752 (N_12752,N_12402,N_12494);
and U12753 (N_12753,N_12445,N_12422);
nand U12754 (N_12754,N_12407,N_12589);
nand U12755 (N_12755,N_12456,N_12400);
nand U12756 (N_12756,N_12438,N_12592);
xor U12757 (N_12757,N_12428,N_12503);
nand U12758 (N_12758,N_12422,N_12460);
nor U12759 (N_12759,N_12422,N_12457);
and U12760 (N_12760,N_12438,N_12589);
or U12761 (N_12761,N_12439,N_12466);
or U12762 (N_12762,N_12583,N_12594);
nand U12763 (N_12763,N_12417,N_12488);
xnor U12764 (N_12764,N_12470,N_12404);
and U12765 (N_12765,N_12588,N_12595);
nand U12766 (N_12766,N_12524,N_12544);
or U12767 (N_12767,N_12591,N_12543);
or U12768 (N_12768,N_12460,N_12537);
nor U12769 (N_12769,N_12551,N_12494);
or U12770 (N_12770,N_12427,N_12518);
nand U12771 (N_12771,N_12505,N_12517);
and U12772 (N_12772,N_12577,N_12430);
or U12773 (N_12773,N_12423,N_12448);
or U12774 (N_12774,N_12527,N_12413);
nor U12775 (N_12775,N_12583,N_12431);
xor U12776 (N_12776,N_12406,N_12509);
nor U12777 (N_12777,N_12517,N_12598);
nand U12778 (N_12778,N_12418,N_12538);
and U12779 (N_12779,N_12481,N_12507);
nand U12780 (N_12780,N_12457,N_12592);
xor U12781 (N_12781,N_12539,N_12536);
nor U12782 (N_12782,N_12495,N_12517);
and U12783 (N_12783,N_12452,N_12529);
and U12784 (N_12784,N_12520,N_12555);
and U12785 (N_12785,N_12589,N_12459);
xnor U12786 (N_12786,N_12414,N_12412);
nor U12787 (N_12787,N_12578,N_12594);
and U12788 (N_12788,N_12527,N_12542);
xnor U12789 (N_12789,N_12507,N_12420);
nand U12790 (N_12790,N_12495,N_12448);
or U12791 (N_12791,N_12486,N_12557);
or U12792 (N_12792,N_12513,N_12413);
nand U12793 (N_12793,N_12445,N_12482);
and U12794 (N_12794,N_12592,N_12551);
or U12795 (N_12795,N_12589,N_12449);
or U12796 (N_12796,N_12491,N_12470);
or U12797 (N_12797,N_12426,N_12595);
or U12798 (N_12798,N_12557,N_12562);
nand U12799 (N_12799,N_12517,N_12473);
and U12800 (N_12800,N_12705,N_12600);
xnor U12801 (N_12801,N_12749,N_12743);
nand U12802 (N_12802,N_12748,N_12653);
or U12803 (N_12803,N_12737,N_12777);
nand U12804 (N_12804,N_12753,N_12784);
and U12805 (N_12805,N_12747,N_12712);
xor U12806 (N_12806,N_12742,N_12615);
and U12807 (N_12807,N_12739,N_12799);
or U12808 (N_12808,N_12625,N_12720);
xnor U12809 (N_12809,N_12762,N_12710);
nor U12810 (N_12810,N_12763,N_12666);
nor U12811 (N_12811,N_12668,N_12791);
nand U12812 (N_12812,N_12620,N_12651);
nand U12813 (N_12813,N_12682,N_12679);
nor U12814 (N_12814,N_12709,N_12632);
or U12815 (N_12815,N_12684,N_12797);
nand U12816 (N_12816,N_12771,N_12675);
and U12817 (N_12817,N_12733,N_12781);
and U12818 (N_12818,N_12678,N_12783);
xor U12819 (N_12819,N_12779,N_12736);
xor U12820 (N_12820,N_12792,N_12640);
xor U12821 (N_12821,N_12772,N_12745);
and U12822 (N_12822,N_12631,N_12760);
and U12823 (N_12823,N_12662,N_12647);
nand U12824 (N_12824,N_12674,N_12624);
or U12825 (N_12825,N_12611,N_12627);
xor U12826 (N_12826,N_12732,N_12610);
xnor U12827 (N_12827,N_12605,N_12708);
nand U12828 (N_12828,N_12667,N_12612);
or U12829 (N_12829,N_12603,N_12622);
xnor U12830 (N_12830,N_12721,N_12673);
nor U12831 (N_12831,N_12774,N_12764);
and U12832 (N_12832,N_12706,N_12656);
nor U12833 (N_12833,N_12703,N_12769);
nor U12834 (N_12834,N_12601,N_12717);
nor U12835 (N_12835,N_12614,N_12677);
nor U12836 (N_12836,N_12759,N_12741);
nor U12837 (N_12837,N_12634,N_12643);
nand U12838 (N_12838,N_12724,N_12685);
xor U12839 (N_12839,N_12711,N_12609);
nor U12840 (N_12840,N_12722,N_12793);
nor U12841 (N_12841,N_12676,N_12746);
xnor U12842 (N_12842,N_12695,N_12617);
xnor U12843 (N_12843,N_12637,N_12790);
or U12844 (N_12844,N_12649,N_12786);
and U12845 (N_12845,N_12796,N_12725);
or U12846 (N_12846,N_12744,N_12604);
xor U12847 (N_12847,N_12715,N_12602);
nand U12848 (N_12848,N_12768,N_12702);
nor U12849 (N_12849,N_12765,N_12619);
or U12850 (N_12850,N_12635,N_12692);
xor U12851 (N_12851,N_12767,N_12645);
nand U12852 (N_12852,N_12795,N_12650);
nor U12853 (N_12853,N_12727,N_12654);
and U12854 (N_12854,N_12752,N_12633);
and U12855 (N_12855,N_12730,N_12608);
and U12856 (N_12856,N_12670,N_12776);
or U12857 (N_12857,N_12680,N_12778);
xor U12858 (N_12858,N_12754,N_12658);
or U12859 (N_12859,N_12788,N_12655);
or U12860 (N_12860,N_12735,N_12638);
nor U12861 (N_12861,N_12636,N_12694);
and U12862 (N_12862,N_12738,N_12704);
or U12863 (N_12863,N_12785,N_12689);
nor U12864 (N_12864,N_12623,N_12621);
xor U12865 (N_12865,N_12669,N_12755);
xnor U12866 (N_12866,N_12629,N_12787);
nor U12867 (N_12867,N_12750,N_12780);
nor U12868 (N_12868,N_12686,N_12690);
xor U12869 (N_12869,N_12726,N_12657);
nand U12870 (N_12870,N_12626,N_12719);
nand U12871 (N_12871,N_12616,N_12699);
xnor U12872 (N_12872,N_12697,N_12641);
xnor U12873 (N_12873,N_12683,N_12652);
and U12874 (N_12874,N_12664,N_12770);
and U12875 (N_12875,N_12701,N_12663);
nor U12876 (N_12876,N_12713,N_12659);
nand U12877 (N_12877,N_12639,N_12698);
or U12878 (N_12878,N_12798,N_12731);
nor U12879 (N_12879,N_12648,N_12606);
nand U12880 (N_12880,N_12734,N_12723);
nor U12881 (N_12881,N_12671,N_12672);
and U12882 (N_12882,N_12618,N_12789);
and U12883 (N_12883,N_12716,N_12714);
and U12884 (N_12884,N_12729,N_12740);
nor U12885 (N_12885,N_12660,N_12758);
xnor U12886 (N_12886,N_12756,N_12681);
and U12887 (N_12887,N_12687,N_12718);
nor U12888 (N_12888,N_12700,N_12628);
nand U12889 (N_12889,N_12696,N_12775);
nand U12890 (N_12890,N_12661,N_12794);
nand U12891 (N_12891,N_12691,N_12707);
nand U12892 (N_12892,N_12613,N_12761);
nor U12893 (N_12893,N_12665,N_12693);
or U12894 (N_12894,N_12728,N_12642);
and U12895 (N_12895,N_12766,N_12757);
xnor U12896 (N_12896,N_12607,N_12751);
or U12897 (N_12897,N_12773,N_12646);
and U12898 (N_12898,N_12688,N_12644);
and U12899 (N_12899,N_12782,N_12630);
or U12900 (N_12900,N_12605,N_12702);
nand U12901 (N_12901,N_12655,N_12714);
or U12902 (N_12902,N_12738,N_12606);
nor U12903 (N_12903,N_12602,N_12769);
or U12904 (N_12904,N_12680,N_12638);
xor U12905 (N_12905,N_12723,N_12729);
or U12906 (N_12906,N_12674,N_12796);
nor U12907 (N_12907,N_12690,N_12739);
or U12908 (N_12908,N_12740,N_12634);
or U12909 (N_12909,N_12677,N_12648);
and U12910 (N_12910,N_12643,N_12699);
nor U12911 (N_12911,N_12759,N_12648);
and U12912 (N_12912,N_12747,N_12650);
xor U12913 (N_12913,N_12605,N_12631);
nor U12914 (N_12914,N_12772,N_12760);
nand U12915 (N_12915,N_12700,N_12621);
nor U12916 (N_12916,N_12729,N_12638);
and U12917 (N_12917,N_12791,N_12786);
or U12918 (N_12918,N_12763,N_12719);
nor U12919 (N_12919,N_12722,N_12737);
xor U12920 (N_12920,N_12628,N_12680);
or U12921 (N_12921,N_12786,N_12713);
nor U12922 (N_12922,N_12651,N_12715);
nand U12923 (N_12923,N_12605,N_12668);
nand U12924 (N_12924,N_12752,N_12746);
nor U12925 (N_12925,N_12701,N_12748);
xor U12926 (N_12926,N_12680,N_12652);
xnor U12927 (N_12927,N_12774,N_12742);
nand U12928 (N_12928,N_12637,N_12632);
nand U12929 (N_12929,N_12649,N_12787);
and U12930 (N_12930,N_12787,N_12707);
nor U12931 (N_12931,N_12762,N_12652);
nand U12932 (N_12932,N_12642,N_12614);
and U12933 (N_12933,N_12758,N_12647);
nor U12934 (N_12934,N_12713,N_12770);
and U12935 (N_12935,N_12651,N_12606);
and U12936 (N_12936,N_12609,N_12656);
nor U12937 (N_12937,N_12769,N_12675);
xnor U12938 (N_12938,N_12760,N_12710);
and U12939 (N_12939,N_12720,N_12600);
xor U12940 (N_12940,N_12775,N_12782);
or U12941 (N_12941,N_12723,N_12743);
nor U12942 (N_12942,N_12702,N_12769);
nor U12943 (N_12943,N_12626,N_12715);
xor U12944 (N_12944,N_12716,N_12751);
nand U12945 (N_12945,N_12604,N_12702);
xor U12946 (N_12946,N_12773,N_12788);
nand U12947 (N_12947,N_12672,N_12724);
nand U12948 (N_12948,N_12696,N_12680);
xnor U12949 (N_12949,N_12769,N_12721);
nand U12950 (N_12950,N_12686,N_12668);
nand U12951 (N_12951,N_12790,N_12656);
xor U12952 (N_12952,N_12605,N_12690);
and U12953 (N_12953,N_12741,N_12736);
nor U12954 (N_12954,N_12649,N_12662);
and U12955 (N_12955,N_12765,N_12754);
nand U12956 (N_12956,N_12734,N_12629);
xor U12957 (N_12957,N_12604,N_12725);
nor U12958 (N_12958,N_12601,N_12640);
nand U12959 (N_12959,N_12614,N_12780);
and U12960 (N_12960,N_12746,N_12744);
nor U12961 (N_12961,N_12608,N_12766);
xnor U12962 (N_12962,N_12703,N_12660);
xor U12963 (N_12963,N_12761,N_12707);
and U12964 (N_12964,N_12746,N_12718);
and U12965 (N_12965,N_12718,N_12607);
and U12966 (N_12966,N_12617,N_12653);
and U12967 (N_12967,N_12739,N_12763);
or U12968 (N_12968,N_12644,N_12664);
and U12969 (N_12969,N_12755,N_12645);
or U12970 (N_12970,N_12604,N_12741);
xnor U12971 (N_12971,N_12660,N_12693);
xor U12972 (N_12972,N_12661,N_12668);
and U12973 (N_12973,N_12784,N_12644);
nand U12974 (N_12974,N_12619,N_12656);
xnor U12975 (N_12975,N_12620,N_12607);
nor U12976 (N_12976,N_12607,N_12713);
and U12977 (N_12977,N_12613,N_12768);
xnor U12978 (N_12978,N_12714,N_12731);
or U12979 (N_12979,N_12711,N_12755);
nand U12980 (N_12980,N_12639,N_12779);
xor U12981 (N_12981,N_12774,N_12783);
and U12982 (N_12982,N_12769,N_12753);
xor U12983 (N_12983,N_12683,N_12743);
nand U12984 (N_12984,N_12620,N_12717);
nor U12985 (N_12985,N_12610,N_12645);
xnor U12986 (N_12986,N_12784,N_12792);
or U12987 (N_12987,N_12701,N_12786);
nand U12988 (N_12988,N_12618,N_12688);
nand U12989 (N_12989,N_12646,N_12626);
nand U12990 (N_12990,N_12781,N_12682);
xnor U12991 (N_12991,N_12666,N_12690);
nand U12992 (N_12992,N_12692,N_12718);
nand U12993 (N_12993,N_12635,N_12639);
and U12994 (N_12994,N_12691,N_12763);
and U12995 (N_12995,N_12610,N_12739);
nor U12996 (N_12996,N_12721,N_12602);
nor U12997 (N_12997,N_12772,N_12650);
nor U12998 (N_12998,N_12681,N_12783);
nor U12999 (N_12999,N_12655,N_12786);
or U13000 (N_13000,N_12858,N_12817);
xor U13001 (N_13001,N_12975,N_12945);
nor U13002 (N_13002,N_12946,N_12922);
xor U13003 (N_13003,N_12883,N_12928);
nor U13004 (N_13004,N_12894,N_12899);
and U13005 (N_13005,N_12997,N_12958);
xor U13006 (N_13006,N_12976,N_12926);
xor U13007 (N_13007,N_12878,N_12921);
or U13008 (N_13008,N_12836,N_12935);
nor U13009 (N_13009,N_12927,N_12850);
or U13010 (N_13010,N_12810,N_12844);
and U13011 (N_13011,N_12845,N_12822);
xor U13012 (N_13012,N_12914,N_12869);
and U13013 (N_13013,N_12989,N_12964);
nand U13014 (N_13014,N_12977,N_12853);
and U13015 (N_13015,N_12875,N_12936);
xor U13016 (N_13016,N_12880,N_12999);
nand U13017 (N_13017,N_12994,N_12983);
and U13018 (N_13018,N_12985,N_12904);
xnor U13019 (N_13019,N_12961,N_12930);
and U13020 (N_13020,N_12944,N_12916);
xnor U13021 (N_13021,N_12959,N_12966);
xnor U13022 (N_13022,N_12950,N_12988);
nor U13023 (N_13023,N_12803,N_12938);
nand U13024 (N_13024,N_12849,N_12973);
xnor U13025 (N_13025,N_12889,N_12837);
and U13026 (N_13026,N_12847,N_12905);
nand U13027 (N_13027,N_12826,N_12925);
and U13028 (N_13028,N_12862,N_12949);
or U13029 (N_13029,N_12998,N_12865);
nor U13030 (N_13030,N_12821,N_12800);
and U13031 (N_13031,N_12972,N_12952);
nand U13032 (N_13032,N_12948,N_12932);
or U13033 (N_13033,N_12830,N_12912);
nand U13034 (N_13034,N_12808,N_12963);
nand U13035 (N_13035,N_12873,N_12868);
nand U13036 (N_13036,N_12891,N_12834);
nand U13037 (N_13037,N_12979,N_12953);
and U13038 (N_13038,N_12902,N_12968);
xor U13039 (N_13039,N_12892,N_12887);
and U13040 (N_13040,N_12813,N_12969);
and U13041 (N_13041,N_12890,N_12896);
and U13042 (N_13042,N_12851,N_12954);
xor U13043 (N_13043,N_12835,N_12801);
nor U13044 (N_13044,N_12960,N_12860);
and U13045 (N_13045,N_12937,N_12993);
and U13046 (N_13046,N_12978,N_12915);
xor U13047 (N_13047,N_12843,N_12841);
or U13048 (N_13048,N_12934,N_12802);
and U13049 (N_13049,N_12917,N_12913);
xnor U13050 (N_13050,N_12876,N_12906);
nor U13051 (N_13051,N_12811,N_12918);
nor U13052 (N_13052,N_12943,N_12819);
nor U13053 (N_13053,N_12939,N_12842);
nor U13054 (N_13054,N_12984,N_12856);
and U13055 (N_13055,N_12804,N_12852);
nand U13056 (N_13056,N_12931,N_12857);
or U13057 (N_13057,N_12827,N_12941);
and U13058 (N_13058,N_12866,N_12861);
nand U13059 (N_13059,N_12848,N_12859);
and U13060 (N_13060,N_12971,N_12920);
and U13061 (N_13061,N_12816,N_12871);
and U13062 (N_13062,N_12846,N_12987);
and U13063 (N_13063,N_12838,N_12806);
and U13064 (N_13064,N_12893,N_12924);
or U13065 (N_13065,N_12990,N_12992);
nor U13066 (N_13066,N_12907,N_12867);
nor U13067 (N_13067,N_12901,N_12809);
nand U13068 (N_13068,N_12974,N_12855);
nand U13069 (N_13069,N_12910,N_12986);
nand U13070 (N_13070,N_12864,N_12940);
nand U13071 (N_13071,N_12957,N_12995);
nand U13072 (N_13072,N_12947,N_12818);
nor U13073 (N_13073,N_12820,N_12923);
nand U13074 (N_13074,N_12933,N_12909);
nand U13075 (N_13075,N_12956,N_12900);
or U13076 (N_13076,N_12903,N_12828);
nand U13077 (N_13077,N_12829,N_12839);
xnor U13078 (N_13078,N_12870,N_12967);
or U13079 (N_13079,N_12807,N_12886);
and U13080 (N_13080,N_12882,N_12897);
or U13081 (N_13081,N_12812,N_12951);
nand U13082 (N_13082,N_12955,N_12823);
nand U13083 (N_13083,N_12898,N_12962);
nor U13084 (N_13084,N_12877,N_12840);
nand U13085 (N_13085,N_12911,N_12991);
xnor U13086 (N_13086,N_12970,N_12824);
nand U13087 (N_13087,N_12815,N_12874);
or U13088 (N_13088,N_12919,N_12863);
and U13089 (N_13089,N_12996,N_12884);
nor U13090 (N_13090,N_12805,N_12895);
and U13091 (N_13091,N_12814,N_12825);
xnor U13092 (N_13092,N_12980,N_12831);
nor U13093 (N_13093,N_12832,N_12981);
nand U13094 (N_13094,N_12872,N_12854);
or U13095 (N_13095,N_12885,N_12879);
nor U13096 (N_13096,N_12881,N_12888);
nor U13097 (N_13097,N_12908,N_12942);
or U13098 (N_13098,N_12833,N_12982);
or U13099 (N_13099,N_12929,N_12965);
or U13100 (N_13100,N_12933,N_12925);
or U13101 (N_13101,N_12994,N_12975);
or U13102 (N_13102,N_12923,N_12979);
and U13103 (N_13103,N_12848,N_12980);
and U13104 (N_13104,N_12832,N_12978);
nor U13105 (N_13105,N_12926,N_12844);
and U13106 (N_13106,N_12865,N_12925);
or U13107 (N_13107,N_12851,N_12816);
nor U13108 (N_13108,N_12961,N_12918);
xor U13109 (N_13109,N_12939,N_12830);
xor U13110 (N_13110,N_12983,N_12912);
and U13111 (N_13111,N_12885,N_12912);
and U13112 (N_13112,N_12924,N_12937);
nand U13113 (N_13113,N_12976,N_12991);
or U13114 (N_13114,N_12870,N_12802);
xor U13115 (N_13115,N_12861,N_12948);
nor U13116 (N_13116,N_12981,N_12954);
nor U13117 (N_13117,N_12872,N_12857);
xnor U13118 (N_13118,N_12808,N_12974);
xor U13119 (N_13119,N_12870,N_12938);
and U13120 (N_13120,N_12822,N_12962);
nor U13121 (N_13121,N_12938,N_12940);
xnor U13122 (N_13122,N_12841,N_12855);
nor U13123 (N_13123,N_12900,N_12964);
nand U13124 (N_13124,N_12951,N_12811);
xnor U13125 (N_13125,N_12824,N_12935);
and U13126 (N_13126,N_12939,N_12903);
nor U13127 (N_13127,N_12820,N_12856);
and U13128 (N_13128,N_12814,N_12894);
and U13129 (N_13129,N_12878,N_12981);
nand U13130 (N_13130,N_12935,N_12922);
and U13131 (N_13131,N_12800,N_12817);
and U13132 (N_13132,N_12969,N_12823);
xnor U13133 (N_13133,N_12876,N_12868);
xnor U13134 (N_13134,N_12839,N_12891);
or U13135 (N_13135,N_12809,N_12810);
and U13136 (N_13136,N_12824,N_12917);
and U13137 (N_13137,N_12995,N_12937);
or U13138 (N_13138,N_12954,N_12982);
or U13139 (N_13139,N_12973,N_12943);
or U13140 (N_13140,N_12828,N_12953);
or U13141 (N_13141,N_12957,N_12916);
xor U13142 (N_13142,N_12901,N_12966);
and U13143 (N_13143,N_12801,N_12862);
or U13144 (N_13144,N_12837,N_12980);
nor U13145 (N_13145,N_12996,N_12909);
or U13146 (N_13146,N_12873,N_12936);
nor U13147 (N_13147,N_12826,N_12954);
nor U13148 (N_13148,N_12998,N_12896);
and U13149 (N_13149,N_12951,N_12948);
xnor U13150 (N_13150,N_12868,N_12810);
or U13151 (N_13151,N_12834,N_12971);
nor U13152 (N_13152,N_12948,N_12946);
and U13153 (N_13153,N_12877,N_12862);
or U13154 (N_13154,N_12984,N_12881);
and U13155 (N_13155,N_12912,N_12906);
xor U13156 (N_13156,N_12813,N_12856);
nand U13157 (N_13157,N_12909,N_12980);
xnor U13158 (N_13158,N_12847,N_12956);
nand U13159 (N_13159,N_12961,N_12999);
xnor U13160 (N_13160,N_12843,N_12861);
xor U13161 (N_13161,N_12812,N_12843);
and U13162 (N_13162,N_12912,N_12821);
nor U13163 (N_13163,N_12978,N_12827);
nand U13164 (N_13164,N_12958,N_12998);
or U13165 (N_13165,N_12894,N_12821);
and U13166 (N_13166,N_12946,N_12837);
and U13167 (N_13167,N_12919,N_12964);
nor U13168 (N_13168,N_12930,N_12876);
nor U13169 (N_13169,N_12947,N_12829);
and U13170 (N_13170,N_12848,N_12999);
or U13171 (N_13171,N_12992,N_12943);
or U13172 (N_13172,N_12835,N_12906);
or U13173 (N_13173,N_12867,N_12991);
xnor U13174 (N_13174,N_12832,N_12874);
nor U13175 (N_13175,N_12894,N_12956);
nand U13176 (N_13176,N_12846,N_12819);
and U13177 (N_13177,N_12958,N_12981);
and U13178 (N_13178,N_12847,N_12881);
xnor U13179 (N_13179,N_12933,N_12974);
xnor U13180 (N_13180,N_12919,N_12965);
or U13181 (N_13181,N_12880,N_12854);
or U13182 (N_13182,N_12862,N_12962);
and U13183 (N_13183,N_12878,N_12961);
or U13184 (N_13184,N_12982,N_12999);
nor U13185 (N_13185,N_12814,N_12888);
nand U13186 (N_13186,N_12858,N_12939);
and U13187 (N_13187,N_12817,N_12888);
xnor U13188 (N_13188,N_12920,N_12969);
or U13189 (N_13189,N_12827,N_12967);
and U13190 (N_13190,N_12802,N_12823);
or U13191 (N_13191,N_12986,N_12961);
nor U13192 (N_13192,N_12913,N_12948);
and U13193 (N_13193,N_12960,N_12968);
and U13194 (N_13194,N_12974,N_12951);
nand U13195 (N_13195,N_12996,N_12943);
nor U13196 (N_13196,N_12899,N_12946);
and U13197 (N_13197,N_12819,N_12870);
xor U13198 (N_13198,N_12981,N_12955);
nor U13199 (N_13199,N_12999,N_12818);
or U13200 (N_13200,N_13082,N_13012);
and U13201 (N_13201,N_13092,N_13088);
xor U13202 (N_13202,N_13046,N_13022);
and U13203 (N_13203,N_13100,N_13049);
nand U13204 (N_13204,N_13039,N_13098);
and U13205 (N_13205,N_13078,N_13140);
nand U13206 (N_13206,N_13043,N_13027);
xor U13207 (N_13207,N_13014,N_13032);
and U13208 (N_13208,N_13040,N_13182);
and U13209 (N_13209,N_13143,N_13139);
or U13210 (N_13210,N_13174,N_13047);
and U13211 (N_13211,N_13054,N_13002);
xor U13212 (N_13212,N_13094,N_13083);
or U13213 (N_13213,N_13133,N_13165);
and U13214 (N_13214,N_13162,N_13086);
xor U13215 (N_13215,N_13087,N_13136);
and U13216 (N_13216,N_13158,N_13144);
and U13217 (N_13217,N_13189,N_13147);
or U13218 (N_13218,N_13085,N_13106);
or U13219 (N_13219,N_13150,N_13091);
and U13220 (N_13220,N_13180,N_13151);
or U13221 (N_13221,N_13058,N_13007);
nor U13222 (N_13222,N_13041,N_13141);
nor U13223 (N_13223,N_13124,N_13123);
nand U13224 (N_13224,N_13060,N_13109);
xor U13225 (N_13225,N_13062,N_13081);
or U13226 (N_13226,N_13108,N_13161);
xor U13227 (N_13227,N_13072,N_13132);
xnor U13228 (N_13228,N_13026,N_13168);
xnor U13229 (N_13229,N_13005,N_13163);
xnor U13230 (N_13230,N_13175,N_13152);
nand U13231 (N_13231,N_13122,N_13053);
nor U13232 (N_13232,N_13125,N_13001);
nor U13233 (N_13233,N_13111,N_13178);
nor U13234 (N_13234,N_13008,N_13167);
and U13235 (N_13235,N_13157,N_13070);
and U13236 (N_13236,N_13142,N_13033);
and U13237 (N_13237,N_13076,N_13114);
or U13238 (N_13238,N_13126,N_13044);
and U13239 (N_13239,N_13154,N_13093);
xnor U13240 (N_13240,N_13057,N_13119);
nand U13241 (N_13241,N_13159,N_13071);
and U13242 (N_13242,N_13055,N_13128);
or U13243 (N_13243,N_13199,N_13160);
or U13244 (N_13244,N_13010,N_13068);
nand U13245 (N_13245,N_13045,N_13117);
and U13246 (N_13246,N_13052,N_13185);
xor U13247 (N_13247,N_13021,N_13192);
xnor U13248 (N_13248,N_13112,N_13110);
nand U13249 (N_13249,N_13149,N_13066);
nor U13250 (N_13250,N_13176,N_13181);
nand U13251 (N_13251,N_13077,N_13197);
and U13252 (N_13252,N_13025,N_13024);
and U13253 (N_13253,N_13193,N_13000);
or U13254 (N_13254,N_13073,N_13015);
xnor U13255 (N_13255,N_13095,N_13031);
xnor U13256 (N_13256,N_13080,N_13156);
nor U13257 (N_13257,N_13016,N_13198);
or U13258 (N_13258,N_13155,N_13051);
nand U13259 (N_13259,N_13067,N_13153);
nor U13260 (N_13260,N_13146,N_13103);
xor U13261 (N_13261,N_13191,N_13089);
xor U13262 (N_13262,N_13101,N_13020);
nor U13263 (N_13263,N_13096,N_13018);
or U13264 (N_13264,N_13035,N_13172);
xor U13265 (N_13265,N_13166,N_13063);
xor U13266 (N_13266,N_13138,N_13116);
or U13267 (N_13267,N_13013,N_13171);
xor U13268 (N_13268,N_13183,N_13127);
or U13269 (N_13269,N_13048,N_13006);
or U13270 (N_13270,N_13042,N_13059);
and U13271 (N_13271,N_13069,N_13164);
xor U13272 (N_13272,N_13099,N_13009);
and U13273 (N_13273,N_13134,N_13090);
nor U13274 (N_13274,N_13148,N_13034);
nand U13275 (N_13275,N_13118,N_13177);
or U13276 (N_13276,N_13194,N_13170);
or U13277 (N_13277,N_13079,N_13135);
and U13278 (N_13278,N_13003,N_13169);
nand U13279 (N_13279,N_13097,N_13105);
or U13280 (N_13280,N_13104,N_13173);
nor U13281 (N_13281,N_13184,N_13061);
or U13282 (N_13282,N_13029,N_13017);
xor U13283 (N_13283,N_13179,N_13121);
nor U13284 (N_13284,N_13004,N_13011);
or U13285 (N_13285,N_13130,N_13065);
and U13286 (N_13286,N_13028,N_13120);
and U13287 (N_13287,N_13030,N_13131);
or U13288 (N_13288,N_13187,N_13115);
nor U13289 (N_13289,N_13102,N_13137);
or U13290 (N_13290,N_13190,N_13188);
and U13291 (N_13291,N_13129,N_13195);
or U13292 (N_13292,N_13050,N_13075);
nor U13293 (N_13293,N_13113,N_13084);
nand U13294 (N_13294,N_13107,N_13023);
and U13295 (N_13295,N_13038,N_13145);
nand U13296 (N_13296,N_13036,N_13019);
or U13297 (N_13297,N_13196,N_13064);
or U13298 (N_13298,N_13186,N_13037);
xor U13299 (N_13299,N_13074,N_13056);
or U13300 (N_13300,N_13046,N_13103);
xnor U13301 (N_13301,N_13179,N_13186);
nor U13302 (N_13302,N_13198,N_13195);
nand U13303 (N_13303,N_13132,N_13008);
xnor U13304 (N_13304,N_13185,N_13099);
nand U13305 (N_13305,N_13060,N_13043);
nor U13306 (N_13306,N_13061,N_13174);
and U13307 (N_13307,N_13122,N_13047);
and U13308 (N_13308,N_13115,N_13133);
nand U13309 (N_13309,N_13182,N_13077);
xor U13310 (N_13310,N_13140,N_13105);
or U13311 (N_13311,N_13025,N_13193);
and U13312 (N_13312,N_13084,N_13017);
or U13313 (N_13313,N_13168,N_13056);
nand U13314 (N_13314,N_13152,N_13141);
or U13315 (N_13315,N_13155,N_13170);
nand U13316 (N_13316,N_13175,N_13108);
nand U13317 (N_13317,N_13041,N_13068);
nand U13318 (N_13318,N_13075,N_13096);
xor U13319 (N_13319,N_13078,N_13153);
or U13320 (N_13320,N_13146,N_13107);
or U13321 (N_13321,N_13140,N_13150);
nor U13322 (N_13322,N_13082,N_13018);
or U13323 (N_13323,N_13146,N_13028);
nand U13324 (N_13324,N_13047,N_13186);
xnor U13325 (N_13325,N_13038,N_13158);
or U13326 (N_13326,N_13175,N_13050);
or U13327 (N_13327,N_13125,N_13051);
or U13328 (N_13328,N_13151,N_13013);
or U13329 (N_13329,N_13039,N_13073);
or U13330 (N_13330,N_13154,N_13173);
and U13331 (N_13331,N_13045,N_13052);
or U13332 (N_13332,N_13160,N_13193);
and U13333 (N_13333,N_13064,N_13021);
xor U13334 (N_13334,N_13040,N_13154);
nand U13335 (N_13335,N_13015,N_13012);
and U13336 (N_13336,N_13113,N_13066);
nand U13337 (N_13337,N_13199,N_13092);
or U13338 (N_13338,N_13149,N_13107);
and U13339 (N_13339,N_13187,N_13008);
nand U13340 (N_13340,N_13034,N_13100);
and U13341 (N_13341,N_13041,N_13048);
nand U13342 (N_13342,N_13040,N_13103);
or U13343 (N_13343,N_13061,N_13113);
nor U13344 (N_13344,N_13056,N_13085);
or U13345 (N_13345,N_13193,N_13059);
or U13346 (N_13346,N_13109,N_13017);
nor U13347 (N_13347,N_13164,N_13161);
and U13348 (N_13348,N_13153,N_13166);
or U13349 (N_13349,N_13046,N_13013);
nor U13350 (N_13350,N_13028,N_13115);
nand U13351 (N_13351,N_13104,N_13143);
and U13352 (N_13352,N_13073,N_13173);
nand U13353 (N_13353,N_13169,N_13149);
xnor U13354 (N_13354,N_13143,N_13116);
nand U13355 (N_13355,N_13102,N_13180);
xnor U13356 (N_13356,N_13176,N_13032);
and U13357 (N_13357,N_13087,N_13115);
xor U13358 (N_13358,N_13166,N_13009);
xnor U13359 (N_13359,N_13105,N_13106);
nor U13360 (N_13360,N_13198,N_13182);
nor U13361 (N_13361,N_13094,N_13146);
xnor U13362 (N_13362,N_13057,N_13146);
nand U13363 (N_13363,N_13120,N_13067);
nor U13364 (N_13364,N_13187,N_13043);
nand U13365 (N_13365,N_13067,N_13190);
nand U13366 (N_13366,N_13151,N_13171);
xor U13367 (N_13367,N_13093,N_13090);
nor U13368 (N_13368,N_13077,N_13119);
or U13369 (N_13369,N_13176,N_13091);
nand U13370 (N_13370,N_13019,N_13147);
or U13371 (N_13371,N_13154,N_13037);
and U13372 (N_13372,N_13129,N_13056);
nor U13373 (N_13373,N_13178,N_13105);
nand U13374 (N_13374,N_13061,N_13121);
xnor U13375 (N_13375,N_13065,N_13090);
nor U13376 (N_13376,N_13127,N_13033);
nand U13377 (N_13377,N_13026,N_13107);
xnor U13378 (N_13378,N_13036,N_13180);
nor U13379 (N_13379,N_13008,N_13062);
and U13380 (N_13380,N_13033,N_13023);
nor U13381 (N_13381,N_13132,N_13043);
nor U13382 (N_13382,N_13186,N_13005);
or U13383 (N_13383,N_13109,N_13127);
and U13384 (N_13384,N_13093,N_13126);
or U13385 (N_13385,N_13147,N_13103);
xor U13386 (N_13386,N_13198,N_13055);
xnor U13387 (N_13387,N_13177,N_13157);
and U13388 (N_13388,N_13099,N_13171);
nand U13389 (N_13389,N_13147,N_13005);
and U13390 (N_13390,N_13041,N_13088);
xor U13391 (N_13391,N_13193,N_13199);
nand U13392 (N_13392,N_13190,N_13066);
or U13393 (N_13393,N_13099,N_13086);
nor U13394 (N_13394,N_13040,N_13000);
nor U13395 (N_13395,N_13141,N_13186);
nand U13396 (N_13396,N_13017,N_13097);
or U13397 (N_13397,N_13169,N_13157);
xnor U13398 (N_13398,N_13153,N_13049);
nor U13399 (N_13399,N_13118,N_13167);
nand U13400 (N_13400,N_13332,N_13315);
nor U13401 (N_13401,N_13364,N_13220);
xor U13402 (N_13402,N_13235,N_13236);
and U13403 (N_13403,N_13371,N_13383);
and U13404 (N_13404,N_13234,N_13312);
and U13405 (N_13405,N_13393,N_13359);
xnor U13406 (N_13406,N_13372,N_13388);
or U13407 (N_13407,N_13333,N_13376);
nor U13408 (N_13408,N_13317,N_13392);
or U13409 (N_13409,N_13322,N_13213);
xor U13410 (N_13410,N_13203,N_13370);
xor U13411 (N_13411,N_13335,N_13296);
or U13412 (N_13412,N_13204,N_13390);
nand U13413 (N_13413,N_13222,N_13255);
xor U13414 (N_13414,N_13395,N_13381);
and U13415 (N_13415,N_13337,N_13346);
and U13416 (N_13416,N_13215,N_13287);
and U13417 (N_13417,N_13365,N_13258);
nor U13418 (N_13418,N_13386,N_13290);
nor U13419 (N_13419,N_13217,N_13301);
or U13420 (N_13420,N_13253,N_13257);
and U13421 (N_13421,N_13309,N_13303);
or U13422 (N_13422,N_13274,N_13262);
nor U13423 (N_13423,N_13248,N_13329);
nand U13424 (N_13424,N_13208,N_13350);
nand U13425 (N_13425,N_13252,N_13230);
xnor U13426 (N_13426,N_13278,N_13345);
and U13427 (N_13427,N_13357,N_13266);
and U13428 (N_13428,N_13354,N_13341);
or U13429 (N_13429,N_13367,N_13307);
nand U13430 (N_13430,N_13308,N_13318);
xor U13431 (N_13431,N_13219,N_13273);
nand U13432 (N_13432,N_13325,N_13200);
nand U13433 (N_13433,N_13327,N_13311);
and U13434 (N_13434,N_13225,N_13216);
nand U13435 (N_13435,N_13326,N_13348);
nor U13436 (N_13436,N_13299,N_13397);
xnor U13437 (N_13437,N_13275,N_13382);
nand U13438 (N_13438,N_13347,N_13368);
nand U13439 (N_13439,N_13277,N_13384);
nand U13440 (N_13440,N_13242,N_13358);
nor U13441 (N_13441,N_13211,N_13391);
and U13442 (N_13442,N_13214,N_13380);
nor U13443 (N_13443,N_13340,N_13209);
nand U13444 (N_13444,N_13334,N_13279);
and U13445 (N_13445,N_13264,N_13302);
nor U13446 (N_13446,N_13286,N_13344);
xor U13447 (N_13447,N_13339,N_13298);
nor U13448 (N_13448,N_13244,N_13378);
nand U13449 (N_13449,N_13269,N_13336);
xnor U13450 (N_13450,N_13228,N_13305);
xnor U13451 (N_13451,N_13362,N_13316);
nand U13452 (N_13452,N_13319,N_13281);
nand U13453 (N_13453,N_13352,N_13377);
nor U13454 (N_13454,N_13379,N_13321);
xnor U13455 (N_13455,N_13342,N_13324);
xnor U13456 (N_13456,N_13261,N_13226);
and U13457 (N_13457,N_13293,N_13265);
nand U13458 (N_13458,N_13238,N_13250);
and U13459 (N_13459,N_13314,N_13224);
and U13460 (N_13460,N_13267,N_13237);
xnor U13461 (N_13461,N_13223,N_13231);
xor U13462 (N_13462,N_13313,N_13243);
nor U13463 (N_13463,N_13291,N_13276);
nor U13464 (N_13464,N_13297,N_13260);
and U13465 (N_13465,N_13233,N_13241);
or U13466 (N_13466,N_13306,N_13251);
and U13467 (N_13467,N_13328,N_13320);
xor U13468 (N_13468,N_13207,N_13280);
nand U13469 (N_13469,N_13353,N_13263);
and U13470 (N_13470,N_13349,N_13221);
xnor U13471 (N_13471,N_13206,N_13284);
and U13472 (N_13472,N_13373,N_13399);
nand U13473 (N_13473,N_13202,N_13394);
nor U13474 (N_13474,N_13396,N_13375);
nor U13475 (N_13475,N_13360,N_13210);
xor U13476 (N_13476,N_13271,N_13323);
nand U13477 (N_13477,N_13256,N_13361);
nand U13478 (N_13478,N_13245,N_13285);
and U13479 (N_13479,N_13363,N_13338);
xnor U13480 (N_13480,N_13398,N_13310);
nand U13481 (N_13481,N_13389,N_13201);
xor U13482 (N_13482,N_13385,N_13205);
and U13483 (N_13483,N_13289,N_13355);
nor U13484 (N_13484,N_13295,N_13331);
xor U13485 (N_13485,N_13239,N_13218);
nor U13486 (N_13486,N_13304,N_13259);
nand U13487 (N_13487,N_13272,N_13366);
xnor U13488 (N_13488,N_13294,N_13270);
nor U13489 (N_13489,N_13247,N_13229);
and U13490 (N_13490,N_13212,N_13268);
nand U13491 (N_13491,N_13240,N_13246);
and U13492 (N_13492,N_13369,N_13288);
xnor U13493 (N_13493,N_13356,N_13351);
or U13494 (N_13494,N_13343,N_13330);
xor U13495 (N_13495,N_13283,N_13374);
and U13496 (N_13496,N_13387,N_13282);
xnor U13497 (N_13497,N_13292,N_13249);
nor U13498 (N_13498,N_13227,N_13232);
nor U13499 (N_13499,N_13254,N_13300);
or U13500 (N_13500,N_13217,N_13204);
nor U13501 (N_13501,N_13333,N_13380);
and U13502 (N_13502,N_13304,N_13364);
nand U13503 (N_13503,N_13270,N_13275);
and U13504 (N_13504,N_13310,N_13252);
or U13505 (N_13505,N_13200,N_13301);
and U13506 (N_13506,N_13325,N_13260);
and U13507 (N_13507,N_13202,N_13330);
xor U13508 (N_13508,N_13265,N_13326);
and U13509 (N_13509,N_13393,N_13282);
nand U13510 (N_13510,N_13346,N_13208);
nor U13511 (N_13511,N_13339,N_13272);
nor U13512 (N_13512,N_13247,N_13341);
xor U13513 (N_13513,N_13266,N_13294);
and U13514 (N_13514,N_13232,N_13245);
nand U13515 (N_13515,N_13324,N_13360);
nor U13516 (N_13516,N_13313,N_13386);
xnor U13517 (N_13517,N_13307,N_13339);
nor U13518 (N_13518,N_13217,N_13308);
xor U13519 (N_13519,N_13245,N_13390);
or U13520 (N_13520,N_13206,N_13211);
and U13521 (N_13521,N_13228,N_13337);
nor U13522 (N_13522,N_13250,N_13251);
xor U13523 (N_13523,N_13217,N_13348);
nand U13524 (N_13524,N_13234,N_13357);
nand U13525 (N_13525,N_13377,N_13208);
or U13526 (N_13526,N_13292,N_13260);
nor U13527 (N_13527,N_13373,N_13389);
nor U13528 (N_13528,N_13235,N_13234);
nor U13529 (N_13529,N_13251,N_13289);
nand U13530 (N_13530,N_13205,N_13261);
nor U13531 (N_13531,N_13200,N_13307);
or U13532 (N_13532,N_13276,N_13250);
nand U13533 (N_13533,N_13305,N_13291);
nand U13534 (N_13534,N_13264,N_13355);
nand U13535 (N_13535,N_13361,N_13246);
xnor U13536 (N_13536,N_13359,N_13325);
or U13537 (N_13537,N_13357,N_13323);
and U13538 (N_13538,N_13201,N_13377);
nor U13539 (N_13539,N_13259,N_13392);
nand U13540 (N_13540,N_13373,N_13267);
or U13541 (N_13541,N_13299,N_13353);
or U13542 (N_13542,N_13207,N_13247);
xor U13543 (N_13543,N_13355,N_13205);
or U13544 (N_13544,N_13395,N_13346);
nand U13545 (N_13545,N_13231,N_13310);
or U13546 (N_13546,N_13226,N_13266);
nor U13547 (N_13547,N_13208,N_13249);
xor U13548 (N_13548,N_13237,N_13296);
and U13549 (N_13549,N_13225,N_13380);
or U13550 (N_13550,N_13385,N_13360);
or U13551 (N_13551,N_13295,N_13373);
and U13552 (N_13552,N_13367,N_13363);
nand U13553 (N_13553,N_13380,N_13398);
nand U13554 (N_13554,N_13363,N_13397);
or U13555 (N_13555,N_13262,N_13246);
or U13556 (N_13556,N_13243,N_13366);
or U13557 (N_13557,N_13349,N_13375);
and U13558 (N_13558,N_13210,N_13385);
nand U13559 (N_13559,N_13264,N_13255);
xor U13560 (N_13560,N_13322,N_13323);
and U13561 (N_13561,N_13222,N_13295);
nor U13562 (N_13562,N_13354,N_13264);
and U13563 (N_13563,N_13298,N_13384);
nand U13564 (N_13564,N_13208,N_13312);
or U13565 (N_13565,N_13337,N_13283);
or U13566 (N_13566,N_13359,N_13384);
nand U13567 (N_13567,N_13223,N_13304);
and U13568 (N_13568,N_13365,N_13268);
and U13569 (N_13569,N_13349,N_13308);
and U13570 (N_13570,N_13263,N_13213);
xor U13571 (N_13571,N_13369,N_13367);
nor U13572 (N_13572,N_13285,N_13223);
or U13573 (N_13573,N_13203,N_13270);
and U13574 (N_13574,N_13266,N_13278);
and U13575 (N_13575,N_13340,N_13288);
nor U13576 (N_13576,N_13246,N_13204);
xnor U13577 (N_13577,N_13371,N_13277);
or U13578 (N_13578,N_13375,N_13299);
and U13579 (N_13579,N_13254,N_13270);
nand U13580 (N_13580,N_13375,N_13226);
xor U13581 (N_13581,N_13374,N_13363);
or U13582 (N_13582,N_13360,N_13289);
or U13583 (N_13583,N_13304,N_13216);
xor U13584 (N_13584,N_13357,N_13392);
nor U13585 (N_13585,N_13311,N_13348);
nand U13586 (N_13586,N_13361,N_13377);
and U13587 (N_13587,N_13383,N_13259);
xnor U13588 (N_13588,N_13391,N_13223);
xnor U13589 (N_13589,N_13232,N_13278);
xnor U13590 (N_13590,N_13218,N_13315);
nor U13591 (N_13591,N_13211,N_13277);
nand U13592 (N_13592,N_13239,N_13292);
and U13593 (N_13593,N_13384,N_13399);
or U13594 (N_13594,N_13229,N_13329);
and U13595 (N_13595,N_13250,N_13360);
xor U13596 (N_13596,N_13359,N_13316);
nand U13597 (N_13597,N_13240,N_13389);
nor U13598 (N_13598,N_13344,N_13238);
or U13599 (N_13599,N_13390,N_13268);
xnor U13600 (N_13600,N_13487,N_13531);
and U13601 (N_13601,N_13527,N_13516);
xnor U13602 (N_13602,N_13561,N_13569);
nor U13603 (N_13603,N_13427,N_13506);
nand U13604 (N_13604,N_13515,N_13567);
and U13605 (N_13605,N_13475,N_13401);
nor U13606 (N_13606,N_13571,N_13538);
nor U13607 (N_13607,N_13444,N_13485);
nand U13608 (N_13608,N_13453,N_13548);
nand U13609 (N_13609,N_13554,N_13517);
and U13610 (N_13610,N_13421,N_13555);
nor U13611 (N_13611,N_13417,N_13513);
nand U13612 (N_13612,N_13454,N_13526);
and U13613 (N_13613,N_13441,N_13519);
or U13614 (N_13614,N_13501,N_13523);
xnor U13615 (N_13615,N_13481,N_13443);
xnor U13616 (N_13616,N_13423,N_13564);
or U13617 (N_13617,N_13546,N_13403);
or U13618 (N_13618,N_13420,N_13514);
nand U13619 (N_13619,N_13438,N_13414);
nor U13620 (N_13620,N_13510,N_13435);
or U13621 (N_13621,N_13479,N_13574);
and U13622 (N_13622,N_13440,N_13432);
nand U13623 (N_13623,N_13568,N_13431);
and U13624 (N_13624,N_13416,N_13412);
nor U13625 (N_13625,N_13558,N_13502);
or U13626 (N_13626,N_13464,N_13525);
and U13627 (N_13627,N_13424,N_13559);
nor U13628 (N_13628,N_13521,N_13422);
nor U13629 (N_13629,N_13596,N_13494);
or U13630 (N_13630,N_13591,N_13542);
nand U13631 (N_13631,N_13406,N_13544);
xnor U13632 (N_13632,N_13592,N_13447);
nor U13633 (N_13633,N_13490,N_13572);
xor U13634 (N_13634,N_13450,N_13587);
and U13635 (N_13635,N_13595,N_13533);
nor U13636 (N_13636,N_13593,N_13570);
xor U13637 (N_13637,N_13573,N_13552);
nor U13638 (N_13638,N_13582,N_13588);
and U13639 (N_13639,N_13549,N_13419);
or U13640 (N_13640,N_13456,N_13476);
and U13641 (N_13641,N_13442,N_13448);
xnor U13642 (N_13642,N_13520,N_13584);
nor U13643 (N_13643,N_13539,N_13409);
or U13644 (N_13644,N_13597,N_13434);
nand U13645 (N_13645,N_13405,N_13497);
xor U13646 (N_13646,N_13451,N_13557);
nand U13647 (N_13647,N_13474,N_13452);
xnor U13648 (N_13648,N_13590,N_13493);
xnor U13649 (N_13649,N_13471,N_13507);
xor U13650 (N_13650,N_13522,N_13551);
nand U13651 (N_13651,N_13484,N_13589);
or U13652 (N_13652,N_13408,N_13524);
nand U13653 (N_13653,N_13425,N_13577);
and U13654 (N_13654,N_13530,N_13581);
nand U13655 (N_13655,N_13511,N_13428);
and U13656 (N_13656,N_13505,N_13537);
xnor U13657 (N_13657,N_13446,N_13585);
or U13658 (N_13658,N_13458,N_13459);
nand U13659 (N_13659,N_13586,N_13534);
nor U13660 (N_13660,N_13565,N_13540);
xor U13661 (N_13661,N_13594,N_13489);
and U13662 (N_13662,N_13402,N_13439);
or U13663 (N_13663,N_13566,N_13461);
nand U13664 (N_13664,N_13430,N_13410);
and U13665 (N_13665,N_13532,N_13478);
nor U13666 (N_13666,N_13598,N_13580);
nand U13667 (N_13667,N_13469,N_13404);
nand U13668 (N_13668,N_13437,N_13529);
xnor U13669 (N_13669,N_13426,N_13407);
or U13670 (N_13670,N_13415,N_13541);
nor U13671 (N_13671,N_13411,N_13528);
xor U13672 (N_13672,N_13449,N_13460);
or U13673 (N_13673,N_13473,N_13433);
and U13674 (N_13674,N_13576,N_13508);
nand U13675 (N_13675,N_13499,N_13536);
or U13676 (N_13676,N_13496,N_13579);
xor U13677 (N_13677,N_13477,N_13482);
and U13678 (N_13678,N_13483,N_13400);
and U13679 (N_13679,N_13470,N_13547);
nor U13680 (N_13680,N_13463,N_13436);
and U13681 (N_13681,N_13465,N_13575);
nor U13682 (N_13682,N_13455,N_13498);
and U13683 (N_13683,N_13495,N_13488);
nand U13684 (N_13684,N_13445,N_13468);
or U13685 (N_13685,N_13429,N_13550);
nor U13686 (N_13686,N_13500,N_13503);
xnor U13687 (N_13687,N_13553,N_13418);
or U13688 (N_13688,N_13562,N_13512);
or U13689 (N_13689,N_13486,N_13556);
or U13690 (N_13690,N_13560,N_13491);
or U13691 (N_13691,N_13545,N_13492);
nor U13692 (N_13692,N_13535,N_13413);
or U13693 (N_13693,N_13466,N_13583);
or U13694 (N_13694,N_13509,N_13467);
xnor U13695 (N_13695,N_13518,N_13599);
or U13696 (N_13696,N_13504,N_13578);
nor U13697 (N_13697,N_13543,N_13563);
xnor U13698 (N_13698,N_13480,N_13462);
nand U13699 (N_13699,N_13472,N_13457);
or U13700 (N_13700,N_13539,N_13450);
or U13701 (N_13701,N_13464,N_13485);
nor U13702 (N_13702,N_13415,N_13544);
and U13703 (N_13703,N_13469,N_13582);
nand U13704 (N_13704,N_13526,N_13432);
nor U13705 (N_13705,N_13505,N_13442);
and U13706 (N_13706,N_13434,N_13467);
or U13707 (N_13707,N_13538,N_13469);
nor U13708 (N_13708,N_13525,N_13585);
and U13709 (N_13709,N_13542,N_13461);
and U13710 (N_13710,N_13429,N_13530);
or U13711 (N_13711,N_13408,N_13508);
or U13712 (N_13712,N_13582,N_13450);
nand U13713 (N_13713,N_13525,N_13428);
or U13714 (N_13714,N_13563,N_13434);
nand U13715 (N_13715,N_13433,N_13424);
nor U13716 (N_13716,N_13414,N_13547);
or U13717 (N_13717,N_13406,N_13442);
and U13718 (N_13718,N_13536,N_13469);
nand U13719 (N_13719,N_13411,N_13403);
and U13720 (N_13720,N_13473,N_13440);
and U13721 (N_13721,N_13430,N_13492);
nand U13722 (N_13722,N_13466,N_13510);
xnor U13723 (N_13723,N_13525,N_13512);
or U13724 (N_13724,N_13406,N_13553);
or U13725 (N_13725,N_13471,N_13533);
or U13726 (N_13726,N_13501,N_13447);
and U13727 (N_13727,N_13591,N_13587);
xor U13728 (N_13728,N_13565,N_13584);
xnor U13729 (N_13729,N_13490,N_13545);
or U13730 (N_13730,N_13457,N_13551);
xnor U13731 (N_13731,N_13408,N_13405);
nand U13732 (N_13732,N_13477,N_13525);
nand U13733 (N_13733,N_13519,N_13445);
or U13734 (N_13734,N_13596,N_13518);
nand U13735 (N_13735,N_13512,N_13549);
or U13736 (N_13736,N_13557,N_13444);
nor U13737 (N_13737,N_13574,N_13458);
nor U13738 (N_13738,N_13404,N_13423);
xor U13739 (N_13739,N_13525,N_13549);
xnor U13740 (N_13740,N_13451,N_13461);
nand U13741 (N_13741,N_13445,N_13421);
nor U13742 (N_13742,N_13520,N_13588);
or U13743 (N_13743,N_13554,N_13483);
nand U13744 (N_13744,N_13445,N_13464);
or U13745 (N_13745,N_13423,N_13427);
nand U13746 (N_13746,N_13575,N_13562);
or U13747 (N_13747,N_13568,N_13469);
xor U13748 (N_13748,N_13410,N_13582);
xnor U13749 (N_13749,N_13550,N_13496);
or U13750 (N_13750,N_13477,N_13563);
and U13751 (N_13751,N_13470,N_13569);
nor U13752 (N_13752,N_13528,N_13443);
or U13753 (N_13753,N_13442,N_13417);
nor U13754 (N_13754,N_13416,N_13401);
xor U13755 (N_13755,N_13592,N_13544);
nor U13756 (N_13756,N_13535,N_13579);
or U13757 (N_13757,N_13436,N_13543);
nor U13758 (N_13758,N_13465,N_13577);
or U13759 (N_13759,N_13545,N_13578);
or U13760 (N_13760,N_13579,N_13557);
xor U13761 (N_13761,N_13532,N_13546);
xnor U13762 (N_13762,N_13405,N_13599);
nor U13763 (N_13763,N_13540,N_13566);
xnor U13764 (N_13764,N_13539,N_13440);
nand U13765 (N_13765,N_13481,N_13488);
nor U13766 (N_13766,N_13561,N_13571);
or U13767 (N_13767,N_13513,N_13432);
xnor U13768 (N_13768,N_13478,N_13470);
or U13769 (N_13769,N_13578,N_13434);
xor U13770 (N_13770,N_13523,N_13406);
xnor U13771 (N_13771,N_13541,N_13418);
xnor U13772 (N_13772,N_13582,N_13486);
nor U13773 (N_13773,N_13421,N_13477);
nand U13774 (N_13774,N_13445,N_13463);
nand U13775 (N_13775,N_13532,N_13567);
nand U13776 (N_13776,N_13539,N_13545);
or U13777 (N_13777,N_13542,N_13478);
nor U13778 (N_13778,N_13578,N_13425);
nor U13779 (N_13779,N_13591,N_13526);
xnor U13780 (N_13780,N_13407,N_13579);
xnor U13781 (N_13781,N_13400,N_13478);
and U13782 (N_13782,N_13416,N_13485);
nor U13783 (N_13783,N_13455,N_13412);
nor U13784 (N_13784,N_13489,N_13595);
and U13785 (N_13785,N_13435,N_13423);
nand U13786 (N_13786,N_13415,N_13434);
and U13787 (N_13787,N_13441,N_13503);
or U13788 (N_13788,N_13526,N_13530);
nand U13789 (N_13789,N_13432,N_13495);
or U13790 (N_13790,N_13531,N_13562);
and U13791 (N_13791,N_13401,N_13473);
nand U13792 (N_13792,N_13465,N_13469);
nand U13793 (N_13793,N_13487,N_13582);
and U13794 (N_13794,N_13467,N_13413);
xor U13795 (N_13795,N_13580,N_13555);
or U13796 (N_13796,N_13456,N_13525);
xnor U13797 (N_13797,N_13412,N_13507);
nor U13798 (N_13798,N_13585,N_13524);
or U13799 (N_13799,N_13552,N_13582);
and U13800 (N_13800,N_13704,N_13636);
nand U13801 (N_13801,N_13645,N_13786);
xnor U13802 (N_13802,N_13741,N_13753);
or U13803 (N_13803,N_13736,N_13605);
and U13804 (N_13804,N_13795,N_13791);
or U13805 (N_13805,N_13799,N_13690);
and U13806 (N_13806,N_13634,N_13647);
nand U13807 (N_13807,N_13610,N_13757);
or U13808 (N_13808,N_13798,N_13728);
xnor U13809 (N_13809,N_13784,N_13670);
and U13810 (N_13810,N_13630,N_13743);
xor U13811 (N_13811,N_13677,N_13653);
or U13812 (N_13812,N_13660,N_13637);
xnor U13813 (N_13813,N_13714,N_13734);
xnor U13814 (N_13814,N_13718,N_13693);
nand U13815 (N_13815,N_13651,N_13613);
nand U13816 (N_13816,N_13742,N_13774);
or U13817 (N_13817,N_13717,N_13655);
nor U13818 (N_13818,N_13681,N_13684);
nand U13819 (N_13819,N_13661,N_13686);
and U13820 (N_13820,N_13797,N_13754);
nor U13821 (N_13821,N_13688,N_13657);
or U13822 (N_13822,N_13648,N_13694);
and U13823 (N_13823,N_13649,N_13671);
and U13824 (N_13824,N_13739,N_13640);
or U13825 (N_13825,N_13773,N_13621);
and U13826 (N_13826,N_13643,N_13745);
nor U13827 (N_13827,N_13765,N_13711);
nand U13828 (N_13828,N_13683,N_13787);
and U13829 (N_13829,N_13723,N_13685);
xnor U13830 (N_13830,N_13738,N_13658);
and U13831 (N_13831,N_13749,N_13703);
and U13832 (N_13832,N_13772,N_13629);
and U13833 (N_13833,N_13789,N_13747);
or U13834 (N_13834,N_13650,N_13779);
xor U13835 (N_13835,N_13733,N_13654);
nor U13836 (N_13836,N_13730,N_13770);
nor U13837 (N_13837,N_13760,N_13708);
nand U13838 (N_13838,N_13682,N_13764);
and U13839 (N_13839,N_13619,N_13755);
nor U13840 (N_13840,N_13776,N_13751);
or U13841 (N_13841,N_13668,N_13792);
nor U13842 (N_13842,N_13627,N_13624);
or U13843 (N_13843,N_13731,N_13740);
xnor U13844 (N_13844,N_13638,N_13665);
or U13845 (N_13845,N_13626,N_13611);
or U13846 (N_13846,N_13608,N_13620);
or U13847 (N_13847,N_13758,N_13622);
xnor U13848 (N_13848,N_13623,N_13782);
or U13849 (N_13849,N_13644,N_13632);
and U13850 (N_13850,N_13631,N_13680);
nand U13851 (N_13851,N_13705,N_13721);
or U13852 (N_13852,N_13635,N_13667);
nand U13853 (N_13853,N_13628,N_13662);
nor U13854 (N_13854,N_13642,N_13724);
nand U13855 (N_13855,N_13687,N_13706);
or U13856 (N_13856,N_13766,N_13676);
nor U13857 (N_13857,N_13794,N_13603);
nor U13858 (N_13858,N_13727,N_13639);
and U13859 (N_13859,N_13725,N_13673);
or U13860 (N_13860,N_13732,N_13615);
or U13861 (N_13861,N_13696,N_13762);
nand U13862 (N_13862,N_13756,N_13771);
nand U13863 (N_13863,N_13710,N_13674);
and U13864 (N_13864,N_13614,N_13726);
and U13865 (N_13865,N_13604,N_13750);
nor U13866 (N_13866,N_13602,N_13692);
and U13867 (N_13867,N_13780,N_13746);
or U13868 (N_13868,N_13607,N_13652);
and U13869 (N_13869,N_13788,N_13783);
xor U13870 (N_13870,N_13695,N_13735);
xnor U13871 (N_13871,N_13664,N_13700);
or U13872 (N_13872,N_13722,N_13663);
and U13873 (N_13873,N_13713,N_13744);
or U13874 (N_13874,N_13600,N_13737);
xnor U13875 (N_13875,N_13625,N_13707);
or U13876 (N_13876,N_13646,N_13748);
and U13877 (N_13877,N_13669,N_13659);
or U13878 (N_13878,N_13633,N_13761);
nand U13879 (N_13879,N_13790,N_13759);
or U13880 (N_13880,N_13715,N_13719);
xnor U13881 (N_13881,N_13678,N_13679);
xnor U13882 (N_13882,N_13793,N_13689);
and U13883 (N_13883,N_13641,N_13763);
or U13884 (N_13884,N_13778,N_13720);
xnor U13885 (N_13885,N_13781,N_13697);
nand U13886 (N_13886,N_13612,N_13609);
or U13887 (N_13887,N_13617,N_13618);
xnor U13888 (N_13888,N_13666,N_13785);
nor U13889 (N_13889,N_13775,N_13712);
nand U13890 (N_13890,N_13691,N_13698);
xnor U13891 (N_13891,N_13656,N_13675);
nand U13892 (N_13892,N_13616,N_13777);
nand U13893 (N_13893,N_13796,N_13716);
and U13894 (N_13894,N_13701,N_13672);
and U13895 (N_13895,N_13699,N_13729);
or U13896 (N_13896,N_13709,N_13768);
xnor U13897 (N_13897,N_13752,N_13767);
xor U13898 (N_13898,N_13769,N_13601);
and U13899 (N_13899,N_13702,N_13606);
nor U13900 (N_13900,N_13693,N_13768);
nor U13901 (N_13901,N_13659,N_13670);
xor U13902 (N_13902,N_13734,N_13796);
nand U13903 (N_13903,N_13764,N_13751);
or U13904 (N_13904,N_13785,N_13738);
xnor U13905 (N_13905,N_13734,N_13743);
xnor U13906 (N_13906,N_13613,N_13762);
or U13907 (N_13907,N_13694,N_13624);
nand U13908 (N_13908,N_13788,N_13761);
and U13909 (N_13909,N_13780,N_13743);
xnor U13910 (N_13910,N_13700,N_13655);
nand U13911 (N_13911,N_13648,N_13603);
and U13912 (N_13912,N_13631,N_13618);
nor U13913 (N_13913,N_13638,N_13712);
nor U13914 (N_13914,N_13711,N_13613);
nor U13915 (N_13915,N_13771,N_13610);
xor U13916 (N_13916,N_13789,N_13750);
nor U13917 (N_13917,N_13738,N_13678);
or U13918 (N_13918,N_13749,N_13612);
nand U13919 (N_13919,N_13770,N_13604);
nand U13920 (N_13920,N_13615,N_13797);
or U13921 (N_13921,N_13754,N_13700);
and U13922 (N_13922,N_13763,N_13720);
xnor U13923 (N_13923,N_13691,N_13635);
or U13924 (N_13924,N_13799,N_13693);
or U13925 (N_13925,N_13640,N_13799);
nor U13926 (N_13926,N_13779,N_13649);
or U13927 (N_13927,N_13754,N_13618);
nor U13928 (N_13928,N_13678,N_13706);
nand U13929 (N_13929,N_13693,N_13623);
nand U13930 (N_13930,N_13760,N_13750);
xor U13931 (N_13931,N_13792,N_13769);
or U13932 (N_13932,N_13714,N_13630);
xnor U13933 (N_13933,N_13658,N_13781);
or U13934 (N_13934,N_13651,N_13752);
xor U13935 (N_13935,N_13642,N_13661);
nand U13936 (N_13936,N_13612,N_13761);
and U13937 (N_13937,N_13750,N_13625);
nor U13938 (N_13938,N_13726,N_13706);
xnor U13939 (N_13939,N_13633,N_13665);
or U13940 (N_13940,N_13780,N_13733);
nor U13941 (N_13941,N_13704,N_13646);
xnor U13942 (N_13942,N_13784,N_13783);
and U13943 (N_13943,N_13624,N_13796);
nand U13944 (N_13944,N_13685,N_13739);
nor U13945 (N_13945,N_13654,N_13716);
xor U13946 (N_13946,N_13753,N_13691);
or U13947 (N_13947,N_13704,N_13740);
or U13948 (N_13948,N_13798,N_13654);
xor U13949 (N_13949,N_13644,N_13640);
and U13950 (N_13950,N_13675,N_13679);
or U13951 (N_13951,N_13659,N_13620);
nor U13952 (N_13952,N_13640,N_13687);
and U13953 (N_13953,N_13656,N_13707);
nand U13954 (N_13954,N_13760,N_13749);
nor U13955 (N_13955,N_13621,N_13624);
and U13956 (N_13956,N_13769,N_13742);
and U13957 (N_13957,N_13604,N_13638);
and U13958 (N_13958,N_13619,N_13777);
nand U13959 (N_13959,N_13683,N_13704);
nand U13960 (N_13960,N_13608,N_13659);
nand U13961 (N_13961,N_13604,N_13752);
xnor U13962 (N_13962,N_13765,N_13618);
nor U13963 (N_13963,N_13773,N_13613);
xor U13964 (N_13964,N_13605,N_13704);
or U13965 (N_13965,N_13701,N_13796);
xnor U13966 (N_13966,N_13681,N_13755);
nand U13967 (N_13967,N_13766,N_13792);
or U13968 (N_13968,N_13708,N_13794);
xnor U13969 (N_13969,N_13617,N_13626);
xor U13970 (N_13970,N_13747,N_13731);
nor U13971 (N_13971,N_13655,N_13778);
and U13972 (N_13972,N_13621,N_13610);
nand U13973 (N_13973,N_13613,N_13603);
nor U13974 (N_13974,N_13777,N_13605);
xnor U13975 (N_13975,N_13696,N_13606);
or U13976 (N_13976,N_13797,N_13644);
nor U13977 (N_13977,N_13666,N_13756);
nand U13978 (N_13978,N_13613,N_13699);
nor U13979 (N_13979,N_13769,N_13662);
or U13980 (N_13980,N_13778,N_13784);
xor U13981 (N_13981,N_13674,N_13684);
or U13982 (N_13982,N_13795,N_13617);
nand U13983 (N_13983,N_13791,N_13618);
nor U13984 (N_13984,N_13776,N_13712);
nand U13985 (N_13985,N_13693,N_13735);
nand U13986 (N_13986,N_13664,N_13689);
nor U13987 (N_13987,N_13630,N_13776);
or U13988 (N_13988,N_13719,N_13782);
nor U13989 (N_13989,N_13671,N_13683);
xnor U13990 (N_13990,N_13625,N_13770);
xor U13991 (N_13991,N_13759,N_13720);
and U13992 (N_13992,N_13708,N_13649);
nand U13993 (N_13993,N_13732,N_13785);
xnor U13994 (N_13994,N_13765,N_13782);
nand U13995 (N_13995,N_13784,N_13660);
nand U13996 (N_13996,N_13664,N_13642);
nand U13997 (N_13997,N_13685,N_13797);
nand U13998 (N_13998,N_13635,N_13641);
nor U13999 (N_13999,N_13634,N_13767);
nand U14000 (N_14000,N_13837,N_13951);
xnor U14001 (N_14001,N_13806,N_13934);
and U14002 (N_14002,N_13980,N_13963);
and U14003 (N_14003,N_13921,N_13836);
nor U14004 (N_14004,N_13924,N_13970);
nand U14005 (N_14005,N_13901,N_13902);
xor U14006 (N_14006,N_13849,N_13813);
and U14007 (N_14007,N_13810,N_13917);
or U14008 (N_14008,N_13882,N_13974);
and U14009 (N_14009,N_13977,N_13877);
nor U14010 (N_14010,N_13843,N_13949);
nor U14011 (N_14011,N_13904,N_13815);
or U14012 (N_14012,N_13985,N_13926);
or U14013 (N_14013,N_13997,N_13862);
or U14014 (N_14014,N_13932,N_13816);
and U14015 (N_14015,N_13938,N_13935);
nand U14016 (N_14016,N_13950,N_13822);
and U14017 (N_14017,N_13819,N_13895);
xnor U14018 (N_14018,N_13920,N_13918);
and U14019 (N_14019,N_13953,N_13878);
xor U14020 (N_14020,N_13820,N_13957);
nand U14021 (N_14021,N_13846,N_13851);
and U14022 (N_14022,N_13907,N_13885);
or U14023 (N_14023,N_13956,N_13898);
nor U14024 (N_14024,N_13839,N_13800);
nor U14025 (N_14025,N_13834,N_13880);
or U14026 (N_14026,N_13841,N_13835);
xnor U14027 (N_14027,N_13884,N_13998);
or U14028 (N_14028,N_13848,N_13826);
nand U14029 (N_14029,N_13940,N_13939);
and U14030 (N_14030,N_13958,N_13908);
xor U14031 (N_14031,N_13899,N_13869);
xnor U14032 (N_14032,N_13812,N_13892);
nor U14033 (N_14033,N_13807,N_13906);
or U14034 (N_14034,N_13801,N_13952);
or U14035 (N_14035,N_13814,N_13919);
nor U14036 (N_14036,N_13829,N_13942);
nand U14037 (N_14037,N_13808,N_13955);
nand U14038 (N_14038,N_13905,N_13911);
nand U14039 (N_14039,N_13865,N_13831);
and U14040 (N_14040,N_13915,N_13881);
nor U14041 (N_14041,N_13978,N_13825);
or U14042 (N_14042,N_13854,N_13943);
or U14043 (N_14043,N_13821,N_13883);
nand U14044 (N_14044,N_13981,N_13967);
xnor U14045 (N_14045,N_13986,N_13954);
nor U14046 (N_14046,N_13993,N_13922);
nand U14047 (N_14047,N_13873,N_13824);
xnor U14048 (N_14048,N_13987,N_13992);
or U14049 (N_14049,N_13976,N_13972);
xor U14050 (N_14050,N_13874,N_13870);
or U14051 (N_14051,N_13979,N_13912);
or U14052 (N_14052,N_13946,N_13844);
nand U14053 (N_14053,N_13893,N_13828);
nor U14054 (N_14054,N_13913,N_13947);
nand U14055 (N_14055,N_13894,N_13975);
nor U14056 (N_14056,N_13944,N_13853);
nor U14057 (N_14057,N_13988,N_13832);
nor U14058 (N_14058,N_13842,N_13966);
or U14059 (N_14059,N_13890,N_13876);
or U14060 (N_14060,N_13996,N_13823);
xor U14061 (N_14061,N_13818,N_13891);
and U14062 (N_14062,N_13941,N_13809);
and U14063 (N_14063,N_13833,N_13838);
xnor U14064 (N_14064,N_13888,N_13968);
xor U14065 (N_14065,N_13864,N_13872);
nor U14066 (N_14066,N_13948,N_13930);
and U14067 (N_14067,N_13945,N_13886);
and U14068 (N_14068,N_13889,N_13802);
nor U14069 (N_14069,N_13961,N_13965);
or U14070 (N_14070,N_13858,N_13868);
and U14071 (N_14071,N_13859,N_13840);
nor U14072 (N_14072,N_13960,N_13857);
and U14073 (N_14073,N_13830,N_13867);
and U14074 (N_14074,N_13982,N_13805);
nand U14075 (N_14075,N_13845,N_13817);
nand U14076 (N_14076,N_13933,N_13804);
nand U14077 (N_14077,N_13896,N_13937);
or U14078 (N_14078,N_13879,N_13929);
xnor U14079 (N_14079,N_13923,N_13875);
and U14080 (N_14080,N_13969,N_13925);
nand U14081 (N_14081,N_13887,N_13811);
or U14082 (N_14082,N_13855,N_13964);
xnor U14083 (N_14083,N_13936,N_13827);
or U14084 (N_14084,N_13995,N_13989);
nand U14085 (N_14085,N_13962,N_13991);
nand U14086 (N_14086,N_13910,N_13860);
nand U14087 (N_14087,N_13871,N_13863);
xor U14088 (N_14088,N_13999,N_13850);
or U14089 (N_14089,N_13971,N_13909);
nand U14090 (N_14090,N_13803,N_13897);
nand U14091 (N_14091,N_13994,N_13931);
nand U14092 (N_14092,N_13852,N_13903);
or U14093 (N_14093,N_13959,N_13866);
nor U14094 (N_14094,N_13847,N_13861);
nand U14095 (N_14095,N_13856,N_13916);
nand U14096 (N_14096,N_13990,N_13973);
or U14097 (N_14097,N_13983,N_13928);
nand U14098 (N_14098,N_13927,N_13984);
or U14099 (N_14099,N_13914,N_13900);
nor U14100 (N_14100,N_13930,N_13906);
or U14101 (N_14101,N_13999,N_13831);
or U14102 (N_14102,N_13946,N_13999);
nor U14103 (N_14103,N_13976,N_13875);
xnor U14104 (N_14104,N_13944,N_13969);
nand U14105 (N_14105,N_13928,N_13874);
nand U14106 (N_14106,N_13889,N_13949);
or U14107 (N_14107,N_13932,N_13949);
nor U14108 (N_14108,N_13998,N_13991);
nor U14109 (N_14109,N_13919,N_13907);
or U14110 (N_14110,N_13871,N_13987);
and U14111 (N_14111,N_13975,N_13961);
or U14112 (N_14112,N_13847,N_13959);
or U14113 (N_14113,N_13945,N_13856);
and U14114 (N_14114,N_13909,N_13870);
or U14115 (N_14115,N_13966,N_13814);
or U14116 (N_14116,N_13981,N_13839);
and U14117 (N_14117,N_13984,N_13851);
and U14118 (N_14118,N_13993,N_13821);
or U14119 (N_14119,N_13978,N_13946);
nand U14120 (N_14120,N_13920,N_13816);
nor U14121 (N_14121,N_13976,N_13868);
or U14122 (N_14122,N_13936,N_13831);
xor U14123 (N_14123,N_13997,N_13881);
nand U14124 (N_14124,N_13987,N_13812);
xor U14125 (N_14125,N_13904,N_13998);
xnor U14126 (N_14126,N_13916,N_13820);
and U14127 (N_14127,N_13982,N_13846);
and U14128 (N_14128,N_13866,N_13902);
nor U14129 (N_14129,N_13962,N_13915);
xor U14130 (N_14130,N_13920,N_13866);
xnor U14131 (N_14131,N_13836,N_13909);
xnor U14132 (N_14132,N_13828,N_13852);
or U14133 (N_14133,N_13929,N_13873);
nand U14134 (N_14134,N_13947,N_13911);
nand U14135 (N_14135,N_13861,N_13875);
and U14136 (N_14136,N_13910,N_13912);
and U14137 (N_14137,N_13940,N_13842);
nor U14138 (N_14138,N_13921,N_13949);
nand U14139 (N_14139,N_13991,N_13867);
xnor U14140 (N_14140,N_13896,N_13902);
nand U14141 (N_14141,N_13830,N_13804);
nand U14142 (N_14142,N_13896,N_13924);
nor U14143 (N_14143,N_13984,N_13942);
nand U14144 (N_14144,N_13828,N_13807);
nor U14145 (N_14145,N_13898,N_13908);
nor U14146 (N_14146,N_13813,N_13904);
nand U14147 (N_14147,N_13925,N_13824);
xor U14148 (N_14148,N_13988,N_13827);
xor U14149 (N_14149,N_13892,N_13881);
and U14150 (N_14150,N_13935,N_13815);
nor U14151 (N_14151,N_13911,N_13972);
xor U14152 (N_14152,N_13840,N_13945);
or U14153 (N_14153,N_13869,N_13875);
and U14154 (N_14154,N_13979,N_13877);
or U14155 (N_14155,N_13976,N_13924);
nand U14156 (N_14156,N_13842,N_13968);
or U14157 (N_14157,N_13812,N_13800);
or U14158 (N_14158,N_13901,N_13867);
or U14159 (N_14159,N_13954,N_13987);
or U14160 (N_14160,N_13989,N_13817);
xor U14161 (N_14161,N_13872,N_13998);
nor U14162 (N_14162,N_13948,N_13978);
and U14163 (N_14163,N_13957,N_13946);
or U14164 (N_14164,N_13885,N_13875);
and U14165 (N_14165,N_13917,N_13880);
or U14166 (N_14166,N_13941,N_13859);
or U14167 (N_14167,N_13982,N_13876);
or U14168 (N_14168,N_13822,N_13895);
and U14169 (N_14169,N_13990,N_13869);
and U14170 (N_14170,N_13909,N_13904);
xor U14171 (N_14171,N_13961,N_13997);
and U14172 (N_14172,N_13951,N_13807);
xnor U14173 (N_14173,N_13935,N_13801);
nor U14174 (N_14174,N_13868,N_13919);
and U14175 (N_14175,N_13916,N_13904);
xnor U14176 (N_14176,N_13937,N_13804);
xnor U14177 (N_14177,N_13953,N_13847);
and U14178 (N_14178,N_13995,N_13808);
xnor U14179 (N_14179,N_13976,N_13889);
xnor U14180 (N_14180,N_13805,N_13939);
nand U14181 (N_14181,N_13859,N_13911);
xnor U14182 (N_14182,N_13843,N_13862);
nor U14183 (N_14183,N_13917,N_13847);
nor U14184 (N_14184,N_13838,N_13898);
and U14185 (N_14185,N_13843,N_13864);
or U14186 (N_14186,N_13802,N_13812);
nor U14187 (N_14187,N_13952,N_13883);
nand U14188 (N_14188,N_13843,N_13858);
xor U14189 (N_14189,N_13912,N_13930);
or U14190 (N_14190,N_13801,N_13876);
nand U14191 (N_14191,N_13994,N_13867);
nor U14192 (N_14192,N_13803,N_13805);
nor U14193 (N_14193,N_13918,N_13961);
and U14194 (N_14194,N_13881,N_13837);
and U14195 (N_14195,N_13872,N_13818);
nor U14196 (N_14196,N_13875,N_13866);
nor U14197 (N_14197,N_13905,N_13955);
and U14198 (N_14198,N_13878,N_13907);
nor U14199 (N_14199,N_13950,N_13910);
nand U14200 (N_14200,N_14115,N_14120);
or U14201 (N_14201,N_14020,N_14182);
and U14202 (N_14202,N_14063,N_14035);
or U14203 (N_14203,N_14065,N_14179);
and U14204 (N_14204,N_14007,N_14085);
xor U14205 (N_14205,N_14172,N_14178);
or U14206 (N_14206,N_14173,N_14117);
nor U14207 (N_14207,N_14052,N_14054);
or U14208 (N_14208,N_14163,N_14145);
nand U14209 (N_14209,N_14156,N_14158);
or U14210 (N_14210,N_14138,N_14045);
xor U14211 (N_14211,N_14022,N_14012);
or U14212 (N_14212,N_14143,N_14177);
nand U14213 (N_14213,N_14036,N_14071);
or U14214 (N_14214,N_14141,N_14095);
nor U14215 (N_14215,N_14099,N_14188);
and U14216 (N_14216,N_14142,N_14058);
or U14217 (N_14217,N_14038,N_14185);
nor U14218 (N_14218,N_14016,N_14018);
nand U14219 (N_14219,N_14186,N_14028);
or U14220 (N_14220,N_14119,N_14109);
xor U14221 (N_14221,N_14032,N_14043);
and U14222 (N_14222,N_14135,N_14030);
xnor U14223 (N_14223,N_14164,N_14023);
nor U14224 (N_14224,N_14195,N_14187);
xnor U14225 (N_14225,N_14066,N_14107);
and U14226 (N_14226,N_14199,N_14064);
or U14227 (N_14227,N_14147,N_14002);
and U14228 (N_14228,N_14046,N_14091);
xnor U14229 (N_14229,N_14034,N_14125);
and U14230 (N_14230,N_14074,N_14031);
or U14231 (N_14231,N_14061,N_14008);
or U14232 (N_14232,N_14001,N_14094);
nand U14233 (N_14233,N_14004,N_14042);
or U14234 (N_14234,N_14152,N_14197);
xor U14235 (N_14235,N_14121,N_14093);
xnor U14236 (N_14236,N_14155,N_14057);
nand U14237 (N_14237,N_14060,N_14111);
nor U14238 (N_14238,N_14056,N_14169);
and U14239 (N_14239,N_14130,N_14067);
nand U14240 (N_14240,N_14171,N_14037);
nor U14241 (N_14241,N_14070,N_14108);
nand U14242 (N_14242,N_14196,N_14026);
nor U14243 (N_14243,N_14017,N_14005);
or U14244 (N_14244,N_14039,N_14009);
nor U14245 (N_14245,N_14087,N_14025);
and U14246 (N_14246,N_14014,N_14180);
nor U14247 (N_14247,N_14090,N_14149);
or U14248 (N_14248,N_14157,N_14134);
nor U14249 (N_14249,N_14132,N_14010);
and U14250 (N_14250,N_14098,N_14154);
or U14251 (N_14251,N_14159,N_14033);
xor U14252 (N_14252,N_14069,N_14165);
or U14253 (N_14253,N_14080,N_14029);
and U14254 (N_14254,N_14047,N_14194);
nor U14255 (N_14255,N_14055,N_14191);
xor U14256 (N_14256,N_14189,N_14162);
or U14257 (N_14257,N_14106,N_14081);
and U14258 (N_14258,N_14190,N_14123);
nor U14259 (N_14259,N_14062,N_14184);
nand U14260 (N_14260,N_14146,N_14024);
xor U14261 (N_14261,N_14088,N_14140);
xor U14262 (N_14262,N_14079,N_14128);
nor U14263 (N_14263,N_14137,N_14041);
nand U14264 (N_14264,N_14096,N_14084);
nand U14265 (N_14265,N_14078,N_14073);
xor U14266 (N_14266,N_14092,N_14110);
nor U14267 (N_14267,N_14124,N_14006);
and U14268 (N_14268,N_14166,N_14175);
xor U14269 (N_14269,N_14100,N_14027);
nor U14270 (N_14270,N_14089,N_14077);
nand U14271 (N_14271,N_14086,N_14198);
nand U14272 (N_14272,N_14104,N_14139);
nor U14273 (N_14273,N_14072,N_14059);
or U14274 (N_14274,N_14116,N_14044);
and U14275 (N_14275,N_14118,N_14183);
nor U14276 (N_14276,N_14129,N_14168);
and U14277 (N_14277,N_14144,N_14151);
or U14278 (N_14278,N_14176,N_14127);
and U14279 (N_14279,N_14076,N_14068);
nand U14280 (N_14280,N_14170,N_14193);
xor U14281 (N_14281,N_14103,N_14075);
and U14282 (N_14282,N_14015,N_14148);
and U14283 (N_14283,N_14019,N_14000);
nand U14284 (N_14284,N_14097,N_14013);
nor U14285 (N_14285,N_14101,N_14167);
nor U14286 (N_14286,N_14048,N_14192);
nand U14287 (N_14287,N_14150,N_14126);
and U14288 (N_14288,N_14083,N_14181);
nor U14289 (N_14289,N_14131,N_14114);
or U14290 (N_14290,N_14136,N_14011);
or U14291 (N_14291,N_14161,N_14105);
and U14292 (N_14292,N_14174,N_14160);
or U14293 (N_14293,N_14040,N_14112);
xor U14294 (N_14294,N_14113,N_14122);
xnor U14295 (N_14295,N_14053,N_14051);
nor U14296 (N_14296,N_14153,N_14102);
nand U14297 (N_14297,N_14021,N_14133);
or U14298 (N_14298,N_14003,N_14049);
and U14299 (N_14299,N_14050,N_14082);
or U14300 (N_14300,N_14135,N_14131);
or U14301 (N_14301,N_14196,N_14086);
xnor U14302 (N_14302,N_14071,N_14046);
xor U14303 (N_14303,N_14196,N_14066);
and U14304 (N_14304,N_14143,N_14051);
nand U14305 (N_14305,N_14083,N_14032);
nor U14306 (N_14306,N_14066,N_14083);
and U14307 (N_14307,N_14177,N_14008);
nor U14308 (N_14308,N_14015,N_14106);
and U14309 (N_14309,N_14175,N_14019);
and U14310 (N_14310,N_14069,N_14090);
nand U14311 (N_14311,N_14148,N_14162);
and U14312 (N_14312,N_14140,N_14035);
nand U14313 (N_14313,N_14012,N_14037);
nor U14314 (N_14314,N_14014,N_14147);
nor U14315 (N_14315,N_14015,N_14013);
xnor U14316 (N_14316,N_14108,N_14187);
nor U14317 (N_14317,N_14068,N_14015);
and U14318 (N_14318,N_14093,N_14009);
or U14319 (N_14319,N_14192,N_14065);
and U14320 (N_14320,N_14081,N_14166);
and U14321 (N_14321,N_14173,N_14164);
nor U14322 (N_14322,N_14031,N_14166);
nor U14323 (N_14323,N_14153,N_14197);
nor U14324 (N_14324,N_14194,N_14087);
nor U14325 (N_14325,N_14181,N_14062);
xnor U14326 (N_14326,N_14124,N_14175);
and U14327 (N_14327,N_14171,N_14177);
nor U14328 (N_14328,N_14138,N_14025);
and U14329 (N_14329,N_14187,N_14023);
or U14330 (N_14330,N_14137,N_14156);
and U14331 (N_14331,N_14070,N_14094);
or U14332 (N_14332,N_14110,N_14013);
or U14333 (N_14333,N_14164,N_14014);
or U14334 (N_14334,N_14104,N_14061);
and U14335 (N_14335,N_14010,N_14130);
or U14336 (N_14336,N_14036,N_14024);
xnor U14337 (N_14337,N_14144,N_14043);
nor U14338 (N_14338,N_14077,N_14147);
nand U14339 (N_14339,N_14151,N_14076);
nor U14340 (N_14340,N_14178,N_14134);
nand U14341 (N_14341,N_14145,N_14147);
or U14342 (N_14342,N_14098,N_14094);
or U14343 (N_14343,N_14083,N_14116);
or U14344 (N_14344,N_14048,N_14026);
nand U14345 (N_14345,N_14143,N_14009);
xnor U14346 (N_14346,N_14069,N_14076);
xnor U14347 (N_14347,N_14024,N_14065);
nand U14348 (N_14348,N_14191,N_14140);
nand U14349 (N_14349,N_14098,N_14187);
nand U14350 (N_14350,N_14128,N_14060);
and U14351 (N_14351,N_14139,N_14029);
nor U14352 (N_14352,N_14088,N_14165);
xnor U14353 (N_14353,N_14140,N_14002);
or U14354 (N_14354,N_14149,N_14051);
and U14355 (N_14355,N_14045,N_14181);
nand U14356 (N_14356,N_14053,N_14115);
or U14357 (N_14357,N_14112,N_14020);
or U14358 (N_14358,N_14022,N_14017);
or U14359 (N_14359,N_14035,N_14176);
nor U14360 (N_14360,N_14018,N_14177);
nor U14361 (N_14361,N_14190,N_14167);
nor U14362 (N_14362,N_14133,N_14086);
xnor U14363 (N_14363,N_14190,N_14145);
xnor U14364 (N_14364,N_14160,N_14079);
xor U14365 (N_14365,N_14098,N_14151);
and U14366 (N_14366,N_14085,N_14123);
and U14367 (N_14367,N_14081,N_14149);
nand U14368 (N_14368,N_14151,N_14049);
nor U14369 (N_14369,N_14044,N_14014);
nand U14370 (N_14370,N_14089,N_14099);
nor U14371 (N_14371,N_14150,N_14028);
or U14372 (N_14372,N_14015,N_14178);
or U14373 (N_14373,N_14079,N_14163);
and U14374 (N_14374,N_14193,N_14126);
xnor U14375 (N_14375,N_14034,N_14186);
xor U14376 (N_14376,N_14193,N_14014);
nand U14377 (N_14377,N_14059,N_14150);
and U14378 (N_14378,N_14190,N_14187);
nor U14379 (N_14379,N_14135,N_14035);
or U14380 (N_14380,N_14095,N_14018);
or U14381 (N_14381,N_14170,N_14053);
or U14382 (N_14382,N_14015,N_14054);
xor U14383 (N_14383,N_14173,N_14044);
nand U14384 (N_14384,N_14085,N_14187);
or U14385 (N_14385,N_14158,N_14166);
and U14386 (N_14386,N_14091,N_14192);
or U14387 (N_14387,N_14146,N_14129);
xor U14388 (N_14388,N_14166,N_14013);
and U14389 (N_14389,N_14105,N_14167);
and U14390 (N_14390,N_14071,N_14123);
and U14391 (N_14391,N_14038,N_14187);
nand U14392 (N_14392,N_14027,N_14042);
or U14393 (N_14393,N_14121,N_14084);
nor U14394 (N_14394,N_14044,N_14119);
or U14395 (N_14395,N_14176,N_14168);
nand U14396 (N_14396,N_14063,N_14090);
nor U14397 (N_14397,N_14189,N_14176);
nand U14398 (N_14398,N_14010,N_14039);
nand U14399 (N_14399,N_14180,N_14054);
nor U14400 (N_14400,N_14259,N_14256);
nor U14401 (N_14401,N_14348,N_14293);
and U14402 (N_14402,N_14308,N_14324);
xnor U14403 (N_14403,N_14353,N_14226);
nor U14404 (N_14404,N_14306,N_14232);
and U14405 (N_14405,N_14282,N_14396);
and U14406 (N_14406,N_14208,N_14260);
or U14407 (N_14407,N_14262,N_14319);
xnor U14408 (N_14408,N_14350,N_14215);
and U14409 (N_14409,N_14337,N_14335);
and U14410 (N_14410,N_14246,N_14371);
xor U14411 (N_14411,N_14300,N_14395);
nor U14412 (N_14412,N_14349,N_14206);
and U14413 (N_14413,N_14228,N_14331);
and U14414 (N_14414,N_14332,N_14330);
and U14415 (N_14415,N_14227,N_14255);
and U14416 (N_14416,N_14356,N_14375);
or U14417 (N_14417,N_14369,N_14296);
or U14418 (N_14418,N_14316,N_14207);
xnor U14419 (N_14419,N_14365,N_14373);
nor U14420 (N_14420,N_14368,N_14270);
nor U14421 (N_14421,N_14276,N_14318);
xnor U14422 (N_14422,N_14242,N_14364);
xor U14423 (N_14423,N_14314,N_14328);
nand U14424 (N_14424,N_14297,N_14252);
and U14425 (N_14425,N_14367,N_14250);
nand U14426 (N_14426,N_14268,N_14392);
nand U14427 (N_14427,N_14239,N_14313);
or U14428 (N_14428,N_14379,N_14346);
xor U14429 (N_14429,N_14281,N_14340);
or U14430 (N_14430,N_14211,N_14283);
or U14431 (N_14431,N_14360,N_14213);
and U14432 (N_14432,N_14298,N_14305);
nand U14433 (N_14433,N_14385,N_14274);
xnor U14434 (N_14434,N_14266,N_14249);
nor U14435 (N_14435,N_14352,N_14389);
nor U14436 (N_14436,N_14220,N_14245);
and U14437 (N_14437,N_14258,N_14240);
nand U14438 (N_14438,N_14272,N_14218);
and U14439 (N_14439,N_14280,N_14388);
and U14440 (N_14440,N_14288,N_14247);
or U14441 (N_14441,N_14370,N_14391);
nor U14442 (N_14442,N_14351,N_14311);
xor U14443 (N_14443,N_14287,N_14285);
and U14444 (N_14444,N_14394,N_14234);
nor U14445 (N_14445,N_14238,N_14248);
and U14446 (N_14446,N_14304,N_14290);
nand U14447 (N_14447,N_14291,N_14320);
xor U14448 (N_14448,N_14386,N_14229);
nand U14449 (N_14449,N_14254,N_14347);
nor U14450 (N_14450,N_14279,N_14237);
nand U14451 (N_14451,N_14358,N_14345);
xor U14452 (N_14452,N_14382,N_14393);
nor U14453 (N_14453,N_14225,N_14200);
or U14454 (N_14454,N_14217,N_14363);
and U14455 (N_14455,N_14244,N_14372);
and U14456 (N_14456,N_14204,N_14212);
xnor U14457 (N_14457,N_14263,N_14310);
and U14458 (N_14458,N_14322,N_14278);
or U14459 (N_14459,N_14292,N_14344);
or U14460 (N_14460,N_14341,N_14334);
nand U14461 (N_14461,N_14203,N_14321);
nor U14462 (N_14462,N_14275,N_14277);
nand U14463 (N_14463,N_14380,N_14210);
and U14464 (N_14464,N_14222,N_14271);
and U14465 (N_14465,N_14294,N_14289);
nor U14466 (N_14466,N_14354,N_14333);
nor U14467 (N_14467,N_14205,N_14267);
nor U14468 (N_14468,N_14261,N_14303);
and U14469 (N_14469,N_14235,N_14301);
or U14470 (N_14470,N_14343,N_14253);
xor U14471 (N_14471,N_14342,N_14378);
nor U14472 (N_14472,N_14284,N_14387);
nand U14473 (N_14473,N_14264,N_14397);
or U14474 (N_14474,N_14336,N_14221);
and U14475 (N_14475,N_14377,N_14241);
or U14476 (N_14476,N_14257,N_14355);
xnor U14477 (N_14477,N_14329,N_14214);
nor U14478 (N_14478,N_14357,N_14265);
nand U14479 (N_14479,N_14376,N_14326);
nand U14480 (N_14480,N_14243,N_14231);
nor U14481 (N_14481,N_14317,N_14323);
nor U14482 (N_14482,N_14299,N_14269);
nand U14483 (N_14483,N_14315,N_14312);
and U14484 (N_14484,N_14202,N_14216);
nor U14485 (N_14485,N_14230,N_14295);
xnor U14486 (N_14486,N_14390,N_14381);
xnor U14487 (N_14487,N_14201,N_14374);
nor U14488 (N_14488,N_14273,N_14233);
or U14489 (N_14489,N_14219,N_14302);
nand U14490 (N_14490,N_14398,N_14362);
nand U14491 (N_14491,N_14236,N_14286);
or U14492 (N_14492,N_14359,N_14383);
and U14493 (N_14493,N_14366,N_14327);
nand U14494 (N_14494,N_14307,N_14209);
and U14495 (N_14495,N_14309,N_14251);
xor U14496 (N_14496,N_14339,N_14399);
xnor U14497 (N_14497,N_14361,N_14224);
nand U14498 (N_14498,N_14338,N_14384);
xor U14499 (N_14499,N_14223,N_14325);
xor U14500 (N_14500,N_14253,N_14366);
xnor U14501 (N_14501,N_14265,N_14384);
xor U14502 (N_14502,N_14371,N_14277);
xor U14503 (N_14503,N_14251,N_14345);
nor U14504 (N_14504,N_14253,N_14237);
nor U14505 (N_14505,N_14347,N_14257);
nand U14506 (N_14506,N_14302,N_14228);
nand U14507 (N_14507,N_14256,N_14205);
nand U14508 (N_14508,N_14243,N_14294);
xnor U14509 (N_14509,N_14261,N_14290);
or U14510 (N_14510,N_14201,N_14344);
nand U14511 (N_14511,N_14368,N_14263);
xor U14512 (N_14512,N_14232,N_14385);
and U14513 (N_14513,N_14312,N_14331);
xnor U14514 (N_14514,N_14211,N_14366);
or U14515 (N_14515,N_14327,N_14289);
xor U14516 (N_14516,N_14314,N_14249);
and U14517 (N_14517,N_14398,N_14393);
and U14518 (N_14518,N_14264,N_14361);
and U14519 (N_14519,N_14223,N_14350);
and U14520 (N_14520,N_14201,N_14313);
xor U14521 (N_14521,N_14313,N_14223);
xor U14522 (N_14522,N_14389,N_14398);
nand U14523 (N_14523,N_14372,N_14280);
nand U14524 (N_14524,N_14208,N_14318);
and U14525 (N_14525,N_14397,N_14378);
xnor U14526 (N_14526,N_14279,N_14338);
nand U14527 (N_14527,N_14307,N_14261);
nor U14528 (N_14528,N_14253,N_14275);
nor U14529 (N_14529,N_14206,N_14364);
nand U14530 (N_14530,N_14376,N_14283);
nor U14531 (N_14531,N_14243,N_14380);
and U14532 (N_14532,N_14226,N_14340);
xnor U14533 (N_14533,N_14309,N_14337);
or U14534 (N_14534,N_14329,N_14286);
nor U14535 (N_14535,N_14357,N_14247);
xnor U14536 (N_14536,N_14247,N_14259);
xor U14537 (N_14537,N_14364,N_14391);
and U14538 (N_14538,N_14324,N_14265);
or U14539 (N_14539,N_14360,N_14329);
nor U14540 (N_14540,N_14235,N_14333);
nor U14541 (N_14541,N_14270,N_14256);
or U14542 (N_14542,N_14384,N_14300);
xor U14543 (N_14543,N_14242,N_14284);
and U14544 (N_14544,N_14254,N_14291);
nand U14545 (N_14545,N_14235,N_14319);
nor U14546 (N_14546,N_14382,N_14333);
nor U14547 (N_14547,N_14351,N_14338);
nand U14548 (N_14548,N_14245,N_14247);
nand U14549 (N_14549,N_14309,N_14296);
and U14550 (N_14550,N_14348,N_14377);
nand U14551 (N_14551,N_14347,N_14276);
xnor U14552 (N_14552,N_14349,N_14224);
nor U14553 (N_14553,N_14233,N_14307);
nand U14554 (N_14554,N_14266,N_14385);
or U14555 (N_14555,N_14286,N_14332);
nor U14556 (N_14556,N_14280,N_14246);
or U14557 (N_14557,N_14219,N_14220);
xor U14558 (N_14558,N_14391,N_14332);
or U14559 (N_14559,N_14290,N_14289);
and U14560 (N_14560,N_14318,N_14322);
or U14561 (N_14561,N_14214,N_14235);
nor U14562 (N_14562,N_14312,N_14261);
or U14563 (N_14563,N_14331,N_14383);
nor U14564 (N_14564,N_14289,N_14271);
nor U14565 (N_14565,N_14261,N_14317);
or U14566 (N_14566,N_14235,N_14203);
and U14567 (N_14567,N_14200,N_14262);
xor U14568 (N_14568,N_14291,N_14302);
or U14569 (N_14569,N_14294,N_14396);
and U14570 (N_14570,N_14267,N_14338);
or U14571 (N_14571,N_14376,N_14293);
nor U14572 (N_14572,N_14384,N_14225);
or U14573 (N_14573,N_14220,N_14224);
xnor U14574 (N_14574,N_14369,N_14241);
and U14575 (N_14575,N_14215,N_14377);
or U14576 (N_14576,N_14271,N_14299);
nor U14577 (N_14577,N_14278,N_14367);
and U14578 (N_14578,N_14202,N_14337);
or U14579 (N_14579,N_14261,N_14348);
nand U14580 (N_14580,N_14312,N_14271);
xnor U14581 (N_14581,N_14211,N_14348);
or U14582 (N_14582,N_14287,N_14314);
xor U14583 (N_14583,N_14313,N_14352);
xnor U14584 (N_14584,N_14386,N_14278);
and U14585 (N_14585,N_14303,N_14206);
nor U14586 (N_14586,N_14347,N_14248);
xor U14587 (N_14587,N_14261,N_14286);
nor U14588 (N_14588,N_14239,N_14237);
and U14589 (N_14589,N_14209,N_14217);
nand U14590 (N_14590,N_14383,N_14340);
nand U14591 (N_14591,N_14348,N_14329);
nor U14592 (N_14592,N_14280,N_14220);
xor U14593 (N_14593,N_14329,N_14278);
nor U14594 (N_14594,N_14310,N_14213);
or U14595 (N_14595,N_14207,N_14328);
and U14596 (N_14596,N_14379,N_14374);
nand U14597 (N_14597,N_14369,N_14335);
and U14598 (N_14598,N_14232,N_14358);
xor U14599 (N_14599,N_14307,N_14295);
or U14600 (N_14600,N_14449,N_14430);
xnor U14601 (N_14601,N_14413,N_14522);
nand U14602 (N_14602,N_14503,N_14498);
nand U14603 (N_14603,N_14462,N_14506);
or U14604 (N_14604,N_14567,N_14452);
and U14605 (N_14605,N_14598,N_14450);
nor U14606 (N_14606,N_14484,N_14436);
xor U14607 (N_14607,N_14599,N_14423);
nand U14608 (N_14608,N_14521,N_14416);
nand U14609 (N_14609,N_14569,N_14494);
nor U14610 (N_14610,N_14568,N_14509);
nor U14611 (N_14611,N_14590,N_14488);
or U14612 (N_14612,N_14508,N_14407);
xor U14613 (N_14613,N_14524,N_14473);
nor U14614 (N_14614,N_14467,N_14469);
and U14615 (N_14615,N_14571,N_14575);
nand U14616 (N_14616,N_14442,N_14441);
or U14617 (N_14617,N_14502,N_14400);
and U14618 (N_14618,N_14585,N_14439);
nand U14619 (N_14619,N_14427,N_14435);
nor U14620 (N_14620,N_14410,N_14543);
nor U14621 (N_14621,N_14472,N_14523);
nand U14622 (N_14622,N_14547,N_14554);
nand U14623 (N_14623,N_14566,N_14564);
and U14624 (N_14624,N_14493,N_14582);
and U14625 (N_14625,N_14565,N_14415);
nor U14626 (N_14626,N_14406,N_14504);
nor U14627 (N_14627,N_14481,N_14588);
nor U14628 (N_14628,N_14425,N_14553);
nand U14629 (N_14629,N_14477,N_14544);
nor U14630 (N_14630,N_14409,N_14587);
nand U14631 (N_14631,N_14478,N_14591);
and U14632 (N_14632,N_14510,N_14448);
or U14633 (N_14633,N_14434,N_14500);
or U14634 (N_14634,N_14556,N_14418);
nor U14635 (N_14635,N_14527,N_14476);
xnor U14636 (N_14636,N_14507,N_14417);
nor U14637 (N_14637,N_14492,N_14520);
and U14638 (N_14638,N_14482,N_14551);
and U14639 (N_14639,N_14437,N_14573);
or U14640 (N_14640,N_14496,N_14411);
or U14641 (N_14641,N_14495,N_14446);
and U14642 (N_14642,N_14589,N_14515);
nor U14643 (N_14643,N_14401,N_14475);
nor U14644 (N_14644,N_14540,N_14432);
nand U14645 (N_14645,N_14546,N_14428);
and U14646 (N_14646,N_14404,N_14445);
nand U14647 (N_14647,N_14451,N_14537);
xnor U14648 (N_14648,N_14586,N_14408);
nand U14649 (N_14649,N_14528,N_14463);
or U14650 (N_14650,N_14516,N_14595);
nor U14651 (N_14651,N_14513,N_14426);
and U14652 (N_14652,N_14489,N_14529);
nand U14653 (N_14653,N_14572,N_14438);
xor U14654 (N_14654,N_14487,N_14542);
and U14655 (N_14655,N_14584,N_14576);
or U14656 (N_14656,N_14447,N_14519);
xor U14657 (N_14657,N_14597,N_14535);
nor U14658 (N_14658,N_14517,N_14431);
or U14659 (N_14659,N_14443,N_14471);
nor U14660 (N_14660,N_14596,N_14460);
and U14661 (N_14661,N_14548,N_14593);
or U14662 (N_14662,N_14552,N_14497);
nand U14663 (N_14663,N_14525,N_14512);
nand U14664 (N_14664,N_14420,N_14479);
xor U14665 (N_14665,N_14444,N_14560);
and U14666 (N_14666,N_14454,N_14433);
nand U14667 (N_14667,N_14501,N_14539);
xnor U14668 (N_14668,N_14559,N_14581);
nand U14669 (N_14669,N_14457,N_14563);
or U14670 (N_14670,N_14424,N_14555);
nor U14671 (N_14671,N_14538,N_14458);
or U14672 (N_14672,N_14403,N_14464);
xnor U14673 (N_14673,N_14534,N_14465);
or U14674 (N_14674,N_14402,N_14419);
or U14675 (N_14675,N_14412,N_14574);
nor U14676 (N_14676,N_14440,N_14526);
xnor U14677 (N_14677,N_14414,N_14461);
xor U14678 (N_14678,N_14533,N_14491);
and U14679 (N_14679,N_14470,N_14511);
or U14680 (N_14680,N_14485,N_14579);
or U14681 (N_14681,N_14421,N_14531);
xnor U14682 (N_14682,N_14558,N_14592);
nor U14683 (N_14683,N_14453,N_14468);
xor U14684 (N_14684,N_14594,N_14459);
nand U14685 (N_14685,N_14505,N_14490);
xnor U14686 (N_14686,N_14561,N_14429);
xnor U14687 (N_14687,N_14536,N_14480);
xnor U14688 (N_14688,N_14466,N_14483);
and U14689 (N_14689,N_14583,N_14549);
and U14690 (N_14690,N_14456,N_14518);
xor U14691 (N_14691,N_14550,N_14541);
and U14692 (N_14692,N_14486,N_14570);
xor U14693 (N_14693,N_14455,N_14532);
or U14694 (N_14694,N_14580,N_14577);
and U14695 (N_14695,N_14562,N_14578);
nor U14696 (N_14696,N_14545,N_14474);
and U14697 (N_14697,N_14499,N_14530);
and U14698 (N_14698,N_14557,N_14405);
or U14699 (N_14699,N_14514,N_14422);
and U14700 (N_14700,N_14584,N_14522);
nand U14701 (N_14701,N_14420,N_14414);
and U14702 (N_14702,N_14412,N_14592);
and U14703 (N_14703,N_14474,N_14565);
and U14704 (N_14704,N_14467,N_14434);
and U14705 (N_14705,N_14539,N_14529);
and U14706 (N_14706,N_14529,N_14422);
or U14707 (N_14707,N_14597,N_14496);
nor U14708 (N_14708,N_14438,N_14536);
and U14709 (N_14709,N_14580,N_14565);
or U14710 (N_14710,N_14579,N_14430);
nand U14711 (N_14711,N_14447,N_14599);
nand U14712 (N_14712,N_14513,N_14430);
nand U14713 (N_14713,N_14598,N_14527);
xor U14714 (N_14714,N_14430,N_14578);
and U14715 (N_14715,N_14594,N_14570);
xor U14716 (N_14716,N_14511,N_14519);
nor U14717 (N_14717,N_14534,N_14567);
nor U14718 (N_14718,N_14580,N_14526);
xnor U14719 (N_14719,N_14417,N_14527);
and U14720 (N_14720,N_14454,N_14545);
nor U14721 (N_14721,N_14585,N_14551);
or U14722 (N_14722,N_14537,N_14530);
xnor U14723 (N_14723,N_14416,N_14564);
or U14724 (N_14724,N_14522,N_14561);
nor U14725 (N_14725,N_14491,N_14492);
nand U14726 (N_14726,N_14527,N_14546);
nand U14727 (N_14727,N_14489,N_14507);
or U14728 (N_14728,N_14584,N_14429);
nand U14729 (N_14729,N_14568,N_14439);
or U14730 (N_14730,N_14584,N_14443);
nand U14731 (N_14731,N_14453,N_14554);
xor U14732 (N_14732,N_14514,N_14565);
nor U14733 (N_14733,N_14506,N_14539);
nand U14734 (N_14734,N_14545,N_14591);
or U14735 (N_14735,N_14468,N_14555);
and U14736 (N_14736,N_14464,N_14526);
or U14737 (N_14737,N_14423,N_14442);
and U14738 (N_14738,N_14425,N_14458);
nand U14739 (N_14739,N_14480,N_14405);
xor U14740 (N_14740,N_14414,N_14432);
xor U14741 (N_14741,N_14465,N_14500);
xnor U14742 (N_14742,N_14466,N_14593);
nand U14743 (N_14743,N_14589,N_14491);
nand U14744 (N_14744,N_14459,N_14404);
nand U14745 (N_14745,N_14562,N_14445);
nor U14746 (N_14746,N_14478,N_14451);
nand U14747 (N_14747,N_14479,N_14542);
nor U14748 (N_14748,N_14477,N_14431);
or U14749 (N_14749,N_14497,N_14414);
xor U14750 (N_14750,N_14560,N_14401);
nand U14751 (N_14751,N_14550,N_14448);
xnor U14752 (N_14752,N_14489,N_14569);
and U14753 (N_14753,N_14572,N_14429);
and U14754 (N_14754,N_14570,N_14527);
xnor U14755 (N_14755,N_14598,N_14405);
xnor U14756 (N_14756,N_14481,N_14421);
xnor U14757 (N_14757,N_14452,N_14557);
or U14758 (N_14758,N_14493,N_14405);
nor U14759 (N_14759,N_14451,N_14572);
and U14760 (N_14760,N_14447,N_14453);
and U14761 (N_14761,N_14528,N_14456);
and U14762 (N_14762,N_14540,N_14440);
or U14763 (N_14763,N_14558,N_14463);
xnor U14764 (N_14764,N_14537,N_14455);
xnor U14765 (N_14765,N_14401,N_14465);
nand U14766 (N_14766,N_14421,N_14472);
and U14767 (N_14767,N_14406,N_14525);
nor U14768 (N_14768,N_14452,N_14518);
xor U14769 (N_14769,N_14595,N_14475);
nand U14770 (N_14770,N_14506,N_14573);
and U14771 (N_14771,N_14553,N_14494);
nand U14772 (N_14772,N_14483,N_14558);
nand U14773 (N_14773,N_14489,N_14405);
and U14774 (N_14774,N_14590,N_14416);
and U14775 (N_14775,N_14474,N_14493);
xor U14776 (N_14776,N_14591,N_14554);
and U14777 (N_14777,N_14599,N_14463);
and U14778 (N_14778,N_14462,N_14459);
and U14779 (N_14779,N_14552,N_14529);
nand U14780 (N_14780,N_14427,N_14519);
or U14781 (N_14781,N_14408,N_14494);
or U14782 (N_14782,N_14422,N_14464);
or U14783 (N_14783,N_14422,N_14596);
xor U14784 (N_14784,N_14521,N_14596);
xor U14785 (N_14785,N_14468,N_14413);
nand U14786 (N_14786,N_14569,N_14467);
or U14787 (N_14787,N_14495,N_14589);
or U14788 (N_14788,N_14540,N_14449);
nor U14789 (N_14789,N_14492,N_14539);
xor U14790 (N_14790,N_14413,N_14488);
xnor U14791 (N_14791,N_14505,N_14542);
nor U14792 (N_14792,N_14404,N_14572);
nor U14793 (N_14793,N_14453,N_14591);
nand U14794 (N_14794,N_14438,N_14479);
xnor U14795 (N_14795,N_14477,N_14517);
and U14796 (N_14796,N_14579,N_14507);
and U14797 (N_14797,N_14561,N_14457);
nor U14798 (N_14798,N_14448,N_14529);
and U14799 (N_14799,N_14574,N_14577);
or U14800 (N_14800,N_14787,N_14658);
and U14801 (N_14801,N_14792,N_14737);
and U14802 (N_14802,N_14609,N_14719);
nor U14803 (N_14803,N_14698,N_14717);
nor U14804 (N_14804,N_14705,N_14613);
nand U14805 (N_14805,N_14751,N_14758);
or U14806 (N_14806,N_14602,N_14670);
or U14807 (N_14807,N_14778,N_14741);
or U14808 (N_14808,N_14684,N_14614);
xor U14809 (N_14809,N_14687,N_14776);
and U14810 (N_14810,N_14706,N_14708);
and U14811 (N_14811,N_14672,N_14699);
nand U14812 (N_14812,N_14761,N_14789);
or U14813 (N_14813,N_14691,N_14653);
nor U14814 (N_14814,N_14606,N_14624);
nor U14815 (N_14815,N_14638,N_14747);
or U14816 (N_14816,N_14635,N_14623);
nor U14817 (N_14817,N_14647,N_14770);
and U14818 (N_14818,N_14600,N_14680);
nor U14819 (N_14819,N_14607,N_14714);
nor U14820 (N_14820,N_14753,N_14671);
nand U14821 (N_14821,N_14669,N_14625);
xor U14822 (N_14822,N_14663,N_14668);
xor U14823 (N_14823,N_14694,N_14674);
nor U14824 (N_14824,N_14750,N_14659);
or U14825 (N_14825,N_14666,N_14718);
nand U14826 (N_14826,N_14745,N_14756);
nand U14827 (N_14827,N_14733,N_14768);
xor U14828 (N_14828,N_14785,N_14738);
or U14829 (N_14829,N_14755,N_14657);
nor U14830 (N_14830,N_14730,N_14743);
xor U14831 (N_14831,N_14752,N_14627);
and U14832 (N_14832,N_14686,N_14610);
and U14833 (N_14833,N_14723,N_14656);
or U14834 (N_14834,N_14702,N_14766);
and U14835 (N_14835,N_14695,N_14618);
or U14836 (N_14836,N_14667,N_14724);
nand U14837 (N_14837,N_14661,N_14744);
or U14838 (N_14838,N_14631,N_14725);
nand U14839 (N_14839,N_14728,N_14736);
or U14840 (N_14840,N_14673,N_14722);
or U14841 (N_14841,N_14664,N_14617);
nand U14842 (N_14842,N_14628,N_14794);
and U14843 (N_14843,N_14742,N_14645);
and U14844 (N_14844,N_14654,N_14710);
nand U14845 (N_14845,N_14780,N_14637);
nand U14846 (N_14846,N_14697,N_14655);
or U14847 (N_14847,N_14641,N_14690);
or U14848 (N_14848,N_14605,N_14693);
nand U14849 (N_14849,N_14779,N_14759);
nor U14850 (N_14850,N_14678,N_14709);
and U14851 (N_14851,N_14760,N_14612);
and U14852 (N_14852,N_14793,N_14773);
nor U14853 (N_14853,N_14757,N_14726);
nand U14854 (N_14854,N_14679,N_14774);
xnor U14855 (N_14855,N_14676,N_14689);
xor U14856 (N_14856,N_14681,N_14767);
xor U14857 (N_14857,N_14712,N_14682);
and U14858 (N_14858,N_14703,N_14762);
or U14859 (N_14859,N_14644,N_14790);
or U14860 (N_14860,N_14615,N_14639);
or U14861 (N_14861,N_14604,N_14772);
nand U14862 (N_14862,N_14603,N_14634);
nor U14863 (N_14863,N_14688,N_14777);
nor U14864 (N_14864,N_14649,N_14721);
nor U14865 (N_14865,N_14707,N_14619);
and U14866 (N_14866,N_14748,N_14675);
xnor U14867 (N_14867,N_14727,N_14652);
nor U14868 (N_14868,N_14795,N_14630);
and U14869 (N_14869,N_14616,N_14611);
nand U14870 (N_14870,N_14796,N_14798);
or U14871 (N_14871,N_14696,N_14739);
nor U14872 (N_14872,N_14683,N_14781);
xor U14873 (N_14873,N_14608,N_14786);
nand U14874 (N_14874,N_14636,N_14601);
nor U14875 (N_14875,N_14662,N_14646);
or U14876 (N_14876,N_14799,N_14685);
nand U14877 (N_14877,N_14765,N_14740);
xnor U14878 (N_14878,N_14620,N_14704);
xor U14879 (N_14879,N_14701,N_14677);
xnor U14880 (N_14880,N_14711,N_14783);
nand U14881 (N_14881,N_14784,N_14665);
nand U14882 (N_14882,N_14651,N_14754);
nor U14883 (N_14883,N_14640,N_14791);
nand U14884 (N_14884,N_14729,N_14629);
xor U14885 (N_14885,N_14788,N_14734);
and U14886 (N_14886,N_14650,N_14716);
or U14887 (N_14887,N_14648,N_14731);
xnor U14888 (N_14888,N_14626,N_14735);
nor U14889 (N_14889,N_14642,N_14633);
or U14890 (N_14890,N_14769,N_14643);
xor U14891 (N_14891,N_14715,N_14797);
or U14892 (N_14892,N_14713,N_14763);
xor U14893 (N_14893,N_14621,N_14771);
xnor U14894 (N_14894,N_14692,N_14632);
nor U14895 (N_14895,N_14749,N_14622);
and U14896 (N_14896,N_14775,N_14660);
or U14897 (N_14897,N_14700,N_14746);
and U14898 (N_14898,N_14764,N_14782);
nor U14899 (N_14899,N_14732,N_14720);
nor U14900 (N_14900,N_14712,N_14789);
xor U14901 (N_14901,N_14722,N_14744);
xor U14902 (N_14902,N_14639,N_14702);
nand U14903 (N_14903,N_14601,N_14778);
nand U14904 (N_14904,N_14741,N_14784);
or U14905 (N_14905,N_14798,N_14748);
nor U14906 (N_14906,N_14705,N_14767);
and U14907 (N_14907,N_14742,N_14736);
nand U14908 (N_14908,N_14789,N_14797);
nand U14909 (N_14909,N_14766,N_14760);
and U14910 (N_14910,N_14633,N_14696);
or U14911 (N_14911,N_14745,N_14686);
or U14912 (N_14912,N_14795,N_14683);
and U14913 (N_14913,N_14689,N_14755);
and U14914 (N_14914,N_14609,N_14659);
and U14915 (N_14915,N_14789,N_14622);
or U14916 (N_14916,N_14611,N_14668);
nand U14917 (N_14917,N_14661,N_14768);
and U14918 (N_14918,N_14682,N_14690);
nand U14919 (N_14919,N_14747,N_14772);
xor U14920 (N_14920,N_14616,N_14770);
nand U14921 (N_14921,N_14763,N_14662);
xor U14922 (N_14922,N_14765,N_14745);
or U14923 (N_14923,N_14746,N_14680);
nor U14924 (N_14924,N_14621,N_14629);
and U14925 (N_14925,N_14705,N_14797);
nand U14926 (N_14926,N_14798,N_14600);
or U14927 (N_14927,N_14671,N_14780);
or U14928 (N_14928,N_14764,N_14631);
and U14929 (N_14929,N_14677,N_14755);
xor U14930 (N_14930,N_14615,N_14691);
xnor U14931 (N_14931,N_14715,N_14793);
nor U14932 (N_14932,N_14669,N_14681);
and U14933 (N_14933,N_14676,N_14636);
nor U14934 (N_14934,N_14687,N_14721);
nor U14935 (N_14935,N_14601,N_14715);
or U14936 (N_14936,N_14710,N_14763);
xor U14937 (N_14937,N_14752,N_14644);
nor U14938 (N_14938,N_14603,N_14783);
nand U14939 (N_14939,N_14692,N_14621);
nand U14940 (N_14940,N_14741,N_14644);
xor U14941 (N_14941,N_14736,N_14733);
or U14942 (N_14942,N_14735,N_14768);
nand U14943 (N_14943,N_14652,N_14766);
nor U14944 (N_14944,N_14676,N_14633);
xnor U14945 (N_14945,N_14667,N_14635);
or U14946 (N_14946,N_14699,N_14726);
nor U14947 (N_14947,N_14745,N_14719);
xnor U14948 (N_14948,N_14631,N_14695);
nand U14949 (N_14949,N_14654,N_14736);
xnor U14950 (N_14950,N_14786,N_14621);
xnor U14951 (N_14951,N_14647,N_14786);
and U14952 (N_14952,N_14716,N_14654);
or U14953 (N_14953,N_14655,N_14715);
and U14954 (N_14954,N_14685,N_14641);
nor U14955 (N_14955,N_14671,N_14645);
nor U14956 (N_14956,N_14720,N_14638);
or U14957 (N_14957,N_14767,N_14686);
xnor U14958 (N_14958,N_14784,N_14760);
xor U14959 (N_14959,N_14609,N_14769);
and U14960 (N_14960,N_14760,N_14712);
and U14961 (N_14961,N_14715,N_14644);
nand U14962 (N_14962,N_14619,N_14641);
xnor U14963 (N_14963,N_14672,N_14638);
or U14964 (N_14964,N_14604,N_14658);
xor U14965 (N_14965,N_14612,N_14671);
nor U14966 (N_14966,N_14642,N_14673);
or U14967 (N_14967,N_14642,N_14626);
nor U14968 (N_14968,N_14643,N_14746);
or U14969 (N_14969,N_14789,N_14780);
nand U14970 (N_14970,N_14629,N_14637);
and U14971 (N_14971,N_14649,N_14704);
nand U14972 (N_14972,N_14670,N_14715);
nor U14973 (N_14973,N_14646,N_14783);
xnor U14974 (N_14974,N_14737,N_14629);
and U14975 (N_14975,N_14765,N_14759);
and U14976 (N_14976,N_14771,N_14701);
nand U14977 (N_14977,N_14762,N_14607);
nand U14978 (N_14978,N_14736,N_14798);
or U14979 (N_14979,N_14631,N_14665);
nor U14980 (N_14980,N_14636,N_14634);
nor U14981 (N_14981,N_14671,N_14708);
and U14982 (N_14982,N_14727,N_14714);
and U14983 (N_14983,N_14606,N_14766);
and U14984 (N_14984,N_14792,N_14672);
nor U14985 (N_14985,N_14668,N_14651);
nand U14986 (N_14986,N_14760,N_14669);
xnor U14987 (N_14987,N_14765,N_14781);
and U14988 (N_14988,N_14679,N_14753);
nand U14989 (N_14989,N_14632,N_14756);
or U14990 (N_14990,N_14612,N_14785);
and U14991 (N_14991,N_14752,N_14772);
xnor U14992 (N_14992,N_14690,N_14783);
nand U14993 (N_14993,N_14604,N_14712);
xnor U14994 (N_14994,N_14645,N_14775);
nand U14995 (N_14995,N_14736,N_14768);
nand U14996 (N_14996,N_14726,N_14651);
xnor U14997 (N_14997,N_14667,N_14717);
nand U14998 (N_14998,N_14703,N_14662);
nor U14999 (N_14999,N_14683,N_14640);
nand U15000 (N_15000,N_14963,N_14933);
nand U15001 (N_15001,N_14828,N_14934);
nor U15002 (N_15002,N_14980,N_14940);
xor U15003 (N_15003,N_14982,N_14915);
and U15004 (N_15004,N_14996,N_14887);
or U15005 (N_15005,N_14895,N_14900);
nor U15006 (N_15006,N_14991,N_14876);
nand U15007 (N_15007,N_14852,N_14962);
nor U15008 (N_15008,N_14959,N_14903);
xnor U15009 (N_15009,N_14997,N_14805);
nor U15010 (N_15010,N_14822,N_14811);
xnor U15011 (N_15011,N_14918,N_14956);
nand U15012 (N_15012,N_14970,N_14836);
or U15013 (N_15013,N_14901,N_14802);
nand U15014 (N_15014,N_14814,N_14830);
nor U15015 (N_15015,N_14928,N_14889);
nor U15016 (N_15016,N_14881,N_14833);
nor U15017 (N_15017,N_14872,N_14841);
xnor U15018 (N_15018,N_14987,N_14923);
nand U15019 (N_15019,N_14864,N_14952);
nand U15020 (N_15020,N_14807,N_14943);
xor U15021 (N_15021,N_14913,N_14868);
xor U15022 (N_15022,N_14862,N_14922);
xor U15023 (N_15023,N_14831,N_14834);
nand U15024 (N_15024,N_14908,N_14914);
or U15025 (N_15025,N_14838,N_14821);
nor U15026 (N_15026,N_14939,N_14815);
or U15027 (N_15027,N_14829,N_14998);
xor U15028 (N_15028,N_14866,N_14861);
nor U15029 (N_15029,N_14867,N_14803);
xor U15030 (N_15030,N_14960,N_14850);
nor U15031 (N_15031,N_14892,N_14825);
nor U15032 (N_15032,N_14857,N_14999);
or U15033 (N_15033,N_14971,N_14869);
nor U15034 (N_15034,N_14818,N_14950);
xor U15035 (N_15035,N_14843,N_14977);
xnor U15036 (N_15036,N_14951,N_14972);
nand U15037 (N_15037,N_14804,N_14975);
xor U15038 (N_15038,N_14816,N_14974);
or U15039 (N_15039,N_14813,N_14845);
and U15040 (N_15040,N_14988,N_14871);
xnor U15041 (N_15041,N_14844,N_14819);
xnor U15042 (N_15042,N_14973,N_14877);
xor U15043 (N_15043,N_14860,N_14809);
nor U15044 (N_15044,N_14954,N_14854);
or U15045 (N_15045,N_14919,N_14808);
and U15046 (N_15046,N_14839,N_14957);
and U15047 (N_15047,N_14968,N_14945);
nor U15048 (N_15048,N_14840,N_14827);
nand U15049 (N_15049,N_14907,N_14880);
and U15050 (N_15050,N_14899,N_14992);
and U15051 (N_15051,N_14931,N_14942);
nand U15052 (N_15052,N_14964,N_14949);
nand U15053 (N_15053,N_14884,N_14883);
or U15054 (N_15054,N_14906,N_14851);
xnor U15055 (N_15055,N_14875,N_14837);
xnor U15056 (N_15056,N_14916,N_14890);
nor U15057 (N_15057,N_14978,N_14925);
xnor U15058 (N_15058,N_14885,N_14948);
or U15059 (N_15059,N_14849,N_14994);
nor U15060 (N_15060,N_14981,N_14835);
nor U15061 (N_15061,N_14966,N_14873);
nor U15062 (N_15062,N_14935,N_14863);
nand U15063 (N_15063,N_14870,N_14946);
xor U15064 (N_15064,N_14979,N_14953);
nand U15065 (N_15065,N_14955,N_14993);
and U15066 (N_15066,N_14891,N_14947);
and U15067 (N_15067,N_14878,N_14911);
and U15068 (N_15068,N_14910,N_14896);
nor U15069 (N_15069,N_14842,N_14858);
nor U15070 (N_15070,N_14920,N_14859);
nand U15071 (N_15071,N_14985,N_14921);
xnor U15072 (N_15072,N_14806,N_14995);
xnor U15073 (N_15073,N_14888,N_14847);
nor U15074 (N_15074,N_14817,N_14824);
and U15075 (N_15075,N_14823,N_14958);
nand U15076 (N_15076,N_14820,N_14905);
and U15077 (N_15077,N_14832,N_14983);
xor U15078 (N_15078,N_14929,N_14826);
or U15079 (N_15079,N_14810,N_14846);
or U15080 (N_15080,N_14853,N_14812);
and U15081 (N_15081,N_14936,N_14926);
or U15082 (N_15082,N_14856,N_14917);
nand U15083 (N_15083,N_14986,N_14961);
nor U15084 (N_15084,N_14904,N_14941);
nor U15085 (N_15085,N_14848,N_14967);
nand U15086 (N_15086,N_14894,N_14879);
or U15087 (N_15087,N_14886,N_14984);
nor U15088 (N_15088,N_14932,N_14893);
or U15089 (N_15089,N_14944,N_14930);
nand U15090 (N_15090,N_14874,N_14912);
xnor U15091 (N_15091,N_14898,N_14927);
nor U15092 (N_15092,N_14976,N_14855);
or U15093 (N_15093,N_14937,N_14801);
xnor U15094 (N_15094,N_14865,N_14965);
xor U15095 (N_15095,N_14909,N_14924);
nand U15096 (N_15096,N_14882,N_14938);
xor U15097 (N_15097,N_14969,N_14902);
or U15098 (N_15098,N_14989,N_14800);
and U15099 (N_15099,N_14897,N_14990);
and U15100 (N_15100,N_14993,N_14981);
nand U15101 (N_15101,N_14809,N_14956);
or U15102 (N_15102,N_14852,N_14885);
and U15103 (N_15103,N_14882,N_14811);
xnor U15104 (N_15104,N_14871,N_14866);
nor U15105 (N_15105,N_14887,N_14861);
nand U15106 (N_15106,N_14848,N_14942);
nand U15107 (N_15107,N_14959,N_14807);
nand U15108 (N_15108,N_14836,N_14895);
nor U15109 (N_15109,N_14965,N_14968);
and U15110 (N_15110,N_14903,N_14957);
nand U15111 (N_15111,N_14910,N_14923);
and U15112 (N_15112,N_14915,N_14853);
xor U15113 (N_15113,N_14823,N_14941);
and U15114 (N_15114,N_14831,N_14848);
xnor U15115 (N_15115,N_14819,N_14824);
nor U15116 (N_15116,N_14821,N_14858);
or U15117 (N_15117,N_14931,N_14926);
nor U15118 (N_15118,N_14923,N_14939);
nand U15119 (N_15119,N_14925,N_14985);
and U15120 (N_15120,N_14887,N_14961);
xor U15121 (N_15121,N_14810,N_14834);
nor U15122 (N_15122,N_14913,N_14818);
or U15123 (N_15123,N_14813,N_14814);
xnor U15124 (N_15124,N_14875,N_14959);
or U15125 (N_15125,N_14920,N_14963);
or U15126 (N_15126,N_14916,N_14825);
nor U15127 (N_15127,N_14974,N_14917);
xor U15128 (N_15128,N_14831,N_14938);
or U15129 (N_15129,N_14880,N_14847);
xnor U15130 (N_15130,N_14960,N_14993);
nor U15131 (N_15131,N_14938,N_14973);
xnor U15132 (N_15132,N_14864,N_14835);
and U15133 (N_15133,N_14946,N_14853);
xnor U15134 (N_15134,N_14906,N_14973);
nand U15135 (N_15135,N_14840,N_14871);
xnor U15136 (N_15136,N_14820,N_14893);
and U15137 (N_15137,N_14803,N_14940);
or U15138 (N_15138,N_14985,N_14974);
and U15139 (N_15139,N_14840,N_14917);
and U15140 (N_15140,N_14871,N_14949);
or U15141 (N_15141,N_14831,N_14837);
nand U15142 (N_15142,N_14872,N_14980);
nand U15143 (N_15143,N_14876,N_14927);
nor U15144 (N_15144,N_14866,N_14996);
nand U15145 (N_15145,N_14999,N_14978);
xnor U15146 (N_15146,N_14872,N_14963);
xor U15147 (N_15147,N_14829,N_14999);
nand U15148 (N_15148,N_14972,N_14859);
nand U15149 (N_15149,N_14845,N_14986);
nor U15150 (N_15150,N_14829,N_14932);
nand U15151 (N_15151,N_14824,N_14864);
and U15152 (N_15152,N_14871,N_14842);
nor U15153 (N_15153,N_14923,N_14977);
nor U15154 (N_15154,N_14871,N_14858);
and U15155 (N_15155,N_14817,N_14860);
and U15156 (N_15156,N_14916,N_14973);
nor U15157 (N_15157,N_14902,N_14915);
or U15158 (N_15158,N_14942,N_14917);
nand U15159 (N_15159,N_14935,N_14870);
xor U15160 (N_15160,N_14971,N_14857);
xnor U15161 (N_15161,N_14889,N_14852);
or U15162 (N_15162,N_14920,N_14857);
nand U15163 (N_15163,N_14842,N_14854);
and U15164 (N_15164,N_14919,N_14905);
nor U15165 (N_15165,N_14803,N_14971);
and U15166 (N_15166,N_14852,N_14826);
or U15167 (N_15167,N_14918,N_14972);
nand U15168 (N_15168,N_14925,N_14861);
or U15169 (N_15169,N_14823,N_14825);
and U15170 (N_15170,N_14975,N_14898);
nor U15171 (N_15171,N_14964,N_14805);
xnor U15172 (N_15172,N_14801,N_14918);
nor U15173 (N_15173,N_14948,N_14987);
xor U15174 (N_15174,N_14953,N_14911);
xor U15175 (N_15175,N_14925,N_14940);
nand U15176 (N_15176,N_14885,N_14856);
xor U15177 (N_15177,N_14877,N_14888);
nor U15178 (N_15178,N_14926,N_14862);
nor U15179 (N_15179,N_14966,N_14930);
and U15180 (N_15180,N_14838,N_14801);
nand U15181 (N_15181,N_14811,N_14896);
and U15182 (N_15182,N_14882,N_14922);
and U15183 (N_15183,N_14947,N_14888);
nand U15184 (N_15184,N_14908,N_14862);
nor U15185 (N_15185,N_14823,N_14931);
xor U15186 (N_15186,N_14965,N_14835);
or U15187 (N_15187,N_14922,N_14893);
and U15188 (N_15188,N_14911,N_14894);
and U15189 (N_15189,N_14803,N_14871);
or U15190 (N_15190,N_14834,N_14929);
or U15191 (N_15191,N_14839,N_14984);
and U15192 (N_15192,N_14992,N_14959);
and U15193 (N_15193,N_14862,N_14890);
xnor U15194 (N_15194,N_14876,N_14999);
or U15195 (N_15195,N_14995,N_14998);
nor U15196 (N_15196,N_14955,N_14996);
xor U15197 (N_15197,N_14930,N_14838);
or U15198 (N_15198,N_14802,N_14895);
nand U15199 (N_15199,N_14855,N_14819);
nand U15200 (N_15200,N_15080,N_15056);
or U15201 (N_15201,N_15127,N_15180);
or U15202 (N_15202,N_15151,N_15114);
or U15203 (N_15203,N_15007,N_15015);
nand U15204 (N_15204,N_15170,N_15154);
nor U15205 (N_15205,N_15098,N_15105);
nor U15206 (N_15206,N_15168,N_15001);
xor U15207 (N_15207,N_15031,N_15062);
nand U15208 (N_15208,N_15198,N_15178);
or U15209 (N_15209,N_15083,N_15125);
nand U15210 (N_15210,N_15057,N_15191);
xor U15211 (N_15211,N_15155,N_15163);
nand U15212 (N_15212,N_15099,N_15009);
nand U15213 (N_15213,N_15085,N_15045);
nand U15214 (N_15214,N_15189,N_15069);
nor U15215 (N_15215,N_15052,N_15013);
and U15216 (N_15216,N_15111,N_15090);
nor U15217 (N_15217,N_15108,N_15164);
nand U15218 (N_15218,N_15188,N_15120);
nor U15219 (N_15219,N_15117,N_15116);
xnor U15220 (N_15220,N_15115,N_15079);
xor U15221 (N_15221,N_15037,N_15134);
and U15222 (N_15222,N_15034,N_15072);
or U15223 (N_15223,N_15076,N_15097);
nor U15224 (N_15224,N_15089,N_15043);
nand U15225 (N_15225,N_15064,N_15035);
or U15226 (N_15226,N_15026,N_15174);
or U15227 (N_15227,N_15122,N_15137);
or U15228 (N_15228,N_15096,N_15158);
nand U15229 (N_15229,N_15106,N_15060);
nand U15230 (N_15230,N_15185,N_15047);
nand U15231 (N_15231,N_15110,N_15138);
xor U15232 (N_15232,N_15132,N_15184);
or U15233 (N_15233,N_15159,N_15103);
nor U15234 (N_15234,N_15156,N_15100);
nor U15235 (N_15235,N_15177,N_15008);
or U15236 (N_15236,N_15140,N_15181);
nand U15237 (N_15237,N_15058,N_15142);
nor U15238 (N_15238,N_15135,N_15084);
or U15239 (N_15239,N_15186,N_15148);
nor U15240 (N_15240,N_15049,N_15006);
or U15241 (N_15241,N_15065,N_15024);
or U15242 (N_15242,N_15141,N_15171);
xor U15243 (N_15243,N_15044,N_15030);
xor U15244 (N_15244,N_15102,N_15126);
xor U15245 (N_15245,N_15153,N_15067);
nand U15246 (N_15246,N_15081,N_15002);
or U15247 (N_15247,N_15162,N_15161);
xnor U15248 (N_15248,N_15165,N_15063);
nor U15249 (N_15249,N_15021,N_15073);
nor U15250 (N_15250,N_15139,N_15143);
and U15251 (N_15251,N_15183,N_15175);
nand U15252 (N_15252,N_15041,N_15051);
or U15253 (N_15253,N_15018,N_15032);
and U15254 (N_15254,N_15119,N_15130);
xor U15255 (N_15255,N_15004,N_15023);
nor U15256 (N_15256,N_15173,N_15082);
nand U15257 (N_15257,N_15123,N_15172);
xor U15258 (N_15258,N_15124,N_15169);
nand U15259 (N_15259,N_15087,N_15112);
nor U15260 (N_15260,N_15027,N_15017);
and U15261 (N_15261,N_15193,N_15094);
or U15262 (N_15262,N_15028,N_15011);
nor U15263 (N_15263,N_15022,N_15197);
nor U15264 (N_15264,N_15086,N_15118);
nand U15265 (N_15265,N_15113,N_15128);
nand U15266 (N_15266,N_15014,N_15092);
nor U15267 (N_15267,N_15131,N_15039);
xor U15268 (N_15268,N_15176,N_15061);
nor U15269 (N_15269,N_15003,N_15012);
and U15270 (N_15270,N_15187,N_15129);
or U15271 (N_15271,N_15109,N_15192);
xnor U15272 (N_15272,N_15025,N_15149);
or U15273 (N_15273,N_15071,N_15196);
or U15274 (N_15274,N_15005,N_15019);
nand U15275 (N_15275,N_15144,N_15088);
and U15276 (N_15276,N_15199,N_15074);
or U15277 (N_15277,N_15033,N_15179);
or U15278 (N_15278,N_15107,N_15195);
nand U15279 (N_15279,N_15010,N_15042);
nor U15280 (N_15280,N_15038,N_15121);
xor U15281 (N_15281,N_15016,N_15101);
or U15282 (N_15282,N_15020,N_15054);
xnor U15283 (N_15283,N_15095,N_15066);
or U15284 (N_15284,N_15046,N_15182);
xor U15285 (N_15285,N_15147,N_15029);
or U15286 (N_15286,N_15040,N_15104);
or U15287 (N_15287,N_15036,N_15157);
nand U15288 (N_15288,N_15048,N_15091);
nor U15289 (N_15289,N_15136,N_15150);
and U15290 (N_15290,N_15194,N_15053);
nor U15291 (N_15291,N_15050,N_15068);
nor U15292 (N_15292,N_15167,N_15160);
or U15293 (N_15293,N_15077,N_15133);
nor U15294 (N_15294,N_15078,N_15000);
nand U15295 (N_15295,N_15152,N_15093);
and U15296 (N_15296,N_15145,N_15059);
xor U15297 (N_15297,N_15190,N_15070);
xor U15298 (N_15298,N_15055,N_15146);
or U15299 (N_15299,N_15166,N_15075);
xor U15300 (N_15300,N_15087,N_15190);
and U15301 (N_15301,N_15124,N_15138);
and U15302 (N_15302,N_15164,N_15075);
nand U15303 (N_15303,N_15153,N_15155);
or U15304 (N_15304,N_15110,N_15140);
xnor U15305 (N_15305,N_15044,N_15130);
and U15306 (N_15306,N_15074,N_15011);
xnor U15307 (N_15307,N_15193,N_15039);
nor U15308 (N_15308,N_15015,N_15089);
xor U15309 (N_15309,N_15164,N_15133);
or U15310 (N_15310,N_15158,N_15167);
and U15311 (N_15311,N_15199,N_15005);
xor U15312 (N_15312,N_15158,N_15114);
nand U15313 (N_15313,N_15040,N_15057);
nand U15314 (N_15314,N_15129,N_15042);
xnor U15315 (N_15315,N_15195,N_15046);
or U15316 (N_15316,N_15178,N_15168);
nand U15317 (N_15317,N_15046,N_15056);
xnor U15318 (N_15318,N_15025,N_15195);
or U15319 (N_15319,N_15101,N_15057);
nand U15320 (N_15320,N_15060,N_15155);
or U15321 (N_15321,N_15083,N_15145);
and U15322 (N_15322,N_15111,N_15193);
or U15323 (N_15323,N_15161,N_15027);
and U15324 (N_15324,N_15146,N_15022);
and U15325 (N_15325,N_15053,N_15035);
and U15326 (N_15326,N_15025,N_15049);
nor U15327 (N_15327,N_15145,N_15025);
nor U15328 (N_15328,N_15084,N_15083);
xor U15329 (N_15329,N_15045,N_15136);
or U15330 (N_15330,N_15096,N_15024);
nand U15331 (N_15331,N_15090,N_15182);
and U15332 (N_15332,N_15083,N_15052);
or U15333 (N_15333,N_15034,N_15085);
xnor U15334 (N_15334,N_15104,N_15166);
nor U15335 (N_15335,N_15121,N_15134);
xnor U15336 (N_15336,N_15147,N_15028);
xor U15337 (N_15337,N_15129,N_15128);
xnor U15338 (N_15338,N_15091,N_15008);
nand U15339 (N_15339,N_15006,N_15197);
or U15340 (N_15340,N_15182,N_15123);
xor U15341 (N_15341,N_15143,N_15025);
or U15342 (N_15342,N_15124,N_15156);
or U15343 (N_15343,N_15078,N_15168);
and U15344 (N_15344,N_15179,N_15177);
nor U15345 (N_15345,N_15009,N_15073);
xnor U15346 (N_15346,N_15139,N_15037);
nand U15347 (N_15347,N_15153,N_15193);
or U15348 (N_15348,N_15019,N_15017);
xor U15349 (N_15349,N_15128,N_15061);
xor U15350 (N_15350,N_15027,N_15136);
nand U15351 (N_15351,N_15171,N_15107);
and U15352 (N_15352,N_15141,N_15137);
nor U15353 (N_15353,N_15083,N_15112);
or U15354 (N_15354,N_15081,N_15185);
nand U15355 (N_15355,N_15130,N_15022);
and U15356 (N_15356,N_15072,N_15094);
or U15357 (N_15357,N_15095,N_15080);
nand U15358 (N_15358,N_15046,N_15175);
xnor U15359 (N_15359,N_15187,N_15138);
or U15360 (N_15360,N_15047,N_15158);
nor U15361 (N_15361,N_15175,N_15044);
or U15362 (N_15362,N_15071,N_15152);
nand U15363 (N_15363,N_15123,N_15060);
and U15364 (N_15364,N_15142,N_15039);
and U15365 (N_15365,N_15066,N_15018);
or U15366 (N_15366,N_15185,N_15062);
xnor U15367 (N_15367,N_15025,N_15087);
or U15368 (N_15368,N_15106,N_15009);
nor U15369 (N_15369,N_15174,N_15150);
xnor U15370 (N_15370,N_15167,N_15077);
or U15371 (N_15371,N_15112,N_15042);
nor U15372 (N_15372,N_15096,N_15109);
nor U15373 (N_15373,N_15079,N_15076);
and U15374 (N_15374,N_15010,N_15143);
or U15375 (N_15375,N_15143,N_15061);
or U15376 (N_15376,N_15111,N_15138);
or U15377 (N_15377,N_15088,N_15032);
xor U15378 (N_15378,N_15117,N_15039);
xor U15379 (N_15379,N_15139,N_15077);
and U15380 (N_15380,N_15033,N_15078);
or U15381 (N_15381,N_15002,N_15017);
or U15382 (N_15382,N_15016,N_15142);
nor U15383 (N_15383,N_15132,N_15160);
nor U15384 (N_15384,N_15069,N_15127);
or U15385 (N_15385,N_15175,N_15132);
xnor U15386 (N_15386,N_15029,N_15154);
and U15387 (N_15387,N_15095,N_15134);
xor U15388 (N_15388,N_15109,N_15079);
xnor U15389 (N_15389,N_15102,N_15119);
or U15390 (N_15390,N_15088,N_15188);
nand U15391 (N_15391,N_15067,N_15010);
or U15392 (N_15392,N_15162,N_15192);
or U15393 (N_15393,N_15175,N_15018);
xor U15394 (N_15394,N_15031,N_15049);
nor U15395 (N_15395,N_15142,N_15108);
and U15396 (N_15396,N_15037,N_15158);
nand U15397 (N_15397,N_15162,N_15032);
xnor U15398 (N_15398,N_15044,N_15100);
or U15399 (N_15399,N_15186,N_15070);
xor U15400 (N_15400,N_15216,N_15305);
or U15401 (N_15401,N_15224,N_15328);
and U15402 (N_15402,N_15315,N_15243);
nand U15403 (N_15403,N_15375,N_15302);
xor U15404 (N_15404,N_15364,N_15272);
nor U15405 (N_15405,N_15311,N_15289);
xor U15406 (N_15406,N_15206,N_15298);
nand U15407 (N_15407,N_15210,N_15260);
or U15408 (N_15408,N_15371,N_15363);
and U15409 (N_15409,N_15285,N_15270);
xnor U15410 (N_15410,N_15335,N_15268);
xnor U15411 (N_15411,N_15265,N_15241);
and U15412 (N_15412,N_15288,N_15303);
xnor U15413 (N_15413,N_15348,N_15217);
nor U15414 (N_15414,N_15365,N_15369);
xnor U15415 (N_15415,N_15221,N_15234);
nand U15416 (N_15416,N_15319,N_15220);
xnor U15417 (N_15417,N_15337,N_15306);
nor U15418 (N_15418,N_15376,N_15238);
and U15419 (N_15419,N_15395,N_15248);
and U15420 (N_15420,N_15331,N_15361);
or U15421 (N_15421,N_15271,N_15384);
nand U15422 (N_15422,N_15326,N_15259);
and U15423 (N_15423,N_15284,N_15380);
and U15424 (N_15424,N_15230,N_15316);
or U15425 (N_15425,N_15332,N_15266);
or U15426 (N_15426,N_15249,N_15281);
or U15427 (N_15427,N_15374,N_15219);
and U15428 (N_15428,N_15334,N_15366);
or U15429 (N_15429,N_15367,N_15354);
xor U15430 (N_15430,N_15252,N_15214);
nand U15431 (N_15431,N_15352,N_15246);
xnor U15432 (N_15432,N_15263,N_15292);
nand U15433 (N_15433,N_15330,N_15229);
xor U15434 (N_15434,N_15360,N_15267);
nand U15435 (N_15435,N_15355,N_15228);
nand U15436 (N_15436,N_15342,N_15282);
and U15437 (N_15437,N_15370,N_15389);
and U15438 (N_15438,N_15207,N_15232);
nand U15439 (N_15439,N_15323,N_15231);
or U15440 (N_15440,N_15225,N_15209);
or U15441 (N_15441,N_15213,N_15353);
or U15442 (N_15442,N_15312,N_15279);
or U15443 (N_15443,N_15222,N_15280);
nor U15444 (N_15444,N_15308,N_15227);
nor U15445 (N_15445,N_15287,N_15347);
xnor U15446 (N_15446,N_15293,N_15318);
xor U15447 (N_15447,N_15327,N_15264);
and U15448 (N_15448,N_15373,N_15394);
nor U15449 (N_15449,N_15340,N_15383);
nor U15450 (N_15450,N_15208,N_15235);
or U15451 (N_15451,N_15237,N_15388);
and U15452 (N_15452,N_15301,N_15275);
xnor U15453 (N_15453,N_15368,N_15346);
or U15454 (N_15454,N_15254,N_15256);
and U15455 (N_15455,N_15325,N_15276);
xor U15456 (N_15456,N_15215,N_15244);
xnor U15457 (N_15457,N_15398,N_15212);
or U15458 (N_15458,N_15290,N_15313);
nor U15459 (N_15459,N_15299,N_15205);
xnor U15460 (N_15460,N_15204,N_15223);
and U15461 (N_15461,N_15286,N_15341);
or U15462 (N_15462,N_15350,N_15251);
and U15463 (N_15463,N_15240,N_15333);
and U15464 (N_15464,N_15203,N_15250);
or U15465 (N_15465,N_15258,N_15317);
and U15466 (N_15466,N_15245,N_15218);
nand U15467 (N_15467,N_15300,N_15283);
and U15468 (N_15468,N_15255,N_15377);
or U15469 (N_15469,N_15320,N_15385);
and U15470 (N_15470,N_15357,N_15202);
nor U15471 (N_15471,N_15322,N_15297);
or U15472 (N_15472,N_15307,N_15321);
xor U15473 (N_15473,N_15304,N_15344);
xnor U15474 (N_15474,N_15349,N_15278);
xor U15475 (N_15475,N_15236,N_15233);
nand U15476 (N_15476,N_15339,N_15392);
and U15477 (N_15477,N_15396,N_15291);
and U15478 (N_15478,N_15269,N_15390);
nor U15479 (N_15479,N_15329,N_15274);
nor U15480 (N_15480,N_15247,N_15356);
and U15481 (N_15481,N_15242,N_15257);
or U15482 (N_15482,N_15273,N_15399);
xor U15483 (N_15483,N_15239,N_15253);
or U15484 (N_15484,N_15358,N_15387);
nor U15485 (N_15485,N_15379,N_15336);
nor U15486 (N_15486,N_15382,N_15296);
nand U15487 (N_15487,N_15378,N_15351);
nand U15488 (N_15488,N_15200,N_15314);
nand U15489 (N_15489,N_15261,N_15226);
xnor U15490 (N_15490,N_15362,N_15391);
nor U15491 (N_15491,N_15211,N_15397);
nand U15492 (N_15492,N_15262,N_15386);
or U15493 (N_15493,N_15359,N_15345);
nor U15494 (N_15494,N_15381,N_15310);
xnor U15495 (N_15495,N_15393,N_15277);
and U15496 (N_15496,N_15324,N_15295);
nor U15497 (N_15497,N_15372,N_15201);
nand U15498 (N_15498,N_15338,N_15309);
and U15499 (N_15499,N_15294,N_15343);
or U15500 (N_15500,N_15200,N_15333);
xnor U15501 (N_15501,N_15321,N_15266);
nor U15502 (N_15502,N_15205,N_15355);
and U15503 (N_15503,N_15337,N_15283);
nor U15504 (N_15504,N_15214,N_15263);
and U15505 (N_15505,N_15356,N_15203);
nand U15506 (N_15506,N_15231,N_15377);
nor U15507 (N_15507,N_15367,N_15381);
nand U15508 (N_15508,N_15384,N_15364);
or U15509 (N_15509,N_15362,N_15246);
nand U15510 (N_15510,N_15276,N_15254);
nor U15511 (N_15511,N_15265,N_15310);
and U15512 (N_15512,N_15266,N_15342);
nand U15513 (N_15513,N_15246,N_15226);
or U15514 (N_15514,N_15348,N_15259);
and U15515 (N_15515,N_15293,N_15255);
and U15516 (N_15516,N_15390,N_15374);
nor U15517 (N_15517,N_15328,N_15391);
and U15518 (N_15518,N_15209,N_15288);
or U15519 (N_15519,N_15214,N_15369);
and U15520 (N_15520,N_15242,N_15366);
nor U15521 (N_15521,N_15235,N_15326);
xnor U15522 (N_15522,N_15256,N_15369);
nor U15523 (N_15523,N_15210,N_15388);
nor U15524 (N_15524,N_15272,N_15399);
xor U15525 (N_15525,N_15357,N_15229);
nand U15526 (N_15526,N_15225,N_15230);
and U15527 (N_15527,N_15288,N_15314);
or U15528 (N_15528,N_15325,N_15352);
nor U15529 (N_15529,N_15365,N_15390);
xnor U15530 (N_15530,N_15341,N_15308);
and U15531 (N_15531,N_15359,N_15381);
nand U15532 (N_15532,N_15290,N_15385);
or U15533 (N_15533,N_15292,N_15295);
xor U15534 (N_15534,N_15342,N_15378);
xnor U15535 (N_15535,N_15379,N_15340);
or U15536 (N_15536,N_15204,N_15304);
nor U15537 (N_15537,N_15346,N_15315);
xnor U15538 (N_15538,N_15369,N_15366);
nand U15539 (N_15539,N_15306,N_15223);
nand U15540 (N_15540,N_15327,N_15274);
and U15541 (N_15541,N_15387,N_15283);
or U15542 (N_15542,N_15272,N_15233);
xor U15543 (N_15543,N_15228,N_15361);
nand U15544 (N_15544,N_15346,N_15326);
and U15545 (N_15545,N_15326,N_15358);
or U15546 (N_15546,N_15398,N_15379);
xnor U15547 (N_15547,N_15380,N_15334);
and U15548 (N_15548,N_15341,N_15226);
xor U15549 (N_15549,N_15243,N_15274);
or U15550 (N_15550,N_15257,N_15320);
or U15551 (N_15551,N_15322,N_15302);
nand U15552 (N_15552,N_15395,N_15266);
nor U15553 (N_15553,N_15361,N_15390);
nand U15554 (N_15554,N_15276,N_15244);
xnor U15555 (N_15555,N_15385,N_15294);
and U15556 (N_15556,N_15393,N_15315);
or U15557 (N_15557,N_15235,N_15348);
xor U15558 (N_15558,N_15243,N_15232);
and U15559 (N_15559,N_15335,N_15295);
nand U15560 (N_15560,N_15371,N_15267);
or U15561 (N_15561,N_15352,N_15301);
and U15562 (N_15562,N_15376,N_15260);
or U15563 (N_15563,N_15212,N_15279);
and U15564 (N_15564,N_15227,N_15217);
nand U15565 (N_15565,N_15206,N_15327);
or U15566 (N_15566,N_15364,N_15360);
nand U15567 (N_15567,N_15317,N_15362);
or U15568 (N_15568,N_15202,N_15209);
or U15569 (N_15569,N_15329,N_15359);
or U15570 (N_15570,N_15303,N_15269);
nand U15571 (N_15571,N_15277,N_15300);
nand U15572 (N_15572,N_15245,N_15349);
nor U15573 (N_15573,N_15257,N_15294);
nand U15574 (N_15574,N_15367,N_15304);
nand U15575 (N_15575,N_15247,N_15344);
or U15576 (N_15576,N_15351,N_15208);
nor U15577 (N_15577,N_15208,N_15215);
nor U15578 (N_15578,N_15215,N_15333);
xnor U15579 (N_15579,N_15204,N_15337);
xor U15580 (N_15580,N_15303,N_15249);
nor U15581 (N_15581,N_15308,N_15289);
nor U15582 (N_15582,N_15312,N_15334);
xor U15583 (N_15583,N_15243,N_15283);
nand U15584 (N_15584,N_15298,N_15209);
nor U15585 (N_15585,N_15213,N_15326);
nor U15586 (N_15586,N_15326,N_15344);
nor U15587 (N_15587,N_15378,N_15259);
and U15588 (N_15588,N_15217,N_15257);
and U15589 (N_15589,N_15301,N_15375);
and U15590 (N_15590,N_15335,N_15350);
nand U15591 (N_15591,N_15281,N_15273);
xnor U15592 (N_15592,N_15359,N_15238);
nand U15593 (N_15593,N_15309,N_15289);
and U15594 (N_15594,N_15285,N_15344);
or U15595 (N_15595,N_15203,N_15379);
and U15596 (N_15596,N_15261,N_15306);
xnor U15597 (N_15597,N_15246,N_15255);
xor U15598 (N_15598,N_15365,N_15326);
nand U15599 (N_15599,N_15207,N_15324);
or U15600 (N_15600,N_15501,N_15436);
or U15601 (N_15601,N_15554,N_15408);
nand U15602 (N_15602,N_15583,N_15472);
and U15603 (N_15603,N_15407,N_15461);
xor U15604 (N_15604,N_15449,N_15468);
xnor U15605 (N_15605,N_15537,N_15568);
xor U15606 (N_15606,N_15434,N_15464);
and U15607 (N_15607,N_15497,N_15591);
xnor U15608 (N_15608,N_15532,N_15420);
xor U15609 (N_15609,N_15540,N_15453);
and U15610 (N_15610,N_15585,N_15596);
nand U15611 (N_15611,N_15418,N_15504);
xor U15612 (N_15612,N_15470,N_15432);
nand U15613 (N_15613,N_15471,N_15482);
xnor U15614 (N_15614,N_15452,N_15409);
or U15615 (N_15615,N_15512,N_15490);
and U15616 (N_15616,N_15435,N_15503);
nand U15617 (N_15617,N_15431,N_15574);
and U15618 (N_15618,N_15410,N_15401);
nor U15619 (N_15619,N_15575,N_15582);
nor U15620 (N_15620,N_15493,N_15522);
nand U15621 (N_15621,N_15424,N_15533);
nor U15622 (N_15622,N_15539,N_15567);
nor U15623 (N_15623,N_15538,N_15473);
nand U15624 (N_15624,N_15589,N_15505);
or U15625 (N_15625,N_15444,N_15515);
xor U15626 (N_15626,N_15403,N_15508);
nand U15627 (N_15627,N_15428,N_15555);
xor U15628 (N_15628,N_15513,N_15477);
nor U15629 (N_15629,N_15523,N_15581);
nor U15630 (N_15630,N_15599,N_15566);
xor U15631 (N_15631,N_15579,N_15463);
nor U15632 (N_15632,N_15536,N_15587);
nor U15633 (N_15633,N_15570,N_15433);
xnor U15634 (N_15634,N_15478,N_15479);
and U15635 (N_15635,N_15443,N_15483);
nand U15636 (N_15636,N_15518,N_15430);
and U15637 (N_15637,N_15400,N_15475);
nor U15638 (N_15638,N_15456,N_15429);
and U15639 (N_15639,N_15507,N_15416);
xor U15640 (N_15640,N_15516,N_15551);
xor U15641 (N_15641,N_15588,N_15531);
and U15642 (N_15642,N_15499,N_15586);
nor U15643 (N_15643,N_15524,N_15469);
nand U15644 (N_15644,N_15406,N_15423);
nand U15645 (N_15645,N_15467,N_15447);
nor U15646 (N_15646,N_15562,N_15534);
or U15647 (N_15647,N_15510,N_15543);
nand U15648 (N_15648,N_15451,N_15550);
or U15649 (N_15649,N_15506,N_15526);
nor U15650 (N_15650,N_15542,N_15549);
xnor U15651 (N_15651,N_15419,N_15577);
nand U15652 (N_15652,N_15553,N_15442);
nor U15653 (N_15653,N_15525,N_15414);
nor U15654 (N_15654,N_15561,N_15421);
or U15655 (N_15655,N_15500,N_15440);
and U15656 (N_15656,N_15489,N_15590);
or U15657 (N_15657,N_15557,N_15564);
nor U15658 (N_15658,N_15474,N_15511);
xor U15659 (N_15659,N_15597,N_15520);
or U15660 (N_15660,N_15572,N_15573);
and U15661 (N_15661,N_15441,N_15446);
xnor U15662 (N_15662,N_15563,N_15584);
and U15663 (N_15663,N_15455,N_15546);
and U15664 (N_15664,N_15495,N_15445);
nor U15665 (N_15665,N_15481,N_15415);
and U15666 (N_15666,N_15496,N_15454);
xnor U15667 (N_15667,N_15422,N_15517);
and U15668 (N_15668,N_15576,N_15498);
nor U15669 (N_15669,N_15411,N_15535);
xor U15670 (N_15670,N_15527,N_15502);
xor U15671 (N_15671,N_15412,N_15488);
xor U15672 (N_15672,N_15460,N_15465);
nand U15673 (N_15673,N_15413,N_15578);
xor U15674 (N_15674,N_15528,N_15598);
nand U15675 (N_15675,N_15565,N_15494);
or U15676 (N_15676,N_15484,N_15558);
or U15677 (N_15677,N_15458,N_15426);
and U15678 (N_15678,N_15548,N_15457);
and U15679 (N_15679,N_15486,N_15437);
and U15680 (N_15680,N_15559,N_15476);
xnor U15681 (N_15681,N_15466,N_15462);
nand U15682 (N_15682,N_15593,N_15519);
or U15683 (N_15683,N_15592,N_15530);
nand U15684 (N_15684,N_15492,N_15402);
or U15685 (N_15685,N_15580,N_15480);
xor U15686 (N_15686,N_15417,N_15404);
nor U15687 (N_15687,N_15487,N_15491);
xnor U15688 (N_15688,N_15514,N_15595);
or U15689 (N_15689,N_15556,N_15547);
or U15690 (N_15690,N_15541,N_15571);
nor U15691 (N_15691,N_15438,N_15448);
and U15692 (N_15692,N_15425,N_15450);
or U15693 (N_15693,N_15545,N_15427);
nand U15694 (N_15694,N_15552,N_15544);
and U15695 (N_15695,N_15521,N_15405);
and U15696 (N_15696,N_15485,N_15459);
nand U15697 (N_15697,N_15560,N_15439);
nand U15698 (N_15698,N_15509,N_15529);
xor U15699 (N_15699,N_15569,N_15594);
or U15700 (N_15700,N_15442,N_15531);
and U15701 (N_15701,N_15557,N_15443);
nand U15702 (N_15702,N_15407,N_15559);
nor U15703 (N_15703,N_15516,N_15502);
nor U15704 (N_15704,N_15423,N_15474);
and U15705 (N_15705,N_15410,N_15578);
nand U15706 (N_15706,N_15464,N_15433);
xor U15707 (N_15707,N_15534,N_15461);
nor U15708 (N_15708,N_15518,N_15442);
xor U15709 (N_15709,N_15468,N_15442);
and U15710 (N_15710,N_15557,N_15430);
xnor U15711 (N_15711,N_15439,N_15479);
nor U15712 (N_15712,N_15442,N_15592);
or U15713 (N_15713,N_15580,N_15584);
and U15714 (N_15714,N_15501,N_15490);
nor U15715 (N_15715,N_15494,N_15577);
nor U15716 (N_15716,N_15547,N_15535);
xnor U15717 (N_15717,N_15505,N_15588);
xor U15718 (N_15718,N_15466,N_15494);
nor U15719 (N_15719,N_15588,N_15571);
and U15720 (N_15720,N_15582,N_15521);
xnor U15721 (N_15721,N_15535,N_15461);
xnor U15722 (N_15722,N_15433,N_15460);
nor U15723 (N_15723,N_15443,N_15479);
nor U15724 (N_15724,N_15437,N_15587);
xor U15725 (N_15725,N_15516,N_15430);
xor U15726 (N_15726,N_15505,N_15411);
nand U15727 (N_15727,N_15554,N_15428);
xor U15728 (N_15728,N_15460,N_15463);
nor U15729 (N_15729,N_15400,N_15593);
nand U15730 (N_15730,N_15549,N_15498);
xnor U15731 (N_15731,N_15519,N_15518);
nor U15732 (N_15732,N_15455,N_15592);
and U15733 (N_15733,N_15504,N_15577);
and U15734 (N_15734,N_15563,N_15470);
nor U15735 (N_15735,N_15407,N_15526);
or U15736 (N_15736,N_15469,N_15486);
nor U15737 (N_15737,N_15567,N_15542);
or U15738 (N_15738,N_15518,N_15594);
xor U15739 (N_15739,N_15574,N_15527);
nand U15740 (N_15740,N_15592,N_15405);
nor U15741 (N_15741,N_15524,N_15599);
nand U15742 (N_15742,N_15592,N_15571);
xor U15743 (N_15743,N_15495,N_15543);
or U15744 (N_15744,N_15552,N_15554);
nor U15745 (N_15745,N_15545,N_15491);
or U15746 (N_15746,N_15597,N_15563);
or U15747 (N_15747,N_15461,N_15493);
xnor U15748 (N_15748,N_15409,N_15568);
nor U15749 (N_15749,N_15441,N_15424);
or U15750 (N_15750,N_15594,N_15552);
nor U15751 (N_15751,N_15580,N_15539);
xor U15752 (N_15752,N_15523,N_15460);
and U15753 (N_15753,N_15535,N_15444);
and U15754 (N_15754,N_15571,N_15578);
nand U15755 (N_15755,N_15591,N_15496);
or U15756 (N_15756,N_15565,N_15554);
nor U15757 (N_15757,N_15436,N_15508);
or U15758 (N_15758,N_15435,N_15418);
and U15759 (N_15759,N_15419,N_15447);
nor U15760 (N_15760,N_15482,N_15424);
and U15761 (N_15761,N_15552,N_15530);
xor U15762 (N_15762,N_15481,N_15509);
nor U15763 (N_15763,N_15506,N_15558);
and U15764 (N_15764,N_15569,N_15527);
xnor U15765 (N_15765,N_15421,N_15526);
and U15766 (N_15766,N_15435,N_15455);
or U15767 (N_15767,N_15405,N_15530);
nand U15768 (N_15768,N_15568,N_15581);
xor U15769 (N_15769,N_15547,N_15433);
nor U15770 (N_15770,N_15532,N_15459);
xnor U15771 (N_15771,N_15507,N_15423);
nand U15772 (N_15772,N_15441,N_15599);
nor U15773 (N_15773,N_15476,N_15426);
nor U15774 (N_15774,N_15404,N_15518);
nor U15775 (N_15775,N_15483,N_15539);
and U15776 (N_15776,N_15438,N_15588);
xor U15777 (N_15777,N_15463,N_15580);
nor U15778 (N_15778,N_15444,N_15510);
and U15779 (N_15779,N_15474,N_15524);
nand U15780 (N_15780,N_15564,N_15597);
nand U15781 (N_15781,N_15578,N_15431);
or U15782 (N_15782,N_15581,N_15462);
nor U15783 (N_15783,N_15403,N_15471);
or U15784 (N_15784,N_15472,N_15592);
or U15785 (N_15785,N_15493,N_15455);
and U15786 (N_15786,N_15490,N_15599);
and U15787 (N_15787,N_15586,N_15458);
nand U15788 (N_15788,N_15578,N_15427);
and U15789 (N_15789,N_15543,N_15401);
nor U15790 (N_15790,N_15478,N_15464);
or U15791 (N_15791,N_15554,N_15466);
nor U15792 (N_15792,N_15574,N_15566);
nand U15793 (N_15793,N_15474,N_15541);
or U15794 (N_15794,N_15544,N_15474);
nand U15795 (N_15795,N_15585,N_15526);
and U15796 (N_15796,N_15560,N_15444);
nand U15797 (N_15797,N_15538,N_15510);
nand U15798 (N_15798,N_15551,N_15544);
nand U15799 (N_15799,N_15507,N_15558);
nand U15800 (N_15800,N_15666,N_15668);
nand U15801 (N_15801,N_15787,N_15675);
or U15802 (N_15802,N_15721,N_15771);
nand U15803 (N_15803,N_15791,N_15713);
or U15804 (N_15804,N_15778,N_15611);
and U15805 (N_15805,N_15730,N_15773);
nor U15806 (N_15806,N_15677,N_15639);
or U15807 (N_15807,N_15687,N_15711);
xnor U15808 (N_15808,N_15732,N_15705);
or U15809 (N_15809,N_15647,N_15609);
nand U15810 (N_15810,N_15694,N_15758);
and U15811 (N_15811,N_15699,N_15784);
or U15812 (N_15812,N_15757,N_15738);
xnor U15813 (N_15813,N_15670,N_15672);
nor U15814 (N_15814,N_15712,N_15616);
and U15815 (N_15815,N_15655,N_15736);
nor U15816 (N_15816,N_15674,N_15688);
nand U15817 (N_15817,N_15697,N_15710);
nand U15818 (N_15818,N_15660,N_15614);
and U15819 (N_15819,N_15799,N_15658);
and U15820 (N_15820,N_15613,N_15605);
xnor U15821 (N_15821,N_15717,N_15622);
and U15822 (N_15822,N_15750,N_15681);
or U15823 (N_15823,N_15715,N_15630);
nor U15824 (N_15824,N_15663,N_15780);
xor U15825 (N_15825,N_15650,N_15608);
or U15826 (N_15826,N_15649,N_15706);
and U15827 (N_15827,N_15689,N_15684);
and U15828 (N_15828,N_15797,N_15770);
or U15829 (N_15829,N_15753,N_15623);
and U15830 (N_15830,N_15762,N_15634);
nand U15831 (N_15831,N_15740,N_15765);
and U15832 (N_15832,N_15610,N_15628);
nor U15833 (N_15833,N_15745,N_15627);
nor U15834 (N_15834,N_15619,N_15748);
and U15835 (N_15835,N_15783,N_15716);
nand U15836 (N_15836,N_15781,N_15662);
nor U15837 (N_15837,N_15648,N_15632);
xnor U15838 (N_15838,N_15708,N_15625);
nand U15839 (N_15839,N_15602,N_15626);
or U15840 (N_15840,N_15743,N_15734);
nand U15841 (N_15841,N_15788,N_15742);
or U15842 (N_15842,N_15604,N_15798);
and U15843 (N_15843,N_15646,N_15794);
and U15844 (N_15844,N_15657,N_15665);
nor U15845 (N_15845,N_15775,N_15659);
or U15846 (N_15846,N_15790,N_15772);
nand U15847 (N_15847,N_15620,N_15737);
and U15848 (N_15848,N_15752,N_15680);
xor U15849 (N_15849,N_15685,N_15618);
or U15850 (N_15850,N_15673,N_15769);
and U15851 (N_15851,N_15703,N_15640);
nand U15852 (N_15852,N_15637,N_15603);
nor U15853 (N_15853,N_15629,N_15723);
nor U15854 (N_15854,N_15661,N_15636);
nand U15855 (N_15855,N_15682,N_15755);
xnor U15856 (N_15856,N_15767,N_15671);
xor U15857 (N_15857,N_15641,N_15759);
xor U15858 (N_15858,N_15692,N_15731);
xor U15859 (N_15859,N_15756,N_15676);
or U15860 (N_15860,N_15701,N_15600);
xnor U15861 (N_15861,N_15669,N_15607);
nand U15862 (N_15862,N_15601,N_15621);
nor U15863 (N_15863,N_15709,N_15792);
or U15864 (N_15864,N_15795,N_15645);
nand U15865 (N_15865,N_15764,N_15631);
nand U15866 (N_15866,N_15763,N_15786);
or U15867 (N_15867,N_15777,N_15683);
xnor U15868 (N_15868,N_15638,N_15739);
and U15869 (N_15869,N_15735,N_15768);
and U15870 (N_15870,N_15667,N_15664);
and U15871 (N_15871,N_15754,N_15643);
nor U15872 (N_15872,N_15774,N_15766);
nor U15873 (N_15873,N_15624,N_15652);
nor U15874 (N_15874,N_15633,N_15690);
nor U15875 (N_15875,N_15744,N_15727);
nor U15876 (N_15876,N_15704,N_15693);
or U15877 (N_15877,N_15733,N_15729);
nand U15878 (N_15878,N_15707,N_15635);
or U15879 (N_15879,N_15718,N_15702);
nand U15880 (N_15880,N_15696,N_15679);
or U15881 (N_15881,N_15700,N_15642);
xor U15882 (N_15882,N_15695,N_15644);
or U15883 (N_15883,N_15698,N_15776);
or U15884 (N_15884,N_15686,N_15615);
nand U15885 (N_15885,N_15722,N_15793);
nand U15886 (N_15886,N_15720,N_15741);
and U15887 (N_15887,N_15785,N_15728);
and U15888 (N_15888,N_15761,N_15719);
or U15889 (N_15889,N_15656,N_15796);
or U15890 (N_15890,N_15782,N_15653);
xor U15891 (N_15891,N_15747,N_15714);
nand U15892 (N_15892,N_15654,N_15751);
nand U15893 (N_15893,N_15779,N_15651);
and U15894 (N_15894,N_15606,N_15678);
nor U15895 (N_15895,N_15749,N_15760);
nor U15896 (N_15896,N_15725,N_15746);
or U15897 (N_15897,N_15724,N_15612);
nand U15898 (N_15898,N_15617,N_15726);
xnor U15899 (N_15899,N_15789,N_15691);
and U15900 (N_15900,N_15629,N_15691);
or U15901 (N_15901,N_15774,N_15645);
nor U15902 (N_15902,N_15780,N_15740);
nor U15903 (N_15903,N_15736,N_15788);
nand U15904 (N_15904,N_15790,N_15603);
nand U15905 (N_15905,N_15712,N_15781);
and U15906 (N_15906,N_15668,N_15634);
nand U15907 (N_15907,N_15777,N_15730);
nor U15908 (N_15908,N_15625,N_15638);
nand U15909 (N_15909,N_15664,N_15662);
xor U15910 (N_15910,N_15671,N_15658);
and U15911 (N_15911,N_15611,N_15640);
nand U15912 (N_15912,N_15616,N_15625);
or U15913 (N_15913,N_15739,N_15793);
nor U15914 (N_15914,N_15750,N_15724);
xor U15915 (N_15915,N_15639,N_15734);
nor U15916 (N_15916,N_15611,N_15783);
nand U15917 (N_15917,N_15664,N_15659);
xor U15918 (N_15918,N_15755,N_15715);
nand U15919 (N_15919,N_15607,N_15722);
and U15920 (N_15920,N_15673,N_15614);
and U15921 (N_15921,N_15665,N_15747);
nor U15922 (N_15922,N_15768,N_15770);
nand U15923 (N_15923,N_15619,N_15711);
xor U15924 (N_15924,N_15611,N_15704);
or U15925 (N_15925,N_15788,N_15671);
nor U15926 (N_15926,N_15756,N_15791);
nand U15927 (N_15927,N_15682,N_15605);
nor U15928 (N_15928,N_15785,N_15680);
xnor U15929 (N_15929,N_15735,N_15747);
or U15930 (N_15930,N_15768,N_15694);
or U15931 (N_15931,N_15775,N_15731);
nand U15932 (N_15932,N_15665,N_15653);
xnor U15933 (N_15933,N_15660,N_15696);
xor U15934 (N_15934,N_15760,N_15627);
nand U15935 (N_15935,N_15612,N_15743);
nor U15936 (N_15936,N_15737,N_15655);
and U15937 (N_15937,N_15773,N_15799);
xnor U15938 (N_15938,N_15755,N_15708);
or U15939 (N_15939,N_15615,N_15681);
and U15940 (N_15940,N_15767,N_15622);
and U15941 (N_15941,N_15656,N_15672);
nand U15942 (N_15942,N_15622,N_15604);
and U15943 (N_15943,N_15656,N_15776);
nand U15944 (N_15944,N_15645,N_15628);
nor U15945 (N_15945,N_15673,N_15606);
xnor U15946 (N_15946,N_15695,N_15639);
or U15947 (N_15947,N_15753,N_15763);
and U15948 (N_15948,N_15761,N_15718);
xnor U15949 (N_15949,N_15699,N_15701);
nor U15950 (N_15950,N_15730,N_15797);
nand U15951 (N_15951,N_15720,N_15666);
xnor U15952 (N_15952,N_15722,N_15654);
xnor U15953 (N_15953,N_15760,N_15797);
or U15954 (N_15954,N_15600,N_15794);
nor U15955 (N_15955,N_15703,N_15603);
and U15956 (N_15956,N_15689,N_15798);
and U15957 (N_15957,N_15688,N_15620);
nor U15958 (N_15958,N_15690,N_15652);
nand U15959 (N_15959,N_15645,N_15689);
xor U15960 (N_15960,N_15640,N_15760);
xor U15961 (N_15961,N_15719,N_15687);
nand U15962 (N_15962,N_15680,N_15668);
nand U15963 (N_15963,N_15646,N_15629);
xor U15964 (N_15964,N_15720,N_15778);
xor U15965 (N_15965,N_15749,N_15675);
nand U15966 (N_15966,N_15736,N_15705);
nor U15967 (N_15967,N_15683,N_15752);
xor U15968 (N_15968,N_15676,N_15608);
nor U15969 (N_15969,N_15717,N_15791);
or U15970 (N_15970,N_15679,N_15758);
and U15971 (N_15971,N_15799,N_15621);
and U15972 (N_15972,N_15782,N_15710);
and U15973 (N_15973,N_15629,N_15765);
nand U15974 (N_15974,N_15727,N_15749);
or U15975 (N_15975,N_15795,N_15610);
xor U15976 (N_15976,N_15759,N_15620);
xnor U15977 (N_15977,N_15783,N_15678);
nand U15978 (N_15978,N_15669,N_15717);
or U15979 (N_15979,N_15754,N_15647);
and U15980 (N_15980,N_15771,N_15608);
or U15981 (N_15981,N_15732,N_15608);
nand U15982 (N_15982,N_15648,N_15775);
and U15983 (N_15983,N_15725,N_15701);
nor U15984 (N_15984,N_15700,N_15684);
or U15985 (N_15985,N_15600,N_15667);
nand U15986 (N_15986,N_15711,N_15720);
or U15987 (N_15987,N_15621,N_15654);
nor U15988 (N_15988,N_15709,N_15606);
xnor U15989 (N_15989,N_15701,N_15615);
nand U15990 (N_15990,N_15664,N_15713);
and U15991 (N_15991,N_15684,N_15602);
nor U15992 (N_15992,N_15616,N_15643);
or U15993 (N_15993,N_15789,N_15604);
nor U15994 (N_15994,N_15786,N_15798);
xor U15995 (N_15995,N_15687,N_15613);
xnor U15996 (N_15996,N_15692,N_15653);
or U15997 (N_15997,N_15639,N_15751);
xor U15998 (N_15998,N_15743,N_15712);
and U15999 (N_15999,N_15651,N_15623);
nand U16000 (N_16000,N_15945,N_15993);
nor U16001 (N_16001,N_15846,N_15951);
nor U16002 (N_16002,N_15849,N_15841);
and U16003 (N_16003,N_15880,N_15861);
and U16004 (N_16004,N_15997,N_15874);
xnor U16005 (N_16005,N_15952,N_15992);
and U16006 (N_16006,N_15838,N_15912);
or U16007 (N_16007,N_15812,N_15872);
xnor U16008 (N_16008,N_15928,N_15976);
xnor U16009 (N_16009,N_15826,N_15831);
xnor U16010 (N_16010,N_15907,N_15863);
nand U16011 (N_16011,N_15851,N_15921);
nand U16012 (N_16012,N_15873,N_15927);
nand U16013 (N_16013,N_15914,N_15837);
nand U16014 (N_16014,N_15821,N_15867);
and U16015 (N_16015,N_15913,N_15991);
nand U16016 (N_16016,N_15978,N_15972);
nand U16017 (N_16017,N_15998,N_15871);
nor U16018 (N_16018,N_15870,N_15816);
xnor U16019 (N_16019,N_15848,N_15930);
and U16020 (N_16020,N_15943,N_15920);
nand U16021 (N_16021,N_15859,N_15917);
xor U16022 (N_16022,N_15832,N_15807);
or U16023 (N_16023,N_15982,N_15967);
nand U16024 (N_16024,N_15809,N_15903);
xnor U16025 (N_16025,N_15990,N_15953);
xnor U16026 (N_16026,N_15802,N_15989);
or U16027 (N_16027,N_15966,N_15987);
and U16028 (N_16028,N_15825,N_15895);
nor U16029 (N_16029,N_15855,N_15941);
xor U16030 (N_16030,N_15915,N_15847);
and U16031 (N_16031,N_15836,N_15877);
nor U16032 (N_16032,N_15957,N_15853);
nand U16033 (N_16033,N_15889,N_15984);
or U16034 (N_16034,N_15822,N_15828);
xnor U16035 (N_16035,N_15891,N_15910);
and U16036 (N_16036,N_15918,N_15902);
and U16037 (N_16037,N_15942,N_15840);
nand U16038 (N_16038,N_15916,N_15850);
and U16039 (N_16039,N_15980,N_15815);
and U16040 (N_16040,N_15904,N_15814);
nand U16041 (N_16041,N_15973,N_15959);
xnor U16042 (N_16042,N_15926,N_15835);
xnor U16043 (N_16043,N_15864,N_15933);
xnor U16044 (N_16044,N_15875,N_15968);
and U16045 (N_16045,N_15883,N_15884);
nand U16046 (N_16046,N_15955,N_15862);
nand U16047 (N_16047,N_15900,N_15857);
or U16048 (N_16048,N_15885,N_15886);
nor U16049 (N_16049,N_15954,N_15813);
or U16050 (N_16050,N_15824,N_15964);
or U16051 (N_16051,N_15881,N_15843);
nand U16052 (N_16052,N_15975,N_15974);
nand U16053 (N_16053,N_15898,N_15839);
and U16054 (N_16054,N_15996,N_15810);
xor U16055 (N_16055,N_15823,N_15808);
nand U16056 (N_16056,N_15932,N_15890);
or U16057 (N_16057,N_15925,N_15858);
nor U16058 (N_16058,N_15946,N_15985);
nand U16059 (N_16059,N_15944,N_15894);
or U16060 (N_16060,N_15937,N_15938);
nand U16061 (N_16061,N_15970,N_15923);
xor U16062 (N_16062,N_15929,N_15827);
nand U16063 (N_16063,N_15844,N_15979);
nor U16064 (N_16064,N_15963,N_15830);
xor U16065 (N_16065,N_15804,N_15866);
and U16066 (N_16066,N_15856,N_15893);
or U16067 (N_16067,N_15892,N_15833);
xnor U16068 (N_16068,N_15800,N_15948);
xnor U16069 (N_16069,N_15962,N_15934);
xnor U16070 (N_16070,N_15956,N_15834);
nand U16071 (N_16071,N_15947,N_15819);
nand U16072 (N_16072,N_15801,N_15977);
and U16073 (N_16073,N_15854,N_15960);
and U16074 (N_16074,N_15888,N_15899);
and U16075 (N_16075,N_15965,N_15896);
xor U16076 (N_16076,N_15887,N_15924);
or U16077 (N_16077,N_15879,N_15983);
nand U16078 (N_16078,N_15922,N_15897);
xor U16079 (N_16079,N_15852,N_15919);
nor U16080 (N_16080,N_15905,N_15869);
and U16081 (N_16081,N_15876,N_15820);
or U16082 (N_16082,N_15994,N_15878);
nand U16083 (N_16083,N_15803,N_15806);
nand U16084 (N_16084,N_15817,N_15969);
xor U16085 (N_16085,N_15865,N_15971);
xor U16086 (N_16086,N_15845,N_15901);
nand U16087 (N_16087,N_15908,N_15909);
nor U16088 (N_16088,N_15860,N_15842);
and U16089 (N_16089,N_15961,N_15981);
or U16090 (N_16090,N_15988,N_15949);
xor U16091 (N_16091,N_15936,N_15818);
xnor U16092 (N_16092,N_15940,N_15911);
xor U16093 (N_16093,N_15829,N_15950);
xor U16094 (N_16094,N_15906,N_15958);
and U16095 (N_16095,N_15931,N_15986);
and U16096 (N_16096,N_15868,N_15999);
nand U16097 (N_16097,N_15882,N_15811);
or U16098 (N_16098,N_15935,N_15805);
nand U16099 (N_16099,N_15939,N_15995);
and U16100 (N_16100,N_15912,N_15965);
or U16101 (N_16101,N_15822,N_15930);
and U16102 (N_16102,N_15911,N_15816);
or U16103 (N_16103,N_15843,N_15986);
nor U16104 (N_16104,N_15803,N_15833);
or U16105 (N_16105,N_15961,N_15861);
nand U16106 (N_16106,N_15995,N_15869);
nor U16107 (N_16107,N_15888,N_15808);
xnor U16108 (N_16108,N_15832,N_15952);
nor U16109 (N_16109,N_15958,N_15864);
or U16110 (N_16110,N_15913,N_15948);
nor U16111 (N_16111,N_15849,N_15951);
nor U16112 (N_16112,N_15875,N_15828);
xor U16113 (N_16113,N_15935,N_15802);
and U16114 (N_16114,N_15973,N_15854);
xor U16115 (N_16115,N_15898,N_15947);
nor U16116 (N_16116,N_15822,N_15811);
nand U16117 (N_16117,N_15991,N_15982);
xnor U16118 (N_16118,N_15951,N_15897);
nor U16119 (N_16119,N_15975,N_15995);
xor U16120 (N_16120,N_15838,N_15873);
and U16121 (N_16121,N_15856,N_15834);
xnor U16122 (N_16122,N_15890,N_15902);
and U16123 (N_16123,N_15956,N_15885);
nor U16124 (N_16124,N_15836,N_15952);
nand U16125 (N_16125,N_15984,N_15965);
xor U16126 (N_16126,N_15941,N_15972);
nor U16127 (N_16127,N_15923,N_15944);
nor U16128 (N_16128,N_15869,N_15824);
or U16129 (N_16129,N_15919,N_15947);
nand U16130 (N_16130,N_15815,N_15999);
or U16131 (N_16131,N_15969,N_15925);
nor U16132 (N_16132,N_15831,N_15898);
xor U16133 (N_16133,N_15930,N_15940);
nand U16134 (N_16134,N_15882,N_15871);
nor U16135 (N_16135,N_15915,N_15817);
or U16136 (N_16136,N_15806,N_15811);
or U16137 (N_16137,N_15806,N_15821);
xor U16138 (N_16138,N_15989,N_15857);
or U16139 (N_16139,N_15901,N_15992);
nand U16140 (N_16140,N_15813,N_15915);
or U16141 (N_16141,N_15929,N_15883);
nand U16142 (N_16142,N_15997,N_15928);
nand U16143 (N_16143,N_15822,N_15953);
and U16144 (N_16144,N_15803,N_15917);
xor U16145 (N_16145,N_15823,N_15924);
xnor U16146 (N_16146,N_15918,N_15996);
xor U16147 (N_16147,N_15941,N_15977);
xor U16148 (N_16148,N_15920,N_15993);
xnor U16149 (N_16149,N_15815,N_15940);
nand U16150 (N_16150,N_15890,N_15861);
nor U16151 (N_16151,N_15803,N_15938);
or U16152 (N_16152,N_15952,N_15932);
nand U16153 (N_16153,N_15874,N_15990);
xor U16154 (N_16154,N_15816,N_15958);
nor U16155 (N_16155,N_15920,N_15894);
nand U16156 (N_16156,N_15973,N_15958);
nor U16157 (N_16157,N_15800,N_15894);
nor U16158 (N_16158,N_15948,N_15939);
nand U16159 (N_16159,N_15970,N_15909);
or U16160 (N_16160,N_15902,N_15842);
or U16161 (N_16161,N_15965,N_15808);
xnor U16162 (N_16162,N_15872,N_15916);
nand U16163 (N_16163,N_15864,N_15871);
xnor U16164 (N_16164,N_15831,N_15877);
nand U16165 (N_16165,N_15901,N_15974);
and U16166 (N_16166,N_15904,N_15824);
nor U16167 (N_16167,N_15970,N_15978);
nand U16168 (N_16168,N_15858,N_15954);
or U16169 (N_16169,N_15856,N_15987);
nand U16170 (N_16170,N_15876,N_15860);
xnor U16171 (N_16171,N_15894,N_15985);
nor U16172 (N_16172,N_15823,N_15990);
nor U16173 (N_16173,N_15881,N_15812);
or U16174 (N_16174,N_15908,N_15992);
or U16175 (N_16175,N_15962,N_15866);
or U16176 (N_16176,N_15891,N_15952);
nor U16177 (N_16177,N_15821,N_15956);
nor U16178 (N_16178,N_15805,N_15966);
or U16179 (N_16179,N_15813,N_15996);
nor U16180 (N_16180,N_15882,N_15830);
or U16181 (N_16181,N_15851,N_15803);
nand U16182 (N_16182,N_15895,N_15887);
nor U16183 (N_16183,N_15817,N_15966);
nand U16184 (N_16184,N_15997,N_15811);
xor U16185 (N_16185,N_15823,N_15827);
nor U16186 (N_16186,N_15802,N_15897);
xor U16187 (N_16187,N_15936,N_15904);
or U16188 (N_16188,N_15952,N_15897);
and U16189 (N_16189,N_15817,N_15954);
nand U16190 (N_16190,N_15849,N_15939);
or U16191 (N_16191,N_15920,N_15863);
nor U16192 (N_16192,N_15902,N_15824);
or U16193 (N_16193,N_15975,N_15981);
and U16194 (N_16194,N_15984,N_15859);
and U16195 (N_16195,N_15935,N_15890);
or U16196 (N_16196,N_15889,N_15918);
xnor U16197 (N_16197,N_15943,N_15843);
and U16198 (N_16198,N_15823,N_15844);
or U16199 (N_16199,N_15816,N_15823);
nor U16200 (N_16200,N_16000,N_16163);
and U16201 (N_16201,N_16020,N_16010);
nor U16202 (N_16202,N_16196,N_16148);
xnor U16203 (N_16203,N_16158,N_16178);
xor U16204 (N_16204,N_16060,N_16189);
nor U16205 (N_16205,N_16066,N_16127);
xnor U16206 (N_16206,N_16011,N_16167);
or U16207 (N_16207,N_16159,N_16099);
nor U16208 (N_16208,N_16086,N_16126);
xor U16209 (N_16209,N_16129,N_16119);
nand U16210 (N_16210,N_16036,N_16078);
and U16211 (N_16211,N_16077,N_16121);
nand U16212 (N_16212,N_16063,N_16059);
or U16213 (N_16213,N_16035,N_16191);
xor U16214 (N_16214,N_16058,N_16161);
or U16215 (N_16215,N_16007,N_16037);
and U16216 (N_16216,N_16061,N_16101);
or U16217 (N_16217,N_16019,N_16053);
or U16218 (N_16218,N_16096,N_16149);
or U16219 (N_16219,N_16081,N_16073);
xor U16220 (N_16220,N_16155,N_16054);
nor U16221 (N_16221,N_16120,N_16156);
nor U16222 (N_16222,N_16193,N_16082);
and U16223 (N_16223,N_16122,N_16188);
nor U16224 (N_16224,N_16017,N_16141);
and U16225 (N_16225,N_16170,N_16046);
or U16226 (N_16226,N_16041,N_16175);
nand U16227 (N_16227,N_16144,N_16045);
or U16228 (N_16228,N_16065,N_16027);
nand U16229 (N_16229,N_16110,N_16147);
nand U16230 (N_16230,N_16113,N_16165);
xnor U16231 (N_16231,N_16042,N_16090);
nand U16232 (N_16232,N_16047,N_16079);
or U16233 (N_16233,N_16140,N_16021);
and U16234 (N_16234,N_16104,N_16107);
nand U16235 (N_16235,N_16176,N_16106);
or U16236 (N_16236,N_16084,N_16003);
nand U16237 (N_16237,N_16118,N_16192);
or U16238 (N_16238,N_16044,N_16013);
or U16239 (N_16239,N_16025,N_16151);
or U16240 (N_16240,N_16031,N_16116);
or U16241 (N_16241,N_16092,N_16069);
nor U16242 (N_16242,N_16185,N_16172);
or U16243 (N_16243,N_16015,N_16135);
nand U16244 (N_16244,N_16049,N_16023);
and U16245 (N_16245,N_16105,N_16150);
nand U16246 (N_16246,N_16139,N_16102);
nand U16247 (N_16247,N_16186,N_16071);
xnor U16248 (N_16248,N_16074,N_16112);
or U16249 (N_16249,N_16085,N_16095);
nor U16250 (N_16250,N_16179,N_16199);
nand U16251 (N_16251,N_16157,N_16062);
and U16252 (N_16252,N_16076,N_16169);
nor U16253 (N_16253,N_16087,N_16108);
or U16254 (N_16254,N_16032,N_16184);
or U16255 (N_16255,N_16088,N_16051);
and U16256 (N_16256,N_16130,N_16030);
nor U16257 (N_16257,N_16123,N_16190);
and U16258 (N_16258,N_16195,N_16162);
xnor U16259 (N_16259,N_16018,N_16138);
and U16260 (N_16260,N_16136,N_16146);
and U16261 (N_16261,N_16057,N_16083);
and U16262 (N_16262,N_16055,N_16145);
xnor U16263 (N_16263,N_16103,N_16029);
nand U16264 (N_16264,N_16174,N_16026);
or U16265 (N_16265,N_16114,N_16001);
or U16266 (N_16266,N_16133,N_16160);
xor U16267 (N_16267,N_16072,N_16153);
nor U16268 (N_16268,N_16094,N_16142);
nor U16269 (N_16269,N_16016,N_16152);
xnor U16270 (N_16270,N_16173,N_16177);
or U16271 (N_16271,N_16034,N_16028);
and U16272 (N_16272,N_16012,N_16002);
nor U16273 (N_16273,N_16194,N_16124);
xor U16274 (N_16274,N_16131,N_16008);
or U16275 (N_16275,N_16070,N_16009);
and U16276 (N_16276,N_16006,N_16109);
nand U16277 (N_16277,N_16068,N_16143);
nor U16278 (N_16278,N_16033,N_16180);
and U16279 (N_16279,N_16154,N_16004);
or U16280 (N_16280,N_16093,N_16091);
nand U16281 (N_16281,N_16022,N_16168);
and U16282 (N_16282,N_16038,N_16098);
or U16283 (N_16283,N_16097,N_16164);
nand U16284 (N_16284,N_16171,N_16183);
nand U16285 (N_16285,N_16080,N_16117);
xor U16286 (N_16286,N_16043,N_16187);
xor U16287 (N_16287,N_16181,N_16040);
or U16288 (N_16288,N_16100,N_16197);
and U16289 (N_16289,N_16115,N_16052);
xnor U16290 (N_16290,N_16128,N_16048);
nor U16291 (N_16291,N_16198,N_16039);
or U16292 (N_16292,N_16134,N_16056);
and U16293 (N_16293,N_16064,N_16132);
xnor U16294 (N_16294,N_16050,N_16111);
or U16295 (N_16295,N_16075,N_16024);
nor U16296 (N_16296,N_16089,N_16125);
and U16297 (N_16297,N_16166,N_16005);
nor U16298 (N_16298,N_16067,N_16014);
and U16299 (N_16299,N_16182,N_16137);
xnor U16300 (N_16300,N_16082,N_16187);
nand U16301 (N_16301,N_16172,N_16005);
nor U16302 (N_16302,N_16104,N_16019);
nor U16303 (N_16303,N_16029,N_16055);
or U16304 (N_16304,N_16186,N_16036);
nand U16305 (N_16305,N_16066,N_16076);
or U16306 (N_16306,N_16117,N_16152);
nand U16307 (N_16307,N_16029,N_16146);
nand U16308 (N_16308,N_16019,N_16027);
nand U16309 (N_16309,N_16003,N_16087);
nor U16310 (N_16310,N_16192,N_16006);
and U16311 (N_16311,N_16051,N_16037);
nor U16312 (N_16312,N_16157,N_16146);
nand U16313 (N_16313,N_16151,N_16198);
xor U16314 (N_16314,N_16072,N_16040);
and U16315 (N_16315,N_16031,N_16181);
and U16316 (N_16316,N_16035,N_16190);
xnor U16317 (N_16317,N_16185,N_16186);
nand U16318 (N_16318,N_16185,N_16190);
and U16319 (N_16319,N_16115,N_16137);
nand U16320 (N_16320,N_16009,N_16136);
xnor U16321 (N_16321,N_16081,N_16126);
and U16322 (N_16322,N_16020,N_16052);
or U16323 (N_16323,N_16004,N_16103);
xnor U16324 (N_16324,N_16183,N_16068);
nand U16325 (N_16325,N_16005,N_16073);
nand U16326 (N_16326,N_16110,N_16028);
xor U16327 (N_16327,N_16101,N_16185);
xnor U16328 (N_16328,N_16054,N_16096);
nand U16329 (N_16329,N_16033,N_16168);
xnor U16330 (N_16330,N_16132,N_16153);
or U16331 (N_16331,N_16157,N_16053);
nand U16332 (N_16332,N_16198,N_16123);
or U16333 (N_16333,N_16169,N_16022);
xnor U16334 (N_16334,N_16022,N_16134);
nand U16335 (N_16335,N_16005,N_16082);
nor U16336 (N_16336,N_16030,N_16095);
xnor U16337 (N_16337,N_16084,N_16172);
xnor U16338 (N_16338,N_16041,N_16164);
nand U16339 (N_16339,N_16005,N_16145);
nand U16340 (N_16340,N_16002,N_16129);
nor U16341 (N_16341,N_16020,N_16163);
and U16342 (N_16342,N_16107,N_16110);
and U16343 (N_16343,N_16020,N_16015);
nor U16344 (N_16344,N_16120,N_16077);
and U16345 (N_16345,N_16020,N_16036);
or U16346 (N_16346,N_16165,N_16173);
nand U16347 (N_16347,N_16001,N_16067);
nand U16348 (N_16348,N_16106,N_16025);
nor U16349 (N_16349,N_16055,N_16166);
and U16350 (N_16350,N_16086,N_16037);
xor U16351 (N_16351,N_16135,N_16060);
nand U16352 (N_16352,N_16088,N_16122);
and U16353 (N_16353,N_16181,N_16032);
xor U16354 (N_16354,N_16179,N_16084);
or U16355 (N_16355,N_16098,N_16099);
nand U16356 (N_16356,N_16117,N_16082);
or U16357 (N_16357,N_16019,N_16046);
or U16358 (N_16358,N_16132,N_16158);
or U16359 (N_16359,N_16049,N_16143);
nor U16360 (N_16360,N_16054,N_16108);
nand U16361 (N_16361,N_16102,N_16199);
nand U16362 (N_16362,N_16197,N_16167);
nor U16363 (N_16363,N_16101,N_16010);
nor U16364 (N_16364,N_16143,N_16054);
and U16365 (N_16365,N_16075,N_16034);
xor U16366 (N_16366,N_16189,N_16038);
or U16367 (N_16367,N_16125,N_16127);
xor U16368 (N_16368,N_16188,N_16175);
xnor U16369 (N_16369,N_16078,N_16157);
nor U16370 (N_16370,N_16016,N_16192);
nor U16371 (N_16371,N_16109,N_16151);
nand U16372 (N_16372,N_16162,N_16171);
nand U16373 (N_16373,N_16187,N_16168);
xnor U16374 (N_16374,N_16024,N_16097);
xor U16375 (N_16375,N_16053,N_16016);
xor U16376 (N_16376,N_16149,N_16044);
and U16377 (N_16377,N_16060,N_16104);
nor U16378 (N_16378,N_16062,N_16053);
xnor U16379 (N_16379,N_16111,N_16173);
xnor U16380 (N_16380,N_16066,N_16064);
nor U16381 (N_16381,N_16072,N_16116);
xor U16382 (N_16382,N_16097,N_16196);
xor U16383 (N_16383,N_16020,N_16123);
and U16384 (N_16384,N_16097,N_16117);
nand U16385 (N_16385,N_16010,N_16177);
nor U16386 (N_16386,N_16126,N_16145);
and U16387 (N_16387,N_16174,N_16018);
nand U16388 (N_16388,N_16142,N_16109);
xnor U16389 (N_16389,N_16192,N_16050);
nand U16390 (N_16390,N_16179,N_16072);
or U16391 (N_16391,N_16154,N_16176);
and U16392 (N_16392,N_16021,N_16060);
nand U16393 (N_16393,N_16072,N_16096);
nand U16394 (N_16394,N_16172,N_16153);
or U16395 (N_16395,N_16199,N_16049);
nor U16396 (N_16396,N_16109,N_16135);
and U16397 (N_16397,N_16030,N_16045);
xor U16398 (N_16398,N_16185,N_16070);
or U16399 (N_16399,N_16004,N_16158);
nand U16400 (N_16400,N_16283,N_16294);
or U16401 (N_16401,N_16254,N_16384);
or U16402 (N_16402,N_16220,N_16211);
xnor U16403 (N_16403,N_16341,N_16206);
xor U16404 (N_16404,N_16389,N_16263);
and U16405 (N_16405,N_16301,N_16380);
or U16406 (N_16406,N_16370,N_16312);
nor U16407 (N_16407,N_16371,N_16266);
nor U16408 (N_16408,N_16375,N_16264);
or U16409 (N_16409,N_16276,N_16340);
xnor U16410 (N_16410,N_16269,N_16396);
nor U16411 (N_16411,N_16212,N_16320);
and U16412 (N_16412,N_16324,N_16280);
nor U16413 (N_16413,N_16267,N_16291);
or U16414 (N_16414,N_16397,N_16367);
or U16415 (N_16415,N_16318,N_16325);
or U16416 (N_16416,N_16272,N_16222);
xnor U16417 (N_16417,N_16306,N_16339);
and U16418 (N_16418,N_16378,N_16246);
nor U16419 (N_16419,N_16303,N_16233);
xnor U16420 (N_16420,N_16241,N_16334);
nand U16421 (N_16421,N_16225,N_16281);
nor U16422 (N_16422,N_16207,N_16361);
nor U16423 (N_16423,N_16293,N_16289);
and U16424 (N_16424,N_16232,N_16290);
nor U16425 (N_16425,N_16231,N_16250);
or U16426 (N_16426,N_16393,N_16376);
nand U16427 (N_16427,N_16282,N_16201);
xor U16428 (N_16428,N_16348,N_16261);
or U16429 (N_16429,N_16239,N_16387);
or U16430 (N_16430,N_16299,N_16309);
nor U16431 (N_16431,N_16379,N_16385);
and U16432 (N_16432,N_16373,N_16286);
or U16433 (N_16433,N_16360,N_16242);
nor U16434 (N_16434,N_16328,N_16288);
nor U16435 (N_16435,N_16221,N_16359);
nor U16436 (N_16436,N_16357,N_16323);
nor U16437 (N_16437,N_16308,N_16298);
nor U16438 (N_16438,N_16236,N_16381);
and U16439 (N_16439,N_16287,N_16268);
and U16440 (N_16440,N_16321,N_16248);
xnor U16441 (N_16441,N_16363,N_16330);
or U16442 (N_16442,N_16329,N_16346);
nand U16443 (N_16443,N_16237,N_16395);
or U16444 (N_16444,N_16202,N_16251);
nor U16445 (N_16445,N_16398,N_16297);
xor U16446 (N_16446,N_16349,N_16295);
xnor U16447 (N_16447,N_16304,N_16392);
nor U16448 (N_16448,N_16256,N_16217);
and U16449 (N_16449,N_16244,N_16333);
nor U16450 (N_16450,N_16240,N_16391);
or U16451 (N_16451,N_16355,N_16270);
xor U16452 (N_16452,N_16238,N_16352);
nand U16453 (N_16453,N_16353,N_16316);
and U16454 (N_16454,N_16215,N_16257);
nor U16455 (N_16455,N_16262,N_16399);
and U16456 (N_16456,N_16394,N_16300);
xor U16457 (N_16457,N_16275,N_16344);
nand U16458 (N_16458,N_16372,N_16203);
and U16459 (N_16459,N_16214,N_16307);
nor U16460 (N_16460,N_16342,N_16235);
or U16461 (N_16461,N_16382,N_16277);
nand U16462 (N_16462,N_16317,N_16362);
nand U16463 (N_16463,N_16279,N_16337);
and U16464 (N_16464,N_16311,N_16219);
or U16465 (N_16465,N_16234,N_16296);
xnor U16466 (N_16466,N_16292,N_16358);
nand U16467 (N_16467,N_16204,N_16265);
nand U16468 (N_16468,N_16255,N_16227);
nor U16469 (N_16469,N_16345,N_16216);
xor U16470 (N_16470,N_16210,N_16327);
and U16471 (N_16471,N_16253,N_16224);
or U16472 (N_16472,N_16315,N_16274);
or U16473 (N_16473,N_16364,N_16271);
or U16474 (N_16474,N_16249,N_16336);
nor U16475 (N_16475,N_16377,N_16205);
or U16476 (N_16476,N_16285,N_16213);
nand U16477 (N_16477,N_16314,N_16259);
or U16478 (N_16478,N_16369,N_16273);
nand U16479 (N_16479,N_16335,N_16356);
nor U16480 (N_16480,N_16319,N_16351);
and U16481 (N_16481,N_16258,N_16247);
xor U16482 (N_16482,N_16305,N_16228);
or U16483 (N_16483,N_16365,N_16218);
nor U16484 (N_16484,N_16322,N_16388);
xnor U16485 (N_16485,N_16326,N_16374);
or U16486 (N_16486,N_16383,N_16260);
xnor U16487 (N_16487,N_16284,N_16332);
xnor U16488 (N_16488,N_16338,N_16331);
or U16489 (N_16489,N_16310,N_16200);
nor U16490 (N_16490,N_16390,N_16368);
nor U16491 (N_16491,N_16354,N_16208);
or U16492 (N_16492,N_16245,N_16350);
xnor U16493 (N_16493,N_16343,N_16226);
or U16494 (N_16494,N_16302,N_16230);
nor U16495 (N_16495,N_16366,N_16313);
or U16496 (N_16496,N_16229,N_16347);
and U16497 (N_16497,N_16278,N_16209);
nor U16498 (N_16498,N_16243,N_16252);
and U16499 (N_16499,N_16223,N_16386);
xnor U16500 (N_16500,N_16210,N_16203);
nor U16501 (N_16501,N_16263,N_16394);
nor U16502 (N_16502,N_16387,N_16231);
and U16503 (N_16503,N_16252,N_16338);
xor U16504 (N_16504,N_16346,N_16298);
nor U16505 (N_16505,N_16227,N_16252);
and U16506 (N_16506,N_16333,N_16252);
xnor U16507 (N_16507,N_16354,N_16284);
xnor U16508 (N_16508,N_16205,N_16211);
and U16509 (N_16509,N_16398,N_16289);
nand U16510 (N_16510,N_16356,N_16391);
nand U16511 (N_16511,N_16368,N_16204);
and U16512 (N_16512,N_16308,N_16367);
nor U16513 (N_16513,N_16372,N_16314);
nor U16514 (N_16514,N_16317,N_16212);
nand U16515 (N_16515,N_16335,N_16314);
and U16516 (N_16516,N_16315,N_16227);
and U16517 (N_16517,N_16316,N_16291);
or U16518 (N_16518,N_16349,N_16231);
and U16519 (N_16519,N_16294,N_16278);
nand U16520 (N_16520,N_16238,N_16344);
nand U16521 (N_16521,N_16203,N_16226);
or U16522 (N_16522,N_16286,N_16309);
nand U16523 (N_16523,N_16387,N_16274);
or U16524 (N_16524,N_16299,N_16352);
and U16525 (N_16525,N_16356,N_16333);
nand U16526 (N_16526,N_16310,N_16352);
and U16527 (N_16527,N_16278,N_16279);
nand U16528 (N_16528,N_16216,N_16200);
or U16529 (N_16529,N_16215,N_16328);
or U16530 (N_16530,N_16278,N_16260);
nor U16531 (N_16531,N_16251,N_16252);
xor U16532 (N_16532,N_16369,N_16243);
xnor U16533 (N_16533,N_16245,N_16326);
nand U16534 (N_16534,N_16224,N_16362);
nand U16535 (N_16535,N_16366,N_16354);
and U16536 (N_16536,N_16356,N_16365);
nor U16537 (N_16537,N_16222,N_16380);
nand U16538 (N_16538,N_16362,N_16233);
xnor U16539 (N_16539,N_16247,N_16261);
xor U16540 (N_16540,N_16295,N_16264);
nor U16541 (N_16541,N_16370,N_16216);
xnor U16542 (N_16542,N_16348,N_16270);
or U16543 (N_16543,N_16396,N_16363);
and U16544 (N_16544,N_16202,N_16321);
nor U16545 (N_16545,N_16296,N_16317);
and U16546 (N_16546,N_16262,N_16355);
nor U16547 (N_16547,N_16377,N_16324);
xnor U16548 (N_16548,N_16239,N_16319);
nand U16549 (N_16549,N_16289,N_16382);
nand U16550 (N_16550,N_16279,N_16375);
nor U16551 (N_16551,N_16240,N_16352);
nand U16552 (N_16552,N_16329,N_16208);
or U16553 (N_16553,N_16203,N_16201);
xnor U16554 (N_16554,N_16303,N_16273);
or U16555 (N_16555,N_16232,N_16331);
nor U16556 (N_16556,N_16256,N_16323);
xnor U16557 (N_16557,N_16340,N_16347);
or U16558 (N_16558,N_16373,N_16321);
xor U16559 (N_16559,N_16274,N_16370);
nor U16560 (N_16560,N_16231,N_16280);
or U16561 (N_16561,N_16289,N_16318);
nor U16562 (N_16562,N_16349,N_16398);
xnor U16563 (N_16563,N_16276,N_16345);
nand U16564 (N_16564,N_16272,N_16240);
xor U16565 (N_16565,N_16298,N_16368);
xnor U16566 (N_16566,N_16372,N_16336);
xnor U16567 (N_16567,N_16337,N_16223);
nor U16568 (N_16568,N_16305,N_16236);
and U16569 (N_16569,N_16274,N_16259);
xor U16570 (N_16570,N_16212,N_16278);
and U16571 (N_16571,N_16388,N_16373);
nand U16572 (N_16572,N_16339,N_16275);
nor U16573 (N_16573,N_16308,N_16225);
or U16574 (N_16574,N_16285,N_16359);
nor U16575 (N_16575,N_16266,N_16229);
or U16576 (N_16576,N_16293,N_16230);
and U16577 (N_16577,N_16253,N_16334);
nor U16578 (N_16578,N_16329,N_16278);
nor U16579 (N_16579,N_16230,N_16271);
xor U16580 (N_16580,N_16263,N_16223);
nor U16581 (N_16581,N_16393,N_16334);
and U16582 (N_16582,N_16391,N_16231);
nor U16583 (N_16583,N_16373,N_16355);
or U16584 (N_16584,N_16386,N_16377);
nor U16585 (N_16585,N_16286,N_16360);
xnor U16586 (N_16586,N_16364,N_16300);
or U16587 (N_16587,N_16279,N_16287);
and U16588 (N_16588,N_16367,N_16277);
and U16589 (N_16589,N_16316,N_16377);
nor U16590 (N_16590,N_16375,N_16298);
nand U16591 (N_16591,N_16239,N_16263);
xor U16592 (N_16592,N_16296,N_16274);
nand U16593 (N_16593,N_16342,N_16269);
or U16594 (N_16594,N_16347,N_16376);
or U16595 (N_16595,N_16375,N_16310);
xnor U16596 (N_16596,N_16328,N_16270);
nand U16597 (N_16597,N_16306,N_16256);
nand U16598 (N_16598,N_16274,N_16339);
and U16599 (N_16599,N_16323,N_16366);
xnor U16600 (N_16600,N_16549,N_16421);
or U16601 (N_16601,N_16414,N_16596);
nor U16602 (N_16602,N_16597,N_16553);
and U16603 (N_16603,N_16494,N_16554);
xnor U16604 (N_16604,N_16493,N_16537);
nor U16605 (N_16605,N_16566,N_16479);
nor U16606 (N_16606,N_16556,N_16503);
xnor U16607 (N_16607,N_16422,N_16403);
nor U16608 (N_16608,N_16518,N_16443);
and U16609 (N_16609,N_16569,N_16438);
and U16610 (N_16610,N_16533,N_16534);
and U16611 (N_16611,N_16436,N_16515);
xor U16612 (N_16612,N_16498,N_16577);
xnor U16613 (N_16613,N_16430,N_16473);
nand U16614 (N_16614,N_16568,N_16470);
xor U16615 (N_16615,N_16405,N_16586);
nor U16616 (N_16616,N_16578,N_16591);
nand U16617 (N_16617,N_16508,N_16565);
nand U16618 (N_16618,N_16447,N_16424);
or U16619 (N_16619,N_16485,N_16408);
xnor U16620 (N_16620,N_16450,N_16462);
nand U16621 (N_16621,N_16567,N_16589);
or U16622 (N_16622,N_16418,N_16522);
nand U16623 (N_16623,N_16541,N_16461);
nand U16624 (N_16624,N_16521,N_16448);
or U16625 (N_16625,N_16435,N_16574);
or U16626 (N_16626,N_16542,N_16579);
xnor U16627 (N_16627,N_16483,N_16445);
nand U16628 (N_16628,N_16573,N_16407);
xnor U16629 (N_16629,N_16571,N_16598);
and U16630 (N_16630,N_16490,N_16527);
xor U16631 (N_16631,N_16491,N_16559);
nor U16632 (N_16632,N_16416,N_16581);
xor U16633 (N_16633,N_16439,N_16444);
or U16634 (N_16634,N_16495,N_16463);
or U16635 (N_16635,N_16562,N_16530);
nor U16636 (N_16636,N_16520,N_16545);
nand U16637 (N_16637,N_16476,N_16497);
xnor U16638 (N_16638,N_16452,N_16551);
xor U16639 (N_16639,N_16441,N_16509);
or U16640 (N_16640,N_16546,N_16477);
nand U16641 (N_16641,N_16594,N_16505);
nand U16642 (N_16642,N_16484,N_16457);
xnor U16643 (N_16643,N_16440,N_16555);
and U16644 (N_16644,N_16507,N_16442);
nor U16645 (N_16645,N_16529,N_16426);
or U16646 (N_16646,N_16464,N_16592);
and U16647 (N_16647,N_16502,N_16486);
xnor U16648 (N_16648,N_16510,N_16532);
or U16649 (N_16649,N_16412,N_16593);
or U16650 (N_16650,N_16504,N_16467);
xor U16651 (N_16651,N_16588,N_16404);
nand U16652 (N_16652,N_16539,N_16482);
nor U16653 (N_16653,N_16516,N_16411);
nor U16654 (N_16654,N_16506,N_16514);
or U16655 (N_16655,N_16512,N_16531);
nor U16656 (N_16656,N_16474,N_16433);
nor U16657 (N_16657,N_16472,N_16400);
or U16658 (N_16658,N_16456,N_16459);
nor U16659 (N_16659,N_16535,N_16402);
and U16660 (N_16660,N_16536,N_16423);
nand U16661 (N_16661,N_16420,N_16587);
xnor U16662 (N_16662,N_16437,N_16468);
nand U16663 (N_16663,N_16451,N_16487);
nand U16664 (N_16664,N_16519,N_16469);
and U16665 (N_16665,N_16471,N_16454);
or U16666 (N_16666,N_16453,N_16434);
or U16667 (N_16667,N_16480,N_16413);
xor U16668 (N_16668,N_16466,N_16460);
and U16669 (N_16669,N_16524,N_16401);
nand U16670 (N_16670,N_16410,N_16557);
nor U16671 (N_16671,N_16580,N_16560);
xor U16672 (N_16672,N_16540,N_16538);
nor U16673 (N_16673,N_16558,N_16432);
xnor U16674 (N_16674,N_16547,N_16419);
or U16675 (N_16675,N_16496,N_16511);
xnor U16676 (N_16676,N_16582,N_16475);
and U16677 (N_16677,N_16492,N_16544);
and U16678 (N_16678,N_16488,N_16425);
and U16679 (N_16679,N_16543,N_16528);
xor U16680 (N_16680,N_16449,N_16564);
and U16681 (N_16681,N_16595,N_16526);
or U16682 (N_16682,N_16409,N_16429);
or U16683 (N_16683,N_16458,N_16513);
xor U16684 (N_16684,N_16575,N_16415);
or U16685 (N_16685,N_16561,N_16499);
or U16686 (N_16686,N_16550,N_16406);
or U16687 (N_16687,N_16599,N_16585);
nor U16688 (N_16688,N_16427,N_16455);
nand U16689 (N_16689,N_16501,N_16563);
or U16690 (N_16690,N_16548,N_16590);
nand U16691 (N_16691,N_16500,N_16465);
and U16692 (N_16692,N_16552,N_16570);
xor U16693 (N_16693,N_16517,N_16576);
xor U16694 (N_16694,N_16583,N_16584);
nor U16695 (N_16695,N_16525,N_16523);
xor U16696 (N_16696,N_16446,N_16431);
and U16697 (N_16697,N_16572,N_16481);
and U16698 (N_16698,N_16428,N_16478);
or U16699 (N_16699,N_16489,N_16417);
or U16700 (N_16700,N_16537,N_16487);
and U16701 (N_16701,N_16471,N_16588);
nor U16702 (N_16702,N_16442,N_16500);
and U16703 (N_16703,N_16538,N_16452);
or U16704 (N_16704,N_16507,N_16416);
or U16705 (N_16705,N_16546,N_16411);
or U16706 (N_16706,N_16548,N_16514);
and U16707 (N_16707,N_16516,N_16455);
nor U16708 (N_16708,N_16573,N_16524);
or U16709 (N_16709,N_16560,N_16566);
and U16710 (N_16710,N_16454,N_16450);
nand U16711 (N_16711,N_16516,N_16521);
and U16712 (N_16712,N_16438,N_16571);
or U16713 (N_16713,N_16452,N_16585);
nor U16714 (N_16714,N_16499,N_16469);
nand U16715 (N_16715,N_16489,N_16564);
and U16716 (N_16716,N_16445,N_16536);
nor U16717 (N_16717,N_16587,N_16470);
and U16718 (N_16718,N_16490,N_16535);
nand U16719 (N_16719,N_16415,N_16446);
nor U16720 (N_16720,N_16538,N_16518);
nand U16721 (N_16721,N_16596,N_16532);
or U16722 (N_16722,N_16459,N_16424);
nor U16723 (N_16723,N_16570,N_16536);
nor U16724 (N_16724,N_16428,N_16429);
nor U16725 (N_16725,N_16499,N_16403);
nand U16726 (N_16726,N_16425,N_16522);
or U16727 (N_16727,N_16401,N_16516);
nor U16728 (N_16728,N_16453,N_16432);
nor U16729 (N_16729,N_16488,N_16523);
or U16730 (N_16730,N_16481,N_16487);
nand U16731 (N_16731,N_16582,N_16411);
and U16732 (N_16732,N_16561,N_16582);
xnor U16733 (N_16733,N_16400,N_16423);
nor U16734 (N_16734,N_16497,N_16536);
and U16735 (N_16735,N_16417,N_16484);
xor U16736 (N_16736,N_16483,N_16593);
nand U16737 (N_16737,N_16564,N_16512);
xor U16738 (N_16738,N_16438,N_16488);
or U16739 (N_16739,N_16496,N_16586);
nand U16740 (N_16740,N_16459,N_16486);
and U16741 (N_16741,N_16580,N_16453);
nand U16742 (N_16742,N_16594,N_16481);
nand U16743 (N_16743,N_16531,N_16574);
nor U16744 (N_16744,N_16547,N_16504);
or U16745 (N_16745,N_16438,N_16492);
and U16746 (N_16746,N_16439,N_16537);
and U16747 (N_16747,N_16449,N_16557);
nand U16748 (N_16748,N_16453,N_16528);
or U16749 (N_16749,N_16430,N_16496);
nor U16750 (N_16750,N_16451,N_16501);
nand U16751 (N_16751,N_16573,N_16405);
xnor U16752 (N_16752,N_16423,N_16480);
or U16753 (N_16753,N_16580,N_16421);
xnor U16754 (N_16754,N_16405,N_16416);
and U16755 (N_16755,N_16537,N_16598);
nand U16756 (N_16756,N_16530,N_16505);
nand U16757 (N_16757,N_16500,N_16512);
nand U16758 (N_16758,N_16536,N_16567);
nand U16759 (N_16759,N_16541,N_16494);
or U16760 (N_16760,N_16453,N_16598);
xnor U16761 (N_16761,N_16525,N_16560);
and U16762 (N_16762,N_16548,N_16439);
or U16763 (N_16763,N_16453,N_16410);
xor U16764 (N_16764,N_16588,N_16563);
nand U16765 (N_16765,N_16417,N_16490);
nand U16766 (N_16766,N_16486,N_16415);
or U16767 (N_16767,N_16465,N_16479);
and U16768 (N_16768,N_16552,N_16595);
nand U16769 (N_16769,N_16405,N_16560);
or U16770 (N_16770,N_16566,N_16445);
or U16771 (N_16771,N_16566,N_16457);
or U16772 (N_16772,N_16518,N_16412);
or U16773 (N_16773,N_16474,N_16558);
or U16774 (N_16774,N_16502,N_16528);
nand U16775 (N_16775,N_16459,N_16505);
or U16776 (N_16776,N_16506,N_16445);
nand U16777 (N_16777,N_16556,N_16500);
nand U16778 (N_16778,N_16533,N_16453);
nor U16779 (N_16779,N_16538,N_16466);
xnor U16780 (N_16780,N_16505,N_16589);
or U16781 (N_16781,N_16530,N_16534);
and U16782 (N_16782,N_16526,N_16456);
nand U16783 (N_16783,N_16467,N_16577);
and U16784 (N_16784,N_16523,N_16505);
xor U16785 (N_16785,N_16416,N_16571);
nand U16786 (N_16786,N_16523,N_16554);
nor U16787 (N_16787,N_16478,N_16589);
nand U16788 (N_16788,N_16572,N_16571);
nand U16789 (N_16789,N_16489,N_16551);
or U16790 (N_16790,N_16489,N_16524);
and U16791 (N_16791,N_16523,N_16501);
nand U16792 (N_16792,N_16490,N_16426);
nor U16793 (N_16793,N_16436,N_16520);
nand U16794 (N_16794,N_16571,N_16504);
nor U16795 (N_16795,N_16533,N_16485);
nand U16796 (N_16796,N_16447,N_16513);
nor U16797 (N_16797,N_16552,N_16525);
or U16798 (N_16798,N_16568,N_16522);
nor U16799 (N_16799,N_16525,N_16405);
xor U16800 (N_16800,N_16602,N_16607);
xnor U16801 (N_16801,N_16730,N_16711);
or U16802 (N_16802,N_16798,N_16773);
nand U16803 (N_16803,N_16768,N_16791);
and U16804 (N_16804,N_16750,N_16685);
xor U16805 (N_16805,N_16705,N_16767);
or U16806 (N_16806,N_16635,N_16659);
nor U16807 (N_16807,N_16669,N_16657);
or U16808 (N_16808,N_16759,N_16620);
nor U16809 (N_16809,N_16727,N_16748);
xor U16810 (N_16810,N_16777,N_16679);
or U16811 (N_16811,N_16761,N_16682);
xnor U16812 (N_16812,N_16680,N_16681);
or U16813 (N_16813,N_16692,N_16612);
nor U16814 (N_16814,N_16751,N_16738);
xor U16815 (N_16815,N_16785,N_16674);
or U16816 (N_16816,N_16735,N_16799);
nand U16817 (N_16817,N_16671,N_16781);
nand U16818 (N_16818,N_16697,N_16629);
nand U16819 (N_16819,N_16639,N_16677);
or U16820 (N_16820,N_16691,N_16630);
xnor U16821 (N_16821,N_16733,N_16737);
and U16822 (N_16822,N_16728,N_16709);
nor U16823 (N_16823,N_16716,N_16690);
or U16824 (N_16824,N_16666,N_16661);
nand U16825 (N_16825,N_16600,N_16601);
nand U16826 (N_16826,N_16622,N_16615);
or U16827 (N_16827,N_16604,N_16694);
xor U16828 (N_16828,N_16747,N_16626);
nor U16829 (N_16829,N_16644,N_16775);
xnor U16830 (N_16830,N_16795,N_16744);
nor U16831 (N_16831,N_16676,N_16743);
nand U16832 (N_16832,N_16776,N_16634);
or U16833 (N_16833,N_16687,N_16723);
nand U16834 (N_16834,N_16782,N_16650);
nand U16835 (N_16835,N_16770,N_16632);
nor U16836 (N_16836,N_16715,N_16794);
or U16837 (N_16837,N_16792,N_16755);
or U16838 (N_16838,N_16712,N_16762);
nor U16839 (N_16839,N_16672,N_16609);
or U16840 (N_16840,N_16613,N_16667);
or U16841 (N_16841,N_16623,N_16724);
or U16842 (N_16842,N_16725,N_16624);
xnor U16843 (N_16843,N_16664,N_16718);
xor U16844 (N_16844,N_16670,N_16722);
nand U16845 (N_16845,N_16696,N_16706);
nand U16846 (N_16846,N_16760,N_16736);
xor U16847 (N_16847,N_16673,N_16688);
nand U16848 (N_16848,N_16766,N_16637);
and U16849 (N_16849,N_16686,N_16636);
nand U16850 (N_16850,N_16764,N_16643);
nand U16851 (N_16851,N_16614,N_16746);
xnor U16852 (N_16852,N_16753,N_16779);
xor U16853 (N_16853,N_16720,N_16771);
nand U16854 (N_16854,N_16787,N_16780);
nand U16855 (N_16855,N_16605,N_16645);
nand U16856 (N_16856,N_16678,N_16708);
or U16857 (N_16857,N_16606,N_16603);
or U16858 (N_16858,N_16660,N_16638);
and U16859 (N_16859,N_16749,N_16621);
and U16860 (N_16860,N_16665,N_16797);
nor U16861 (N_16861,N_16610,N_16689);
nand U16862 (N_16862,N_16658,N_16683);
or U16863 (N_16863,N_16729,N_16765);
and U16864 (N_16864,N_16662,N_16628);
and U16865 (N_16865,N_16653,N_16633);
nand U16866 (N_16866,N_16778,N_16789);
nand U16867 (N_16867,N_16611,N_16754);
nor U16868 (N_16868,N_16651,N_16702);
or U16869 (N_16869,N_16758,N_16756);
nand U16870 (N_16870,N_16793,N_16668);
nor U16871 (N_16871,N_16741,N_16700);
nor U16872 (N_16872,N_16769,N_16619);
nand U16873 (N_16873,N_16652,N_16675);
or U16874 (N_16874,N_16648,N_16790);
xor U16875 (N_16875,N_16788,N_16726);
nand U16876 (N_16876,N_16752,N_16663);
and U16877 (N_16877,N_16704,N_16647);
nand U16878 (N_16878,N_16701,N_16734);
xnor U16879 (N_16879,N_16745,N_16608);
nor U16880 (N_16880,N_16641,N_16693);
or U16881 (N_16881,N_16627,N_16721);
nand U16882 (N_16882,N_16640,N_16618);
nor U16883 (N_16883,N_16649,N_16786);
xnor U16884 (N_16884,N_16713,N_16784);
xor U16885 (N_16885,N_16631,N_16717);
and U16886 (N_16886,N_16783,N_16763);
nand U16887 (N_16887,N_16684,N_16654);
xnor U16888 (N_16888,N_16707,N_16757);
and U16889 (N_16889,N_16740,N_16796);
nor U16890 (N_16890,N_16739,N_16699);
and U16891 (N_16891,N_16695,N_16625);
and U16892 (N_16892,N_16719,N_16772);
nor U16893 (N_16893,N_16714,N_16774);
xor U16894 (N_16894,N_16742,N_16731);
and U16895 (N_16895,N_16642,N_16732);
nor U16896 (N_16896,N_16646,N_16698);
or U16897 (N_16897,N_16655,N_16616);
or U16898 (N_16898,N_16656,N_16703);
xor U16899 (N_16899,N_16710,N_16617);
xnor U16900 (N_16900,N_16685,N_16604);
and U16901 (N_16901,N_16667,N_16627);
xnor U16902 (N_16902,N_16774,N_16748);
nor U16903 (N_16903,N_16677,N_16787);
and U16904 (N_16904,N_16795,N_16747);
nand U16905 (N_16905,N_16674,N_16661);
or U16906 (N_16906,N_16768,N_16740);
and U16907 (N_16907,N_16663,N_16727);
or U16908 (N_16908,N_16703,N_16767);
and U16909 (N_16909,N_16694,N_16678);
or U16910 (N_16910,N_16671,N_16787);
nor U16911 (N_16911,N_16753,N_16784);
or U16912 (N_16912,N_16791,N_16661);
or U16913 (N_16913,N_16752,N_16609);
and U16914 (N_16914,N_16686,N_16661);
and U16915 (N_16915,N_16768,N_16688);
or U16916 (N_16916,N_16634,N_16726);
or U16917 (N_16917,N_16777,N_16640);
and U16918 (N_16918,N_16610,N_16703);
or U16919 (N_16919,N_16688,N_16700);
and U16920 (N_16920,N_16692,N_16690);
and U16921 (N_16921,N_16789,N_16797);
or U16922 (N_16922,N_16725,N_16656);
or U16923 (N_16923,N_16601,N_16751);
nand U16924 (N_16924,N_16612,N_16747);
xor U16925 (N_16925,N_16635,N_16716);
xnor U16926 (N_16926,N_16602,N_16650);
or U16927 (N_16927,N_16795,N_16646);
nand U16928 (N_16928,N_16684,N_16620);
nand U16929 (N_16929,N_16719,N_16624);
xnor U16930 (N_16930,N_16783,N_16669);
and U16931 (N_16931,N_16662,N_16733);
nand U16932 (N_16932,N_16697,N_16615);
xnor U16933 (N_16933,N_16734,N_16697);
xnor U16934 (N_16934,N_16683,N_16678);
xor U16935 (N_16935,N_16646,N_16729);
and U16936 (N_16936,N_16781,N_16603);
nand U16937 (N_16937,N_16753,N_16716);
and U16938 (N_16938,N_16718,N_16786);
and U16939 (N_16939,N_16795,N_16745);
nand U16940 (N_16940,N_16652,N_16678);
xor U16941 (N_16941,N_16790,N_16611);
and U16942 (N_16942,N_16656,N_16733);
nand U16943 (N_16943,N_16786,N_16739);
nor U16944 (N_16944,N_16659,N_16684);
or U16945 (N_16945,N_16716,N_16735);
xor U16946 (N_16946,N_16624,N_16699);
nor U16947 (N_16947,N_16770,N_16678);
nor U16948 (N_16948,N_16690,N_16741);
nor U16949 (N_16949,N_16642,N_16679);
and U16950 (N_16950,N_16626,N_16648);
xnor U16951 (N_16951,N_16757,N_16657);
nor U16952 (N_16952,N_16759,N_16799);
xnor U16953 (N_16953,N_16653,N_16701);
and U16954 (N_16954,N_16643,N_16662);
nor U16955 (N_16955,N_16681,N_16637);
and U16956 (N_16956,N_16624,N_16729);
xnor U16957 (N_16957,N_16638,N_16735);
nor U16958 (N_16958,N_16678,N_16778);
xor U16959 (N_16959,N_16606,N_16741);
xnor U16960 (N_16960,N_16672,N_16665);
xor U16961 (N_16961,N_16628,N_16636);
nor U16962 (N_16962,N_16674,N_16679);
and U16963 (N_16963,N_16735,N_16625);
xnor U16964 (N_16964,N_16787,N_16773);
nand U16965 (N_16965,N_16631,N_16795);
and U16966 (N_16966,N_16649,N_16690);
or U16967 (N_16967,N_16648,N_16761);
nand U16968 (N_16968,N_16725,N_16685);
nand U16969 (N_16969,N_16664,N_16612);
or U16970 (N_16970,N_16769,N_16611);
nand U16971 (N_16971,N_16696,N_16788);
or U16972 (N_16972,N_16617,N_16739);
or U16973 (N_16973,N_16649,N_16727);
or U16974 (N_16974,N_16639,N_16651);
or U16975 (N_16975,N_16757,N_16631);
nor U16976 (N_16976,N_16658,N_16736);
xor U16977 (N_16977,N_16740,N_16639);
nor U16978 (N_16978,N_16647,N_16654);
nor U16979 (N_16979,N_16654,N_16662);
or U16980 (N_16980,N_16712,N_16755);
and U16981 (N_16981,N_16710,N_16767);
xnor U16982 (N_16982,N_16613,N_16796);
and U16983 (N_16983,N_16669,N_16653);
nand U16984 (N_16984,N_16663,N_16622);
and U16985 (N_16985,N_16681,N_16677);
nand U16986 (N_16986,N_16603,N_16704);
nand U16987 (N_16987,N_16726,N_16605);
nor U16988 (N_16988,N_16632,N_16789);
or U16989 (N_16989,N_16703,N_16734);
and U16990 (N_16990,N_16610,N_16765);
nand U16991 (N_16991,N_16746,N_16734);
nand U16992 (N_16992,N_16734,N_16720);
nand U16993 (N_16993,N_16721,N_16620);
nand U16994 (N_16994,N_16684,N_16672);
or U16995 (N_16995,N_16777,N_16697);
nor U16996 (N_16996,N_16728,N_16703);
xnor U16997 (N_16997,N_16675,N_16771);
or U16998 (N_16998,N_16699,N_16796);
nor U16999 (N_16999,N_16634,N_16649);
nor U17000 (N_17000,N_16988,N_16968);
nor U17001 (N_17001,N_16880,N_16923);
or U17002 (N_17002,N_16827,N_16935);
nand U17003 (N_17003,N_16895,N_16953);
nand U17004 (N_17004,N_16901,N_16841);
and U17005 (N_17005,N_16931,N_16810);
xor U17006 (N_17006,N_16892,N_16878);
xor U17007 (N_17007,N_16936,N_16884);
or U17008 (N_17008,N_16918,N_16964);
xor U17009 (N_17009,N_16991,N_16938);
or U17010 (N_17010,N_16856,N_16854);
xnor U17011 (N_17011,N_16825,N_16847);
xor U17012 (N_17012,N_16898,N_16849);
and U17013 (N_17013,N_16843,N_16829);
nand U17014 (N_17014,N_16870,N_16906);
or U17015 (N_17015,N_16925,N_16820);
and U17016 (N_17016,N_16881,N_16919);
or U17017 (N_17017,N_16816,N_16814);
and U17018 (N_17018,N_16962,N_16807);
nand U17019 (N_17019,N_16994,N_16812);
or U17020 (N_17020,N_16973,N_16972);
nand U17021 (N_17021,N_16838,N_16800);
and U17022 (N_17022,N_16940,N_16956);
or U17023 (N_17023,N_16937,N_16943);
and U17024 (N_17024,N_16821,N_16939);
nand U17025 (N_17025,N_16866,N_16928);
and U17026 (N_17026,N_16833,N_16883);
xor U17027 (N_17027,N_16999,N_16864);
nand U17028 (N_17028,N_16828,N_16886);
nand U17029 (N_17029,N_16987,N_16945);
xor U17030 (N_17030,N_16970,N_16868);
and U17031 (N_17031,N_16808,N_16875);
and U17032 (N_17032,N_16934,N_16922);
nor U17033 (N_17033,N_16948,N_16913);
nand U17034 (N_17034,N_16904,N_16845);
xnor U17035 (N_17035,N_16839,N_16946);
and U17036 (N_17036,N_16984,N_16831);
nor U17037 (N_17037,N_16846,N_16813);
xor U17038 (N_17038,N_16977,N_16914);
xnor U17039 (N_17039,N_16975,N_16835);
or U17040 (N_17040,N_16852,N_16888);
and U17041 (N_17041,N_16836,N_16907);
xor U17042 (N_17042,N_16860,N_16992);
or U17043 (N_17043,N_16911,N_16997);
xnor U17044 (N_17044,N_16905,N_16855);
or U17045 (N_17045,N_16861,N_16877);
nor U17046 (N_17046,N_16874,N_16912);
and U17047 (N_17047,N_16853,N_16957);
nor U17048 (N_17048,N_16899,N_16891);
and U17049 (N_17049,N_16989,N_16986);
or U17050 (N_17050,N_16885,N_16961);
nand U17051 (N_17051,N_16993,N_16871);
nand U17052 (N_17052,N_16932,N_16978);
and U17053 (N_17053,N_16817,N_16941);
and U17054 (N_17054,N_16894,N_16903);
or U17055 (N_17055,N_16867,N_16806);
or U17056 (N_17056,N_16859,N_16837);
xnor U17057 (N_17057,N_16804,N_16842);
and U17058 (N_17058,N_16980,N_16832);
nor U17059 (N_17059,N_16869,N_16840);
or U17060 (N_17060,N_16927,N_16926);
xor U17061 (N_17061,N_16920,N_16983);
xnor U17062 (N_17062,N_16818,N_16950);
or U17063 (N_17063,N_16917,N_16960);
or U17064 (N_17064,N_16955,N_16876);
or U17065 (N_17065,N_16805,N_16981);
or U17066 (N_17066,N_16889,N_16809);
and U17067 (N_17067,N_16900,N_16998);
nor U17068 (N_17068,N_16976,N_16982);
and U17069 (N_17069,N_16965,N_16974);
or U17070 (N_17070,N_16930,N_16803);
nand U17071 (N_17071,N_16834,N_16949);
xor U17072 (N_17072,N_16951,N_16959);
nor U17073 (N_17073,N_16908,N_16879);
xnor U17074 (N_17074,N_16995,N_16858);
or U17075 (N_17075,N_16963,N_16979);
and U17076 (N_17076,N_16873,N_16826);
nand U17077 (N_17077,N_16863,N_16933);
nor U17078 (N_17078,N_16848,N_16958);
and U17079 (N_17079,N_16896,N_16872);
nand U17080 (N_17080,N_16851,N_16942);
nor U17081 (N_17081,N_16811,N_16890);
or U17082 (N_17082,N_16844,N_16865);
and U17083 (N_17083,N_16954,N_16952);
and U17084 (N_17084,N_16801,N_16893);
xor U17085 (N_17085,N_16857,N_16944);
nor U17086 (N_17086,N_16990,N_16815);
xnor U17087 (N_17087,N_16985,N_16882);
and U17088 (N_17088,N_16910,N_16830);
and U17089 (N_17089,N_16897,N_16969);
xor U17090 (N_17090,N_16929,N_16916);
nand U17091 (N_17091,N_16824,N_16909);
xnor U17092 (N_17092,N_16971,N_16996);
nor U17093 (N_17093,N_16966,N_16823);
or U17094 (N_17094,N_16924,N_16802);
nor U17095 (N_17095,N_16819,N_16887);
or U17096 (N_17096,N_16967,N_16850);
or U17097 (N_17097,N_16902,N_16822);
nand U17098 (N_17098,N_16921,N_16947);
and U17099 (N_17099,N_16862,N_16915);
nor U17100 (N_17100,N_16870,N_16818);
nand U17101 (N_17101,N_16935,N_16917);
and U17102 (N_17102,N_16988,N_16917);
xor U17103 (N_17103,N_16850,N_16825);
and U17104 (N_17104,N_16981,N_16839);
xor U17105 (N_17105,N_16821,N_16809);
xnor U17106 (N_17106,N_16967,N_16859);
nor U17107 (N_17107,N_16967,N_16840);
or U17108 (N_17108,N_16990,N_16855);
nor U17109 (N_17109,N_16955,N_16960);
nand U17110 (N_17110,N_16908,N_16871);
nor U17111 (N_17111,N_16937,N_16819);
nor U17112 (N_17112,N_16816,N_16933);
xor U17113 (N_17113,N_16954,N_16919);
nand U17114 (N_17114,N_16874,N_16944);
and U17115 (N_17115,N_16820,N_16877);
xnor U17116 (N_17116,N_16847,N_16816);
and U17117 (N_17117,N_16879,N_16952);
and U17118 (N_17118,N_16938,N_16962);
xnor U17119 (N_17119,N_16915,N_16958);
or U17120 (N_17120,N_16943,N_16808);
nand U17121 (N_17121,N_16956,N_16861);
or U17122 (N_17122,N_16988,N_16997);
nand U17123 (N_17123,N_16977,N_16925);
nor U17124 (N_17124,N_16878,N_16967);
nand U17125 (N_17125,N_16903,N_16835);
xor U17126 (N_17126,N_16831,N_16930);
and U17127 (N_17127,N_16860,N_16977);
xor U17128 (N_17128,N_16914,N_16898);
and U17129 (N_17129,N_16911,N_16815);
nor U17130 (N_17130,N_16848,N_16943);
xor U17131 (N_17131,N_16981,N_16869);
nand U17132 (N_17132,N_16982,N_16826);
and U17133 (N_17133,N_16829,N_16987);
and U17134 (N_17134,N_16943,N_16880);
or U17135 (N_17135,N_16856,N_16903);
nand U17136 (N_17136,N_16921,N_16956);
nand U17137 (N_17137,N_16873,N_16848);
and U17138 (N_17138,N_16939,N_16848);
and U17139 (N_17139,N_16872,N_16848);
nand U17140 (N_17140,N_16914,N_16917);
and U17141 (N_17141,N_16938,N_16992);
nand U17142 (N_17142,N_16927,N_16832);
nand U17143 (N_17143,N_16864,N_16876);
and U17144 (N_17144,N_16977,N_16993);
or U17145 (N_17145,N_16998,N_16804);
xor U17146 (N_17146,N_16847,N_16905);
nand U17147 (N_17147,N_16958,N_16907);
and U17148 (N_17148,N_16855,N_16805);
and U17149 (N_17149,N_16872,N_16903);
xnor U17150 (N_17150,N_16937,N_16914);
xor U17151 (N_17151,N_16955,N_16901);
nor U17152 (N_17152,N_16873,N_16863);
nor U17153 (N_17153,N_16996,N_16942);
nand U17154 (N_17154,N_16809,N_16986);
nand U17155 (N_17155,N_16863,N_16989);
and U17156 (N_17156,N_16946,N_16871);
nor U17157 (N_17157,N_16837,N_16916);
nor U17158 (N_17158,N_16860,N_16989);
nor U17159 (N_17159,N_16836,N_16999);
nand U17160 (N_17160,N_16853,N_16803);
or U17161 (N_17161,N_16878,N_16882);
nor U17162 (N_17162,N_16817,N_16982);
or U17163 (N_17163,N_16968,N_16966);
or U17164 (N_17164,N_16846,N_16946);
and U17165 (N_17165,N_16854,N_16886);
or U17166 (N_17166,N_16997,N_16888);
and U17167 (N_17167,N_16851,N_16922);
nand U17168 (N_17168,N_16873,N_16989);
xor U17169 (N_17169,N_16976,N_16860);
xor U17170 (N_17170,N_16891,N_16863);
nand U17171 (N_17171,N_16918,N_16949);
xor U17172 (N_17172,N_16830,N_16873);
xnor U17173 (N_17173,N_16868,N_16940);
or U17174 (N_17174,N_16822,N_16938);
and U17175 (N_17175,N_16964,N_16950);
or U17176 (N_17176,N_16970,N_16958);
xnor U17177 (N_17177,N_16893,N_16839);
nor U17178 (N_17178,N_16971,N_16915);
and U17179 (N_17179,N_16811,N_16910);
or U17180 (N_17180,N_16897,N_16916);
nor U17181 (N_17181,N_16897,N_16805);
nand U17182 (N_17182,N_16892,N_16896);
and U17183 (N_17183,N_16952,N_16883);
xnor U17184 (N_17184,N_16955,N_16997);
nor U17185 (N_17185,N_16936,N_16891);
xor U17186 (N_17186,N_16980,N_16825);
or U17187 (N_17187,N_16875,N_16996);
xor U17188 (N_17188,N_16854,N_16957);
nand U17189 (N_17189,N_16820,N_16913);
nand U17190 (N_17190,N_16904,N_16956);
xnor U17191 (N_17191,N_16939,N_16956);
and U17192 (N_17192,N_16949,N_16816);
nand U17193 (N_17193,N_16824,N_16931);
xor U17194 (N_17194,N_16957,N_16904);
nand U17195 (N_17195,N_16923,N_16935);
nand U17196 (N_17196,N_16944,N_16940);
xor U17197 (N_17197,N_16997,N_16846);
nor U17198 (N_17198,N_16994,N_16967);
and U17199 (N_17199,N_16866,N_16858);
nand U17200 (N_17200,N_17015,N_17181);
xor U17201 (N_17201,N_17113,N_17052);
or U17202 (N_17202,N_17062,N_17119);
and U17203 (N_17203,N_17196,N_17092);
xnor U17204 (N_17204,N_17093,N_17033);
or U17205 (N_17205,N_17109,N_17095);
and U17206 (N_17206,N_17107,N_17155);
or U17207 (N_17207,N_17054,N_17043);
xnor U17208 (N_17208,N_17182,N_17164);
or U17209 (N_17209,N_17058,N_17129);
nand U17210 (N_17210,N_17016,N_17106);
nor U17211 (N_17211,N_17032,N_17151);
xor U17212 (N_17212,N_17108,N_17040);
and U17213 (N_17213,N_17169,N_17031);
and U17214 (N_17214,N_17019,N_17004);
nand U17215 (N_17215,N_17179,N_17075);
nand U17216 (N_17216,N_17088,N_17023);
or U17217 (N_17217,N_17039,N_17166);
xnor U17218 (N_17218,N_17057,N_17186);
or U17219 (N_17219,N_17174,N_17190);
xnor U17220 (N_17220,N_17146,N_17120);
xnor U17221 (N_17221,N_17139,N_17042);
or U17222 (N_17222,N_17197,N_17020);
and U17223 (N_17223,N_17158,N_17098);
xor U17224 (N_17224,N_17142,N_17066);
xor U17225 (N_17225,N_17002,N_17150);
xor U17226 (N_17226,N_17105,N_17018);
nand U17227 (N_17227,N_17000,N_17188);
nor U17228 (N_17228,N_17017,N_17104);
xor U17229 (N_17229,N_17148,N_17135);
nor U17230 (N_17230,N_17102,N_17101);
nand U17231 (N_17231,N_17091,N_17086);
nand U17232 (N_17232,N_17007,N_17035);
nor U17233 (N_17233,N_17128,N_17021);
xnor U17234 (N_17234,N_17048,N_17080);
or U17235 (N_17235,N_17085,N_17143);
nor U17236 (N_17236,N_17083,N_17122);
xor U17237 (N_17237,N_17140,N_17127);
nand U17238 (N_17238,N_17082,N_17159);
nand U17239 (N_17239,N_17126,N_17116);
or U17240 (N_17240,N_17081,N_17157);
nand U17241 (N_17241,N_17074,N_17024);
and U17242 (N_17242,N_17100,N_17046);
or U17243 (N_17243,N_17010,N_17059);
xor U17244 (N_17244,N_17121,N_17027);
nor U17245 (N_17245,N_17044,N_17089);
xnor U17246 (N_17246,N_17110,N_17094);
nor U17247 (N_17247,N_17034,N_17029);
or U17248 (N_17248,N_17191,N_17193);
nor U17249 (N_17249,N_17096,N_17036);
or U17250 (N_17250,N_17051,N_17005);
or U17251 (N_17251,N_17008,N_17192);
and U17252 (N_17252,N_17115,N_17041);
xor U17253 (N_17253,N_17198,N_17171);
nor U17254 (N_17254,N_17117,N_17145);
or U17255 (N_17255,N_17177,N_17162);
and U17256 (N_17256,N_17047,N_17199);
nand U17257 (N_17257,N_17194,N_17136);
xor U17258 (N_17258,N_17103,N_17141);
nor U17259 (N_17259,N_17087,N_17003);
xnor U17260 (N_17260,N_17178,N_17056);
and U17261 (N_17261,N_17167,N_17001);
and U17262 (N_17262,N_17138,N_17124);
or U17263 (N_17263,N_17184,N_17133);
or U17264 (N_17264,N_17061,N_17183);
nand U17265 (N_17265,N_17045,N_17175);
and U17266 (N_17266,N_17065,N_17006);
or U17267 (N_17267,N_17154,N_17025);
nor U17268 (N_17268,N_17067,N_17070);
or U17269 (N_17269,N_17185,N_17079);
and U17270 (N_17270,N_17147,N_17189);
or U17271 (N_17271,N_17160,N_17195);
xnor U17272 (N_17272,N_17077,N_17013);
xor U17273 (N_17273,N_17030,N_17161);
or U17274 (N_17274,N_17187,N_17028);
xnor U17275 (N_17275,N_17172,N_17011);
or U17276 (N_17276,N_17073,N_17163);
xnor U17277 (N_17277,N_17038,N_17125);
nor U17278 (N_17278,N_17132,N_17037);
xor U17279 (N_17279,N_17055,N_17176);
and U17280 (N_17280,N_17168,N_17097);
nor U17281 (N_17281,N_17009,N_17123);
nor U17282 (N_17282,N_17152,N_17114);
or U17283 (N_17283,N_17180,N_17165);
xor U17284 (N_17284,N_17144,N_17090);
nor U17285 (N_17285,N_17173,N_17049);
nor U17286 (N_17286,N_17170,N_17137);
and U17287 (N_17287,N_17068,N_17026);
or U17288 (N_17288,N_17156,N_17084);
or U17289 (N_17289,N_17134,N_17131);
xnor U17290 (N_17290,N_17063,N_17099);
nand U17291 (N_17291,N_17060,N_17053);
xor U17292 (N_17292,N_17118,N_17153);
xnor U17293 (N_17293,N_17069,N_17078);
and U17294 (N_17294,N_17149,N_17012);
xor U17295 (N_17295,N_17072,N_17112);
xor U17296 (N_17296,N_17050,N_17071);
xnor U17297 (N_17297,N_17014,N_17064);
and U17298 (N_17298,N_17130,N_17022);
nand U17299 (N_17299,N_17111,N_17076);
or U17300 (N_17300,N_17069,N_17057);
nand U17301 (N_17301,N_17028,N_17060);
nor U17302 (N_17302,N_17096,N_17073);
xnor U17303 (N_17303,N_17118,N_17181);
nor U17304 (N_17304,N_17131,N_17003);
nand U17305 (N_17305,N_17005,N_17089);
nand U17306 (N_17306,N_17131,N_17088);
nand U17307 (N_17307,N_17166,N_17016);
xnor U17308 (N_17308,N_17079,N_17129);
nand U17309 (N_17309,N_17047,N_17128);
nor U17310 (N_17310,N_17043,N_17186);
xor U17311 (N_17311,N_17008,N_17060);
nand U17312 (N_17312,N_17198,N_17043);
nor U17313 (N_17313,N_17177,N_17104);
nand U17314 (N_17314,N_17171,N_17003);
nand U17315 (N_17315,N_17097,N_17095);
nand U17316 (N_17316,N_17065,N_17036);
or U17317 (N_17317,N_17122,N_17106);
xor U17318 (N_17318,N_17041,N_17050);
and U17319 (N_17319,N_17190,N_17130);
xnor U17320 (N_17320,N_17026,N_17028);
nand U17321 (N_17321,N_17109,N_17188);
and U17322 (N_17322,N_17149,N_17033);
nand U17323 (N_17323,N_17032,N_17196);
and U17324 (N_17324,N_17173,N_17085);
nand U17325 (N_17325,N_17130,N_17178);
or U17326 (N_17326,N_17014,N_17013);
nor U17327 (N_17327,N_17084,N_17185);
nand U17328 (N_17328,N_17096,N_17149);
or U17329 (N_17329,N_17024,N_17032);
nor U17330 (N_17330,N_17119,N_17083);
nor U17331 (N_17331,N_17082,N_17033);
nor U17332 (N_17332,N_17109,N_17008);
and U17333 (N_17333,N_17119,N_17043);
nand U17334 (N_17334,N_17140,N_17093);
nand U17335 (N_17335,N_17189,N_17028);
or U17336 (N_17336,N_17156,N_17161);
xor U17337 (N_17337,N_17092,N_17035);
nand U17338 (N_17338,N_17040,N_17081);
nor U17339 (N_17339,N_17039,N_17163);
nand U17340 (N_17340,N_17016,N_17090);
nor U17341 (N_17341,N_17092,N_17098);
nand U17342 (N_17342,N_17103,N_17148);
nor U17343 (N_17343,N_17119,N_17032);
nand U17344 (N_17344,N_17079,N_17043);
nand U17345 (N_17345,N_17035,N_17037);
and U17346 (N_17346,N_17059,N_17179);
nor U17347 (N_17347,N_17083,N_17124);
nor U17348 (N_17348,N_17062,N_17049);
and U17349 (N_17349,N_17065,N_17074);
nor U17350 (N_17350,N_17183,N_17015);
or U17351 (N_17351,N_17114,N_17126);
xnor U17352 (N_17352,N_17118,N_17086);
and U17353 (N_17353,N_17189,N_17044);
nor U17354 (N_17354,N_17147,N_17091);
or U17355 (N_17355,N_17103,N_17050);
nand U17356 (N_17356,N_17118,N_17017);
and U17357 (N_17357,N_17084,N_17049);
xnor U17358 (N_17358,N_17152,N_17161);
or U17359 (N_17359,N_17170,N_17093);
nand U17360 (N_17360,N_17150,N_17057);
xor U17361 (N_17361,N_17114,N_17096);
or U17362 (N_17362,N_17184,N_17162);
and U17363 (N_17363,N_17143,N_17079);
nor U17364 (N_17364,N_17055,N_17187);
nand U17365 (N_17365,N_17196,N_17178);
and U17366 (N_17366,N_17079,N_17179);
nand U17367 (N_17367,N_17056,N_17055);
nand U17368 (N_17368,N_17067,N_17177);
nor U17369 (N_17369,N_17153,N_17120);
and U17370 (N_17370,N_17170,N_17034);
or U17371 (N_17371,N_17118,N_17023);
xnor U17372 (N_17372,N_17028,N_17092);
xnor U17373 (N_17373,N_17022,N_17193);
nor U17374 (N_17374,N_17093,N_17057);
or U17375 (N_17375,N_17082,N_17182);
xor U17376 (N_17376,N_17122,N_17023);
and U17377 (N_17377,N_17136,N_17123);
nor U17378 (N_17378,N_17031,N_17033);
and U17379 (N_17379,N_17100,N_17087);
or U17380 (N_17380,N_17164,N_17005);
and U17381 (N_17381,N_17108,N_17187);
xor U17382 (N_17382,N_17148,N_17172);
nand U17383 (N_17383,N_17183,N_17107);
nand U17384 (N_17384,N_17042,N_17161);
nand U17385 (N_17385,N_17132,N_17145);
xnor U17386 (N_17386,N_17066,N_17022);
xor U17387 (N_17387,N_17074,N_17182);
nor U17388 (N_17388,N_17135,N_17044);
or U17389 (N_17389,N_17078,N_17178);
nand U17390 (N_17390,N_17140,N_17067);
xnor U17391 (N_17391,N_17122,N_17073);
and U17392 (N_17392,N_17134,N_17055);
nor U17393 (N_17393,N_17060,N_17066);
nand U17394 (N_17394,N_17143,N_17091);
nor U17395 (N_17395,N_17075,N_17146);
nand U17396 (N_17396,N_17099,N_17178);
xnor U17397 (N_17397,N_17192,N_17031);
or U17398 (N_17398,N_17139,N_17022);
nand U17399 (N_17399,N_17135,N_17150);
xnor U17400 (N_17400,N_17223,N_17317);
nand U17401 (N_17401,N_17355,N_17333);
or U17402 (N_17402,N_17205,N_17284);
xnor U17403 (N_17403,N_17294,N_17263);
and U17404 (N_17404,N_17329,N_17296);
xnor U17405 (N_17405,N_17328,N_17270);
xor U17406 (N_17406,N_17356,N_17206);
nor U17407 (N_17407,N_17334,N_17342);
or U17408 (N_17408,N_17299,N_17245);
xor U17409 (N_17409,N_17221,N_17248);
nand U17410 (N_17410,N_17235,N_17277);
xnor U17411 (N_17411,N_17272,N_17226);
nand U17412 (N_17412,N_17351,N_17394);
or U17413 (N_17413,N_17255,N_17393);
or U17414 (N_17414,N_17241,N_17281);
and U17415 (N_17415,N_17321,N_17327);
nand U17416 (N_17416,N_17256,N_17212);
nand U17417 (N_17417,N_17259,N_17332);
xor U17418 (N_17418,N_17219,N_17319);
and U17419 (N_17419,N_17340,N_17210);
or U17420 (N_17420,N_17268,N_17373);
nand U17421 (N_17421,N_17273,N_17335);
and U17422 (N_17422,N_17252,N_17365);
and U17423 (N_17423,N_17280,N_17295);
and U17424 (N_17424,N_17282,N_17388);
nand U17425 (N_17425,N_17378,N_17303);
nand U17426 (N_17426,N_17361,N_17369);
and U17427 (N_17427,N_17208,N_17311);
nor U17428 (N_17428,N_17374,N_17238);
and U17429 (N_17429,N_17204,N_17387);
xor U17430 (N_17430,N_17211,N_17398);
xor U17431 (N_17431,N_17309,N_17331);
nand U17432 (N_17432,N_17290,N_17292);
nor U17433 (N_17433,N_17260,N_17242);
or U17434 (N_17434,N_17217,N_17392);
and U17435 (N_17435,N_17315,N_17379);
nand U17436 (N_17436,N_17289,N_17276);
nand U17437 (N_17437,N_17322,N_17370);
or U17438 (N_17438,N_17341,N_17354);
and U17439 (N_17439,N_17213,N_17330);
nand U17440 (N_17440,N_17215,N_17269);
and U17441 (N_17441,N_17337,N_17318);
nor U17442 (N_17442,N_17357,N_17375);
xor U17443 (N_17443,N_17232,N_17266);
and U17444 (N_17444,N_17310,N_17262);
xor U17445 (N_17445,N_17229,N_17222);
or U17446 (N_17446,N_17291,N_17267);
xnor U17447 (N_17447,N_17233,N_17350);
or U17448 (N_17448,N_17344,N_17390);
xnor U17449 (N_17449,N_17326,N_17293);
and U17450 (N_17450,N_17325,N_17249);
and U17451 (N_17451,N_17367,N_17381);
nand U17452 (N_17452,N_17384,N_17336);
nand U17453 (N_17453,N_17275,N_17389);
xor U17454 (N_17454,N_17320,N_17231);
and U17455 (N_17455,N_17253,N_17352);
nand U17456 (N_17456,N_17363,N_17230);
and U17457 (N_17457,N_17368,N_17225);
xnor U17458 (N_17458,N_17323,N_17224);
xor U17459 (N_17459,N_17371,N_17302);
xor U17460 (N_17460,N_17271,N_17385);
nand U17461 (N_17461,N_17250,N_17261);
nand U17462 (N_17462,N_17244,N_17397);
xnor U17463 (N_17463,N_17377,N_17220);
nor U17464 (N_17464,N_17307,N_17339);
nor U17465 (N_17465,N_17236,N_17301);
nand U17466 (N_17466,N_17288,N_17300);
or U17467 (N_17467,N_17264,N_17316);
nand U17468 (N_17468,N_17243,N_17346);
nand U17469 (N_17469,N_17338,N_17201);
and U17470 (N_17470,N_17254,N_17274);
or U17471 (N_17471,N_17366,N_17251);
nand U17472 (N_17472,N_17283,N_17306);
nor U17473 (N_17473,N_17237,N_17234);
nand U17474 (N_17474,N_17218,N_17380);
nor U17475 (N_17475,N_17396,N_17214);
xor U17476 (N_17476,N_17358,N_17324);
and U17477 (N_17477,N_17209,N_17246);
and U17478 (N_17478,N_17298,N_17376);
and U17479 (N_17479,N_17258,N_17359);
and U17480 (N_17480,N_17399,N_17349);
and U17481 (N_17481,N_17239,N_17216);
nand U17482 (N_17482,N_17313,N_17362);
nand U17483 (N_17483,N_17360,N_17395);
or U17484 (N_17484,N_17257,N_17278);
nor U17485 (N_17485,N_17353,N_17383);
xnor U17486 (N_17486,N_17312,N_17347);
and U17487 (N_17487,N_17203,N_17305);
and U17488 (N_17488,N_17279,N_17202);
nand U17489 (N_17489,N_17200,N_17227);
and U17490 (N_17490,N_17314,N_17386);
nand U17491 (N_17491,N_17304,N_17207);
nor U17492 (N_17492,N_17391,N_17265);
or U17493 (N_17493,N_17372,N_17247);
and U17494 (N_17494,N_17308,N_17382);
or U17495 (N_17495,N_17364,N_17343);
or U17496 (N_17496,N_17348,N_17286);
nand U17497 (N_17497,N_17287,N_17345);
xnor U17498 (N_17498,N_17285,N_17240);
xnor U17499 (N_17499,N_17228,N_17297);
and U17500 (N_17500,N_17288,N_17226);
nand U17501 (N_17501,N_17390,N_17367);
or U17502 (N_17502,N_17209,N_17386);
nor U17503 (N_17503,N_17386,N_17221);
nand U17504 (N_17504,N_17241,N_17282);
and U17505 (N_17505,N_17201,N_17229);
xor U17506 (N_17506,N_17200,N_17312);
nand U17507 (N_17507,N_17222,N_17374);
xor U17508 (N_17508,N_17218,N_17288);
nand U17509 (N_17509,N_17216,N_17240);
and U17510 (N_17510,N_17208,N_17396);
or U17511 (N_17511,N_17283,N_17303);
and U17512 (N_17512,N_17245,N_17319);
nor U17513 (N_17513,N_17273,N_17389);
nor U17514 (N_17514,N_17220,N_17208);
and U17515 (N_17515,N_17214,N_17318);
nor U17516 (N_17516,N_17362,N_17340);
nand U17517 (N_17517,N_17382,N_17216);
xnor U17518 (N_17518,N_17204,N_17344);
or U17519 (N_17519,N_17226,N_17284);
and U17520 (N_17520,N_17353,N_17272);
and U17521 (N_17521,N_17358,N_17293);
xnor U17522 (N_17522,N_17202,N_17376);
nand U17523 (N_17523,N_17242,N_17207);
nand U17524 (N_17524,N_17265,N_17285);
xor U17525 (N_17525,N_17348,N_17311);
and U17526 (N_17526,N_17217,N_17387);
xor U17527 (N_17527,N_17273,N_17314);
nand U17528 (N_17528,N_17227,N_17360);
nand U17529 (N_17529,N_17280,N_17326);
nor U17530 (N_17530,N_17228,N_17206);
and U17531 (N_17531,N_17222,N_17227);
xor U17532 (N_17532,N_17345,N_17209);
nor U17533 (N_17533,N_17345,N_17330);
nor U17534 (N_17534,N_17375,N_17317);
nand U17535 (N_17535,N_17357,N_17326);
xnor U17536 (N_17536,N_17217,N_17390);
or U17537 (N_17537,N_17363,N_17241);
or U17538 (N_17538,N_17203,N_17332);
nand U17539 (N_17539,N_17365,N_17288);
nand U17540 (N_17540,N_17384,N_17273);
and U17541 (N_17541,N_17301,N_17251);
xor U17542 (N_17542,N_17252,N_17379);
xor U17543 (N_17543,N_17257,N_17273);
or U17544 (N_17544,N_17368,N_17232);
nand U17545 (N_17545,N_17218,N_17254);
and U17546 (N_17546,N_17290,N_17364);
xnor U17547 (N_17547,N_17368,N_17227);
xnor U17548 (N_17548,N_17260,N_17209);
nand U17549 (N_17549,N_17261,N_17352);
xnor U17550 (N_17550,N_17363,N_17339);
nand U17551 (N_17551,N_17292,N_17227);
or U17552 (N_17552,N_17292,N_17397);
xor U17553 (N_17553,N_17245,N_17214);
and U17554 (N_17554,N_17374,N_17273);
xnor U17555 (N_17555,N_17240,N_17352);
xnor U17556 (N_17556,N_17230,N_17244);
and U17557 (N_17557,N_17399,N_17352);
nor U17558 (N_17558,N_17379,N_17320);
xor U17559 (N_17559,N_17241,N_17255);
and U17560 (N_17560,N_17278,N_17383);
nand U17561 (N_17561,N_17293,N_17377);
nand U17562 (N_17562,N_17342,N_17270);
nor U17563 (N_17563,N_17372,N_17315);
and U17564 (N_17564,N_17388,N_17325);
or U17565 (N_17565,N_17392,N_17374);
xnor U17566 (N_17566,N_17229,N_17209);
nor U17567 (N_17567,N_17205,N_17203);
or U17568 (N_17568,N_17256,N_17239);
xnor U17569 (N_17569,N_17334,N_17301);
xnor U17570 (N_17570,N_17234,N_17348);
nor U17571 (N_17571,N_17386,N_17279);
nand U17572 (N_17572,N_17371,N_17283);
xor U17573 (N_17573,N_17258,N_17307);
and U17574 (N_17574,N_17330,N_17333);
nand U17575 (N_17575,N_17346,N_17234);
and U17576 (N_17576,N_17337,N_17266);
nor U17577 (N_17577,N_17265,N_17225);
nor U17578 (N_17578,N_17334,N_17203);
nor U17579 (N_17579,N_17321,N_17230);
nor U17580 (N_17580,N_17234,N_17375);
or U17581 (N_17581,N_17376,N_17281);
and U17582 (N_17582,N_17340,N_17386);
or U17583 (N_17583,N_17372,N_17201);
or U17584 (N_17584,N_17392,N_17203);
nor U17585 (N_17585,N_17201,N_17284);
nor U17586 (N_17586,N_17338,N_17371);
and U17587 (N_17587,N_17316,N_17326);
xor U17588 (N_17588,N_17262,N_17326);
or U17589 (N_17589,N_17357,N_17365);
nor U17590 (N_17590,N_17354,N_17258);
xnor U17591 (N_17591,N_17342,N_17288);
or U17592 (N_17592,N_17296,N_17225);
or U17593 (N_17593,N_17289,N_17311);
nor U17594 (N_17594,N_17207,N_17339);
nor U17595 (N_17595,N_17204,N_17366);
xnor U17596 (N_17596,N_17275,N_17252);
nor U17597 (N_17597,N_17382,N_17275);
nor U17598 (N_17598,N_17342,N_17289);
and U17599 (N_17599,N_17235,N_17228);
xor U17600 (N_17600,N_17412,N_17420);
and U17601 (N_17601,N_17590,N_17469);
and U17602 (N_17602,N_17425,N_17526);
nand U17603 (N_17603,N_17500,N_17575);
xor U17604 (N_17604,N_17539,N_17553);
or U17605 (N_17605,N_17536,N_17414);
or U17606 (N_17606,N_17451,N_17475);
or U17607 (N_17607,N_17548,N_17540);
xnor U17608 (N_17608,N_17525,N_17458);
nor U17609 (N_17609,N_17545,N_17503);
or U17610 (N_17610,N_17421,N_17441);
nor U17611 (N_17611,N_17440,N_17442);
nor U17612 (N_17612,N_17597,N_17416);
nand U17613 (N_17613,N_17494,N_17462);
or U17614 (N_17614,N_17417,N_17479);
xor U17615 (N_17615,N_17562,N_17543);
or U17616 (N_17616,N_17507,N_17559);
or U17617 (N_17617,N_17404,N_17487);
nand U17618 (N_17618,N_17484,N_17413);
nor U17619 (N_17619,N_17527,N_17497);
nor U17620 (N_17620,N_17529,N_17549);
and U17621 (N_17621,N_17589,N_17521);
nand U17622 (N_17622,N_17599,N_17501);
xnor U17623 (N_17623,N_17431,N_17502);
nand U17624 (N_17624,N_17505,N_17450);
and U17625 (N_17625,N_17433,N_17568);
or U17626 (N_17626,N_17513,N_17415);
or U17627 (N_17627,N_17511,N_17522);
or U17628 (N_17628,N_17483,N_17532);
nor U17629 (N_17629,N_17504,N_17499);
and U17630 (N_17630,N_17470,N_17580);
and U17631 (N_17631,N_17574,N_17436);
nand U17632 (N_17632,N_17556,N_17535);
nor U17633 (N_17633,N_17476,N_17403);
nand U17634 (N_17634,N_17578,N_17498);
nor U17635 (N_17635,N_17456,N_17508);
or U17636 (N_17636,N_17554,N_17520);
and U17637 (N_17637,N_17591,N_17444);
or U17638 (N_17638,N_17424,N_17409);
nor U17639 (N_17639,N_17512,N_17465);
nand U17640 (N_17640,N_17588,N_17496);
nand U17641 (N_17641,N_17472,N_17452);
and U17642 (N_17642,N_17432,N_17422);
nor U17643 (N_17643,N_17405,N_17555);
or U17644 (N_17644,N_17473,N_17427);
and U17645 (N_17645,N_17552,N_17466);
nand U17646 (N_17646,N_17402,N_17524);
nor U17647 (N_17647,N_17445,N_17565);
or U17648 (N_17648,N_17534,N_17460);
or U17649 (N_17649,N_17530,N_17448);
or U17650 (N_17650,N_17546,N_17506);
or U17651 (N_17651,N_17523,N_17485);
and U17652 (N_17652,N_17592,N_17429);
and U17653 (N_17653,N_17482,N_17544);
or U17654 (N_17654,N_17514,N_17517);
nand U17655 (N_17655,N_17573,N_17426);
and U17656 (N_17656,N_17576,N_17594);
nor U17657 (N_17657,N_17454,N_17410);
and U17658 (N_17658,N_17557,N_17437);
nand U17659 (N_17659,N_17583,N_17558);
or U17660 (N_17660,N_17490,N_17489);
nand U17661 (N_17661,N_17449,N_17519);
xnor U17662 (N_17662,N_17551,N_17510);
nor U17663 (N_17663,N_17480,N_17538);
and U17664 (N_17664,N_17537,N_17581);
or U17665 (N_17665,N_17481,N_17515);
xor U17666 (N_17666,N_17459,N_17407);
nor U17667 (N_17667,N_17474,N_17492);
or U17668 (N_17668,N_17438,N_17509);
and U17669 (N_17669,N_17443,N_17430);
nor U17670 (N_17670,N_17406,N_17518);
xnor U17671 (N_17671,N_17547,N_17563);
nor U17672 (N_17672,N_17572,N_17457);
or U17673 (N_17673,N_17486,N_17477);
or U17674 (N_17674,N_17418,N_17435);
nand U17675 (N_17675,N_17491,N_17587);
and U17676 (N_17676,N_17439,N_17408);
nand U17677 (N_17677,N_17495,N_17595);
nand U17678 (N_17678,N_17579,N_17478);
nor U17679 (N_17679,N_17455,N_17400);
nand U17680 (N_17680,N_17434,N_17453);
and U17681 (N_17681,N_17423,N_17564);
or U17682 (N_17682,N_17528,N_17560);
nand U17683 (N_17683,N_17566,N_17446);
or U17684 (N_17684,N_17533,N_17596);
xnor U17685 (N_17685,N_17577,N_17428);
nor U17686 (N_17686,N_17488,N_17550);
or U17687 (N_17687,N_17593,N_17471);
xor U17688 (N_17688,N_17464,N_17586);
and U17689 (N_17689,N_17493,N_17531);
and U17690 (N_17690,N_17542,N_17463);
or U17691 (N_17691,N_17569,N_17401);
nand U17692 (N_17692,N_17467,N_17516);
xnor U17693 (N_17693,N_17419,N_17570);
and U17694 (N_17694,N_17411,N_17584);
nor U17695 (N_17695,N_17447,N_17582);
or U17696 (N_17696,N_17571,N_17468);
xnor U17697 (N_17697,N_17585,N_17561);
or U17698 (N_17698,N_17567,N_17598);
nand U17699 (N_17699,N_17541,N_17461);
nor U17700 (N_17700,N_17494,N_17410);
xor U17701 (N_17701,N_17506,N_17509);
nor U17702 (N_17702,N_17449,N_17562);
xor U17703 (N_17703,N_17569,N_17404);
and U17704 (N_17704,N_17562,N_17440);
xnor U17705 (N_17705,N_17477,N_17529);
or U17706 (N_17706,N_17581,N_17501);
or U17707 (N_17707,N_17553,N_17597);
xor U17708 (N_17708,N_17456,N_17547);
or U17709 (N_17709,N_17568,N_17445);
or U17710 (N_17710,N_17427,N_17411);
or U17711 (N_17711,N_17486,N_17501);
nand U17712 (N_17712,N_17595,N_17550);
xor U17713 (N_17713,N_17561,N_17513);
xor U17714 (N_17714,N_17460,N_17459);
xnor U17715 (N_17715,N_17411,N_17444);
and U17716 (N_17716,N_17432,N_17539);
and U17717 (N_17717,N_17444,N_17461);
xnor U17718 (N_17718,N_17557,N_17440);
and U17719 (N_17719,N_17418,N_17533);
or U17720 (N_17720,N_17477,N_17450);
xor U17721 (N_17721,N_17497,N_17572);
nor U17722 (N_17722,N_17434,N_17494);
nor U17723 (N_17723,N_17510,N_17524);
nor U17724 (N_17724,N_17458,N_17586);
nor U17725 (N_17725,N_17478,N_17538);
or U17726 (N_17726,N_17440,N_17469);
and U17727 (N_17727,N_17571,N_17435);
or U17728 (N_17728,N_17407,N_17518);
nor U17729 (N_17729,N_17450,N_17516);
xor U17730 (N_17730,N_17596,N_17552);
xor U17731 (N_17731,N_17542,N_17401);
nor U17732 (N_17732,N_17429,N_17498);
xnor U17733 (N_17733,N_17503,N_17493);
nor U17734 (N_17734,N_17486,N_17498);
xor U17735 (N_17735,N_17464,N_17491);
and U17736 (N_17736,N_17411,N_17491);
and U17737 (N_17737,N_17458,N_17491);
xnor U17738 (N_17738,N_17476,N_17590);
or U17739 (N_17739,N_17593,N_17445);
nand U17740 (N_17740,N_17471,N_17582);
nor U17741 (N_17741,N_17438,N_17484);
nor U17742 (N_17742,N_17424,N_17595);
xor U17743 (N_17743,N_17499,N_17417);
nor U17744 (N_17744,N_17513,N_17464);
and U17745 (N_17745,N_17451,N_17427);
or U17746 (N_17746,N_17442,N_17490);
nor U17747 (N_17747,N_17529,N_17433);
and U17748 (N_17748,N_17468,N_17463);
nand U17749 (N_17749,N_17507,N_17586);
and U17750 (N_17750,N_17499,N_17570);
xnor U17751 (N_17751,N_17498,N_17534);
xnor U17752 (N_17752,N_17545,N_17401);
or U17753 (N_17753,N_17478,N_17408);
xnor U17754 (N_17754,N_17580,N_17546);
and U17755 (N_17755,N_17449,N_17506);
or U17756 (N_17756,N_17586,N_17476);
xnor U17757 (N_17757,N_17492,N_17456);
nor U17758 (N_17758,N_17461,N_17417);
and U17759 (N_17759,N_17409,N_17548);
or U17760 (N_17760,N_17433,N_17465);
xnor U17761 (N_17761,N_17572,N_17504);
and U17762 (N_17762,N_17506,N_17513);
or U17763 (N_17763,N_17459,N_17468);
nand U17764 (N_17764,N_17500,N_17548);
and U17765 (N_17765,N_17482,N_17481);
xor U17766 (N_17766,N_17418,N_17519);
and U17767 (N_17767,N_17587,N_17400);
nand U17768 (N_17768,N_17466,N_17595);
nand U17769 (N_17769,N_17452,N_17432);
xor U17770 (N_17770,N_17424,N_17480);
nor U17771 (N_17771,N_17425,N_17436);
xor U17772 (N_17772,N_17550,N_17421);
nor U17773 (N_17773,N_17522,N_17530);
and U17774 (N_17774,N_17516,N_17437);
or U17775 (N_17775,N_17430,N_17585);
or U17776 (N_17776,N_17448,N_17536);
nor U17777 (N_17777,N_17540,N_17437);
and U17778 (N_17778,N_17587,N_17415);
and U17779 (N_17779,N_17473,N_17444);
nor U17780 (N_17780,N_17465,N_17422);
nand U17781 (N_17781,N_17429,N_17551);
nor U17782 (N_17782,N_17538,N_17437);
nor U17783 (N_17783,N_17441,N_17599);
nor U17784 (N_17784,N_17571,N_17486);
and U17785 (N_17785,N_17503,N_17513);
xor U17786 (N_17786,N_17584,N_17441);
nand U17787 (N_17787,N_17523,N_17510);
and U17788 (N_17788,N_17406,N_17578);
or U17789 (N_17789,N_17471,N_17431);
or U17790 (N_17790,N_17538,N_17470);
nor U17791 (N_17791,N_17523,N_17513);
nand U17792 (N_17792,N_17420,N_17577);
xor U17793 (N_17793,N_17439,N_17406);
and U17794 (N_17794,N_17411,N_17539);
and U17795 (N_17795,N_17574,N_17440);
and U17796 (N_17796,N_17417,N_17523);
and U17797 (N_17797,N_17494,N_17594);
nor U17798 (N_17798,N_17549,N_17538);
xnor U17799 (N_17799,N_17442,N_17498);
nand U17800 (N_17800,N_17789,N_17716);
nand U17801 (N_17801,N_17684,N_17608);
nor U17802 (N_17802,N_17743,N_17739);
nor U17803 (N_17803,N_17711,N_17647);
nand U17804 (N_17804,N_17650,N_17610);
and U17805 (N_17805,N_17694,N_17685);
nand U17806 (N_17806,N_17756,N_17677);
or U17807 (N_17807,N_17662,N_17629);
or U17808 (N_17808,N_17776,N_17651);
nand U17809 (N_17809,N_17660,N_17753);
xor U17810 (N_17810,N_17736,N_17670);
xnor U17811 (N_17811,N_17751,N_17656);
xor U17812 (N_17812,N_17764,N_17715);
and U17813 (N_17813,N_17772,N_17795);
xnor U17814 (N_17814,N_17672,N_17737);
and U17815 (N_17815,N_17667,N_17769);
and U17816 (N_17816,N_17642,N_17696);
and U17817 (N_17817,N_17773,N_17771);
xor U17818 (N_17818,N_17678,N_17701);
xnor U17819 (N_17819,N_17750,N_17774);
xnor U17820 (N_17820,N_17641,N_17767);
nand U17821 (N_17821,N_17787,N_17698);
or U17822 (N_17822,N_17635,N_17652);
and U17823 (N_17823,N_17683,N_17665);
xor U17824 (N_17824,N_17605,N_17690);
nor U17825 (N_17825,N_17655,N_17617);
nor U17826 (N_17826,N_17797,N_17676);
nor U17827 (N_17827,N_17618,N_17719);
nor U17828 (N_17828,N_17745,N_17796);
xor U17829 (N_17829,N_17788,N_17661);
and U17830 (N_17830,N_17693,N_17744);
nor U17831 (N_17831,N_17620,N_17634);
and U17832 (N_17832,N_17637,N_17695);
xor U17833 (N_17833,N_17704,N_17758);
or U17834 (N_17834,N_17631,N_17724);
or U17835 (N_17835,N_17606,N_17786);
and U17836 (N_17836,N_17682,N_17626);
and U17837 (N_17837,N_17628,N_17609);
xor U17838 (N_17838,N_17777,N_17746);
nand U17839 (N_17839,N_17738,N_17791);
or U17840 (N_17840,N_17666,N_17681);
or U17841 (N_17841,N_17752,N_17679);
or U17842 (N_17842,N_17755,N_17705);
nor U17843 (N_17843,N_17760,N_17707);
and U17844 (N_17844,N_17768,N_17708);
or U17845 (N_17845,N_17747,N_17790);
nor U17846 (N_17846,N_17793,N_17675);
and U17847 (N_17847,N_17636,N_17785);
or U17848 (N_17848,N_17633,N_17680);
nor U17849 (N_17849,N_17603,N_17614);
or U17850 (N_17850,N_17639,N_17730);
or U17851 (N_17851,N_17691,N_17688);
nand U17852 (N_17852,N_17714,N_17733);
nand U17853 (N_17853,N_17709,N_17703);
or U17854 (N_17854,N_17762,N_17646);
and U17855 (N_17855,N_17754,N_17741);
nand U17856 (N_17856,N_17783,N_17657);
nand U17857 (N_17857,N_17731,N_17697);
xor U17858 (N_17858,N_17799,N_17638);
or U17859 (N_17859,N_17602,N_17726);
nand U17860 (N_17860,N_17723,N_17612);
and U17861 (N_17861,N_17601,N_17607);
nor U17862 (N_17862,N_17706,N_17669);
nand U17863 (N_17863,N_17692,N_17710);
and U17864 (N_17864,N_17780,N_17770);
nor U17865 (N_17865,N_17654,N_17713);
nor U17866 (N_17866,N_17664,N_17761);
or U17867 (N_17867,N_17632,N_17686);
or U17868 (N_17868,N_17748,N_17616);
xor U17869 (N_17869,N_17625,N_17643);
or U17870 (N_17870,N_17640,N_17749);
and U17871 (N_17871,N_17627,N_17781);
or U17872 (N_17872,N_17792,N_17778);
nand U17873 (N_17873,N_17630,N_17734);
or U17874 (N_17874,N_17673,N_17763);
and U17875 (N_17875,N_17622,N_17611);
or U17876 (N_17876,N_17712,N_17732);
xnor U17877 (N_17877,N_17623,N_17663);
and U17878 (N_17878,N_17619,N_17782);
nor U17879 (N_17879,N_17794,N_17728);
nor U17880 (N_17880,N_17721,N_17645);
nor U17881 (N_17881,N_17735,N_17798);
nand U17882 (N_17882,N_17765,N_17740);
or U17883 (N_17883,N_17700,N_17600);
xnor U17884 (N_17884,N_17615,N_17779);
xnor U17885 (N_17885,N_17613,N_17659);
or U17886 (N_17886,N_17757,N_17759);
nor U17887 (N_17887,N_17621,N_17775);
nor U17888 (N_17888,N_17687,N_17702);
nor U17889 (N_17889,N_17644,N_17653);
and U17890 (N_17890,N_17725,N_17742);
nor U17891 (N_17891,N_17766,N_17648);
and U17892 (N_17892,N_17784,N_17729);
and U17893 (N_17893,N_17699,N_17722);
xnor U17894 (N_17894,N_17720,N_17718);
nand U17895 (N_17895,N_17624,N_17658);
or U17896 (N_17896,N_17727,N_17649);
nor U17897 (N_17897,N_17604,N_17674);
nand U17898 (N_17898,N_17668,N_17717);
or U17899 (N_17899,N_17671,N_17689);
nand U17900 (N_17900,N_17629,N_17627);
and U17901 (N_17901,N_17773,N_17676);
nand U17902 (N_17902,N_17673,N_17787);
nand U17903 (N_17903,N_17697,N_17743);
or U17904 (N_17904,N_17664,N_17651);
nand U17905 (N_17905,N_17778,N_17679);
or U17906 (N_17906,N_17795,N_17790);
xnor U17907 (N_17907,N_17741,N_17641);
nand U17908 (N_17908,N_17627,N_17794);
or U17909 (N_17909,N_17640,N_17662);
and U17910 (N_17910,N_17614,N_17679);
xor U17911 (N_17911,N_17717,N_17629);
xnor U17912 (N_17912,N_17641,N_17687);
nand U17913 (N_17913,N_17735,N_17643);
and U17914 (N_17914,N_17689,N_17702);
and U17915 (N_17915,N_17724,N_17689);
and U17916 (N_17916,N_17663,N_17703);
nand U17917 (N_17917,N_17747,N_17732);
and U17918 (N_17918,N_17614,N_17694);
and U17919 (N_17919,N_17683,N_17711);
nand U17920 (N_17920,N_17733,N_17727);
nor U17921 (N_17921,N_17723,N_17708);
and U17922 (N_17922,N_17615,N_17784);
nor U17923 (N_17923,N_17610,N_17792);
nor U17924 (N_17924,N_17610,N_17645);
nor U17925 (N_17925,N_17677,N_17692);
nand U17926 (N_17926,N_17710,N_17752);
nand U17927 (N_17927,N_17685,N_17627);
nor U17928 (N_17928,N_17704,N_17764);
nand U17929 (N_17929,N_17612,N_17651);
nand U17930 (N_17930,N_17667,N_17719);
or U17931 (N_17931,N_17626,N_17604);
xor U17932 (N_17932,N_17661,N_17727);
xor U17933 (N_17933,N_17704,N_17678);
xor U17934 (N_17934,N_17698,N_17692);
or U17935 (N_17935,N_17628,N_17602);
nand U17936 (N_17936,N_17773,N_17613);
nor U17937 (N_17937,N_17697,N_17689);
and U17938 (N_17938,N_17630,N_17787);
or U17939 (N_17939,N_17793,N_17720);
and U17940 (N_17940,N_17794,N_17741);
or U17941 (N_17941,N_17610,N_17602);
xor U17942 (N_17942,N_17643,N_17660);
nor U17943 (N_17943,N_17685,N_17681);
nand U17944 (N_17944,N_17658,N_17703);
nor U17945 (N_17945,N_17670,N_17707);
and U17946 (N_17946,N_17671,N_17684);
nor U17947 (N_17947,N_17608,N_17776);
nand U17948 (N_17948,N_17708,N_17704);
xor U17949 (N_17949,N_17646,N_17630);
and U17950 (N_17950,N_17600,N_17774);
nor U17951 (N_17951,N_17674,N_17713);
nor U17952 (N_17952,N_17684,N_17698);
nor U17953 (N_17953,N_17626,N_17621);
nor U17954 (N_17954,N_17678,N_17641);
nor U17955 (N_17955,N_17621,N_17773);
and U17956 (N_17956,N_17636,N_17714);
nor U17957 (N_17957,N_17686,N_17698);
xnor U17958 (N_17958,N_17671,N_17630);
nand U17959 (N_17959,N_17644,N_17632);
and U17960 (N_17960,N_17655,N_17744);
nand U17961 (N_17961,N_17777,N_17755);
xnor U17962 (N_17962,N_17769,N_17638);
nor U17963 (N_17963,N_17617,N_17726);
and U17964 (N_17964,N_17684,N_17615);
or U17965 (N_17965,N_17715,N_17681);
and U17966 (N_17966,N_17738,N_17799);
nor U17967 (N_17967,N_17790,N_17687);
or U17968 (N_17968,N_17792,N_17783);
and U17969 (N_17969,N_17679,N_17601);
nor U17970 (N_17970,N_17791,N_17760);
xor U17971 (N_17971,N_17675,N_17726);
nor U17972 (N_17972,N_17608,N_17749);
and U17973 (N_17973,N_17774,N_17698);
and U17974 (N_17974,N_17741,N_17663);
xnor U17975 (N_17975,N_17796,N_17668);
nor U17976 (N_17976,N_17700,N_17786);
or U17977 (N_17977,N_17636,N_17606);
or U17978 (N_17978,N_17675,N_17620);
nand U17979 (N_17979,N_17629,N_17730);
or U17980 (N_17980,N_17606,N_17728);
and U17981 (N_17981,N_17653,N_17761);
nor U17982 (N_17982,N_17678,N_17787);
nor U17983 (N_17983,N_17792,N_17638);
and U17984 (N_17984,N_17790,N_17642);
and U17985 (N_17985,N_17625,N_17674);
nand U17986 (N_17986,N_17753,N_17792);
xnor U17987 (N_17987,N_17669,N_17755);
xnor U17988 (N_17988,N_17707,N_17720);
nor U17989 (N_17989,N_17714,N_17787);
nand U17990 (N_17990,N_17788,N_17702);
or U17991 (N_17991,N_17670,N_17784);
nor U17992 (N_17992,N_17678,N_17637);
and U17993 (N_17993,N_17714,N_17605);
and U17994 (N_17994,N_17649,N_17642);
or U17995 (N_17995,N_17719,N_17658);
xnor U17996 (N_17996,N_17782,N_17699);
or U17997 (N_17997,N_17791,N_17795);
or U17998 (N_17998,N_17601,N_17658);
xnor U17999 (N_17999,N_17605,N_17794);
nor U18000 (N_18000,N_17888,N_17853);
nor U18001 (N_18001,N_17873,N_17878);
nor U18002 (N_18002,N_17988,N_17854);
and U18003 (N_18003,N_17892,N_17927);
xor U18004 (N_18004,N_17964,N_17805);
nand U18005 (N_18005,N_17812,N_17863);
xnor U18006 (N_18006,N_17976,N_17852);
xor U18007 (N_18007,N_17827,N_17908);
xnor U18008 (N_18008,N_17830,N_17826);
or U18009 (N_18009,N_17929,N_17965);
xor U18010 (N_18010,N_17836,N_17921);
nor U18011 (N_18011,N_17926,N_17834);
or U18012 (N_18012,N_17981,N_17881);
and U18013 (N_18013,N_17814,N_17983);
nand U18014 (N_18014,N_17950,N_17867);
and U18015 (N_18015,N_17809,N_17932);
nor U18016 (N_18016,N_17954,N_17987);
xnor U18017 (N_18017,N_17810,N_17831);
or U18018 (N_18018,N_17840,N_17894);
or U18019 (N_18019,N_17869,N_17974);
and U18020 (N_18020,N_17984,N_17957);
nand U18021 (N_18021,N_17937,N_17913);
nand U18022 (N_18022,N_17887,N_17914);
and U18023 (N_18023,N_17821,N_17850);
and U18024 (N_18024,N_17906,N_17963);
or U18025 (N_18025,N_17872,N_17910);
nor U18026 (N_18026,N_17896,N_17962);
or U18027 (N_18027,N_17995,N_17866);
nor U18028 (N_18028,N_17855,N_17979);
or U18029 (N_18029,N_17862,N_17839);
and U18030 (N_18030,N_17816,N_17970);
and U18031 (N_18031,N_17843,N_17832);
or U18032 (N_18032,N_17898,N_17828);
nor U18033 (N_18033,N_17999,N_17930);
xnor U18034 (N_18034,N_17919,N_17980);
nand U18035 (N_18035,N_17907,N_17800);
nand U18036 (N_18036,N_17891,N_17815);
nand U18037 (N_18037,N_17938,N_17918);
nand U18038 (N_18038,N_17996,N_17939);
nand U18039 (N_18039,N_17895,N_17959);
nand U18040 (N_18040,N_17877,N_17953);
or U18041 (N_18041,N_17993,N_17817);
and U18042 (N_18042,N_17911,N_17972);
xnor U18043 (N_18043,N_17923,N_17956);
or U18044 (N_18044,N_17942,N_17917);
nand U18045 (N_18045,N_17803,N_17941);
or U18046 (N_18046,N_17811,N_17997);
nor U18047 (N_18047,N_17819,N_17856);
xor U18048 (N_18048,N_17905,N_17936);
nor U18049 (N_18049,N_17935,N_17876);
xnor U18050 (N_18050,N_17848,N_17945);
or U18051 (N_18051,N_17813,N_17902);
and U18052 (N_18052,N_17928,N_17849);
or U18053 (N_18053,N_17851,N_17880);
xor U18054 (N_18054,N_17897,N_17958);
or U18055 (N_18055,N_17870,N_17871);
nand U18056 (N_18056,N_17847,N_17801);
xor U18057 (N_18057,N_17889,N_17934);
and U18058 (N_18058,N_17944,N_17890);
xnor U18059 (N_18059,N_17885,N_17947);
nand U18060 (N_18060,N_17971,N_17882);
nor U18061 (N_18061,N_17909,N_17933);
or U18062 (N_18062,N_17808,N_17865);
xnor U18063 (N_18063,N_17904,N_17903);
xnor U18064 (N_18064,N_17899,N_17820);
nor U18065 (N_18065,N_17874,N_17994);
nand U18066 (N_18066,N_17916,N_17841);
or U18067 (N_18067,N_17859,N_17967);
nand U18068 (N_18068,N_17920,N_17824);
nor U18069 (N_18069,N_17857,N_17949);
and U18070 (N_18070,N_17802,N_17833);
and U18071 (N_18071,N_17925,N_17837);
xor U18072 (N_18072,N_17946,N_17991);
or U18073 (N_18073,N_17943,N_17931);
and U18074 (N_18074,N_17900,N_17985);
nand U18075 (N_18075,N_17924,N_17982);
nor U18076 (N_18076,N_17879,N_17845);
or U18077 (N_18077,N_17915,N_17978);
or U18078 (N_18078,N_17975,N_17977);
or U18079 (N_18079,N_17806,N_17948);
xor U18080 (N_18080,N_17823,N_17912);
xor U18081 (N_18081,N_17966,N_17940);
xor U18082 (N_18082,N_17858,N_17992);
nand U18083 (N_18083,N_17968,N_17864);
or U18084 (N_18084,N_17969,N_17893);
or U18085 (N_18085,N_17818,N_17835);
or U18086 (N_18086,N_17861,N_17838);
nand U18087 (N_18087,N_17807,N_17883);
or U18088 (N_18088,N_17842,N_17901);
nand U18089 (N_18089,N_17922,N_17955);
nand U18090 (N_18090,N_17822,N_17884);
or U18091 (N_18091,N_17844,N_17960);
nand U18092 (N_18092,N_17952,N_17829);
xor U18093 (N_18093,N_17825,N_17804);
or U18094 (N_18094,N_17951,N_17868);
nor U18095 (N_18095,N_17886,N_17986);
nand U18096 (N_18096,N_17998,N_17973);
or U18097 (N_18097,N_17961,N_17860);
xnor U18098 (N_18098,N_17990,N_17846);
xor U18099 (N_18099,N_17989,N_17875);
nor U18100 (N_18100,N_17900,N_17878);
nand U18101 (N_18101,N_17974,N_17874);
nor U18102 (N_18102,N_17949,N_17966);
nor U18103 (N_18103,N_17949,N_17874);
or U18104 (N_18104,N_17968,N_17948);
nor U18105 (N_18105,N_17862,N_17928);
or U18106 (N_18106,N_17927,N_17911);
nor U18107 (N_18107,N_17912,N_17915);
xor U18108 (N_18108,N_17877,N_17917);
nor U18109 (N_18109,N_17808,N_17871);
or U18110 (N_18110,N_17812,N_17992);
or U18111 (N_18111,N_17870,N_17944);
xnor U18112 (N_18112,N_17858,N_17883);
and U18113 (N_18113,N_17833,N_17940);
xnor U18114 (N_18114,N_17854,N_17815);
xnor U18115 (N_18115,N_17854,N_17912);
or U18116 (N_18116,N_17964,N_17992);
nor U18117 (N_18117,N_17945,N_17835);
xnor U18118 (N_18118,N_17892,N_17828);
nor U18119 (N_18119,N_17962,N_17800);
xnor U18120 (N_18120,N_17814,N_17890);
nor U18121 (N_18121,N_17866,N_17870);
or U18122 (N_18122,N_17930,N_17813);
nor U18123 (N_18123,N_17975,N_17904);
nand U18124 (N_18124,N_17848,N_17937);
and U18125 (N_18125,N_17856,N_17953);
and U18126 (N_18126,N_17946,N_17910);
nand U18127 (N_18127,N_17870,N_17911);
and U18128 (N_18128,N_17885,N_17878);
and U18129 (N_18129,N_17930,N_17960);
nand U18130 (N_18130,N_17969,N_17864);
and U18131 (N_18131,N_17903,N_17996);
nor U18132 (N_18132,N_17816,N_17835);
or U18133 (N_18133,N_17832,N_17871);
or U18134 (N_18134,N_17918,N_17852);
xnor U18135 (N_18135,N_17939,N_17995);
nand U18136 (N_18136,N_17980,N_17979);
nand U18137 (N_18137,N_17958,N_17887);
xor U18138 (N_18138,N_17911,N_17918);
nor U18139 (N_18139,N_17989,N_17990);
nor U18140 (N_18140,N_17831,N_17963);
and U18141 (N_18141,N_17888,N_17950);
or U18142 (N_18142,N_17850,N_17948);
and U18143 (N_18143,N_17958,N_17906);
xor U18144 (N_18144,N_17925,N_17820);
nand U18145 (N_18145,N_17814,N_17864);
nor U18146 (N_18146,N_17984,N_17802);
xor U18147 (N_18147,N_17996,N_17975);
nor U18148 (N_18148,N_17902,N_17808);
nor U18149 (N_18149,N_17835,N_17897);
nor U18150 (N_18150,N_17926,N_17831);
and U18151 (N_18151,N_17927,N_17966);
nand U18152 (N_18152,N_17842,N_17862);
nor U18153 (N_18153,N_17888,N_17915);
and U18154 (N_18154,N_17929,N_17838);
nand U18155 (N_18155,N_17876,N_17891);
xor U18156 (N_18156,N_17969,N_17878);
nor U18157 (N_18157,N_17964,N_17878);
nand U18158 (N_18158,N_17950,N_17858);
and U18159 (N_18159,N_17938,N_17925);
xor U18160 (N_18160,N_17902,N_17865);
and U18161 (N_18161,N_17934,N_17953);
and U18162 (N_18162,N_17820,N_17885);
or U18163 (N_18163,N_17803,N_17860);
nand U18164 (N_18164,N_17869,N_17859);
nand U18165 (N_18165,N_17862,N_17906);
and U18166 (N_18166,N_17891,N_17803);
and U18167 (N_18167,N_17932,N_17958);
or U18168 (N_18168,N_17884,N_17857);
nand U18169 (N_18169,N_17950,N_17975);
or U18170 (N_18170,N_17973,N_17904);
and U18171 (N_18171,N_17800,N_17985);
and U18172 (N_18172,N_17921,N_17801);
xor U18173 (N_18173,N_17961,N_17979);
and U18174 (N_18174,N_17849,N_17865);
or U18175 (N_18175,N_17968,N_17852);
xnor U18176 (N_18176,N_17888,N_17941);
and U18177 (N_18177,N_17845,N_17909);
nand U18178 (N_18178,N_17995,N_17914);
nor U18179 (N_18179,N_17804,N_17987);
and U18180 (N_18180,N_17872,N_17964);
xnor U18181 (N_18181,N_17844,N_17808);
and U18182 (N_18182,N_17934,N_17993);
nand U18183 (N_18183,N_17880,N_17986);
and U18184 (N_18184,N_17988,N_17842);
nand U18185 (N_18185,N_17861,N_17915);
and U18186 (N_18186,N_17838,N_17924);
nand U18187 (N_18187,N_17878,N_17973);
nand U18188 (N_18188,N_17873,N_17828);
or U18189 (N_18189,N_17817,N_17855);
and U18190 (N_18190,N_17959,N_17828);
or U18191 (N_18191,N_17923,N_17834);
and U18192 (N_18192,N_17864,N_17822);
or U18193 (N_18193,N_17862,N_17856);
and U18194 (N_18194,N_17899,N_17827);
or U18195 (N_18195,N_17993,N_17923);
nor U18196 (N_18196,N_17952,N_17809);
xnor U18197 (N_18197,N_17999,N_17929);
nand U18198 (N_18198,N_17916,N_17991);
or U18199 (N_18199,N_17954,N_17991);
nand U18200 (N_18200,N_18013,N_18111);
and U18201 (N_18201,N_18156,N_18099);
and U18202 (N_18202,N_18195,N_18078);
xnor U18203 (N_18203,N_18105,N_18198);
or U18204 (N_18204,N_18102,N_18016);
nor U18205 (N_18205,N_18171,N_18147);
and U18206 (N_18206,N_18154,N_18043);
or U18207 (N_18207,N_18123,N_18030);
nand U18208 (N_18208,N_18057,N_18139);
or U18209 (N_18209,N_18100,N_18091);
or U18210 (N_18210,N_18064,N_18117);
xnor U18211 (N_18211,N_18025,N_18132);
xor U18212 (N_18212,N_18088,N_18039);
nor U18213 (N_18213,N_18143,N_18140);
nor U18214 (N_18214,N_18017,N_18131);
xnor U18215 (N_18215,N_18138,N_18197);
nand U18216 (N_18216,N_18062,N_18001);
xnor U18217 (N_18217,N_18021,N_18187);
nand U18218 (N_18218,N_18049,N_18061);
or U18219 (N_18219,N_18066,N_18141);
and U18220 (N_18220,N_18028,N_18050);
nand U18221 (N_18221,N_18087,N_18189);
nand U18222 (N_18222,N_18127,N_18182);
nand U18223 (N_18223,N_18083,N_18038);
nand U18224 (N_18224,N_18056,N_18145);
or U18225 (N_18225,N_18177,N_18137);
xnor U18226 (N_18226,N_18014,N_18086);
xor U18227 (N_18227,N_18065,N_18183);
xor U18228 (N_18228,N_18047,N_18175);
or U18229 (N_18229,N_18036,N_18018);
nand U18230 (N_18230,N_18090,N_18045);
and U18231 (N_18231,N_18020,N_18008);
nor U18232 (N_18232,N_18063,N_18075);
xnor U18233 (N_18233,N_18181,N_18134);
or U18234 (N_18234,N_18098,N_18160);
nand U18235 (N_18235,N_18034,N_18186);
xor U18236 (N_18236,N_18178,N_18084);
or U18237 (N_18237,N_18000,N_18104);
xor U18238 (N_18238,N_18003,N_18113);
and U18239 (N_18239,N_18068,N_18071);
nand U18240 (N_18240,N_18172,N_18110);
and U18241 (N_18241,N_18081,N_18136);
xnor U18242 (N_18242,N_18094,N_18184);
xnor U18243 (N_18243,N_18118,N_18115);
nor U18244 (N_18244,N_18085,N_18158);
or U18245 (N_18245,N_18126,N_18193);
xnor U18246 (N_18246,N_18167,N_18133);
or U18247 (N_18247,N_18159,N_18048);
nor U18248 (N_18248,N_18191,N_18109);
and U18249 (N_18249,N_18031,N_18112);
xor U18250 (N_18250,N_18157,N_18180);
and U18251 (N_18251,N_18149,N_18166);
nor U18252 (N_18252,N_18174,N_18176);
or U18253 (N_18253,N_18169,N_18027);
and U18254 (N_18254,N_18097,N_18029);
xnor U18255 (N_18255,N_18161,N_18080);
nand U18256 (N_18256,N_18116,N_18070);
xor U18257 (N_18257,N_18032,N_18054);
xnor U18258 (N_18258,N_18144,N_18192);
xor U18259 (N_18259,N_18199,N_18124);
xor U18260 (N_18260,N_18120,N_18101);
and U18261 (N_18261,N_18194,N_18188);
and U18262 (N_18262,N_18055,N_18072);
and U18263 (N_18263,N_18009,N_18150);
or U18264 (N_18264,N_18173,N_18058);
or U18265 (N_18265,N_18073,N_18135);
nor U18266 (N_18266,N_18023,N_18155);
and U18267 (N_18267,N_18067,N_18095);
nor U18268 (N_18268,N_18106,N_18096);
and U18269 (N_18269,N_18046,N_18015);
nand U18270 (N_18270,N_18128,N_18179);
nor U18271 (N_18271,N_18185,N_18146);
nand U18272 (N_18272,N_18004,N_18060);
xnor U18273 (N_18273,N_18165,N_18044);
nor U18274 (N_18274,N_18130,N_18006);
and U18275 (N_18275,N_18122,N_18026);
nand U18276 (N_18276,N_18079,N_18162);
nor U18277 (N_18277,N_18024,N_18074);
and U18278 (N_18278,N_18196,N_18107);
or U18279 (N_18279,N_18119,N_18168);
nor U18280 (N_18280,N_18033,N_18190);
nor U18281 (N_18281,N_18129,N_18163);
and U18282 (N_18282,N_18069,N_18164);
xnor U18283 (N_18283,N_18037,N_18153);
or U18284 (N_18284,N_18053,N_18042);
and U18285 (N_18285,N_18092,N_18082);
nor U18286 (N_18286,N_18035,N_18148);
and U18287 (N_18287,N_18052,N_18010);
xor U18288 (N_18288,N_18114,N_18002);
xnor U18289 (N_18289,N_18103,N_18151);
xor U18290 (N_18290,N_18059,N_18121);
and U18291 (N_18291,N_18019,N_18125);
and U18292 (N_18292,N_18040,N_18051);
xor U18293 (N_18293,N_18152,N_18012);
nor U18294 (N_18294,N_18093,N_18089);
and U18295 (N_18295,N_18007,N_18041);
xnor U18296 (N_18296,N_18170,N_18022);
and U18297 (N_18297,N_18108,N_18077);
and U18298 (N_18298,N_18005,N_18011);
xnor U18299 (N_18299,N_18076,N_18142);
and U18300 (N_18300,N_18097,N_18108);
and U18301 (N_18301,N_18164,N_18081);
nand U18302 (N_18302,N_18046,N_18074);
nor U18303 (N_18303,N_18105,N_18065);
nand U18304 (N_18304,N_18021,N_18008);
or U18305 (N_18305,N_18062,N_18187);
nand U18306 (N_18306,N_18175,N_18130);
nand U18307 (N_18307,N_18166,N_18191);
xor U18308 (N_18308,N_18172,N_18038);
nor U18309 (N_18309,N_18102,N_18173);
nor U18310 (N_18310,N_18107,N_18190);
and U18311 (N_18311,N_18043,N_18082);
nand U18312 (N_18312,N_18090,N_18006);
nand U18313 (N_18313,N_18045,N_18195);
or U18314 (N_18314,N_18050,N_18026);
and U18315 (N_18315,N_18196,N_18189);
or U18316 (N_18316,N_18173,N_18198);
nor U18317 (N_18317,N_18075,N_18080);
nor U18318 (N_18318,N_18047,N_18187);
and U18319 (N_18319,N_18061,N_18147);
nor U18320 (N_18320,N_18024,N_18002);
xor U18321 (N_18321,N_18117,N_18032);
xnor U18322 (N_18322,N_18133,N_18009);
nand U18323 (N_18323,N_18156,N_18018);
and U18324 (N_18324,N_18189,N_18019);
and U18325 (N_18325,N_18163,N_18165);
xnor U18326 (N_18326,N_18077,N_18192);
nor U18327 (N_18327,N_18108,N_18153);
and U18328 (N_18328,N_18139,N_18155);
nand U18329 (N_18329,N_18186,N_18113);
and U18330 (N_18330,N_18129,N_18161);
nand U18331 (N_18331,N_18046,N_18064);
nand U18332 (N_18332,N_18171,N_18046);
or U18333 (N_18333,N_18015,N_18107);
and U18334 (N_18334,N_18070,N_18127);
or U18335 (N_18335,N_18168,N_18005);
nor U18336 (N_18336,N_18047,N_18143);
or U18337 (N_18337,N_18194,N_18124);
xor U18338 (N_18338,N_18055,N_18075);
or U18339 (N_18339,N_18023,N_18033);
xor U18340 (N_18340,N_18194,N_18060);
and U18341 (N_18341,N_18081,N_18019);
xnor U18342 (N_18342,N_18145,N_18159);
nor U18343 (N_18343,N_18148,N_18030);
nand U18344 (N_18344,N_18072,N_18014);
nand U18345 (N_18345,N_18117,N_18118);
nor U18346 (N_18346,N_18109,N_18179);
xor U18347 (N_18347,N_18193,N_18146);
xnor U18348 (N_18348,N_18100,N_18151);
xnor U18349 (N_18349,N_18122,N_18197);
and U18350 (N_18350,N_18192,N_18101);
xnor U18351 (N_18351,N_18014,N_18153);
and U18352 (N_18352,N_18098,N_18152);
nor U18353 (N_18353,N_18088,N_18147);
nand U18354 (N_18354,N_18077,N_18025);
or U18355 (N_18355,N_18129,N_18027);
and U18356 (N_18356,N_18038,N_18169);
nor U18357 (N_18357,N_18053,N_18050);
xor U18358 (N_18358,N_18015,N_18059);
xnor U18359 (N_18359,N_18193,N_18078);
xnor U18360 (N_18360,N_18145,N_18177);
nand U18361 (N_18361,N_18060,N_18093);
or U18362 (N_18362,N_18193,N_18127);
xnor U18363 (N_18363,N_18081,N_18055);
and U18364 (N_18364,N_18100,N_18165);
or U18365 (N_18365,N_18176,N_18055);
xnor U18366 (N_18366,N_18160,N_18157);
nand U18367 (N_18367,N_18178,N_18159);
nor U18368 (N_18368,N_18128,N_18065);
nand U18369 (N_18369,N_18118,N_18030);
and U18370 (N_18370,N_18050,N_18045);
nand U18371 (N_18371,N_18121,N_18067);
xor U18372 (N_18372,N_18169,N_18051);
and U18373 (N_18373,N_18043,N_18114);
and U18374 (N_18374,N_18003,N_18029);
nand U18375 (N_18375,N_18040,N_18190);
nand U18376 (N_18376,N_18159,N_18064);
or U18377 (N_18377,N_18143,N_18104);
or U18378 (N_18378,N_18169,N_18072);
or U18379 (N_18379,N_18036,N_18115);
or U18380 (N_18380,N_18106,N_18017);
and U18381 (N_18381,N_18040,N_18034);
or U18382 (N_18382,N_18133,N_18057);
and U18383 (N_18383,N_18001,N_18154);
or U18384 (N_18384,N_18060,N_18197);
nand U18385 (N_18385,N_18164,N_18167);
nand U18386 (N_18386,N_18134,N_18074);
or U18387 (N_18387,N_18007,N_18016);
nor U18388 (N_18388,N_18158,N_18082);
and U18389 (N_18389,N_18131,N_18068);
nand U18390 (N_18390,N_18125,N_18085);
nand U18391 (N_18391,N_18121,N_18076);
nand U18392 (N_18392,N_18111,N_18014);
nand U18393 (N_18393,N_18002,N_18068);
or U18394 (N_18394,N_18016,N_18108);
and U18395 (N_18395,N_18099,N_18032);
or U18396 (N_18396,N_18049,N_18000);
and U18397 (N_18397,N_18121,N_18084);
or U18398 (N_18398,N_18001,N_18092);
nand U18399 (N_18399,N_18020,N_18119);
nor U18400 (N_18400,N_18237,N_18231);
xnor U18401 (N_18401,N_18239,N_18264);
nand U18402 (N_18402,N_18394,N_18391);
nand U18403 (N_18403,N_18277,N_18349);
nor U18404 (N_18404,N_18355,N_18281);
nor U18405 (N_18405,N_18322,N_18221);
nor U18406 (N_18406,N_18293,N_18360);
nor U18407 (N_18407,N_18223,N_18262);
nand U18408 (N_18408,N_18256,N_18213);
nand U18409 (N_18409,N_18362,N_18284);
and U18410 (N_18410,N_18308,N_18326);
nand U18411 (N_18411,N_18300,N_18319);
nand U18412 (N_18412,N_18283,N_18383);
nor U18413 (N_18413,N_18229,N_18333);
nor U18414 (N_18414,N_18358,N_18218);
or U18415 (N_18415,N_18343,N_18235);
xnor U18416 (N_18416,N_18219,N_18357);
and U18417 (N_18417,N_18305,N_18296);
xor U18418 (N_18418,N_18201,N_18271);
or U18419 (N_18419,N_18253,N_18205);
nand U18420 (N_18420,N_18382,N_18311);
nor U18421 (N_18421,N_18268,N_18246);
xnor U18422 (N_18422,N_18209,N_18393);
nor U18423 (N_18423,N_18352,N_18368);
xnor U18424 (N_18424,N_18377,N_18230);
and U18425 (N_18425,N_18367,N_18238);
xor U18426 (N_18426,N_18353,N_18243);
and U18427 (N_18427,N_18233,N_18265);
nor U18428 (N_18428,N_18370,N_18299);
xor U18429 (N_18429,N_18346,N_18335);
nand U18430 (N_18430,N_18347,N_18303);
xnor U18431 (N_18431,N_18388,N_18228);
nand U18432 (N_18432,N_18312,N_18385);
or U18433 (N_18433,N_18325,N_18316);
nand U18434 (N_18434,N_18376,N_18288);
and U18435 (N_18435,N_18345,N_18395);
xor U18436 (N_18436,N_18216,N_18236);
xnor U18437 (N_18437,N_18240,N_18204);
xor U18438 (N_18438,N_18329,N_18287);
nor U18439 (N_18439,N_18289,N_18356);
nor U18440 (N_18440,N_18298,N_18371);
nand U18441 (N_18441,N_18290,N_18307);
xor U18442 (N_18442,N_18399,N_18211);
nand U18443 (N_18443,N_18252,N_18304);
or U18444 (N_18444,N_18279,N_18226);
nand U18445 (N_18445,N_18320,N_18274);
or U18446 (N_18446,N_18285,N_18351);
xor U18447 (N_18447,N_18222,N_18203);
or U18448 (N_18448,N_18234,N_18280);
xnor U18449 (N_18449,N_18380,N_18255);
or U18450 (N_18450,N_18270,N_18225);
or U18451 (N_18451,N_18373,N_18224);
nor U18452 (N_18452,N_18344,N_18328);
xor U18453 (N_18453,N_18334,N_18369);
xnor U18454 (N_18454,N_18331,N_18310);
nor U18455 (N_18455,N_18286,N_18241);
nor U18456 (N_18456,N_18242,N_18327);
nor U18457 (N_18457,N_18206,N_18227);
or U18458 (N_18458,N_18390,N_18260);
or U18459 (N_18459,N_18378,N_18337);
or U18460 (N_18460,N_18323,N_18294);
nor U18461 (N_18461,N_18245,N_18215);
nand U18462 (N_18462,N_18220,N_18263);
or U18463 (N_18463,N_18292,N_18217);
nand U18464 (N_18464,N_18254,N_18324);
nor U18465 (N_18465,N_18363,N_18365);
nand U18466 (N_18466,N_18361,N_18295);
or U18467 (N_18467,N_18297,N_18374);
nand U18468 (N_18468,N_18272,N_18381);
or U18469 (N_18469,N_18318,N_18384);
or U18470 (N_18470,N_18302,N_18207);
and U18471 (N_18471,N_18250,N_18332);
and U18472 (N_18472,N_18232,N_18269);
nor U18473 (N_18473,N_18266,N_18366);
xor U18474 (N_18474,N_18359,N_18372);
and U18475 (N_18475,N_18282,N_18336);
and U18476 (N_18476,N_18214,N_18330);
xnor U18477 (N_18477,N_18202,N_18314);
nand U18478 (N_18478,N_18387,N_18200);
nand U18479 (N_18479,N_18348,N_18317);
xor U18480 (N_18480,N_18244,N_18212);
xor U18481 (N_18481,N_18210,N_18321);
and U18482 (N_18482,N_18340,N_18309);
nand U18483 (N_18483,N_18278,N_18276);
and U18484 (N_18484,N_18291,N_18398);
nand U18485 (N_18485,N_18386,N_18261);
xor U18486 (N_18486,N_18257,N_18364);
or U18487 (N_18487,N_18350,N_18259);
or U18488 (N_18488,N_18392,N_18273);
nand U18489 (N_18489,N_18267,N_18249);
or U18490 (N_18490,N_18301,N_18354);
xnor U18491 (N_18491,N_18251,N_18315);
nor U18492 (N_18492,N_18258,N_18397);
or U18493 (N_18493,N_18375,N_18306);
nand U18494 (N_18494,N_18339,N_18208);
nor U18495 (N_18495,N_18313,N_18248);
nand U18496 (N_18496,N_18379,N_18275);
and U18497 (N_18497,N_18338,N_18341);
xor U18498 (N_18498,N_18247,N_18342);
xor U18499 (N_18499,N_18396,N_18389);
nor U18500 (N_18500,N_18370,N_18358);
nand U18501 (N_18501,N_18200,N_18215);
or U18502 (N_18502,N_18203,N_18340);
and U18503 (N_18503,N_18229,N_18306);
nor U18504 (N_18504,N_18322,N_18315);
nor U18505 (N_18505,N_18382,N_18305);
or U18506 (N_18506,N_18239,N_18289);
and U18507 (N_18507,N_18202,N_18389);
and U18508 (N_18508,N_18398,N_18371);
or U18509 (N_18509,N_18235,N_18387);
and U18510 (N_18510,N_18257,N_18242);
nand U18511 (N_18511,N_18273,N_18237);
xor U18512 (N_18512,N_18215,N_18391);
nand U18513 (N_18513,N_18366,N_18209);
or U18514 (N_18514,N_18253,N_18281);
xnor U18515 (N_18515,N_18361,N_18377);
and U18516 (N_18516,N_18311,N_18203);
nor U18517 (N_18517,N_18397,N_18309);
or U18518 (N_18518,N_18389,N_18347);
or U18519 (N_18519,N_18391,N_18225);
nand U18520 (N_18520,N_18368,N_18210);
xnor U18521 (N_18521,N_18375,N_18300);
nor U18522 (N_18522,N_18312,N_18307);
nor U18523 (N_18523,N_18394,N_18281);
or U18524 (N_18524,N_18235,N_18388);
nor U18525 (N_18525,N_18215,N_18322);
nand U18526 (N_18526,N_18339,N_18364);
xor U18527 (N_18527,N_18334,N_18397);
nor U18528 (N_18528,N_18369,N_18306);
or U18529 (N_18529,N_18321,N_18251);
nand U18530 (N_18530,N_18216,N_18246);
xor U18531 (N_18531,N_18220,N_18360);
or U18532 (N_18532,N_18311,N_18234);
xor U18533 (N_18533,N_18264,N_18257);
nor U18534 (N_18534,N_18291,N_18339);
nor U18535 (N_18535,N_18353,N_18302);
or U18536 (N_18536,N_18249,N_18203);
nor U18537 (N_18537,N_18372,N_18373);
xnor U18538 (N_18538,N_18293,N_18255);
nor U18539 (N_18539,N_18274,N_18292);
nor U18540 (N_18540,N_18261,N_18293);
and U18541 (N_18541,N_18219,N_18267);
or U18542 (N_18542,N_18223,N_18315);
nand U18543 (N_18543,N_18395,N_18324);
and U18544 (N_18544,N_18214,N_18254);
or U18545 (N_18545,N_18395,N_18367);
nor U18546 (N_18546,N_18327,N_18260);
and U18547 (N_18547,N_18292,N_18375);
nor U18548 (N_18548,N_18381,N_18334);
and U18549 (N_18549,N_18374,N_18244);
nor U18550 (N_18550,N_18282,N_18393);
and U18551 (N_18551,N_18229,N_18384);
or U18552 (N_18552,N_18304,N_18262);
and U18553 (N_18553,N_18287,N_18367);
nor U18554 (N_18554,N_18266,N_18394);
xor U18555 (N_18555,N_18241,N_18214);
and U18556 (N_18556,N_18357,N_18337);
nand U18557 (N_18557,N_18320,N_18270);
xor U18558 (N_18558,N_18392,N_18251);
nor U18559 (N_18559,N_18331,N_18211);
or U18560 (N_18560,N_18351,N_18291);
and U18561 (N_18561,N_18360,N_18316);
or U18562 (N_18562,N_18253,N_18369);
or U18563 (N_18563,N_18361,N_18391);
xnor U18564 (N_18564,N_18320,N_18245);
and U18565 (N_18565,N_18262,N_18328);
and U18566 (N_18566,N_18284,N_18371);
and U18567 (N_18567,N_18309,N_18359);
and U18568 (N_18568,N_18346,N_18317);
and U18569 (N_18569,N_18318,N_18237);
and U18570 (N_18570,N_18202,N_18265);
nand U18571 (N_18571,N_18367,N_18340);
and U18572 (N_18572,N_18356,N_18205);
xor U18573 (N_18573,N_18307,N_18211);
nor U18574 (N_18574,N_18228,N_18345);
xor U18575 (N_18575,N_18309,N_18322);
xnor U18576 (N_18576,N_18364,N_18399);
and U18577 (N_18577,N_18233,N_18348);
or U18578 (N_18578,N_18285,N_18256);
nand U18579 (N_18579,N_18240,N_18290);
nand U18580 (N_18580,N_18362,N_18248);
nor U18581 (N_18581,N_18284,N_18367);
or U18582 (N_18582,N_18219,N_18221);
and U18583 (N_18583,N_18301,N_18389);
or U18584 (N_18584,N_18395,N_18387);
xnor U18585 (N_18585,N_18370,N_18364);
nand U18586 (N_18586,N_18273,N_18309);
and U18587 (N_18587,N_18279,N_18351);
or U18588 (N_18588,N_18301,N_18336);
and U18589 (N_18589,N_18333,N_18381);
xnor U18590 (N_18590,N_18338,N_18240);
nor U18591 (N_18591,N_18330,N_18353);
nand U18592 (N_18592,N_18310,N_18267);
xnor U18593 (N_18593,N_18208,N_18334);
and U18594 (N_18594,N_18332,N_18218);
nor U18595 (N_18595,N_18387,N_18295);
xor U18596 (N_18596,N_18226,N_18219);
xnor U18597 (N_18597,N_18389,N_18392);
xnor U18598 (N_18598,N_18379,N_18283);
or U18599 (N_18599,N_18309,N_18278);
or U18600 (N_18600,N_18447,N_18511);
nor U18601 (N_18601,N_18505,N_18545);
nor U18602 (N_18602,N_18406,N_18509);
xnor U18603 (N_18603,N_18476,N_18413);
xnor U18604 (N_18604,N_18484,N_18566);
nand U18605 (N_18605,N_18424,N_18423);
nand U18606 (N_18606,N_18588,N_18530);
nand U18607 (N_18607,N_18575,N_18448);
nor U18608 (N_18608,N_18453,N_18458);
or U18609 (N_18609,N_18435,N_18425);
xnor U18610 (N_18610,N_18446,N_18443);
nand U18611 (N_18611,N_18433,N_18570);
xnor U18612 (N_18612,N_18401,N_18591);
xnor U18613 (N_18613,N_18494,N_18547);
xnor U18614 (N_18614,N_18518,N_18539);
nand U18615 (N_18615,N_18506,N_18421);
nand U18616 (N_18616,N_18531,N_18422);
nor U18617 (N_18617,N_18479,N_18498);
nor U18618 (N_18618,N_18553,N_18542);
xnor U18619 (N_18619,N_18420,N_18578);
nor U18620 (N_18620,N_18429,N_18525);
nand U18621 (N_18621,N_18457,N_18538);
and U18622 (N_18622,N_18452,N_18430);
or U18623 (N_18623,N_18580,N_18596);
xor U18624 (N_18624,N_18400,N_18587);
nand U18625 (N_18625,N_18559,N_18486);
xnor U18626 (N_18626,N_18541,N_18502);
and U18627 (N_18627,N_18589,N_18516);
nor U18628 (N_18628,N_18440,N_18480);
or U18629 (N_18629,N_18515,N_18426);
and U18630 (N_18630,N_18455,N_18584);
or U18631 (N_18631,N_18472,N_18565);
xor U18632 (N_18632,N_18546,N_18599);
or U18633 (N_18633,N_18558,N_18490);
xnor U18634 (N_18634,N_18464,N_18454);
and U18635 (N_18635,N_18532,N_18534);
xnor U18636 (N_18636,N_18549,N_18543);
nor U18637 (N_18637,N_18590,N_18417);
nor U18638 (N_18638,N_18436,N_18451);
xor U18639 (N_18639,N_18507,N_18465);
nor U18640 (N_18640,N_18571,N_18548);
xor U18641 (N_18641,N_18520,N_18526);
nor U18642 (N_18642,N_18499,N_18551);
or U18643 (N_18643,N_18597,N_18527);
xnor U18644 (N_18644,N_18483,N_18434);
nand U18645 (N_18645,N_18510,N_18556);
nand U18646 (N_18646,N_18528,N_18439);
xor U18647 (N_18647,N_18475,N_18474);
nand U18648 (N_18648,N_18459,N_18462);
and U18649 (N_18649,N_18467,N_18415);
xor U18650 (N_18650,N_18573,N_18592);
and U18651 (N_18651,N_18557,N_18550);
and U18652 (N_18652,N_18432,N_18470);
nor U18653 (N_18653,N_18536,N_18410);
or U18654 (N_18654,N_18405,N_18561);
nand U18655 (N_18655,N_18529,N_18402);
xnor U18656 (N_18656,N_18574,N_18572);
or U18657 (N_18657,N_18593,N_18552);
or U18658 (N_18658,N_18576,N_18524);
or U18659 (N_18659,N_18504,N_18427);
xnor U18660 (N_18660,N_18523,N_18428);
and U18661 (N_18661,N_18404,N_18583);
or U18662 (N_18662,N_18469,N_18412);
nand U18663 (N_18663,N_18477,N_18514);
xnor U18664 (N_18664,N_18537,N_18585);
xnor U18665 (N_18665,N_18568,N_18560);
nor U18666 (N_18666,N_18416,N_18577);
and U18667 (N_18667,N_18460,N_18468);
nor U18668 (N_18668,N_18473,N_18437);
or U18669 (N_18669,N_18438,N_18533);
nor U18670 (N_18670,N_18579,N_18567);
or U18671 (N_18671,N_18522,N_18450);
nor U18672 (N_18672,N_18488,N_18595);
xnor U18673 (N_18673,N_18419,N_18493);
or U18674 (N_18674,N_18471,N_18508);
and U18675 (N_18675,N_18540,N_18408);
xnor U18676 (N_18676,N_18482,N_18594);
nor U18677 (N_18677,N_18418,N_18555);
xor U18678 (N_18678,N_18466,N_18513);
nand U18679 (N_18679,N_18562,N_18487);
or U18680 (N_18680,N_18569,N_18444);
and U18681 (N_18681,N_18461,N_18449);
and U18682 (N_18682,N_18586,N_18500);
and U18683 (N_18683,N_18582,N_18503);
xnor U18684 (N_18684,N_18492,N_18414);
xnor U18685 (N_18685,N_18544,N_18598);
and U18686 (N_18686,N_18512,N_18564);
and U18687 (N_18687,N_18491,N_18485);
nor U18688 (N_18688,N_18407,N_18501);
or U18689 (N_18689,N_18496,N_18519);
and U18690 (N_18690,N_18442,N_18554);
and U18691 (N_18691,N_18517,N_18456);
xnor U18692 (N_18692,N_18411,N_18481);
nor U18693 (N_18693,N_18495,N_18445);
nor U18694 (N_18694,N_18441,N_18489);
xnor U18695 (N_18695,N_18497,N_18563);
or U18696 (N_18696,N_18463,N_18478);
nand U18697 (N_18697,N_18431,N_18581);
and U18698 (N_18698,N_18521,N_18409);
and U18699 (N_18699,N_18535,N_18403);
nor U18700 (N_18700,N_18533,N_18512);
nand U18701 (N_18701,N_18527,N_18461);
nor U18702 (N_18702,N_18486,N_18558);
nor U18703 (N_18703,N_18592,N_18404);
nand U18704 (N_18704,N_18416,N_18531);
nor U18705 (N_18705,N_18586,N_18599);
nand U18706 (N_18706,N_18545,N_18523);
nand U18707 (N_18707,N_18475,N_18564);
nor U18708 (N_18708,N_18414,N_18575);
and U18709 (N_18709,N_18500,N_18584);
nor U18710 (N_18710,N_18437,N_18495);
and U18711 (N_18711,N_18512,N_18547);
nor U18712 (N_18712,N_18561,N_18594);
and U18713 (N_18713,N_18409,N_18439);
nor U18714 (N_18714,N_18572,N_18454);
nor U18715 (N_18715,N_18579,N_18583);
or U18716 (N_18716,N_18439,N_18561);
and U18717 (N_18717,N_18549,N_18522);
xor U18718 (N_18718,N_18421,N_18502);
and U18719 (N_18719,N_18459,N_18431);
and U18720 (N_18720,N_18527,N_18443);
and U18721 (N_18721,N_18571,N_18404);
xor U18722 (N_18722,N_18582,N_18562);
nand U18723 (N_18723,N_18505,N_18564);
nand U18724 (N_18724,N_18438,N_18580);
nor U18725 (N_18725,N_18456,N_18406);
nor U18726 (N_18726,N_18515,N_18525);
and U18727 (N_18727,N_18428,N_18404);
xor U18728 (N_18728,N_18400,N_18466);
nor U18729 (N_18729,N_18427,N_18590);
or U18730 (N_18730,N_18505,N_18401);
and U18731 (N_18731,N_18423,N_18414);
nor U18732 (N_18732,N_18492,N_18583);
and U18733 (N_18733,N_18455,N_18483);
nor U18734 (N_18734,N_18489,N_18515);
and U18735 (N_18735,N_18473,N_18555);
nand U18736 (N_18736,N_18565,N_18406);
xor U18737 (N_18737,N_18463,N_18526);
xor U18738 (N_18738,N_18584,N_18597);
or U18739 (N_18739,N_18483,N_18467);
and U18740 (N_18740,N_18410,N_18455);
nor U18741 (N_18741,N_18511,N_18555);
and U18742 (N_18742,N_18500,N_18591);
or U18743 (N_18743,N_18428,N_18579);
or U18744 (N_18744,N_18501,N_18505);
nand U18745 (N_18745,N_18541,N_18589);
xor U18746 (N_18746,N_18560,N_18472);
and U18747 (N_18747,N_18443,N_18529);
xnor U18748 (N_18748,N_18595,N_18480);
and U18749 (N_18749,N_18447,N_18419);
nor U18750 (N_18750,N_18577,N_18434);
xnor U18751 (N_18751,N_18450,N_18527);
nor U18752 (N_18752,N_18478,N_18487);
or U18753 (N_18753,N_18584,N_18518);
nor U18754 (N_18754,N_18443,N_18500);
or U18755 (N_18755,N_18407,N_18485);
and U18756 (N_18756,N_18433,N_18417);
and U18757 (N_18757,N_18497,N_18561);
nand U18758 (N_18758,N_18515,N_18484);
or U18759 (N_18759,N_18574,N_18536);
xnor U18760 (N_18760,N_18578,N_18539);
nor U18761 (N_18761,N_18514,N_18447);
xor U18762 (N_18762,N_18502,N_18519);
nand U18763 (N_18763,N_18495,N_18514);
and U18764 (N_18764,N_18514,N_18435);
nor U18765 (N_18765,N_18421,N_18514);
nor U18766 (N_18766,N_18501,N_18427);
or U18767 (N_18767,N_18549,N_18557);
or U18768 (N_18768,N_18567,N_18547);
xnor U18769 (N_18769,N_18577,N_18470);
xnor U18770 (N_18770,N_18574,N_18556);
and U18771 (N_18771,N_18590,N_18459);
or U18772 (N_18772,N_18565,N_18588);
nand U18773 (N_18773,N_18443,N_18576);
xor U18774 (N_18774,N_18512,N_18408);
xnor U18775 (N_18775,N_18533,N_18457);
or U18776 (N_18776,N_18589,N_18447);
or U18777 (N_18777,N_18595,N_18560);
xnor U18778 (N_18778,N_18412,N_18403);
and U18779 (N_18779,N_18539,N_18423);
xnor U18780 (N_18780,N_18485,N_18575);
nand U18781 (N_18781,N_18410,N_18522);
nor U18782 (N_18782,N_18555,N_18421);
xnor U18783 (N_18783,N_18511,N_18475);
xnor U18784 (N_18784,N_18497,N_18597);
nand U18785 (N_18785,N_18446,N_18536);
or U18786 (N_18786,N_18419,N_18428);
nor U18787 (N_18787,N_18572,N_18583);
nand U18788 (N_18788,N_18567,N_18406);
xor U18789 (N_18789,N_18456,N_18440);
and U18790 (N_18790,N_18453,N_18566);
nor U18791 (N_18791,N_18541,N_18574);
and U18792 (N_18792,N_18424,N_18586);
nand U18793 (N_18793,N_18501,N_18445);
or U18794 (N_18794,N_18546,N_18425);
nand U18795 (N_18795,N_18518,N_18427);
nor U18796 (N_18796,N_18592,N_18502);
xnor U18797 (N_18797,N_18412,N_18440);
nand U18798 (N_18798,N_18593,N_18465);
nor U18799 (N_18799,N_18559,N_18592);
and U18800 (N_18800,N_18791,N_18780);
or U18801 (N_18801,N_18715,N_18743);
nor U18802 (N_18802,N_18720,N_18699);
or U18803 (N_18803,N_18733,N_18796);
nor U18804 (N_18804,N_18654,N_18724);
nand U18805 (N_18805,N_18760,N_18615);
and U18806 (N_18806,N_18783,N_18766);
nand U18807 (N_18807,N_18757,N_18711);
xnor U18808 (N_18808,N_18764,N_18647);
and U18809 (N_18809,N_18799,N_18776);
nand U18810 (N_18810,N_18605,N_18696);
nand U18811 (N_18811,N_18701,N_18621);
xor U18812 (N_18812,N_18606,N_18744);
or U18813 (N_18813,N_18629,N_18669);
and U18814 (N_18814,N_18792,N_18727);
nand U18815 (N_18815,N_18738,N_18681);
nor U18816 (N_18816,N_18616,N_18667);
and U18817 (N_18817,N_18765,N_18666);
nor U18818 (N_18818,N_18725,N_18748);
or U18819 (N_18819,N_18772,N_18702);
or U18820 (N_18820,N_18689,N_18630);
xnor U18821 (N_18821,N_18678,N_18710);
and U18822 (N_18822,N_18661,N_18688);
nor U18823 (N_18823,N_18745,N_18742);
or U18824 (N_18824,N_18665,N_18610);
nor U18825 (N_18825,N_18603,N_18693);
nor U18826 (N_18826,N_18761,N_18750);
and U18827 (N_18827,N_18718,N_18746);
nand U18828 (N_18828,N_18769,N_18713);
or U18829 (N_18829,N_18762,N_18653);
nand U18830 (N_18830,N_18676,N_18614);
xor U18831 (N_18831,N_18698,N_18790);
nor U18832 (N_18832,N_18708,N_18719);
or U18833 (N_18833,N_18721,N_18753);
and U18834 (N_18834,N_18684,N_18623);
nor U18835 (N_18835,N_18691,N_18779);
nor U18836 (N_18836,N_18728,N_18797);
xnor U18837 (N_18837,N_18655,N_18798);
nand U18838 (N_18838,N_18700,N_18604);
or U18839 (N_18839,N_18767,N_18634);
xor U18840 (N_18840,N_18686,N_18709);
and U18841 (N_18841,N_18652,N_18638);
and U18842 (N_18842,N_18730,N_18671);
nor U18843 (N_18843,N_18751,N_18775);
or U18844 (N_18844,N_18703,N_18754);
or U18845 (N_18845,N_18626,N_18664);
or U18846 (N_18846,N_18613,N_18777);
and U18847 (N_18847,N_18736,N_18706);
nor U18848 (N_18848,N_18619,N_18651);
nor U18849 (N_18849,N_18707,N_18646);
nand U18850 (N_18850,N_18643,N_18645);
or U18851 (N_18851,N_18697,N_18758);
nand U18852 (N_18852,N_18773,N_18795);
and U18853 (N_18853,N_18668,N_18657);
or U18854 (N_18854,N_18625,N_18732);
and U18855 (N_18855,N_18704,N_18624);
nand U18856 (N_18856,N_18726,N_18607);
xor U18857 (N_18857,N_18723,N_18692);
or U18858 (N_18858,N_18612,N_18774);
nand U18859 (N_18859,N_18714,N_18785);
nor U18860 (N_18860,N_18771,N_18722);
nand U18861 (N_18861,N_18602,N_18794);
xnor U18862 (N_18862,N_18685,N_18755);
xor U18863 (N_18863,N_18781,N_18675);
or U18864 (N_18864,N_18729,N_18737);
nand U18865 (N_18865,N_18636,N_18632);
nand U18866 (N_18866,N_18747,N_18673);
nand U18867 (N_18867,N_18768,N_18677);
nor U18868 (N_18868,N_18752,N_18735);
nor U18869 (N_18869,N_18611,N_18658);
xor U18870 (N_18870,N_18749,N_18734);
xnor U18871 (N_18871,N_18617,N_18784);
nor U18872 (N_18872,N_18694,N_18631);
and U18873 (N_18873,N_18712,N_18670);
xnor U18874 (N_18874,N_18672,N_18674);
nor U18875 (N_18875,N_18618,N_18770);
nand U18876 (N_18876,N_18648,N_18622);
xor U18877 (N_18877,N_18627,N_18789);
nand U18878 (N_18878,N_18662,N_18786);
and U18879 (N_18879,N_18608,N_18639);
xor U18880 (N_18880,N_18659,N_18650);
or U18881 (N_18881,N_18649,N_18601);
xor U18882 (N_18882,N_18628,N_18609);
nand U18883 (N_18883,N_18782,N_18687);
nand U18884 (N_18884,N_18683,N_18716);
nand U18885 (N_18885,N_18787,N_18778);
nand U18886 (N_18886,N_18637,N_18680);
nand U18887 (N_18887,N_18640,N_18690);
xnor U18888 (N_18888,N_18756,N_18642);
nor U18889 (N_18889,N_18644,N_18656);
or U18890 (N_18890,N_18759,N_18641);
nor U18891 (N_18891,N_18740,N_18679);
xor U18892 (N_18892,N_18763,N_18705);
nor U18893 (N_18893,N_18793,N_18633);
and U18894 (N_18894,N_18741,N_18600);
nand U18895 (N_18895,N_18695,N_18788);
and U18896 (N_18896,N_18663,N_18660);
nand U18897 (N_18897,N_18731,N_18635);
and U18898 (N_18898,N_18620,N_18682);
nand U18899 (N_18899,N_18739,N_18717);
and U18900 (N_18900,N_18733,N_18679);
nand U18901 (N_18901,N_18718,N_18787);
and U18902 (N_18902,N_18735,N_18718);
and U18903 (N_18903,N_18647,N_18681);
and U18904 (N_18904,N_18746,N_18751);
nand U18905 (N_18905,N_18711,N_18743);
and U18906 (N_18906,N_18621,N_18717);
nand U18907 (N_18907,N_18734,N_18783);
or U18908 (N_18908,N_18774,N_18738);
xnor U18909 (N_18909,N_18789,N_18618);
nand U18910 (N_18910,N_18689,N_18666);
or U18911 (N_18911,N_18704,N_18707);
xor U18912 (N_18912,N_18715,N_18604);
xnor U18913 (N_18913,N_18691,N_18660);
or U18914 (N_18914,N_18719,N_18670);
or U18915 (N_18915,N_18753,N_18656);
xnor U18916 (N_18916,N_18684,N_18793);
and U18917 (N_18917,N_18630,N_18790);
or U18918 (N_18918,N_18704,N_18637);
nor U18919 (N_18919,N_18713,N_18667);
and U18920 (N_18920,N_18799,N_18714);
and U18921 (N_18921,N_18785,N_18721);
or U18922 (N_18922,N_18700,N_18790);
nand U18923 (N_18923,N_18715,N_18777);
xnor U18924 (N_18924,N_18741,N_18725);
nand U18925 (N_18925,N_18696,N_18791);
xor U18926 (N_18926,N_18656,N_18663);
and U18927 (N_18927,N_18602,N_18744);
xnor U18928 (N_18928,N_18678,N_18753);
or U18929 (N_18929,N_18682,N_18651);
nor U18930 (N_18930,N_18697,N_18742);
or U18931 (N_18931,N_18687,N_18681);
and U18932 (N_18932,N_18615,N_18726);
xnor U18933 (N_18933,N_18641,N_18653);
nand U18934 (N_18934,N_18626,N_18600);
and U18935 (N_18935,N_18769,N_18793);
nand U18936 (N_18936,N_18797,N_18794);
nand U18937 (N_18937,N_18748,N_18770);
nand U18938 (N_18938,N_18768,N_18788);
and U18939 (N_18939,N_18611,N_18654);
xnor U18940 (N_18940,N_18731,N_18727);
or U18941 (N_18941,N_18775,N_18608);
nor U18942 (N_18942,N_18764,N_18745);
nand U18943 (N_18943,N_18717,N_18759);
xor U18944 (N_18944,N_18754,N_18680);
and U18945 (N_18945,N_18773,N_18729);
and U18946 (N_18946,N_18610,N_18748);
and U18947 (N_18947,N_18732,N_18692);
nand U18948 (N_18948,N_18717,N_18667);
or U18949 (N_18949,N_18776,N_18708);
nand U18950 (N_18950,N_18696,N_18775);
and U18951 (N_18951,N_18768,N_18724);
and U18952 (N_18952,N_18734,N_18738);
or U18953 (N_18953,N_18698,N_18788);
or U18954 (N_18954,N_18726,N_18756);
nor U18955 (N_18955,N_18729,N_18711);
or U18956 (N_18956,N_18753,N_18625);
nor U18957 (N_18957,N_18767,N_18777);
nand U18958 (N_18958,N_18707,N_18696);
nor U18959 (N_18959,N_18639,N_18632);
xor U18960 (N_18960,N_18688,N_18742);
xor U18961 (N_18961,N_18609,N_18686);
nor U18962 (N_18962,N_18769,N_18738);
or U18963 (N_18963,N_18724,N_18665);
or U18964 (N_18964,N_18758,N_18705);
and U18965 (N_18965,N_18674,N_18709);
nor U18966 (N_18966,N_18625,N_18606);
and U18967 (N_18967,N_18638,N_18726);
or U18968 (N_18968,N_18638,N_18615);
and U18969 (N_18969,N_18799,N_18703);
xor U18970 (N_18970,N_18706,N_18630);
xnor U18971 (N_18971,N_18778,N_18690);
or U18972 (N_18972,N_18679,N_18768);
and U18973 (N_18973,N_18766,N_18685);
nand U18974 (N_18974,N_18713,N_18749);
nand U18975 (N_18975,N_18736,N_18694);
xnor U18976 (N_18976,N_18714,N_18763);
or U18977 (N_18977,N_18605,N_18784);
and U18978 (N_18978,N_18757,N_18780);
and U18979 (N_18979,N_18774,N_18652);
nand U18980 (N_18980,N_18678,N_18625);
xnor U18981 (N_18981,N_18642,N_18711);
or U18982 (N_18982,N_18613,N_18658);
xor U18983 (N_18983,N_18794,N_18776);
xor U18984 (N_18984,N_18722,N_18708);
and U18985 (N_18985,N_18632,N_18709);
or U18986 (N_18986,N_18687,N_18797);
and U18987 (N_18987,N_18772,N_18725);
nor U18988 (N_18988,N_18736,N_18784);
and U18989 (N_18989,N_18694,N_18696);
xnor U18990 (N_18990,N_18623,N_18768);
and U18991 (N_18991,N_18702,N_18608);
nor U18992 (N_18992,N_18754,N_18776);
xor U18993 (N_18993,N_18741,N_18754);
and U18994 (N_18994,N_18663,N_18686);
or U18995 (N_18995,N_18602,N_18675);
nor U18996 (N_18996,N_18668,N_18744);
or U18997 (N_18997,N_18776,N_18737);
nand U18998 (N_18998,N_18718,N_18733);
and U18999 (N_18999,N_18745,N_18791);
or U19000 (N_19000,N_18834,N_18990);
or U19001 (N_19001,N_18823,N_18881);
or U19002 (N_19002,N_18835,N_18871);
and U19003 (N_19003,N_18978,N_18849);
xor U19004 (N_19004,N_18960,N_18907);
and U19005 (N_19005,N_18864,N_18906);
xor U19006 (N_19006,N_18962,N_18952);
xnor U19007 (N_19007,N_18931,N_18930);
xnor U19008 (N_19008,N_18969,N_18892);
nor U19009 (N_19009,N_18925,N_18987);
and U19010 (N_19010,N_18832,N_18877);
or U19011 (N_19011,N_18827,N_18846);
nand U19012 (N_19012,N_18997,N_18979);
and U19013 (N_19013,N_18982,N_18850);
nor U19014 (N_19014,N_18995,N_18961);
nand U19015 (N_19015,N_18919,N_18911);
or U19016 (N_19016,N_18836,N_18860);
nand U19017 (N_19017,N_18870,N_18803);
or U19018 (N_19018,N_18989,N_18927);
xor U19019 (N_19019,N_18838,N_18888);
nor U19020 (N_19020,N_18894,N_18856);
nor U19021 (N_19021,N_18980,N_18947);
or U19022 (N_19022,N_18878,N_18861);
nor U19023 (N_19023,N_18913,N_18921);
nor U19024 (N_19024,N_18976,N_18844);
nand U19025 (N_19025,N_18967,N_18944);
or U19026 (N_19026,N_18998,N_18889);
nor U19027 (N_19027,N_18984,N_18981);
nand U19028 (N_19028,N_18886,N_18950);
or U19029 (N_19029,N_18959,N_18807);
or U19030 (N_19030,N_18821,N_18988);
and U19031 (N_19031,N_18831,N_18893);
xor U19032 (N_19032,N_18983,N_18882);
and U19033 (N_19033,N_18940,N_18866);
xnor U19034 (N_19034,N_18946,N_18945);
or U19035 (N_19035,N_18942,N_18905);
and U19036 (N_19036,N_18862,N_18923);
nand U19037 (N_19037,N_18966,N_18926);
nor U19038 (N_19038,N_18841,N_18973);
and U19039 (N_19039,N_18898,N_18891);
nand U19040 (N_19040,N_18805,N_18879);
or U19041 (N_19041,N_18824,N_18852);
nor U19042 (N_19042,N_18922,N_18874);
and U19043 (N_19043,N_18817,N_18855);
or U19044 (N_19044,N_18853,N_18816);
xnor U19045 (N_19045,N_18801,N_18932);
xnor U19046 (N_19046,N_18820,N_18804);
or U19047 (N_19047,N_18943,N_18915);
nor U19048 (N_19048,N_18867,N_18939);
and U19049 (N_19049,N_18955,N_18808);
nor U19050 (N_19050,N_18847,N_18840);
nor U19051 (N_19051,N_18992,N_18941);
nor U19052 (N_19052,N_18970,N_18818);
nor U19053 (N_19053,N_18956,N_18986);
or U19054 (N_19054,N_18937,N_18901);
nor U19055 (N_19055,N_18929,N_18876);
xnor U19056 (N_19056,N_18918,N_18996);
nand U19057 (N_19057,N_18813,N_18900);
or U19058 (N_19058,N_18828,N_18934);
nor U19059 (N_19059,N_18916,N_18935);
and U19060 (N_19060,N_18974,N_18897);
nand U19061 (N_19061,N_18958,N_18809);
nor U19062 (N_19062,N_18806,N_18826);
and U19063 (N_19063,N_18910,N_18914);
xor U19064 (N_19064,N_18993,N_18857);
nor U19065 (N_19065,N_18890,N_18972);
nand U19066 (N_19066,N_18953,N_18924);
and U19067 (N_19067,N_18868,N_18903);
or U19068 (N_19068,N_18928,N_18965);
nor U19069 (N_19069,N_18920,N_18895);
nor U19070 (N_19070,N_18971,N_18833);
xnor U19071 (N_19071,N_18896,N_18802);
xor U19072 (N_19072,N_18908,N_18933);
nand U19073 (N_19073,N_18800,N_18872);
nor U19074 (N_19074,N_18951,N_18912);
nor U19075 (N_19075,N_18985,N_18839);
and U19076 (N_19076,N_18873,N_18954);
xor U19077 (N_19077,N_18975,N_18884);
nand U19078 (N_19078,N_18851,N_18863);
or U19079 (N_19079,N_18909,N_18829);
nor U19080 (N_19080,N_18994,N_18999);
and U19081 (N_19081,N_18938,N_18865);
nor U19082 (N_19082,N_18957,N_18858);
xnor U19083 (N_19083,N_18880,N_18814);
and U19084 (N_19084,N_18883,N_18991);
nand U19085 (N_19085,N_18843,N_18904);
or U19086 (N_19086,N_18842,N_18810);
xnor U19087 (N_19087,N_18968,N_18899);
or U19088 (N_19088,N_18869,N_18948);
nand U19089 (N_19089,N_18854,N_18936);
or U19090 (N_19090,N_18815,N_18949);
xnor U19091 (N_19091,N_18819,N_18875);
nor U19092 (N_19092,N_18825,N_18963);
and U19093 (N_19093,N_18977,N_18845);
and U19094 (N_19094,N_18830,N_18812);
xor U19095 (N_19095,N_18811,N_18848);
nand U19096 (N_19096,N_18859,N_18887);
and U19097 (N_19097,N_18964,N_18902);
or U19098 (N_19098,N_18822,N_18837);
nand U19099 (N_19099,N_18917,N_18885);
and U19100 (N_19100,N_18941,N_18863);
xnor U19101 (N_19101,N_18831,N_18948);
and U19102 (N_19102,N_18893,N_18876);
and U19103 (N_19103,N_18802,N_18881);
nand U19104 (N_19104,N_18867,N_18917);
xor U19105 (N_19105,N_18894,N_18934);
xor U19106 (N_19106,N_18974,N_18935);
nand U19107 (N_19107,N_18826,N_18973);
xor U19108 (N_19108,N_18824,N_18951);
or U19109 (N_19109,N_18823,N_18959);
nor U19110 (N_19110,N_18914,N_18900);
and U19111 (N_19111,N_18846,N_18941);
nand U19112 (N_19112,N_18830,N_18801);
or U19113 (N_19113,N_18936,N_18960);
xor U19114 (N_19114,N_18824,N_18877);
nor U19115 (N_19115,N_18840,N_18976);
and U19116 (N_19116,N_18937,N_18858);
and U19117 (N_19117,N_18847,N_18823);
xnor U19118 (N_19118,N_18991,N_18852);
xnor U19119 (N_19119,N_18947,N_18934);
and U19120 (N_19120,N_18857,N_18984);
nor U19121 (N_19121,N_18959,N_18800);
nor U19122 (N_19122,N_18920,N_18957);
nand U19123 (N_19123,N_18949,N_18812);
nand U19124 (N_19124,N_18860,N_18829);
nor U19125 (N_19125,N_18977,N_18994);
nand U19126 (N_19126,N_18858,N_18844);
nor U19127 (N_19127,N_18867,N_18884);
xnor U19128 (N_19128,N_18905,N_18811);
nor U19129 (N_19129,N_18805,N_18997);
and U19130 (N_19130,N_18882,N_18970);
xnor U19131 (N_19131,N_18953,N_18894);
or U19132 (N_19132,N_18911,N_18880);
and U19133 (N_19133,N_18807,N_18882);
or U19134 (N_19134,N_18844,N_18803);
nor U19135 (N_19135,N_18811,N_18807);
or U19136 (N_19136,N_18984,N_18818);
nand U19137 (N_19137,N_18868,N_18832);
nand U19138 (N_19138,N_18918,N_18997);
nor U19139 (N_19139,N_18993,N_18836);
and U19140 (N_19140,N_18910,N_18884);
xor U19141 (N_19141,N_18902,N_18838);
xor U19142 (N_19142,N_18911,N_18991);
nor U19143 (N_19143,N_18916,N_18891);
nand U19144 (N_19144,N_18864,N_18862);
nor U19145 (N_19145,N_18848,N_18940);
and U19146 (N_19146,N_18824,N_18949);
nand U19147 (N_19147,N_18899,N_18885);
nand U19148 (N_19148,N_18935,N_18894);
nor U19149 (N_19149,N_18914,N_18904);
nor U19150 (N_19150,N_18988,N_18815);
nand U19151 (N_19151,N_18992,N_18915);
and U19152 (N_19152,N_18888,N_18886);
nand U19153 (N_19153,N_18808,N_18837);
nor U19154 (N_19154,N_18926,N_18813);
and U19155 (N_19155,N_18838,N_18965);
nand U19156 (N_19156,N_18821,N_18817);
xnor U19157 (N_19157,N_18882,N_18857);
nand U19158 (N_19158,N_18884,N_18860);
nor U19159 (N_19159,N_18986,N_18856);
or U19160 (N_19160,N_18835,N_18802);
and U19161 (N_19161,N_18958,N_18801);
and U19162 (N_19162,N_18847,N_18944);
or U19163 (N_19163,N_18849,N_18832);
xnor U19164 (N_19164,N_18984,N_18894);
or U19165 (N_19165,N_18862,N_18898);
xnor U19166 (N_19166,N_18945,N_18979);
or U19167 (N_19167,N_18806,N_18964);
nor U19168 (N_19168,N_18873,N_18972);
or U19169 (N_19169,N_18932,N_18857);
nor U19170 (N_19170,N_18872,N_18964);
nand U19171 (N_19171,N_18931,N_18835);
nand U19172 (N_19172,N_18887,N_18924);
nand U19173 (N_19173,N_18876,N_18952);
and U19174 (N_19174,N_18958,N_18882);
nand U19175 (N_19175,N_18808,N_18803);
nor U19176 (N_19176,N_18893,N_18805);
xnor U19177 (N_19177,N_18886,N_18921);
or U19178 (N_19178,N_18823,N_18809);
or U19179 (N_19179,N_18997,N_18812);
or U19180 (N_19180,N_18928,N_18857);
or U19181 (N_19181,N_18804,N_18916);
nand U19182 (N_19182,N_18902,N_18853);
xnor U19183 (N_19183,N_18974,N_18885);
nand U19184 (N_19184,N_18976,N_18938);
and U19185 (N_19185,N_18818,N_18890);
and U19186 (N_19186,N_18801,N_18850);
nor U19187 (N_19187,N_18824,N_18990);
or U19188 (N_19188,N_18943,N_18981);
nor U19189 (N_19189,N_18909,N_18974);
or U19190 (N_19190,N_18916,N_18825);
xor U19191 (N_19191,N_18919,N_18870);
nor U19192 (N_19192,N_18889,N_18961);
or U19193 (N_19193,N_18819,N_18818);
nand U19194 (N_19194,N_18957,N_18930);
or U19195 (N_19195,N_18950,N_18947);
nand U19196 (N_19196,N_18889,N_18914);
nor U19197 (N_19197,N_18902,N_18922);
or U19198 (N_19198,N_18910,N_18856);
xnor U19199 (N_19199,N_18877,N_18869);
and U19200 (N_19200,N_19150,N_19112);
nand U19201 (N_19201,N_19199,N_19120);
xor U19202 (N_19202,N_19029,N_19187);
xnor U19203 (N_19203,N_19031,N_19050);
and U19204 (N_19204,N_19122,N_19066);
nand U19205 (N_19205,N_19076,N_19111);
or U19206 (N_19206,N_19190,N_19065);
and U19207 (N_19207,N_19098,N_19093);
nand U19208 (N_19208,N_19023,N_19035);
or U19209 (N_19209,N_19056,N_19138);
xnor U19210 (N_19210,N_19154,N_19007);
nand U19211 (N_19211,N_19020,N_19036);
nor U19212 (N_19212,N_19025,N_19040);
xnor U19213 (N_19213,N_19133,N_19169);
nand U19214 (N_19214,N_19081,N_19090);
nand U19215 (N_19215,N_19057,N_19083);
nor U19216 (N_19216,N_19004,N_19127);
nand U19217 (N_19217,N_19192,N_19185);
nor U19218 (N_19218,N_19195,N_19148);
or U19219 (N_19219,N_19032,N_19074);
or U19220 (N_19220,N_19028,N_19003);
or U19221 (N_19221,N_19097,N_19108);
nor U19222 (N_19222,N_19100,N_19165);
nand U19223 (N_19223,N_19082,N_19049);
xnor U19224 (N_19224,N_19151,N_19062);
or U19225 (N_19225,N_19037,N_19153);
and U19226 (N_19226,N_19172,N_19181);
nor U19227 (N_19227,N_19184,N_19183);
or U19228 (N_19228,N_19136,N_19053);
and U19229 (N_19229,N_19134,N_19188);
nor U19230 (N_19230,N_19140,N_19061);
nor U19231 (N_19231,N_19171,N_19010);
or U19232 (N_19232,N_19147,N_19086);
nor U19233 (N_19233,N_19158,N_19119);
nand U19234 (N_19234,N_19177,N_19033);
and U19235 (N_19235,N_19071,N_19016);
nand U19236 (N_19236,N_19149,N_19135);
and U19237 (N_19237,N_19042,N_19159);
or U19238 (N_19238,N_19052,N_19030);
and U19239 (N_19239,N_19123,N_19026);
nor U19240 (N_19240,N_19193,N_19069);
and U19241 (N_19241,N_19005,N_19045);
or U19242 (N_19242,N_19106,N_19131);
xor U19243 (N_19243,N_19046,N_19179);
nor U19244 (N_19244,N_19137,N_19144);
and U19245 (N_19245,N_19019,N_19164);
xnor U19246 (N_19246,N_19099,N_19104);
and U19247 (N_19247,N_19006,N_19008);
xor U19248 (N_19248,N_19160,N_19072);
xnor U19249 (N_19249,N_19067,N_19121);
nor U19250 (N_19250,N_19156,N_19048);
nor U19251 (N_19251,N_19178,N_19110);
nor U19252 (N_19252,N_19196,N_19091);
and U19253 (N_19253,N_19087,N_19014);
and U19254 (N_19254,N_19115,N_19182);
xnor U19255 (N_19255,N_19012,N_19168);
or U19256 (N_19256,N_19064,N_19039);
and U19257 (N_19257,N_19034,N_19130);
xnor U19258 (N_19258,N_19145,N_19013);
nand U19259 (N_19259,N_19051,N_19162);
nand U19260 (N_19260,N_19024,N_19022);
nor U19261 (N_19261,N_19092,N_19079);
and U19262 (N_19262,N_19094,N_19078);
and U19263 (N_19263,N_19103,N_19089);
or U19264 (N_19264,N_19043,N_19001);
or U19265 (N_19265,N_19139,N_19125);
or U19266 (N_19266,N_19174,N_19070);
nand U19267 (N_19267,N_19021,N_19068);
xor U19268 (N_19268,N_19161,N_19117);
xnor U19269 (N_19269,N_19102,N_19059);
nand U19270 (N_19270,N_19143,N_19085);
nand U19271 (N_19271,N_19038,N_19197);
or U19272 (N_19272,N_19186,N_19060);
xnor U19273 (N_19273,N_19166,N_19101);
and U19274 (N_19274,N_19084,N_19096);
nor U19275 (N_19275,N_19054,N_19132);
xor U19276 (N_19276,N_19107,N_19194);
and U19277 (N_19277,N_19167,N_19088);
and U19278 (N_19278,N_19015,N_19146);
xor U19279 (N_19279,N_19163,N_19017);
nor U19280 (N_19280,N_19000,N_19128);
nor U19281 (N_19281,N_19155,N_19129);
nand U19282 (N_19282,N_19113,N_19027);
xor U19283 (N_19283,N_19189,N_19047);
xnor U19284 (N_19284,N_19063,N_19124);
nor U19285 (N_19285,N_19073,N_19105);
nand U19286 (N_19286,N_19011,N_19141);
nor U19287 (N_19287,N_19191,N_19142);
nand U19288 (N_19288,N_19116,N_19114);
nor U19289 (N_19289,N_19175,N_19157);
nand U19290 (N_19290,N_19109,N_19152);
or U19291 (N_19291,N_19095,N_19018);
nor U19292 (N_19292,N_19075,N_19058);
nor U19293 (N_19293,N_19044,N_19055);
xnor U19294 (N_19294,N_19118,N_19198);
nand U19295 (N_19295,N_19002,N_19080);
nor U19296 (N_19296,N_19126,N_19176);
and U19297 (N_19297,N_19173,N_19077);
nand U19298 (N_19298,N_19041,N_19009);
and U19299 (N_19299,N_19180,N_19170);
nor U19300 (N_19300,N_19162,N_19013);
or U19301 (N_19301,N_19095,N_19079);
nor U19302 (N_19302,N_19064,N_19065);
nor U19303 (N_19303,N_19137,N_19076);
and U19304 (N_19304,N_19189,N_19071);
or U19305 (N_19305,N_19024,N_19157);
nand U19306 (N_19306,N_19113,N_19105);
and U19307 (N_19307,N_19120,N_19049);
and U19308 (N_19308,N_19175,N_19115);
or U19309 (N_19309,N_19068,N_19069);
and U19310 (N_19310,N_19199,N_19097);
or U19311 (N_19311,N_19182,N_19085);
xor U19312 (N_19312,N_19091,N_19143);
and U19313 (N_19313,N_19169,N_19178);
xor U19314 (N_19314,N_19163,N_19108);
xor U19315 (N_19315,N_19191,N_19123);
nor U19316 (N_19316,N_19166,N_19011);
nor U19317 (N_19317,N_19118,N_19190);
or U19318 (N_19318,N_19121,N_19155);
nand U19319 (N_19319,N_19135,N_19039);
nand U19320 (N_19320,N_19121,N_19073);
nor U19321 (N_19321,N_19166,N_19057);
and U19322 (N_19322,N_19062,N_19120);
xor U19323 (N_19323,N_19002,N_19011);
or U19324 (N_19324,N_19108,N_19194);
or U19325 (N_19325,N_19118,N_19009);
or U19326 (N_19326,N_19008,N_19063);
or U19327 (N_19327,N_19111,N_19104);
xnor U19328 (N_19328,N_19088,N_19146);
nand U19329 (N_19329,N_19161,N_19119);
or U19330 (N_19330,N_19111,N_19115);
nor U19331 (N_19331,N_19174,N_19103);
or U19332 (N_19332,N_19028,N_19158);
and U19333 (N_19333,N_19040,N_19117);
nor U19334 (N_19334,N_19025,N_19103);
nor U19335 (N_19335,N_19035,N_19017);
and U19336 (N_19336,N_19112,N_19129);
nor U19337 (N_19337,N_19024,N_19042);
and U19338 (N_19338,N_19077,N_19186);
nor U19339 (N_19339,N_19017,N_19031);
nor U19340 (N_19340,N_19123,N_19043);
or U19341 (N_19341,N_19100,N_19096);
and U19342 (N_19342,N_19165,N_19145);
or U19343 (N_19343,N_19046,N_19090);
and U19344 (N_19344,N_19155,N_19094);
and U19345 (N_19345,N_19079,N_19003);
and U19346 (N_19346,N_19055,N_19061);
or U19347 (N_19347,N_19099,N_19129);
xnor U19348 (N_19348,N_19113,N_19157);
nor U19349 (N_19349,N_19064,N_19116);
nor U19350 (N_19350,N_19048,N_19040);
nand U19351 (N_19351,N_19091,N_19187);
xnor U19352 (N_19352,N_19032,N_19106);
or U19353 (N_19353,N_19183,N_19000);
xnor U19354 (N_19354,N_19170,N_19004);
nand U19355 (N_19355,N_19047,N_19082);
or U19356 (N_19356,N_19132,N_19135);
nor U19357 (N_19357,N_19087,N_19016);
xor U19358 (N_19358,N_19119,N_19111);
or U19359 (N_19359,N_19189,N_19179);
and U19360 (N_19360,N_19146,N_19112);
or U19361 (N_19361,N_19059,N_19032);
nor U19362 (N_19362,N_19148,N_19078);
nand U19363 (N_19363,N_19147,N_19134);
nand U19364 (N_19364,N_19079,N_19122);
or U19365 (N_19365,N_19128,N_19165);
nor U19366 (N_19366,N_19021,N_19149);
nor U19367 (N_19367,N_19166,N_19177);
or U19368 (N_19368,N_19035,N_19081);
or U19369 (N_19369,N_19159,N_19118);
and U19370 (N_19370,N_19002,N_19121);
nand U19371 (N_19371,N_19045,N_19128);
or U19372 (N_19372,N_19119,N_19054);
or U19373 (N_19373,N_19066,N_19194);
nor U19374 (N_19374,N_19036,N_19028);
nor U19375 (N_19375,N_19001,N_19126);
xor U19376 (N_19376,N_19109,N_19111);
and U19377 (N_19377,N_19174,N_19068);
nand U19378 (N_19378,N_19105,N_19038);
or U19379 (N_19379,N_19164,N_19027);
nor U19380 (N_19380,N_19098,N_19166);
xnor U19381 (N_19381,N_19115,N_19009);
or U19382 (N_19382,N_19032,N_19199);
and U19383 (N_19383,N_19080,N_19071);
and U19384 (N_19384,N_19151,N_19025);
and U19385 (N_19385,N_19129,N_19017);
and U19386 (N_19386,N_19128,N_19199);
nor U19387 (N_19387,N_19062,N_19055);
nand U19388 (N_19388,N_19166,N_19042);
nor U19389 (N_19389,N_19195,N_19018);
xnor U19390 (N_19390,N_19169,N_19089);
nor U19391 (N_19391,N_19027,N_19122);
xor U19392 (N_19392,N_19107,N_19182);
or U19393 (N_19393,N_19055,N_19008);
or U19394 (N_19394,N_19117,N_19045);
or U19395 (N_19395,N_19184,N_19020);
nor U19396 (N_19396,N_19196,N_19074);
or U19397 (N_19397,N_19032,N_19004);
xnor U19398 (N_19398,N_19130,N_19122);
nor U19399 (N_19399,N_19073,N_19065);
nand U19400 (N_19400,N_19370,N_19291);
nor U19401 (N_19401,N_19391,N_19327);
xnor U19402 (N_19402,N_19280,N_19259);
nand U19403 (N_19403,N_19384,N_19271);
or U19404 (N_19404,N_19237,N_19215);
and U19405 (N_19405,N_19371,N_19216);
nand U19406 (N_19406,N_19240,N_19356);
xnor U19407 (N_19407,N_19267,N_19312);
nand U19408 (N_19408,N_19263,N_19253);
xor U19409 (N_19409,N_19339,N_19392);
xnor U19410 (N_19410,N_19347,N_19288);
and U19411 (N_19411,N_19234,N_19287);
nand U19412 (N_19412,N_19285,N_19309);
nor U19413 (N_19413,N_19290,N_19310);
or U19414 (N_19414,N_19250,N_19213);
and U19415 (N_19415,N_19218,N_19251);
and U19416 (N_19416,N_19390,N_19334);
nor U19417 (N_19417,N_19329,N_19346);
nor U19418 (N_19418,N_19266,N_19387);
nor U19419 (N_19419,N_19324,N_19393);
xnor U19420 (N_19420,N_19252,N_19340);
xor U19421 (N_19421,N_19206,N_19281);
nand U19422 (N_19422,N_19325,N_19269);
xor U19423 (N_19423,N_19395,N_19223);
or U19424 (N_19424,N_19283,N_19233);
or U19425 (N_19425,N_19374,N_19232);
xor U19426 (N_19426,N_19294,N_19338);
nor U19427 (N_19427,N_19228,N_19236);
nand U19428 (N_19428,N_19335,N_19397);
and U19429 (N_19429,N_19368,N_19214);
and U19430 (N_19430,N_19224,N_19209);
nor U19431 (N_19431,N_19201,N_19320);
nor U19432 (N_19432,N_19270,N_19332);
nand U19433 (N_19433,N_19382,N_19345);
nand U19434 (N_19434,N_19377,N_19372);
nand U19435 (N_19435,N_19272,N_19292);
and U19436 (N_19436,N_19373,N_19348);
xor U19437 (N_19437,N_19254,N_19255);
xnor U19438 (N_19438,N_19378,N_19319);
nor U19439 (N_19439,N_19304,N_19256);
nor U19440 (N_19440,N_19248,N_19361);
nor U19441 (N_19441,N_19313,N_19200);
nor U19442 (N_19442,N_19260,N_19308);
and U19443 (N_19443,N_19221,N_19311);
nor U19444 (N_19444,N_19351,N_19398);
and U19445 (N_19445,N_19273,N_19362);
and U19446 (N_19446,N_19314,N_19386);
and U19447 (N_19447,N_19336,N_19366);
xor U19448 (N_19448,N_19249,N_19241);
nor U19449 (N_19449,N_19350,N_19303);
nor U19450 (N_19450,N_19278,N_19330);
nand U19451 (N_19451,N_19204,N_19217);
nand U19452 (N_19452,N_19379,N_19326);
or U19453 (N_19453,N_19355,N_19245);
nand U19454 (N_19454,N_19360,N_19305);
nand U19455 (N_19455,N_19363,N_19293);
xor U19456 (N_19456,N_19396,N_19297);
or U19457 (N_19457,N_19277,N_19227);
or U19458 (N_19458,N_19383,N_19202);
nand U19459 (N_19459,N_19220,N_19229);
nand U19460 (N_19460,N_19295,N_19357);
and U19461 (N_19461,N_19265,N_19344);
xor U19462 (N_19462,N_19301,N_19289);
or U19463 (N_19463,N_19230,N_19210);
or U19464 (N_19464,N_19364,N_19274);
and U19465 (N_19465,N_19337,N_19333);
nor U19466 (N_19466,N_19238,N_19211);
or U19467 (N_19467,N_19321,N_19231);
xnor U19468 (N_19468,N_19322,N_19208);
nor U19469 (N_19469,N_19367,N_19296);
nor U19470 (N_19470,N_19316,N_19389);
xnor U19471 (N_19471,N_19318,N_19235);
nor U19472 (N_19472,N_19342,N_19261);
nor U19473 (N_19473,N_19205,N_19225);
and U19474 (N_19474,N_19307,N_19258);
and U19475 (N_19475,N_19212,N_19388);
nand U19476 (N_19476,N_19222,N_19331);
xnor U19477 (N_19477,N_19376,N_19246);
nor U19478 (N_19478,N_19323,N_19306);
or U19479 (N_19479,N_19247,N_19243);
nor U19480 (N_19480,N_19399,N_19341);
nor U19481 (N_19481,N_19359,N_19275);
xor U19482 (N_19482,N_19257,N_19207);
or U19483 (N_19483,N_19244,N_19375);
and U19484 (N_19484,N_19239,N_19242);
xnor U19485 (N_19485,N_19299,N_19381);
nand U19486 (N_19486,N_19226,N_19264);
or U19487 (N_19487,N_19385,N_19268);
xor U19488 (N_19488,N_19349,N_19365);
nor U19489 (N_19489,N_19300,N_19394);
or U19490 (N_19490,N_19282,N_19380);
nand U19491 (N_19491,N_19328,N_19315);
xor U19492 (N_19492,N_19317,N_19358);
nor U19493 (N_19493,N_19369,N_19302);
or U19494 (N_19494,N_19262,N_19352);
or U19495 (N_19495,N_19203,N_19343);
nand U19496 (N_19496,N_19284,N_19286);
and U19497 (N_19497,N_19276,N_19353);
nand U19498 (N_19498,N_19279,N_19219);
xor U19499 (N_19499,N_19298,N_19354);
and U19500 (N_19500,N_19352,N_19388);
nand U19501 (N_19501,N_19318,N_19308);
and U19502 (N_19502,N_19344,N_19289);
nand U19503 (N_19503,N_19359,N_19272);
xor U19504 (N_19504,N_19315,N_19210);
or U19505 (N_19505,N_19397,N_19371);
nor U19506 (N_19506,N_19268,N_19219);
nand U19507 (N_19507,N_19200,N_19334);
nor U19508 (N_19508,N_19353,N_19216);
nor U19509 (N_19509,N_19369,N_19238);
or U19510 (N_19510,N_19285,N_19385);
xor U19511 (N_19511,N_19378,N_19377);
xnor U19512 (N_19512,N_19302,N_19247);
xnor U19513 (N_19513,N_19267,N_19226);
or U19514 (N_19514,N_19342,N_19344);
nor U19515 (N_19515,N_19344,N_19234);
xnor U19516 (N_19516,N_19365,N_19212);
xnor U19517 (N_19517,N_19359,N_19244);
xor U19518 (N_19518,N_19217,N_19346);
nor U19519 (N_19519,N_19271,N_19219);
nor U19520 (N_19520,N_19281,N_19306);
nand U19521 (N_19521,N_19305,N_19316);
and U19522 (N_19522,N_19332,N_19215);
or U19523 (N_19523,N_19227,N_19274);
xnor U19524 (N_19524,N_19293,N_19276);
nand U19525 (N_19525,N_19235,N_19345);
and U19526 (N_19526,N_19258,N_19204);
nand U19527 (N_19527,N_19396,N_19332);
nor U19528 (N_19528,N_19246,N_19210);
or U19529 (N_19529,N_19348,N_19310);
xnor U19530 (N_19530,N_19309,N_19322);
xnor U19531 (N_19531,N_19389,N_19269);
nor U19532 (N_19532,N_19263,N_19360);
nor U19533 (N_19533,N_19237,N_19343);
and U19534 (N_19534,N_19378,N_19360);
nand U19535 (N_19535,N_19220,N_19271);
or U19536 (N_19536,N_19214,N_19209);
nand U19537 (N_19537,N_19275,N_19263);
nor U19538 (N_19538,N_19327,N_19366);
and U19539 (N_19539,N_19370,N_19268);
nand U19540 (N_19540,N_19379,N_19249);
nor U19541 (N_19541,N_19230,N_19221);
or U19542 (N_19542,N_19346,N_19236);
or U19543 (N_19543,N_19263,N_19244);
xnor U19544 (N_19544,N_19307,N_19303);
xnor U19545 (N_19545,N_19252,N_19391);
nand U19546 (N_19546,N_19384,N_19206);
nor U19547 (N_19547,N_19391,N_19377);
xnor U19548 (N_19548,N_19287,N_19248);
nor U19549 (N_19549,N_19206,N_19209);
xnor U19550 (N_19550,N_19224,N_19249);
or U19551 (N_19551,N_19389,N_19337);
and U19552 (N_19552,N_19324,N_19230);
nor U19553 (N_19553,N_19245,N_19282);
or U19554 (N_19554,N_19204,N_19348);
nand U19555 (N_19555,N_19303,N_19373);
xnor U19556 (N_19556,N_19241,N_19296);
xnor U19557 (N_19557,N_19329,N_19334);
nor U19558 (N_19558,N_19274,N_19268);
nand U19559 (N_19559,N_19299,N_19239);
nor U19560 (N_19560,N_19385,N_19237);
or U19561 (N_19561,N_19383,N_19382);
nor U19562 (N_19562,N_19327,N_19399);
and U19563 (N_19563,N_19287,N_19326);
xor U19564 (N_19564,N_19207,N_19391);
nor U19565 (N_19565,N_19350,N_19372);
nor U19566 (N_19566,N_19298,N_19362);
xnor U19567 (N_19567,N_19340,N_19346);
xor U19568 (N_19568,N_19269,N_19341);
and U19569 (N_19569,N_19230,N_19272);
xor U19570 (N_19570,N_19353,N_19248);
nand U19571 (N_19571,N_19310,N_19352);
nor U19572 (N_19572,N_19302,N_19271);
or U19573 (N_19573,N_19327,N_19357);
nand U19574 (N_19574,N_19370,N_19376);
or U19575 (N_19575,N_19387,N_19294);
and U19576 (N_19576,N_19327,N_19204);
or U19577 (N_19577,N_19242,N_19226);
nor U19578 (N_19578,N_19331,N_19288);
and U19579 (N_19579,N_19234,N_19338);
xnor U19580 (N_19580,N_19246,N_19374);
or U19581 (N_19581,N_19264,N_19347);
and U19582 (N_19582,N_19300,N_19332);
xnor U19583 (N_19583,N_19305,N_19351);
and U19584 (N_19584,N_19278,N_19329);
and U19585 (N_19585,N_19291,N_19350);
nand U19586 (N_19586,N_19273,N_19350);
or U19587 (N_19587,N_19331,N_19322);
nor U19588 (N_19588,N_19361,N_19229);
or U19589 (N_19589,N_19224,N_19374);
and U19590 (N_19590,N_19269,N_19309);
nand U19591 (N_19591,N_19311,N_19306);
and U19592 (N_19592,N_19283,N_19396);
nand U19593 (N_19593,N_19210,N_19240);
and U19594 (N_19594,N_19209,N_19354);
or U19595 (N_19595,N_19278,N_19283);
or U19596 (N_19596,N_19280,N_19207);
or U19597 (N_19597,N_19223,N_19308);
nand U19598 (N_19598,N_19346,N_19304);
nand U19599 (N_19599,N_19362,N_19334);
or U19600 (N_19600,N_19442,N_19528);
nor U19601 (N_19601,N_19495,N_19587);
xnor U19602 (N_19602,N_19417,N_19501);
nand U19603 (N_19603,N_19449,N_19582);
nor U19604 (N_19604,N_19540,N_19592);
and U19605 (N_19605,N_19552,N_19597);
or U19606 (N_19606,N_19457,N_19469);
nand U19607 (N_19607,N_19524,N_19508);
xor U19608 (N_19608,N_19547,N_19583);
nor U19609 (N_19609,N_19473,N_19565);
xor U19610 (N_19610,N_19496,N_19415);
and U19611 (N_19611,N_19408,N_19472);
xor U19612 (N_19612,N_19579,N_19533);
or U19613 (N_19613,N_19514,N_19414);
nor U19614 (N_19614,N_19537,N_19439);
nand U19615 (N_19615,N_19440,N_19541);
and U19616 (N_19616,N_19577,N_19578);
and U19617 (N_19617,N_19598,N_19551);
nand U19618 (N_19618,N_19484,N_19557);
xor U19619 (N_19619,N_19492,N_19490);
or U19620 (N_19620,N_19544,N_19482);
or U19621 (N_19621,N_19402,N_19571);
nand U19622 (N_19622,N_19568,N_19520);
and U19623 (N_19623,N_19521,N_19530);
nor U19624 (N_19624,N_19455,N_19412);
nand U19625 (N_19625,N_19574,N_19462);
nor U19626 (N_19626,N_19599,N_19554);
nor U19627 (N_19627,N_19487,N_19588);
and U19628 (N_19628,N_19543,N_19448);
xor U19629 (N_19629,N_19411,N_19536);
or U19630 (N_19630,N_19546,N_19403);
or U19631 (N_19631,N_19447,N_19507);
nor U19632 (N_19632,N_19566,N_19575);
xor U19633 (N_19633,N_19405,N_19419);
or U19634 (N_19634,N_19561,N_19517);
nor U19635 (N_19635,N_19460,N_19453);
and U19636 (N_19636,N_19452,N_19426);
nand U19637 (N_19637,N_19585,N_19576);
and U19638 (N_19638,N_19589,N_19503);
nor U19639 (N_19639,N_19502,N_19489);
nand U19640 (N_19640,N_19459,N_19534);
xnor U19641 (N_19641,N_19400,N_19564);
nor U19642 (N_19642,N_19545,N_19468);
nand U19643 (N_19643,N_19478,N_19481);
or U19644 (N_19644,N_19515,N_19525);
nand U19645 (N_19645,N_19477,N_19416);
or U19646 (N_19646,N_19569,N_19479);
or U19647 (N_19647,N_19433,N_19444);
and U19648 (N_19648,N_19538,N_19466);
nor U19649 (N_19649,N_19532,N_19458);
and U19650 (N_19650,N_19559,N_19553);
nand U19651 (N_19651,N_19596,N_19527);
and U19652 (N_19652,N_19435,N_19456);
nor U19653 (N_19653,N_19558,N_19590);
nand U19654 (N_19654,N_19573,N_19471);
nand U19655 (N_19655,N_19465,N_19486);
and U19656 (N_19656,N_19421,N_19483);
nor U19657 (N_19657,N_19406,N_19498);
xor U19658 (N_19658,N_19427,N_19429);
and U19659 (N_19659,N_19556,N_19511);
or U19660 (N_19660,N_19488,N_19494);
nand U19661 (N_19661,N_19470,N_19423);
or U19662 (N_19662,N_19497,N_19594);
nor U19663 (N_19663,N_19461,N_19441);
and U19664 (N_19664,N_19567,N_19531);
nor U19665 (N_19665,N_19504,N_19542);
or U19666 (N_19666,N_19550,N_19560);
xor U19667 (N_19667,N_19450,N_19432);
nor U19668 (N_19668,N_19445,N_19430);
and U19669 (N_19669,N_19424,N_19493);
nand U19670 (N_19670,N_19467,N_19518);
or U19671 (N_19671,N_19500,N_19431);
nand U19672 (N_19672,N_19513,N_19475);
or U19673 (N_19673,N_19474,N_19401);
nand U19674 (N_19674,N_19464,N_19436);
or U19675 (N_19675,N_19404,N_19437);
xor U19676 (N_19676,N_19491,N_19584);
nand U19677 (N_19677,N_19410,N_19522);
nor U19678 (N_19678,N_19454,N_19512);
nor U19679 (N_19679,N_19506,N_19463);
or U19680 (N_19680,N_19420,N_19519);
or U19681 (N_19681,N_19593,N_19570);
nand U19682 (N_19682,N_19529,N_19418);
and U19683 (N_19683,N_19446,N_19516);
nor U19684 (N_19684,N_19555,N_19409);
nor U19685 (N_19685,N_19422,N_19451);
nand U19686 (N_19686,N_19476,N_19581);
nor U19687 (N_19687,N_19428,N_19549);
xnor U19688 (N_19688,N_19563,N_19425);
nor U19689 (N_19689,N_19505,N_19510);
nor U19690 (N_19690,N_19443,N_19580);
nand U19691 (N_19691,N_19572,N_19438);
nor U19692 (N_19692,N_19526,N_19413);
or U19693 (N_19693,N_19485,N_19434);
nand U19694 (N_19694,N_19480,N_19586);
nor U19695 (N_19695,N_19499,N_19509);
xor U19696 (N_19696,N_19407,N_19548);
xor U19697 (N_19697,N_19595,N_19535);
nand U19698 (N_19698,N_19562,N_19539);
nand U19699 (N_19699,N_19523,N_19591);
xor U19700 (N_19700,N_19534,N_19530);
or U19701 (N_19701,N_19503,N_19405);
nand U19702 (N_19702,N_19519,N_19514);
or U19703 (N_19703,N_19596,N_19598);
and U19704 (N_19704,N_19586,N_19577);
or U19705 (N_19705,N_19420,N_19567);
and U19706 (N_19706,N_19528,N_19435);
nor U19707 (N_19707,N_19468,N_19511);
nand U19708 (N_19708,N_19506,N_19473);
or U19709 (N_19709,N_19416,N_19430);
nor U19710 (N_19710,N_19479,N_19484);
or U19711 (N_19711,N_19574,N_19448);
nand U19712 (N_19712,N_19496,N_19533);
nand U19713 (N_19713,N_19496,N_19445);
nor U19714 (N_19714,N_19487,N_19424);
and U19715 (N_19715,N_19539,N_19422);
or U19716 (N_19716,N_19586,N_19477);
xnor U19717 (N_19717,N_19584,N_19432);
nand U19718 (N_19718,N_19542,N_19572);
nor U19719 (N_19719,N_19404,N_19543);
xor U19720 (N_19720,N_19548,N_19515);
xor U19721 (N_19721,N_19498,N_19554);
nor U19722 (N_19722,N_19561,N_19538);
nor U19723 (N_19723,N_19555,N_19491);
and U19724 (N_19724,N_19481,N_19402);
or U19725 (N_19725,N_19411,N_19456);
nor U19726 (N_19726,N_19433,N_19591);
nor U19727 (N_19727,N_19445,N_19568);
nor U19728 (N_19728,N_19451,N_19597);
nor U19729 (N_19729,N_19493,N_19558);
or U19730 (N_19730,N_19505,N_19597);
nor U19731 (N_19731,N_19445,N_19454);
nor U19732 (N_19732,N_19549,N_19532);
and U19733 (N_19733,N_19593,N_19557);
xor U19734 (N_19734,N_19401,N_19586);
or U19735 (N_19735,N_19407,N_19459);
nor U19736 (N_19736,N_19493,N_19406);
nand U19737 (N_19737,N_19483,N_19451);
and U19738 (N_19738,N_19482,N_19499);
xor U19739 (N_19739,N_19557,N_19576);
xor U19740 (N_19740,N_19588,N_19549);
nand U19741 (N_19741,N_19572,N_19480);
or U19742 (N_19742,N_19401,N_19574);
or U19743 (N_19743,N_19433,N_19597);
or U19744 (N_19744,N_19410,N_19544);
and U19745 (N_19745,N_19507,N_19511);
and U19746 (N_19746,N_19499,N_19438);
and U19747 (N_19747,N_19598,N_19588);
nand U19748 (N_19748,N_19472,N_19484);
and U19749 (N_19749,N_19474,N_19407);
xnor U19750 (N_19750,N_19506,N_19492);
xor U19751 (N_19751,N_19501,N_19418);
nor U19752 (N_19752,N_19529,N_19484);
and U19753 (N_19753,N_19471,N_19578);
nor U19754 (N_19754,N_19499,N_19498);
and U19755 (N_19755,N_19565,N_19427);
nand U19756 (N_19756,N_19437,N_19509);
nand U19757 (N_19757,N_19400,N_19413);
xnor U19758 (N_19758,N_19457,N_19431);
and U19759 (N_19759,N_19573,N_19440);
nand U19760 (N_19760,N_19410,N_19514);
nand U19761 (N_19761,N_19552,N_19513);
and U19762 (N_19762,N_19508,N_19585);
xor U19763 (N_19763,N_19506,N_19471);
and U19764 (N_19764,N_19426,N_19511);
nor U19765 (N_19765,N_19476,N_19580);
nand U19766 (N_19766,N_19514,N_19533);
nand U19767 (N_19767,N_19457,N_19571);
or U19768 (N_19768,N_19516,N_19483);
nor U19769 (N_19769,N_19570,N_19568);
and U19770 (N_19770,N_19561,N_19421);
nand U19771 (N_19771,N_19509,N_19431);
xnor U19772 (N_19772,N_19488,N_19549);
and U19773 (N_19773,N_19444,N_19531);
nand U19774 (N_19774,N_19406,N_19590);
nor U19775 (N_19775,N_19576,N_19517);
xnor U19776 (N_19776,N_19504,N_19462);
and U19777 (N_19777,N_19589,N_19441);
xor U19778 (N_19778,N_19589,N_19536);
xor U19779 (N_19779,N_19502,N_19517);
and U19780 (N_19780,N_19535,N_19486);
and U19781 (N_19781,N_19540,N_19494);
nor U19782 (N_19782,N_19596,N_19560);
xor U19783 (N_19783,N_19549,N_19582);
or U19784 (N_19784,N_19596,N_19460);
or U19785 (N_19785,N_19546,N_19499);
nand U19786 (N_19786,N_19563,N_19460);
xnor U19787 (N_19787,N_19486,N_19577);
and U19788 (N_19788,N_19496,N_19560);
xor U19789 (N_19789,N_19576,N_19458);
nand U19790 (N_19790,N_19507,N_19523);
and U19791 (N_19791,N_19428,N_19408);
or U19792 (N_19792,N_19438,N_19460);
xnor U19793 (N_19793,N_19551,N_19505);
nor U19794 (N_19794,N_19544,N_19454);
xor U19795 (N_19795,N_19597,N_19590);
and U19796 (N_19796,N_19462,N_19465);
nand U19797 (N_19797,N_19475,N_19481);
xnor U19798 (N_19798,N_19435,N_19481);
nand U19799 (N_19799,N_19537,N_19556);
or U19800 (N_19800,N_19640,N_19781);
nor U19801 (N_19801,N_19793,N_19641);
nand U19802 (N_19802,N_19647,N_19690);
and U19803 (N_19803,N_19736,N_19693);
nand U19804 (N_19804,N_19764,N_19623);
nor U19805 (N_19805,N_19710,N_19774);
nor U19806 (N_19806,N_19633,N_19709);
xor U19807 (N_19807,N_19691,N_19695);
and U19808 (N_19808,N_19632,N_19790);
nor U19809 (N_19809,N_19732,N_19605);
and U19810 (N_19810,N_19777,N_19752);
nand U19811 (N_19811,N_19608,N_19675);
nor U19812 (N_19812,N_19787,N_19775);
nand U19813 (N_19813,N_19614,N_19689);
nand U19814 (N_19814,N_19639,N_19666);
and U19815 (N_19815,N_19779,N_19656);
nand U19816 (N_19816,N_19663,N_19621);
or U19817 (N_19817,N_19660,N_19626);
and U19818 (N_19818,N_19734,N_19701);
nand U19819 (N_19819,N_19707,N_19763);
nor U19820 (N_19820,N_19737,N_19697);
and U19821 (N_19821,N_19791,N_19742);
or U19822 (N_19822,N_19622,N_19636);
nand U19823 (N_19823,N_19624,N_19783);
and U19824 (N_19824,N_19798,N_19699);
nor U19825 (N_19825,N_19661,N_19761);
xnor U19826 (N_19826,N_19718,N_19782);
and U19827 (N_19827,N_19756,N_19627);
nand U19828 (N_19828,N_19745,N_19744);
or U19829 (N_19829,N_19651,N_19601);
nor U19830 (N_19830,N_19754,N_19748);
nor U19831 (N_19831,N_19679,N_19658);
nand U19832 (N_19832,N_19746,N_19696);
xnor U19833 (N_19833,N_19673,N_19767);
and U19834 (N_19834,N_19616,N_19716);
or U19835 (N_19835,N_19676,N_19725);
nor U19836 (N_19836,N_19778,N_19794);
and U19837 (N_19837,N_19788,N_19770);
or U19838 (N_19838,N_19652,N_19719);
nor U19839 (N_19839,N_19740,N_19618);
xor U19840 (N_19840,N_19750,N_19708);
nor U19841 (N_19841,N_19796,N_19702);
or U19842 (N_19842,N_19706,N_19698);
nor U19843 (N_19843,N_19712,N_19692);
or U19844 (N_19844,N_19771,N_19721);
and U19845 (N_19845,N_19646,N_19635);
nand U19846 (N_19846,N_19600,N_19751);
and U19847 (N_19847,N_19776,N_19664);
nor U19848 (N_19848,N_19747,N_19773);
or U19849 (N_19849,N_19795,N_19681);
and U19850 (N_19850,N_19717,N_19680);
xor U19851 (N_19851,N_19602,N_19653);
nand U19852 (N_19852,N_19772,N_19685);
nand U19853 (N_19853,N_19606,N_19743);
or U19854 (N_19854,N_19667,N_19643);
and U19855 (N_19855,N_19769,N_19741);
and U19856 (N_19856,N_19759,N_19753);
nor U19857 (N_19857,N_19659,N_19728);
nor U19858 (N_19858,N_19611,N_19687);
and U19859 (N_19859,N_19784,N_19722);
nor U19860 (N_19860,N_19649,N_19713);
nor U19861 (N_19861,N_19671,N_19644);
nand U19862 (N_19862,N_19715,N_19637);
and U19863 (N_19863,N_19720,N_19762);
or U19864 (N_19864,N_19780,N_19688);
xnor U19865 (N_19865,N_19609,N_19645);
xor U19866 (N_19866,N_19631,N_19683);
nand U19867 (N_19867,N_19677,N_19765);
nand U19868 (N_19868,N_19657,N_19766);
nand U19869 (N_19869,N_19630,N_19655);
or U19870 (N_19870,N_19629,N_19755);
nor U19871 (N_19871,N_19704,N_19792);
nor U19872 (N_19872,N_19726,N_19738);
xnor U19873 (N_19873,N_19603,N_19604);
nand U19874 (N_19874,N_19768,N_19705);
and U19875 (N_19875,N_19799,N_19711);
nor U19876 (N_19876,N_19638,N_19615);
xnor U19877 (N_19877,N_19613,N_19634);
nor U19878 (N_19878,N_19723,N_19694);
nor U19879 (N_19879,N_19730,N_19731);
and U19880 (N_19880,N_19735,N_19654);
and U19881 (N_19881,N_19733,N_19672);
or U19882 (N_19882,N_19703,N_19686);
nor U19883 (N_19883,N_19758,N_19669);
nand U19884 (N_19884,N_19642,N_19665);
xnor U19885 (N_19885,N_19684,N_19724);
nand U19886 (N_19886,N_19650,N_19668);
or U19887 (N_19887,N_19625,N_19757);
and U19888 (N_19888,N_19674,N_19700);
and U19889 (N_19889,N_19648,N_19789);
nand U19890 (N_19890,N_19682,N_19714);
nand U19891 (N_19891,N_19797,N_19617);
nand U19892 (N_19892,N_19620,N_19760);
nor U19893 (N_19893,N_19662,N_19785);
nor U19894 (N_19894,N_19749,N_19628);
and U19895 (N_19895,N_19739,N_19619);
nand U19896 (N_19896,N_19670,N_19729);
nor U19897 (N_19897,N_19610,N_19727);
xnor U19898 (N_19898,N_19612,N_19786);
and U19899 (N_19899,N_19607,N_19678);
or U19900 (N_19900,N_19739,N_19646);
nand U19901 (N_19901,N_19741,N_19699);
nor U19902 (N_19902,N_19795,N_19621);
nand U19903 (N_19903,N_19651,N_19720);
and U19904 (N_19904,N_19731,N_19682);
nor U19905 (N_19905,N_19613,N_19632);
and U19906 (N_19906,N_19778,N_19726);
xnor U19907 (N_19907,N_19623,N_19669);
or U19908 (N_19908,N_19644,N_19701);
and U19909 (N_19909,N_19735,N_19731);
and U19910 (N_19910,N_19797,N_19683);
nand U19911 (N_19911,N_19769,N_19648);
xnor U19912 (N_19912,N_19603,N_19694);
nand U19913 (N_19913,N_19661,N_19646);
nand U19914 (N_19914,N_19627,N_19664);
nand U19915 (N_19915,N_19771,N_19637);
nor U19916 (N_19916,N_19785,N_19620);
or U19917 (N_19917,N_19748,N_19627);
xnor U19918 (N_19918,N_19673,N_19731);
nand U19919 (N_19919,N_19780,N_19773);
or U19920 (N_19920,N_19665,N_19617);
nand U19921 (N_19921,N_19788,N_19716);
or U19922 (N_19922,N_19780,N_19662);
nor U19923 (N_19923,N_19792,N_19630);
nor U19924 (N_19924,N_19779,N_19732);
xor U19925 (N_19925,N_19634,N_19619);
and U19926 (N_19926,N_19664,N_19758);
or U19927 (N_19927,N_19606,N_19699);
nand U19928 (N_19928,N_19724,N_19734);
nand U19929 (N_19929,N_19736,N_19742);
or U19930 (N_19930,N_19712,N_19750);
nand U19931 (N_19931,N_19610,N_19739);
nand U19932 (N_19932,N_19601,N_19711);
and U19933 (N_19933,N_19743,N_19642);
nand U19934 (N_19934,N_19795,N_19700);
xnor U19935 (N_19935,N_19660,N_19722);
and U19936 (N_19936,N_19765,N_19688);
nand U19937 (N_19937,N_19618,N_19667);
nor U19938 (N_19938,N_19665,N_19772);
nand U19939 (N_19939,N_19747,N_19669);
xnor U19940 (N_19940,N_19796,N_19767);
and U19941 (N_19941,N_19777,N_19766);
xnor U19942 (N_19942,N_19702,N_19750);
xor U19943 (N_19943,N_19613,N_19759);
or U19944 (N_19944,N_19671,N_19721);
or U19945 (N_19945,N_19673,N_19651);
nor U19946 (N_19946,N_19623,N_19771);
and U19947 (N_19947,N_19682,N_19746);
nor U19948 (N_19948,N_19716,N_19740);
xor U19949 (N_19949,N_19622,N_19646);
or U19950 (N_19950,N_19714,N_19783);
nor U19951 (N_19951,N_19697,N_19625);
and U19952 (N_19952,N_19673,N_19763);
xnor U19953 (N_19953,N_19647,N_19681);
nor U19954 (N_19954,N_19792,N_19600);
nor U19955 (N_19955,N_19750,N_19730);
xor U19956 (N_19956,N_19674,N_19789);
nor U19957 (N_19957,N_19621,N_19742);
and U19958 (N_19958,N_19780,N_19628);
or U19959 (N_19959,N_19667,N_19697);
xor U19960 (N_19960,N_19799,N_19724);
or U19961 (N_19961,N_19623,N_19785);
and U19962 (N_19962,N_19652,N_19613);
xor U19963 (N_19963,N_19710,N_19676);
or U19964 (N_19964,N_19638,N_19653);
nor U19965 (N_19965,N_19666,N_19616);
or U19966 (N_19966,N_19614,N_19643);
and U19967 (N_19967,N_19731,N_19687);
or U19968 (N_19968,N_19711,N_19665);
and U19969 (N_19969,N_19750,N_19630);
xor U19970 (N_19970,N_19655,N_19736);
or U19971 (N_19971,N_19798,N_19658);
nor U19972 (N_19972,N_19644,N_19780);
xnor U19973 (N_19973,N_19678,N_19787);
and U19974 (N_19974,N_19693,N_19710);
nor U19975 (N_19975,N_19765,N_19742);
xnor U19976 (N_19976,N_19741,N_19607);
and U19977 (N_19977,N_19669,N_19765);
and U19978 (N_19978,N_19714,N_19603);
or U19979 (N_19979,N_19697,N_19727);
or U19980 (N_19980,N_19705,N_19726);
nand U19981 (N_19981,N_19759,N_19713);
nor U19982 (N_19982,N_19736,N_19689);
nor U19983 (N_19983,N_19762,N_19733);
nor U19984 (N_19984,N_19666,N_19769);
nand U19985 (N_19985,N_19643,N_19606);
and U19986 (N_19986,N_19640,N_19706);
xnor U19987 (N_19987,N_19785,N_19631);
and U19988 (N_19988,N_19739,N_19673);
nor U19989 (N_19989,N_19624,N_19754);
xnor U19990 (N_19990,N_19716,N_19753);
xnor U19991 (N_19991,N_19602,N_19690);
or U19992 (N_19992,N_19693,N_19780);
and U19993 (N_19993,N_19642,N_19797);
nand U19994 (N_19994,N_19688,N_19794);
nand U19995 (N_19995,N_19625,N_19715);
and U19996 (N_19996,N_19600,N_19648);
nand U19997 (N_19997,N_19775,N_19638);
or U19998 (N_19998,N_19730,N_19767);
nor U19999 (N_19999,N_19754,N_19717);
nand U20000 (N_20000,N_19911,N_19977);
and U20001 (N_20001,N_19863,N_19907);
or U20002 (N_20002,N_19832,N_19898);
xnor U20003 (N_20003,N_19974,N_19865);
nand U20004 (N_20004,N_19846,N_19842);
nor U20005 (N_20005,N_19983,N_19910);
xor U20006 (N_20006,N_19932,N_19915);
nor U20007 (N_20007,N_19858,N_19962);
nand U20008 (N_20008,N_19945,N_19881);
or U20009 (N_20009,N_19871,N_19981);
nand U20010 (N_20010,N_19990,N_19987);
nand U20011 (N_20011,N_19892,N_19928);
nor U20012 (N_20012,N_19843,N_19994);
or U20013 (N_20013,N_19817,N_19824);
and U20014 (N_20014,N_19938,N_19851);
xor U20015 (N_20015,N_19922,N_19968);
nand U20016 (N_20016,N_19982,N_19804);
nor U20017 (N_20017,N_19921,N_19926);
nand U20018 (N_20018,N_19836,N_19813);
xor U20019 (N_20019,N_19805,N_19976);
xnor U20020 (N_20020,N_19855,N_19985);
or U20021 (N_20021,N_19853,N_19908);
nand U20022 (N_20022,N_19952,N_19848);
or U20023 (N_20023,N_19943,N_19902);
or U20024 (N_20024,N_19829,N_19859);
and U20025 (N_20025,N_19850,N_19840);
or U20026 (N_20026,N_19978,N_19884);
nand U20027 (N_20027,N_19866,N_19991);
xor U20028 (N_20028,N_19827,N_19870);
and U20029 (N_20029,N_19988,N_19946);
nand U20030 (N_20030,N_19961,N_19971);
xor U20031 (N_20031,N_19935,N_19862);
nand U20032 (N_20032,N_19839,N_19880);
xor U20033 (N_20033,N_19960,N_19888);
or U20034 (N_20034,N_19822,N_19959);
and U20035 (N_20035,N_19833,N_19802);
nand U20036 (N_20036,N_19944,N_19820);
or U20037 (N_20037,N_19901,N_19891);
nand U20038 (N_20038,N_19807,N_19984);
and U20039 (N_20039,N_19861,N_19810);
or U20040 (N_20040,N_19919,N_19890);
xor U20041 (N_20041,N_19951,N_19803);
or U20042 (N_20042,N_19864,N_19996);
nor U20043 (N_20043,N_19999,N_19811);
and U20044 (N_20044,N_19818,N_19878);
xor U20045 (N_20045,N_19877,N_19808);
nand U20046 (N_20046,N_19812,N_19847);
xnor U20047 (N_20047,N_19947,N_19967);
or U20048 (N_20048,N_19950,N_19815);
xnor U20049 (N_20049,N_19954,N_19949);
or U20050 (N_20050,N_19966,N_19916);
and U20051 (N_20051,N_19904,N_19939);
nand U20052 (N_20052,N_19800,N_19831);
xor U20053 (N_20053,N_19814,N_19889);
or U20054 (N_20054,N_19972,N_19887);
or U20055 (N_20055,N_19912,N_19895);
nor U20056 (N_20056,N_19975,N_19809);
nand U20057 (N_20057,N_19899,N_19992);
nand U20058 (N_20058,N_19868,N_19825);
xnor U20059 (N_20059,N_19924,N_19925);
xor U20060 (N_20060,N_19823,N_19828);
and U20061 (N_20061,N_19874,N_19964);
nand U20062 (N_20062,N_19906,N_19980);
and U20063 (N_20063,N_19849,N_19927);
and U20064 (N_20064,N_19869,N_19821);
and U20065 (N_20065,N_19860,N_19963);
nand U20066 (N_20066,N_19893,N_19897);
or U20067 (N_20067,N_19937,N_19979);
nand U20068 (N_20068,N_19956,N_19886);
and U20069 (N_20069,N_19896,N_19857);
xor U20070 (N_20070,N_19969,N_19883);
nand U20071 (N_20071,N_19905,N_19918);
and U20072 (N_20072,N_19929,N_19819);
and U20073 (N_20073,N_19852,N_19955);
and U20074 (N_20074,N_19993,N_19838);
or U20075 (N_20075,N_19933,N_19894);
or U20076 (N_20076,N_19917,N_19854);
nor U20077 (N_20077,N_19885,N_19873);
nor U20078 (N_20078,N_19806,N_19882);
and U20079 (N_20079,N_19875,N_19934);
or U20080 (N_20080,N_19948,N_19970);
or U20081 (N_20081,N_19930,N_19923);
and U20082 (N_20082,N_19989,N_19953);
or U20083 (N_20083,N_19997,N_19998);
nor U20084 (N_20084,N_19872,N_19973);
xnor U20085 (N_20085,N_19913,N_19826);
nor U20086 (N_20086,N_19995,N_19986);
or U20087 (N_20087,N_19936,N_19834);
and U20088 (N_20088,N_19942,N_19958);
nand U20089 (N_20089,N_19801,N_19844);
nand U20090 (N_20090,N_19835,N_19957);
or U20091 (N_20091,N_19867,N_19941);
nand U20092 (N_20092,N_19914,N_19900);
nand U20093 (N_20093,N_19841,N_19931);
nor U20094 (N_20094,N_19920,N_19940);
and U20095 (N_20095,N_19856,N_19845);
nor U20096 (N_20096,N_19837,N_19816);
nand U20097 (N_20097,N_19876,N_19830);
and U20098 (N_20098,N_19903,N_19965);
and U20099 (N_20099,N_19909,N_19879);
nor U20100 (N_20100,N_19898,N_19869);
nor U20101 (N_20101,N_19962,N_19853);
nand U20102 (N_20102,N_19833,N_19917);
xnor U20103 (N_20103,N_19930,N_19811);
and U20104 (N_20104,N_19994,N_19802);
nor U20105 (N_20105,N_19899,N_19859);
or U20106 (N_20106,N_19860,N_19869);
nor U20107 (N_20107,N_19912,N_19862);
and U20108 (N_20108,N_19865,N_19960);
and U20109 (N_20109,N_19902,N_19934);
nor U20110 (N_20110,N_19856,N_19832);
or U20111 (N_20111,N_19825,N_19889);
nand U20112 (N_20112,N_19977,N_19954);
nor U20113 (N_20113,N_19924,N_19819);
and U20114 (N_20114,N_19926,N_19835);
or U20115 (N_20115,N_19844,N_19936);
nand U20116 (N_20116,N_19838,N_19971);
or U20117 (N_20117,N_19832,N_19957);
or U20118 (N_20118,N_19937,N_19810);
or U20119 (N_20119,N_19949,N_19922);
or U20120 (N_20120,N_19903,N_19850);
xor U20121 (N_20121,N_19821,N_19806);
xor U20122 (N_20122,N_19995,N_19937);
or U20123 (N_20123,N_19961,N_19822);
nor U20124 (N_20124,N_19930,N_19835);
and U20125 (N_20125,N_19837,N_19951);
xor U20126 (N_20126,N_19982,N_19850);
and U20127 (N_20127,N_19965,N_19822);
or U20128 (N_20128,N_19979,N_19840);
and U20129 (N_20129,N_19899,N_19837);
nor U20130 (N_20130,N_19957,N_19947);
nand U20131 (N_20131,N_19878,N_19874);
nand U20132 (N_20132,N_19930,N_19810);
nand U20133 (N_20133,N_19897,N_19956);
and U20134 (N_20134,N_19928,N_19976);
or U20135 (N_20135,N_19895,N_19840);
xnor U20136 (N_20136,N_19842,N_19852);
nor U20137 (N_20137,N_19905,N_19896);
xnor U20138 (N_20138,N_19801,N_19892);
nor U20139 (N_20139,N_19886,N_19835);
xor U20140 (N_20140,N_19920,N_19988);
or U20141 (N_20141,N_19934,N_19879);
nor U20142 (N_20142,N_19955,N_19850);
nand U20143 (N_20143,N_19810,N_19927);
nand U20144 (N_20144,N_19891,N_19985);
and U20145 (N_20145,N_19908,N_19971);
nand U20146 (N_20146,N_19816,N_19812);
and U20147 (N_20147,N_19973,N_19918);
nand U20148 (N_20148,N_19822,N_19823);
or U20149 (N_20149,N_19800,N_19822);
or U20150 (N_20150,N_19885,N_19923);
and U20151 (N_20151,N_19964,N_19906);
and U20152 (N_20152,N_19822,N_19884);
nor U20153 (N_20153,N_19915,N_19838);
xnor U20154 (N_20154,N_19884,N_19962);
xnor U20155 (N_20155,N_19865,N_19901);
nor U20156 (N_20156,N_19898,N_19878);
xnor U20157 (N_20157,N_19888,N_19861);
xor U20158 (N_20158,N_19927,N_19835);
and U20159 (N_20159,N_19923,N_19962);
and U20160 (N_20160,N_19960,N_19935);
and U20161 (N_20161,N_19995,N_19999);
or U20162 (N_20162,N_19842,N_19923);
or U20163 (N_20163,N_19964,N_19977);
and U20164 (N_20164,N_19864,N_19846);
nand U20165 (N_20165,N_19870,N_19954);
or U20166 (N_20166,N_19931,N_19998);
and U20167 (N_20167,N_19852,N_19918);
or U20168 (N_20168,N_19992,N_19972);
nor U20169 (N_20169,N_19941,N_19939);
nor U20170 (N_20170,N_19910,N_19878);
and U20171 (N_20171,N_19910,N_19876);
and U20172 (N_20172,N_19972,N_19896);
or U20173 (N_20173,N_19999,N_19970);
nand U20174 (N_20174,N_19840,N_19911);
and U20175 (N_20175,N_19970,N_19862);
or U20176 (N_20176,N_19939,N_19993);
xor U20177 (N_20177,N_19971,N_19960);
nand U20178 (N_20178,N_19950,N_19833);
or U20179 (N_20179,N_19815,N_19838);
and U20180 (N_20180,N_19932,N_19865);
and U20181 (N_20181,N_19928,N_19934);
and U20182 (N_20182,N_19957,N_19874);
nand U20183 (N_20183,N_19802,N_19851);
and U20184 (N_20184,N_19822,N_19947);
xor U20185 (N_20185,N_19888,N_19979);
or U20186 (N_20186,N_19863,N_19914);
and U20187 (N_20187,N_19861,N_19864);
and U20188 (N_20188,N_19818,N_19931);
nor U20189 (N_20189,N_19917,N_19914);
nand U20190 (N_20190,N_19857,N_19877);
or U20191 (N_20191,N_19958,N_19902);
or U20192 (N_20192,N_19918,N_19878);
and U20193 (N_20193,N_19876,N_19955);
nand U20194 (N_20194,N_19904,N_19871);
nand U20195 (N_20195,N_19980,N_19907);
or U20196 (N_20196,N_19873,N_19933);
xnor U20197 (N_20197,N_19838,N_19943);
nor U20198 (N_20198,N_19988,N_19908);
or U20199 (N_20199,N_19967,N_19823);
nor U20200 (N_20200,N_20075,N_20007);
nor U20201 (N_20201,N_20164,N_20087);
nand U20202 (N_20202,N_20049,N_20023);
xnor U20203 (N_20203,N_20041,N_20010);
xnor U20204 (N_20204,N_20106,N_20163);
nand U20205 (N_20205,N_20191,N_20005);
nor U20206 (N_20206,N_20172,N_20099);
xor U20207 (N_20207,N_20004,N_20183);
nor U20208 (N_20208,N_20112,N_20174);
nand U20209 (N_20209,N_20159,N_20044);
nand U20210 (N_20210,N_20143,N_20134);
nand U20211 (N_20211,N_20131,N_20025);
nor U20212 (N_20212,N_20062,N_20119);
nand U20213 (N_20213,N_20029,N_20127);
nand U20214 (N_20214,N_20167,N_20192);
nand U20215 (N_20215,N_20126,N_20154);
or U20216 (N_20216,N_20080,N_20083);
nor U20217 (N_20217,N_20050,N_20196);
nand U20218 (N_20218,N_20139,N_20036);
nor U20219 (N_20219,N_20101,N_20030);
nand U20220 (N_20220,N_20130,N_20078);
and U20221 (N_20221,N_20000,N_20152);
or U20222 (N_20222,N_20091,N_20058);
nor U20223 (N_20223,N_20012,N_20182);
nor U20224 (N_20224,N_20002,N_20125);
nor U20225 (N_20225,N_20055,N_20117);
nand U20226 (N_20226,N_20035,N_20177);
or U20227 (N_20227,N_20198,N_20063);
xor U20228 (N_20228,N_20129,N_20011);
nand U20229 (N_20229,N_20077,N_20047);
xnor U20230 (N_20230,N_20060,N_20095);
nor U20231 (N_20231,N_20024,N_20020);
nand U20232 (N_20232,N_20108,N_20179);
nand U20233 (N_20233,N_20115,N_20169);
and U20234 (N_20234,N_20039,N_20155);
xnor U20235 (N_20235,N_20145,N_20079);
or U20236 (N_20236,N_20040,N_20071);
nand U20237 (N_20237,N_20031,N_20181);
or U20238 (N_20238,N_20034,N_20017);
xor U20239 (N_20239,N_20173,N_20180);
and U20240 (N_20240,N_20133,N_20138);
nand U20241 (N_20241,N_20082,N_20001);
nor U20242 (N_20242,N_20021,N_20072);
xnor U20243 (N_20243,N_20161,N_20042);
or U20244 (N_20244,N_20160,N_20088);
nand U20245 (N_20245,N_20136,N_20140);
or U20246 (N_20246,N_20018,N_20090);
and U20247 (N_20247,N_20059,N_20027);
or U20248 (N_20248,N_20051,N_20195);
or U20249 (N_20249,N_20084,N_20066);
and U20250 (N_20250,N_20046,N_20003);
xnor U20251 (N_20251,N_20188,N_20199);
nand U20252 (N_20252,N_20067,N_20038);
nor U20253 (N_20253,N_20022,N_20093);
xnor U20254 (N_20254,N_20086,N_20026);
nand U20255 (N_20255,N_20185,N_20081);
and U20256 (N_20256,N_20132,N_20114);
xor U20257 (N_20257,N_20054,N_20176);
nand U20258 (N_20258,N_20110,N_20121);
or U20259 (N_20259,N_20171,N_20118);
or U20260 (N_20260,N_20057,N_20184);
xnor U20261 (N_20261,N_20070,N_20149);
xnor U20262 (N_20262,N_20197,N_20098);
xnor U20263 (N_20263,N_20168,N_20170);
and U20264 (N_20264,N_20105,N_20104);
xnor U20265 (N_20265,N_20189,N_20089);
nand U20266 (N_20266,N_20153,N_20151);
and U20267 (N_20267,N_20096,N_20165);
nor U20268 (N_20268,N_20056,N_20146);
xnor U20269 (N_20269,N_20009,N_20094);
nand U20270 (N_20270,N_20064,N_20113);
and U20271 (N_20271,N_20085,N_20019);
nor U20272 (N_20272,N_20137,N_20068);
nor U20273 (N_20273,N_20156,N_20178);
nor U20274 (N_20274,N_20037,N_20193);
nor U20275 (N_20275,N_20016,N_20013);
or U20276 (N_20276,N_20190,N_20045);
nand U20277 (N_20277,N_20158,N_20076);
nand U20278 (N_20278,N_20128,N_20141);
or U20279 (N_20279,N_20175,N_20074);
or U20280 (N_20280,N_20150,N_20166);
nand U20281 (N_20281,N_20048,N_20102);
and U20282 (N_20282,N_20028,N_20015);
nor U20283 (N_20283,N_20135,N_20186);
nand U20284 (N_20284,N_20073,N_20032);
xnor U20285 (N_20285,N_20157,N_20103);
nor U20286 (N_20286,N_20187,N_20109);
xnor U20287 (N_20287,N_20124,N_20194);
nand U20288 (N_20288,N_20120,N_20008);
nand U20289 (N_20289,N_20043,N_20052);
xnor U20290 (N_20290,N_20061,N_20006);
nand U20291 (N_20291,N_20097,N_20147);
xor U20292 (N_20292,N_20092,N_20142);
or U20293 (N_20293,N_20014,N_20123);
nor U20294 (N_20294,N_20122,N_20162);
or U20295 (N_20295,N_20053,N_20148);
nand U20296 (N_20296,N_20065,N_20107);
xor U20297 (N_20297,N_20033,N_20144);
or U20298 (N_20298,N_20069,N_20116);
nand U20299 (N_20299,N_20100,N_20111);
nor U20300 (N_20300,N_20079,N_20069);
and U20301 (N_20301,N_20020,N_20132);
and U20302 (N_20302,N_20069,N_20016);
nand U20303 (N_20303,N_20089,N_20114);
nor U20304 (N_20304,N_20185,N_20048);
nand U20305 (N_20305,N_20118,N_20181);
nor U20306 (N_20306,N_20006,N_20040);
and U20307 (N_20307,N_20146,N_20195);
nor U20308 (N_20308,N_20186,N_20166);
xnor U20309 (N_20309,N_20195,N_20138);
and U20310 (N_20310,N_20124,N_20081);
xnor U20311 (N_20311,N_20140,N_20119);
xor U20312 (N_20312,N_20070,N_20169);
nor U20313 (N_20313,N_20196,N_20034);
and U20314 (N_20314,N_20092,N_20000);
nand U20315 (N_20315,N_20080,N_20118);
and U20316 (N_20316,N_20037,N_20067);
xor U20317 (N_20317,N_20158,N_20090);
nand U20318 (N_20318,N_20149,N_20109);
xnor U20319 (N_20319,N_20179,N_20000);
xor U20320 (N_20320,N_20064,N_20166);
nor U20321 (N_20321,N_20074,N_20003);
nand U20322 (N_20322,N_20092,N_20007);
and U20323 (N_20323,N_20133,N_20161);
or U20324 (N_20324,N_20081,N_20169);
or U20325 (N_20325,N_20076,N_20016);
nand U20326 (N_20326,N_20073,N_20117);
and U20327 (N_20327,N_20184,N_20163);
nand U20328 (N_20328,N_20127,N_20191);
nand U20329 (N_20329,N_20024,N_20160);
xnor U20330 (N_20330,N_20000,N_20108);
and U20331 (N_20331,N_20058,N_20165);
and U20332 (N_20332,N_20084,N_20192);
xor U20333 (N_20333,N_20032,N_20059);
xor U20334 (N_20334,N_20046,N_20111);
and U20335 (N_20335,N_20138,N_20135);
or U20336 (N_20336,N_20083,N_20132);
and U20337 (N_20337,N_20085,N_20181);
nor U20338 (N_20338,N_20131,N_20146);
nor U20339 (N_20339,N_20165,N_20086);
nand U20340 (N_20340,N_20074,N_20041);
nor U20341 (N_20341,N_20102,N_20181);
and U20342 (N_20342,N_20123,N_20167);
nor U20343 (N_20343,N_20134,N_20181);
xor U20344 (N_20344,N_20006,N_20092);
nand U20345 (N_20345,N_20140,N_20029);
nor U20346 (N_20346,N_20050,N_20068);
nand U20347 (N_20347,N_20081,N_20059);
xnor U20348 (N_20348,N_20108,N_20089);
or U20349 (N_20349,N_20010,N_20045);
xor U20350 (N_20350,N_20171,N_20019);
nand U20351 (N_20351,N_20084,N_20089);
xor U20352 (N_20352,N_20105,N_20037);
xor U20353 (N_20353,N_20051,N_20178);
nor U20354 (N_20354,N_20074,N_20019);
xor U20355 (N_20355,N_20127,N_20159);
nor U20356 (N_20356,N_20194,N_20193);
nand U20357 (N_20357,N_20125,N_20111);
nand U20358 (N_20358,N_20072,N_20027);
nor U20359 (N_20359,N_20009,N_20132);
nand U20360 (N_20360,N_20009,N_20096);
nor U20361 (N_20361,N_20054,N_20067);
and U20362 (N_20362,N_20025,N_20105);
nor U20363 (N_20363,N_20021,N_20034);
xor U20364 (N_20364,N_20123,N_20105);
nor U20365 (N_20365,N_20196,N_20132);
or U20366 (N_20366,N_20141,N_20058);
nand U20367 (N_20367,N_20145,N_20118);
nor U20368 (N_20368,N_20006,N_20119);
xnor U20369 (N_20369,N_20030,N_20140);
or U20370 (N_20370,N_20104,N_20087);
and U20371 (N_20371,N_20174,N_20107);
nand U20372 (N_20372,N_20043,N_20003);
xor U20373 (N_20373,N_20048,N_20134);
nor U20374 (N_20374,N_20176,N_20168);
nor U20375 (N_20375,N_20092,N_20131);
or U20376 (N_20376,N_20045,N_20193);
nand U20377 (N_20377,N_20043,N_20125);
or U20378 (N_20378,N_20161,N_20129);
nor U20379 (N_20379,N_20096,N_20052);
and U20380 (N_20380,N_20169,N_20162);
and U20381 (N_20381,N_20027,N_20160);
or U20382 (N_20382,N_20145,N_20067);
or U20383 (N_20383,N_20039,N_20068);
xnor U20384 (N_20384,N_20183,N_20039);
or U20385 (N_20385,N_20126,N_20170);
nor U20386 (N_20386,N_20123,N_20099);
and U20387 (N_20387,N_20105,N_20143);
xnor U20388 (N_20388,N_20063,N_20161);
nor U20389 (N_20389,N_20042,N_20048);
xor U20390 (N_20390,N_20146,N_20173);
or U20391 (N_20391,N_20141,N_20171);
xnor U20392 (N_20392,N_20166,N_20105);
or U20393 (N_20393,N_20031,N_20005);
or U20394 (N_20394,N_20197,N_20142);
nand U20395 (N_20395,N_20142,N_20079);
nor U20396 (N_20396,N_20087,N_20194);
or U20397 (N_20397,N_20133,N_20077);
and U20398 (N_20398,N_20162,N_20161);
or U20399 (N_20399,N_20183,N_20106);
or U20400 (N_20400,N_20264,N_20388);
or U20401 (N_20401,N_20378,N_20320);
nand U20402 (N_20402,N_20216,N_20255);
nand U20403 (N_20403,N_20376,N_20251);
nand U20404 (N_20404,N_20291,N_20287);
nor U20405 (N_20405,N_20288,N_20217);
nand U20406 (N_20406,N_20286,N_20235);
xor U20407 (N_20407,N_20354,N_20219);
and U20408 (N_20408,N_20359,N_20360);
or U20409 (N_20409,N_20230,N_20395);
nor U20410 (N_20410,N_20386,N_20365);
xor U20411 (N_20411,N_20331,N_20348);
xor U20412 (N_20412,N_20353,N_20200);
nand U20413 (N_20413,N_20220,N_20275);
nor U20414 (N_20414,N_20299,N_20390);
and U20415 (N_20415,N_20269,N_20345);
or U20416 (N_20416,N_20308,N_20284);
nand U20417 (N_20417,N_20322,N_20392);
nor U20418 (N_20418,N_20270,N_20384);
and U20419 (N_20419,N_20358,N_20207);
xor U20420 (N_20420,N_20243,N_20257);
xnor U20421 (N_20421,N_20351,N_20326);
nor U20422 (N_20422,N_20215,N_20300);
and U20423 (N_20423,N_20250,N_20206);
and U20424 (N_20424,N_20314,N_20312);
xor U20425 (N_20425,N_20245,N_20328);
nand U20426 (N_20426,N_20397,N_20349);
and U20427 (N_20427,N_20362,N_20285);
nor U20428 (N_20428,N_20262,N_20315);
and U20429 (N_20429,N_20234,N_20325);
nand U20430 (N_20430,N_20382,N_20339);
nand U20431 (N_20431,N_20311,N_20398);
nor U20432 (N_20432,N_20294,N_20394);
nor U20433 (N_20433,N_20340,N_20265);
or U20434 (N_20434,N_20272,N_20356);
nand U20435 (N_20435,N_20327,N_20304);
xor U20436 (N_20436,N_20347,N_20253);
nor U20437 (N_20437,N_20364,N_20301);
xnor U20438 (N_20438,N_20307,N_20346);
nand U20439 (N_20439,N_20361,N_20377);
nor U20440 (N_20440,N_20324,N_20278);
xor U20441 (N_20441,N_20256,N_20369);
nor U20442 (N_20442,N_20259,N_20247);
or U20443 (N_20443,N_20231,N_20309);
or U20444 (N_20444,N_20252,N_20204);
xnor U20445 (N_20445,N_20292,N_20274);
nor U20446 (N_20446,N_20332,N_20375);
nor U20447 (N_20447,N_20336,N_20289);
xnor U20448 (N_20448,N_20306,N_20226);
xnor U20449 (N_20449,N_20316,N_20258);
and U20450 (N_20450,N_20303,N_20203);
and U20451 (N_20451,N_20225,N_20380);
nor U20452 (N_20452,N_20233,N_20281);
and U20453 (N_20453,N_20260,N_20343);
nor U20454 (N_20454,N_20205,N_20367);
nand U20455 (N_20455,N_20282,N_20271);
and U20456 (N_20456,N_20268,N_20244);
nor U20457 (N_20457,N_20273,N_20222);
nand U20458 (N_20458,N_20279,N_20373);
nor U20459 (N_20459,N_20391,N_20333);
xnor U20460 (N_20460,N_20341,N_20210);
nor U20461 (N_20461,N_20298,N_20218);
and U20462 (N_20462,N_20385,N_20280);
and U20463 (N_20463,N_20379,N_20383);
and U20464 (N_20464,N_20357,N_20393);
or U20465 (N_20465,N_20370,N_20318);
nand U20466 (N_20466,N_20329,N_20371);
nand U20467 (N_20467,N_20366,N_20229);
xnor U20468 (N_20468,N_20236,N_20302);
xor U20469 (N_20469,N_20232,N_20399);
or U20470 (N_20470,N_20323,N_20290);
nand U20471 (N_20471,N_20223,N_20317);
nand U20472 (N_20472,N_20296,N_20240);
and U20473 (N_20473,N_20335,N_20254);
xnor U20474 (N_20474,N_20212,N_20267);
and U20475 (N_20475,N_20350,N_20224);
nand U20476 (N_20476,N_20237,N_20368);
nand U20477 (N_20477,N_20246,N_20330);
nand U20478 (N_20478,N_20201,N_20313);
or U20479 (N_20479,N_20305,N_20372);
or U20480 (N_20480,N_20261,N_20293);
or U20481 (N_20481,N_20310,N_20342);
or U20482 (N_20482,N_20213,N_20277);
nand U20483 (N_20483,N_20297,N_20239);
xor U20484 (N_20484,N_20266,N_20338);
or U20485 (N_20485,N_20295,N_20276);
nor U20486 (N_20486,N_20248,N_20214);
and U20487 (N_20487,N_20321,N_20283);
nand U20488 (N_20488,N_20352,N_20334);
or U20489 (N_20489,N_20228,N_20249);
or U20490 (N_20490,N_20337,N_20263);
nor U20491 (N_20491,N_20242,N_20344);
nand U20492 (N_20492,N_20238,N_20211);
and U20493 (N_20493,N_20227,N_20241);
or U20494 (N_20494,N_20355,N_20221);
or U20495 (N_20495,N_20209,N_20374);
or U20496 (N_20496,N_20389,N_20363);
xnor U20497 (N_20497,N_20319,N_20208);
nand U20498 (N_20498,N_20396,N_20387);
xor U20499 (N_20499,N_20202,N_20381);
or U20500 (N_20500,N_20285,N_20264);
nor U20501 (N_20501,N_20367,N_20236);
xor U20502 (N_20502,N_20243,N_20332);
nand U20503 (N_20503,N_20278,N_20274);
xnor U20504 (N_20504,N_20398,N_20249);
and U20505 (N_20505,N_20295,N_20265);
nor U20506 (N_20506,N_20391,N_20358);
nand U20507 (N_20507,N_20299,N_20350);
nor U20508 (N_20508,N_20335,N_20337);
nor U20509 (N_20509,N_20333,N_20336);
nor U20510 (N_20510,N_20346,N_20398);
nor U20511 (N_20511,N_20241,N_20333);
xnor U20512 (N_20512,N_20279,N_20231);
nor U20513 (N_20513,N_20224,N_20365);
and U20514 (N_20514,N_20381,N_20271);
nor U20515 (N_20515,N_20328,N_20252);
xnor U20516 (N_20516,N_20305,N_20348);
nand U20517 (N_20517,N_20360,N_20328);
xnor U20518 (N_20518,N_20226,N_20297);
nand U20519 (N_20519,N_20233,N_20259);
nor U20520 (N_20520,N_20264,N_20386);
nor U20521 (N_20521,N_20320,N_20297);
nor U20522 (N_20522,N_20255,N_20353);
or U20523 (N_20523,N_20369,N_20380);
nand U20524 (N_20524,N_20277,N_20327);
and U20525 (N_20525,N_20295,N_20317);
and U20526 (N_20526,N_20308,N_20382);
nor U20527 (N_20527,N_20242,N_20365);
nor U20528 (N_20528,N_20346,N_20255);
nand U20529 (N_20529,N_20328,N_20359);
nand U20530 (N_20530,N_20379,N_20201);
xor U20531 (N_20531,N_20264,N_20279);
or U20532 (N_20532,N_20246,N_20299);
nor U20533 (N_20533,N_20220,N_20399);
and U20534 (N_20534,N_20215,N_20287);
nor U20535 (N_20535,N_20287,N_20381);
nor U20536 (N_20536,N_20207,N_20222);
and U20537 (N_20537,N_20272,N_20390);
nor U20538 (N_20538,N_20222,N_20352);
and U20539 (N_20539,N_20307,N_20239);
nand U20540 (N_20540,N_20330,N_20393);
or U20541 (N_20541,N_20268,N_20201);
or U20542 (N_20542,N_20343,N_20259);
nor U20543 (N_20543,N_20315,N_20368);
nor U20544 (N_20544,N_20211,N_20232);
or U20545 (N_20545,N_20348,N_20221);
and U20546 (N_20546,N_20255,N_20288);
xnor U20547 (N_20547,N_20285,N_20273);
nand U20548 (N_20548,N_20266,N_20309);
nand U20549 (N_20549,N_20272,N_20269);
or U20550 (N_20550,N_20343,N_20299);
nor U20551 (N_20551,N_20334,N_20381);
nand U20552 (N_20552,N_20309,N_20326);
and U20553 (N_20553,N_20276,N_20209);
and U20554 (N_20554,N_20398,N_20310);
and U20555 (N_20555,N_20366,N_20296);
or U20556 (N_20556,N_20305,N_20294);
or U20557 (N_20557,N_20399,N_20344);
nor U20558 (N_20558,N_20366,N_20212);
nor U20559 (N_20559,N_20335,N_20212);
and U20560 (N_20560,N_20224,N_20201);
nand U20561 (N_20561,N_20391,N_20292);
and U20562 (N_20562,N_20381,N_20352);
and U20563 (N_20563,N_20366,N_20379);
nor U20564 (N_20564,N_20254,N_20238);
nor U20565 (N_20565,N_20202,N_20375);
xnor U20566 (N_20566,N_20359,N_20299);
nor U20567 (N_20567,N_20393,N_20305);
nor U20568 (N_20568,N_20220,N_20226);
or U20569 (N_20569,N_20362,N_20373);
xnor U20570 (N_20570,N_20230,N_20265);
xnor U20571 (N_20571,N_20378,N_20297);
and U20572 (N_20572,N_20255,N_20253);
nor U20573 (N_20573,N_20397,N_20331);
xor U20574 (N_20574,N_20342,N_20341);
or U20575 (N_20575,N_20370,N_20222);
nand U20576 (N_20576,N_20354,N_20355);
and U20577 (N_20577,N_20283,N_20335);
xnor U20578 (N_20578,N_20275,N_20387);
or U20579 (N_20579,N_20356,N_20252);
or U20580 (N_20580,N_20317,N_20208);
xor U20581 (N_20581,N_20380,N_20253);
and U20582 (N_20582,N_20273,N_20201);
or U20583 (N_20583,N_20388,N_20372);
or U20584 (N_20584,N_20357,N_20325);
nor U20585 (N_20585,N_20315,N_20380);
or U20586 (N_20586,N_20348,N_20372);
and U20587 (N_20587,N_20239,N_20217);
nand U20588 (N_20588,N_20241,N_20266);
nand U20589 (N_20589,N_20334,N_20290);
or U20590 (N_20590,N_20357,N_20391);
nor U20591 (N_20591,N_20244,N_20284);
or U20592 (N_20592,N_20253,N_20343);
or U20593 (N_20593,N_20292,N_20315);
and U20594 (N_20594,N_20373,N_20345);
xor U20595 (N_20595,N_20346,N_20205);
and U20596 (N_20596,N_20361,N_20278);
and U20597 (N_20597,N_20379,N_20355);
and U20598 (N_20598,N_20294,N_20369);
and U20599 (N_20599,N_20295,N_20282);
and U20600 (N_20600,N_20400,N_20440);
nand U20601 (N_20601,N_20490,N_20423);
nand U20602 (N_20602,N_20510,N_20596);
nand U20603 (N_20603,N_20404,N_20581);
xor U20604 (N_20604,N_20543,N_20557);
nor U20605 (N_20605,N_20410,N_20413);
and U20606 (N_20606,N_20443,N_20494);
xnor U20607 (N_20607,N_20473,N_20564);
nand U20608 (N_20608,N_20480,N_20548);
xor U20609 (N_20609,N_20587,N_20426);
xnor U20610 (N_20610,N_20445,N_20512);
and U20611 (N_20611,N_20500,N_20477);
nor U20612 (N_20612,N_20537,N_20415);
nor U20613 (N_20613,N_20536,N_20460);
nand U20614 (N_20614,N_20567,N_20449);
or U20615 (N_20615,N_20513,N_20552);
nand U20616 (N_20616,N_20458,N_20503);
or U20617 (N_20617,N_20402,N_20424);
nand U20618 (N_20618,N_20556,N_20565);
or U20619 (N_20619,N_20527,N_20493);
xnor U20620 (N_20620,N_20584,N_20588);
and U20621 (N_20621,N_20511,N_20519);
and U20622 (N_20622,N_20482,N_20474);
or U20623 (N_20623,N_20592,N_20535);
or U20624 (N_20624,N_20574,N_20428);
nor U20625 (N_20625,N_20419,N_20521);
xor U20626 (N_20626,N_20447,N_20448);
nand U20627 (N_20627,N_20444,N_20469);
and U20628 (N_20628,N_20522,N_20576);
nor U20629 (N_20629,N_20405,N_20439);
xnor U20630 (N_20630,N_20438,N_20485);
nor U20631 (N_20631,N_20463,N_20496);
nor U20632 (N_20632,N_20505,N_20590);
nor U20633 (N_20633,N_20561,N_20540);
nor U20634 (N_20634,N_20544,N_20579);
and U20635 (N_20635,N_20403,N_20499);
nand U20636 (N_20636,N_20491,N_20441);
and U20637 (N_20637,N_20433,N_20504);
nor U20638 (N_20638,N_20450,N_20572);
nor U20639 (N_20639,N_20578,N_20570);
nand U20640 (N_20640,N_20515,N_20597);
nor U20641 (N_20641,N_20516,N_20585);
nand U20642 (N_20642,N_20541,N_20569);
xor U20643 (N_20643,N_20435,N_20528);
nor U20644 (N_20644,N_20492,N_20429);
or U20645 (N_20645,N_20593,N_20401);
and U20646 (N_20646,N_20533,N_20420);
nor U20647 (N_20647,N_20451,N_20580);
nand U20648 (N_20648,N_20506,N_20560);
and U20649 (N_20649,N_20464,N_20408);
or U20650 (N_20650,N_20471,N_20598);
and U20651 (N_20651,N_20434,N_20425);
nand U20652 (N_20652,N_20465,N_20432);
or U20653 (N_20653,N_20509,N_20546);
nand U20654 (N_20654,N_20483,N_20455);
nor U20655 (N_20655,N_20411,N_20551);
xor U20656 (N_20656,N_20478,N_20530);
and U20657 (N_20657,N_20582,N_20472);
nand U20658 (N_20658,N_20542,N_20418);
nor U20659 (N_20659,N_20599,N_20436);
or U20660 (N_20660,N_20431,N_20550);
and U20661 (N_20661,N_20417,N_20422);
nor U20662 (N_20662,N_20442,N_20467);
xnor U20663 (N_20663,N_20547,N_20456);
nor U20664 (N_20664,N_20412,N_20575);
xnor U20665 (N_20665,N_20437,N_20476);
nor U20666 (N_20666,N_20414,N_20555);
or U20667 (N_20667,N_20487,N_20514);
or U20668 (N_20668,N_20534,N_20486);
nand U20669 (N_20669,N_20517,N_20508);
and U20670 (N_20670,N_20457,N_20497);
and U20671 (N_20671,N_20566,N_20571);
nor U20672 (N_20672,N_20454,N_20529);
or U20673 (N_20673,N_20518,N_20532);
xnor U20674 (N_20674,N_20531,N_20524);
nor U20675 (N_20675,N_20538,N_20452);
xnor U20676 (N_20676,N_20558,N_20525);
xnor U20677 (N_20677,N_20553,N_20591);
and U20678 (N_20678,N_20539,N_20583);
and U20679 (N_20679,N_20549,N_20520);
nor U20680 (N_20680,N_20554,N_20468);
nor U20681 (N_20681,N_20495,N_20523);
or U20682 (N_20682,N_20459,N_20416);
nand U20683 (N_20683,N_20479,N_20430);
xor U20684 (N_20684,N_20409,N_20507);
nand U20685 (N_20685,N_20545,N_20526);
nor U20686 (N_20686,N_20462,N_20577);
xor U20687 (N_20687,N_20421,N_20475);
or U20688 (N_20688,N_20501,N_20407);
nor U20689 (N_20689,N_20595,N_20466);
nand U20690 (N_20690,N_20461,N_20559);
and U20691 (N_20691,N_20589,N_20453);
xor U20692 (N_20692,N_20563,N_20446);
nand U20693 (N_20693,N_20470,N_20406);
and U20694 (N_20694,N_20573,N_20502);
nand U20695 (N_20695,N_20488,N_20427);
xnor U20696 (N_20696,N_20484,N_20489);
xnor U20697 (N_20697,N_20498,N_20586);
or U20698 (N_20698,N_20594,N_20568);
or U20699 (N_20699,N_20481,N_20562);
or U20700 (N_20700,N_20478,N_20579);
and U20701 (N_20701,N_20427,N_20532);
nor U20702 (N_20702,N_20534,N_20509);
nor U20703 (N_20703,N_20441,N_20429);
nor U20704 (N_20704,N_20497,N_20404);
nor U20705 (N_20705,N_20433,N_20517);
or U20706 (N_20706,N_20428,N_20464);
or U20707 (N_20707,N_20439,N_20564);
nand U20708 (N_20708,N_20565,N_20455);
nand U20709 (N_20709,N_20463,N_20594);
nand U20710 (N_20710,N_20514,N_20410);
xor U20711 (N_20711,N_20548,N_20467);
and U20712 (N_20712,N_20529,N_20561);
or U20713 (N_20713,N_20463,N_20558);
xor U20714 (N_20714,N_20471,N_20478);
or U20715 (N_20715,N_20426,N_20460);
or U20716 (N_20716,N_20548,N_20457);
nor U20717 (N_20717,N_20430,N_20429);
nor U20718 (N_20718,N_20513,N_20434);
and U20719 (N_20719,N_20565,N_20479);
nor U20720 (N_20720,N_20417,N_20479);
and U20721 (N_20721,N_20535,N_20445);
and U20722 (N_20722,N_20501,N_20512);
xnor U20723 (N_20723,N_20575,N_20555);
xnor U20724 (N_20724,N_20405,N_20442);
xor U20725 (N_20725,N_20448,N_20542);
nor U20726 (N_20726,N_20511,N_20442);
xnor U20727 (N_20727,N_20483,N_20519);
xor U20728 (N_20728,N_20528,N_20408);
nand U20729 (N_20729,N_20400,N_20453);
or U20730 (N_20730,N_20588,N_20408);
and U20731 (N_20731,N_20522,N_20456);
nand U20732 (N_20732,N_20582,N_20467);
or U20733 (N_20733,N_20418,N_20471);
nor U20734 (N_20734,N_20469,N_20459);
xnor U20735 (N_20735,N_20505,N_20506);
xnor U20736 (N_20736,N_20557,N_20431);
and U20737 (N_20737,N_20596,N_20468);
nor U20738 (N_20738,N_20432,N_20414);
and U20739 (N_20739,N_20439,N_20414);
and U20740 (N_20740,N_20574,N_20456);
nor U20741 (N_20741,N_20424,N_20513);
nand U20742 (N_20742,N_20416,N_20533);
or U20743 (N_20743,N_20519,N_20436);
or U20744 (N_20744,N_20401,N_20478);
nor U20745 (N_20745,N_20457,N_20597);
nor U20746 (N_20746,N_20442,N_20568);
xnor U20747 (N_20747,N_20422,N_20451);
nor U20748 (N_20748,N_20546,N_20573);
or U20749 (N_20749,N_20549,N_20450);
nor U20750 (N_20750,N_20486,N_20475);
or U20751 (N_20751,N_20552,N_20476);
or U20752 (N_20752,N_20486,N_20520);
xor U20753 (N_20753,N_20523,N_20414);
and U20754 (N_20754,N_20550,N_20475);
and U20755 (N_20755,N_20598,N_20457);
nor U20756 (N_20756,N_20566,N_20584);
or U20757 (N_20757,N_20405,N_20463);
nor U20758 (N_20758,N_20420,N_20441);
nor U20759 (N_20759,N_20477,N_20580);
and U20760 (N_20760,N_20568,N_20407);
and U20761 (N_20761,N_20559,N_20515);
and U20762 (N_20762,N_20496,N_20407);
nand U20763 (N_20763,N_20461,N_20540);
and U20764 (N_20764,N_20521,N_20427);
or U20765 (N_20765,N_20425,N_20532);
nor U20766 (N_20766,N_20523,N_20496);
nor U20767 (N_20767,N_20561,N_20553);
or U20768 (N_20768,N_20577,N_20435);
nand U20769 (N_20769,N_20526,N_20459);
nor U20770 (N_20770,N_20471,N_20422);
nand U20771 (N_20771,N_20403,N_20576);
xor U20772 (N_20772,N_20566,N_20515);
nor U20773 (N_20773,N_20509,N_20503);
xnor U20774 (N_20774,N_20444,N_20424);
nand U20775 (N_20775,N_20531,N_20587);
xor U20776 (N_20776,N_20531,N_20526);
xnor U20777 (N_20777,N_20587,N_20595);
nand U20778 (N_20778,N_20404,N_20597);
nor U20779 (N_20779,N_20429,N_20418);
nor U20780 (N_20780,N_20561,N_20519);
or U20781 (N_20781,N_20489,N_20440);
or U20782 (N_20782,N_20466,N_20415);
and U20783 (N_20783,N_20592,N_20577);
or U20784 (N_20784,N_20559,N_20530);
and U20785 (N_20785,N_20552,N_20490);
nand U20786 (N_20786,N_20470,N_20440);
nor U20787 (N_20787,N_20520,N_20544);
nor U20788 (N_20788,N_20405,N_20552);
xor U20789 (N_20789,N_20435,N_20462);
nor U20790 (N_20790,N_20558,N_20489);
xor U20791 (N_20791,N_20526,N_20574);
and U20792 (N_20792,N_20590,N_20572);
and U20793 (N_20793,N_20418,N_20499);
and U20794 (N_20794,N_20412,N_20442);
or U20795 (N_20795,N_20476,N_20427);
and U20796 (N_20796,N_20490,N_20483);
or U20797 (N_20797,N_20563,N_20518);
or U20798 (N_20798,N_20507,N_20597);
nor U20799 (N_20799,N_20577,N_20486);
or U20800 (N_20800,N_20644,N_20658);
nor U20801 (N_20801,N_20655,N_20793);
nand U20802 (N_20802,N_20746,N_20770);
or U20803 (N_20803,N_20774,N_20630);
or U20804 (N_20804,N_20738,N_20651);
and U20805 (N_20805,N_20724,N_20685);
and U20806 (N_20806,N_20610,N_20768);
nor U20807 (N_20807,N_20723,N_20784);
or U20808 (N_20808,N_20600,N_20669);
xnor U20809 (N_20809,N_20755,N_20684);
xnor U20810 (N_20810,N_20683,N_20725);
xnor U20811 (N_20811,N_20795,N_20673);
and U20812 (N_20812,N_20675,N_20615);
nor U20813 (N_20813,N_20639,N_20711);
xor U20814 (N_20814,N_20659,N_20796);
nor U20815 (N_20815,N_20717,N_20649);
or U20816 (N_20816,N_20732,N_20601);
nand U20817 (N_20817,N_20751,N_20665);
nand U20818 (N_20818,N_20642,N_20771);
and U20819 (N_20819,N_20616,N_20676);
and U20820 (N_20820,N_20663,N_20643);
nor U20821 (N_20821,N_20691,N_20757);
nor U20822 (N_20822,N_20668,N_20650);
nor U20823 (N_20823,N_20689,N_20662);
nor U20824 (N_20824,N_20710,N_20750);
nand U20825 (N_20825,N_20704,N_20635);
and U20826 (N_20826,N_20677,N_20678);
and U20827 (N_20827,N_20604,N_20721);
or U20828 (N_20828,N_20703,N_20797);
nor U20829 (N_20829,N_20603,N_20674);
and U20830 (N_20830,N_20682,N_20666);
xnor U20831 (N_20831,N_20608,N_20758);
xnor U20832 (N_20832,N_20798,N_20799);
nor U20833 (N_20833,N_20740,N_20762);
and U20834 (N_20834,N_20748,N_20617);
or U20835 (N_20835,N_20744,N_20606);
and U20836 (N_20836,N_20694,N_20705);
nor U20837 (N_20837,N_20772,N_20625);
or U20838 (N_20838,N_20759,N_20773);
nand U20839 (N_20839,N_20714,N_20712);
nand U20840 (N_20840,N_20775,N_20715);
nor U20841 (N_20841,N_20672,N_20618);
nand U20842 (N_20842,N_20646,N_20629);
and U20843 (N_20843,N_20726,N_20602);
nand U20844 (N_20844,N_20638,N_20729);
xnor U20845 (N_20845,N_20735,N_20698);
or U20846 (N_20846,N_20731,N_20754);
nor U20847 (N_20847,N_20756,N_20791);
xnor U20848 (N_20848,N_20713,N_20769);
or U20849 (N_20849,N_20624,N_20728);
nand U20850 (N_20850,N_20765,N_20645);
nor U20851 (N_20851,N_20782,N_20776);
nand U20852 (N_20852,N_20745,N_20742);
nand U20853 (N_20853,N_20741,N_20671);
or U20854 (N_20854,N_20778,N_20620);
xor U20855 (N_20855,N_20609,N_20623);
or U20856 (N_20856,N_20730,N_20767);
xor U20857 (N_20857,N_20652,N_20743);
xnor U20858 (N_20858,N_20794,N_20785);
nand U20859 (N_20859,N_20780,N_20718);
nand U20860 (N_20860,N_20637,N_20697);
nor U20861 (N_20861,N_20640,N_20627);
nand U20862 (N_20862,N_20747,N_20708);
and U20863 (N_20863,N_20612,N_20693);
xor U20864 (N_20864,N_20701,N_20690);
and U20865 (N_20865,N_20699,N_20733);
nor U20866 (N_20866,N_20790,N_20786);
and U20867 (N_20867,N_20692,N_20722);
nor U20868 (N_20868,N_20760,N_20619);
xor U20869 (N_20869,N_20761,N_20680);
and U20870 (N_20870,N_20613,N_20660);
and U20871 (N_20871,N_20653,N_20661);
nor U20872 (N_20872,N_20688,N_20766);
and U20873 (N_20873,N_20706,N_20641);
xor U20874 (N_20874,N_20752,N_20779);
nand U20875 (N_20875,N_20719,N_20686);
or U20876 (N_20876,N_20687,N_20777);
and U20877 (N_20877,N_20707,N_20628);
nand U20878 (N_20878,N_20654,N_20605);
or U20879 (N_20879,N_20621,N_20626);
nor U20880 (N_20880,N_20667,N_20737);
nand U20881 (N_20881,N_20695,N_20788);
and U20882 (N_20882,N_20679,N_20631);
or U20883 (N_20883,N_20736,N_20781);
nor U20884 (N_20884,N_20696,N_20792);
or U20885 (N_20885,N_20787,N_20636);
and U20886 (N_20886,N_20700,N_20734);
or U20887 (N_20887,N_20789,N_20763);
and U20888 (N_20888,N_20633,N_20753);
nand U20889 (N_20889,N_20783,N_20764);
xor U20890 (N_20890,N_20670,N_20656);
and U20891 (N_20891,N_20607,N_20727);
xor U20892 (N_20892,N_20739,N_20614);
and U20893 (N_20893,N_20716,N_20622);
nor U20894 (N_20894,N_20702,N_20657);
nand U20895 (N_20895,N_20634,N_20749);
or U20896 (N_20896,N_20709,N_20632);
nand U20897 (N_20897,N_20611,N_20720);
and U20898 (N_20898,N_20664,N_20648);
or U20899 (N_20899,N_20647,N_20681);
or U20900 (N_20900,N_20622,N_20757);
nor U20901 (N_20901,N_20790,N_20712);
or U20902 (N_20902,N_20760,N_20645);
xor U20903 (N_20903,N_20779,N_20731);
nand U20904 (N_20904,N_20662,N_20674);
or U20905 (N_20905,N_20707,N_20718);
nor U20906 (N_20906,N_20678,N_20705);
or U20907 (N_20907,N_20775,N_20712);
and U20908 (N_20908,N_20718,N_20675);
nor U20909 (N_20909,N_20735,N_20733);
or U20910 (N_20910,N_20794,N_20655);
xnor U20911 (N_20911,N_20644,N_20634);
xor U20912 (N_20912,N_20687,N_20749);
or U20913 (N_20913,N_20722,N_20723);
nor U20914 (N_20914,N_20730,N_20755);
nand U20915 (N_20915,N_20730,N_20658);
nor U20916 (N_20916,N_20638,N_20615);
xnor U20917 (N_20917,N_20715,N_20710);
nor U20918 (N_20918,N_20732,N_20782);
and U20919 (N_20919,N_20765,N_20653);
or U20920 (N_20920,N_20730,N_20776);
and U20921 (N_20921,N_20603,N_20782);
or U20922 (N_20922,N_20627,N_20610);
xnor U20923 (N_20923,N_20696,N_20786);
nand U20924 (N_20924,N_20656,N_20614);
or U20925 (N_20925,N_20699,N_20670);
or U20926 (N_20926,N_20621,N_20603);
and U20927 (N_20927,N_20799,N_20656);
or U20928 (N_20928,N_20636,N_20688);
and U20929 (N_20929,N_20764,N_20703);
xnor U20930 (N_20930,N_20626,N_20770);
nor U20931 (N_20931,N_20632,N_20611);
and U20932 (N_20932,N_20764,N_20752);
or U20933 (N_20933,N_20682,N_20628);
nand U20934 (N_20934,N_20770,N_20666);
nand U20935 (N_20935,N_20782,N_20792);
nor U20936 (N_20936,N_20684,N_20630);
or U20937 (N_20937,N_20698,N_20717);
nand U20938 (N_20938,N_20602,N_20675);
xnor U20939 (N_20939,N_20639,N_20634);
or U20940 (N_20940,N_20675,N_20746);
nor U20941 (N_20941,N_20756,N_20708);
and U20942 (N_20942,N_20625,N_20777);
and U20943 (N_20943,N_20750,N_20689);
and U20944 (N_20944,N_20647,N_20704);
xnor U20945 (N_20945,N_20639,N_20778);
xor U20946 (N_20946,N_20631,N_20640);
nand U20947 (N_20947,N_20617,N_20679);
or U20948 (N_20948,N_20640,N_20715);
and U20949 (N_20949,N_20666,N_20719);
and U20950 (N_20950,N_20606,N_20736);
or U20951 (N_20951,N_20743,N_20671);
nand U20952 (N_20952,N_20708,N_20697);
nor U20953 (N_20953,N_20654,N_20717);
or U20954 (N_20954,N_20694,N_20792);
or U20955 (N_20955,N_20636,N_20723);
xor U20956 (N_20956,N_20640,N_20750);
nand U20957 (N_20957,N_20705,N_20790);
nand U20958 (N_20958,N_20733,N_20737);
or U20959 (N_20959,N_20796,N_20705);
xnor U20960 (N_20960,N_20799,N_20627);
nand U20961 (N_20961,N_20625,N_20694);
xnor U20962 (N_20962,N_20658,N_20789);
nor U20963 (N_20963,N_20604,N_20636);
xor U20964 (N_20964,N_20712,N_20797);
and U20965 (N_20965,N_20630,N_20611);
or U20966 (N_20966,N_20609,N_20730);
xnor U20967 (N_20967,N_20700,N_20675);
or U20968 (N_20968,N_20681,N_20699);
xor U20969 (N_20969,N_20771,N_20732);
xor U20970 (N_20970,N_20620,N_20685);
nand U20971 (N_20971,N_20654,N_20691);
xor U20972 (N_20972,N_20647,N_20650);
nand U20973 (N_20973,N_20764,N_20777);
and U20974 (N_20974,N_20789,N_20710);
xor U20975 (N_20975,N_20737,N_20699);
or U20976 (N_20976,N_20620,N_20756);
nor U20977 (N_20977,N_20615,N_20616);
and U20978 (N_20978,N_20708,N_20623);
or U20979 (N_20979,N_20792,N_20640);
and U20980 (N_20980,N_20642,N_20649);
nand U20981 (N_20981,N_20689,N_20664);
nand U20982 (N_20982,N_20678,N_20760);
nand U20983 (N_20983,N_20762,N_20654);
and U20984 (N_20984,N_20699,N_20766);
nor U20985 (N_20985,N_20720,N_20724);
or U20986 (N_20986,N_20693,N_20771);
xnor U20987 (N_20987,N_20722,N_20765);
or U20988 (N_20988,N_20737,N_20721);
nor U20989 (N_20989,N_20734,N_20733);
xnor U20990 (N_20990,N_20630,N_20783);
nor U20991 (N_20991,N_20616,N_20653);
nor U20992 (N_20992,N_20744,N_20632);
or U20993 (N_20993,N_20712,N_20758);
and U20994 (N_20994,N_20639,N_20720);
or U20995 (N_20995,N_20792,N_20740);
nand U20996 (N_20996,N_20790,N_20640);
nor U20997 (N_20997,N_20636,N_20788);
nand U20998 (N_20998,N_20783,N_20795);
nand U20999 (N_20999,N_20682,N_20707);
xnor U21000 (N_21000,N_20809,N_20987);
and U21001 (N_21001,N_20918,N_20922);
nor U21002 (N_21002,N_20976,N_20823);
nor U21003 (N_21003,N_20863,N_20831);
or U21004 (N_21004,N_20912,N_20819);
nor U21005 (N_21005,N_20920,N_20965);
or U21006 (N_21006,N_20854,N_20967);
and U21007 (N_21007,N_20807,N_20905);
and U21008 (N_21008,N_20964,N_20891);
nand U21009 (N_21009,N_20958,N_20968);
and U21010 (N_21010,N_20861,N_20804);
or U21011 (N_21011,N_20882,N_20981);
and U21012 (N_21012,N_20837,N_20896);
xor U21013 (N_21013,N_20811,N_20887);
nand U21014 (N_21014,N_20917,N_20915);
nand U21015 (N_21015,N_20963,N_20827);
nand U21016 (N_21016,N_20980,N_20865);
nand U21017 (N_21017,N_20991,N_20890);
xnor U21018 (N_21018,N_20849,N_20936);
nand U21019 (N_21019,N_20808,N_20805);
xor U21020 (N_21020,N_20952,N_20934);
nand U21021 (N_21021,N_20972,N_20971);
nor U21022 (N_21022,N_20862,N_20950);
nand U21023 (N_21023,N_20913,N_20892);
nor U21024 (N_21024,N_20904,N_20875);
and U21025 (N_21025,N_20982,N_20914);
and U21026 (N_21026,N_20803,N_20951);
xor U21027 (N_21027,N_20969,N_20801);
nand U21028 (N_21028,N_20903,N_20906);
nor U21029 (N_21029,N_20844,N_20990);
nand U21030 (N_21030,N_20864,N_20929);
xnor U21031 (N_21031,N_20909,N_20928);
nor U21032 (N_21032,N_20894,N_20910);
nor U21033 (N_21033,N_20886,N_20860);
and U21034 (N_21034,N_20870,N_20851);
and U21035 (N_21035,N_20871,N_20821);
and U21036 (N_21036,N_20866,N_20979);
nor U21037 (N_21037,N_20828,N_20856);
nand U21038 (N_21038,N_20802,N_20924);
or U21039 (N_21039,N_20883,N_20825);
and U21040 (N_21040,N_20984,N_20927);
and U21041 (N_21041,N_20822,N_20841);
nand U21042 (N_21042,N_20975,N_20817);
nand U21043 (N_21043,N_20930,N_20932);
nor U21044 (N_21044,N_20824,N_20816);
and U21045 (N_21045,N_20940,N_20810);
and U21046 (N_21046,N_20868,N_20954);
nor U21047 (N_21047,N_20955,N_20937);
and U21048 (N_21048,N_20995,N_20983);
or U21049 (N_21049,N_20842,N_20998);
xnor U21050 (N_21050,N_20847,N_20876);
xnor U21051 (N_21051,N_20889,N_20843);
xor U21052 (N_21052,N_20884,N_20839);
and U21053 (N_21053,N_20901,N_20908);
nand U21054 (N_21054,N_20859,N_20872);
xor U21055 (N_21055,N_20953,N_20939);
nand U21056 (N_21056,N_20878,N_20978);
xnor U21057 (N_21057,N_20948,N_20966);
nand U21058 (N_21058,N_20997,N_20925);
xor U21059 (N_21059,N_20855,N_20941);
or U21060 (N_21060,N_20919,N_20833);
and U21061 (N_21061,N_20974,N_20916);
nand U21062 (N_21062,N_20994,N_20880);
and U21063 (N_21063,N_20931,N_20897);
nor U21064 (N_21064,N_20869,N_20946);
nand U21065 (N_21065,N_20900,N_20806);
nor U21066 (N_21066,N_20988,N_20840);
nand U21067 (N_21067,N_20942,N_20800);
and U21068 (N_21068,N_20973,N_20834);
and U21069 (N_21069,N_20830,N_20874);
and U21070 (N_21070,N_20813,N_20999);
or U21071 (N_21071,N_20838,N_20898);
xor U21072 (N_21072,N_20961,N_20899);
and U21073 (N_21073,N_20858,N_20885);
nand U21074 (N_21074,N_20846,N_20970);
or U21075 (N_21075,N_20826,N_20949);
nand U21076 (N_21076,N_20850,N_20815);
and U21077 (N_21077,N_20877,N_20992);
or U21078 (N_21078,N_20832,N_20814);
or U21079 (N_21079,N_20923,N_20911);
or U21080 (N_21080,N_20845,N_20935);
and U21081 (N_21081,N_20836,N_20956);
nor U21082 (N_21082,N_20895,N_20902);
xor U21083 (N_21083,N_20957,N_20959);
nor U21084 (N_21084,N_20921,N_20820);
or U21085 (N_21085,N_20944,N_20907);
xor U21086 (N_21086,N_20960,N_20835);
xor U21087 (N_21087,N_20933,N_20945);
nor U21088 (N_21088,N_20947,N_20853);
and U21089 (N_21089,N_20881,N_20812);
xor U21090 (N_21090,N_20857,N_20996);
nand U21091 (N_21091,N_20985,N_20926);
nor U21092 (N_21092,N_20962,N_20989);
xor U21093 (N_21093,N_20873,N_20867);
and U21094 (N_21094,N_20818,N_20852);
xnor U21095 (N_21095,N_20848,N_20888);
or U21096 (N_21096,N_20943,N_20986);
or U21097 (N_21097,N_20879,N_20893);
nor U21098 (N_21098,N_20938,N_20993);
xor U21099 (N_21099,N_20829,N_20977);
nand U21100 (N_21100,N_20877,N_20840);
xor U21101 (N_21101,N_20909,N_20829);
nor U21102 (N_21102,N_20805,N_20879);
xor U21103 (N_21103,N_20869,N_20972);
and U21104 (N_21104,N_20881,N_20953);
or U21105 (N_21105,N_20928,N_20848);
and U21106 (N_21106,N_20903,N_20932);
and U21107 (N_21107,N_20943,N_20963);
nor U21108 (N_21108,N_20913,N_20884);
or U21109 (N_21109,N_20840,N_20916);
nor U21110 (N_21110,N_20940,N_20895);
and U21111 (N_21111,N_20832,N_20846);
or U21112 (N_21112,N_20833,N_20963);
and U21113 (N_21113,N_20844,N_20943);
or U21114 (N_21114,N_20803,N_20944);
or U21115 (N_21115,N_20908,N_20872);
or U21116 (N_21116,N_20844,N_20832);
or U21117 (N_21117,N_20800,N_20821);
nand U21118 (N_21118,N_20916,N_20800);
nor U21119 (N_21119,N_20894,N_20912);
nor U21120 (N_21120,N_20811,N_20869);
and U21121 (N_21121,N_20947,N_20849);
xnor U21122 (N_21122,N_20876,N_20820);
xor U21123 (N_21123,N_20935,N_20852);
nand U21124 (N_21124,N_20811,N_20839);
nand U21125 (N_21125,N_20957,N_20826);
or U21126 (N_21126,N_20905,N_20993);
and U21127 (N_21127,N_20993,N_20958);
and U21128 (N_21128,N_20847,N_20875);
nor U21129 (N_21129,N_20806,N_20884);
nand U21130 (N_21130,N_20986,N_20907);
nand U21131 (N_21131,N_20955,N_20813);
nand U21132 (N_21132,N_20934,N_20924);
nor U21133 (N_21133,N_20900,N_20844);
xor U21134 (N_21134,N_20999,N_20800);
nand U21135 (N_21135,N_20829,N_20862);
or U21136 (N_21136,N_20924,N_20842);
nand U21137 (N_21137,N_20803,N_20962);
and U21138 (N_21138,N_20923,N_20892);
nor U21139 (N_21139,N_20964,N_20925);
nand U21140 (N_21140,N_20933,N_20900);
or U21141 (N_21141,N_20916,N_20848);
nand U21142 (N_21142,N_20861,N_20919);
or U21143 (N_21143,N_20804,N_20997);
and U21144 (N_21144,N_20914,N_20907);
nand U21145 (N_21145,N_20944,N_20988);
xor U21146 (N_21146,N_20913,N_20831);
nand U21147 (N_21147,N_20817,N_20935);
nand U21148 (N_21148,N_20935,N_20925);
nor U21149 (N_21149,N_20930,N_20978);
xnor U21150 (N_21150,N_20874,N_20847);
or U21151 (N_21151,N_20998,N_20982);
and U21152 (N_21152,N_20959,N_20935);
nor U21153 (N_21153,N_20848,N_20941);
nand U21154 (N_21154,N_20810,N_20837);
nand U21155 (N_21155,N_20853,N_20891);
or U21156 (N_21156,N_20810,N_20938);
and U21157 (N_21157,N_20949,N_20951);
xnor U21158 (N_21158,N_20807,N_20982);
xnor U21159 (N_21159,N_20827,N_20837);
or U21160 (N_21160,N_20876,N_20802);
or U21161 (N_21161,N_20814,N_20856);
and U21162 (N_21162,N_20814,N_20899);
and U21163 (N_21163,N_20990,N_20850);
xor U21164 (N_21164,N_20897,N_20936);
or U21165 (N_21165,N_20827,N_20856);
nand U21166 (N_21166,N_20927,N_20898);
or U21167 (N_21167,N_20932,N_20869);
nand U21168 (N_21168,N_20885,N_20896);
and U21169 (N_21169,N_20917,N_20851);
nand U21170 (N_21170,N_20872,N_20869);
nand U21171 (N_21171,N_20922,N_20894);
nand U21172 (N_21172,N_20919,N_20944);
xor U21173 (N_21173,N_20838,N_20875);
nor U21174 (N_21174,N_20995,N_20899);
nand U21175 (N_21175,N_20813,N_20899);
and U21176 (N_21176,N_20879,N_20911);
nor U21177 (N_21177,N_20831,N_20908);
or U21178 (N_21178,N_20892,N_20916);
or U21179 (N_21179,N_20911,N_20845);
and U21180 (N_21180,N_20914,N_20929);
nor U21181 (N_21181,N_20818,N_20957);
or U21182 (N_21182,N_20842,N_20893);
or U21183 (N_21183,N_20950,N_20834);
or U21184 (N_21184,N_20862,N_20803);
xor U21185 (N_21185,N_20996,N_20863);
nand U21186 (N_21186,N_20984,N_20896);
or U21187 (N_21187,N_20812,N_20983);
nor U21188 (N_21188,N_20946,N_20951);
nor U21189 (N_21189,N_20871,N_20830);
or U21190 (N_21190,N_20954,N_20981);
and U21191 (N_21191,N_20935,N_20837);
nand U21192 (N_21192,N_20969,N_20897);
nand U21193 (N_21193,N_20834,N_20989);
nor U21194 (N_21194,N_20901,N_20879);
nand U21195 (N_21195,N_20846,N_20949);
or U21196 (N_21196,N_20955,N_20883);
xor U21197 (N_21197,N_20804,N_20911);
or U21198 (N_21198,N_20845,N_20858);
nand U21199 (N_21199,N_20818,N_20955);
and U21200 (N_21200,N_21083,N_21054);
nor U21201 (N_21201,N_21002,N_21060);
nor U21202 (N_21202,N_21096,N_21148);
or U21203 (N_21203,N_21072,N_21068);
and U21204 (N_21204,N_21025,N_21061);
or U21205 (N_21205,N_21126,N_21034);
nor U21206 (N_21206,N_21197,N_21160);
nand U21207 (N_21207,N_21145,N_21161);
or U21208 (N_21208,N_21142,N_21192);
nor U21209 (N_21209,N_21110,N_21182);
nand U21210 (N_21210,N_21094,N_21144);
and U21211 (N_21211,N_21097,N_21093);
xnor U21212 (N_21212,N_21042,N_21066);
and U21213 (N_21213,N_21092,N_21167);
nor U21214 (N_21214,N_21033,N_21012);
or U21215 (N_21215,N_21069,N_21084);
and U21216 (N_21216,N_21130,N_21059);
or U21217 (N_21217,N_21117,N_21121);
nand U21218 (N_21218,N_21151,N_21147);
nand U21219 (N_21219,N_21005,N_21062);
nand U21220 (N_21220,N_21177,N_21189);
or U21221 (N_21221,N_21188,N_21043);
xor U21222 (N_21222,N_21050,N_21137);
nor U21223 (N_21223,N_21198,N_21075);
and U21224 (N_21224,N_21074,N_21052);
xnor U21225 (N_21225,N_21187,N_21150);
nor U21226 (N_21226,N_21138,N_21128);
nand U21227 (N_21227,N_21009,N_21114);
nand U21228 (N_21228,N_21171,N_21024);
and U21229 (N_21229,N_21018,N_21124);
nor U21230 (N_21230,N_21141,N_21176);
nand U21231 (N_21231,N_21175,N_21032);
and U21232 (N_21232,N_21155,N_21090);
or U21233 (N_21233,N_21038,N_21157);
or U21234 (N_21234,N_21104,N_21030);
and U21235 (N_21235,N_21179,N_21115);
nand U21236 (N_21236,N_21078,N_21131);
xnor U21237 (N_21237,N_21085,N_21191);
or U21238 (N_21238,N_21116,N_21106);
nand U21239 (N_21239,N_21140,N_21149);
nand U21240 (N_21240,N_21112,N_21058);
xnor U21241 (N_21241,N_21098,N_21111);
xnor U21242 (N_21242,N_21100,N_21132);
and U21243 (N_21243,N_21017,N_21057);
xor U21244 (N_21244,N_21180,N_21186);
or U21245 (N_21245,N_21045,N_21026);
nand U21246 (N_21246,N_21135,N_21051);
or U21247 (N_21247,N_21036,N_21071);
nand U21248 (N_21248,N_21029,N_21159);
and U21249 (N_21249,N_21101,N_21185);
or U21250 (N_21250,N_21063,N_21136);
nor U21251 (N_21251,N_21056,N_21119);
or U21252 (N_21252,N_21195,N_21156);
nor U21253 (N_21253,N_21162,N_21079);
nor U21254 (N_21254,N_21196,N_21047);
and U21255 (N_21255,N_21133,N_21073);
nand U21256 (N_21256,N_21003,N_21006);
nand U21257 (N_21257,N_21163,N_21129);
or U21258 (N_21258,N_21123,N_21103);
nand U21259 (N_21259,N_21055,N_21190);
or U21260 (N_21260,N_21020,N_21080);
nand U21261 (N_21261,N_21081,N_21070);
or U21262 (N_21262,N_21076,N_21022);
xnor U21263 (N_21263,N_21122,N_21049);
nand U21264 (N_21264,N_21108,N_21077);
xnor U21265 (N_21265,N_21019,N_21164);
nor U21266 (N_21266,N_21010,N_21153);
xnor U21267 (N_21267,N_21194,N_21152);
nor U21268 (N_21268,N_21125,N_21143);
nand U21269 (N_21269,N_21014,N_21102);
nor U21270 (N_21270,N_21178,N_21016);
or U21271 (N_21271,N_21001,N_21053);
nand U21272 (N_21272,N_21013,N_21172);
nor U21273 (N_21273,N_21168,N_21086);
xor U21274 (N_21274,N_21113,N_21048);
or U21275 (N_21275,N_21146,N_21105);
nand U21276 (N_21276,N_21087,N_21134);
nor U21277 (N_21277,N_21064,N_21099);
nand U21278 (N_21278,N_21088,N_21000);
xnor U21279 (N_21279,N_21139,N_21082);
nor U21280 (N_21280,N_21165,N_21028);
nand U21281 (N_21281,N_21166,N_21023);
nor U21282 (N_21282,N_21181,N_21184);
nor U21283 (N_21283,N_21011,N_21040);
nor U21284 (N_21284,N_21193,N_21035);
xnor U21285 (N_21285,N_21169,N_21008);
nor U21286 (N_21286,N_21118,N_21065);
nand U21287 (N_21287,N_21031,N_21120);
nor U21288 (N_21288,N_21044,N_21091);
or U21289 (N_21289,N_21158,N_21067);
and U21290 (N_21290,N_21183,N_21039);
xnor U21291 (N_21291,N_21095,N_21015);
xor U21292 (N_21292,N_21199,N_21127);
or U21293 (N_21293,N_21173,N_21037);
nand U21294 (N_21294,N_21021,N_21089);
xnor U21295 (N_21295,N_21109,N_21007);
and U21296 (N_21296,N_21170,N_21027);
xnor U21297 (N_21297,N_21041,N_21107);
nand U21298 (N_21298,N_21046,N_21154);
nor U21299 (N_21299,N_21004,N_21174);
nor U21300 (N_21300,N_21181,N_21023);
xor U21301 (N_21301,N_21184,N_21090);
or U21302 (N_21302,N_21152,N_21060);
or U21303 (N_21303,N_21119,N_21121);
or U21304 (N_21304,N_21140,N_21125);
and U21305 (N_21305,N_21089,N_21166);
or U21306 (N_21306,N_21063,N_21112);
or U21307 (N_21307,N_21029,N_21017);
nor U21308 (N_21308,N_21047,N_21012);
or U21309 (N_21309,N_21178,N_21050);
nor U21310 (N_21310,N_21018,N_21177);
or U21311 (N_21311,N_21172,N_21085);
or U21312 (N_21312,N_21178,N_21120);
nor U21313 (N_21313,N_21098,N_21175);
nand U21314 (N_21314,N_21144,N_21063);
or U21315 (N_21315,N_21068,N_21048);
nor U21316 (N_21316,N_21109,N_21161);
nor U21317 (N_21317,N_21150,N_21122);
nor U21318 (N_21318,N_21197,N_21009);
nor U21319 (N_21319,N_21037,N_21017);
and U21320 (N_21320,N_21018,N_21094);
nor U21321 (N_21321,N_21050,N_21071);
or U21322 (N_21322,N_21175,N_21115);
and U21323 (N_21323,N_21075,N_21049);
and U21324 (N_21324,N_21006,N_21022);
xnor U21325 (N_21325,N_21067,N_21182);
nand U21326 (N_21326,N_21111,N_21174);
and U21327 (N_21327,N_21002,N_21036);
and U21328 (N_21328,N_21164,N_21024);
nor U21329 (N_21329,N_21028,N_21100);
or U21330 (N_21330,N_21051,N_21132);
nand U21331 (N_21331,N_21040,N_21013);
xor U21332 (N_21332,N_21101,N_21071);
or U21333 (N_21333,N_21107,N_21182);
nand U21334 (N_21334,N_21170,N_21118);
and U21335 (N_21335,N_21039,N_21100);
xnor U21336 (N_21336,N_21105,N_21118);
nand U21337 (N_21337,N_21121,N_21180);
nor U21338 (N_21338,N_21033,N_21072);
and U21339 (N_21339,N_21035,N_21066);
xor U21340 (N_21340,N_21024,N_21013);
nor U21341 (N_21341,N_21137,N_21124);
or U21342 (N_21342,N_21180,N_21034);
or U21343 (N_21343,N_21088,N_21085);
or U21344 (N_21344,N_21004,N_21162);
nor U21345 (N_21345,N_21176,N_21005);
xor U21346 (N_21346,N_21081,N_21169);
and U21347 (N_21347,N_21169,N_21069);
xnor U21348 (N_21348,N_21171,N_21090);
or U21349 (N_21349,N_21031,N_21081);
and U21350 (N_21350,N_21013,N_21078);
nand U21351 (N_21351,N_21176,N_21085);
nor U21352 (N_21352,N_21018,N_21048);
and U21353 (N_21353,N_21136,N_21133);
nor U21354 (N_21354,N_21039,N_21129);
nand U21355 (N_21355,N_21096,N_21137);
nand U21356 (N_21356,N_21048,N_21009);
xnor U21357 (N_21357,N_21161,N_21150);
or U21358 (N_21358,N_21125,N_21156);
nor U21359 (N_21359,N_21018,N_21102);
nand U21360 (N_21360,N_21128,N_21029);
xor U21361 (N_21361,N_21020,N_21032);
xnor U21362 (N_21362,N_21006,N_21165);
nand U21363 (N_21363,N_21143,N_21062);
and U21364 (N_21364,N_21073,N_21177);
nor U21365 (N_21365,N_21113,N_21053);
or U21366 (N_21366,N_21103,N_21021);
or U21367 (N_21367,N_21021,N_21189);
xor U21368 (N_21368,N_21146,N_21093);
nor U21369 (N_21369,N_21045,N_21189);
nor U21370 (N_21370,N_21192,N_21185);
nand U21371 (N_21371,N_21146,N_21175);
nor U21372 (N_21372,N_21074,N_21199);
nor U21373 (N_21373,N_21002,N_21105);
or U21374 (N_21374,N_21018,N_21076);
and U21375 (N_21375,N_21094,N_21067);
nor U21376 (N_21376,N_21152,N_21046);
xor U21377 (N_21377,N_21060,N_21028);
or U21378 (N_21378,N_21182,N_21099);
or U21379 (N_21379,N_21020,N_21175);
or U21380 (N_21380,N_21169,N_21082);
or U21381 (N_21381,N_21127,N_21098);
nand U21382 (N_21382,N_21190,N_21028);
xnor U21383 (N_21383,N_21176,N_21095);
xor U21384 (N_21384,N_21133,N_21166);
and U21385 (N_21385,N_21137,N_21023);
xor U21386 (N_21386,N_21059,N_21042);
xnor U21387 (N_21387,N_21113,N_21024);
or U21388 (N_21388,N_21195,N_21039);
xor U21389 (N_21389,N_21111,N_21057);
and U21390 (N_21390,N_21191,N_21115);
nand U21391 (N_21391,N_21160,N_21093);
xor U21392 (N_21392,N_21120,N_21152);
nor U21393 (N_21393,N_21063,N_21188);
nor U21394 (N_21394,N_21103,N_21141);
or U21395 (N_21395,N_21019,N_21134);
and U21396 (N_21396,N_21003,N_21036);
nor U21397 (N_21397,N_21156,N_21175);
and U21398 (N_21398,N_21170,N_21072);
and U21399 (N_21399,N_21113,N_21094);
or U21400 (N_21400,N_21269,N_21214);
xnor U21401 (N_21401,N_21202,N_21237);
nand U21402 (N_21402,N_21326,N_21345);
nor U21403 (N_21403,N_21266,N_21350);
and U21404 (N_21404,N_21298,N_21381);
nand U21405 (N_21405,N_21275,N_21323);
nor U21406 (N_21406,N_21282,N_21384);
nand U21407 (N_21407,N_21376,N_21394);
or U21408 (N_21408,N_21255,N_21335);
and U21409 (N_21409,N_21277,N_21316);
and U21410 (N_21410,N_21289,N_21311);
nand U21411 (N_21411,N_21330,N_21365);
xnor U21412 (N_21412,N_21377,N_21346);
nand U21413 (N_21413,N_21355,N_21211);
nand U21414 (N_21414,N_21262,N_21363);
nor U21415 (N_21415,N_21370,N_21294);
nand U21416 (N_21416,N_21299,N_21386);
nand U21417 (N_21417,N_21343,N_21268);
xnor U21418 (N_21418,N_21221,N_21371);
or U21419 (N_21419,N_21264,N_21312);
and U21420 (N_21420,N_21375,N_21334);
xnor U21421 (N_21421,N_21230,N_21388);
nand U21422 (N_21422,N_21314,N_21246);
nand U21423 (N_21423,N_21295,N_21219);
nor U21424 (N_21424,N_21260,N_21297);
and U21425 (N_21425,N_21217,N_21296);
and U21426 (N_21426,N_21367,N_21396);
and U21427 (N_21427,N_21245,N_21322);
nand U21428 (N_21428,N_21391,N_21228);
nor U21429 (N_21429,N_21382,N_21291);
or U21430 (N_21430,N_21247,N_21373);
and U21431 (N_21431,N_21204,N_21398);
nor U21432 (N_21432,N_21313,N_21288);
or U21433 (N_21433,N_21324,N_21364);
nand U21434 (N_21434,N_21281,N_21252);
xnor U21435 (N_21435,N_21347,N_21331);
nor U21436 (N_21436,N_21307,N_21265);
or U21437 (N_21437,N_21248,N_21380);
and U21438 (N_21438,N_21250,N_21328);
nor U21439 (N_21439,N_21320,N_21368);
or U21440 (N_21440,N_21359,N_21318);
nor U21441 (N_21441,N_21261,N_21271);
xnor U21442 (N_21442,N_21226,N_21249);
or U21443 (N_21443,N_21293,N_21227);
xnor U21444 (N_21444,N_21222,N_21236);
xor U21445 (N_21445,N_21257,N_21310);
nand U21446 (N_21446,N_21270,N_21284);
nand U21447 (N_21447,N_21306,N_21209);
and U21448 (N_21448,N_21354,N_21292);
and U21449 (N_21449,N_21254,N_21353);
or U21450 (N_21450,N_21344,N_21378);
or U21451 (N_21451,N_21285,N_21304);
nor U21452 (N_21452,N_21361,N_21369);
or U21453 (N_21453,N_21348,N_21256);
nor U21454 (N_21454,N_21286,N_21232);
xnor U21455 (N_21455,N_21223,N_21205);
and U21456 (N_21456,N_21383,N_21327);
nor U21457 (N_21457,N_21215,N_21243);
nand U21458 (N_21458,N_21379,N_21220);
nor U21459 (N_21459,N_21374,N_21397);
and U21460 (N_21460,N_21352,N_21360);
nand U21461 (N_21461,N_21319,N_21200);
nor U21462 (N_21462,N_21238,N_21302);
xnor U21463 (N_21463,N_21267,N_21329);
and U21464 (N_21464,N_21213,N_21362);
nand U21465 (N_21465,N_21372,N_21358);
or U21466 (N_21466,N_21225,N_21216);
or U21467 (N_21467,N_21259,N_21272);
nor U21468 (N_21468,N_21392,N_21399);
and U21469 (N_21469,N_21393,N_21241);
and U21470 (N_21470,N_21212,N_21201);
xnor U21471 (N_21471,N_21303,N_21340);
or U21472 (N_21472,N_21279,N_21276);
nor U21473 (N_21473,N_21233,N_21305);
or U21474 (N_21474,N_21385,N_21253);
nor U21475 (N_21475,N_21315,N_21332);
and U21476 (N_21476,N_21309,N_21240);
nor U21477 (N_21477,N_21356,N_21321);
and U21478 (N_21478,N_21387,N_21283);
xnor U21479 (N_21479,N_21244,N_21251);
or U21480 (N_21480,N_21301,N_21287);
xnor U21481 (N_21481,N_21300,N_21258);
nand U21482 (N_21482,N_21336,N_21333);
or U21483 (N_21483,N_21337,N_21280);
nand U21484 (N_21484,N_21389,N_21308);
nand U21485 (N_21485,N_21239,N_21341);
xor U21486 (N_21486,N_21210,N_21325);
or U21487 (N_21487,N_21395,N_21339);
or U21488 (N_21488,N_21278,N_21208);
nor U21489 (N_21489,N_21224,N_21206);
or U21490 (N_21490,N_21317,N_21351);
nand U21491 (N_21491,N_21235,N_21338);
xnor U21492 (N_21492,N_21349,N_21242);
or U21493 (N_21493,N_21234,N_21231);
and U21494 (N_21494,N_21273,N_21274);
and U21495 (N_21495,N_21366,N_21263);
nand U21496 (N_21496,N_21203,N_21342);
nand U21497 (N_21497,N_21207,N_21290);
nor U21498 (N_21498,N_21390,N_21357);
or U21499 (N_21499,N_21229,N_21218);
nor U21500 (N_21500,N_21382,N_21216);
nand U21501 (N_21501,N_21269,N_21286);
xnor U21502 (N_21502,N_21247,N_21370);
and U21503 (N_21503,N_21220,N_21355);
nor U21504 (N_21504,N_21210,N_21267);
nand U21505 (N_21505,N_21313,N_21274);
and U21506 (N_21506,N_21331,N_21282);
nand U21507 (N_21507,N_21201,N_21364);
and U21508 (N_21508,N_21371,N_21278);
or U21509 (N_21509,N_21308,N_21372);
and U21510 (N_21510,N_21374,N_21381);
and U21511 (N_21511,N_21276,N_21350);
nor U21512 (N_21512,N_21371,N_21232);
and U21513 (N_21513,N_21204,N_21255);
xor U21514 (N_21514,N_21290,N_21368);
and U21515 (N_21515,N_21209,N_21225);
and U21516 (N_21516,N_21304,N_21209);
xnor U21517 (N_21517,N_21329,N_21380);
or U21518 (N_21518,N_21282,N_21206);
and U21519 (N_21519,N_21317,N_21203);
or U21520 (N_21520,N_21311,N_21376);
nor U21521 (N_21521,N_21368,N_21224);
nor U21522 (N_21522,N_21223,N_21391);
nand U21523 (N_21523,N_21371,N_21314);
or U21524 (N_21524,N_21301,N_21387);
nand U21525 (N_21525,N_21367,N_21207);
xnor U21526 (N_21526,N_21265,N_21253);
nand U21527 (N_21527,N_21244,N_21362);
or U21528 (N_21528,N_21287,N_21374);
or U21529 (N_21529,N_21241,N_21205);
and U21530 (N_21530,N_21297,N_21231);
and U21531 (N_21531,N_21355,N_21224);
and U21532 (N_21532,N_21336,N_21280);
nor U21533 (N_21533,N_21237,N_21228);
xor U21534 (N_21534,N_21203,N_21219);
xnor U21535 (N_21535,N_21360,N_21263);
and U21536 (N_21536,N_21328,N_21275);
xor U21537 (N_21537,N_21291,N_21255);
xor U21538 (N_21538,N_21349,N_21284);
nor U21539 (N_21539,N_21214,N_21301);
xor U21540 (N_21540,N_21221,N_21233);
nor U21541 (N_21541,N_21394,N_21209);
xnor U21542 (N_21542,N_21324,N_21346);
nand U21543 (N_21543,N_21240,N_21393);
or U21544 (N_21544,N_21378,N_21204);
nand U21545 (N_21545,N_21216,N_21367);
or U21546 (N_21546,N_21336,N_21235);
or U21547 (N_21547,N_21203,N_21279);
and U21548 (N_21548,N_21201,N_21259);
nor U21549 (N_21549,N_21320,N_21217);
xnor U21550 (N_21550,N_21297,N_21370);
nand U21551 (N_21551,N_21379,N_21297);
and U21552 (N_21552,N_21224,N_21295);
and U21553 (N_21553,N_21239,N_21303);
nand U21554 (N_21554,N_21322,N_21253);
xor U21555 (N_21555,N_21369,N_21232);
and U21556 (N_21556,N_21268,N_21345);
and U21557 (N_21557,N_21202,N_21382);
nand U21558 (N_21558,N_21354,N_21353);
nand U21559 (N_21559,N_21282,N_21280);
or U21560 (N_21560,N_21353,N_21277);
nand U21561 (N_21561,N_21323,N_21288);
and U21562 (N_21562,N_21352,N_21256);
xnor U21563 (N_21563,N_21237,N_21391);
and U21564 (N_21564,N_21302,N_21203);
and U21565 (N_21565,N_21293,N_21259);
nand U21566 (N_21566,N_21304,N_21309);
and U21567 (N_21567,N_21215,N_21257);
or U21568 (N_21568,N_21384,N_21328);
xor U21569 (N_21569,N_21364,N_21260);
nor U21570 (N_21570,N_21298,N_21220);
and U21571 (N_21571,N_21215,N_21306);
or U21572 (N_21572,N_21217,N_21299);
xor U21573 (N_21573,N_21251,N_21242);
xor U21574 (N_21574,N_21228,N_21223);
nor U21575 (N_21575,N_21397,N_21293);
nor U21576 (N_21576,N_21256,N_21394);
or U21577 (N_21577,N_21284,N_21377);
and U21578 (N_21578,N_21226,N_21251);
nand U21579 (N_21579,N_21236,N_21207);
or U21580 (N_21580,N_21374,N_21232);
and U21581 (N_21581,N_21323,N_21261);
or U21582 (N_21582,N_21393,N_21314);
nor U21583 (N_21583,N_21329,N_21294);
xor U21584 (N_21584,N_21360,N_21212);
or U21585 (N_21585,N_21370,N_21378);
xnor U21586 (N_21586,N_21245,N_21204);
nor U21587 (N_21587,N_21269,N_21224);
xor U21588 (N_21588,N_21389,N_21238);
or U21589 (N_21589,N_21294,N_21292);
nor U21590 (N_21590,N_21250,N_21246);
nor U21591 (N_21591,N_21293,N_21384);
or U21592 (N_21592,N_21291,N_21281);
nand U21593 (N_21593,N_21347,N_21250);
or U21594 (N_21594,N_21367,N_21374);
nand U21595 (N_21595,N_21351,N_21292);
nor U21596 (N_21596,N_21323,N_21332);
xor U21597 (N_21597,N_21278,N_21342);
and U21598 (N_21598,N_21313,N_21241);
or U21599 (N_21599,N_21292,N_21238);
or U21600 (N_21600,N_21558,N_21442);
xnor U21601 (N_21601,N_21572,N_21561);
nand U21602 (N_21602,N_21461,N_21438);
nand U21603 (N_21603,N_21517,N_21486);
xor U21604 (N_21604,N_21509,N_21400);
nor U21605 (N_21605,N_21418,N_21571);
and U21606 (N_21606,N_21427,N_21547);
or U21607 (N_21607,N_21406,N_21435);
nor U21608 (N_21608,N_21412,N_21451);
and U21609 (N_21609,N_21529,N_21465);
nor U21610 (N_21610,N_21496,N_21523);
xor U21611 (N_21611,N_21432,N_21456);
or U21612 (N_21612,N_21501,N_21440);
xor U21613 (N_21613,N_21505,N_21441);
nand U21614 (N_21614,N_21549,N_21524);
nand U21615 (N_21615,N_21459,N_21512);
and U21616 (N_21616,N_21522,N_21447);
nand U21617 (N_21617,N_21526,N_21428);
nor U21618 (N_21618,N_21493,N_21453);
xor U21619 (N_21619,N_21516,N_21472);
nor U21620 (N_21620,N_21504,N_21596);
nand U21621 (N_21621,N_21467,N_21463);
and U21622 (N_21622,N_21570,N_21552);
and U21623 (N_21623,N_21528,N_21539);
nor U21624 (N_21624,N_21581,N_21525);
nand U21625 (N_21625,N_21573,N_21407);
nand U21626 (N_21626,N_21550,N_21468);
nand U21627 (N_21627,N_21479,N_21536);
and U21628 (N_21628,N_21584,N_21568);
nor U21629 (N_21629,N_21578,N_21426);
xor U21630 (N_21630,N_21531,N_21591);
nor U21631 (N_21631,N_21404,N_21436);
and U21632 (N_21632,N_21458,N_21494);
xnor U21633 (N_21633,N_21508,N_21433);
nor U21634 (N_21634,N_21579,N_21597);
or U21635 (N_21635,N_21446,N_21588);
or U21636 (N_21636,N_21490,N_21474);
or U21637 (N_21637,N_21445,N_21476);
xor U21638 (N_21638,N_21566,N_21594);
and U21639 (N_21639,N_21518,N_21425);
or U21640 (N_21640,N_21534,N_21492);
xor U21641 (N_21641,N_21520,N_21478);
xor U21642 (N_21642,N_21545,N_21537);
or U21643 (N_21643,N_21500,N_21498);
nor U21644 (N_21644,N_21460,N_21555);
and U21645 (N_21645,N_21402,N_21541);
nand U21646 (N_21646,N_21421,N_21533);
and U21647 (N_21647,N_21429,N_21564);
nor U21648 (N_21648,N_21491,N_21530);
xor U21649 (N_21649,N_21489,N_21416);
and U21650 (N_21650,N_21585,N_21544);
or U21651 (N_21651,N_21538,N_21405);
nor U21652 (N_21652,N_21471,N_21444);
and U21653 (N_21653,N_21583,N_21473);
nand U21654 (N_21654,N_21466,N_21419);
nor U21655 (N_21655,N_21510,N_21414);
nor U21656 (N_21656,N_21546,N_21592);
nor U21657 (N_21657,N_21515,N_21417);
nand U21658 (N_21658,N_21502,N_21401);
xor U21659 (N_21659,N_21477,N_21475);
or U21660 (N_21660,N_21587,N_21514);
nor U21661 (N_21661,N_21411,N_21422);
and U21662 (N_21662,N_21434,N_21487);
xor U21663 (N_21663,N_21582,N_21495);
nor U21664 (N_21664,N_21548,N_21497);
nand U21665 (N_21665,N_21469,N_21565);
nand U21666 (N_21666,N_21410,N_21452);
nor U21667 (N_21667,N_21511,N_21482);
xnor U21668 (N_21668,N_21424,N_21507);
nor U21669 (N_21669,N_21521,N_21430);
nand U21670 (N_21670,N_21562,N_21576);
or U21671 (N_21671,N_21535,N_21559);
nor U21672 (N_21672,N_21553,N_21543);
xor U21673 (N_21673,N_21551,N_21563);
or U21674 (N_21674,N_21437,N_21464);
and U21675 (N_21675,N_21590,N_21577);
nand U21676 (N_21676,N_21403,N_21560);
nand U21677 (N_21677,N_21575,N_21540);
nor U21678 (N_21678,N_21443,N_21409);
nor U21679 (N_21679,N_21503,N_21449);
or U21680 (N_21680,N_21470,N_21462);
and U21681 (N_21681,N_21485,N_21448);
or U21682 (N_21682,N_21413,N_21574);
or U21683 (N_21683,N_21589,N_21519);
or U21684 (N_21684,N_21513,N_21408);
nand U21685 (N_21685,N_21484,N_21557);
or U21686 (N_21686,N_21488,N_21542);
xnor U21687 (N_21687,N_21454,N_21567);
and U21688 (N_21688,N_21598,N_21455);
xnor U21689 (N_21689,N_21439,N_21480);
nand U21690 (N_21690,N_21423,N_21481);
or U21691 (N_21691,N_21415,N_21580);
and U21692 (N_21692,N_21527,N_21420);
or U21693 (N_21693,N_21595,N_21431);
or U21694 (N_21694,N_21457,N_21450);
nand U21695 (N_21695,N_21556,N_21532);
xnor U21696 (N_21696,N_21554,N_21593);
xor U21697 (N_21697,N_21586,N_21506);
nor U21698 (N_21698,N_21483,N_21569);
nor U21699 (N_21699,N_21499,N_21599);
nand U21700 (N_21700,N_21487,N_21414);
and U21701 (N_21701,N_21556,N_21463);
nor U21702 (N_21702,N_21453,N_21562);
nor U21703 (N_21703,N_21468,N_21440);
and U21704 (N_21704,N_21505,N_21407);
nor U21705 (N_21705,N_21500,N_21574);
nor U21706 (N_21706,N_21588,N_21585);
xnor U21707 (N_21707,N_21495,N_21571);
and U21708 (N_21708,N_21423,N_21555);
nor U21709 (N_21709,N_21469,N_21594);
nand U21710 (N_21710,N_21563,N_21571);
xnor U21711 (N_21711,N_21524,N_21578);
xor U21712 (N_21712,N_21488,N_21499);
xnor U21713 (N_21713,N_21597,N_21420);
nand U21714 (N_21714,N_21554,N_21482);
nor U21715 (N_21715,N_21573,N_21510);
xor U21716 (N_21716,N_21577,N_21476);
xnor U21717 (N_21717,N_21426,N_21509);
nor U21718 (N_21718,N_21551,N_21482);
nor U21719 (N_21719,N_21499,N_21495);
xnor U21720 (N_21720,N_21460,N_21485);
or U21721 (N_21721,N_21542,N_21536);
xor U21722 (N_21722,N_21501,N_21524);
nand U21723 (N_21723,N_21569,N_21440);
nand U21724 (N_21724,N_21518,N_21420);
and U21725 (N_21725,N_21553,N_21476);
or U21726 (N_21726,N_21402,N_21584);
nor U21727 (N_21727,N_21548,N_21585);
nor U21728 (N_21728,N_21589,N_21427);
and U21729 (N_21729,N_21455,N_21452);
and U21730 (N_21730,N_21572,N_21519);
xnor U21731 (N_21731,N_21407,N_21521);
nor U21732 (N_21732,N_21485,N_21521);
and U21733 (N_21733,N_21492,N_21407);
nor U21734 (N_21734,N_21485,N_21429);
or U21735 (N_21735,N_21547,N_21428);
and U21736 (N_21736,N_21430,N_21542);
nor U21737 (N_21737,N_21427,N_21544);
and U21738 (N_21738,N_21582,N_21426);
or U21739 (N_21739,N_21568,N_21479);
or U21740 (N_21740,N_21587,N_21429);
or U21741 (N_21741,N_21519,N_21577);
nand U21742 (N_21742,N_21420,N_21413);
nand U21743 (N_21743,N_21415,N_21482);
nand U21744 (N_21744,N_21437,N_21424);
and U21745 (N_21745,N_21508,N_21441);
nand U21746 (N_21746,N_21401,N_21430);
nor U21747 (N_21747,N_21454,N_21403);
xnor U21748 (N_21748,N_21526,N_21543);
xnor U21749 (N_21749,N_21578,N_21582);
and U21750 (N_21750,N_21527,N_21567);
nand U21751 (N_21751,N_21485,N_21536);
nand U21752 (N_21752,N_21549,N_21595);
nor U21753 (N_21753,N_21543,N_21552);
nor U21754 (N_21754,N_21403,N_21462);
nand U21755 (N_21755,N_21549,N_21571);
nand U21756 (N_21756,N_21418,N_21402);
nand U21757 (N_21757,N_21529,N_21478);
xnor U21758 (N_21758,N_21542,N_21438);
xnor U21759 (N_21759,N_21431,N_21578);
xnor U21760 (N_21760,N_21530,N_21506);
and U21761 (N_21761,N_21428,N_21568);
and U21762 (N_21762,N_21448,N_21409);
or U21763 (N_21763,N_21521,N_21580);
and U21764 (N_21764,N_21453,N_21555);
or U21765 (N_21765,N_21406,N_21541);
nor U21766 (N_21766,N_21458,N_21484);
nand U21767 (N_21767,N_21446,N_21596);
xnor U21768 (N_21768,N_21420,N_21501);
nor U21769 (N_21769,N_21501,N_21565);
xnor U21770 (N_21770,N_21556,N_21424);
xor U21771 (N_21771,N_21582,N_21513);
or U21772 (N_21772,N_21426,N_21547);
xor U21773 (N_21773,N_21425,N_21521);
nor U21774 (N_21774,N_21471,N_21418);
or U21775 (N_21775,N_21501,N_21550);
and U21776 (N_21776,N_21408,N_21556);
nor U21777 (N_21777,N_21422,N_21447);
and U21778 (N_21778,N_21425,N_21537);
and U21779 (N_21779,N_21587,N_21576);
or U21780 (N_21780,N_21517,N_21530);
nand U21781 (N_21781,N_21592,N_21574);
and U21782 (N_21782,N_21407,N_21483);
xor U21783 (N_21783,N_21445,N_21405);
or U21784 (N_21784,N_21483,N_21476);
nor U21785 (N_21785,N_21455,N_21448);
or U21786 (N_21786,N_21417,N_21513);
and U21787 (N_21787,N_21592,N_21438);
nor U21788 (N_21788,N_21558,N_21456);
nand U21789 (N_21789,N_21569,N_21583);
nor U21790 (N_21790,N_21510,N_21565);
nand U21791 (N_21791,N_21569,N_21467);
and U21792 (N_21792,N_21551,N_21525);
or U21793 (N_21793,N_21543,N_21423);
xnor U21794 (N_21794,N_21541,N_21511);
xnor U21795 (N_21795,N_21587,N_21533);
nor U21796 (N_21796,N_21449,N_21522);
nor U21797 (N_21797,N_21477,N_21553);
nand U21798 (N_21798,N_21416,N_21503);
nand U21799 (N_21799,N_21474,N_21405);
xnor U21800 (N_21800,N_21601,N_21735);
or U21801 (N_21801,N_21622,N_21676);
and U21802 (N_21802,N_21606,N_21715);
nand U21803 (N_21803,N_21757,N_21618);
nand U21804 (N_21804,N_21798,N_21600);
nor U21805 (N_21805,N_21660,N_21634);
xor U21806 (N_21806,N_21771,N_21609);
nand U21807 (N_21807,N_21701,N_21780);
nand U21808 (N_21808,N_21756,N_21604);
nor U21809 (N_21809,N_21643,N_21773);
nand U21810 (N_21810,N_21742,N_21686);
and U21811 (N_21811,N_21629,N_21646);
or U21812 (N_21812,N_21746,N_21799);
nor U21813 (N_21813,N_21627,N_21640);
xnor U21814 (N_21814,N_21795,N_21767);
xnor U21815 (N_21815,N_21741,N_21680);
and U21816 (N_21816,N_21752,N_21671);
or U21817 (N_21817,N_21655,N_21781);
and U21818 (N_21818,N_21648,N_21726);
or U21819 (N_21819,N_21690,N_21751);
nand U21820 (N_21820,N_21638,N_21650);
xnor U21821 (N_21821,N_21739,N_21761);
nand U21822 (N_21822,N_21717,N_21685);
nand U21823 (N_21823,N_21796,N_21617);
nand U21824 (N_21824,N_21718,N_21793);
or U21825 (N_21825,N_21612,N_21694);
and U21826 (N_21826,N_21631,N_21794);
xor U21827 (N_21827,N_21788,N_21791);
and U21828 (N_21828,N_21697,N_21696);
nand U21829 (N_21829,N_21673,N_21709);
nand U21830 (N_21830,N_21623,N_21614);
nor U21831 (N_21831,N_21667,N_21719);
nor U21832 (N_21832,N_21626,N_21783);
nand U21833 (N_21833,N_21691,N_21654);
and U21834 (N_21834,N_21641,N_21682);
xor U21835 (N_21835,N_21663,N_21786);
or U21836 (N_21836,N_21679,N_21698);
nand U21837 (N_21837,N_21695,N_21714);
xnor U21838 (N_21838,N_21722,N_21675);
xor U21839 (N_21839,N_21745,N_21760);
nand U21840 (N_21840,N_21615,N_21613);
and U21841 (N_21841,N_21787,N_21738);
nor U21842 (N_21842,N_21774,N_21672);
or U21843 (N_21843,N_21723,N_21743);
nor U21844 (N_21844,N_21630,N_21724);
nand U21845 (N_21845,N_21677,N_21731);
or U21846 (N_21846,N_21633,N_21705);
nand U21847 (N_21847,N_21748,N_21716);
or U21848 (N_21848,N_21602,N_21713);
xnor U21849 (N_21849,N_21610,N_21620);
nand U21850 (N_21850,N_21710,N_21693);
and U21851 (N_21851,N_21644,N_21645);
nand U21852 (N_21852,N_21737,N_21624);
xor U21853 (N_21853,N_21608,N_21632);
nor U21854 (N_21854,N_21721,N_21764);
and U21855 (N_21855,N_21747,N_21668);
nand U21856 (N_21856,N_21734,N_21605);
or U21857 (N_21857,N_21736,N_21750);
xor U21858 (N_21858,N_21711,N_21670);
nand U21859 (N_21859,N_21683,N_21636);
xor U21860 (N_21860,N_21759,N_21789);
and U21861 (N_21861,N_21728,N_21755);
nor U21862 (N_21862,N_21775,N_21687);
or U21863 (N_21863,N_21628,N_21625);
or U21864 (N_21864,N_21635,N_21706);
and U21865 (N_21865,N_21653,N_21708);
nand U21866 (N_21866,N_21702,N_21712);
xnor U21867 (N_21867,N_21753,N_21616);
or U21868 (N_21868,N_21647,N_21664);
and U21869 (N_21869,N_21784,N_21749);
or U21870 (N_21870,N_21790,N_21656);
xor U21871 (N_21871,N_21700,N_21652);
nand U21872 (N_21872,N_21666,N_21649);
nor U21873 (N_21873,N_21657,N_21669);
xnor U21874 (N_21874,N_21619,N_21665);
or U21875 (N_21875,N_21772,N_21681);
or U21876 (N_21876,N_21744,N_21707);
nor U21877 (N_21877,N_21797,N_21779);
and U21878 (N_21878,N_21642,N_21692);
and U21879 (N_21879,N_21699,N_21611);
or U21880 (N_21880,N_21729,N_21770);
nand U21881 (N_21881,N_21765,N_21792);
nor U21882 (N_21882,N_21659,N_21678);
nor U21883 (N_21883,N_21651,N_21674);
or U21884 (N_21884,N_21703,N_21658);
or U21885 (N_21885,N_21684,N_21732);
nand U21886 (N_21886,N_21740,N_21766);
xor U21887 (N_21887,N_21603,N_21758);
nand U21888 (N_21888,N_21607,N_21776);
nor U21889 (N_21889,N_21754,N_21769);
xor U21890 (N_21890,N_21768,N_21785);
and U21891 (N_21891,N_21763,N_21621);
and U21892 (N_21892,N_21733,N_21662);
or U21893 (N_21893,N_21778,N_21661);
xnor U21894 (N_21894,N_21762,N_21704);
and U21895 (N_21895,N_21637,N_21720);
nor U21896 (N_21896,N_21782,N_21730);
nand U21897 (N_21897,N_21639,N_21777);
xor U21898 (N_21898,N_21725,N_21688);
or U21899 (N_21899,N_21727,N_21689);
xor U21900 (N_21900,N_21661,N_21618);
and U21901 (N_21901,N_21697,N_21750);
xor U21902 (N_21902,N_21792,N_21750);
nand U21903 (N_21903,N_21621,N_21710);
nand U21904 (N_21904,N_21741,N_21644);
xnor U21905 (N_21905,N_21775,N_21780);
and U21906 (N_21906,N_21683,N_21630);
nor U21907 (N_21907,N_21613,N_21750);
or U21908 (N_21908,N_21601,N_21734);
xor U21909 (N_21909,N_21794,N_21705);
nor U21910 (N_21910,N_21608,N_21727);
or U21911 (N_21911,N_21670,N_21624);
or U21912 (N_21912,N_21782,N_21635);
nor U21913 (N_21913,N_21789,N_21701);
xor U21914 (N_21914,N_21726,N_21691);
xnor U21915 (N_21915,N_21788,N_21610);
nand U21916 (N_21916,N_21660,N_21690);
or U21917 (N_21917,N_21670,N_21635);
and U21918 (N_21918,N_21687,N_21754);
xor U21919 (N_21919,N_21738,N_21691);
xor U21920 (N_21920,N_21728,N_21604);
xnor U21921 (N_21921,N_21679,N_21626);
or U21922 (N_21922,N_21697,N_21732);
or U21923 (N_21923,N_21780,N_21739);
nand U21924 (N_21924,N_21638,N_21688);
xnor U21925 (N_21925,N_21700,N_21671);
xnor U21926 (N_21926,N_21687,N_21710);
or U21927 (N_21927,N_21706,N_21771);
or U21928 (N_21928,N_21673,N_21666);
xor U21929 (N_21929,N_21742,N_21636);
or U21930 (N_21930,N_21610,N_21790);
and U21931 (N_21931,N_21659,N_21774);
nor U21932 (N_21932,N_21700,N_21766);
xnor U21933 (N_21933,N_21751,N_21775);
nand U21934 (N_21934,N_21615,N_21788);
nor U21935 (N_21935,N_21693,N_21756);
or U21936 (N_21936,N_21667,N_21727);
nand U21937 (N_21937,N_21665,N_21664);
nor U21938 (N_21938,N_21630,N_21709);
xor U21939 (N_21939,N_21617,N_21738);
and U21940 (N_21940,N_21600,N_21619);
nand U21941 (N_21941,N_21606,N_21672);
and U21942 (N_21942,N_21712,N_21722);
and U21943 (N_21943,N_21606,N_21767);
and U21944 (N_21944,N_21711,N_21687);
or U21945 (N_21945,N_21786,N_21753);
or U21946 (N_21946,N_21667,N_21770);
and U21947 (N_21947,N_21665,N_21682);
nand U21948 (N_21948,N_21714,N_21697);
xor U21949 (N_21949,N_21674,N_21742);
nand U21950 (N_21950,N_21716,N_21623);
or U21951 (N_21951,N_21636,N_21605);
or U21952 (N_21952,N_21698,N_21616);
nand U21953 (N_21953,N_21658,N_21689);
xor U21954 (N_21954,N_21687,N_21717);
or U21955 (N_21955,N_21640,N_21777);
xor U21956 (N_21956,N_21704,N_21736);
nor U21957 (N_21957,N_21772,N_21655);
nand U21958 (N_21958,N_21649,N_21646);
nor U21959 (N_21959,N_21785,N_21745);
or U21960 (N_21960,N_21716,N_21713);
nand U21961 (N_21961,N_21759,N_21731);
xor U21962 (N_21962,N_21724,N_21773);
nor U21963 (N_21963,N_21627,N_21683);
or U21964 (N_21964,N_21763,N_21739);
xor U21965 (N_21965,N_21720,N_21639);
xor U21966 (N_21966,N_21663,N_21731);
or U21967 (N_21967,N_21627,N_21723);
xnor U21968 (N_21968,N_21684,N_21613);
nor U21969 (N_21969,N_21750,N_21756);
nor U21970 (N_21970,N_21705,N_21739);
and U21971 (N_21971,N_21718,N_21625);
nor U21972 (N_21972,N_21699,N_21666);
xor U21973 (N_21973,N_21610,N_21632);
nand U21974 (N_21974,N_21673,N_21629);
and U21975 (N_21975,N_21644,N_21725);
xor U21976 (N_21976,N_21719,N_21671);
xor U21977 (N_21977,N_21780,N_21639);
nand U21978 (N_21978,N_21779,N_21642);
and U21979 (N_21979,N_21733,N_21759);
nor U21980 (N_21980,N_21607,N_21762);
xor U21981 (N_21981,N_21665,N_21635);
nor U21982 (N_21982,N_21647,N_21711);
or U21983 (N_21983,N_21635,N_21755);
or U21984 (N_21984,N_21674,N_21652);
nor U21985 (N_21985,N_21775,N_21704);
nand U21986 (N_21986,N_21656,N_21761);
xnor U21987 (N_21987,N_21799,N_21709);
or U21988 (N_21988,N_21600,N_21723);
xor U21989 (N_21989,N_21701,N_21722);
nand U21990 (N_21990,N_21601,N_21714);
or U21991 (N_21991,N_21654,N_21713);
or U21992 (N_21992,N_21699,N_21745);
and U21993 (N_21993,N_21614,N_21703);
and U21994 (N_21994,N_21689,N_21786);
nor U21995 (N_21995,N_21640,N_21754);
nor U21996 (N_21996,N_21637,N_21638);
or U21997 (N_21997,N_21768,N_21762);
and U21998 (N_21998,N_21647,N_21693);
xnor U21999 (N_21999,N_21625,N_21719);
and U22000 (N_22000,N_21893,N_21825);
xor U22001 (N_22001,N_21938,N_21979);
and U22002 (N_22002,N_21864,N_21830);
xnor U22003 (N_22003,N_21919,N_21849);
and U22004 (N_22004,N_21930,N_21933);
and U22005 (N_22005,N_21977,N_21943);
nor U22006 (N_22006,N_21904,N_21875);
nor U22007 (N_22007,N_21816,N_21845);
nand U22008 (N_22008,N_21998,N_21906);
xor U22009 (N_22009,N_21807,N_21950);
or U22010 (N_22010,N_21912,N_21987);
xor U22011 (N_22011,N_21899,N_21853);
nand U22012 (N_22012,N_21868,N_21862);
nand U22013 (N_22013,N_21841,N_21993);
and U22014 (N_22014,N_21890,N_21801);
xnor U22015 (N_22015,N_21903,N_21958);
nand U22016 (N_22016,N_21964,N_21896);
nand U22017 (N_22017,N_21866,N_21983);
or U22018 (N_22018,N_21872,N_21995);
or U22019 (N_22019,N_21895,N_21985);
nand U22020 (N_22020,N_21833,N_21994);
and U22021 (N_22021,N_21902,N_21852);
and U22022 (N_22022,N_21926,N_21911);
or U22023 (N_22023,N_21855,N_21886);
or U22024 (N_22024,N_21851,N_21867);
nor U22025 (N_22025,N_21821,N_21885);
and U22026 (N_22026,N_21808,N_21806);
nand U22027 (N_22027,N_21837,N_21952);
nand U22028 (N_22028,N_21978,N_21914);
nor U22029 (N_22029,N_21870,N_21887);
nor U22030 (N_22030,N_21850,N_21939);
and U22031 (N_22031,N_21961,N_21948);
xor U22032 (N_22032,N_21999,N_21913);
or U22033 (N_22033,N_21920,N_21874);
or U22034 (N_22034,N_21947,N_21921);
or U22035 (N_22035,N_21932,N_21972);
nor U22036 (N_22036,N_21826,N_21846);
or U22037 (N_22037,N_21836,N_21829);
nand U22038 (N_22038,N_21842,N_21934);
nor U22039 (N_22039,N_21854,N_21888);
nor U22040 (N_22040,N_21857,N_21949);
xor U22041 (N_22041,N_21869,N_21892);
xor U22042 (N_22042,N_21882,N_21881);
nor U22043 (N_22043,N_21944,N_21884);
nor U22044 (N_22044,N_21856,N_21988);
nand U22045 (N_22045,N_21820,N_21937);
nand U22046 (N_22046,N_21844,N_21828);
and U22047 (N_22047,N_21861,N_21980);
nand U22048 (N_22048,N_21838,N_21936);
and U22049 (N_22049,N_21971,N_21905);
and U22050 (N_22050,N_21834,N_21992);
nand U22051 (N_22051,N_21898,N_21942);
nor U22052 (N_22052,N_21839,N_21923);
and U22053 (N_22053,N_21945,N_21946);
nand U22054 (N_22054,N_21929,N_21907);
xor U22055 (N_22055,N_21840,N_21959);
and U22056 (N_22056,N_21809,N_21873);
xnor U22057 (N_22057,N_21910,N_21917);
nor U22058 (N_22058,N_21865,N_21883);
or U22059 (N_22059,N_21966,N_21990);
and U22060 (N_22060,N_21811,N_21812);
and U22061 (N_22061,N_21957,N_21941);
or U22062 (N_22062,N_21974,N_21805);
nor U22063 (N_22063,N_21813,N_21877);
and U22064 (N_22064,N_21880,N_21817);
nand U22065 (N_22065,N_21814,N_21860);
or U22066 (N_22066,N_21963,N_21991);
and U22067 (N_22067,N_21800,N_21815);
and U22068 (N_22068,N_21975,N_21891);
nor U22069 (N_22069,N_21940,N_21847);
nand U22070 (N_22070,N_21965,N_21824);
nand U22071 (N_22071,N_21897,N_21924);
nand U22072 (N_22072,N_21968,N_21810);
and U22073 (N_22073,N_21822,N_21908);
and U22074 (N_22074,N_21960,N_21954);
xnor U22075 (N_22075,N_21915,N_21843);
nor U22076 (N_22076,N_21935,N_21819);
and U22077 (N_22077,N_21928,N_21970);
nor U22078 (N_22078,N_21989,N_21848);
and U22079 (N_22079,N_21918,N_21876);
or U22080 (N_22080,N_21802,N_21900);
nor U22081 (N_22081,N_21916,N_21889);
and U22082 (N_22082,N_21956,N_21969);
or U22083 (N_22083,N_21976,N_21901);
nand U22084 (N_22084,N_21984,N_21927);
and U22085 (N_22085,N_21871,N_21955);
nor U22086 (N_22086,N_21962,N_21804);
nor U22087 (N_22087,N_21858,N_21859);
xnor U22088 (N_22088,N_21967,N_21909);
or U22089 (N_22089,N_21831,N_21981);
nor U22090 (N_22090,N_21835,N_21951);
xnor U22091 (N_22091,N_21818,N_21879);
and U22092 (N_22092,N_21925,N_21823);
nand U22093 (N_22093,N_21973,N_21996);
nor U22094 (N_22094,N_21827,N_21931);
nand U22095 (N_22095,N_21953,N_21878);
or U22096 (N_22096,N_21982,N_21832);
or U22097 (N_22097,N_21986,N_21894);
nor U22098 (N_22098,N_21863,N_21922);
nand U22099 (N_22099,N_21997,N_21803);
or U22100 (N_22100,N_21853,N_21913);
nor U22101 (N_22101,N_21970,N_21875);
nand U22102 (N_22102,N_21837,N_21879);
nand U22103 (N_22103,N_21933,N_21915);
or U22104 (N_22104,N_21979,N_21848);
or U22105 (N_22105,N_21872,N_21930);
and U22106 (N_22106,N_21800,N_21922);
or U22107 (N_22107,N_21916,N_21912);
and U22108 (N_22108,N_21946,N_21910);
or U22109 (N_22109,N_21806,N_21869);
nor U22110 (N_22110,N_21856,N_21995);
nor U22111 (N_22111,N_21879,N_21895);
or U22112 (N_22112,N_21929,N_21930);
nand U22113 (N_22113,N_21876,N_21857);
and U22114 (N_22114,N_21996,N_21942);
or U22115 (N_22115,N_21992,N_21953);
xnor U22116 (N_22116,N_21978,N_21815);
or U22117 (N_22117,N_21860,N_21872);
and U22118 (N_22118,N_21861,N_21827);
nand U22119 (N_22119,N_21932,N_21807);
xor U22120 (N_22120,N_21834,N_21876);
nor U22121 (N_22121,N_21975,N_21994);
xnor U22122 (N_22122,N_21968,N_21938);
and U22123 (N_22123,N_21986,N_21890);
nor U22124 (N_22124,N_21986,N_21844);
nor U22125 (N_22125,N_21972,N_21975);
or U22126 (N_22126,N_21996,N_21993);
and U22127 (N_22127,N_21859,N_21857);
and U22128 (N_22128,N_21821,N_21850);
or U22129 (N_22129,N_21813,N_21816);
nand U22130 (N_22130,N_21921,N_21840);
nor U22131 (N_22131,N_21893,N_21866);
nor U22132 (N_22132,N_21898,N_21903);
xor U22133 (N_22133,N_21857,N_21823);
and U22134 (N_22134,N_21867,N_21956);
or U22135 (N_22135,N_21922,N_21852);
xnor U22136 (N_22136,N_21993,N_21951);
xor U22137 (N_22137,N_21998,N_21953);
or U22138 (N_22138,N_21859,N_21819);
and U22139 (N_22139,N_21825,N_21877);
nand U22140 (N_22140,N_21941,N_21853);
nand U22141 (N_22141,N_21855,N_21836);
and U22142 (N_22142,N_21859,N_21905);
xor U22143 (N_22143,N_21961,N_21899);
xnor U22144 (N_22144,N_21800,N_21865);
and U22145 (N_22145,N_21926,N_21886);
and U22146 (N_22146,N_21931,N_21992);
or U22147 (N_22147,N_21858,N_21967);
xnor U22148 (N_22148,N_21818,N_21877);
nand U22149 (N_22149,N_21820,N_21907);
nand U22150 (N_22150,N_21852,N_21821);
xnor U22151 (N_22151,N_21830,N_21946);
nor U22152 (N_22152,N_21862,N_21808);
and U22153 (N_22153,N_21897,N_21992);
and U22154 (N_22154,N_21801,N_21874);
xnor U22155 (N_22155,N_21854,N_21959);
nor U22156 (N_22156,N_21881,N_21826);
xnor U22157 (N_22157,N_21907,N_21993);
nand U22158 (N_22158,N_21898,N_21998);
nor U22159 (N_22159,N_21832,N_21854);
nand U22160 (N_22160,N_21867,N_21884);
nand U22161 (N_22161,N_21857,N_21936);
nand U22162 (N_22162,N_21998,N_21873);
xnor U22163 (N_22163,N_21832,N_21844);
or U22164 (N_22164,N_21854,N_21861);
xnor U22165 (N_22165,N_21968,N_21893);
or U22166 (N_22166,N_21908,N_21941);
or U22167 (N_22167,N_21833,N_21818);
nand U22168 (N_22168,N_21813,N_21978);
xor U22169 (N_22169,N_21976,N_21925);
or U22170 (N_22170,N_21897,N_21978);
and U22171 (N_22171,N_21897,N_21809);
or U22172 (N_22172,N_21960,N_21953);
or U22173 (N_22173,N_21827,N_21944);
xnor U22174 (N_22174,N_21994,N_21814);
or U22175 (N_22175,N_21819,N_21947);
and U22176 (N_22176,N_21886,N_21948);
or U22177 (N_22177,N_21813,N_21833);
and U22178 (N_22178,N_21966,N_21957);
and U22179 (N_22179,N_21920,N_21873);
nand U22180 (N_22180,N_21915,N_21905);
and U22181 (N_22181,N_21978,N_21908);
or U22182 (N_22182,N_21860,N_21955);
xor U22183 (N_22183,N_21991,N_21808);
or U22184 (N_22184,N_21996,N_21951);
nand U22185 (N_22185,N_21868,N_21829);
xnor U22186 (N_22186,N_21982,N_21837);
nor U22187 (N_22187,N_21974,N_21891);
xor U22188 (N_22188,N_21904,N_21865);
xor U22189 (N_22189,N_21917,N_21983);
or U22190 (N_22190,N_21843,N_21852);
xnor U22191 (N_22191,N_21857,N_21812);
or U22192 (N_22192,N_21902,N_21807);
nor U22193 (N_22193,N_21988,N_21916);
xnor U22194 (N_22194,N_21833,N_21958);
nor U22195 (N_22195,N_21966,N_21857);
nor U22196 (N_22196,N_21924,N_21938);
xnor U22197 (N_22197,N_21913,N_21908);
xor U22198 (N_22198,N_21887,N_21923);
nor U22199 (N_22199,N_21857,N_21848);
nand U22200 (N_22200,N_22083,N_22026);
and U22201 (N_22201,N_22098,N_22027);
xnor U22202 (N_22202,N_22131,N_22156);
and U22203 (N_22203,N_22069,N_22063);
nor U22204 (N_22204,N_22175,N_22196);
and U22205 (N_22205,N_22085,N_22088);
nand U22206 (N_22206,N_22151,N_22080);
or U22207 (N_22207,N_22001,N_22003);
or U22208 (N_22208,N_22153,N_22181);
nand U22209 (N_22209,N_22000,N_22178);
nor U22210 (N_22210,N_22115,N_22091);
or U22211 (N_22211,N_22145,N_22070);
nand U22212 (N_22212,N_22055,N_22007);
nand U22213 (N_22213,N_22140,N_22173);
nor U22214 (N_22214,N_22104,N_22167);
nor U22215 (N_22215,N_22134,N_22022);
or U22216 (N_22216,N_22004,N_22165);
xnor U22217 (N_22217,N_22176,N_22159);
nor U22218 (N_22218,N_22142,N_22092);
nor U22219 (N_22219,N_22146,N_22136);
nand U22220 (N_22220,N_22141,N_22170);
nor U22221 (N_22221,N_22038,N_22013);
or U22222 (N_22222,N_22034,N_22191);
nor U22223 (N_22223,N_22157,N_22002);
or U22224 (N_22224,N_22014,N_22152);
or U22225 (N_22225,N_22184,N_22194);
xor U22226 (N_22226,N_22109,N_22024);
or U22227 (N_22227,N_22020,N_22139);
nor U22228 (N_22228,N_22072,N_22094);
and U22229 (N_22229,N_22075,N_22037);
or U22230 (N_22230,N_22016,N_22060);
and U22231 (N_22231,N_22086,N_22025);
or U22232 (N_22232,N_22147,N_22127);
or U22233 (N_22233,N_22130,N_22084);
xor U22234 (N_22234,N_22179,N_22028);
nor U22235 (N_22235,N_22113,N_22066);
and U22236 (N_22236,N_22067,N_22076);
and U22237 (N_22237,N_22090,N_22121);
xor U22238 (N_22238,N_22133,N_22163);
nand U22239 (N_22239,N_22015,N_22044);
nand U22240 (N_22240,N_22123,N_22008);
and U22241 (N_22241,N_22089,N_22033);
xnor U22242 (N_22242,N_22190,N_22122);
nand U22243 (N_22243,N_22198,N_22050);
xnor U22244 (N_22244,N_22096,N_22172);
nand U22245 (N_22245,N_22171,N_22197);
and U22246 (N_22246,N_22029,N_22005);
nand U22247 (N_22247,N_22103,N_22192);
and U22248 (N_22248,N_22112,N_22185);
nand U22249 (N_22249,N_22035,N_22023);
nor U22250 (N_22250,N_22186,N_22100);
xnor U22251 (N_22251,N_22054,N_22078);
nor U22252 (N_22252,N_22071,N_22074);
nand U22253 (N_22253,N_22118,N_22124);
and U22254 (N_22254,N_22011,N_22052);
and U22255 (N_22255,N_22174,N_22059);
nor U22256 (N_22256,N_22051,N_22077);
and U22257 (N_22257,N_22188,N_22047);
or U22258 (N_22258,N_22177,N_22128);
nor U22259 (N_22259,N_22125,N_22079);
and U22260 (N_22260,N_22160,N_22155);
or U22261 (N_22261,N_22148,N_22036);
or U22262 (N_22262,N_22065,N_22187);
xnor U22263 (N_22263,N_22138,N_22099);
xnor U22264 (N_22264,N_22114,N_22082);
nor U22265 (N_22265,N_22199,N_22144);
xnor U22266 (N_22266,N_22043,N_22009);
and U22267 (N_22267,N_22010,N_22046);
nor U22268 (N_22268,N_22166,N_22012);
nor U22269 (N_22269,N_22117,N_22087);
xnor U22270 (N_22270,N_22097,N_22108);
xor U22271 (N_22271,N_22149,N_22183);
and U22272 (N_22272,N_22111,N_22162);
nor U22273 (N_22273,N_22068,N_22006);
xnor U22274 (N_22274,N_22093,N_22031);
and U22275 (N_22275,N_22018,N_22169);
nor U22276 (N_22276,N_22040,N_22030);
nand U22277 (N_22277,N_22064,N_22158);
or U22278 (N_22278,N_22189,N_22135);
nand U22279 (N_22279,N_22150,N_22195);
and U22280 (N_22280,N_22019,N_22039);
nor U22281 (N_22281,N_22061,N_22058);
and U22282 (N_22282,N_22129,N_22057);
nor U22283 (N_22283,N_22062,N_22107);
or U22284 (N_22284,N_22081,N_22182);
or U22285 (N_22285,N_22042,N_22073);
or U22286 (N_22286,N_22120,N_22041);
nor U22287 (N_22287,N_22017,N_22161);
xnor U22288 (N_22288,N_22116,N_22180);
nor U22289 (N_22289,N_22110,N_22154);
nor U22290 (N_22290,N_22021,N_22056);
or U22291 (N_22291,N_22137,N_22049);
nor U22292 (N_22292,N_22032,N_22164);
nor U22293 (N_22293,N_22168,N_22102);
and U22294 (N_22294,N_22132,N_22045);
nand U22295 (N_22295,N_22048,N_22101);
xnor U22296 (N_22296,N_22143,N_22105);
xor U22297 (N_22297,N_22095,N_22126);
nand U22298 (N_22298,N_22053,N_22193);
nor U22299 (N_22299,N_22106,N_22119);
xnor U22300 (N_22300,N_22154,N_22141);
xnor U22301 (N_22301,N_22016,N_22062);
nand U22302 (N_22302,N_22027,N_22003);
or U22303 (N_22303,N_22135,N_22076);
or U22304 (N_22304,N_22120,N_22184);
nand U22305 (N_22305,N_22144,N_22048);
nand U22306 (N_22306,N_22048,N_22194);
or U22307 (N_22307,N_22041,N_22155);
and U22308 (N_22308,N_22132,N_22164);
xor U22309 (N_22309,N_22061,N_22132);
and U22310 (N_22310,N_22193,N_22121);
nand U22311 (N_22311,N_22098,N_22174);
nor U22312 (N_22312,N_22039,N_22195);
nor U22313 (N_22313,N_22101,N_22116);
xnor U22314 (N_22314,N_22095,N_22039);
nand U22315 (N_22315,N_22062,N_22012);
nor U22316 (N_22316,N_22186,N_22037);
nand U22317 (N_22317,N_22055,N_22137);
xnor U22318 (N_22318,N_22091,N_22083);
or U22319 (N_22319,N_22162,N_22021);
nand U22320 (N_22320,N_22053,N_22018);
or U22321 (N_22321,N_22167,N_22034);
nor U22322 (N_22322,N_22005,N_22173);
nand U22323 (N_22323,N_22160,N_22177);
xnor U22324 (N_22324,N_22069,N_22052);
or U22325 (N_22325,N_22093,N_22092);
nor U22326 (N_22326,N_22077,N_22067);
and U22327 (N_22327,N_22164,N_22063);
nand U22328 (N_22328,N_22092,N_22123);
nand U22329 (N_22329,N_22165,N_22091);
nor U22330 (N_22330,N_22026,N_22081);
or U22331 (N_22331,N_22069,N_22086);
nand U22332 (N_22332,N_22050,N_22199);
nor U22333 (N_22333,N_22041,N_22166);
or U22334 (N_22334,N_22159,N_22122);
nor U22335 (N_22335,N_22178,N_22162);
or U22336 (N_22336,N_22120,N_22107);
or U22337 (N_22337,N_22111,N_22157);
nand U22338 (N_22338,N_22035,N_22169);
and U22339 (N_22339,N_22100,N_22044);
xor U22340 (N_22340,N_22040,N_22113);
nor U22341 (N_22341,N_22055,N_22132);
nor U22342 (N_22342,N_22011,N_22081);
or U22343 (N_22343,N_22074,N_22038);
nand U22344 (N_22344,N_22157,N_22182);
nand U22345 (N_22345,N_22017,N_22015);
nand U22346 (N_22346,N_22022,N_22050);
xnor U22347 (N_22347,N_22077,N_22172);
nand U22348 (N_22348,N_22121,N_22129);
xor U22349 (N_22349,N_22019,N_22069);
or U22350 (N_22350,N_22184,N_22078);
nor U22351 (N_22351,N_22118,N_22188);
nor U22352 (N_22352,N_22088,N_22169);
nor U22353 (N_22353,N_22124,N_22073);
or U22354 (N_22354,N_22183,N_22032);
xnor U22355 (N_22355,N_22093,N_22120);
nand U22356 (N_22356,N_22180,N_22184);
nand U22357 (N_22357,N_22003,N_22037);
and U22358 (N_22358,N_22121,N_22043);
nor U22359 (N_22359,N_22172,N_22158);
nand U22360 (N_22360,N_22150,N_22175);
nor U22361 (N_22361,N_22131,N_22063);
and U22362 (N_22362,N_22196,N_22029);
nand U22363 (N_22363,N_22184,N_22090);
or U22364 (N_22364,N_22022,N_22031);
nor U22365 (N_22365,N_22078,N_22084);
or U22366 (N_22366,N_22031,N_22138);
and U22367 (N_22367,N_22158,N_22117);
or U22368 (N_22368,N_22128,N_22153);
nand U22369 (N_22369,N_22011,N_22063);
or U22370 (N_22370,N_22033,N_22050);
and U22371 (N_22371,N_22107,N_22171);
nor U22372 (N_22372,N_22180,N_22117);
nand U22373 (N_22373,N_22031,N_22048);
nor U22374 (N_22374,N_22025,N_22141);
xnor U22375 (N_22375,N_22049,N_22118);
and U22376 (N_22376,N_22175,N_22066);
nand U22377 (N_22377,N_22150,N_22137);
and U22378 (N_22378,N_22088,N_22029);
or U22379 (N_22379,N_22061,N_22139);
or U22380 (N_22380,N_22167,N_22147);
nor U22381 (N_22381,N_22074,N_22064);
and U22382 (N_22382,N_22038,N_22125);
nor U22383 (N_22383,N_22114,N_22118);
xnor U22384 (N_22384,N_22015,N_22073);
and U22385 (N_22385,N_22098,N_22189);
and U22386 (N_22386,N_22049,N_22052);
or U22387 (N_22387,N_22023,N_22155);
xnor U22388 (N_22388,N_22090,N_22192);
and U22389 (N_22389,N_22037,N_22052);
nor U22390 (N_22390,N_22156,N_22145);
xor U22391 (N_22391,N_22199,N_22153);
nand U22392 (N_22392,N_22067,N_22039);
and U22393 (N_22393,N_22067,N_22187);
nor U22394 (N_22394,N_22129,N_22117);
xnor U22395 (N_22395,N_22056,N_22170);
and U22396 (N_22396,N_22045,N_22077);
nor U22397 (N_22397,N_22091,N_22194);
and U22398 (N_22398,N_22144,N_22113);
and U22399 (N_22399,N_22137,N_22174);
nor U22400 (N_22400,N_22323,N_22295);
xor U22401 (N_22401,N_22334,N_22240);
and U22402 (N_22402,N_22338,N_22322);
and U22403 (N_22403,N_22202,N_22301);
and U22404 (N_22404,N_22362,N_22248);
xnor U22405 (N_22405,N_22216,N_22274);
nor U22406 (N_22406,N_22206,N_22311);
nand U22407 (N_22407,N_22374,N_22222);
nor U22408 (N_22408,N_22269,N_22384);
or U22409 (N_22409,N_22379,N_22282);
and U22410 (N_22410,N_22310,N_22306);
nand U22411 (N_22411,N_22387,N_22368);
nand U22412 (N_22412,N_22352,N_22313);
or U22413 (N_22413,N_22326,N_22315);
or U22414 (N_22414,N_22256,N_22314);
xnor U22415 (N_22415,N_22217,N_22383);
nor U22416 (N_22416,N_22258,N_22287);
nor U22417 (N_22417,N_22354,N_22249);
and U22418 (N_22418,N_22307,N_22343);
nor U22419 (N_22419,N_22209,N_22283);
nor U22420 (N_22420,N_22382,N_22257);
and U22421 (N_22421,N_22388,N_22223);
or U22422 (N_22422,N_22275,N_22215);
nand U22423 (N_22423,N_22289,N_22318);
or U22424 (N_22424,N_22228,N_22244);
and U22425 (N_22425,N_22226,N_22279);
nand U22426 (N_22426,N_22270,N_22359);
xnor U22427 (N_22427,N_22300,N_22355);
xor U22428 (N_22428,N_22308,N_22224);
and U22429 (N_22429,N_22357,N_22364);
xnor U22430 (N_22430,N_22261,N_22397);
nor U22431 (N_22431,N_22356,N_22320);
xnor U22432 (N_22432,N_22360,N_22381);
xor U22433 (N_22433,N_22238,N_22259);
nand U22434 (N_22434,N_22376,N_22264);
xnor U22435 (N_22435,N_22278,N_22237);
xor U22436 (N_22436,N_22235,N_22394);
nand U22437 (N_22437,N_22299,N_22207);
nand U22438 (N_22438,N_22366,N_22317);
and U22439 (N_22439,N_22273,N_22233);
xnor U22440 (N_22440,N_22241,N_22230);
nand U22441 (N_22441,N_22292,N_22212);
or U22442 (N_22442,N_22236,N_22377);
and U22443 (N_22443,N_22304,N_22333);
or U22444 (N_22444,N_22312,N_22336);
or U22445 (N_22445,N_22211,N_22385);
or U22446 (N_22446,N_22329,N_22332);
and U22447 (N_22447,N_22243,N_22272);
xor U22448 (N_22448,N_22203,N_22227);
nor U22449 (N_22449,N_22277,N_22386);
xor U22450 (N_22450,N_22219,N_22390);
xnor U22451 (N_22451,N_22225,N_22361);
nand U22452 (N_22452,N_22245,N_22208);
nor U22453 (N_22453,N_22288,N_22345);
or U22454 (N_22454,N_22284,N_22391);
xnor U22455 (N_22455,N_22378,N_22303);
and U22456 (N_22456,N_22204,N_22239);
nand U22457 (N_22457,N_22297,N_22337);
xnor U22458 (N_22458,N_22268,N_22213);
or U22459 (N_22459,N_22395,N_22370);
nand U22460 (N_22460,N_22363,N_22265);
nor U22461 (N_22461,N_22266,N_22302);
nand U22462 (N_22462,N_22260,N_22324);
xnor U22463 (N_22463,N_22296,N_22339);
nor U22464 (N_22464,N_22335,N_22325);
and U22465 (N_22465,N_22305,N_22246);
nor U22466 (N_22466,N_22393,N_22348);
or U22467 (N_22467,N_22350,N_22252);
and U22468 (N_22468,N_22291,N_22342);
nand U22469 (N_22469,N_22263,N_22330);
nor U22470 (N_22470,N_22247,N_22371);
nor U22471 (N_22471,N_22271,N_22328);
nor U22472 (N_22472,N_22367,N_22276);
or U22473 (N_22473,N_22229,N_22220);
or U22474 (N_22474,N_22255,N_22218);
or U22475 (N_22475,N_22293,N_22232);
xnor U22476 (N_22476,N_22353,N_22375);
xnor U22477 (N_22477,N_22205,N_22262);
and U22478 (N_22478,N_22331,N_22221);
or U22479 (N_22479,N_22316,N_22231);
nand U22480 (N_22480,N_22399,N_22250);
nor U22481 (N_22481,N_22286,N_22294);
nand U22482 (N_22482,N_22341,N_22234);
nor U22483 (N_22483,N_22389,N_22372);
nor U22484 (N_22484,N_22242,N_22365);
nor U22485 (N_22485,N_22254,N_22280);
nand U22486 (N_22486,N_22347,N_22253);
nor U22487 (N_22487,N_22210,N_22396);
nand U22488 (N_22488,N_22290,N_22340);
xnor U22489 (N_22489,N_22349,N_22327);
nor U22490 (N_22490,N_22358,N_22351);
or U22491 (N_22491,N_22214,N_22369);
or U22492 (N_22492,N_22380,N_22200);
and U22493 (N_22493,N_22201,N_22267);
or U22494 (N_22494,N_22392,N_22298);
and U22495 (N_22495,N_22281,N_22321);
or U22496 (N_22496,N_22344,N_22285);
or U22497 (N_22497,N_22398,N_22309);
nor U22498 (N_22498,N_22251,N_22346);
nand U22499 (N_22499,N_22373,N_22319);
and U22500 (N_22500,N_22297,N_22267);
nor U22501 (N_22501,N_22323,N_22273);
nor U22502 (N_22502,N_22359,N_22260);
and U22503 (N_22503,N_22341,N_22385);
xor U22504 (N_22504,N_22210,N_22292);
nand U22505 (N_22505,N_22293,N_22262);
and U22506 (N_22506,N_22362,N_22306);
or U22507 (N_22507,N_22272,N_22248);
and U22508 (N_22508,N_22336,N_22268);
nor U22509 (N_22509,N_22312,N_22307);
xor U22510 (N_22510,N_22341,N_22392);
or U22511 (N_22511,N_22240,N_22210);
nand U22512 (N_22512,N_22369,N_22364);
nor U22513 (N_22513,N_22219,N_22307);
xor U22514 (N_22514,N_22392,N_22380);
nor U22515 (N_22515,N_22212,N_22215);
xor U22516 (N_22516,N_22222,N_22370);
and U22517 (N_22517,N_22261,N_22346);
nor U22518 (N_22518,N_22250,N_22276);
nand U22519 (N_22519,N_22240,N_22305);
nor U22520 (N_22520,N_22319,N_22221);
and U22521 (N_22521,N_22344,N_22279);
xor U22522 (N_22522,N_22214,N_22207);
or U22523 (N_22523,N_22387,N_22284);
and U22524 (N_22524,N_22227,N_22368);
or U22525 (N_22525,N_22373,N_22385);
and U22526 (N_22526,N_22291,N_22293);
and U22527 (N_22527,N_22282,N_22237);
nand U22528 (N_22528,N_22312,N_22347);
nand U22529 (N_22529,N_22373,N_22340);
xor U22530 (N_22530,N_22394,N_22265);
nand U22531 (N_22531,N_22262,N_22299);
and U22532 (N_22532,N_22364,N_22390);
or U22533 (N_22533,N_22248,N_22370);
nor U22534 (N_22534,N_22317,N_22310);
or U22535 (N_22535,N_22257,N_22222);
nand U22536 (N_22536,N_22322,N_22309);
or U22537 (N_22537,N_22370,N_22283);
nor U22538 (N_22538,N_22306,N_22335);
and U22539 (N_22539,N_22388,N_22390);
nand U22540 (N_22540,N_22375,N_22357);
xnor U22541 (N_22541,N_22329,N_22207);
and U22542 (N_22542,N_22286,N_22290);
xnor U22543 (N_22543,N_22384,N_22379);
xnor U22544 (N_22544,N_22360,N_22388);
nand U22545 (N_22545,N_22325,N_22203);
nor U22546 (N_22546,N_22390,N_22212);
or U22547 (N_22547,N_22251,N_22252);
xor U22548 (N_22548,N_22284,N_22249);
nor U22549 (N_22549,N_22255,N_22377);
nand U22550 (N_22550,N_22350,N_22335);
or U22551 (N_22551,N_22395,N_22353);
nand U22552 (N_22552,N_22290,N_22323);
xnor U22553 (N_22553,N_22393,N_22215);
and U22554 (N_22554,N_22200,N_22295);
xnor U22555 (N_22555,N_22312,N_22230);
or U22556 (N_22556,N_22212,N_22388);
xor U22557 (N_22557,N_22318,N_22235);
nand U22558 (N_22558,N_22350,N_22216);
nor U22559 (N_22559,N_22242,N_22381);
and U22560 (N_22560,N_22283,N_22330);
nand U22561 (N_22561,N_22344,N_22226);
nor U22562 (N_22562,N_22388,N_22323);
and U22563 (N_22563,N_22215,N_22288);
nor U22564 (N_22564,N_22243,N_22202);
or U22565 (N_22565,N_22371,N_22377);
or U22566 (N_22566,N_22286,N_22234);
nand U22567 (N_22567,N_22232,N_22335);
xnor U22568 (N_22568,N_22311,N_22372);
xor U22569 (N_22569,N_22263,N_22284);
nand U22570 (N_22570,N_22243,N_22294);
xnor U22571 (N_22571,N_22247,N_22216);
and U22572 (N_22572,N_22276,N_22232);
or U22573 (N_22573,N_22207,N_22370);
and U22574 (N_22574,N_22388,N_22373);
or U22575 (N_22575,N_22213,N_22354);
or U22576 (N_22576,N_22298,N_22250);
nor U22577 (N_22577,N_22315,N_22271);
and U22578 (N_22578,N_22274,N_22380);
or U22579 (N_22579,N_22356,N_22222);
and U22580 (N_22580,N_22375,N_22319);
and U22581 (N_22581,N_22328,N_22297);
and U22582 (N_22582,N_22328,N_22295);
nand U22583 (N_22583,N_22213,N_22360);
nand U22584 (N_22584,N_22310,N_22315);
nand U22585 (N_22585,N_22373,N_22278);
and U22586 (N_22586,N_22296,N_22317);
or U22587 (N_22587,N_22332,N_22389);
nor U22588 (N_22588,N_22241,N_22286);
nor U22589 (N_22589,N_22394,N_22324);
or U22590 (N_22590,N_22392,N_22286);
xnor U22591 (N_22591,N_22277,N_22326);
and U22592 (N_22592,N_22215,N_22282);
xnor U22593 (N_22593,N_22266,N_22231);
nand U22594 (N_22594,N_22203,N_22302);
nor U22595 (N_22595,N_22336,N_22298);
and U22596 (N_22596,N_22323,N_22376);
nor U22597 (N_22597,N_22261,N_22260);
or U22598 (N_22598,N_22362,N_22224);
xor U22599 (N_22599,N_22213,N_22274);
xnor U22600 (N_22600,N_22585,N_22533);
xnor U22601 (N_22601,N_22425,N_22518);
nand U22602 (N_22602,N_22475,N_22422);
and U22603 (N_22603,N_22599,N_22462);
nor U22604 (N_22604,N_22589,N_22441);
xor U22605 (N_22605,N_22579,N_22549);
or U22606 (N_22606,N_22497,N_22471);
nor U22607 (N_22607,N_22574,N_22440);
and U22608 (N_22608,N_22584,N_22464);
xor U22609 (N_22609,N_22438,N_22448);
and U22610 (N_22610,N_22528,N_22598);
nand U22611 (N_22611,N_22444,N_22500);
and U22612 (N_22612,N_22530,N_22534);
nor U22613 (N_22613,N_22516,N_22482);
and U22614 (N_22614,N_22423,N_22478);
nand U22615 (N_22615,N_22526,N_22419);
xnor U22616 (N_22616,N_22555,N_22401);
xor U22617 (N_22617,N_22541,N_22458);
nand U22618 (N_22618,N_22537,N_22506);
nand U22619 (N_22619,N_22512,N_22453);
xor U22620 (N_22620,N_22472,N_22413);
or U22621 (N_22621,N_22569,N_22576);
and U22622 (N_22622,N_22470,N_22532);
or U22623 (N_22623,N_22492,N_22446);
nand U22624 (N_22624,N_22447,N_22496);
or U22625 (N_22625,N_22578,N_22522);
nor U22626 (N_22626,N_22494,N_22568);
and U22627 (N_22627,N_22595,N_22567);
nand U22628 (N_22628,N_22424,N_22406);
nand U22629 (N_22629,N_22524,N_22416);
nor U22630 (N_22630,N_22434,N_22490);
nor U22631 (N_22631,N_22433,N_22485);
nor U22632 (N_22632,N_22501,N_22411);
or U22633 (N_22633,N_22479,N_22581);
xnor U22634 (N_22634,N_22551,N_22591);
nor U22635 (N_22635,N_22525,N_22539);
and U22636 (N_22636,N_22410,N_22429);
xnor U22637 (N_22637,N_22445,N_22417);
nor U22638 (N_22638,N_22597,N_22587);
xnor U22639 (N_22639,N_22450,N_22443);
or U22640 (N_22640,N_22586,N_22542);
nand U22641 (N_22641,N_22502,N_22442);
nor U22642 (N_22642,N_22439,N_22565);
and U22643 (N_22643,N_22566,N_22503);
nand U22644 (N_22644,N_22531,N_22452);
and U22645 (N_22645,N_22428,N_22409);
nor U22646 (N_22646,N_22505,N_22513);
xnor U22647 (N_22647,N_22557,N_22572);
nor U22648 (N_22648,N_22449,N_22457);
nand U22649 (N_22649,N_22493,N_22405);
nor U22650 (N_22650,N_22556,N_22466);
or U22651 (N_22651,N_22498,N_22412);
nand U22652 (N_22652,N_22538,N_22517);
nor U22653 (N_22653,N_22536,N_22420);
and U22654 (N_22654,N_22582,N_22511);
or U22655 (N_22655,N_22495,N_22529);
xor U22656 (N_22656,N_22546,N_22510);
xor U22657 (N_22657,N_22575,N_22460);
nand U22658 (N_22658,N_22594,N_22402);
or U22659 (N_22659,N_22459,N_22454);
nor U22660 (N_22660,N_22560,N_22437);
nand U22661 (N_22661,N_22580,N_22456);
nor U22662 (N_22662,N_22507,N_22476);
nor U22663 (N_22663,N_22588,N_22469);
xor U22664 (N_22664,N_22483,N_22535);
or U22665 (N_22665,N_22543,N_22468);
or U22666 (N_22666,N_22415,N_22486);
nor U22667 (N_22667,N_22547,N_22421);
nand U22668 (N_22668,N_22489,N_22583);
or U22669 (N_22669,N_22514,N_22552);
xnor U22670 (N_22670,N_22559,N_22550);
nand U22671 (N_22671,N_22571,N_22484);
and U22672 (N_22672,N_22563,N_22431);
xnor U22673 (N_22673,N_22573,N_22408);
xor U22674 (N_22674,N_22488,N_22593);
and U22675 (N_22675,N_22521,N_22548);
or U22676 (N_22676,N_22558,N_22561);
nand U22677 (N_22677,N_22465,N_22487);
or U22678 (N_22678,N_22430,N_22400);
and U22679 (N_22679,N_22520,N_22407);
xnor U22680 (N_22680,N_22426,N_22461);
and U22681 (N_22681,N_22554,N_22515);
nor U22682 (N_22682,N_22523,N_22481);
nand U22683 (N_22683,N_22509,N_22467);
and U22684 (N_22684,N_22577,N_22477);
nor U22685 (N_22685,N_22480,N_22474);
xor U22686 (N_22686,N_22570,N_22463);
nand U22687 (N_22687,N_22491,N_22404);
nor U22688 (N_22688,N_22436,N_22435);
nor U22689 (N_22689,N_22418,N_22499);
or U22690 (N_22690,N_22519,N_22473);
nor U22691 (N_22691,N_22564,N_22590);
nand U22692 (N_22692,N_22553,N_22403);
and U22693 (N_22693,N_22427,N_22432);
nand U22694 (N_22694,N_22455,N_22592);
xor U22695 (N_22695,N_22527,N_22544);
xnor U22696 (N_22696,N_22596,N_22508);
or U22697 (N_22697,N_22414,N_22504);
xnor U22698 (N_22698,N_22451,N_22540);
and U22699 (N_22699,N_22562,N_22545);
xnor U22700 (N_22700,N_22527,N_22526);
nor U22701 (N_22701,N_22458,N_22572);
xor U22702 (N_22702,N_22449,N_22437);
or U22703 (N_22703,N_22539,N_22508);
and U22704 (N_22704,N_22595,N_22494);
xor U22705 (N_22705,N_22588,N_22591);
nor U22706 (N_22706,N_22419,N_22516);
nand U22707 (N_22707,N_22450,N_22599);
nand U22708 (N_22708,N_22584,N_22423);
xnor U22709 (N_22709,N_22469,N_22473);
or U22710 (N_22710,N_22482,N_22578);
xnor U22711 (N_22711,N_22528,N_22457);
xnor U22712 (N_22712,N_22549,N_22487);
nor U22713 (N_22713,N_22425,N_22525);
or U22714 (N_22714,N_22593,N_22511);
and U22715 (N_22715,N_22427,N_22407);
nand U22716 (N_22716,N_22511,N_22546);
or U22717 (N_22717,N_22493,N_22428);
nor U22718 (N_22718,N_22423,N_22517);
nor U22719 (N_22719,N_22569,N_22560);
nor U22720 (N_22720,N_22469,N_22557);
nand U22721 (N_22721,N_22473,N_22489);
and U22722 (N_22722,N_22489,N_22511);
or U22723 (N_22723,N_22514,N_22473);
or U22724 (N_22724,N_22461,N_22582);
xnor U22725 (N_22725,N_22497,N_22406);
nand U22726 (N_22726,N_22463,N_22420);
and U22727 (N_22727,N_22483,N_22400);
xnor U22728 (N_22728,N_22599,N_22583);
xnor U22729 (N_22729,N_22555,N_22587);
xor U22730 (N_22730,N_22574,N_22568);
xnor U22731 (N_22731,N_22462,N_22529);
and U22732 (N_22732,N_22519,N_22452);
and U22733 (N_22733,N_22583,N_22463);
or U22734 (N_22734,N_22429,N_22539);
nand U22735 (N_22735,N_22560,N_22446);
or U22736 (N_22736,N_22459,N_22587);
nand U22737 (N_22737,N_22414,N_22483);
xnor U22738 (N_22738,N_22570,N_22556);
nor U22739 (N_22739,N_22500,N_22530);
nor U22740 (N_22740,N_22554,N_22477);
xnor U22741 (N_22741,N_22587,N_22550);
xor U22742 (N_22742,N_22573,N_22453);
nor U22743 (N_22743,N_22578,N_22588);
xor U22744 (N_22744,N_22582,N_22465);
nor U22745 (N_22745,N_22445,N_22404);
nor U22746 (N_22746,N_22489,N_22437);
nor U22747 (N_22747,N_22585,N_22423);
nor U22748 (N_22748,N_22576,N_22525);
nand U22749 (N_22749,N_22574,N_22406);
xnor U22750 (N_22750,N_22491,N_22504);
nand U22751 (N_22751,N_22447,N_22599);
nor U22752 (N_22752,N_22438,N_22428);
and U22753 (N_22753,N_22541,N_22507);
xnor U22754 (N_22754,N_22498,N_22547);
xnor U22755 (N_22755,N_22440,N_22470);
xor U22756 (N_22756,N_22531,N_22550);
or U22757 (N_22757,N_22578,N_22497);
xnor U22758 (N_22758,N_22595,N_22500);
nand U22759 (N_22759,N_22562,N_22500);
or U22760 (N_22760,N_22506,N_22436);
or U22761 (N_22761,N_22521,N_22448);
and U22762 (N_22762,N_22583,N_22508);
or U22763 (N_22763,N_22481,N_22432);
nand U22764 (N_22764,N_22425,N_22443);
nand U22765 (N_22765,N_22530,N_22539);
or U22766 (N_22766,N_22588,N_22531);
nand U22767 (N_22767,N_22476,N_22492);
nor U22768 (N_22768,N_22576,N_22515);
xnor U22769 (N_22769,N_22463,N_22419);
and U22770 (N_22770,N_22452,N_22560);
and U22771 (N_22771,N_22458,N_22598);
and U22772 (N_22772,N_22422,N_22447);
and U22773 (N_22773,N_22520,N_22439);
xor U22774 (N_22774,N_22515,N_22538);
or U22775 (N_22775,N_22410,N_22416);
nor U22776 (N_22776,N_22433,N_22546);
nor U22777 (N_22777,N_22473,N_22432);
and U22778 (N_22778,N_22503,N_22572);
nor U22779 (N_22779,N_22470,N_22515);
nor U22780 (N_22780,N_22406,N_22415);
nor U22781 (N_22781,N_22544,N_22456);
nor U22782 (N_22782,N_22593,N_22515);
nand U22783 (N_22783,N_22477,N_22404);
nand U22784 (N_22784,N_22430,N_22465);
xor U22785 (N_22785,N_22523,N_22497);
or U22786 (N_22786,N_22438,N_22573);
nor U22787 (N_22787,N_22424,N_22450);
nand U22788 (N_22788,N_22424,N_22544);
nand U22789 (N_22789,N_22404,N_22416);
or U22790 (N_22790,N_22579,N_22560);
nand U22791 (N_22791,N_22506,N_22491);
nor U22792 (N_22792,N_22581,N_22518);
nand U22793 (N_22793,N_22579,N_22541);
xnor U22794 (N_22794,N_22408,N_22593);
xnor U22795 (N_22795,N_22458,N_22464);
nand U22796 (N_22796,N_22475,N_22562);
nor U22797 (N_22797,N_22477,N_22591);
or U22798 (N_22798,N_22453,N_22418);
or U22799 (N_22799,N_22435,N_22597);
and U22800 (N_22800,N_22700,N_22738);
and U22801 (N_22801,N_22642,N_22773);
nand U22802 (N_22802,N_22695,N_22718);
xor U22803 (N_22803,N_22617,N_22768);
nor U22804 (N_22804,N_22765,N_22601);
nand U22805 (N_22805,N_22648,N_22677);
nand U22806 (N_22806,N_22781,N_22722);
and U22807 (N_22807,N_22797,N_22697);
and U22808 (N_22808,N_22782,N_22669);
and U22809 (N_22809,N_22796,N_22712);
or U22810 (N_22810,N_22736,N_22769);
nor U22811 (N_22811,N_22659,N_22683);
or U22812 (N_22812,N_22685,N_22649);
or U22813 (N_22813,N_22614,N_22671);
nand U22814 (N_22814,N_22689,N_22670);
or U22815 (N_22815,N_22682,N_22772);
and U22816 (N_22816,N_22710,N_22643);
or U22817 (N_22817,N_22748,N_22739);
xnor U22818 (N_22818,N_22656,N_22666);
or U22819 (N_22819,N_22779,N_22668);
nand U22820 (N_22820,N_22663,N_22654);
xor U22821 (N_22821,N_22693,N_22618);
and U22822 (N_22822,N_22747,N_22639);
or U22823 (N_22823,N_22730,N_22713);
xor U22824 (N_22824,N_22717,N_22758);
nand U22825 (N_22825,N_22799,N_22719);
and U22826 (N_22826,N_22625,N_22667);
xor U22827 (N_22827,N_22792,N_22664);
xor U22828 (N_22828,N_22752,N_22637);
nand U22829 (N_22829,N_22749,N_22774);
nor U22830 (N_22830,N_22658,N_22626);
nor U22831 (N_22831,N_22657,N_22771);
xor U22832 (N_22832,N_22651,N_22731);
or U22833 (N_22833,N_22624,N_22699);
xnor U22834 (N_22834,N_22628,N_22737);
or U22835 (N_22835,N_22784,N_22704);
or U22836 (N_22836,N_22761,N_22673);
nand U22837 (N_22837,N_22726,N_22616);
or U22838 (N_22838,N_22687,N_22759);
and U22839 (N_22839,N_22607,N_22764);
nor U22840 (N_22840,N_22729,N_22679);
or U22841 (N_22841,N_22775,N_22696);
xnor U22842 (N_22842,N_22611,N_22684);
xnor U22843 (N_22843,N_22635,N_22785);
nor U22844 (N_22844,N_22640,N_22794);
xor U22845 (N_22845,N_22692,N_22798);
xnor U22846 (N_22846,N_22606,N_22688);
xnor U22847 (N_22847,N_22707,N_22778);
xnor U22848 (N_22848,N_22647,N_22740);
and U22849 (N_22849,N_22724,N_22706);
or U22850 (N_22850,N_22727,N_22620);
nand U22851 (N_22851,N_22690,N_22742);
or U22852 (N_22852,N_22615,N_22762);
and U22853 (N_22853,N_22608,N_22708);
or U22854 (N_22854,N_22653,N_22680);
or U22855 (N_22855,N_22750,N_22788);
nand U22856 (N_22856,N_22665,N_22753);
or U22857 (N_22857,N_22686,N_22645);
nor U22858 (N_22858,N_22709,N_22627);
and U22859 (N_22859,N_22732,N_22770);
nor U22860 (N_22860,N_22723,N_22791);
nand U22861 (N_22861,N_22734,N_22623);
xor U22862 (N_22862,N_22603,N_22698);
and U22863 (N_22863,N_22678,N_22681);
nand U22864 (N_22864,N_22605,N_22725);
or U22865 (N_22865,N_22609,N_22760);
xnor U22866 (N_22866,N_22789,N_22720);
xor U22867 (N_22867,N_22650,N_22741);
and U22868 (N_22868,N_22610,N_22672);
or U22869 (N_22869,N_22641,N_22613);
nor U22870 (N_22870,N_22600,N_22780);
and U22871 (N_22871,N_22602,N_22795);
nor U22872 (N_22872,N_22745,N_22676);
and U22873 (N_22873,N_22646,N_22644);
and U22874 (N_22874,N_22702,N_22751);
xnor U22875 (N_22875,N_22754,N_22691);
nand U22876 (N_22876,N_22660,N_22735);
nor U22877 (N_22877,N_22756,N_22636);
nor U22878 (N_22878,N_22743,N_22790);
nor U22879 (N_22879,N_22662,N_22629);
nand U22880 (N_22880,N_22793,N_22728);
nor U22881 (N_22881,N_22783,N_22757);
or U22882 (N_22882,N_22711,N_22675);
or U22883 (N_22883,N_22612,N_22634);
nor U22884 (N_22884,N_22621,N_22787);
nand U22885 (N_22885,N_22604,N_22674);
xor U22886 (N_22886,N_22733,N_22786);
and U22887 (N_22887,N_22777,N_22776);
and U22888 (N_22888,N_22619,N_22721);
nor U22889 (N_22889,N_22622,N_22652);
nor U22890 (N_22890,N_22633,N_22755);
nand U22891 (N_22891,N_22714,N_22638);
or U22892 (N_22892,N_22715,N_22655);
xnor U22893 (N_22893,N_22746,N_22716);
nor U22894 (N_22894,N_22661,N_22705);
xnor U22895 (N_22895,N_22632,N_22694);
nand U22896 (N_22896,N_22766,N_22631);
and U22897 (N_22897,N_22744,N_22703);
xnor U22898 (N_22898,N_22763,N_22767);
or U22899 (N_22899,N_22630,N_22701);
nand U22900 (N_22900,N_22679,N_22663);
and U22901 (N_22901,N_22604,N_22606);
xor U22902 (N_22902,N_22649,N_22700);
or U22903 (N_22903,N_22602,N_22698);
nor U22904 (N_22904,N_22629,N_22717);
xor U22905 (N_22905,N_22713,N_22637);
xor U22906 (N_22906,N_22674,N_22743);
or U22907 (N_22907,N_22773,N_22781);
nand U22908 (N_22908,N_22728,N_22667);
nor U22909 (N_22909,N_22733,N_22667);
xor U22910 (N_22910,N_22791,N_22738);
xnor U22911 (N_22911,N_22758,N_22786);
or U22912 (N_22912,N_22781,N_22658);
and U22913 (N_22913,N_22654,N_22785);
xnor U22914 (N_22914,N_22671,N_22680);
nand U22915 (N_22915,N_22618,N_22640);
nand U22916 (N_22916,N_22744,N_22691);
and U22917 (N_22917,N_22623,N_22758);
nand U22918 (N_22918,N_22659,N_22751);
and U22919 (N_22919,N_22648,N_22745);
xnor U22920 (N_22920,N_22693,N_22630);
nor U22921 (N_22921,N_22627,N_22628);
or U22922 (N_22922,N_22659,N_22788);
or U22923 (N_22923,N_22716,N_22628);
nor U22924 (N_22924,N_22637,N_22612);
nor U22925 (N_22925,N_22637,N_22734);
nor U22926 (N_22926,N_22756,N_22706);
nor U22927 (N_22927,N_22774,N_22756);
or U22928 (N_22928,N_22735,N_22626);
xnor U22929 (N_22929,N_22716,N_22717);
or U22930 (N_22930,N_22779,N_22687);
nor U22931 (N_22931,N_22696,N_22627);
xnor U22932 (N_22932,N_22605,N_22629);
or U22933 (N_22933,N_22717,N_22752);
or U22934 (N_22934,N_22640,N_22730);
and U22935 (N_22935,N_22709,N_22695);
xnor U22936 (N_22936,N_22729,N_22742);
xor U22937 (N_22937,N_22691,N_22626);
and U22938 (N_22938,N_22769,N_22681);
nor U22939 (N_22939,N_22666,N_22734);
xnor U22940 (N_22940,N_22795,N_22616);
nand U22941 (N_22941,N_22710,N_22704);
and U22942 (N_22942,N_22662,N_22659);
or U22943 (N_22943,N_22723,N_22767);
xor U22944 (N_22944,N_22798,N_22650);
and U22945 (N_22945,N_22771,N_22617);
nand U22946 (N_22946,N_22714,N_22684);
nand U22947 (N_22947,N_22766,N_22681);
nor U22948 (N_22948,N_22637,N_22759);
xor U22949 (N_22949,N_22730,N_22666);
and U22950 (N_22950,N_22630,N_22700);
and U22951 (N_22951,N_22742,N_22611);
nand U22952 (N_22952,N_22655,N_22616);
and U22953 (N_22953,N_22603,N_22704);
nand U22954 (N_22954,N_22762,N_22744);
nand U22955 (N_22955,N_22736,N_22619);
and U22956 (N_22956,N_22778,N_22729);
nor U22957 (N_22957,N_22777,N_22601);
or U22958 (N_22958,N_22613,N_22608);
nand U22959 (N_22959,N_22799,N_22664);
nand U22960 (N_22960,N_22652,N_22753);
xor U22961 (N_22961,N_22620,N_22742);
nor U22962 (N_22962,N_22725,N_22675);
xnor U22963 (N_22963,N_22788,N_22798);
and U22964 (N_22964,N_22785,N_22744);
and U22965 (N_22965,N_22659,N_22743);
and U22966 (N_22966,N_22644,N_22729);
and U22967 (N_22967,N_22627,N_22642);
or U22968 (N_22968,N_22675,N_22667);
nand U22969 (N_22969,N_22650,N_22746);
nand U22970 (N_22970,N_22759,N_22636);
nand U22971 (N_22971,N_22715,N_22736);
xnor U22972 (N_22972,N_22708,N_22676);
and U22973 (N_22973,N_22783,N_22637);
or U22974 (N_22974,N_22627,N_22725);
nor U22975 (N_22975,N_22656,N_22645);
or U22976 (N_22976,N_22632,N_22626);
nand U22977 (N_22977,N_22623,N_22683);
nand U22978 (N_22978,N_22714,N_22744);
or U22979 (N_22979,N_22739,N_22774);
and U22980 (N_22980,N_22755,N_22661);
nand U22981 (N_22981,N_22664,N_22709);
nand U22982 (N_22982,N_22667,N_22657);
nand U22983 (N_22983,N_22779,N_22702);
xnor U22984 (N_22984,N_22605,N_22643);
and U22985 (N_22985,N_22671,N_22679);
nor U22986 (N_22986,N_22657,N_22712);
and U22987 (N_22987,N_22751,N_22687);
nand U22988 (N_22988,N_22673,N_22774);
or U22989 (N_22989,N_22733,N_22773);
nand U22990 (N_22990,N_22655,N_22665);
and U22991 (N_22991,N_22732,N_22681);
nor U22992 (N_22992,N_22727,N_22785);
and U22993 (N_22993,N_22690,N_22783);
nand U22994 (N_22994,N_22652,N_22791);
or U22995 (N_22995,N_22610,N_22765);
or U22996 (N_22996,N_22677,N_22687);
xor U22997 (N_22997,N_22711,N_22633);
nor U22998 (N_22998,N_22649,N_22743);
or U22999 (N_22999,N_22662,N_22637);
and U23000 (N_23000,N_22845,N_22835);
and U23001 (N_23001,N_22940,N_22859);
and U23002 (N_23002,N_22929,N_22837);
or U23003 (N_23003,N_22867,N_22802);
and U23004 (N_23004,N_22925,N_22995);
and U23005 (N_23005,N_22877,N_22904);
nor U23006 (N_23006,N_22818,N_22976);
nor U23007 (N_23007,N_22833,N_22896);
and U23008 (N_23008,N_22879,N_22924);
nor U23009 (N_23009,N_22905,N_22963);
and U23010 (N_23010,N_22913,N_22987);
nor U23011 (N_23011,N_22914,N_22897);
nor U23012 (N_23012,N_22858,N_22942);
and U23013 (N_23013,N_22803,N_22964);
xor U23014 (N_23014,N_22884,N_22809);
nand U23015 (N_23015,N_22825,N_22861);
nor U23016 (N_23016,N_22908,N_22923);
and U23017 (N_23017,N_22930,N_22812);
or U23018 (N_23018,N_22902,N_22873);
nand U23019 (N_23019,N_22842,N_22891);
xor U23020 (N_23020,N_22814,N_22811);
or U23021 (N_23021,N_22815,N_22821);
or U23022 (N_23022,N_22996,N_22838);
and U23023 (N_23023,N_22903,N_22881);
nand U23024 (N_23024,N_22848,N_22950);
nand U23025 (N_23025,N_22936,N_22979);
nor U23026 (N_23026,N_22952,N_22933);
and U23027 (N_23027,N_22941,N_22959);
xor U23028 (N_23028,N_22946,N_22882);
and U23029 (N_23029,N_22975,N_22851);
or U23030 (N_23030,N_22868,N_22980);
nor U23031 (N_23031,N_22869,N_22917);
and U23032 (N_23032,N_22834,N_22958);
and U23033 (N_23033,N_22938,N_22919);
or U23034 (N_23034,N_22824,N_22910);
xnor U23035 (N_23035,N_22943,N_22816);
or U23036 (N_23036,N_22874,N_22830);
xnor U23037 (N_23037,N_22954,N_22886);
nor U23038 (N_23038,N_22887,N_22895);
nor U23039 (N_23039,N_22932,N_22931);
or U23040 (N_23040,N_22900,N_22988);
or U23041 (N_23041,N_22850,N_22991);
xnor U23042 (N_23042,N_22928,N_22955);
xor U23043 (N_23043,N_22860,N_22819);
nand U23044 (N_23044,N_22981,N_22966);
and U23045 (N_23045,N_22957,N_22915);
nor U23046 (N_23046,N_22918,N_22986);
and U23047 (N_23047,N_22994,N_22898);
nor U23048 (N_23048,N_22927,N_22989);
xor U23049 (N_23049,N_22998,N_22862);
or U23050 (N_23050,N_22856,N_22890);
nor U23051 (N_23051,N_22870,N_22984);
or U23052 (N_23052,N_22956,N_22899);
or U23053 (N_23053,N_22926,N_22885);
nand U23054 (N_23054,N_22973,N_22852);
or U23055 (N_23055,N_22997,N_22935);
xor U23056 (N_23056,N_22863,N_22800);
or U23057 (N_23057,N_22962,N_22916);
and U23058 (N_23058,N_22965,N_22846);
or U23059 (N_23059,N_22921,N_22970);
nand U23060 (N_23060,N_22808,N_22827);
nor U23061 (N_23061,N_22912,N_22883);
nand U23062 (N_23062,N_22967,N_22826);
and U23063 (N_23063,N_22971,N_22872);
or U23064 (N_23064,N_22960,N_22836);
and U23065 (N_23065,N_22847,N_22961);
and U23066 (N_23066,N_22880,N_22985);
nor U23067 (N_23067,N_22878,N_22969);
xor U23068 (N_23068,N_22937,N_22944);
xor U23069 (N_23069,N_22990,N_22901);
and U23070 (N_23070,N_22977,N_22853);
nor U23071 (N_23071,N_22934,N_22951);
xnor U23072 (N_23072,N_22828,N_22823);
nor U23073 (N_23073,N_22855,N_22841);
or U23074 (N_23074,N_22953,N_22947);
nor U23075 (N_23075,N_22894,N_22871);
or U23076 (N_23076,N_22822,N_22864);
or U23077 (N_23077,N_22807,N_22840);
nand U23078 (N_23078,N_22906,N_22999);
or U23079 (N_23079,N_22865,N_22839);
nor U23080 (N_23080,N_22857,N_22854);
nor U23081 (N_23081,N_22939,N_22810);
nand U23082 (N_23082,N_22876,N_22866);
or U23083 (N_23083,N_22922,N_22911);
nor U23084 (N_23084,N_22843,N_22893);
nor U23085 (N_23085,N_22805,N_22817);
xnor U23086 (N_23086,N_22978,N_22804);
nor U23087 (N_23087,N_22993,N_22945);
nor U23088 (N_23088,N_22968,N_22948);
nand U23089 (N_23089,N_22801,N_22982);
and U23090 (N_23090,N_22844,N_22909);
or U23091 (N_23091,N_22849,N_22949);
and U23092 (N_23092,N_22832,N_22992);
nand U23093 (N_23093,N_22820,N_22974);
nor U23094 (N_23094,N_22875,N_22831);
xor U23095 (N_23095,N_22892,N_22829);
or U23096 (N_23096,N_22907,N_22813);
nor U23097 (N_23097,N_22920,N_22889);
xnor U23098 (N_23098,N_22888,N_22806);
nor U23099 (N_23099,N_22983,N_22972);
nor U23100 (N_23100,N_22840,N_22947);
and U23101 (N_23101,N_22802,N_22882);
and U23102 (N_23102,N_22881,N_22866);
xnor U23103 (N_23103,N_22874,N_22986);
xor U23104 (N_23104,N_22971,N_22813);
nor U23105 (N_23105,N_22873,N_22910);
nand U23106 (N_23106,N_22819,N_22919);
xnor U23107 (N_23107,N_22959,N_22922);
nor U23108 (N_23108,N_22853,N_22948);
nand U23109 (N_23109,N_22880,N_22850);
and U23110 (N_23110,N_22958,N_22883);
or U23111 (N_23111,N_22830,N_22902);
xnor U23112 (N_23112,N_22929,N_22941);
or U23113 (N_23113,N_22941,N_22885);
nand U23114 (N_23114,N_22888,N_22948);
or U23115 (N_23115,N_22845,N_22976);
and U23116 (N_23116,N_22827,N_22824);
and U23117 (N_23117,N_22892,N_22879);
or U23118 (N_23118,N_22820,N_22813);
nand U23119 (N_23119,N_22919,N_22914);
nor U23120 (N_23120,N_22835,N_22859);
nand U23121 (N_23121,N_22862,N_22973);
nor U23122 (N_23122,N_22927,N_22898);
nand U23123 (N_23123,N_22980,N_22978);
or U23124 (N_23124,N_22918,N_22835);
xnor U23125 (N_23125,N_22951,N_22854);
xor U23126 (N_23126,N_22831,N_22902);
nand U23127 (N_23127,N_22982,N_22991);
nor U23128 (N_23128,N_22878,N_22838);
or U23129 (N_23129,N_22933,N_22882);
or U23130 (N_23130,N_22822,N_22981);
xor U23131 (N_23131,N_22860,N_22914);
xnor U23132 (N_23132,N_22853,N_22946);
or U23133 (N_23133,N_22886,N_22961);
and U23134 (N_23134,N_22853,N_22961);
xnor U23135 (N_23135,N_22850,N_22833);
nor U23136 (N_23136,N_22990,N_22981);
nand U23137 (N_23137,N_22804,N_22990);
xor U23138 (N_23138,N_22994,N_22893);
nand U23139 (N_23139,N_22877,N_22989);
or U23140 (N_23140,N_22931,N_22881);
nand U23141 (N_23141,N_22967,N_22893);
nor U23142 (N_23142,N_22944,N_22831);
and U23143 (N_23143,N_22938,N_22907);
and U23144 (N_23144,N_22985,N_22948);
or U23145 (N_23145,N_22963,N_22871);
nand U23146 (N_23146,N_22984,N_22932);
nand U23147 (N_23147,N_22803,N_22933);
or U23148 (N_23148,N_22903,N_22877);
nand U23149 (N_23149,N_22979,N_22997);
or U23150 (N_23150,N_22989,N_22956);
nand U23151 (N_23151,N_22892,N_22802);
and U23152 (N_23152,N_22958,N_22846);
nand U23153 (N_23153,N_22896,N_22879);
xor U23154 (N_23154,N_22853,N_22817);
and U23155 (N_23155,N_22898,N_22888);
and U23156 (N_23156,N_22919,N_22908);
nor U23157 (N_23157,N_22970,N_22842);
and U23158 (N_23158,N_22956,N_22969);
or U23159 (N_23159,N_22862,N_22893);
nor U23160 (N_23160,N_22886,N_22967);
and U23161 (N_23161,N_22994,N_22813);
and U23162 (N_23162,N_22980,N_22881);
or U23163 (N_23163,N_22811,N_22945);
or U23164 (N_23164,N_22811,N_22898);
nor U23165 (N_23165,N_22801,N_22966);
or U23166 (N_23166,N_22801,N_22920);
xor U23167 (N_23167,N_22914,N_22855);
xor U23168 (N_23168,N_22974,N_22937);
nand U23169 (N_23169,N_22892,N_22917);
nand U23170 (N_23170,N_22852,N_22912);
and U23171 (N_23171,N_22821,N_22830);
xor U23172 (N_23172,N_22956,N_22893);
nor U23173 (N_23173,N_22995,N_22802);
nand U23174 (N_23174,N_22888,N_22899);
xnor U23175 (N_23175,N_22985,N_22823);
nor U23176 (N_23176,N_22960,N_22990);
xor U23177 (N_23177,N_22873,N_22861);
nand U23178 (N_23178,N_22815,N_22918);
nand U23179 (N_23179,N_22885,N_22804);
xor U23180 (N_23180,N_22822,N_22890);
or U23181 (N_23181,N_22938,N_22979);
and U23182 (N_23182,N_22846,N_22867);
and U23183 (N_23183,N_22818,N_22828);
xor U23184 (N_23184,N_22879,N_22968);
and U23185 (N_23185,N_22956,N_22839);
xor U23186 (N_23186,N_22891,N_22992);
and U23187 (N_23187,N_22896,N_22986);
and U23188 (N_23188,N_22897,N_22825);
and U23189 (N_23189,N_22887,N_22888);
nor U23190 (N_23190,N_22883,N_22972);
nor U23191 (N_23191,N_22853,N_22900);
or U23192 (N_23192,N_22869,N_22946);
nand U23193 (N_23193,N_22853,N_22952);
and U23194 (N_23194,N_22870,N_22902);
or U23195 (N_23195,N_22848,N_22953);
or U23196 (N_23196,N_22971,N_22966);
nand U23197 (N_23197,N_22892,N_22833);
xnor U23198 (N_23198,N_22937,N_22852);
or U23199 (N_23199,N_22859,N_22962);
nor U23200 (N_23200,N_23017,N_23027);
nor U23201 (N_23201,N_23086,N_23112);
or U23202 (N_23202,N_23128,N_23108);
nand U23203 (N_23203,N_23154,N_23015);
and U23204 (N_23204,N_23087,N_23130);
and U23205 (N_23205,N_23095,N_23030);
and U23206 (N_23206,N_23094,N_23120);
nor U23207 (N_23207,N_23136,N_23054);
or U23208 (N_23208,N_23193,N_23036);
xor U23209 (N_23209,N_23060,N_23038);
and U23210 (N_23210,N_23135,N_23126);
xor U23211 (N_23211,N_23171,N_23146);
nand U23212 (N_23212,N_23149,N_23153);
or U23213 (N_23213,N_23031,N_23152);
nand U23214 (N_23214,N_23023,N_23144);
and U23215 (N_23215,N_23110,N_23026);
and U23216 (N_23216,N_23088,N_23091);
nand U23217 (N_23217,N_23151,N_23082);
nand U23218 (N_23218,N_23113,N_23143);
nor U23219 (N_23219,N_23070,N_23150);
nor U23220 (N_23220,N_23174,N_23142);
nor U23221 (N_23221,N_23049,N_23185);
xnor U23222 (N_23222,N_23055,N_23067);
xnor U23223 (N_23223,N_23040,N_23119);
nand U23224 (N_23224,N_23177,N_23047);
nor U23225 (N_23225,N_23106,N_23034);
xor U23226 (N_23226,N_23008,N_23168);
nor U23227 (N_23227,N_23050,N_23039);
xnor U23228 (N_23228,N_23041,N_23084);
nand U23229 (N_23229,N_23102,N_23187);
nand U23230 (N_23230,N_23134,N_23073);
nand U23231 (N_23231,N_23190,N_23096);
and U23232 (N_23232,N_23021,N_23122);
nor U23233 (N_23233,N_23160,N_23057);
nor U23234 (N_23234,N_23103,N_23127);
nor U23235 (N_23235,N_23059,N_23183);
nand U23236 (N_23236,N_23001,N_23139);
or U23237 (N_23237,N_23098,N_23131);
and U23238 (N_23238,N_23148,N_23129);
and U23239 (N_23239,N_23158,N_23077);
xor U23240 (N_23240,N_23051,N_23018);
and U23241 (N_23241,N_23081,N_23186);
or U23242 (N_23242,N_23033,N_23022);
and U23243 (N_23243,N_23125,N_23156);
or U23244 (N_23244,N_23014,N_23191);
and U23245 (N_23245,N_23074,N_23024);
xor U23246 (N_23246,N_23012,N_23192);
xnor U23247 (N_23247,N_23184,N_23002);
or U23248 (N_23248,N_23044,N_23043);
or U23249 (N_23249,N_23180,N_23011);
and U23250 (N_23250,N_23104,N_23181);
nor U23251 (N_23251,N_23111,N_23075);
nor U23252 (N_23252,N_23164,N_23078);
or U23253 (N_23253,N_23035,N_23197);
or U23254 (N_23254,N_23006,N_23046);
nor U23255 (N_23255,N_23132,N_23198);
nand U23256 (N_23256,N_23037,N_23083);
nand U23257 (N_23257,N_23071,N_23165);
or U23258 (N_23258,N_23173,N_23056);
or U23259 (N_23259,N_23053,N_23009);
and U23260 (N_23260,N_23116,N_23005);
and U23261 (N_23261,N_23194,N_23080);
nor U23262 (N_23262,N_23137,N_23166);
xnor U23263 (N_23263,N_23032,N_23161);
or U23264 (N_23264,N_23175,N_23118);
or U23265 (N_23265,N_23147,N_23007);
nand U23266 (N_23266,N_23117,N_23016);
or U23267 (N_23267,N_23072,N_23019);
and U23268 (N_23268,N_23155,N_23107);
or U23269 (N_23269,N_23061,N_23097);
nand U23270 (N_23270,N_23099,N_23188);
and U23271 (N_23271,N_23114,N_23068);
and U23272 (N_23272,N_23189,N_23090);
xor U23273 (N_23273,N_23100,N_23101);
and U23274 (N_23274,N_23092,N_23138);
and U23275 (N_23275,N_23124,N_23163);
or U23276 (N_23276,N_23025,N_23093);
nand U23277 (N_23277,N_23176,N_23066);
nand U23278 (N_23278,N_23199,N_23195);
nor U23279 (N_23279,N_23079,N_23157);
nor U23280 (N_23280,N_23020,N_23109);
nor U23281 (N_23281,N_23048,N_23076);
nand U23282 (N_23282,N_23115,N_23123);
or U23283 (N_23283,N_23058,N_23169);
xnor U23284 (N_23284,N_23162,N_23121);
nor U23285 (N_23285,N_23170,N_23029);
nand U23286 (N_23286,N_23196,N_23004);
or U23287 (N_23287,N_23062,N_23089);
nand U23288 (N_23288,N_23010,N_23028);
nand U23289 (N_23289,N_23167,N_23178);
xor U23290 (N_23290,N_23085,N_23042);
nand U23291 (N_23291,N_23069,N_23179);
nor U23292 (N_23292,N_23063,N_23172);
or U23293 (N_23293,N_23045,N_23000);
nand U23294 (N_23294,N_23052,N_23159);
nand U23295 (N_23295,N_23182,N_23064);
or U23296 (N_23296,N_23145,N_23065);
nor U23297 (N_23297,N_23003,N_23141);
xnor U23298 (N_23298,N_23105,N_23140);
nor U23299 (N_23299,N_23013,N_23133);
xor U23300 (N_23300,N_23160,N_23117);
and U23301 (N_23301,N_23152,N_23179);
and U23302 (N_23302,N_23133,N_23069);
nor U23303 (N_23303,N_23130,N_23111);
and U23304 (N_23304,N_23023,N_23179);
xor U23305 (N_23305,N_23111,N_23006);
xnor U23306 (N_23306,N_23073,N_23160);
and U23307 (N_23307,N_23043,N_23038);
xnor U23308 (N_23308,N_23097,N_23113);
nand U23309 (N_23309,N_23064,N_23129);
xnor U23310 (N_23310,N_23192,N_23064);
nor U23311 (N_23311,N_23119,N_23156);
and U23312 (N_23312,N_23191,N_23023);
and U23313 (N_23313,N_23150,N_23092);
xor U23314 (N_23314,N_23060,N_23138);
xor U23315 (N_23315,N_23035,N_23101);
or U23316 (N_23316,N_23006,N_23147);
or U23317 (N_23317,N_23102,N_23037);
nor U23318 (N_23318,N_23102,N_23118);
nand U23319 (N_23319,N_23024,N_23169);
and U23320 (N_23320,N_23020,N_23142);
nor U23321 (N_23321,N_23026,N_23116);
xnor U23322 (N_23322,N_23097,N_23149);
and U23323 (N_23323,N_23071,N_23028);
nor U23324 (N_23324,N_23105,N_23048);
xor U23325 (N_23325,N_23194,N_23068);
xnor U23326 (N_23326,N_23112,N_23108);
nand U23327 (N_23327,N_23037,N_23131);
or U23328 (N_23328,N_23151,N_23099);
nor U23329 (N_23329,N_23138,N_23043);
nand U23330 (N_23330,N_23048,N_23037);
and U23331 (N_23331,N_23014,N_23037);
nand U23332 (N_23332,N_23016,N_23137);
nor U23333 (N_23333,N_23112,N_23043);
nor U23334 (N_23334,N_23135,N_23143);
nor U23335 (N_23335,N_23155,N_23163);
xnor U23336 (N_23336,N_23186,N_23033);
nand U23337 (N_23337,N_23073,N_23067);
xor U23338 (N_23338,N_23160,N_23063);
and U23339 (N_23339,N_23096,N_23097);
nand U23340 (N_23340,N_23198,N_23190);
nor U23341 (N_23341,N_23166,N_23170);
nand U23342 (N_23342,N_23020,N_23183);
nand U23343 (N_23343,N_23196,N_23163);
xnor U23344 (N_23344,N_23032,N_23158);
nor U23345 (N_23345,N_23124,N_23086);
and U23346 (N_23346,N_23195,N_23077);
nor U23347 (N_23347,N_23147,N_23001);
and U23348 (N_23348,N_23144,N_23194);
or U23349 (N_23349,N_23038,N_23029);
or U23350 (N_23350,N_23027,N_23062);
or U23351 (N_23351,N_23056,N_23126);
nor U23352 (N_23352,N_23081,N_23030);
nand U23353 (N_23353,N_23039,N_23080);
nand U23354 (N_23354,N_23164,N_23185);
or U23355 (N_23355,N_23051,N_23067);
and U23356 (N_23356,N_23012,N_23110);
or U23357 (N_23357,N_23103,N_23085);
xor U23358 (N_23358,N_23154,N_23060);
or U23359 (N_23359,N_23179,N_23164);
xnor U23360 (N_23360,N_23189,N_23152);
nand U23361 (N_23361,N_23161,N_23112);
nand U23362 (N_23362,N_23079,N_23013);
nand U23363 (N_23363,N_23055,N_23126);
and U23364 (N_23364,N_23155,N_23192);
xor U23365 (N_23365,N_23156,N_23090);
and U23366 (N_23366,N_23159,N_23124);
or U23367 (N_23367,N_23148,N_23011);
xor U23368 (N_23368,N_23180,N_23130);
or U23369 (N_23369,N_23065,N_23155);
xor U23370 (N_23370,N_23098,N_23011);
nand U23371 (N_23371,N_23173,N_23150);
and U23372 (N_23372,N_23041,N_23133);
and U23373 (N_23373,N_23151,N_23025);
and U23374 (N_23374,N_23062,N_23041);
or U23375 (N_23375,N_23194,N_23139);
nor U23376 (N_23376,N_23122,N_23045);
or U23377 (N_23377,N_23045,N_23002);
and U23378 (N_23378,N_23029,N_23043);
or U23379 (N_23379,N_23162,N_23028);
nand U23380 (N_23380,N_23010,N_23148);
nor U23381 (N_23381,N_23172,N_23155);
and U23382 (N_23382,N_23069,N_23111);
or U23383 (N_23383,N_23145,N_23100);
xnor U23384 (N_23384,N_23178,N_23164);
and U23385 (N_23385,N_23183,N_23058);
nor U23386 (N_23386,N_23036,N_23150);
xnor U23387 (N_23387,N_23064,N_23007);
or U23388 (N_23388,N_23160,N_23092);
nand U23389 (N_23389,N_23163,N_23112);
nand U23390 (N_23390,N_23139,N_23146);
xor U23391 (N_23391,N_23030,N_23067);
nor U23392 (N_23392,N_23018,N_23191);
and U23393 (N_23393,N_23009,N_23189);
xnor U23394 (N_23394,N_23083,N_23047);
xnor U23395 (N_23395,N_23193,N_23083);
xnor U23396 (N_23396,N_23000,N_23140);
and U23397 (N_23397,N_23038,N_23152);
nand U23398 (N_23398,N_23081,N_23188);
nor U23399 (N_23399,N_23063,N_23175);
nand U23400 (N_23400,N_23223,N_23269);
and U23401 (N_23401,N_23317,N_23278);
nor U23402 (N_23402,N_23312,N_23396);
nor U23403 (N_23403,N_23287,N_23282);
nor U23404 (N_23404,N_23356,N_23375);
nor U23405 (N_23405,N_23235,N_23342);
xor U23406 (N_23406,N_23306,N_23368);
xnor U23407 (N_23407,N_23211,N_23297);
xnor U23408 (N_23408,N_23380,N_23343);
and U23409 (N_23409,N_23213,N_23288);
and U23410 (N_23410,N_23279,N_23332);
nand U23411 (N_23411,N_23327,N_23243);
or U23412 (N_23412,N_23337,N_23253);
nand U23413 (N_23413,N_23298,N_23314);
nor U23414 (N_23414,N_23203,N_23336);
or U23415 (N_23415,N_23238,N_23260);
nand U23416 (N_23416,N_23261,N_23284);
nand U23417 (N_23417,N_23385,N_23276);
xnor U23418 (N_23418,N_23383,N_23248);
nor U23419 (N_23419,N_23398,N_23271);
and U23420 (N_23420,N_23267,N_23228);
and U23421 (N_23421,N_23300,N_23244);
and U23422 (N_23422,N_23371,N_23222);
nor U23423 (N_23423,N_23226,N_23346);
nor U23424 (N_23424,N_23331,N_23325);
xnor U23425 (N_23425,N_23334,N_23349);
xor U23426 (N_23426,N_23264,N_23361);
and U23427 (N_23427,N_23273,N_23240);
and U23428 (N_23428,N_23257,N_23233);
nand U23429 (N_23429,N_23286,N_23251);
xor U23430 (N_23430,N_23270,N_23230);
and U23431 (N_23431,N_23341,N_23387);
nor U23432 (N_23432,N_23234,N_23354);
or U23433 (N_23433,N_23378,N_23367);
nand U23434 (N_23434,N_23239,N_23392);
nor U23435 (N_23435,N_23201,N_23340);
or U23436 (N_23436,N_23218,N_23256);
nor U23437 (N_23437,N_23345,N_23301);
and U23438 (N_23438,N_23305,N_23379);
and U23439 (N_23439,N_23289,N_23229);
or U23440 (N_23440,N_23299,N_23370);
nor U23441 (N_23441,N_23389,N_23309);
xnor U23442 (N_23442,N_23362,N_23372);
or U23443 (N_23443,N_23212,N_23364);
nand U23444 (N_23444,N_23281,N_23200);
or U23445 (N_23445,N_23291,N_23250);
nand U23446 (N_23446,N_23311,N_23295);
and U23447 (N_23447,N_23399,N_23376);
or U23448 (N_23448,N_23318,N_23326);
nor U23449 (N_23449,N_23363,N_23394);
nand U23450 (N_23450,N_23263,N_23366);
or U23451 (N_23451,N_23358,N_23381);
and U23452 (N_23452,N_23210,N_23237);
nor U23453 (N_23453,N_23302,N_23227);
and U23454 (N_23454,N_23274,N_23333);
nor U23455 (N_23455,N_23391,N_23268);
and U23456 (N_23456,N_23204,N_23283);
nand U23457 (N_23457,N_23280,N_23277);
nand U23458 (N_23458,N_23252,N_23231);
xor U23459 (N_23459,N_23206,N_23216);
xor U23460 (N_23460,N_23307,N_23255);
nand U23461 (N_23461,N_23209,N_23330);
nand U23462 (N_23462,N_23397,N_23232);
and U23463 (N_23463,N_23339,N_23369);
or U23464 (N_23464,N_23324,N_23338);
nand U23465 (N_23465,N_23225,N_23208);
and U23466 (N_23466,N_23220,N_23348);
nand U23467 (N_23467,N_23246,N_23328);
and U23468 (N_23468,N_23329,N_23353);
or U23469 (N_23469,N_23303,N_23245);
and U23470 (N_23470,N_23320,N_23315);
nor U23471 (N_23471,N_23242,N_23377);
nor U23472 (N_23472,N_23236,N_23304);
xnor U23473 (N_23473,N_23296,N_23322);
nor U23474 (N_23474,N_23347,N_23247);
nor U23475 (N_23475,N_23382,N_23365);
xnor U23476 (N_23476,N_23224,N_23360);
and U23477 (N_23477,N_23214,N_23266);
nor U23478 (N_23478,N_23205,N_23386);
xnor U23479 (N_23479,N_23393,N_23316);
nand U23480 (N_23480,N_23265,N_23241);
nand U23481 (N_23481,N_23313,N_23321);
and U23482 (N_23482,N_23215,N_23308);
xnor U23483 (N_23483,N_23290,N_23373);
or U23484 (N_23484,N_23350,N_23221);
and U23485 (N_23485,N_23395,N_23352);
nand U23486 (N_23486,N_23275,N_23272);
and U23487 (N_23487,N_23355,N_23207);
nand U23488 (N_23488,N_23294,N_23258);
nor U23489 (N_23489,N_23219,N_23292);
or U23490 (N_23490,N_23310,N_23293);
or U23491 (N_23491,N_23344,N_23249);
nand U23492 (N_23492,N_23384,N_23351);
xnor U23493 (N_23493,N_23217,N_23262);
nor U23494 (N_23494,N_23390,N_23202);
nor U23495 (N_23495,N_23359,N_23285);
nand U23496 (N_23496,N_23254,N_23374);
nand U23497 (N_23497,N_23357,N_23259);
xnor U23498 (N_23498,N_23323,N_23335);
nand U23499 (N_23499,N_23319,N_23388);
and U23500 (N_23500,N_23207,N_23323);
or U23501 (N_23501,N_23324,N_23211);
nor U23502 (N_23502,N_23301,N_23305);
or U23503 (N_23503,N_23250,N_23248);
nor U23504 (N_23504,N_23395,N_23376);
nor U23505 (N_23505,N_23290,N_23282);
nand U23506 (N_23506,N_23250,N_23293);
nor U23507 (N_23507,N_23206,N_23282);
nand U23508 (N_23508,N_23258,N_23321);
nand U23509 (N_23509,N_23230,N_23395);
and U23510 (N_23510,N_23221,N_23203);
and U23511 (N_23511,N_23206,N_23242);
xor U23512 (N_23512,N_23390,N_23225);
nand U23513 (N_23513,N_23398,N_23371);
xor U23514 (N_23514,N_23362,N_23398);
and U23515 (N_23515,N_23359,N_23220);
nor U23516 (N_23516,N_23286,N_23244);
and U23517 (N_23517,N_23227,N_23265);
nor U23518 (N_23518,N_23396,N_23362);
nand U23519 (N_23519,N_23355,N_23288);
or U23520 (N_23520,N_23212,N_23358);
nor U23521 (N_23521,N_23313,N_23373);
and U23522 (N_23522,N_23260,N_23243);
and U23523 (N_23523,N_23393,N_23305);
nor U23524 (N_23524,N_23276,N_23327);
or U23525 (N_23525,N_23257,N_23253);
nor U23526 (N_23526,N_23340,N_23280);
xnor U23527 (N_23527,N_23279,N_23226);
and U23528 (N_23528,N_23382,N_23363);
nor U23529 (N_23529,N_23249,N_23210);
xor U23530 (N_23530,N_23376,N_23341);
or U23531 (N_23531,N_23374,N_23319);
nand U23532 (N_23532,N_23202,N_23216);
or U23533 (N_23533,N_23244,N_23221);
or U23534 (N_23534,N_23236,N_23264);
nor U23535 (N_23535,N_23225,N_23312);
and U23536 (N_23536,N_23390,N_23228);
nor U23537 (N_23537,N_23390,N_23215);
nor U23538 (N_23538,N_23347,N_23354);
and U23539 (N_23539,N_23295,N_23220);
or U23540 (N_23540,N_23347,N_23238);
nand U23541 (N_23541,N_23248,N_23249);
or U23542 (N_23542,N_23302,N_23253);
xor U23543 (N_23543,N_23266,N_23287);
xor U23544 (N_23544,N_23305,N_23203);
and U23545 (N_23545,N_23359,N_23202);
nand U23546 (N_23546,N_23256,N_23306);
or U23547 (N_23547,N_23346,N_23309);
nor U23548 (N_23548,N_23335,N_23347);
nor U23549 (N_23549,N_23370,N_23382);
nand U23550 (N_23550,N_23315,N_23298);
nor U23551 (N_23551,N_23379,N_23252);
xnor U23552 (N_23552,N_23208,N_23327);
or U23553 (N_23553,N_23315,N_23274);
xnor U23554 (N_23554,N_23329,N_23215);
xnor U23555 (N_23555,N_23285,N_23386);
and U23556 (N_23556,N_23217,N_23304);
nand U23557 (N_23557,N_23349,N_23247);
or U23558 (N_23558,N_23305,N_23306);
and U23559 (N_23559,N_23327,N_23353);
nand U23560 (N_23560,N_23265,N_23300);
xnor U23561 (N_23561,N_23201,N_23249);
nor U23562 (N_23562,N_23214,N_23236);
nor U23563 (N_23563,N_23225,N_23265);
or U23564 (N_23564,N_23295,N_23286);
and U23565 (N_23565,N_23361,N_23273);
nor U23566 (N_23566,N_23332,N_23340);
or U23567 (N_23567,N_23296,N_23343);
nand U23568 (N_23568,N_23339,N_23212);
and U23569 (N_23569,N_23324,N_23365);
or U23570 (N_23570,N_23356,N_23235);
xnor U23571 (N_23571,N_23297,N_23254);
or U23572 (N_23572,N_23252,N_23313);
nor U23573 (N_23573,N_23292,N_23308);
nor U23574 (N_23574,N_23306,N_23340);
nor U23575 (N_23575,N_23399,N_23201);
nand U23576 (N_23576,N_23225,N_23263);
nor U23577 (N_23577,N_23360,N_23222);
nor U23578 (N_23578,N_23383,N_23286);
nor U23579 (N_23579,N_23332,N_23378);
and U23580 (N_23580,N_23201,N_23312);
xnor U23581 (N_23581,N_23242,N_23282);
nor U23582 (N_23582,N_23350,N_23208);
xor U23583 (N_23583,N_23331,N_23359);
nor U23584 (N_23584,N_23254,N_23220);
nor U23585 (N_23585,N_23335,N_23318);
xor U23586 (N_23586,N_23234,N_23215);
xor U23587 (N_23587,N_23357,N_23358);
or U23588 (N_23588,N_23365,N_23393);
and U23589 (N_23589,N_23328,N_23254);
nand U23590 (N_23590,N_23232,N_23257);
or U23591 (N_23591,N_23326,N_23336);
nand U23592 (N_23592,N_23351,N_23331);
and U23593 (N_23593,N_23288,N_23214);
xor U23594 (N_23594,N_23328,N_23200);
and U23595 (N_23595,N_23356,N_23202);
nand U23596 (N_23596,N_23300,N_23225);
nand U23597 (N_23597,N_23276,N_23346);
nand U23598 (N_23598,N_23201,N_23325);
nand U23599 (N_23599,N_23223,N_23359);
xnor U23600 (N_23600,N_23402,N_23477);
and U23601 (N_23601,N_23418,N_23485);
xnor U23602 (N_23602,N_23447,N_23554);
xnor U23603 (N_23603,N_23422,N_23490);
nand U23604 (N_23604,N_23453,N_23449);
and U23605 (N_23605,N_23511,N_23563);
or U23606 (N_23606,N_23591,N_23462);
nand U23607 (N_23607,N_23437,N_23537);
and U23608 (N_23608,N_23484,N_23542);
nor U23609 (N_23609,N_23510,N_23444);
xor U23610 (N_23610,N_23565,N_23558);
or U23611 (N_23611,N_23552,N_23503);
xnor U23612 (N_23612,N_23434,N_23566);
nand U23613 (N_23613,N_23506,N_23545);
or U23614 (N_23614,N_23487,N_23592);
nor U23615 (N_23615,N_23499,N_23569);
nor U23616 (N_23616,N_23457,N_23573);
nand U23617 (N_23617,N_23517,N_23536);
and U23618 (N_23618,N_23436,N_23471);
nor U23619 (N_23619,N_23439,N_23411);
and U23620 (N_23620,N_23570,N_23519);
nand U23621 (N_23621,N_23562,N_23526);
xor U23622 (N_23622,N_23438,N_23578);
xor U23623 (N_23623,N_23448,N_23488);
nand U23624 (N_23624,N_23498,N_23473);
nor U23625 (N_23625,N_23424,N_23483);
nand U23626 (N_23626,N_23482,N_23456);
xor U23627 (N_23627,N_23446,N_23597);
or U23628 (N_23628,N_23400,N_23515);
nor U23629 (N_23629,N_23486,N_23599);
nor U23630 (N_23630,N_23523,N_23472);
and U23631 (N_23631,N_23412,N_23533);
and U23632 (N_23632,N_23481,N_23460);
or U23633 (N_23633,N_23403,N_23427);
and U23634 (N_23634,N_23568,N_23549);
or U23635 (N_23635,N_23464,N_23546);
nor U23636 (N_23636,N_23580,N_23497);
and U23637 (N_23637,N_23532,N_23587);
nand U23638 (N_23638,N_23458,N_23491);
nor U23639 (N_23639,N_23494,N_23540);
or U23640 (N_23640,N_23445,N_23431);
nand U23641 (N_23641,N_23596,N_23544);
nand U23642 (N_23642,N_23455,N_23441);
nor U23643 (N_23643,N_23572,N_23430);
nand U23644 (N_23644,N_23474,N_23551);
or U23645 (N_23645,N_23534,N_23454);
nor U23646 (N_23646,N_23550,N_23495);
nor U23647 (N_23647,N_23588,N_23579);
xnor U23648 (N_23648,N_23442,N_23443);
nand U23649 (N_23649,N_23440,N_23425);
nor U23650 (N_23650,N_23529,N_23571);
xor U23651 (N_23651,N_23469,N_23567);
or U23652 (N_23652,N_23527,N_23404);
or U23653 (N_23653,N_23593,N_23470);
nand U23654 (N_23654,N_23595,N_23507);
nand U23655 (N_23655,N_23475,N_23520);
xor U23656 (N_23656,N_23557,N_23508);
and U23657 (N_23657,N_23407,N_23419);
xor U23658 (N_23658,N_23426,N_23502);
nand U23659 (N_23659,N_23589,N_23463);
nand U23660 (N_23660,N_23416,N_23528);
and U23661 (N_23661,N_23465,N_23423);
or U23662 (N_23662,N_23435,N_23594);
nor U23663 (N_23663,N_23581,N_23535);
nor U23664 (N_23664,N_23512,N_23466);
or U23665 (N_23665,N_23459,N_23417);
nor U23666 (N_23666,N_23433,N_23553);
nand U23667 (N_23667,N_23509,N_23518);
or U23668 (N_23668,N_23561,N_23452);
nand U23669 (N_23669,N_23539,N_23413);
xnor U23670 (N_23670,N_23432,N_23501);
or U23671 (N_23671,N_23401,N_23555);
xor U23672 (N_23672,N_23489,N_23504);
or U23673 (N_23673,N_23450,N_23548);
xor U23674 (N_23674,N_23451,N_23409);
nand U23675 (N_23675,N_23428,N_23421);
and U23676 (N_23676,N_23556,N_23598);
and U23677 (N_23677,N_23467,N_23590);
and U23678 (N_23678,N_23586,N_23525);
nor U23679 (N_23679,N_23479,N_23584);
nand U23680 (N_23680,N_23524,N_23415);
nand U23681 (N_23681,N_23564,N_23530);
xnor U23682 (N_23682,N_23576,N_23585);
nand U23683 (N_23683,N_23575,N_23405);
nor U23684 (N_23684,N_23429,N_23478);
or U23685 (N_23685,N_23521,N_23547);
or U23686 (N_23686,N_23414,N_23505);
xnor U23687 (N_23687,N_23493,N_23468);
nor U23688 (N_23688,N_23461,N_23420);
and U23689 (N_23689,N_23577,N_23500);
or U23690 (N_23690,N_23406,N_23543);
and U23691 (N_23691,N_23560,N_23513);
and U23692 (N_23692,N_23559,N_23522);
xor U23693 (N_23693,N_23574,N_23582);
or U23694 (N_23694,N_23408,N_23496);
xor U23695 (N_23695,N_23410,N_23476);
nand U23696 (N_23696,N_23480,N_23514);
nor U23697 (N_23697,N_23492,N_23516);
and U23698 (N_23698,N_23538,N_23531);
xor U23699 (N_23699,N_23583,N_23541);
and U23700 (N_23700,N_23403,N_23540);
nor U23701 (N_23701,N_23433,N_23572);
and U23702 (N_23702,N_23543,N_23540);
nand U23703 (N_23703,N_23599,N_23461);
nor U23704 (N_23704,N_23516,N_23480);
or U23705 (N_23705,N_23522,N_23486);
and U23706 (N_23706,N_23482,N_23558);
and U23707 (N_23707,N_23474,N_23546);
and U23708 (N_23708,N_23524,N_23556);
nand U23709 (N_23709,N_23577,N_23505);
nand U23710 (N_23710,N_23555,N_23402);
xor U23711 (N_23711,N_23487,N_23572);
or U23712 (N_23712,N_23451,N_23489);
nor U23713 (N_23713,N_23589,N_23474);
or U23714 (N_23714,N_23589,N_23484);
and U23715 (N_23715,N_23485,N_23583);
xor U23716 (N_23716,N_23425,N_23556);
nor U23717 (N_23717,N_23482,N_23471);
nor U23718 (N_23718,N_23423,N_23440);
xnor U23719 (N_23719,N_23525,N_23499);
and U23720 (N_23720,N_23417,N_23513);
nor U23721 (N_23721,N_23511,N_23427);
nor U23722 (N_23722,N_23459,N_23561);
nand U23723 (N_23723,N_23562,N_23530);
or U23724 (N_23724,N_23543,N_23581);
and U23725 (N_23725,N_23595,N_23408);
nand U23726 (N_23726,N_23527,N_23583);
or U23727 (N_23727,N_23429,N_23427);
nand U23728 (N_23728,N_23473,N_23458);
xnor U23729 (N_23729,N_23516,N_23533);
nand U23730 (N_23730,N_23431,N_23497);
nor U23731 (N_23731,N_23460,N_23577);
and U23732 (N_23732,N_23541,N_23514);
or U23733 (N_23733,N_23570,N_23448);
or U23734 (N_23734,N_23445,N_23447);
nor U23735 (N_23735,N_23424,N_23409);
nand U23736 (N_23736,N_23536,N_23404);
xnor U23737 (N_23737,N_23487,N_23467);
nor U23738 (N_23738,N_23572,N_23452);
or U23739 (N_23739,N_23413,N_23453);
nor U23740 (N_23740,N_23410,N_23433);
xor U23741 (N_23741,N_23490,N_23479);
xor U23742 (N_23742,N_23575,N_23579);
nand U23743 (N_23743,N_23496,N_23551);
and U23744 (N_23744,N_23492,N_23420);
xnor U23745 (N_23745,N_23547,N_23573);
or U23746 (N_23746,N_23568,N_23547);
xnor U23747 (N_23747,N_23591,N_23434);
and U23748 (N_23748,N_23486,N_23560);
nand U23749 (N_23749,N_23408,N_23401);
nand U23750 (N_23750,N_23534,N_23430);
nand U23751 (N_23751,N_23436,N_23592);
xnor U23752 (N_23752,N_23469,N_23481);
and U23753 (N_23753,N_23498,N_23517);
nand U23754 (N_23754,N_23502,N_23596);
nor U23755 (N_23755,N_23567,N_23512);
nor U23756 (N_23756,N_23449,N_23519);
nand U23757 (N_23757,N_23465,N_23531);
or U23758 (N_23758,N_23463,N_23541);
or U23759 (N_23759,N_23460,N_23408);
nor U23760 (N_23760,N_23597,N_23554);
nand U23761 (N_23761,N_23451,N_23599);
and U23762 (N_23762,N_23537,N_23456);
xor U23763 (N_23763,N_23493,N_23583);
or U23764 (N_23764,N_23580,N_23479);
nor U23765 (N_23765,N_23568,N_23472);
and U23766 (N_23766,N_23454,N_23420);
nor U23767 (N_23767,N_23579,N_23563);
xor U23768 (N_23768,N_23561,N_23566);
or U23769 (N_23769,N_23435,N_23466);
and U23770 (N_23770,N_23534,N_23504);
xor U23771 (N_23771,N_23502,N_23579);
nor U23772 (N_23772,N_23447,N_23520);
or U23773 (N_23773,N_23536,N_23512);
nor U23774 (N_23774,N_23438,N_23538);
nand U23775 (N_23775,N_23406,N_23519);
or U23776 (N_23776,N_23587,N_23544);
nand U23777 (N_23777,N_23488,N_23558);
and U23778 (N_23778,N_23529,N_23553);
and U23779 (N_23779,N_23571,N_23580);
nor U23780 (N_23780,N_23429,N_23528);
nor U23781 (N_23781,N_23473,N_23502);
and U23782 (N_23782,N_23503,N_23589);
or U23783 (N_23783,N_23468,N_23530);
and U23784 (N_23784,N_23498,N_23446);
xor U23785 (N_23785,N_23466,N_23414);
or U23786 (N_23786,N_23431,N_23441);
nor U23787 (N_23787,N_23594,N_23585);
nand U23788 (N_23788,N_23435,N_23456);
nand U23789 (N_23789,N_23429,N_23596);
and U23790 (N_23790,N_23406,N_23594);
nand U23791 (N_23791,N_23581,N_23420);
or U23792 (N_23792,N_23550,N_23551);
nor U23793 (N_23793,N_23510,N_23569);
and U23794 (N_23794,N_23592,N_23556);
or U23795 (N_23795,N_23597,N_23559);
and U23796 (N_23796,N_23515,N_23414);
nor U23797 (N_23797,N_23436,N_23431);
nand U23798 (N_23798,N_23539,N_23581);
nand U23799 (N_23799,N_23442,N_23572);
and U23800 (N_23800,N_23783,N_23606);
nand U23801 (N_23801,N_23752,N_23779);
xor U23802 (N_23802,N_23726,N_23786);
xnor U23803 (N_23803,N_23664,N_23702);
and U23804 (N_23804,N_23703,N_23647);
xnor U23805 (N_23805,N_23709,N_23673);
xnor U23806 (N_23806,N_23616,N_23775);
nand U23807 (N_23807,N_23639,N_23623);
nor U23808 (N_23808,N_23684,N_23628);
or U23809 (N_23809,N_23655,N_23765);
nand U23810 (N_23810,N_23609,N_23778);
xnor U23811 (N_23811,N_23781,N_23652);
xnor U23812 (N_23812,N_23690,N_23794);
nor U23813 (N_23813,N_23671,N_23665);
xor U23814 (N_23814,N_23651,N_23791);
nor U23815 (N_23815,N_23677,N_23725);
or U23816 (N_23816,N_23611,N_23612);
nor U23817 (N_23817,N_23658,N_23679);
xor U23818 (N_23818,N_23715,N_23625);
nand U23819 (N_23819,N_23635,N_23678);
or U23820 (N_23820,N_23618,N_23650);
nor U23821 (N_23821,N_23713,N_23761);
nor U23822 (N_23822,N_23714,N_23742);
or U23823 (N_23823,N_23728,N_23766);
and U23824 (N_23824,N_23774,N_23797);
nand U23825 (N_23825,N_23600,N_23683);
xor U23826 (N_23826,N_23691,N_23785);
nand U23827 (N_23827,N_23780,N_23687);
nand U23828 (N_23828,N_23755,N_23634);
nor U23829 (N_23829,N_23748,N_23749);
and U23830 (N_23830,N_23719,N_23692);
nor U23831 (N_23831,N_23796,N_23740);
and U23832 (N_23832,N_23686,N_23694);
xor U23833 (N_23833,N_23729,N_23696);
and U23834 (N_23834,N_23646,N_23723);
xnor U23835 (N_23835,N_23769,N_23633);
or U23836 (N_23836,N_23770,N_23727);
and U23837 (N_23837,N_23631,N_23667);
or U23838 (N_23838,N_23680,N_23777);
nor U23839 (N_23839,N_23733,N_23627);
nor U23840 (N_23840,N_23784,N_23695);
or U23841 (N_23841,N_23669,N_23782);
nor U23842 (N_23842,N_23649,N_23632);
or U23843 (N_23843,N_23614,N_23798);
nor U23844 (N_23844,N_23660,N_23689);
and U23845 (N_23845,N_23648,N_23710);
or U23846 (N_23846,N_23699,N_23734);
and U23847 (N_23847,N_23672,N_23663);
and U23848 (N_23848,N_23736,N_23708);
xnor U23849 (N_23849,N_23707,N_23753);
nand U23850 (N_23850,N_23762,N_23763);
or U23851 (N_23851,N_23744,N_23739);
nand U23852 (N_23852,N_23746,N_23773);
and U23853 (N_23853,N_23682,N_23705);
nor U23854 (N_23854,N_23629,N_23654);
nor U23855 (N_23855,N_23668,N_23772);
or U23856 (N_23856,N_23756,N_23608);
nand U23857 (N_23857,N_23704,N_23701);
xor U23858 (N_23858,N_23792,N_23789);
xor U23859 (N_23859,N_23767,N_23768);
nor U23860 (N_23860,N_23624,N_23693);
and U23861 (N_23861,N_23697,N_23617);
nand U23862 (N_23862,N_23661,N_23716);
nand U23863 (N_23863,N_23670,N_23735);
nand U23864 (N_23864,N_23720,N_23657);
and U23865 (N_23865,N_23771,N_23745);
nand U23866 (N_23866,N_23681,N_23741);
or U23867 (N_23867,N_23604,N_23737);
xnor U23868 (N_23868,N_23607,N_23666);
nand U23869 (N_23869,N_23717,N_23675);
nor U23870 (N_23870,N_23622,N_23738);
nand U23871 (N_23871,N_23640,N_23637);
and U23872 (N_23872,N_23712,N_23601);
or U23873 (N_23873,N_23711,N_23662);
xor U23874 (N_23874,N_23721,N_23630);
or U23875 (N_23875,N_23638,N_23731);
and U23876 (N_23876,N_23641,N_23643);
xor U23877 (N_23877,N_23760,N_23764);
nor U23878 (N_23878,N_23653,N_23730);
nor U23879 (N_23879,N_23636,N_23602);
and U23880 (N_23880,N_23732,N_23795);
xor U23881 (N_23881,N_23757,N_23700);
nor U23882 (N_23882,N_23706,N_23620);
nor U23883 (N_23883,N_23610,N_23698);
xor U23884 (N_23884,N_23776,N_23747);
and U23885 (N_23885,N_23645,N_23724);
nor U23886 (N_23886,N_23743,N_23799);
nor U23887 (N_23887,N_23659,N_23619);
or U23888 (N_23888,N_23758,N_23793);
or U23889 (N_23889,N_23603,N_23751);
or U23890 (N_23890,N_23674,N_23750);
nor U23891 (N_23891,N_23787,N_23718);
nand U23892 (N_23892,N_23759,N_23621);
or U23893 (N_23893,N_23644,N_23754);
or U23894 (N_23894,N_23722,N_23615);
or U23895 (N_23895,N_23685,N_23790);
xor U23896 (N_23896,N_23642,N_23688);
xnor U23897 (N_23897,N_23788,N_23626);
xnor U23898 (N_23898,N_23605,N_23613);
or U23899 (N_23899,N_23656,N_23676);
nand U23900 (N_23900,N_23748,N_23633);
xor U23901 (N_23901,N_23681,N_23675);
nor U23902 (N_23902,N_23675,N_23769);
and U23903 (N_23903,N_23679,N_23713);
nand U23904 (N_23904,N_23681,N_23690);
or U23905 (N_23905,N_23600,N_23623);
nor U23906 (N_23906,N_23662,N_23721);
and U23907 (N_23907,N_23733,N_23643);
xor U23908 (N_23908,N_23674,N_23788);
nand U23909 (N_23909,N_23798,N_23675);
xnor U23910 (N_23910,N_23603,N_23600);
and U23911 (N_23911,N_23753,N_23754);
nand U23912 (N_23912,N_23757,N_23617);
or U23913 (N_23913,N_23686,N_23658);
nor U23914 (N_23914,N_23625,N_23657);
nor U23915 (N_23915,N_23725,N_23631);
nand U23916 (N_23916,N_23770,N_23613);
xnor U23917 (N_23917,N_23762,N_23632);
nor U23918 (N_23918,N_23667,N_23726);
xnor U23919 (N_23919,N_23697,N_23616);
nor U23920 (N_23920,N_23605,N_23731);
nor U23921 (N_23921,N_23774,N_23761);
nor U23922 (N_23922,N_23658,N_23639);
nand U23923 (N_23923,N_23662,N_23670);
nor U23924 (N_23924,N_23624,N_23696);
or U23925 (N_23925,N_23686,N_23689);
xnor U23926 (N_23926,N_23759,N_23662);
or U23927 (N_23927,N_23764,N_23783);
and U23928 (N_23928,N_23620,N_23603);
nand U23929 (N_23929,N_23735,N_23716);
or U23930 (N_23930,N_23657,N_23783);
and U23931 (N_23931,N_23759,N_23625);
or U23932 (N_23932,N_23727,N_23762);
nor U23933 (N_23933,N_23794,N_23684);
or U23934 (N_23934,N_23739,N_23651);
nand U23935 (N_23935,N_23704,N_23653);
nand U23936 (N_23936,N_23649,N_23694);
nor U23937 (N_23937,N_23661,N_23637);
or U23938 (N_23938,N_23664,N_23760);
or U23939 (N_23939,N_23694,N_23761);
or U23940 (N_23940,N_23736,N_23697);
xor U23941 (N_23941,N_23669,N_23640);
nand U23942 (N_23942,N_23616,N_23700);
nand U23943 (N_23943,N_23661,N_23640);
and U23944 (N_23944,N_23688,N_23701);
and U23945 (N_23945,N_23750,N_23655);
or U23946 (N_23946,N_23702,N_23633);
nor U23947 (N_23947,N_23644,N_23752);
and U23948 (N_23948,N_23759,N_23688);
xnor U23949 (N_23949,N_23694,N_23712);
nor U23950 (N_23950,N_23728,N_23659);
nor U23951 (N_23951,N_23637,N_23693);
and U23952 (N_23952,N_23635,N_23661);
xor U23953 (N_23953,N_23630,N_23613);
or U23954 (N_23954,N_23697,N_23609);
and U23955 (N_23955,N_23773,N_23713);
nand U23956 (N_23956,N_23631,N_23604);
nand U23957 (N_23957,N_23732,N_23780);
or U23958 (N_23958,N_23733,N_23794);
and U23959 (N_23959,N_23780,N_23631);
or U23960 (N_23960,N_23712,N_23774);
xor U23961 (N_23961,N_23616,N_23785);
or U23962 (N_23962,N_23690,N_23626);
or U23963 (N_23963,N_23762,N_23761);
nor U23964 (N_23964,N_23727,N_23732);
xor U23965 (N_23965,N_23746,N_23720);
and U23966 (N_23966,N_23720,N_23620);
or U23967 (N_23967,N_23711,N_23758);
nor U23968 (N_23968,N_23685,N_23626);
nor U23969 (N_23969,N_23674,N_23799);
or U23970 (N_23970,N_23612,N_23771);
nand U23971 (N_23971,N_23625,N_23794);
and U23972 (N_23972,N_23704,N_23767);
xor U23973 (N_23973,N_23626,N_23784);
nor U23974 (N_23974,N_23666,N_23761);
and U23975 (N_23975,N_23735,N_23624);
and U23976 (N_23976,N_23694,N_23753);
xor U23977 (N_23977,N_23605,N_23672);
nand U23978 (N_23978,N_23697,N_23767);
xor U23979 (N_23979,N_23692,N_23696);
nand U23980 (N_23980,N_23738,N_23749);
xor U23981 (N_23981,N_23729,N_23649);
or U23982 (N_23982,N_23615,N_23778);
nor U23983 (N_23983,N_23685,N_23614);
xnor U23984 (N_23984,N_23771,N_23707);
and U23985 (N_23985,N_23710,N_23714);
xnor U23986 (N_23986,N_23720,N_23747);
nor U23987 (N_23987,N_23682,N_23620);
and U23988 (N_23988,N_23630,N_23722);
nor U23989 (N_23989,N_23701,N_23672);
nand U23990 (N_23990,N_23669,N_23732);
nor U23991 (N_23991,N_23710,N_23687);
nand U23992 (N_23992,N_23612,N_23623);
nand U23993 (N_23993,N_23641,N_23762);
and U23994 (N_23994,N_23799,N_23645);
xor U23995 (N_23995,N_23676,N_23744);
and U23996 (N_23996,N_23701,N_23629);
nor U23997 (N_23997,N_23788,N_23613);
or U23998 (N_23998,N_23634,N_23745);
and U23999 (N_23999,N_23742,N_23724);
xor U24000 (N_24000,N_23970,N_23963);
and U24001 (N_24001,N_23918,N_23803);
or U24002 (N_24002,N_23875,N_23956);
xor U24003 (N_24003,N_23929,N_23884);
nor U24004 (N_24004,N_23838,N_23914);
nor U24005 (N_24005,N_23943,N_23821);
nand U24006 (N_24006,N_23874,N_23895);
and U24007 (N_24007,N_23991,N_23890);
or U24008 (N_24008,N_23863,N_23945);
nand U24009 (N_24009,N_23962,N_23902);
nand U24010 (N_24010,N_23815,N_23912);
and U24011 (N_24011,N_23953,N_23961);
or U24012 (N_24012,N_23930,N_23971);
nand U24013 (N_24013,N_23968,N_23995);
xor U24014 (N_24014,N_23949,N_23833);
nand U24015 (N_24015,N_23985,N_23829);
and U24016 (N_24016,N_23831,N_23851);
and U24017 (N_24017,N_23915,N_23801);
xnor U24018 (N_24018,N_23871,N_23869);
xor U24019 (N_24019,N_23976,N_23954);
xor U24020 (N_24020,N_23834,N_23897);
nand U24021 (N_24021,N_23901,N_23951);
nor U24022 (N_24022,N_23823,N_23909);
or U24023 (N_24023,N_23920,N_23841);
nand U24024 (N_24024,N_23883,N_23986);
and U24025 (N_24025,N_23804,N_23880);
or U24026 (N_24026,N_23973,N_23950);
xor U24027 (N_24027,N_23820,N_23982);
nor U24028 (N_24028,N_23933,N_23817);
nand U24029 (N_24029,N_23844,N_23958);
and U24030 (N_24030,N_23928,N_23827);
nor U24031 (N_24031,N_23892,N_23845);
nor U24032 (N_24032,N_23936,N_23842);
or U24033 (N_24033,N_23819,N_23975);
and U24034 (N_24034,N_23980,N_23835);
nor U24035 (N_24035,N_23927,N_23964);
nor U24036 (N_24036,N_23843,N_23868);
or U24037 (N_24037,N_23857,N_23886);
xor U24038 (N_24038,N_23940,N_23810);
xnor U24039 (N_24039,N_23917,N_23919);
and U24040 (N_24040,N_23987,N_23881);
and U24041 (N_24041,N_23898,N_23896);
and U24042 (N_24042,N_23922,N_23889);
and U24043 (N_24043,N_23867,N_23997);
and U24044 (N_24044,N_23865,N_23807);
or U24045 (N_24045,N_23992,N_23887);
or U24046 (N_24046,N_23984,N_23802);
nand U24047 (N_24047,N_23910,N_23818);
and U24048 (N_24048,N_23941,N_23861);
xor U24049 (N_24049,N_23937,N_23826);
or U24050 (N_24050,N_23935,N_23952);
nor U24051 (N_24051,N_23931,N_23977);
or U24052 (N_24052,N_23988,N_23888);
and U24053 (N_24053,N_23830,N_23806);
nor U24054 (N_24054,N_23858,N_23907);
xnor U24055 (N_24055,N_23876,N_23814);
and U24056 (N_24056,N_23942,N_23972);
xor U24057 (N_24057,N_23855,N_23948);
nand U24058 (N_24058,N_23966,N_23938);
or U24059 (N_24059,N_23854,N_23866);
and U24060 (N_24060,N_23900,N_23990);
nor U24061 (N_24061,N_23878,N_23944);
or U24062 (N_24062,N_23836,N_23947);
nor U24063 (N_24063,N_23899,N_23864);
and U24064 (N_24064,N_23960,N_23811);
nor U24065 (N_24065,N_23906,N_23939);
nand U24066 (N_24066,N_23911,N_23913);
nor U24067 (N_24067,N_23860,N_23916);
and U24068 (N_24068,N_23994,N_23983);
or U24069 (N_24069,N_23840,N_23856);
nand U24070 (N_24070,N_23999,N_23849);
nor U24071 (N_24071,N_23959,N_23925);
or U24072 (N_24072,N_23904,N_23816);
or U24073 (N_24073,N_23923,N_23839);
xnor U24074 (N_24074,N_23921,N_23946);
xnor U24075 (N_24075,N_23846,N_23837);
nand U24076 (N_24076,N_23893,N_23993);
xnor U24077 (N_24077,N_23872,N_23885);
nor U24078 (N_24078,N_23974,N_23873);
and U24079 (N_24079,N_23828,N_23998);
or U24080 (N_24080,N_23808,N_23850);
nor U24081 (N_24081,N_23969,N_23877);
xor U24082 (N_24082,N_23813,N_23894);
nor U24083 (N_24083,N_23848,N_23908);
nor U24084 (N_24084,N_23979,N_23852);
nand U24085 (N_24085,N_23809,N_23926);
and U24086 (N_24086,N_23989,N_23822);
and U24087 (N_24087,N_23832,N_23800);
or U24088 (N_24088,N_23957,N_23824);
nor U24089 (N_24089,N_23805,N_23812);
nor U24090 (N_24090,N_23825,N_23879);
xor U24091 (N_24091,N_23905,N_23859);
nor U24092 (N_24092,N_23924,N_23862);
nor U24093 (N_24093,N_23955,N_23932);
or U24094 (N_24094,N_23903,N_23891);
nor U24095 (N_24095,N_23978,N_23965);
and U24096 (N_24096,N_23967,N_23996);
nor U24097 (N_24097,N_23853,N_23934);
nor U24098 (N_24098,N_23870,N_23981);
nand U24099 (N_24099,N_23882,N_23847);
xor U24100 (N_24100,N_23892,N_23907);
or U24101 (N_24101,N_23847,N_23928);
or U24102 (N_24102,N_23890,N_23811);
nand U24103 (N_24103,N_23890,N_23937);
or U24104 (N_24104,N_23961,N_23918);
or U24105 (N_24105,N_23837,N_23981);
nor U24106 (N_24106,N_23956,N_23864);
and U24107 (N_24107,N_23938,N_23888);
and U24108 (N_24108,N_23924,N_23881);
xor U24109 (N_24109,N_23814,N_23952);
and U24110 (N_24110,N_23863,N_23927);
nand U24111 (N_24111,N_23919,N_23866);
nor U24112 (N_24112,N_23873,N_23920);
and U24113 (N_24113,N_23945,N_23806);
nand U24114 (N_24114,N_23824,N_23875);
xnor U24115 (N_24115,N_23830,N_23837);
xnor U24116 (N_24116,N_23851,N_23857);
nand U24117 (N_24117,N_23931,N_23984);
or U24118 (N_24118,N_23802,N_23889);
nand U24119 (N_24119,N_23825,N_23851);
and U24120 (N_24120,N_23969,N_23880);
xnor U24121 (N_24121,N_23850,N_23895);
and U24122 (N_24122,N_23943,N_23947);
nor U24123 (N_24123,N_23969,N_23934);
nand U24124 (N_24124,N_23812,N_23874);
and U24125 (N_24125,N_23856,N_23973);
nor U24126 (N_24126,N_23942,N_23920);
nor U24127 (N_24127,N_23925,N_23834);
xnor U24128 (N_24128,N_23921,N_23839);
xnor U24129 (N_24129,N_23895,N_23919);
and U24130 (N_24130,N_23901,N_23987);
xor U24131 (N_24131,N_23975,N_23893);
and U24132 (N_24132,N_23932,N_23824);
nor U24133 (N_24133,N_23910,N_23930);
nor U24134 (N_24134,N_23887,N_23892);
or U24135 (N_24135,N_23872,N_23863);
xnor U24136 (N_24136,N_23921,N_23822);
xor U24137 (N_24137,N_23931,N_23918);
nor U24138 (N_24138,N_23940,N_23876);
nand U24139 (N_24139,N_23810,N_23833);
and U24140 (N_24140,N_23960,N_23961);
xor U24141 (N_24141,N_23802,N_23832);
nor U24142 (N_24142,N_23901,N_23869);
xor U24143 (N_24143,N_23893,N_23921);
nand U24144 (N_24144,N_23881,N_23807);
nand U24145 (N_24145,N_23807,N_23986);
or U24146 (N_24146,N_23921,N_23938);
nor U24147 (N_24147,N_23826,N_23954);
nor U24148 (N_24148,N_23800,N_23902);
and U24149 (N_24149,N_23948,N_23839);
and U24150 (N_24150,N_23980,N_23996);
nand U24151 (N_24151,N_23904,N_23911);
or U24152 (N_24152,N_23956,N_23980);
or U24153 (N_24153,N_23966,N_23916);
xnor U24154 (N_24154,N_23870,N_23935);
nor U24155 (N_24155,N_23895,N_23816);
nand U24156 (N_24156,N_23886,N_23811);
or U24157 (N_24157,N_23911,N_23870);
nor U24158 (N_24158,N_23884,N_23896);
xnor U24159 (N_24159,N_23914,N_23901);
xnor U24160 (N_24160,N_23962,N_23805);
xor U24161 (N_24161,N_23981,N_23908);
xor U24162 (N_24162,N_23814,N_23998);
nand U24163 (N_24163,N_23898,N_23876);
and U24164 (N_24164,N_23931,N_23824);
nor U24165 (N_24165,N_23951,N_23855);
xor U24166 (N_24166,N_23969,N_23993);
xor U24167 (N_24167,N_23950,N_23849);
xor U24168 (N_24168,N_23837,N_23861);
and U24169 (N_24169,N_23897,N_23814);
xnor U24170 (N_24170,N_23879,N_23951);
nor U24171 (N_24171,N_23951,N_23838);
nand U24172 (N_24172,N_23877,N_23836);
xnor U24173 (N_24173,N_23936,N_23923);
and U24174 (N_24174,N_23942,N_23869);
and U24175 (N_24175,N_23887,N_23837);
and U24176 (N_24176,N_23987,N_23979);
xnor U24177 (N_24177,N_23819,N_23888);
xor U24178 (N_24178,N_23808,N_23894);
and U24179 (N_24179,N_23870,N_23855);
and U24180 (N_24180,N_23976,N_23994);
xor U24181 (N_24181,N_23811,N_23807);
and U24182 (N_24182,N_23873,N_23942);
nor U24183 (N_24183,N_23910,N_23996);
nor U24184 (N_24184,N_23879,N_23850);
xor U24185 (N_24185,N_23808,N_23972);
nor U24186 (N_24186,N_23855,N_23974);
nor U24187 (N_24187,N_23855,N_23979);
nand U24188 (N_24188,N_23801,N_23907);
and U24189 (N_24189,N_23852,N_23854);
or U24190 (N_24190,N_23986,N_23922);
and U24191 (N_24191,N_23971,N_23909);
and U24192 (N_24192,N_23877,N_23951);
and U24193 (N_24193,N_23943,N_23977);
nand U24194 (N_24194,N_23951,N_23824);
nor U24195 (N_24195,N_23843,N_23971);
nor U24196 (N_24196,N_23826,N_23939);
nor U24197 (N_24197,N_23950,N_23997);
nor U24198 (N_24198,N_23973,N_23868);
or U24199 (N_24199,N_23968,N_23831);
xnor U24200 (N_24200,N_24195,N_24142);
and U24201 (N_24201,N_24113,N_24043);
xnor U24202 (N_24202,N_24114,N_24032);
xnor U24203 (N_24203,N_24129,N_24019);
and U24204 (N_24204,N_24126,N_24028);
and U24205 (N_24205,N_24150,N_24029);
xnor U24206 (N_24206,N_24115,N_24141);
xnor U24207 (N_24207,N_24057,N_24151);
or U24208 (N_24208,N_24054,N_24030);
or U24209 (N_24209,N_24153,N_24134);
nor U24210 (N_24210,N_24133,N_24066);
nor U24211 (N_24211,N_24042,N_24087);
xor U24212 (N_24212,N_24177,N_24060);
nor U24213 (N_24213,N_24199,N_24014);
nand U24214 (N_24214,N_24034,N_24040);
xnor U24215 (N_24215,N_24073,N_24025);
nand U24216 (N_24216,N_24069,N_24007);
and U24217 (N_24217,N_24003,N_24031);
nor U24218 (N_24218,N_24139,N_24172);
and U24219 (N_24219,N_24051,N_24100);
xnor U24220 (N_24220,N_24059,N_24197);
or U24221 (N_24221,N_24154,N_24187);
or U24222 (N_24222,N_24170,N_24103);
and U24223 (N_24223,N_24157,N_24053);
xnor U24224 (N_24224,N_24167,N_24198);
nor U24225 (N_24225,N_24109,N_24077);
nor U24226 (N_24226,N_24145,N_24144);
nor U24227 (N_24227,N_24106,N_24118);
nand U24228 (N_24228,N_24178,N_24192);
nand U24229 (N_24229,N_24135,N_24191);
xnor U24230 (N_24230,N_24127,N_24140);
nand U24231 (N_24231,N_24183,N_24188);
nand U24232 (N_24232,N_24093,N_24189);
and U24233 (N_24233,N_24194,N_24062);
nand U24234 (N_24234,N_24041,N_24011);
nand U24235 (N_24235,N_24095,N_24065);
nand U24236 (N_24236,N_24076,N_24009);
nor U24237 (N_24237,N_24048,N_24174);
nand U24238 (N_24238,N_24067,N_24044);
and U24239 (N_24239,N_24016,N_24180);
xor U24240 (N_24240,N_24146,N_24184);
or U24241 (N_24241,N_24185,N_24173);
nand U24242 (N_24242,N_24006,N_24190);
nor U24243 (N_24243,N_24101,N_24027);
and U24244 (N_24244,N_24038,N_24084);
or U24245 (N_24245,N_24010,N_24008);
xnor U24246 (N_24246,N_24026,N_24130);
nand U24247 (N_24247,N_24110,N_24022);
xor U24248 (N_24248,N_24089,N_24148);
and U24249 (N_24249,N_24020,N_24002);
nand U24250 (N_24250,N_24164,N_24107);
or U24251 (N_24251,N_24165,N_24169);
and U24252 (N_24252,N_24179,N_24005);
nor U24253 (N_24253,N_24155,N_24074);
nand U24254 (N_24254,N_24098,N_24166);
nand U24255 (N_24255,N_24125,N_24162);
nor U24256 (N_24256,N_24132,N_24099);
xnor U24257 (N_24257,N_24102,N_24147);
or U24258 (N_24258,N_24108,N_24097);
xor U24259 (N_24259,N_24049,N_24119);
or U24260 (N_24260,N_24045,N_24021);
or U24261 (N_24261,N_24122,N_24096);
nor U24262 (N_24262,N_24120,N_24082);
or U24263 (N_24263,N_24012,N_24112);
or U24264 (N_24264,N_24075,N_24160);
or U24265 (N_24265,N_24013,N_24128);
and U24266 (N_24266,N_24090,N_24071);
xor U24267 (N_24267,N_24033,N_24104);
xnor U24268 (N_24268,N_24046,N_24158);
nor U24269 (N_24269,N_24037,N_24092);
and U24270 (N_24270,N_24000,N_24036);
or U24271 (N_24271,N_24001,N_24161);
or U24272 (N_24272,N_24064,N_24117);
and U24273 (N_24273,N_24081,N_24105);
or U24274 (N_24274,N_24137,N_24079);
and U24275 (N_24275,N_24072,N_24080);
and U24276 (N_24276,N_24152,N_24156);
or U24277 (N_24277,N_24159,N_24078);
nand U24278 (N_24278,N_24091,N_24083);
xor U24279 (N_24279,N_24186,N_24193);
or U24280 (N_24280,N_24182,N_24047);
and U24281 (N_24281,N_24068,N_24136);
and U24282 (N_24282,N_24138,N_24023);
or U24283 (N_24283,N_24124,N_24168);
nor U24284 (N_24284,N_24052,N_24111);
and U24285 (N_24285,N_24176,N_24058);
or U24286 (N_24286,N_24131,N_24039);
and U24287 (N_24287,N_24063,N_24018);
nand U24288 (N_24288,N_24181,N_24175);
xnor U24289 (N_24289,N_24086,N_24085);
and U24290 (N_24290,N_24171,N_24055);
nor U24291 (N_24291,N_24035,N_24024);
nor U24292 (N_24292,N_24149,N_24050);
nand U24293 (N_24293,N_24094,N_24163);
or U24294 (N_24294,N_24015,N_24123);
nor U24295 (N_24295,N_24056,N_24196);
xor U24296 (N_24296,N_24088,N_24061);
xnor U24297 (N_24297,N_24121,N_24004);
nor U24298 (N_24298,N_24143,N_24017);
nand U24299 (N_24299,N_24116,N_24070);
nand U24300 (N_24300,N_24073,N_24168);
or U24301 (N_24301,N_24069,N_24045);
and U24302 (N_24302,N_24192,N_24027);
xnor U24303 (N_24303,N_24052,N_24099);
or U24304 (N_24304,N_24166,N_24022);
xnor U24305 (N_24305,N_24100,N_24140);
or U24306 (N_24306,N_24144,N_24010);
nor U24307 (N_24307,N_24040,N_24091);
nand U24308 (N_24308,N_24172,N_24029);
nand U24309 (N_24309,N_24153,N_24146);
and U24310 (N_24310,N_24067,N_24173);
and U24311 (N_24311,N_24166,N_24081);
xor U24312 (N_24312,N_24141,N_24081);
and U24313 (N_24313,N_24067,N_24007);
xor U24314 (N_24314,N_24101,N_24178);
xor U24315 (N_24315,N_24108,N_24118);
nand U24316 (N_24316,N_24188,N_24150);
nand U24317 (N_24317,N_24154,N_24174);
or U24318 (N_24318,N_24193,N_24156);
nor U24319 (N_24319,N_24109,N_24118);
nor U24320 (N_24320,N_24165,N_24112);
or U24321 (N_24321,N_24162,N_24174);
or U24322 (N_24322,N_24022,N_24156);
and U24323 (N_24323,N_24074,N_24075);
nor U24324 (N_24324,N_24024,N_24165);
nor U24325 (N_24325,N_24097,N_24113);
xor U24326 (N_24326,N_24087,N_24150);
xor U24327 (N_24327,N_24096,N_24059);
and U24328 (N_24328,N_24091,N_24141);
and U24329 (N_24329,N_24010,N_24064);
nand U24330 (N_24330,N_24016,N_24168);
nor U24331 (N_24331,N_24136,N_24160);
and U24332 (N_24332,N_24070,N_24041);
nor U24333 (N_24333,N_24128,N_24006);
nor U24334 (N_24334,N_24162,N_24175);
and U24335 (N_24335,N_24013,N_24171);
or U24336 (N_24336,N_24096,N_24027);
or U24337 (N_24337,N_24037,N_24135);
xnor U24338 (N_24338,N_24164,N_24017);
and U24339 (N_24339,N_24059,N_24039);
xnor U24340 (N_24340,N_24181,N_24031);
or U24341 (N_24341,N_24117,N_24137);
xor U24342 (N_24342,N_24144,N_24024);
or U24343 (N_24343,N_24159,N_24006);
nor U24344 (N_24344,N_24095,N_24004);
or U24345 (N_24345,N_24194,N_24060);
nor U24346 (N_24346,N_24010,N_24150);
and U24347 (N_24347,N_24052,N_24157);
nor U24348 (N_24348,N_24085,N_24128);
or U24349 (N_24349,N_24027,N_24195);
nand U24350 (N_24350,N_24025,N_24061);
xor U24351 (N_24351,N_24190,N_24141);
nand U24352 (N_24352,N_24073,N_24003);
and U24353 (N_24353,N_24077,N_24148);
or U24354 (N_24354,N_24164,N_24095);
and U24355 (N_24355,N_24100,N_24148);
and U24356 (N_24356,N_24022,N_24016);
nand U24357 (N_24357,N_24198,N_24045);
nor U24358 (N_24358,N_24180,N_24066);
or U24359 (N_24359,N_24105,N_24160);
and U24360 (N_24360,N_24018,N_24070);
nor U24361 (N_24361,N_24183,N_24029);
xor U24362 (N_24362,N_24023,N_24147);
and U24363 (N_24363,N_24018,N_24164);
nor U24364 (N_24364,N_24047,N_24008);
nand U24365 (N_24365,N_24076,N_24105);
nor U24366 (N_24366,N_24163,N_24148);
or U24367 (N_24367,N_24035,N_24158);
and U24368 (N_24368,N_24079,N_24100);
or U24369 (N_24369,N_24034,N_24131);
or U24370 (N_24370,N_24030,N_24011);
nand U24371 (N_24371,N_24165,N_24083);
xor U24372 (N_24372,N_24005,N_24174);
nor U24373 (N_24373,N_24071,N_24163);
nor U24374 (N_24374,N_24127,N_24102);
nand U24375 (N_24375,N_24170,N_24030);
nand U24376 (N_24376,N_24173,N_24169);
or U24377 (N_24377,N_24081,N_24069);
and U24378 (N_24378,N_24096,N_24161);
or U24379 (N_24379,N_24132,N_24100);
and U24380 (N_24380,N_24101,N_24185);
or U24381 (N_24381,N_24004,N_24013);
or U24382 (N_24382,N_24033,N_24188);
nor U24383 (N_24383,N_24078,N_24061);
nor U24384 (N_24384,N_24075,N_24072);
nand U24385 (N_24385,N_24129,N_24080);
nand U24386 (N_24386,N_24049,N_24008);
and U24387 (N_24387,N_24093,N_24026);
nor U24388 (N_24388,N_24131,N_24161);
nand U24389 (N_24389,N_24059,N_24167);
nor U24390 (N_24390,N_24056,N_24026);
nand U24391 (N_24391,N_24017,N_24193);
nand U24392 (N_24392,N_24110,N_24125);
nand U24393 (N_24393,N_24088,N_24017);
nand U24394 (N_24394,N_24171,N_24199);
nor U24395 (N_24395,N_24142,N_24162);
nand U24396 (N_24396,N_24170,N_24198);
xnor U24397 (N_24397,N_24079,N_24149);
nor U24398 (N_24398,N_24035,N_24123);
and U24399 (N_24399,N_24134,N_24058);
and U24400 (N_24400,N_24252,N_24355);
or U24401 (N_24401,N_24296,N_24345);
nor U24402 (N_24402,N_24305,N_24306);
xnor U24403 (N_24403,N_24336,N_24277);
and U24404 (N_24404,N_24325,N_24267);
nand U24405 (N_24405,N_24317,N_24213);
nor U24406 (N_24406,N_24241,N_24331);
xor U24407 (N_24407,N_24366,N_24367);
and U24408 (N_24408,N_24398,N_24399);
and U24409 (N_24409,N_24257,N_24223);
nand U24410 (N_24410,N_24339,N_24315);
and U24411 (N_24411,N_24395,N_24372);
and U24412 (N_24412,N_24392,N_24322);
and U24413 (N_24413,N_24236,N_24300);
xor U24414 (N_24414,N_24260,N_24338);
and U24415 (N_24415,N_24365,N_24280);
or U24416 (N_24416,N_24230,N_24253);
xnor U24417 (N_24417,N_24337,N_24308);
nand U24418 (N_24418,N_24389,N_24310);
nor U24419 (N_24419,N_24341,N_24218);
and U24420 (N_24420,N_24266,N_24272);
or U24421 (N_24421,N_24360,N_24297);
nor U24422 (N_24422,N_24309,N_24353);
and U24423 (N_24423,N_24209,N_24381);
and U24424 (N_24424,N_24323,N_24385);
nand U24425 (N_24425,N_24294,N_24374);
xor U24426 (N_24426,N_24231,N_24344);
nor U24427 (N_24427,N_24319,N_24240);
or U24428 (N_24428,N_24330,N_24214);
nor U24429 (N_24429,N_24248,N_24351);
nand U24430 (N_24430,N_24215,N_24256);
nor U24431 (N_24431,N_24270,N_24282);
and U24432 (N_24432,N_24269,N_24249);
xnor U24433 (N_24433,N_24333,N_24283);
nor U24434 (N_24434,N_24238,N_24329);
nor U24435 (N_24435,N_24335,N_24304);
nand U24436 (N_24436,N_24312,N_24364);
and U24437 (N_24437,N_24350,N_24288);
nor U24438 (N_24438,N_24358,N_24377);
xnor U24439 (N_24439,N_24378,N_24244);
or U24440 (N_24440,N_24320,N_24390);
or U24441 (N_24441,N_24397,N_24203);
or U24442 (N_24442,N_24217,N_24202);
xnor U24443 (N_24443,N_24207,N_24262);
or U24444 (N_24444,N_24212,N_24334);
nand U24445 (N_24445,N_24289,N_24234);
or U24446 (N_24446,N_24268,N_24384);
or U24447 (N_24447,N_24382,N_24255);
and U24448 (N_24448,N_24259,N_24293);
nor U24449 (N_24449,N_24233,N_24396);
or U24450 (N_24450,N_24328,N_24318);
nor U24451 (N_24451,N_24301,N_24298);
nor U24452 (N_24452,N_24387,N_24376);
xnor U24453 (N_24453,N_24229,N_24232);
xor U24454 (N_24454,N_24324,N_24278);
nand U24455 (N_24455,N_24311,N_24356);
and U24456 (N_24456,N_24352,N_24379);
xor U24457 (N_24457,N_24292,N_24205);
and U24458 (N_24458,N_24219,N_24204);
and U24459 (N_24459,N_24242,N_24380);
and U24460 (N_24460,N_24285,N_24250);
or U24461 (N_24461,N_24275,N_24220);
xor U24462 (N_24462,N_24287,N_24394);
or U24463 (N_24463,N_24246,N_24274);
xor U24464 (N_24464,N_24299,N_24375);
and U24465 (N_24465,N_24206,N_24201);
or U24466 (N_24466,N_24263,N_24222);
and U24467 (N_24467,N_24225,N_24290);
nor U24468 (N_24468,N_24370,N_24346);
nor U24469 (N_24469,N_24342,N_24261);
nand U24470 (N_24470,N_24314,N_24227);
or U24471 (N_24471,N_24295,N_24332);
xnor U24472 (N_24472,N_24326,N_24254);
and U24473 (N_24473,N_24369,N_24359);
nor U24474 (N_24474,N_24363,N_24362);
and U24475 (N_24475,N_24349,N_24237);
or U24476 (N_24476,N_24200,N_24216);
xor U24477 (N_24477,N_24313,N_24226);
and U24478 (N_24478,N_24373,N_24302);
nand U24479 (N_24479,N_24211,N_24273);
nand U24480 (N_24480,N_24235,N_24357);
and U24481 (N_24481,N_24271,N_24286);
and U24482 (N_24482,N_24347,N_24340);
nor U24483 (N_24483,N_24258,N_24265);
or U24484 (N_24484,N_24354,N_24327);
xor U24485 (N_24485,N_24388,N_24245);
xor U24486 (N_24486,N_24284,N_24321);
nor U24487 (N_24487,N_24210,N_24343);
xor U24488 (N_24488,N_24279,N_24316);
xor U24489 (N_24489,N_24243,N_24391);
and U24490 (N_24490,N_24224,N_24393);
xnor U24491 (N_24491,N_24208,N_24281);
nor U24492 (N_24492,N_24228,N_24239);
nor U24493 (N_24493,N_24368,N_24251);
or U24494 (N_24494,N_24386,N_24264);
and U24495 (N_24495,N_24291,N_24361);
and U24496 (N_24496,N_24247,N_24307);
or U24497 (N_24497,N_24221,N_24303);
nand U24498 (N_24498,N_24276,N_24348);
xnor U24499 (N_24499,N_24383,N_24371);
nand U24500 (N_24500,N_24397,N_24257);
nor U24501 (N_24501,N_24278,N_24224);
nor U24502 (N_24502,N_24319,N_24250);
nor U24503 (N_24503,N_24270,N_24243);
and U24504 (N_24504,N_24267,N_24313);
nand U24505 (N_24505,N_24255,N_24263);
and U24506 (N_24506,N_24362,N_24325);
nand U24507 (N_24507,N_24390,N_24235);
nand U24508 (N_24508,N_24348,N_24204);
nor U24509 (N_24509,N_24302,N_24354);
and U24510 (N_24510,N_24207,N_24293);
xor U24511 (N_24511,N_24271,N_24355);
and U24512 (N_24512,N_24283,N_24261);
nor U24513 (N_24513,N_24258,N_24261);
xor U24514 (N_24514,N_24396,N_24245);
and U24515 (N_24515,N_24382,N_24270);
xnor U24516 (N_24516,N_24333,N_24371);
or U24517 (N_24517,N_24264,N_24301);
nor U24518 (N_24518,N_24297,N_24237);
xnor U24519 (N_24519,N_24214,N_24259);
and U24520 (N_24520,N_24367,N_24213);
nand U24521 (N_24521,N_24303,N_24396);
nor U24522 (N_24522,N_24372,N_24298);
or U24523 (N_24523,N_24200,N_24242);
nand U24524 (N_24524,N_24390,N_24208);
xnor U24525 (N_24525,N_24288,N_24270);
nor U24526 (N_24526,N_24221,N_24332);
and U24527 (N_24527,N_24350,N_24247);
or U24528 (N_24528,N_24227,N_24353);
and U24529 (N_24529,N_24256,N_24347);
nand U24530 (N_24530,N_24311,N_24386);
nor U24531 (N_24531,N_24395,N_24247);
nand U24532 (N_24532,N_24374,N_24284);
nor U24533 (N_24533,N_24270,N_24373);
xnor U24534 (N_24534,N_24371,N_24380);
nand U24535 (N_24535,N_24270,N_24364);
and U24536 (N_24536,N_24221,N_24322);
xnor U24537 (N_24537,N_24299,N_24218);
xor U24538 (N_24538,N_24229,N_24322);
xor U24539 (N_24539,N_24207,N_24317);
and U24540 (N_24540,N_24369,N_24345);
nand U24541 (N_24541,N_24217,N_24282);
and U24542 (N_24542,N_24255,N_24347);
xor U24543 (N_24543,N_24387,N_24383);
or U24544 (N_24544,N_24307,N_24358);
nand U24545 (N_24545,N_24375,N_24244);
nor U24546 (N_24546,N_24343,N_24248);
xnor U24547 (N_24547,N_24371,N_24353);
and U24548 (N_24548,N_24210,N_24325);
xor U24549 (N_24549,N_24290,N_24257);
xnor U24550 (N_24550,N_24270,N_24381);
xor U24551 (N_24551,N_24267,N_24211);
or U24552 (N_24552,N_24279,N_24259);
or U24553 (N_24553,N_24214,N_24205);
or U24554 (N_24554,N_24353,N_24379);
nor U24555 (N_24555,N_24210,N_24345);
or U24556 (N_24556,N_24221,N_24230);
nor U24557 (N_24557,N_24357,N_24393);
xnor U24558 (N_24558,N_24393,N_24283);
or U24559 (N_24559,N_24265,N_24203);
and U24560 (N_24560,N_24394,N_24263);
nor U24561 (N_24561,N_24313,N_24388);
nand U24562 (N_24562,N_24219,N_24217);
nor U24563 (N_24563,N_24361,N_24282);
or U24564 (N_24564,N_24350,N_24333);
xor U24565 (N_24565,N_24325,N_24205);
nor U24566 (N_24566,N_24232,N_24373);
nand U24567 (N_24567,N_24395,N_24209);
or U24568 (N_24568,N_24227,N_24287);
nor U24569 (N_24569,N_24377,N_24391);
nor U24570 (N_24570,N_24201,N_24228);
nand U24571 (N_24571,N_24216,N_24301);
nor U24572 (N_24572,N_24211,N_24272);
and U24573 (N_24573,N_24339,N_24278);
or U24574 (N_24574,N_24336,N_24359);
xor U24575 (N_24575,N_24215,N_24326);
nor U24576 (N_24576,N_24368,N_24262);
nor U24577 (N_24577,N_24312,N_24241);
and U24578 (N_24578,N_24268,N_24307);
nor U24579 (N_24579,N_24393,N_24385);
or U24580 (N_24580,N_24386,N_24324);
and U24581 (N_24581,N_24298,N_24254);
nand U24582 (N_24582,N_24295,N_24225);
and U24583 (N_24583,N_24268,N_24283);
xnor U24584 (N_24584,N_24264,N_24256);
nand U24585 (N_24585,N_24311,N_24291);
and U24586 (N_24586,N_24250,N_24351);
or U24587 (N_24587,N_24280,N_24289);
or U24588 (N_24588,N_24217,N_24286);
or U24589 (N_24589,N_24221,N_24245);
xor U24590 (N_24590,N_24309,N_24340);
and U24591 (N_24591,N_24349,N_24245);
nor U24592 (N_24592,N_24305,N_24231);
and U24593 (N_24593,N_24259,N_24230);
nand U24594 (N_24594,N_24234,N_24374);
nor U24595 (N_24595,N_24219,N_24241);
and U24596 (N_24596,N_24297,N_24364);
nor U24597 (N_24597,N_24210,N_24302);
and U24598 (N_24598,N_24249,N_24370);
or U24599 (N_24599,N_24347,N_24337);
and U24600 (N_24600,N_24536,N_24497);
nand U24601 (N_24601,N_24479,N_24577);
and U24602 (N_24602,N_24509,N_24563);
and U24603 (N_24603,N_24470,N_24535);
nand U24604 (N_24604,N_24538,N_24430);
or U24605 (N_24605,N_24585,N_24566);
nand U24606 (N_24606,N_24544,N_24458);
nand U24607 (N_24607,N_24416,N_24593);
nor U24608 (N_24608,N_24418,N_24568);
xnor U24609 (N_24609,N_24446,N_24511);
and U24610 (N_24610,N_24594,N_24477);
nand U24611 (N_24611,N_24414,N_24423);
xnor U24612 (N_24612,N_24412,N_24533);
and U24613 (N_24613,N_24512,N_24441);
and U24614 (N_24614,N_24401,N_24518);
nor U24615 (N_24615,N_24539,N_24467);
xnor U24616 (N_24616,N_24495,N_24514);
nor U24617 (N_24617,N_24435,N_24491);
nand U24618 (N_24618,N_24567,N_24540);
and U24619 (N_24619,N_24506,N_24400);
nand U24620 (N_24620,N_24598,N_24550);
or U24621 (N_24621,N_24419,N_24437);
xor U24622 (N_24622,N_24422,N_24442);
or U24623 (N_24623,N_24478,N_24503);
nor U24624 (N_24624,N_24586,N_24500);
or U24625 (N_24625,N_24452,N_24426);
nand U24626 (N_24626,N_24561,N_24556);
or U24627 (N_24627,N_24529,N_24570);
xnor U24628 (N_24628,N_24582,N_24517);
nor U24629 (N_24629,N_24428,N_24432);
nand U24630 (N_24630,N_24413,N_24531);
nand U24631 (N_24631,N_24417,N_24499);
nor U24632 (N_24632,N_24486,N_24436);
nor U24633 (N_24633,N_24520,N_24579);
nor U24634 (N_24634,N_24508,N_24553);
xnor U24635 (N_24635,N_24543,N_24434);
xnor U24636 (N_24636,N_24421,N_24445);
or U24637 (N_24637,N_24547,N_24440);
xor U24638 (N_24638,N_24496,N_24504);
nand U24639 (N_24639,N_24410,N_24466);
nand U24640 (N_24640,N_24492,N_24560);
and U24641 (N_24641,N_24589,N_24494);
and U24642 (N_24642,N_24469,N_24498);
or U24643 (N_24643,N_24532,N_24415);
nor U24644 (N_24644,N_24562,N_24578);
xor U24645 (N_24645,N_24451,N_24405);
xnor U24646 (N_24646,N_24480,N_24475);
and U24647 (N_24647,N_24459,N_24580);
and U24648 (N_24648,N_24404,N_24559);
nor U24649 (N_24649,N_24493,N_24552);
nor U24650 (N_24650,N_24527,N_24461);
xor U24651 (N_24651,N_24403,N_24505);
or U24652 (N_24652,N_24574,N_24546);
or U24653 (N_24653,N_24502,N_24484);
nand U24654 (N_24654,N_24472,N_24464);
xor U24655 (N_24655,N_24474,N_24481);
xor U24656 (N_24656,N_24558,N_24462);
or U24657 (N_24657,N_24429,N_24427);
and U24658 (N_24658,N_24599,N_24490);
or U24659 (N_24659,N_24411,N_24473);
nor U24660 (N_24660,N_24551,N_24534);
or U24661 (N_24661,N_24488,N_24528);
nor U24662 (N_24662,N_24571,N_24530);
nor U24663 (N_24663,N_24408,N_24522);
nor U24664 (N_24664,N_24450,N_24460);
or U24665 (N_24665,N_24595,N_24483);
or U24666 (N_24666,N_24541,N_24448);
nor U24667 (N_24667,N_24485,N_24471);
and U24668 (N_24668,N_24468,N_24510);
xnor U24669 (N_24669,N_24545,N_24521);
or U24670 (N_24670,N_24564,N_24519);
or U24671 (N_24671,N_24537,N_24592);
nor U24672 (N_24672,N_24548,N_24569);
nor U24673 (N_24673,N_24542,N_24583);
and U24674 (N_24674,N_24439,N_24596);
and U24675 (N_24675,N_24489,N_24438);
nand U24676 (N_24676,N_24425,N_24409);
and U24677 (N_24677,N_24476,N_24406);
nor U24678 (N_24678,N_24407,N_24575);
xor U24679 (N_24679,N_24555,N_24424);
nand U24680 (N_24680,N_24576,N_24565);
nand U24681 (N_24681,N_24420,N_24525);
or U24682 (N_24682,N_24524,N_24588);
or U24683 (N_24683,N_24431,N_24573);
xnor U24684 (N_24684,N_24402,N_24557);
nor U24685 (N_24685,N_24591,N_24597);
or U24686 (N_24686,N_24549,N_24515);
or U24687 (N_24687,N_24482,N_24523);
or U24688 (N_24688,N_24454,N_24447);
xor U24689 (N_24689,N_24455,N_24449);
nand U24690 (N_24690,N_24457,N_24465);
nor U24691 (N_24691,N_24526,N_24456);
nor U24692 (N_24692,N_24587,N_24590);
nand U24693 (N_24693,N_24554,N_24487);
or U24694 (N_24694,N_24443,N_24507);
nor U24695 (N_24695,N_24516,N_24501);
xnor U24696 (N_24696,N_24584,N_24433);
and U24697 (N_24697,N_24463,N_24513);
nor U24698 (N_24698,N_24453,N_24581);
xor U24699 (N_24699,N_24444,N_24572);
nand U24700 (N_24700,N_24455,N_24521);
or U24701 (N_24701,N_24496,N_24532);
nor U24702 (N_24702,N_24522,N_24448);
nor U24703 (N_24703,N_24585,N_24543);
or U24704 (N_24704,N_24540,N_24440);
xnor U24705 (N_24705,N_24407,N_24586);
and U24706 (N_24706,N_24533,N_24490);
and U24707 (N_24707,N_24550,N_24507);
or U24708 (N_24708,N_24404,N_24567);
and U24709 (N_24709,N_24519,N_24579);
and U24710 (N_24710,N_24466,N_24487);
nand U24711 (N_24711,N_24499,N_24583);
nor U24712 (N_24712,N_24517,N_24536);
and U24713 (N_24713,N_24451,N_24553);
nor U24714 (N_24714,N_24531,N_24457);
nor U24715 (N_24715,N_24598,N_24483);
xor U24716 (N_24716,N_24568,N_24404);
nor U24717 (N_24717,N_24529,N_24557);
nor U24718 (N_24718,N_24593,N_24505);
nand U24719 (N_24719,N_24437,N_24407);
xnor U24720 (N_24720,N_24488,N_24429);
and U24721 (N_24721,N_24560,N_24467);
and U24722 (N_24722,N_24569,N_24544);
and U24723 (N_24723,N_24457,N_24477);
or U24724 (N_24724,N_24435,N_24514);
nor U24725 (N_24725,N_24477,N_24565);
nor U24726 (N_24726,N_24411,N_24488);
or U24727 (N_24727,N_24538,N_24599);
xnor U24728 (N_24728,N_24588,N_24533);
xor U24729 (N_24729,N_24520,N_24427);
nand U24730 (N_24730,N_24554,N_24450);
and U24731 (N_24731,N_24588,N_24451);
nor U24732 (N_24732,N_24423,N_24587);
and U24733 (N_24733,N_24571,N_24491);
nor U24734 (N_24734,N_24565,N_24460);
or U24735 (N_24735,N_24460,N_24470);
xnor U24736 (N_24736,N_24426,N_24432);
nor U24737 (N_24737,N_24400,N_24451);
nor U24738 (N_24738,N_24569,N_24551);
and U24739 (N_24739,N_24493,N_24536);
nor U24740 (N_24740,N_24446,N_24467);
and U24741 (N_24741,N_24535,N_24487);
nand U24742 (N_24742,N_24441,N_24403);
or U24743 (N_24743,N_24530,N_24481);
nor U24744 (N_24744,N_24555,N_24462);
nor U24745 (N_24745,N_24528,N_24437);
or U24746 (N_24746,N_24531,N_24472);
nand U24747 (N_24747,N_24519,N_24422);
nand U24748 (N_24748,N_24524,N_24423);
nand U24749 (N_24749,N_24532,N_24596);
nor U24750 (N_24750,N_24503,N_24512);
nor U24751 (N_24751,N_24511,N_24460);
and U24752 (N_24752,N_24513,N_24570);
xnor U24753 (N_24753,N_24531,N_24528);
or U24754 (N_24754,N_24408,N_24586);
nor U24755 (N_24755,N_24497,N_24481);
nor U24756 (N_24756,N_24526,N_24583);
nor U24757 (N_24757,N_24426,N_24442);
nand U24758 (N_24758,N_24546,N_24557);
nand U24759 (N_24759,N_24535,N_24531);
xnor U24760 (N_24760,N_24461,N_24411);
and U24761 (N_24761,N_24462,N_24456);
and U24762 (N_24762,N_24589,N_24478);
or U24763 (N_24763,N_24426,N_24576);
nor U24764 (N_24764,N_24469,N_24503);
nand U24765 (N_24765,N_24536,N_24529);
nand U24766 (N_24766,N_24588,N_24571);
or U24767 (N_24767,N_24525,N_24444);
and U24768 (N_24768,N_24458,N_24442);
or U24769 (N_24769,N_24407,N_24534);
nand U24770 (N_24770,N_24581,N_24462);
or U24771 (N_24771,N_24512,N_24580);
xor U24772 (N_24772,N_24580,N_24404);
nand U24773 (N_24773,N_24494,N_24587);
nor U24774 (N_24774,N_24475,N_24568);
nor U24775 (N_24775,N_24563,N_24562);
nor U24776 (N_24776,N_24434,N_24460);
and U24777 (N_24777,N_24535,N_24428);
xor U24778 (N_24778,N_24450,N_24501);
and U24779 (N_24779,N_24435,N_24524);
nand U24780 (N_24780,N_24538,N_24453);
nor U24781 (N_24781,N_24589,N_24410);
xnor U24782 (N_24782,N_24481,N_24435);
or U24783 (N_24783,N_24547,N_24575);
xnor U24784 (N_24784,N_24563,N_24419);
or U24785 (N_24785,N_24557,N_24492);
and U24786 (N_24786,N_24441,N_24471);
and U24787 (N_24787,N_24528,N_24579);
and U24788 (N_24788,N_24450,N_24587);
and U24789 (N_24789,N_24499,N_24536);
nor U24790 (N_24790,N_24487,N_24566);
and U24791 (N_24791,N_24589,N_24488);
xor U24792 (N_24792,N_24568,N_24547);
xnor U24793 (N_24793,N_24408,N_24513);
nor U24794 (N_24794,N_24546,N_24585);
and U24795 (N_24795,N_24456,N_24563);
xor U24796 (N_24796,N_24468,N_24492);
nor U24797 (N_24797,N_24561,N_24509);
xnor U24798 (N_24798,N_24439,N_24589);
nand U24799 (N_24799,N_24486,N_24520);
and U24800 (N_24800,N_24612,N_24760);
nor U24801 (N_24801,N_24615,N_24781);
or U24802 (N_24802,N_24769,N_24716);
xnor U24803 (N_24803,N_24604,N_24703);
nor U24804 (N_24804,N_24680,N_24623);
and U24805 (N_24805,N_24658,N_24639);
nor U24806 (N_24806,N_24793,N_24713);
and U24807 (N_24807,N_24678,N_24682);
xor U24808 (N_24808,N_24690,N_24730);
and U24809 (N_24809,N_24752,N_24662);
and U24810 (N_24810,N_24686,N_24633);
xor U24811 (N_24811,N_24607,N_24627);
nor U24812 (N_24812,N_24700,N_24715);
nand U24813 (N_24813,N_24726,N_24704);
nand U24814 (N_24814,N_24702,N_24799);
nor U24815 (N_24815,N_24605,N_24744);
or U24816 (N_24816,N_24635,N_24624);
nor U24817 (N_24817,N_24733,N_24628);
nor U24818 (N_24818,N_24750,N_24746);
nand U24819 (N_24819,N_24664,N_24653);
nor U24820 (N_24820,N_24668,N_24785);
and U24821 (N_24821,N_24729,N_24663);
and U24822 (N_24822,N_24641,N_24728);
or U24823 (N_24823,N_24606,N_24698);
nand U24824 (N_24824,N_24631,N_24707);
or U24825 (N_24825,N_24676,N_24789);
or U24826 (N_24826,N_24667,N_24650);
xor U24827 (N_24827,N_24669,N_24642);
or U24828 (N_24828,N_24688,N_24780);
or U24829 (N_24829,N_24665,N_24717);
xnor U24830 (N_24830,N_24768,N_24741);
xor U24831 (N_24831,N_24720,N_24613);
nor U24832 (N_24832,N_24779,N_24685);
nand U24833 (N_24833,N_24721,N_24766);
nand U24834 (N_24834,N_24655,N_24791);
and U24835 (N_24835,N_24652,N_24687);
nor U24836 (N_24836,N_24699,N_24681);
nor U24837 (N_24837,N_24727,N_24626);
nor U24838 (N_24838,N_24740,N_24784);
or U24839 (N_24839,N_24666,N_24731);
and U24840 (N_24840,N_24625,N_24646);
xnor U24841 (N_24841,N_24755,N_24745);
nand U24842 (N_24842,N_24660,N_24651);
and U24843 (N_24843,N_24659,N_24759);
and U24844 (N_24844,N_24767,N_24754);
and U24845 (N_24845,N_24679,N_24683);
and U24846 (N_24846,N_24748,N_24692);
xnor U24847 (N_24847,N_24725,N_24647);
nand U24848 (N_24848,N_24697,N_24790);
or U24849 (N_24849,N_24691,N_24674);
nand U24850 (N_24850,N_24693,N_24775);
xor U24851 (N_24851,N_24718,N_24708);
and U24852 (N_24852,N_24621,N_24645);
nand U24853 (N_24853,N_24787,N_24735);
and U24854 (N_24854,N_24763,N_24603);
xnor U24855 (N_24855,N_24712,N_24638);
xor U24856 (N_24856,N_24762,N_24709);
xor U24857 (N_24857,N_24694,N_24643);
nand U24858 (N_24858,N_24701,N_24634);
xnor U24859 (N_24859,N_24788,N_24714);
xnor U24860 (N_24860,N_24777,N_24757);
xor U24861 (N_24861,N_24614,N_24742);
nand U24862 (N_24862,N_24786,N_24747);
xnor U24863 (N_24863,N_24739,N_24719);
or U24864 (N_24864,N_24602,N_24619);
nor U24865 (N_24865,N_24797,N_24618);
xnor U24866 (N_24866,N_24776,N_24629);
and U24867 (N_24867,N_24636,N_24611);
and U24868 (N_24868,N_24657,N_24770);
nor U24869 (N_24869,N_24616,N_24796);
xor U24870 (N_24870,N_24795,N_24782);
or U24871 (N_24871,N_24600,N_24783);
xor U24872 (N_24872,N_24671,N_24749);
and U24873 (N_24873,N_24772,N_24723);
or U24874 (N_24874,N_24711,N_24738);
nor U24875 (N_24875,N_24798,N_24737);
nor U24876 (N_24876,N_24771,N_24656);
and U24877 (N_24877,N_24610,N_24644);
and U24878 (N_24878,N_24758,N_24695);
xnor U24879 (N_24879,N_24753,N_24608);
nand U24880 (N_24880,N_24609,N_24632);
nand U24881 (N_24881,N_24620,N_24764);
nand U24882 (N_24882,N_24705,N_24696);
and U24883 (N_24883,N_24672,N_24601);
nand U24884 (N_24884,N_24675,N_24649);
nor U24885 (N_24885,N_24773,N_24734);
or U24886 (N_24886,N_24689,N_24722);
xor U24887 (N_24887,N_24654,N_24736);
and U24888 (N_24888,N_24630,N_24617);
nor U24889 (N_24889,N_24684,N_24640);
nand U24890 (N_24890,N_24732,N_24706);
xor U24891 (N_24891,N_24751,N_24661);
xnor U24892 (N_24892,N_24622,N_24710);
or U24893 (N_24893,N_24792,N_24774);
nand U24894 (N_24894,N_24673,N_24794);
or U24895 (N_24895,N_24761,N_24670);
nor U24896 (N_24896,N_24765,N_24743);
nor U24897 (N_24897,N_24724,N_24648);
nor U24898 (N_24898,N_24677,N_24756);
nor U24899 (N_24899,N_24778,N_24637);
xnor U24900 (N_24900,N_24722,N_24743);
nor U24901 (N_24901,N_24737,N_24604);
or U24902 (N_24902,N_24773,N_24658);
xnor U24903 (N_24903,N_24641,N_24722);
nand U24904 (N_24904,N_24724,N_24612);
or U24905 (N_24905,N_24781,N_24680);
or U24906 (N_24906,N_24790,N_24729);
xor U24907 (N_24907,N_24682,N_24649);
xor U24908 (N_24908,N_24680,N_24634);
and U24909 (N_24909,N_24745,N_24703);
or U24910 (N_24910,N_24630,N_24764);
xnor U24911 (N_24911,N_24703,N_24669);
xor U24912 (N_24912,N_24749,N_24637);
or U24913 (N_24913,N_24648,N_24656);
xor U24914 (N_24914,N_24678,N_24668);
nor U24915 (N_24915,N_24761,N_24665);
nand U24916 (N_24916,N_24654,N_24650);
and U24917 (N_24917,N_24700,N_24678);
nor U24918 (N_24918,N_24755,N_24792);
xor U24919 (N_24919,N_24714,N_24606);
and U24920 (N_24920,N_24761,N_24745);
and U24921 (N_24921,N_24708,N_24698);
nor U24922 (N_24922,N_24690,N_24792);
and U24923 (N_24923,N_24653,N_24796);
or U24924 (N_24924,N_24686,N_24758);
xor U24925 (N_24925,N_24695,N_24716);
and U24926 (N_24926,N_24655,N_24691);
or U24927 (N_24927,N_24751,N_24742);
xor U24928 (N_24928,N_24638,N_24654);
xnor U24929 (N_24929,N_24617,N_24755);
and U24930 (N_24930,N_24785,N_24773);
and U24931 (N_24931,N_24778,N_24794);
or U24932 (N_24932,N_24668,N_24738);
xnor U24933 (N_24933,N_24647,N_24653);
and U24934 (N_24934,N_24626,N_24796);
xor U24935 (N_24935,N_24650,N_24644);
or U24936 (N_24936,N_24768,N_24714);
nor U24937 (N_24937,N_24638,N_24772);
nand U24938 (N_24938,N_24653,N_24678);
xor U24939 (N_24939,N_24756,N_24686);
nor U24940 (N_24940,N_24611,N_24723);
and U24941 (N_24941,N_24601,N_24738);
nand U24942 (N_24942,N_24700,N_24781);
or U24943 (N_24943,N_24684,N_24645);
nor U24944 (N_24944,N_24724,N_24679);
nor U24945 (N_24945,N_24767,N_24738);
xnor U24946 (N_24946,N_24684,N_24611);
and U24947 (N_24947,N_24708,N_24663);
or U24948 (N_24948,N_24619,N_24799);
xor U24949 (N_24949,N_24751,N_24752);
nor U24950 (N_24950,N_24763,N_24646);
or U24951 (N_24951,N_24746,N_24648);
or U24952 (N_24952,N_24707,N_24661);
xor U24953 (N_24953,N_24641,N_24663);
nor U24954 (N_24954,N_24782,N_24742);
or U24955 (N_24955,N_24695,N_24788);
nor U24956 (N_24956,N_24620,N_24690);
or U24957 (N_24957,N_24634,N_24647);
nor U24958 (N_24958,N_24652,N_24665);
or U24959 (N_24959,N_24751,N_24630);
and U24960 (N_24960,N_24752,N_24690);
nor U24961 (N_24961,N_24634,N_24754);
or U24962 (N_24962,N_24689,N_24720);
and U24963 (N_24963,N_24741,N_24766);
nor U24964 (N_24964,N_24691,N_24743);
and U24965 (N_24965,N_24778,N_24766);
or U24966 (N_24966,N_24776,N_24649);
nand U24967 (N_24967,N_24624,N_24612);
and U24968 (N_24968,N_24610,N_24622);
and U24969 (N_24969,N_24655,N_24665);
xor U24970 (N_24970,N_24628,N_24623);
and U24971 (N_24971,N_24611,N_24783);
xor U24972 (N_24972,N_24719,N_24715);
and U24973 (N_24973,N_24643,N_24655);
xnor U24974 (N_24974,N_24743,N_24648);
xor U24975 (N_24975,N_24701,N_24732);
xnor U24976 (N_24976,N_24738,N_24667);
and U24977 (N_24977,N_24693,N_24737);
nor U24978 (N_24978,N_24701,N_24721);
nor U24979 (N_24979,N_24638,N_24721);
nor U24980 (N_24980,N_24768,N_24628);
and U24981 (N_24981,N_24767,N_24783);
and U24982 (N_24982,N_24641,N_24747);
xnor U24983 (N_24983,N_24611,N_24614);
xnor U24984 (N_24984,N_24719,N_24736);
or U24985 (N_24985,N_24710,N_24723);
and U24986 (N_24986,N_24624,N_24659);
or U24987 (N_24987,N_24626,N_24774);
or U24988 (N_24988,N_24698,N_24652);
xor U24989 (N_24989,N_24636,N_24635);
xor U24990 (N_24990,N_24775,N_24649);
or U24991 (N_24991,N_24769,N_24613);
nand U24992 (N_24992,N_24731,N_24678);
xnor U24993 (N_24993,N_24728,N_24633);
nor U24994 (N_24994,N_24757,N_24614);
or U24995 (N_24995,N_24640,N_24697);
and U24996 (N_24996,N_24680,N_24794);
xor U24997 (N_24997,N_24761,N_24635);
xor U24998 (N_24998,N_24653,N_24645);
xor U24999 (N_24999,N_24686,N_24701);
nor U25000 (N_25000,N_24959,N_24896);
nor U25001 (N_25001,N_24884,N_24857);
xor U25002 (N_25002,N_24991,N_24881);
xor U25003 (N_25003,N_24973,N_24967);
nor U25004 (N_25004,N_24862,N_24990);
and U25005 (N_25005,N_24870,N_24968);
and U25006 (N_25006,N_24957,N_24951);
xnor U25007 (N_25007,N_24978,N_24874);
and U25008 (N_25008,N_24989,N_24969);
nor U25009 (N_25009,N_24812,N_24813);
xnor U25010 (N_25010,N_24810,N_24849);
xor U25011 (N_25011,N_24992,N_24828);
xnor U25012 (N_25012,N_24816,N_24966);
and U25013 (N_25013,N_24859,N_24909);
nand U25014 (N_25014,N_24893,N_24863);
or U25015 (N_25015,N_24977,N_24956);
and U25016 (N_25016,N_24904,N_24811);
or U25017 (N_25017,N_24926,N_24885);
xnor U25018 (N_25018,N_24901,N_24800);
nand U25019 (N_25019,N_24984,N_24808);
nor U25020 (N_25020,N_24936,N_24839);
xor U25021 (N_25021,N_24850,N_24981);
nand U25022 (N_25022,N_24910,N_24925);
nor U25023 (N_25023,N_24891,N_24847);
xor U25024 (N_25024,N_24994,N_24948);
nor U25025 (N_25025,N_24982,N_24905);
nand U25026 (N_25026,N_24840,N_24916);
and U25027 (N_25027,N_24950,N_24817);
xnor U25028 (N_25028,N_24887,N_24941);
and U25029 (N_25029,N_24979,N_24815);
and U25030 (N_25030,N_24932,N_24807);
xnor U25031 (N_25031,N_24927,N_24976);
and U25032 (N_25032,N_24928,N_24879);
nand U25033 (N_25033,N_24802,N_24983);
nand U25034 (N_25034,N_24939,N_24987);
and U25035 (N_25035,N_24876,N_24906);
xnor U25036 (N_25036,N_24903,N_24820);
or U25037 (N_25037,N_24919,N_24843);
or U25038 (N_25038,N_24902,N_24921);
or U25039 (N_25039,N_24853,N_24866);
and U25040 (N_25040,N_24934,N_24917);
xnor U25041 (N_25041,N_24940,N_24995);
nand U25042 (N_25042,N_24875,N_24865);
or U25043 (N_25043,N_24846,N_24942);
nand U25044 (N_25044,N_24999,N_24837);
nand U25045 (N_25045,N_24914,N_24821);
and U25046 (N_25046,N_24898,N_24868);
or U25047 (N_25047,N_24915,N_24964);
and U25048 (N_25048,N_24897,N_24972);
xnor U25049 (N_25049,N_24908,N_24835);
xor U25050 (N_25050,N_24924,N_24923);
or U25051 (N_25051,N_24831,N_24971);
nand U25052 (N_25052,N_24848,N_24899);
and U25053 (N_25053,N_24830,N_24986);
or U25054 (N_25054,N_24827,N_24814);
and U25055 (N_25055,N_24851,N_24993);
nor U25056 (N_25056,N_24829,N_24877);
and U25057 (N_25057,N_24854,N_24911);
xnor U25058 (N_25058,N_24935,N_24996);
or U25059 (N_25059,N_24900,N_24861);
or U25060 (N_25060,N_24801,N_24842);
and U25061 (N_25061,N_24892,N_24920);
and U25062 (N_25062,N_24947,N_24946);
and U25063 (N_25063,N_24985,N_24883);
xor U25064 (N_25064,N_24895,N_24980);
nor U25065 (N_25065,N_24955,N_24867);
or U25066 (N_25066,N_24852,N_24871);
xnor U25067 (N_25067,N_24889,N_24878);
and U25068 (N_25068,N_24945,N_24818);
nor U25069 (N_25069,N_24949,N_24844);
and U25070 (N_25070,N_24933,N_24890);
nand U25071 (N_25071,N_24804,N_24819);
nand U25072 (N_25072,N_24922,N_24834);
nor U25073 (N_25073,N_24825,N_24912);
and U25074 (N_25074,N_24974,N_24886);
xor U25075 (N_25075,N_24832,N_24826);
nor U25076 (N_25076,N_24860,N_24894);
or U25077 (N_25077,N_24962,N_24869);
nand U25078 (N_25078,N_24931,N_24856);
or U25079 (N_25079,N_24988,N_24970);
nor U25080 (N_25080,N_24913,N_24809);
nor U25081 (N_25081,N_24805,N_24803);
and U25082 (N_25082,N_24873,N_24975);
nor U25083 (N_25083,N_24838,N_24888);
nor U25084 (N_25084,N_24944,N_24997);
or U25085 (N_25085,N_24963,N_24961);
and U25086 (N_25086,N_24806,N_24937);
nor U25087 (N_25087,N_24858,N_24864);
and U25088 (N_25088,N_24907,N_24930);
nand U25089 (N_25089,N_24822,N_24954);
nand U25090 (N_25090,N_24823,N_24938);
nor U25091 (N_25091,N_24880,N_24958);
xor U25092 (N_25092,N_24960,N_24953);
nor U25093 (N_25093,N_24952,N_24965);
or U25094 (N_25094,N_24998,N_24824);
xnor U25095 (N_25095,N_24833,N_24918);
nand U25096 (N_25096,N_24845,N_24836);
xor U25097 (N_25097,N_24872,N_24943);
nor U25098 (N_25098,N_24841,N_24882);
nand U25099 (N_25099,N_24929,N_24855);
and U25100 (N_25100,N_24880,N_24933);
nand U25101 (N_25101,N_24944,N_24845);
or U25102 (N_25102,N_24930,N_24807);
or U25103 (N_25103,N_24860,N_24972);
nor U25104 (N_25104,N_24885,N_24956);
nor U25105 (N_25105,N_24801,N_24807);
or U25106 (N_25106,N_24951,N_24908);
nor U25107 (N_25107,N_24803,N_24942);
xnor U25108 (N_25108,N_24816,N_24849);
nor U25109 (N_25109,N_24905,N_24913);
nand U25110 (N_25110,N_24985,N_24943);
and U25111 (N_25111,N_24970,N_24986);
xnor U25112 (N_25112,N_24926,N_24864);
xor U25113 (N_25113,N_24912,N_24892);
and U25114 (N_25114,N_24982,N_24974);
and U25115 (N_25115,N_24980,N_24807);
and U25116 (N_25116,N_24985,N_24807);
nor U25117 (N_25117,N_24929,N_24893);
xnor U25118 (N_25118,N_24807,N_24914);
and U25119 (N_25119,N_24851,N_24946);
xnor U25120 (N_25120,N_24812,N_24840);
or U25121 (N_25121,N_24845,N_24809);
nor U25122 (N_25122,N_24818,N_24813);
and U25123 (N_25123,N_24902,N_24910);
or U25124 (N_25124,N_24878,N_24811);
nand U25125 (N_25125,N_24858,N_24922);
or U25126 (N_25126,N_24827,N_24961);
nand U25127 (N_25127,N_24982,N_24853);
nand U25128 (N_25128,N_24937,N_24945);
and U25129 (N_25129,N_24974,N_24981);
xor U25130 (N_25130,N_24850,N_24870);
nand U25131 (N_25131,N_24914,N_24938);
xnor U25132 (N_25132,N_24825,N_24889);
and U25133 (N_25133,N_24938,N_24972);
nor U25134 (N_25134,N_24907,N_24953);
and U25135 (N_25135,N_24985,N_24955);
or U25136 (N_25136,N_24843,N_24855);
nand U25137 (N_25137,N_24964,N_24860);
or U25138 (N_25138,N_24960,N_24918);
or U25139 (N_25139,N_24964,N_24802);
nand U25140 (N_25140,N_24933,N_24840);
nand U25141 (N_25141,N_24828,N_24857);
xor U25142 (N_25142,N_24818,N_24917);
nor U25143 (N_25143,N_24899,N_24831);
nor U25144 (N_25144,N_24850,N_24943);
or U25145 (N_25145,N_24912,N_24837);
or U25146 (N_25146,N_24909,N_24861);
nor U25147 (N_25147,N_24840,N_24837);
nor U25148 (N_25148,N_24870,N_24987);
nand U25149 (N_25149,N_24934,N_24943);
or U25150 (N_25150,N_24917,N_24895);
xnor U25151 (N_25151,N_24858,N_24803);
nand U25152 (N_25152,N_24890,N_24840);
xor U25153 (N_25153,N_24847,N_24900);
and U25154 (N_25154,N_24896,N_24884);
xor U25155 (N_25155,N_24802,N_24904);
xnor U25156 (N_25156,N_24808,N_24830);
nand U25157 (N_25157,N_24948,N_24936);
and U25158 (N_25158,N_24927,N_24991);
nor U25159 (N_25159,N_24948,N_24989);
xor U25160 (N_25160,N_24927,N_24987);
xor U25161 (N_25161,N_24811,N_24980);
nand U25162 (N_25162,N_24808,N_24928);
nand U25163 (N_25163,N_24918,N_24907);
and U25164 (N_25164,N_24871,N_24822);
nand U25165 (N_25165,N_24905,N_24801);
nand U25166 (N_25166,N_24967,N_24937);
or U25167 (N_25167,N_24933,N_24884);
xor U25168 (N_25168,N_24916,N_24878);
and U25169 (N_25169,N_24849,N_24813);
and U25170 (N_25170,N_24827,N_24955);
and U25171 (N_25171,N_24906,N_24997);
xnor U25172 (N_25172,N_24831,N_24824);
xor U25173 (N_25173,N_24803,N_24895);
or U25174 (N_25174,N_24918,N_24959);
or U25175 (N_25175,N_24924,N_24939);
and U25176 (N_25176,N_24931,N_24800);
nor U25177 (N_25177,N_24875,N_24850);
xor U25178 (N_25178,N_24893,N_24895);
and U25179 (N_25179,N_24906,N_24825);
xor U25180 (N_25180,N_24986,N_24878);
nor U25181 (N_25181,N_24974,N_24818);
or U25182 (N_25182,N_24957,N_24814);
and U25183 (N_25183,N_24884,N_24914);
nand U25184 (N_25184,N_24889,N_24855);
nor U25185 (N_25185,N_24830,N_24954);
and U25186 (N_25186,N_24846,N_24803);
nor U25187 (N_25187,N_24954,N_24986);
and U25188 (N_25188,N_24865,N_24890);
or U25189 (N_25189,N_24961,N_24854);
and U25190 (N_25190,N_24972,N_24929);
or U25191 (N_25191,N_24805,N_24854);
nor U25192 (N_25192,N_24939,N_24963);
nor U25193 (N_25193,N_24916,N_24952);
nor U25194 (N_25194,N_24892,N_24937);
nor U25195 (N_25195,N_24801,N_24887);
and U25196 (N_25196,N_24959,N_24812);
or U25197 (N_25197,N_24909,N_24888);
nor U25198 (N_25198,N_24817,N_24818);
or U25199 (N_25199,N_24805,N_24836);
nand U25200 (N_25200,N_25127,N_25119);
and U25201 (N_25201,N_25148,N_25114);
nor U25202 (N_25202,N_25049,N_25039);
nand U25203 (N_25203,N_25053,N_25069);
nand U25204 (N_25204,N_25028,N_25124);
xor U25205 (N_25205,N_25099,N_25160);
or U25206 (N_25206,N_25094,N_25137);
nand U25207 (N_25207,N_25169,N_25187);
or U25208 (N_25208,N_25075,N_25154);
or U25209 (N_25209,N_25034,N_25171);
nor U25210 (N_25210,N_25164,N_25022);
nor U25211 (N_25211,N_25087,N_25091);
or U25212 (N_25212,N_25088,N_25122);
nor U25213 (N_25213,N_25002,N_25000);
xnor U25214 (N_25214,N_25141,N_25048);
nand U25215 (N_25215,N_25071,N_25018);
nand U25216 (N_25216,N_25168,N_25131);
or U25217 (N_25217,N_25103,N_25068);
xor U25218 (N_25218,N_25078,N_25150);
and U25219 (N_25219,N_25090,N_25085);
nor U25220 (N_25220,N_25092,N_25023);
nand U25221 (N_25221,N_25024,N_25035);
xor U25222 (N_25222,N_25045,N_25192);
nor U25223 (N_25223,N_25152,N_25153);
xor U25224 (N_25224,N_25161,N_25107);
xor U25225 (N_25225,N_25005,N_25194);
nor U25226 (N_25226,N_25142,N_25033);
or U25227 (N_25227,N_25101,N_25112);
or U25228 (N_25228,N_25042,N_25040);
nand U25229 (N_25229,N_25066,N_25146);
xnor U25230 (N_25230,N_25063,N_25104);
xnor U25231 (N_25231,N_25003,N_25166);
or U25232 (N_25232,N_25081,N_25108);
and U25233 (N_25233,N_25004,N_25084);
or U25234 (N_25234,N_25062,N_25181);
and U25235 (N_25235,N_25100,N_25126);
nor U25236 (N_25236,N_25032,N_25138);
nor U25237 (N_25237,N_25155,N_25109);
xor U25238 (N_25238,N_25129,N_25193);
or U25239 (N_25239,N_25174,N_25056);
nor U25240 (N_25240,N_25076,N_25008);
xnor U25241 (N_25241,N_25183,N_25089);
nor U25242 (N_25242,N_25013,N_25149);
and U25243 (N_25243,N_25098,N_25030);
xnor U25244 (N_25244,N_25135,N_25180);
or U25245 (N_25245,N_25050,N_25134);
nand U25246 (N_25246,N_25133,N_25041);
or U25247 (N_25247,N_25176,N_25027);
and U25248 (N_25248,N_25191,N_25009);
nand U25249 (N_25249,N_25199,N_25029);
or U25250 (N_25250,N_25197,N_25059);
xor U25251 (N_25251,N_25070,N_25057);
or U25252 (N_25252,N_25026,N_25110);
nand U25253 (N_25253,N_25061,N_25172);
xor U25254 (N_25254,N_25095,N_25118);
xnor U25255 (N_25255,N_25182,N_25060);
and U25256 (N_25256,N_25198,N_25007);
and U25257 (N_25257,N_25055,N_25188);
xnor U25258 (N_25258,N_25116,N_25177);
nand U25259 (N_25259,N_25143,N_25178);
nor U25260 (N_25260,N_25051,N_25046);
nand U25261 (N_25261,N_25031,N_25189);
nor U25262 (N_25262,N_25147,N_25117);
xor U25263 (N_25263,N_25132,N_25025);
or U25264 (N_25264,N_25020,N_25190);
nor U25265 (N_25265,N_25157,N_25083);
and U25266 (N_25266,N_25120,N_25130);
xnor U25267 (N_25267,N_25052,N_25111);
and U25268 (N_25268,N_25011,N_25006);
xor U25269 (N_25269,N_25077,N_25021);
and U25270 (N_25270,N_25058,N_25065);
and U25271 (N_25271,N_25047,N_25170);
xnor U25272 (N_25272,N_25082,N_25017);
nor U25273 (N_25273,N_25093,N_25015);
nand U25274 (N_25274,N_25037,N_25128);
xor U25275 (N_25275,N_25139,N_25145);
or U25276 (N_25276,N_25184,N_25067);
or U25277 (N_25277,N_25136,N_25165);
xnor U25278 (N_25278,N_25072,N_25156);
nand U25279 (N_25279,N_25151,N_25105);
nor U25280 (N_25280,N_25086,N_25175);
nand U25281 (N_25281,N_25097,N_25162);
xor U25282 (N_25282,N_25173,N_25106);
and U25283 (N_25283,N_25159,N_25179);
nand U25284 (N_25284,N_25038,N_25036);
xor U25285 (N_25285,N_25115,N_25012);
and U25286 (N_25286,N_25079,N_25096);
nor U25287 (N_25287,N_25186,N_25125);
nor U25288 (N_25288,N_25016,N_25010);
or U25289 (N_25289,N_25074,N_25140);
and U25290 (N_25290,N_25064,N_25144);
and U25291 (N_25291,N_25001,N_25044);
and U25292 (N_25292,N_25196,N_25158);
nand U25293 (N_25293,N_25073,N_25080);
xnor U25294 (N_25294,N_25102,N_25167);
nor U25295 (N_25295,N_25163,N_25043);
and U25296 (N_25296,N_25123,N_25014);
and U25297 (N_25297,N_25054,N_25121);
xor U25298 (N_25298,N_25113,N_25195);
and U25299 (N_25299,N_25019,N_25185);
or U25300 (N_25300,N_25118,N_25024);
or U25301 (N_25301,N_25016,N_25029);
nand U25302 (N_25302,N_25188,N_25175);
xor U25303 (N_25303,N_25113,N_25072);
or U25304 (N_25304,N_25111,N_25104);
and U25305 (N_25305,N_25113,N_25010);
and U25306 (N_25306,N_25135,N_25036);
nand U25307 (N_25307,N_25183,N_25187);
nand U25308 (N_25308,N_25012,N_25196);
and U25309 (N_25309,N_25085,N_25116);
xor U25310 (N_25310,N_25064,N_25019);
or U25311 (N_25311,N_25020,N_25129);
xor U25312 (N_25312,N_25141,N_25096);
and U25313 (N_25313,N_25195,N_25077);
and U25314 (N_25314,N_25120,N_25030);
or U25315 (N_25315,N_25026,N_25059);
or U25316 (N_25316,N_25192,N_25169);
nor U25317 (N_25317,N_25036,N_25021);
or U25318 (N_25318,N_25012,N_25168);
or U25319 (N_25319,N_25037,N_25068);
nor U25320 (N_25320,N_25166,N_25007);
and U25321 (N_25321,N_25172,N_25153);
nand U25322 (N_25322,N_25086,N_25127);
or U25323 (N_25323,N_25090,N_25150);
and U25324 (N_25324,N_25086,N_25133);
xor U25325 (N_25325,N_25003,N_25037);
xnor U25326 (N_25326,N_25104,N_25092);
nor U25327 (N_25327,N_25068,N_25010);
or U25328 (N_25328,N_25004,N_25018);
nand U25329 (N_25329,N_25164,N_25027);
or U25330 (N_25330,N_25157,N_25107);
nand U25331 (N_25331,N_25185,N_25045);
nand U25332 (N_25332,N_25185,N_25056);
nand U25333 (N_25333,N_25068,N_25073);
xnor U25334 (N_25334,N_25077,N_25010);
or U25335 (N_25335,N_25106,N_25080);
xnor U25336 (N_25336,N_25165,N_25042);
nand U25337 (N_25337,N_25144,N_25156);
xor U25338 (N_25338,N_25173,N_25158);
nand U25339 (N_25339,N_25010,N_25091);
nor U25340 (N_25340,N_25114,N_25141);
and U25341 (N_25341,N_25154,N_25080);
xor U25342 (N_25342,N_25111,N_25053);
nor U25343 (N_25343,N_25014,N_25001);
and U25344 (N_25344,N_25199,N_25192);
and U25345 (N_25345,N_25005,N_25179);
or U25346 (N_25346,N_25002,N_25062);
xnor U25347 (N_25347,N_25107,N_25087);
and U25348 (N_25348,N_25015,N_25146);
and U25349 (N_25349,N_25158,N_25071);
and U25350 (N_25350,N_25163,N_25174);
nand U25351 (N_25351,N_25117,N_25106);
xor U25352 (N_25352,N_25027,N_25007);
nand U25353 (N_25353,N_25138,N_25024);
xor U25354 (N_25354,N_25041,N_25033);
nand U25355 (N_25355,N_25083,N_25120);
nor U25356 (N_25356,N_25184,N_25022);
xor U25357 (N_25357,N_25169,N_25049);
or U25358 (N_25358,N_25170,N_25103);
nor U25359 (N_25359,N_25159,N_25153);
nand U25360 (N_25360,N_25009,N_25038);
and U25361 (N_25361,N_25094,N_25125);
xnor U25362 (N_25362,N_25031,N_25009);
nand U25363 (N_25363,N_25011,N_25105);
and U25364 (N_25364,N_25010,N_25147);
or U25365 (N_25365,N_25128,N_25097);
or U25366 (N_25366,N_25091,N_25026);
xnor U25367 (N_25367,N_25128,N_25079);
xnor U25368 (N_25368,N_25050,N_25084);
xnor U25369 (N_25369,N_25046,N_25083);
nor U25370 (N_25370,N_25027,N_25091);
nor U25371 (N_25371,N_25053,N_25132);
nand U25372 (N_25372,N_25155,N_25084);
xnor U25373 (N_25373,N_25108,N_25167);
or U25374 (N_25374,N_25179,N_25156);
and U25375 (N_25375,N_25088,N_25000);
xor U25376 (N_25376,N_25000,N_25175);
nand U25377 (N_25377,N_25044,N_25125);
xor U25378 (N_25378,N_25086,N_25123);
nand U25379 (N_25379,N_25141,N_25191);
or U25380 (N_25380,N_25099,N_25045);
xor U25381 (N_25381,N_25129,N_25110);
xor U25382 (N_25382,N_25197,N_25042);
nand U25383 (N_25383,N_25056,N_25081);
nand U25384 (N_25384,N_25034,N_25128);
nor U25385 (N_25385,N_25177,N_25048);
nand U25386 (N_25386,N_25103,N_25168);
xor U25387 (N_25387,N_25101,N_25135);
nor U25388 (N_25388,N_25009,N_25059);
and U25389 (N_25389,N_25165,N_25117);
xor U25390 (N_25390,N_25035,N_25113);
nand U25391 (N_25391,N_25090,N_25113);
or U25392 (N_25392,N_25076,N_25031);
or U25393 (N_25393,N_25100,N_25039);
and U25394 (N_25394,N_25192,N_25191);
nand U25395 (N_25395,N_25147,N_25096);
and U25396 (N_25396,N_25001,N_25127);
and U25397 (N_25397,N_25070,N_25120);
nand U25398 (N_25398,N_25079,N_25132);
nand U25399 (N_25399,N_25001,N_25176);
nor U25400 (N_25400,N_25303,N_25305);
xnor U25401 (N_25401,N_25315,N_25270);
or U25402 (N_25402,N_25298,N_25360);
nand U25403 (N_25403,N_25377,N_25371);
nand U25404 (N_25404,N_25275,N_25258);
and U25405 (N_25405,N_25257,N_25224);
nor U25406 (N_25406,N_25314,N_25326);
and U25407 (N_25407,N_25240,N_25344);
nor U25408 (N_25408,N_25312,N_25288);
xor U25409 (N_25409,N_25286,N_25376);
and U25410 (N_25410,N_25217,N_25277);
and U25411 (N_25411,N_25320,N_25244);
nand U25412 (N_25412,N_25334,N_25278);
and U25413 (N_25413,N_25285,N_25398);
nand U25414 (N_25414,N_25226,N_25323);
and U25415 (N_25415,N_25297,N_25392);
xnor U25416 (N_25416,N_25389,N_25336);
nand U25417 (N_25417,N_25221,N_25200);
or U25418 (N_25418,N_25208,N_25386);
xnor U25419 (N_25419,N_25212,N_25296);
and U25420 (N_25420,N_25317,N_25375);
nand U25421 (N_25421,N_25372,N_25316);
nand U25422 (N_25422,N_25263,N_25370);
xor U25423 (N_25423,N_25337,N_25255);
nand U25424 (N_25424,N_25391,N_25361);
nor U25425 (N_25425,N_25246,N_25333);
and U25426 (N_25426,N_25249,N_25346);
and U25427 (N_25427,N_25207,N_25247);
and U25428 (N_25428,N_25262,N_25385);
and U25429 (N_25429,N_25382,N_25243);
nor U25430 (N_25430,N_25281,N_25374);
or U25431 (N_25431,N_25219,N_25397);
or U25432 (N_25432,N_25345,N_25353);
xnor U25433 (N_25433,N_25310,N_25299);
nand U25434 (N_25434,N_25248,N_25307);
and U25435 (N_25435,N_25289,N_25313);
and U25436 (N_25436,N_25276,N_25261);
xnor U25437 (N_25437,N_25206,N_25339);
nand U25438 (N_25438,N_25352,N_25379);
nand U25439 (N_25439,N_25381,N_25232);
or U25440 (N_25440,N_25302,N_25273);
and U25441 (N_25441,N_25215,N_25209);
or U25442 (N_25442,N_25220,N_25335);
nor U25443 (N_25443,N_25292,N_25253);
and U25444 (N_25444,N_25311,N_25390);
and U25445 (N_25445,N_25349,N_25396);
or U25446 (N_25446,N_25205,N_25380);
xor U25447 (N_25447,N_25282,N_25300);
nor U25448 (N_25448,N_25254,N_25214);
xnor U25449 (N_25449,N_25319,N_25354);
and U25450 (N_25450,N_25264,N_25306);
xor U25451 (N_25451,N_25235,N_25357);
or U25452 (N_25452,N_25259,N_25387);
and U25453 (N_25453,N_25395,N_25393);
nor U25454 (N_25454,N_25364,N_25222);
nand U25455 (N_25455,N_25267,N_25227);
nor U25456 (N_25456,N_25301,N_25236);
nand U25457 (N_25457,N_25328,N_25228);
and U25458 (N_25458,N_25373,N_25308);
or U25459 (N_25459,N_25213,N_25238);
and U25460 (N_25460,N_25330,N_25241);
xor U25461 (N_25461,N_25237,N_25351);
xnor U25462 (N_25462,N_25309,N_25342);
xnor U25463 (N_25463,N_25202,N_25204);
nand U25464 (N_25464,N_25368,N_25321);
xor U25465 (N_25465,N_25340,N_25291);
nor U25466 (N_25466,N_25318,N_25304);
xnor U25467 (N_25467,N_25239,N_25329);
and U25468 (N_25468,N_25295,N_25347);
nand U25469 (N_25469,N_25230,N_25211);
and U25470 (N_25470,N_25324,N_25201);
or U25471 (N_25471,N_25274,N_25269);
nor U25472 (N_25472,N_25355,N_25362);
and U25473 (N_25473,N_25225,N_25294);
or U25474 (N_25474,N_25283,N_25325);
or U25475 (N_25475,N_25272,N_25203);
nor U25476 (N_25476,N_25266,N_25358);
xor U25477 (N_25477,N_25338,N_25363);
or U25478 (N_25478,N_25287,N_25280);
and U25479 (N_25479,N_25234,N_25210);
nor U25480 (N_25480,N_25367,N_25383);
xnor U25481 (N_25481,N_25218,N_25331);
nand U25482 (N_25482,N_25231,N_25260);
nand U25483 (N_25483,N_25216,N_25271);
nor U25484 (N_25484,N_25268,N_25341);
or U25485 (N_25485,N_25279,N_25356);
and U25486 (N_25486,N_25332,N_25327);
and U25487 (N_25487,N_25322,N_25366);
nor U25488 (N_25488,N_25256,N_25245);
nand U25489 (N_25489,N_25394,N_25233);
xor U25490 (N_25490,N_25365,N_25343);
nor U25491 (N_25491,N_25223,N_25251);
nand U25492 (N_25492,N_25359,N_25290);
nor U25493 (N_25493,N_25242,N_25284);
nor U25494 (N_25494,N_25252,N_25293);
nand U25495 (N_25495,N_25229,N_25378);
nand U25496 (N_25496,N_25384,N_25348);
xor U25497 (N_25497,N_25388,N_25265);
or U25498 (N_25498,N_25369,N_25350);
xnor U25499 (N_25499,N_25250,N_25399);
and U25500 (N_25500,N_25269,N_25249);
nand U25501 (N_25501,N_25319,N_25209);
nand U25502 (N_25502,N_25390,N_25336);
or U25503 (N_25503,N_25209,N_25218);
nor U25504 (N_25504,N_25217,N_25278);
and U25505 (N_25505,N_25353,N_25203);
xnor U25506 (N_25506,N_25372,N_25270);
and U25507 (N_25507,N_25233,N_25310);
and U25508 (N_25508,N_25320,N_25232);
nor U25509 (N_25509,N_25291,N_25273);
nand U25510 (N_25510,N_25263,N_25389);
nand U25511 (N_25511,N_25247,N_25237);
xor U25512 (N_25512,N_25227,N_25280);
and U25513 (N_25513,N_25277,N_25216);
nand U25514 (N_25514,N_25387,N_25252);
nand U25515 (N_25515,N_25340,N_25374);
or U25516 (N_25516,N_25378,N_25360);
nor U25517 (N_25517,N_25218,N_25343);
and U25518 (N_25518,N_25336,N_25378);
nor U25519 (N_25519,N_25206,N_25214);
nor U25520 (N_25520,N_25304,N_25387);
and U25521 (N_25521,N_25376,N_25375);
xor U25522 (N_25522,N_25211,N_25301);
nor U25523 (N_25523,N_25263,N_25363);
nand U25524 (N_25524,N_25201,N_25240);
and U25525 (N_25525,N_25295,N_25298);
or U25526 (N_25526,N_25278,N_25233);
or U25527 (N_25527,N_25393,N_25201);
xnor U25528 (N_25528,N_25266,N_25241);
or U25529 (N_25529,N_25250,N_25222);
nand U25530 (N_25530,N_25269,N_25309);
xnor U25531 (N_25531,N_25240,N_25282);
and U25532 (N_25532,N_25362,N_25212);
or U25533 (N_25533,N_25379,N_25335);
and U25534 (N_25534,N_25367,N_25300);
nor U25535 (N_25535,N_25395,N_25364);
and U25536 (N_25536,N_25369,N_25316);
nand U25537 (N_25537,N_25362,N_25232);
nor U25538 (N_25538,N_25375,N_25363);
and U25539 (N_25539,N_25300,N_25361);
nor U25540 (N_25540,N_25371,N_25232);
or U25541 (N_25541,N_25260,N_25379);
xnor U25542 (N_25542,N_25304,N_25275);
and U25543 (N_25543,N_25316,N_25363);
xnor U25544 (N_25544,N_25386,N_25353);
xnor U25545 (N_25545,N_25341,N_25305);
nand U25546 (N_25546,N_25272,N_25375);
nand U25547 (N_25547,N_25278,N_25280);
nor U25548 (N_25548,N_25276,N_25268);
or U25549 (N_25549,N_25385,N_25316);
nor U25550 (N_25550,N_25367,N_25255);
nor U25551 (N_25551,N_25274,N_25363);
and U25552 (N_25552,N_25286,N_25234);
and U25553 (N_25553,N_25303,N_25217);
nand U25554 (N_25554,N_25352,N_25222);
xnor U25555 (N_25555,N_25337,N_25231);
or U25556 (N_25556,N_25360,N_25275);
nand U25557 (N_25557,N_25364,N_25312);
or U25558 (N_25558,N_25363,N_25376);
and U25559 (N_25559,N_25237,N_25285);
xnor U25560 (N_25560,N_25362,N_25271);
or U25561 (N_25561,N_25370,N_25260);
nor U25562 (N_25562,N_25254,N_25292);
or U25563 (N_25563,N_25225,N_25364);
or U25564 (N_25564,N_25294,N_25221);
nor U25565 (N_25565,N_25290,N_25382);
or U25566 (N_25566,N_25395,N_25228);
nand U25567 (N_25567,N_25267,N_25372);
nand U25568 (N_25568,N_25262,N_25349);
xnor U25569 (N_25569,N_25345,N_25210);
or U25570 (N_25570,N_25226,N_25262);
or U25571 (N_25571,N_25319,N_25301);
nor U25572 (N_25572,N_25385,N_25220);
xnor U25573 (N_25573,N_25302,N_25274);
and U25574 (N_25574,N_25201,N_25260);
nor U25575 (N_25575,N_25300,N_25215);
or U25576 (N_25576,N_25250,N_25394);
or U25577 (N_25577,N_25389,N_25296);
xor U25578 (N_25578,N_25272,N_25390);
nand U25579 (N_25579,N_25250,N_25334);
xor U25580 (N_25580,N_25219,N_25202);
nand U25581 (N_25581,N_25388,N_25230);
nand U25582 (N_25582,N_25237,N_25345);
nand U25583 (N_25583,N_25235,N_25345);
nor U25584 (N_25584,N_25302,N_25206);
and U25585 (N_25585,N_25287,N_25253);
nor U25586 (N_25586,N_25259,N_25220);
or U25587 (N_25587,N_25258,N_25294);
xnor U25588 (N_25588,N_25244,N_25286);
xnor U25589 (N_25589,N_25396,N_25302);
xnor U25590 (N_25590,N_25310,N_25282);
or U25591 (N_25591,N_25248,N_25275);
or U25592 (N_25592,N_25314,N_25360);
xnor U25593 (N_25593,N_25382,N_25226);
nand U25594 (N_25594,N_25202,N_25266);
xor U25595 (N_25595,N_25359,N_25396);
xnor U25596 (N_25596,N_25317,N_25333);
xor U25597 (N_25597,N_25251,N_25315);
nand U25598 (N_25598,N_25342,N_25293);
xnor U25599 (N_25599,N_25304,N_25289);
nor U25600 (N_25600,N_25505,N_25495);
xor U25601 (N_25601,N_25428,N_25536);
xnor U25602 (N_25602,N_25487,N_25427);
or U25603 (N_25603,N_25527,N_25537);
nand U25604 (N_25604,N_25540,N_25489);
and U25605 (N_25605,N_25504,N_25480);
or U25606 (N_25606,N_25596,N_25564);
xnor U25607 (N_25607,N_25499,N_25508);
nor U25608 (N_25608,N_25409,N_25490);
and U25609 (N_25609,N_25416,N_25454);
xnor U25610 (N_25610,N_25545,N_25436);
nand U25611 (N_25611,N_25519,N_25503);
and U25612 (N_25612,N_25595,N_25535);
or U25613 (N_25613,N_25412,N_25533);
and U25614 (N_25614,N_25463,N_25541);
nor U25615 (N_25615,N_25452,N_25522);
or U25616 (N_25616,N_25547,N_25440);
nor U25617 (N_25617,N_25500,N_25481);
and U25618 (N_25618,N_25478,N_25560);
and U25619 (N_25619,N_25476,N_25462);
and U25620 (N_25620,N_25557,N_25467);
and U25621 (N_25621,N_25403,N_25405);
and U25622 (N_25622,N_25441,N_25474);
nand U25623 (N_25623,N_25431,N_25471);
xnor U25624 (N_25624,N_25599,N_25413);
and U25625 (N_25625,N_25479,N_25584);
or U25626 (N_25626,N_25475,N_25451);
nor U25627 (N_25627,N_25573,N_25552);
xnor U25628 (N_25628,N_25445,N_25432);
xor U25629 (N_25629,N_25528,N_25472);
nand U25630 (N_25630,N_25502,N_25424);
nor U25631 (N_25631,N_25443,N_25497);
xor U25632 (N_25632,N_25469,N_25466);
xor U25633 (N_25633,N_25583,N_25542);
xnor U25634 (N_25634,N_25568,N_25516);
xnor U25635 (N_25635,N_25418,N_25523);
nor U25636 (N_25636,N_25592,N_25470);
nor U25637 (N_25637,N_25585,N_25407);
and U25638 (N_25638,N_25579,N_25422);
and U25639 (N_25639,N_25556,N_25483);
and U25640 (N_25640,N_25498,N_25555);
or U25641 (N_25641,N_25509,N_25526);
or U25642 (N_25642,N_25520,N_25414);
or U25643 (N_25643,N_25465,N_25434);
nor U25644 (N_25644,N_25561,N_25510);
nand U25645 (N_25645,N_25532,N_25529);
nor U25646 (N_25646,N_25587,N_25461);
nor U25647 (N_25647,N_25486,N_25513);
xnor U25648 (N_25648,N_25419,N_25507);
or U25649 (N_25649,N_25586,N_25578);
or U25650 (N_25650,N_25521,N_25459);
nor U25651 (N_25651,N_25446,N_25493);
xor U25652 (N_25652,N_25455,N_25571);
xor U25653 (N_25653,N_25518,N_25566);
xor U25654 (N_25654,N_25442,N_25544);
xor U25655 (N_25655,N_25515,N_25411);
nor U25656 (N_25656,N_25488,N_25400);
and U25657 (N_25657,N_25538,N_25581);
nand U25658 (N_25658,N_25572,N_25525);
nand U25659 (N_25659,N_25570,N_25464);
nand U25660 (N_25660,N_25562,N_25429);
xnor U25661 (N_25661,N_25420,N_25531);
nand U25662 (N_25662,N_25404,N_25491);
nor U25663 (N_25663,N_25577,N_25546);
xor U25664 (N_25664,N_25473,N_25460);
or U25665 (N_25665,N_25551,N_25550);
nor U25666 (N_25666,N_25597,N_25453);
or U25667 (N_25667,N_25468,N_25548);
nand U25668 (N_25668,N_25589,N_25494);
nand U25669 (N_25669,N_25558,N_25482);
and U25670 (N_25670,N_25447,N_25430);
nand U25671 (N_25671,N_25421,N_25458);
nor U25672 (N_25672,N_25524,N_25456);
xor U25673 (N_25673,N_25569,N_25574);
nand U25674 (N_25674,N_25580,N_25444);
nor U25675 (N_25675,N_25539,N_25594);
or U25676 (N_25676,N_25415,N_25433);
or U25677 (N_25677,N_25582,N_25511);
xor U25678 (N_25678,N_25553,N_25588);
and U25679 (N_25679,N_25534,N_25496);
xnor U25680 (N_25680,N_25426,N_25457);
or U25681 (N_25681,N_25449,N_25450);
or U25682 (N_25682,N_25590,N_25417);
or U25683 (N_25683,N_25425,N_25554);
nor U25684 (N_25684,N_25543,N_25565);
and U25685 (N_25685,N_25506,N_25477);
and U25686 (N_25686,N_25406,N_25517);
xnor U25687 (N_25687,N_25501,N_25576);
and U25688 (N_25688,N_25401,N_25485);
xor U25689 (N_25689,N_25438,N_25591);
or U25690 (N_25690,N_25514,N_25549);
nand U25691 (N_25691,N_25410,N_25593);
xor U25692 (N_25692,N_25575,N_25559);
nand U25693 (N_25693,N_25439,N_25563);
or U25694 (N_25694,N_25492,N_25448);
xor U25695 (N_25695,N_25435,N_25512);
nand U25696 (N_25696,N_25484,N_25408);
or U25697 (N_25697,N_25423,N_25530);
or U25698 (N_25698,N_25437,N_25598);
nor U25699 (N_25699,N_25567,N_25402);
or U25700 (N_25700,N_25598,N_25585);
and U25701 (N_25701,N_25423,N_25465);
and U25702 (N_25702,N_25493,N_25406);
nor U25703 (N_25703,N_25465,N_25466);
xor U25704 (N_25704,N_25552,N_25483);
or U25705 (N_25705,N_25431,N_25556);
or U25706 (N_25706,N_25476,N_25441);
and U25707 (N_25707,N_25432,N_25485);
nor U25708 (N_25708,N_25468,N_25414);
xnor U25709 (N_25709,N_25424,N_25513);
nand U25710 (N_25710,N_25544,N_25486);
nor U25711 (N_25711,N_25410,N_25589);
or U25712 (N_25712,N_25435,N_25401);
nor U25713 (N_25713,N_25461,N_25576);
nand U25714 (N_25714,N_25558,N_25551);
nor U25715 (N_25715,N_25451,N_25493);
or U25716 (N_25716,N_25541,N_25429);
nand U25717 (N_25717,N_25407,N_25411);
nor U25718 (N_25718,N_25458,N_25430);
or U25719 (N_25719,N_25537,N_25443);
or U25720 (N_25720,N_25520,N_25411);
nor U25721 (N_25721,N_25519,N_25529);
and U25722 (N_25722,N_25515,N_25475);
nor U25723 (N_25723,N_25516,N_25584);
nor U25724 (N_25724,N_25550,N_25557);
and U25725 (N_25725,N_25556,N_25485);
nor U25726 (N_25726,N_25539,N_25574);
or U25727 (N_25727,N_25579,N_25455);
xor U25728 (N_25728,N_25533,N_25497);
or U25729 (N_25729,N_25464,N_25537);
or U25730 (N_25730,N_25570,N_25489);
xor U25731 (N_25731,N_25449,N_25595);
nor U25732 (N_25732,N_25412,N_25410);
and U25733 (N_25733,N_25496,N_25407);
xor U25734 (N_25734,N_25533,N_25504);
nor U25735 (N_25735,N_25413,N_25596);
and U25736 (N_25736,N_25572,N_25475);
nand U25737 (N_25737,N_25532,N_25442);
and U25738 (N_25738,N_25417,N_25493);
or U25739 (N_25739,N_25419,N_25498);
nand U25740 (N_25740,N_25437,N_25512);
and U25741 (N_25741,N_25570,N_25412);
nor U25742 (N_25742,N_25433,N_25590);
nor U25743 (N_25743,N_25495,N_25468);
nor U25744 (N_25744,N_25401,N_25571);
nand U25745 (N_25745,N_25515,N_25498);
nor U25746 (N_25746,N_25543,N_25439);
nand U25747 (N_25747,N_25530,N_25464);
or U25748 (N_25748,N_25499,N_25552);
nand U25749 (N_25749,N_25509,N_25476);
xor U25750 (N_25750,N_25564,N_25404);
and U25751 (N_25751,N_25455,N_25442);
nor U25752 (N_25752,N_25422,N_25494);
and U25753 (N_25753,N_25543,N_25450);
nor U25754 (N_25754,N_25471,N_25592);
and U25755 (N_25755,N_25420,N_25427);
nor U25756 (N_25756,N_25538,N_25483);
nor U25757 (N_25757,N_25457,N_25536);
xnor U25758 (N_25758,N_25585,N_25489);
xnor U25759 (N_25759,N_25498,N_25597);
nor U25760 (N_25760,N_25525,N_25416);
nand U25761 (N_25761,N_25569,N_25480);
nor U25762 (N_25762,N_25413,N_25567);
nor U25763 (N_25763,N_25444,N_25462);
xor U25764 (N_25764,N_25591,N_25479);
nand U25765 (N_25765,N_25537,N_25515);
and U25766 (N_25766,N_25513,N_25525);
nand U25767 (N_25767,N_25419,N_25582);
or U25768 (N_25768,N_25584,N_25544);
nor U25769 (N_25769,N_25455,N_25430);
or U25770 (N_25770,N_25427,N_25471);
nand U25771 (N_25771,N_25480,N_25527);
nor U25772 (N_25772,N_25470,N_25570);
or U25773 (N_25773,N_25570,N_25427);
xnor U25774 (N_25774,N_25509,N_25555);
xnor U25775 (N_25775,N_25470,N_25447);
nor U25776 (N_25776,N_25469,N_25508);
nor U25777 (N_25777,N_25432,N_25426);
and U25778 (N_25778,N_25498,N_25545);
and U25779 (N_25779,N_25477,N_25511);
or U25780 (N_25780,N_25573,N_25595);
nand U25781 (N_25781,N_25594,N_25508);
or U25782 (N_25782,N_25414,N_25429);
or U25783 (N_25783,N_25596,N_25432);
xor U25784 (N_25784,N_25488,N_25559);
or U25785 (N_25785,N_25593,N_25506);
or U25786 (N_25786,N_25434,N_25534);
nor U25787 (N_25787,N_25434,N_25541);
nand U25788 (N_25788,N_25509,N_25582);
xnor U25789 (N_25789,N_25580,N_25557);
and U25790 (N_25790,N_25485,N_25527);
and U25791 (N_25791,N_25453,N_25437);
xnor U25792 (N_25792,N_25531,N_25472);
xor U25793 (N_25793,N_25468,N_25514);
nand U25794 (N_25794,N_25527,N_25449);
xor U25795 (N_25795,N_25592,N_25466);
xor U25796 (N_25796,N_25476,N_25423);
nand U25797 (N_25797,N_25426,N_25427);
and U25798 (N_25798,N_25452,N_25498);
and U25799 (N_25799,N_25525,N_25586);
nor U25800 (N_25800,N_25769,N_25748);
xnor U25801 (N_25801,N_25799,N_25798);
nand U25802 (N_25802,N_25603,N_25786);
nor U25803 (N_25803,N_25773,N_25790);
xor U25804 (N_25804,N_25725,N_25616);
nor U25805 (N_25805,N_25765,N_25683);
and U25806 (N_25806,N_25779,N_25707);
or U25807 (N_25807,N_25635,N_25699);
or U25808 (N_25808,N_25768,N_25688);
nor U25809 (N_25809,N_25728,N_25702);
nand U25810 (N_25810,N_25690,N_25706);
nand U25811 (N_25811,N_25734,N_25682);
xor U25812 (N_25812,N_25742,N_25747);
and U25813 (N_25813,N_25648,N_25626);
xnor U25814 (N_25814,N_25746,N_25713);
xnor U25815 (N_25815,N_25757,N_25723);
and U25816 (N_25816,N_25697,N_25676);
nor U25817 (N_25817,N_25647,N_25624);
nor U25818 (N_25818,N_25760,N_25633);
and U25819 (N_25819,N_25639,N_25736);
or U25820 (N_25820,N_25774,N_25698);
nand U25821 (N_25821,N_25735,N_25733);
nand U25822 (N_25822,N_25703,N_25659);
nor U25823 (N_25823,N_25792,N_25615);
nor U25824 (N_25824,N_25791,N_25680);
and U25825 (N_25825,N_25672,N_25681);
xor U25826 (N_25826,N_25700,N_25674);
nand U25827 (N_25827,N_25645,N_25623);
nand U25828 (N_25828,N_25695,N_25711);
or U25829 (N_25829,N_25709,N_25715);
nand U25830 (N_25830,N_25718,N_25669);
and U25831 (N_25831,N_25606,N_25777);
nor U25832 (N_25832,N_25617,N_25668);
nor U25833 (N_25833,N_25692,N_25664);
xnor U25834 (N_25834,N_25795,N_25771);
nor U25835 (N_25835,N_25620,N_25727);
nor U25836 (N_25836,N_25696,N_25724);
or U25837 (N_25837,N_25776,N_25694);
xnor U25838 (N_25838,N_25646,N_25675);
or U25839 (N_25839,N_25666,N_25759);
and U25840 (N_25840,N_25766,N_25763);
xor U25841 (N_25841,N_25729,N_25778);
xnor U25842 (N_25842,N_25640,N_25752);
nand U25843 (N_25843,N_25652,N_25601);
nor U25844 (N_25844,N_25783,N_25780);
nand U25845 (N_25845,N_25761,N_25644);
xor U25846 (N_25846,N_25684,N_25632);
nor U25847 (N_25847,N_25641,N_25621);
and U25848 (N_25848,N_25732,N_25726);
or U25849 (N_25849,N_25661,N_25784);
nor U25850 (N_25850,N_25797,N_25653);
or U25851 (N_25851,N_25691,N_25753);
and U25852 (N_25852,N_25751,N_25637);
nand U25853 (N_25853,N_25638,N_25730);
nor U25854 (N_25854,N_25755,N_25610);
xnor U25855 (N_25855,N_25712,N_25628);
or U25856 (N_25856,N_25673,N_25701);
nor U25857 (N_25857,N_25657,N_25739);
nor U25858 (N_25858,N_25775,N_25740);
xnor U25859 (N_25859,N_25785,N_25794);
and U25860 (N_25860,N_25642,N_25649);
and U25861 (N_25861,N_25714,N_25654);
nor U25862 (N_25862,N_25630,N_25720);
and U25863 (N_25863,N_25631,N_25658);
nor U25864 (N_25864,N_25600,N_25722);
xnor U25865 (N_25865,N_25781,N_25744);
nand U25866 (N_25866,N_25665,N_25670);
or U25867 (N_25867,N_25618,N_25741);
or U25868 (N_25868,N_25685,N_25737);
or U25869 (N_25869,N_25710,N_25708);
nand U25870 (N_25870,N_25750,N_25749);
nor U25871 (N_25871,N_25602,N_25619);
nand U25872 (N_25872,N_25756,N_25745);
or U25873 (N_25873,N_25754,N_25796);
nand U25874 (N_25874,N_25655,N_25678);
and U25875 (N_25875,N_25704,N_25625);
or U25876 (N_25876,N_25721,N_25660);
and U25877 (N_25877,N_25716,N_25787);
or U25878 (N_25878,N_25605,N_25738);
nand U25879 (N_25879,N_25650,N_25613);
nand U25880 (N_25880,N_25687,N_25608);
or U25881 (N_25881,N_25671,N_25767);
xnor U25882 (N_25882,N_25743,N_25609);
nor U25883 (N_25883,N_25770,N_25789);
or U25884 (N_25884,N_25636,N_25679);
nor U25885 (N_25885,N_25627,N_25622);
xnor U25886 (N_25886,N_25612,N_25693);
nand U25887 (N_25887,N_25788,N_25764);
or U25888 (N_25888,N_25651,N_25689);
nor U25889 (N_25889,N_25643,N_25686);
nor U25890 (N_25890,N_25793,N_25629);
or U25891 (N_25891,N_25782,N_25667);
and U25892 (N_25892,N_25731,N_25611);
nand U25893 (N_25893,N_25663,N_25607);
and U25894 (N_25894,N_25758,N_25719);
nand U25895 (N_25895,N_25614,N_25662);
or U25896 (N_25896,N_25677,N_25656);
nand U25897 (N_25897,N_25604,N_25705);
and U25898 (N_25898,N_25634,N_25772);
nor U25899 (N_25899,N_25762,N_25717);
and U25900 (N_25900,N_25796,N_25799);
nor U25901 (N_25901,N_25633,N_25663);
and U25902 (N_25902,N_25760,N_25646);
nand U25903 (N_25903,N_25603,N_25772);
nor U25904 (N_25904,N_25671,N_25793);
and U25905 (N_25905,N_25643,N_25754);
nor U25906 (N_25906,N_25766,N_25787);
and U25907 (N_25907,N_25747,N_25620);
nor U25908 (N_25908,N_25704,N_25669);
xor U25909 (N_25909,N_25792,N_25726);
or U25910 (N_25910,N_25745,N_25672);
xor U25911 (N_25911,N_25777,N_25761);
nor U25912 (N_25912,N_25773,N_25664);
xnor U25913 (N_25913,N_25644,N_25607);
or U25914 (N_25914,N_25709,N_25682);
xnor U25915 (N_25915,N_25680,N_25751);
nor U25916 (N_25916,N_25667,N_25687);
xnor U25917 (N_25917,N_25747,N_25739);
or U25918 (N_25918,N_25707,N_25723);
nand U25919 (N_25919,N_25689,N_25742);
and U25920 (N_25920,N_25691,N_25730);
xnor U25921 (N_25921,N_25614,N_25792);
or U25922 (N_25922,N_25638,N_25795);
nand U25923 (N_25923,N_25791,N_25722);
xnor U25924 (N_25924,N_25765,N_25702);
nor U25925 (N_25925,N_25668,N_25630);
or U25926 (N_25926,N_25621,N_25717);
or U25927 (N_25927,N_25775,N_25690);
or U25928 (N_25928,N_25682,N_25601);
and U25929 (N_25929,N_25600,N_25630);
or U25930 (N_25930,N_25641,N_25620);
xor U25931 (N_25931,N_25646,N_25692);
or U25932 (N_25932,N_25662,N_25640);
xor U25933 (N_25933,N_25653,N_25661);
and U25934 (N_25934,N_25777,N_25675);
or U25935 (N_25935,N_25618,N_25693);
nor U25936 (N_25936,N_25726,N_25712);
and U25937 (N_25937,N_25709,N_25723);
or U25938 (N_25938,N_25663,N_25723);
or U25939 (N_25939,N_25690,N_25692);
or U25940 (N_25940,N_25610,N_25752);
and U25941 (N_25941,N_25653,N_25681);
xor U25942 (N_25942,N_25776,N_25601);
nor U25943 (N_25943,N_25729,N_25652);
nor U25944 (N_25944,N_25718,N_25631);
or U25945 (N_25945,N_25641,N_25739);
or U25946 (N_25946,N_25778,N_25765);
or U25947 (N_25947,N_25735,N_25602);
nor U25948 (N_25948,N_25616,N_25788);
xor U25949 (N_25949,N_25674,N_25714);
nor U25950 (N_25950,N_25756,N_25611);
nand U25951 (N_25951,N_25794,N_25687);
xnor U25952 (N_25952,N_25747,N_25657);
and U25953 (N_25953,N_25650,N_25616);
or U25954 (N_25954,N_25637,N_25794);
or U25955 (N_25955,N_25726,N_25624);
and U25956 (N_25956,N_25708,N_25702);
or U25957 (N_25957,N_25624,N_25603);
xnor U25958 (N_25958,N_25617,N_25687);
nor U25959 (N_25959,N_25680,N_25632);
nand U25960 (N_25960,N_25645,N_25664);
or U25961 (N_25961,N_25682,N_25703);
and U25962 (N_25962,N_25670,N_25626);
nor U25963 (N_25963,N_25773,N_25732);
and U25964 (N_25964,N_25639,N_25698);
or U25965 (N_25965,N_25652,N_25728);
xnor U25966 (N_25966,N_25670,N_25730);
xnor U25967 (N_25967,N_25709,N_25787);
xnor U25968 (N_25968,N_25672,N_25720);
nand U25969 (N_25969,N_25777,N_25741);
nor U25970 (N_25970,N_25659,N_25697);
nand U25971 (N_25971,N_25673,N_25671);
or U25972 (N_25972,N_25664,N_25782);
xor U25973 (N_25973,N_25712,N_25757);
and U25974 (N_25974,N_25627,N_25743);
nor U25975 (N_25975,N_25650,N_25776);
and U25976 (N_25976,N_25719,N_25674);
xor U25977 (N_25977,N_25621,N_25682);
or U25978 (N_25978,N_25636,N_25668);
and U25979 (N_25979,N_25671,N_25734);
xnor U25980 (N_25980,N_25754,N_25639);
and U25981 (N_25981,N_25610,N_25726);
or U25982 (N_25982,N_25789,N_25724);
xor U25983 (N_25983,N_25795,N_25716);
xnor U25984 (N_25984,N_25705,N_25688);
and U25985 (N_25985,N_25746,N_25744);
or U25986 (N_25986,N_25706,N_25672);
nor U25987 (N_25987,N_25725,N_25644);
and U25988 (N_25988,N_25672,N_25608);
and U25989 (N_25989,N_25777,N_25794);
xnor U25990 (N_25990,N_25757,N_25651);
or U25991 (N_25991,N_25766,N_25741);
or U25992 (N_25992,N_25703,N_25779);
nor U25993 (N_25993,N_25644,N_25737);
and U25994 (N_25994,N_25659,N_25670);
and U25995 (N_25995,N_25643,N_25791);
xnor U25996 (N_25996,N_25771,N_25720);
nand U25997 (N_25997,N_25776,N_25686);
nor U25998 (N_25998,N_25731,N_25618);
xor U25999 (N_25999,N_25680,N_25709);
nand U26000 (N_26000,N_25888,N_25962);
and U26001 (N_26001,N_25850,N_25947);
nor U26002 (N_26002,N_25907,N_25840);
and U26003 (N_26003,N_25893,N_25940);
or U26004 (N_26004,N_25913,N_25928);
and U26005 (N_26005,N_25939,N_25892);
nand U26006 (N_26006,N_25812,N_25944);
or U26007 (N_26007,N_25848,N_25980);
nor U26008 (N_26008,N_25831,N_25919);
nor U26009 (N_26009,N_25992,N_25955);
xnor U26010 (N_26010,N_25968,N_25924);
xnor U26011 (N_26011,N_25828,N_25846);
nand U26012 (N_26012,N_25881,N_25922);
nor U26013 (N_26013,N_25986,N_25832);
nand U26014 (N_26014,N_25925,N_25958);
or U26015 (N_26015,N_25971,N_25963);
and U26016 (N_26016,N_25884,N_25886);
xnor U26017 (N_26017,N_25960,N_25863);
xor U26018 (N_26018,N_25943,N_25981);
nand U26019 (N_26019,N_25899,N_25987);
nand U26020 (N_26020,N_25949,N_25852);
and U26021 (N_26021,N_25938,N_25844);
nand U26022 (N_26022,N_25900,N_25834);
nor U26023 (N_26023,N_25880,N_25904);
nor U26024 (N_26024,N_25942,N_25821);
xnor U26025 (N_26025,N_25862,N_25946);
xor U26026 (N_26026,N_25923,N_25935);
nor U26027 (N_26027,N_25894,N_25906);
nor U26028 (N_26028,N_25898,N_25809);
or U26029 (N_26029,N_25908,N_25857);
xnor U26030 (N_26030,N_25841,N_25835);
nand U26031 (N_26031,N_25807,N_25895);
nor U26032 (N_26032,N_25909,N_25972);
xor U26033 (N_26033,N_25990,N_25948);
or U26034 (N_26034,N_25825,N_25875);
nor U26035 (N_26035,N_25830,N_25803);
nand U26036 (N_26036,N_25931,N_25956);
nor U26037 (N_26037,N_25811,N_25824);
nand U26038 (N_26038,N_25977,N_25921);
xnor U26039 (N_26039,N_25983,N_25854);
or U26040 (N_26040,N_25842,N_25897);
or U26041 (N_26041,N_25856,N_25820);
and U26042 (N_26042,N_25861,N_25851);
and U26043 (N_26043,N_25966,N_25952);
or U26044 (N_26044,N_25890,N_25896);
nand U26045 (N_26045,N_25975,N_25988);
xnor U26046 (N_26046,N_25813,N_25937);
nand U26047 (N_26047,N_25858,N_25934);
and U26048 (N_26048,N_25871,N_25860);
nor U26049 (N_26049,N_25822,N_25802);
xnor U26050 (N_26050,N_25887,N_25801);
xor U26051 (N_26051,N_25853,N_25866);
xor U26052 (N_26052,N_25878,N_25819);
nor U26053 (N_26053,N_25838,N_25978);
xnor U26054 (N_26054,N_25965,N_25815);
xor U26055 (N_26055,N_25826,N_25999);
nor U26056 (N_26056,N_25976,N_25870);
nand U26057 (N_26057,N_25855,N_25984);
nor U26058 (N_26058,N_25915,N_25874);
nor U26059 (N_26059,N_25941,N_25912);
nor U26060 (N_26060,N_25936,N_25998);
and U26061 (N_26061,N_25927,N_25969);
and U26062 (N_26062,N_25989,N_25910);
or U26063 (N_26063,N_25816,N_25877);
nor U26064 (N_26064,N_25993,N_25905);
nand U26065 (N_26065,N_25979,N_25845);
or U26066 (N_26066,N_25810,N_25885);
nor U26067 (N_26067,N_25843,N_25873);
xor U26068 (N_26068,N_25929,N_25859);
nand U26069 (N_26069,N_25836,N_25997);
nand U26070 (N_26070,N_25953,N_25974);
xor U26071 (N_26071,N_25973,N_25945);
or U26072 (N_26072,N_25982,N_25805);
nor U26073 (N_26073,N_25903,N_25818);
or U26074 (N_26074,N_25957,N_25911);
nand U26075 (N_26075,N_25823,N_25800);
nand U26076 (N_26076,N_25926,N_25901);
and U26077 (N_26077,N_25829,N_25876);
nand U26078 (N_26078,N_25837,N_25964);
and U26079 (N_26079,N_25916,N_25864);
and U26080 (N_26080,N_25920,N_25996);
or U26081 (N_26081,N_25951,N_25932);
and U26082 (N_26082,N_25872,N_25869);
or U26083 (N_26083,N_25847,N_25930);
xor U26084 (N_26084,N_25849,N_25961);
xor U26085 (N_26085,N_25865,N_25994);
nor U26086 (N_26086,N_25950,N_25914);
xnor U26087 (N_26087,N_25879,N_25917);
nand U26088 (N_26088,N_25868,N_25954);
nor U26089 (N_26089,N_25804,N_25833);
or U26090 (N_26090,N_25839,N_25902);
and U26091 (N_26091,N_25806,N_25933);
and U26092 (N_26092,N_25883,N_25891);
and U26093 (N_26093,N_25808,N_25995);
and U26094 (N_26094,N_25889,N_25991);
nand U26095 (N_26095,N_25817,N_25867);
or U26096 (N_26096,N_25814,N_25882);
nor U26097 (N_26097,N_25959,N_25985);
and U26098 (N_26098,N_25967,N_25827);
or U26099 (N_26099,N_25970,N_25918);
nand U26100 (N_26100,N_25875,N_25833);
nand U26101 (N_26101,N_25816,N_25979);
or U26102 (N_26102,N_25892,N_25926);
nand U26103 (N_26103,N_25869,N_25941);
xnor U26104 (N_26104,N_25924,N_25941);
or U26105 (N_26105,N_25859,N_25939);
nand U26106 (N_26106,N_25928,N_25909);
xnor U26107 (N_26107,N_25845,N_25887);
nor U26108 (N_26108,N_25913,N_25948);
nand U26109 (N_26109,N_25924,N_25913);
and U26110 (N_26110,N_25990,N_25823);
xor U26111 (N_26111,N_25999,N_25823);
xor U26112 (N_26112,N_25996,N_25985);
xnor U26113 (N_26113,N_25996,N_25922);
and U26114 (N_26114,N_25882,N_25857);
xnor U26115 (N_26115,N_25817,N_25900);
xor U26116 (N_26116,N_25901,N_25835);
or U26117 (N_26117,N_25831,N_25966);
xor U26118 (N_26118,N_25961,N_25940);
nand U26119 (N_26119,N_25910,N_25942);
and U26120 (N_26120,N_25941,N_25978);
nand U26121 (N_26121,N_25817,N_25829);
xor U26122 (N_26122,N_25951,N_25802);
xor U26123 (N_26123,N_25987,N_25839);
and U26124 (N_26124,N_25968,N_25881);
nand U26125 (N_26125,N_25900,N_25920);
nor U26126 (N_26126,N_25829,N_25894);
nand U26127 (N_26127,N_25912,N_25935);
nor U26128 (N_26128,N_25915,N_25983);
or U26129 (N_26129,N_25820,N_25878);
xnor U26130 (N_26130,N_25866,N_25969);
xor U26131 (N_26131,N_25873,N_25856);
or U26132 (N_26132,N_25854,N_25996);
nor U26133 (N_26133,N_25810,N_25890);
xnor U26134 (N_26134,N_25959,N_25962);
nor U26135 (N_26135,N_25821,N_25866);
and U26136 (N_26136,N_25899,N_25847);
and U26137 (N_26137,N_25953,N_25975);
or U26138 (N_26138,N_25824,N_25909);
nand U26139 (N_26139,N_25862,N_25897);
nor U26140 (N_26140,N_25977,N_25932);
nand U26141 (N_26141,N_25967,N_25918);
and U26142 (N_26142,N_25975,N_25926);
and U26143 (N_26143,N_25996,N_25988);
and U26144 (N_26144,N_25902,N_25817);
nand U26145 (N_26145,N_25864,N_25806);
nand U26146 (N_26146,N_25858,N_25917);
nand U26147 (N_26147,N_25971,N_25923);
xor U26148 (N_26148,N_25897,N_25854);
nor U26149 (N_26149,N_25917,N_25922);
or U26150 (N_26150,N_25822,N_25974);
nor U26151 (N_26151,N_25919,N_25856);
or U26152 (N_26152,N_25853,N_25896);
nor U26153 (N_26153,N_25937,N_25886);
nor U26154 (N_26154,N_25801,N_25880);
and U26155 (N_26155,N_25863,N_25925);
xnor U26156 (N_26156,N_25999,N_25907);
and U26157 (N_26157,N_25999,N_25846);
xor U26158 (N_26158,N_25914,N_25916);
nand U26159 (N_26159,N_25965,N_25824);
nand U26160 (N_26160,N_25995,N_25911);
or U26161 (N_26161,N_25980,N_25859);
nor U26162 (N_26162,N_25971,N_25818);
or U26163 (N_26163,N_25912,N_25909);
and U26164 (N_26164,N_25800,N_25998);
or U26165 (N_26165,N_25858,N_25902);
xor U26166 (N_26166,N_25982,N_25926);
or U26167 (N_26167,N_25849,N_25956);
nand U26168 (N_26168,N_25930,N_25806);
xnor U26169 (N_26169,N_25958,N_25942);
nand U26170 (N_26170,N_25836,N_25865);
nor U26171 (N_26171,N_25871,N_25817);
and U26172 (N_26172,N_25843,N_25951);
and U26173 (N_26173,N_25959,N_25817);
xnor U26174 (N_26174,N_25811,N_25805);
nand U26175 (N_26175,N_25890,N_25889);
or U26176 (N_26176,N_25914,N_25986);
and U26177 (N_26177,N_25938,N_25919);
nor U26178 (N_26178,N_25934,N_25977);
nor U26179 (N_26179,N_25880,N_25919);
nor U26180 (N_26180,N_25879,N_25878);
xor U26181 (N_26181,N_25849,N_25808);
or U26182 (N_26182,N_25974,N_25823);
and U26183 (N_26183,N_25881,N_25843);
and U26184 (N_26184,N_25846,N_25965);
xnor U26185 (N_26185,N_25949,N_25819);
nor U26186 (N_26186,N_25979,N_25873);
nand U26187 (N_26187,N_25921,N_25956);
and U26188 (N_26188,N_25883,N_25913);
nand U26189 (N_26189,N_25826,N_25872);
xor U26190 (N_26190,N_25931,N_25865);
nand U26191 (N_26191,N_25877,N_25997);
nand U26192 (N_26192,N_25915,N_25825);
or U26193 (N_26193,N_25893,N_25994);
and U26194 (N_26194,N_25937,N_25995);
xor U26195 (N_26195,N_25997,N_25917);
nand U26196 (N_26196,N_25876,N_25938);
xor U26197 (N_26197,N_25889,N_25810);
xnor U26198 (N_26198,N_25970,N_25897);
nor U26199 (N_26199,N_25938,N_25966);
and U26200 (N_26200,N_26013,N_26094);
and U26201 (N_26201,N_26102,N_26155);
and U26202 (N_26202,N_26179,N_26165);
nand U26203 (N_26203,N_26105,N_26017);
and U26204 (N_26204,N_26098,N_26198);
nand U26205 (N_26205,N_26116,N_26129);
nand U26206 (N_26206,N_26025,N_26135);
and U26207 (N_26207,N_26036,N_26002);
nand U26208 (N_26208,N_26111,N_26178);
nand U26209 (N_26209,N_26166,N_26056);
or U26210 (N_26210,N_26106,N_26019);
and U26211 (N_26211,N_26124,N_26108);
nand U26212 (N_26212,N_26188,N_26113);
or U26213 (N_26213,N_26031,N_26157);
nand U26214 (N_26214,N_26103,N_26029);
xnor U26215 (N_26215,N_26021,N_26136);
and U26216 (N_26216,N_26080,N_26092);
nor U26217 (N_26217,N_26154,N_26130);
and U26218 (N_26218,N_26189,N_26164);
xor U26219 (N_26219,N_26152,N_26186);
or U26220 (N_26220,N_26060,N_26173);
nand U26221 (N_26221,N_26147,N_26073);
xnor U26222 (N_26222,N_26145,N_26096);
nand U26223 (N_26223,N_26054,N_26159);
nor U26224 (N_26224,N_26127,N_26045);
or U26225 (N_26225,N_26182,N_26168);
xor U26226 (N_26226,N_26091,N_26199);
xor U26227 (N_26227,N_26062,N_26052);
or U26228 (N_26228,N_26187,N_26191);
xnor U26229 (N_26229,N_26089,N_26044);
xor U26230 (N_26230,N_26023,N_26151);
and U26231 (N_26231,N_26140,N_26163);
nand U26232 (N_26232,N_26051,N_26049);
and U26233 (N_26233,N_26082,N_26121);
nor U26234 (N_26234,N_26131,N_26171);
nand U26235 (N_26235,N_26150,N_26067);
xnor U26236 (N_26236,N_26156,N_26195);
xor U26237 (N_26237,N_26088,N_26010);
nand U26238 (N_26238,N_26120,N_26058);
or U26239 (N_26239,N_26185,N_26117);
xnor U26240 (N_26240,N_26181,N_26100);
or U26241 (N_26241,N_26123,N_26196);
nand U26242 (N_26242,N_26132,N_26176);
xor U26243 (N_26243,N_26142,N_26146);
and U26244 (N_26244,N_26072,N_26133);
or U26245 (N_26245,N_26030,N_26055);
xor U26246 (N_26246,N_26001,N_26149);
nor U26247 (N_26247,N_26079,N_26107);
and U26248 (N_26248,N_26034,N_26035);
nor U26249 (N_26249,N_26144,N_26071);
nand U26250 (N_26250,N_26048,N_26183);
and U26251 (N_26251,N_26193,N_26084);
nor U26252 (N_26252,N_26043,N_26046);
xnor U26253 (N_26253,N_26053,N_26125);
nor U26254 (N_26254,N_26172,N_26119);
and U26255 (N_26255,N_26170,N_26077);
and U26256 (N_26256,N_26007,N_26024);
nand U26257 (N_26257,N_26097,N_26038);
and U26258 (N_26258,N_26169,N_26032);
nor U26259 (N_26259,N_26099,N_26190);
xnor U26260 (N_26260,N_26141,N_26042);
and U26261 (N_26261,N_26061,N_26014);
and U26262 (N_26262,N_26095,N_26112);
nand U26263 (N_26263,N_26040,N_26128);
or U26264 (N_26264,N_26011,N_26134);
and U26265 (N_26265,N_26066,N_26109);
nor U26266 (N_26266,N_26167,N_26003);
nor U26267 (N_26267,N_26047,N_26000);
xor U26268 (N_26268,N_26020,N_26118);
nor U26269 (N_26269,N_26086,N_26064);
and U26270 (N_26270,N_26005,N_26085);
and U26271 (N_26271,N_26158,N_26033);
and U26272 (N_26272,N_26162,N_26065);
xnor U26273 (N_26273,N_26153,N_26139);
and U26274 (N_26274,N_26093,N_26039);
and U26275 (N_26275,N_26104,N_26012);
nor U26276 (N_26276,N_26122,N_26160);
nand U26277 (N_26277,N_26197,N_26137);
or U26278 (N_26278,N_26074,N_26114);
xor U26279 (N_26279,N_26018,N_26192);
xor U26280 (N_26280,N_26059,N_26115);
xor U26281 (N_26281,N_26050,N_26028);
nor U26282 (N_26282,N_26177,N_26069);
and U26283 (N_26283,N_26174,N_26083);
and U26284 (N_26284,N_26022,N_26090);
and U26285 (N_26285,N_26075,N_26126);
or U26286 (N_26286,N_26148,N_26087);
nor U26287 (N_26287,N_26194,N_26006);
nand U26288 (N_26288,N_26070,N_26009);
and U26289 (N_26289,N_26008,N_26078);
nor U26290 (N_26290,N_26068,N_26015);
or U26291 (N_26291,N_26027,N_26138);
nor U26292 (N_26292,N_26143,N_26004);
xnor U26293 (N_26293,N_26041,N_26180);
xnor U26294 (N_26294,N_26110,N_26161);
xor U26295 (N_26295,N_26026,N_26016);
or U26296 (N_26296,N_26175,N_26037);
nand U26297 (N_26297,N_26063,N_26057);
nand U26298 (N_26298,N_26076,N_26101);
and U26299 (N_26299,N_26081,N_26184);
or U26300 (N_26300,N_26171,N_26036);
or U26301 (N_26301,N_26171,N_26120);
nand U26302 (N_26302,N_26123,N_26114);
and U26303 (N_26303,N_26049,N_26110);
or U26304 (N_26304,N_26050,N_26043);
xor U26305 (N_26305,N_26021,N_26116);
nor U26306 (N_26306,N_26134,N_26183);
nand U26307 (N_26307,N_26121,N_26193);
nor U26308 (N_26308,N_26172,N_26161);
or U26309 (N_26309,N_26193,N_26013);
nand U26310 (N_26310,N_26012,N_26086);
nor U26311 (N_26311,N_26170,N_26031);
and U26312 (N_26312,N_26046,N_26037);
xor U26313 (N_26313,N_26164,N_26135);
nor U26314 (N_26314,N_26120,N_26156);
nand U26315 (N_26315,N_26010,N_26119);
xor U26316 (N_26316,N_26084,N_26023);
and U26317 (N_26317,N_26182,N_26007);
and U26318 (N_26318,N_26148,N_26053);
nor U26319 (N_26319,N_26185,N_26129);
xnor U26320 (N_26320,N_26162,N_26165);
or U26321 (N_26321,N_26050,N_26081);
xnor U26322 (N_26322,N_26109,N_26177);
and U26323 (N_26323,N_26008,N_26010);
nor U26324 (N_26324,N_26097,N_26134);
nor U26325 (N_26325,N_26163,N_26038);
or U26326 (N_26326,N_26195,N_26137);
nand U26327 (N_26327,N_26106,N_26144);
nor U26328 (N_26328,N_26191,N_26045);
nor U26329 (N_26329,N_26192,N_26094);
xnor U26330 (N_26330,N_26009,N_26180);
and U26331 (N_26331,N_26090,N_26011);
nor U26332 (N_26332,N_26038,N_26103);
and U26333 (N_26333,N_26008,N_26188);
xnor U26334 (N_26334,N_26029,N_26056);
nand U26335 (N_26335,N_26121,N_26153);
or U26336 (N_26336,N_26123,N_26135);
nand U26337 (N_26337,N_26130,N_26007);
and U26338 (N_26338,N_26103,N_26197);
xor U26339 (N_26339,N_26075,N_26073);
nand U26340 (N_26340,N_26196,N_26144);
and U26341 (N_26341,N_26051,N_26010);
or U26342 (N_26342,N_26091,N_26152);
nor U26343 (N_26343,N_26157,N_26020);
or U26344 (N_26344,N_26172,N_26112);
xor U26345 (N_26345,N_26025,N_26157);
nand U26346 (N_26346,N_26010,N_26121);
xnor U26347 (N_26347,N_26189,N_26167);
and U26348 (N_26348,N_26047,N_26113);
xor U26349 (N_26349,N_26154,N_26155);
xnor U26350 (N_26350,N_26103,N_26043);
xnor U26351 (N_26351,N_26137,N_26058);
nor U26352 (N_26352,N_26124,N_26040);
xor U26353 (N_26353,N_26095,N_26174);
or U26354 (N_26354,N_26087,N_26162);
nand U26355 (N_26355,N_26138,N_26049);
nand U26356 (N_26356,N_26167,N_26001);
xnor U26357 (N_26357,N_26084,N_26133);
nor U26358 (N_26358,N_26188,N_26090);
nor U26359 (N_26359,N_26019,N_26149);
or U26360 (N_26360,N_26152,N_26183);
and U26361 (N_26361,N_26157,N_26096);
nor U26362 (N_26362,N_26071,N_26021);
nor U26363 (N_26363,N_26188,N_26103);
or U26364 (N_26364,N_26120,N_26146);
nand U26365 (N_26365,N_26012,N_26151);
xor U26366 (N_26366,N_26182,N_26141);
or U26367 (N_26367,N_26093,N_26163);
and U26368 (N_26368,N_26072,N_26033);
xnor U26369 (N_26369,N_26076,N_26058);
or U26370 (N_26370,N_26085,N_26156);
xnor U26371 (N_26371,N_26102,N_26031);
or U26372 (N_26372,N_26177,N_26102);
xor U26373 (N_26373,N_26086,N_26075);
nand U26374 (N_26374,N_26103,N_26066);
nand U26375 (N_26375,N_26130,N_26097);
and U26376 (N_26376,N_26023,N_26061);
nor U26377 (N_26377,N_26007,N_26132);
or U26378 (N_26378,N_26074,N_26020);
nor U26379 (N_26379,N_26052,N_26053);
or U26380 (N_26380,N_26187,N_26122);
and U26381 (N_26381,N_26021,N_26034);
nor U26382 (N_26382,N_26055,N_26127);
or U26383 (N_26383,N_26192,N_26027);
xnor U26384 (N_26384,N_26155,N_26043);
nor U26385 (N_26385,N_26052,N_26096);
nand U26386 (N_26386,N_26195,N_26104);
xor U26387 (N_26387,N_26179,N_26194);
xnor U26388 (N_26388,N_26124,N_26177);
xor U26389 (N_26389,N_26071,N_26075);
and U26390 (N_26390,N_26191,N_26013);
xnor U26391 (N_26391,N_26004,N_26180);
nor U26392 (N_26392,N_26131,N_26145);
and U26393 (N_26393,N_26195,N_26044);
nand U26394 (N_26394,N_26010,N_26111);
or U26395 (N_26395,N_26115,N_26026);
or U26396 (N_26396,N_26037,N_26106);
xor U26397 (N_26397,N_26022,N_26192);
or U26398 (N_26398,N_26088,N_26043);
or U26399 (N_26399,N_26067,N_26047);
nand U26400 (N_26400,N_26216,N_26300);
nor U26401 (N_26401,N_26323,N_26388);
nor U26402 (N_26402,N_26353,N_26286);
xnor U26403 (N_26403,N_26281,N_26365);
nand U26404 (N_26404,N_26368,N_26253);
or U26405 (N_26405,N_26264,N_26260);
xnor U26406 (N_26406,N_26283,N_26372);
nor U26407 (N_26407,N_26382,N_26312);
xnor U26408 (N_26408,N_26374,N_26200);
nor U26409 (N_26409,N_26322,N_26328);
and U26410 (N_26410,N_26309,N_26239);
nand U26411 (N_26411,N_26303,N_26273);
and U26412 (N_26412,N_26241,N_26232);
nor U26413 (N_26413,N_26222,N_26361);
and U26414 (N_26414,N_26327,N_26261);
xnor U26415 (N_26415,N_26265,N_26363);
nand U26416 (N_26416,N_26201,N_26316);
and U26417 (N_26417,N_26224,N_26396);
nand U26418 (N_26418,N_26331,N_26211);
or U26419 (N_26419,N_26267,N_26231);
and U26420 (N_26420,N_26397,N_26226);
or U26421 (N_26421,N_26377,N_26223);
or U26422 (N_26422,N_26252,N_26367);
and U26423 (N_26423,N_26301,N_26259);
xor U26424 (N_26424,N_26371,N_26330);
xor U26425 (N_26425,N_26317,N_26390);
nand U26426 (N_26426,N_26237,N_26333);
and U26427 (N_26427,N_26255,N_26315);
and U26428 (N_26428,N_26227,N_26369);
nor U26429 (N_26429,N_26215,N_26251);
nand U26430 (N_26430,N_26299,N_26348);
xnor U26431 (N_26431,N_26319,N_26268);
nor U26432 (N_26432,N_26336,N_26393);
nand U26433 (N_26433,N_26359,N_26389);
nand U26434 (N_26434,N_26258,N_26356);
or U26435 (N_26435,N_26357,N_26230);
xnor U26436 (N_26436,N_26362,N_26320);
and U26437 (N_26437,N_26240,N_26249);
or U26438 (N_26438,N_26335,N_26292);
and U26439 (N_26439,N_26288,N_26271);
xnor U26440 (N_26440,N_26314,N_26394);
or U26441 (N_26441,N_26349,N_26272);
or U26442 (N_26442,N_26373,N_26280);
xnor U26443 (N_26443,N_26399,N_26340);
or U26444 (N_26444,N_26246,N_26392);
or U26445 (N_26445,N_26282,N_26234);
nand U26446 (N_26446,N_26269,N_26277);
xor U26447 (N_26447,N_26346,N_26384);
xnor U26448 (N_26448,N_26209,N_26302);
and U26449 (N_26449,N_26360,N_26307);
xnor U26450 (N_26450,N_26318,N_26354);
and U26451 (N_26451,N_26311,N_26257);
nor U26452 (N_26452,N_26380,N_26350);
nand U26453 (N_26453,N_26274,N_26305);
and U26454 (N_26454,N_26262,N_26308);
nor U26455 (N_26455,N_26364,N_26334);
nand U26456 (N_26456,N_26296,N_26376);
xor U26457 (N_26457,N_26342,N_26235);
nand U26458 (N_26458,N_26297,N_26290);
or U26459 (N_26459,N_26366,N_26245);
and U26460 (N_26460,N_26217,N_26387);
xnor U26461 (N_26461,N_26219,N_26338);
nor U26462 (N_26462,N_26236,N_26250);
nor U26463 (N_26463,N_26341,N_26284);
or U26464 (N_26464,N_26210,N_26378);
or U26465 (N_26465,N_26370,N_26293);
nand U26466 (N_26466,N_26381,N_26276);
nand U26467 (N_26467,N_26229,N_26221);
xor U26468 (N_26468,N_26306,N_26298);
nor U26469 (N_26469,N_26332,N_26395);
and U26470 (N_26470,N_26337,N_26206);
nor U26471 (N_26471,N_26385,N_26321);
and U26472 (N_26472,N_26345,N_26285);
xor U26473 (N_26473,N_26352,N_26263);
nand U26474 (N_26474,N_26228,N_26351);
nor U26475 (N_26475,N_26244,N_26202);
and U26476 (N_26476,N_26242,N_26208);
and U26477 (N_26477,N_26238,N_26325);
nand U26478 (N_26478,N_26375,N_26289);
xor U26479 (N_26479,N_26247,N_26324);
nand U26480 (N_26480,N_26339,N_26275);
xor U26481 (N_26481,N_26344,N_26270);
xnor U26482 (N_26482,N_26291,N_26310);
nor U26483 (N_26483,N_26220,N_26207);
nor U26484 (N_26484,N_26266,N_26347);
or U26485 (N_26485,N_26326,N_26218);
or U26486 (N_26486,N_26343,N_26304);
nand U26487 (N_26487,N_26243,N_26358);
and U26488 (N_26488,N_26248,N_26233);
and U26489 (N_26489,N_26386,N_26225);
nand U26490 (N_26490,N_26383,N_26212);
and U26491 (N_26491,N_26391,N_26256);
nor U26492 (N_26492,N_26287,N_26254);
nand U26493 (N_26493,N_26214,N_26205);
nand U26494 (N_26494,N_26379,N_26355);
nor U26495 (N_26495,N_26398,N_26213);
nand U26496 (N_26496,N_26313,N_26204);
xnor U26497 (N_26497,N_26294,N_26329);
or U26498 (N_26498,N_26278,N_26295);
nor U26499 (N_26499,N_26279,N_26203);
xnor U26500 (N_26500,N_26314,N_26233);
xnor U26501 (N_26501,N_26306,N_26360);
and U26502 (N_26502,N_26277,N_26241);
xnor U26503 (N_26503,N_26279,N_26275);
and U26504 (N_26504,N_26207,N_26341);
nor U26505 (N_26505,N_26212,N_26264);
and U26506 (N_26506,N_26321,N_26319);
nand U26507 (N_26507,N_26326,N_26235);
nand U26508 (N_26508,N_26226,N_26246);
or U26509 (N_26509,N_26309,N_26298);
nor U26510 (N_26510,N_26226,N_26256);
nor U26511 (N_26511,N_26309,N_26394);
nor U26512 (N_26512,N_26226,N_26248);
xor U26513 (N_26513,N_26379,N_26350);
and U26514 (N_26514,N_26259,N_26383);
and U26515 (N_26515,N_26221,N_26348);
or U26516 (N_26516,N_26378,N_26249);
and U26517 (N_26517,N_26221,N_26246);
xor U26518 (N_26518,N_26387,N_26397);
nand U26519 (N_26519,N_26369,N_26363);
or U26520 (N_26520,N_26357,N_26388);
nand U26521 (N_26521,N_26372,N_26379);
and U26522 (N_26522,N_26267,N_26331);
nor U26523 (N_26523,N_26303,N_26325);
nand U26524 (N_26524,N_26303,N_26313);
nand U26525 (N_26525,N_26304,N_26253);
nor U26526 (N_26526,N_26208,N_26238);
nand U26527 (N_26527,N_26330,N_26392);
nor U26528 (N_26528,N_26393,N_26254);
and U26529 (N_26529,N_26343,N_26215);
and U26530 (N_26530,N_26302,N_26277);
xor U26531 (N_26531,N_26359,N_26373);
or U26532 (N_26532,N_26211,N_26241);
nor U26533 (N_26533,N_26262,N_26267);
nor U26534 (N_26534,N_26218,N_26354);
nand U26535 (N_26535,N_26365,N_26243);
and U26536 (N_26536,N_26234,N_26244);
or U26537 (N_26537,N_26339,N_26363);
or U26538 (N_26538,N_26317,N_26264);
nor U26539 (N_26539,N_26285,N_26222);
xnor U26540 (N_26540,N_26368,N_26398);
or U26541 (N_26541,N_26319,N_26355);
nand U26542 (N_26542,N_26236,N_26280);
or U26543 (N_26543,N_26306,N_26376);
and U26544 (N_26544,N_26268,N_26385);
or U26545 (N_26545,N_26376,N_26246);
or U26546 (N_26546,N_26259,N_26217);
or U26547 (N_26547,N_26315,N_26276);
and U26548 (N_26548,N_26346,N_26326);
nor U26549 (N_26549,N_26210,N_26350);
nor U26550 (N_26550,N_26332,N_26221);
nor U26551 (N_26551,N_26377,N_26289);
xor U26552 (N_26552,N_26285,N_26239);
nand U26553 (N_26553,N_26206,N_26261);
xnor U26554 (N_26554,N_26367,N_26274);
nor U26555 (N_26555,N_26348,N_26331);
nand U26556 (N_26556,N_26393,N_26200);
nand U26557 (N_26557,N_26296,N_26334);
xor U26558 (N_26558,N_26260,N_26237);
or U26559 (N_26559,N_26394,N_26330);
and U26560 (N_26560,N_26388,N_26352);
nor U26561 (N_26561,N_26234,N_26361);
or U26562 (N_26562,N_26215,N_26292);
nand U26563 (N_26563,N_26268,N_26355);
nor U26564 (N_26564,N_26244,N_26352);
xnor U26565 (N_26565,N_26396,N_26205);
and U26566 (N_26566,N_26255,N_26388);
xnor U26567 (N_26567,N_26372,N_26261);
or U26568 (N_26568,N_26344,N_26315);
nand U26569 (N_26569,N_26267,N_26388);
or U26570 (N_26570,N_26285,N_26261);
xnor U26571 (N_26571,N_26220,N_26359);
and U26572 (N_26572,N_26220,N_26235);
nor U26573 (N_26573,N_26242,N_26341);
nand U26574 (N_26574,N_26247,N_26273);
xnor U26575 (N_26575,N_26238,N_26304);
nor U26576 (N_26576,N_26359,N_26234);
nor U26577 (N_26577,N_26314,N_26345);
nand U26578 (N_26578,N_26247,N_26274);
or U26579 (N_26579,N_26240,N_26311);
and U26580 (N_26580,N_26307,N_26210);
and U26581 (N_26581,N_26332,N_26247);
or U26582 (N_26582,N_26249,N_26372);
and U26583 (N_26583,N_26370,N_26396);
or U26584 (N_26584,N_26230,N_26240);
nor U26585 (N_26585,N_26396,N_26318);
xnor U26586 (N_26586,N_26218,N_26380);
nand U26587 (N_26587,N_26376,N_26297);
xor U26588 (N_26588,N_26357,N_26223);
nand U26589 (N_26589,N_26297,N_26315);
or U26590 (N_26590,N_26372,N_26216);
nand U26591 (N_26591,N_26398,N_26384);
xnor U26592 (N_26592,N_26203,N_26234);
or U26593 (N_26593,N_26244,N_26347);
nor U26594 (N_26594,N_26312,N_26213);
or U26595 (N_26595,N_26334,N_26317);
or U26596 (N_26596,N_26246,N_26264);
and U26597 (N_26597,N_26388,N_26280);
nor U26598 (N_26598,N_26397,N_26239);
nand U26599 (N_26599,N_26279,N_26316);
and U26600 (N_26600,N_26571,N_26411);
and U26601 (N_26601,N_26503,N_26500);
and U26602 (N_26602,N_26446,N_26496);
nor U26603 (N_26603,N_26516,N_26450);
nor U26604 (N_26604,N_26572,N_26524);
or U26605 (N_26605,N_26580,N_26559);
nand U26606 (N_26606,N_26465,N_26471);
nor U26607 (N_26607,N_26528,N_26579);
or U26608 (N_26608,N_26475,N_26593);
xor U26609 (N_26609,N_26456,N_26412);
xnor U26610 (N_26610,N_26551,N_26512);
xor U26611 (N_26611,N_26509,N_26440);
nand U26612 (N_26612,N_26462,N_26419);
xnor U26613 (N_26613,N_26598,N_26532);
nand U26614 (N_26614,N_26545,N_26511);
or U26615 (N_26615,N_26531,N_26549);
and U26616 (N_26616,N_26562,N_26480);
or U26617 (N_26617,N_26569,N_26555);
or U26618 (N_26618,N_26515,N_26560);
or U26619 (N_26619,N_26510,N_26589);
nor U26620 (N_26620,N_26498,N_26402);
or U26621 (N_26621,N_26526,N_26586);
or U26622 (N_26622,N_26430,N_26433);
xnor U26623 (N_26623,N_26418,N_26595);
nand U26624 (N_26624,N_26408,N_26557);
xor U26625 (N_26625,N_26507,N_26492);
and U26626 (N_26626,N_26468,N_26493);
xor U26627 (N_26627,N_26548,N_26485);
and U26628 (N_26628,N_26484,N_26592);
nor U26629 (N_26629,N_26550,N_26570);
nor U26630 (N_26630,N_26554,N_26467);
and U26631 (N_26631,N_26466,N_26442);
or U26632 (N_26632,N_26596,N_26414);
nand U26633 (N_26633,N_26438,N_26536);
or U26634 (N_26634,N_26499,N_26444);
nand U26635 (N_26635,N_26481,N_26424);
xnor U26636 (N_26636,N_26537,N_26514);
xor U26637 (N_26637,N_26472,N_26504);
or U26638 (N_26638,N_26533,N_26530);
or U26639 (N_26639,N_26425,N_26461);
nor U26640 (N_26640,N_26590,N_26587);
nand U26641 (N_26641,N_26435,N_26487);
or U26642 (N_26642,N_26522,N_26473);
or U26643 (N_26643,N_26458,N_26495);
xor U26644 (N_26644,N_26575,N_26553);
xor U26645 (N_26645,N_26523,N_26561);
xor U26646 (N_26646,N_26483,N_26409);
and U26647 (N_26647,N_26547,N_26567);
and U26648 (N_26648,N_26420,N_26599);
nand U26649 (N_26649,N_26489,N_26581);
xor U26650 (N_26650,N_26427,N_26459);
xnor U26651 (N_26651,N_26460,N_26543);
nand U26652 (N_26652,N_26422,N_26470);
xnor U26653 (N_26653,N_26431,N_26474);
xnor U26654 (N_26654,N_26404,N_26464);
nor U26655 (N_26655,N_26454,N_26502);
xnor U26656 (N_26656,N_26513,N_26568);
xor U26657 (N_26657,N_26573,N_26546);
or U26658 (N_26658,N_26416,N_26479);
or U26659 (N_26659,N_26541,N_26517);
or U26660 (N_26660,N_26584,N_26539);
nor U26661 (N_26661,N_26577,N_26476);
xnor U26662 (N_26662,N_26413,N_26558);
or U26663 (N_26663,N_26400,N_26439);
or U26664 (N_26664,N_26597,N_26486);
nor U26665 (N_26665,N_26451,N_26437);
xnor U26666 (N_26666,N_26565,N_26574);
nor U26667 (N_26667,N_26552,N_26428);
and U26668 (N_26668,N_26529,N_26519);
or U26669 (N_26669,N_26429,N_26525);
nor U26670 (N_26670,N_26491,N_26407);
nor U26671 (N_26671,N_26564,N_26477);
nor U26672 (N_26672,N_26453,N_26578);
nor U26673 (N_26673,N_26585,N_26521);
xor U26674 (N_26674,N_26576,N_26406);
or U26675 (N_26675,N_26520,N_26455);
and U26676 (N_26676,N_26482,N_26506);
xnor U26677 (N_26677,N_26591,N_26463);
and U26678 (N_26678,N_26497,N_26423);
nand U26679 (N_26679,N_26566,N_26544);
or U26680 (N_26680,N_26441,N_26556);
xnor U26681 (N_26681,N_26436,N_26449);
xnor U26682 (N_26682,N_26563,N_26421);
xnor U26683 (N_26683,N_26594,N_26505);
nand U26684 (N_26684,N_26494,N_26445);
nor U26685 (N_26685,N_26405,N_26583);
nand U26686 (N_26686,N_26434,N_26403);
or U26687 (N_26687,N_26518,N_26582);
xnor U26688 (N_26688,N_26501,N_26448);
nand U26689 (N_26689,N_26415,N_26469);
and U26690 (N_26690,N_26417,N_26527);
nor U26691 (N_26691,N_26540,N_26432);
xnor U26692 (N_26692,N_26478,N_26508);
and U26693 (N_26693,N_26410,N_26401);
xnor U26694 (N_26694,N_26443,N_26588);
nand U26695 (N_26695,N_26457,N_26542);
nand U26696 (N_26696,N_26490,N_26452);
or U26697 (N_26697,N_26426,N_26447);
or U26698 (N_26698,N_26488,N_26535);
and U26699 (N_26699,N_26538,N_26534);
or U26700 (N_26700,N_26511,N_26495);
xnor U26701 (N_26701,N_26427,N_26519);
or U26702 (N_26702,N_26439,N_26489);
nand U26703 (N_26703,N_26510,N_26502);
or U26704 (N_26704,N_26546,N_26525);
nand U26705 (N_26705,N_26504,N_26573);
or U26706 (N_26706,N_26526,N_26599);
xnor U26707 (N_26707,N_26518,N_26592);
and U26708 (N_26708,N_26523,N_26428);
nor U26709 (N_26709,N_26488,N_26456);
and U26710 (N_26710,N_26472,N_26441);
nand U26711 (N_26711,N_26543,N_26428);
nand U26712 (N_26712,N_26528,N_26566);
xor U26713 (N_26713,N_26478,N_26520);
or U26714 (N_26714,N_26431,N_26430);
or U26715 (N_26715,N_26423,N_26590);
and U26716 (N_26716,N_26455,N_26435);
and U26717 (N_26717,N_26525,N_26473);
nor U26718 (N_26718,N_26456,N_26424);
nand U26719 (N_26719,N_26444,N_26500);
or U26720 (N_26720,N_26499,N_26419);
nor U26721 (N_26721,N_26582,N_26492);
and U26722 (N_26722,N_26578,N_26564);
or U26723 (N_26723,N_26412,N_26574);
xnor U26724 (N_26724,N_26530,N_26495);
nand U26725 (N_26725,N_26545,N_26469);
nand U26726 (N_26726,N_26535,N_26539);
or U26727 (N_26727,N_26532,N_26497);
or U26728 (N_26728,N_26522,N_26520);
or U26729 (N_26729,N_26554,N_26447);
or U26730 (N_26730,N_26425,N_26498);
xor U26731 (N_26731,N_26502,N_26574);
xnor U26732 (N_26732,N_26566,N_26575);
nand U26733 (N_26733,N_26596,N_26599);
xor U26734 (N_26734,N_26514,N_26564);
and U26735 (N_26735,N_26477,N_26595);
nor U26736 (N_26736,N_26428,N_26569);
nand U26737 (N_26737,N_26524,N_26589);
xnor U26738 (N_26738,N_26552,N_26493);
xnor U26739 (N_26739,N_26421,N_26577);
or U26740 (N_26740,N_26482,N_26435);
nand U26741 (N_26741,N_26539,N_26543);
nor U26742 (N_26742,N_26542,N_26408);
nor U26743 (N_26743,N_26469,N_26450);
or U26744 (N_26744,N_26519,N_26470);
nand U26745 (N_26745,N_26412,N_26478);
nand U26746 (N_26746,N_26464,N_26456);
and U26747 (N_26747,N_26478,N_26455);
xor U26748 (N_26748,N_26441,N_26589);
xnor U26749 (N_26749,N_26561,N_26450);
and U26750 (N_26750,N_26538,N_26576);
and U26751 (N_26751,N_26568,N_26510);
nand U26752 (N_26752,N_26582,N_26425);
and U26753 (N_26753,N_26549,N_26595);
or U26754 (N_26754,N_26422,N_26400);
nor U26755 (N_26755,N_26414,N_26498);
xnor U26756 (N_26756,N_26408,N_26434);
nor U26757 (N_26757,N_26585,N_26542);
nor U26758 (N_26758,N_26599,N_26460);
xnor U26759 (N_26759,N_26496,N_26423);
or U26760 (N_26760,N_26510,N_26410);
and U26761 (N_26761,N_26463,N_26507);
nand U26762 (N_26762,N_26420,N_26558);
nor U26763 (N_26763,N_26508,N_26443);
or U26764 (N_26764,N_26441,N_26563);
xnor U26765 (N_26765,N_26422,N_26460);
or U26766 (N_26766,N_26555,N_26540);
nand U26767 (N_26767,N_26452,N_26466);
or U26768 (N_26768,N_26598,N_26408);
and U26769 (N_26769,N_26569,N_26496);
and U26770 (N_26770,N_26452,N_26511);
or U26771 (N_26771,N_26594,N_26565);
or U26772 (N_26772,N_26542,N_26528);
nand U26773 (N_26773,N_26510,N_26421);
nor U26774 (N_26774,N_26458,N_26426);
or U26775 (N_26775,N_26565,N_26527);
nand U26776 (N_26776,N_26500,N_26533);
and U26777 (N_26777,N_26441,N_26560);
or U26778 (N_26778,N_26549,N_26426);
and U26779 (N_26779,N_26570,N_26599);
and U26780 (N_26780,N_26489,N_26543);
and U26781 (N_26781,N_26553,N_26455);
nor U26782 (N_26782,N_26589,N_26514);
nor U26783 (N_26783,N_26425,N_26411);
nand U26784 (N_26784,N_26450,N_26458);
nor U26785 (N_26785,N_26534,N_26537);
nand U26786 (N_26786,N_26571,N_26580);
xor U26787 (N_26787,N_26472,N_26409);
and U26788 (N_26788,N_26452,N_26460);
or U26789 (N_26789,N_26411,N_26466);
nor U26790 (N_26790,N_26492,N_26490);
and U26791 (N_26791,N_26572,N_26448);
xor U26792 (N_26792,N_26551,N_26403);
nor U26793 (N_26793,N_26502,N_26538);
xnor U26794 (N_26794,N_26550,N_26481);
nor U26795 (N_26795,N_26475,N_26583);
nor U26796 (N_26796,N_26524,N_26442);
nand U26797 (N_26797,N_26556,N_26471);
nor U26798 (N_26798,N_26460,N_26583);
nor U26799 (N_26799,N_26544,N_26486);
and U26800 (N_26800,N_26627,N_26755);
xnor U26801 (N_26801,N_26645,N_26653);
or U26802 (N_26802,N_26779,N_26658);
nor U26803 (N_26803,N_26763,N_26778);
nor U26804 (N_26804,N_26785,N_26744);
xnor U26805 (N_26805,N_26752,N_26776);
xnor U26806 (N_26806,N_26650,N_26663);
nand U26807 (N_26807,N_26718,N_26758);
nand U26808 (N_26808,N_26739,N_26713);
xnor U26809 (N_26809,N_26679,N_26680);
or U26810 (N_26810,N_26724,N_26742);
nor U26811 (N_26811,N_26764,N_26635);
nand U26812 (N_26812,N_26659,N_26794);
nor U26813 (N_26813,N_26719,N_26600);
nor U26814 (N_26814,N_26722,N_26604);
nand U26815 (N_26815,N_26672,N_26620);
nand U26816 (N_26816,N_26691,N_26687);
and U26817 (N_26817,N_26768,N_26716);
nand U26818 (N_26818,N_26648,N_26607);
nand U26819 (N_26819,N_26662,N_26669);
or U26820 (N_26820,N_26692,N_26732);
xor U26821 (N_26821,N_26685,N_26619);
and U26822 (N_26822,N_26723,N_26655);
and U26823 (N_26823,N_26780,N_26786);
xnor U26824 (N_26824,N_26652,N_26668);
nor U26825 (N_26825,N_26751,N_26769);
nand U26826 (N_26826,N_26753,N_26711);
nand U26827 (N_26827,N_26788,N_26613);
nand U26828 (N_26828,N_26651,N_26703);
nand U26829 (N_26829,N_26731,N_26702);
and U26830 (N_26830,N_26757,N_26606);
and U26831 (N_26831,N_26643,N_26735);
xor U26832 (N_26832,N_26701,N_26721);
nand U26833 (N_26833,N_26693,N_26792);
and U26834 (N_26834,N_26700,N_26644);
xor U26835 (N_26835,N_26623,N_26773);
and U26836 (N_26836,N_26725,N_26690);
nand U26837 (N_26837,N_26682,N_26730);
nor U26838 (N_26838,N_26720,N_26614);
nor U26839 (N_26839,N_26664,N_26689);
nand U26840 (N_26840,N_26781,N_26748);
nand U26841 (N_26841,N_26697,N_26640);
nor U26842 (N_26842,N_26741,N_26631);
nor U26843 (N_26843,N_26617,N_26601);
nand U26844 (N_26844,N_26775,N_26667);
xor U26845 (N_26845,N_26630,N_26746);
xor U26846 (N_26846,N_26777,N_26639);
or U26847 (N_26847,N_26634,N_26770);
nor U26848 (N_26848,N_26743,N_26622);
or U26849 (N_26849,N_26710,N_26675);
or U26850 (N_26850,N_26698,N_26608);
nor U26851 (N_26851,N_26628,N_26671);
and U26852 (N_26852,N_26784,N_26745);
nor U26853 (N_26853,N_26616,N_26656);
nand U26854 (N_26854,N_26765,N_26626);
xor U26855 (N_26855,N_26712,N_26766);
or U26856 (N_26856,N_26760,N_26674);
nor U26857 (N_26857,N_26795,N_26704);
nor U26858 (N_26858,N_26734,N_26797);
and U26859 (N_26859,N_26611,N_26705);
nand U26860 (N_26860,N_26615,N_26633);
nand U26861 (N_26861,N_26796,N_26688);
nor U26862 (N_26862,N_26750,N_26609);
and U26863 (N_26863,N_26625,N_26787);
nor U26864 (N_26864,N_26673,N_26657);
nand U26865 (N_26865,N_26738,N_26605);
or U26866 (N_26866,N_26684,N_26762);
nor U26867 (N_26867,N_26660,N_26676);
nor U26868 (N_26868,N_26761,N_26798);
nand U26869 (N_26869,N_26799,N_26726);
or U26870 (N_26870,N_26636,N_26632);
xnor U26871 (N_26871,N_26666,N_26646);
xnor U26872 (N_26872,N_26772,N_26681);
or U26873 (N_26873,N_26696,N_26733);
and U26874 (N_26874,N_26677,N_26654);
nor U26875 (N_26875,N_26694,N_26740);
and U26876 (N_26876,N_26717,N_26642);
xor U26877 (N_26877,N_26665,N_26649);
nor U26878 (N_26878,N_26624,N_26759);
or U26879 (N_26879,N_26737,N_26728);
and U26880 (N_26880,N_26603,N_26791);
or U26881 (N_26881,N_26638,N_26621);
nor U26882 (N_26882,N_26729,N_26783);
and U26883 (N_26883,N_26683,N_26709);
or U26884 (N_26884,N_26686,N_26637);
and U26885 (N_26885,N_26610,N_26747);
nor U26886 (N_26886,N_26793,N_26708);
nand U26887 (N_26887,N_26782,N_26789);
nor U26888 (N_26888,N_26699,N_26727);
nand U26889 (N_26889,N_26661,N_26771);
nor U26890 (N_26890,N_26641,N_26647);
or U26891 (N_26891,N_26678,N_26790);
or U26892 (N_26892,N_26714,N_26774);
nor U26893 (N_26893,N_26754,N_26756);
or U26894 (N_26894,N_26618,N_26749);
or U26895 (N_26895,N_26767,N_26715);
nand U26896 (N_26896,N_26707,N_26695);
nand U26897 (N_26897,N_26629,N_26602);
nor U26898 (N_26898,N_26736,N_26612);
nand U26899 (N_26899,N_26670,N_26706);
nor U26900 (N_26900,N_26798,N_26707);
or U26901 (N_26901,N_26763,N_26720);
nor U26902 (N_26902,N_26774,N_26612);
and U26903 (N_26903,N_26610,N_26681);
and U26904 (N_26904,N_26748,N_26789);
or U26905 (N_26905,N_26762,N_26604);
or U26906 (N_26906,N_26605,N_26622);
nand U26907 (N_26907,N_26736,N_26678);
nor U26908 (N_26908,N_26796,N_26719);
nand U26909 (N_26909,N_26728,N_26640);
nor U26910 (N_26910,N_26776,N_26789);
nand U26911 (N_26911,N_26664,N_26654);
xor U26912 (N_26912,N_26680,N_26606);
and U26913 (N_26913,N_26676,N_26712);
nor U26914 (N_26914,N_26633,N_26765);
and U26915 (N_26915,N_26710,N_26696);
xor U26916 (N_26916,N_26743,N_26678);
nor U26917 (N_26917,N_26716,N_26668);
or U26918 (N_26918,N_26601,N_26727);
xnor U26919 (N_26919,N_26745,N_26638);
and U26920 (N_26920,N_26710,N_26712);
nor U26921 (N_26921,N_26662,N_26674);
or U26922 (N_26922,N_26606,N_26746);
xnor U26923 (N_26923,N_26792,N_26728);
nand U26924 (N_26924,N_26649,N_26707);
or U26925 (N_26925,N_26655,N_26743);
and U26926 (N_26926,N_26749,N_26716);
xnor U26927 (N_26927,N_26753,N_26771);
nand U26928 (N_26928,N_26742,N_26745);
nor U26929 (N_26929,N_26785,N_26762);
or U26930 (N_26930,N_26773,N_26739);
or U26931 (N_26931,N_26631,N_26674);
xnor U26932 (N_26932,N_26747,N_26795);
nor U26933 (N_26933,N_26646,N_26702);
or U26934 (N_26934,N_26690,N_26674);
or U26935 (N_26935,N_26663,N_26641);
or U26936 (N_26936,N_26672,N_26717);
or U26937 (N_26937,N_26669,N_26645);
xor U26938 (N_26938,N_26672,N_26782);
or U26939 (N_26939,N_26695,N_26679);
xnor U26940 (N_26940,N_26740,N_26646);
and U26941 (N_26941,N_26724,N_26670);
xor U26942 (N_26942,N_26678,N_26676);
nand U26943 (N_26943,N_26782,N_26662);
or U26944 (N_26944,N_26702,N_26732);
or U26945 (N_26945,N_26753,N_26700);
nor U26946 (N_26946,N_26750,N_26786);
or U26947 (N_26947,N_26771,N_26721);
or U26948 (N_26948,N_26678,N_26711);
and U26949 (N_26949,N_26628,N_26673);
and U26950 (N_26950,N_26734,N_26768);
or U26951 (N_26951,N_26754,N_26788);
xor U26952 (N_26952,N_26737,N_26676);
xnor U26953 (N_26953,N_26704,N_26784);
or U26954 (N_26954,N_26669,N_26647);
nand U26955 (N_26955,N_26686,N_26782);
nor U26956 (N_26956,N_26768,N_26697);
and U26957 (N_26957,N_26615,N_26649);
and U26958 (N_26958,N_26717,N_26675);
xnor U26959 (N_26959,N_26632,N_26621);
and U26960 (N_26960,N_26797,N_26714);
xnor U26961 (N_26961,N_26648,N_26778);
or U26962 (N_26962,N_26743,N_26617);
and U26963 (N_26963,N_26774,N_26747);
xor U26964 (N_26964,N_26713,N_26634);
or U26965 (N_26965,N_26769,N_26685);
and U26966 (N_26966,N_26659,N_26633);
nor U26967 (N_26967,N_26735,N_26603);
xor U26968 (N_26968,N_26745,N_26611);
xor U26969 (N_26969,N_26724,N_26702);
and U26970 (N_26970,N_26681,N_26709);
or U26971 (N_26971,N_26711,N_26658);
nor U26972 (N_26972,N_26609,N_26698);
xor U26973 (N_26973,N_26663,N_26798);
and U26974 (N_26974,N_26637,N_26638);
nand U26975 (N_26975,N_26737,N_26708);
xnor U26976 (N_26976,N_26744,N_26745);
nand U26977 (N_26977,N_26625,N_26668);
nand U26978 (N_26978,N_26757,N_26774);
or U26979 (N_26979,N_26742,N_26645);
xnor U26980 (N_26980,N_26641,N_26776);
nor U26981 (N_26981,N_26699,N_26760);
and U26982 (N_26982,N_26648,N_26721);
or U26983 (N_26983,N_26768,N_26753);
and U26984 (N_26984,N_26606,N_26631);
nor U26985 (N_26985,N_26630,N_26673);
and U26986 (N_26986,N_26609,N_26717);
or U26987 (N_26987,N_26681,N_26790);
nor U26988 (N_26988,N_26713,N_26699);
and U26989 (N_26989,N_26746,N_26749);
and U26990 (N_26990,N_26717,N_26632);
or U26991 (N_26991,N_26642,N_26729);
and U26992 (N_26992,N_26726,N_26736);
nand U26993 (N_26993,N_26743,N_26639);
or U26994 (N_26994,N_26604,N_26763);
and U26995 (N_26995,N_26779,N_26626);
or U26996 (N_26996,N_26715,N_26658);
xnor U26997 (N_26997,N_26773,N_26747);
or U26998 (N_26998,N_26729,N_26782);
xor U26999 (N_26999,N_26734,N_26670);
xor U27000 (N_27000,N_26822,N_26826);
nor U27001 (N_27001,N_26889,N_26868);
and U27002 (N_27002,N_26871,N_26817);
and U27003 (N_27003,N_26959,N_26840);
xor U27004 (N_27004,N_26916,N_26965);
xnor U27005 (N_27005,N_26980,N_26851);
nand U27006 (N_27006,N_26897,N_26816);
nor U27007 (N_27007,N_26932,N_26973);
and U27008 (N_27008,N_26934,N_26859);
xor U27009 (N_27009,N_26903,N_26946);
xnor U27010 (N_27010,N_26907,N_26865);
xor U27011 (N_27011,N_26918,N_26929);
nor U27012 (N_27012,N_26983,N_26823);
xor U27013 (N_27013,N_26938,N_26812);
or U27014 (N_27014,N_26847,N_26874);
nor U27015 (N_27015,N_26839,N_26952);
and U27016 (N_27016,N_26977,N_26923);
or U27017 (N_27017,N_26811,N_26920);
and U27018 (N_27018,N_26935,N_26971);
nor U27019 (N_27019,N_26872,N_26902);
xnor U27020 (N_27020,N_26953,N_26901);
xor U27021 (N_27021,N_26854,N_26915);
nor U27022 (N_27022,N_26857,N_26877);
or U27023 (N_27023,N_26995,N_26849);
nand U27024 (N_27024,N_26895,N_26866);
and U27025 (N_27025,N_26886,N_26821);
xnor U27026 (N_27026,N_26986,N_26982);
nand U27027 (N_27027,N_26800,N_26917);
xnor U27028 (N_27028,N_26900,N_26969);
nor U27029 (N_27029,N_26820,N_26996);
nor U27030 (N_27030,N_26803,N_26848);
nor U27031 (N_27031,N_26975,N_26926);
nor U27032 (N_27032,N_26940,N_26884);
nand U27033 (N_27033,N_26984,N_26968);
nor U27034 (N_27034,N_26955,N_26908);
xor U27035 (N_27035,N_26972,N_26813);
xor U27036 (N_27036,N_26939,N_26924);
nand U27037 (N_27037,N_26862,N_26948);
nand U27038 (N_27038,N_26852,N_26802);
nand U27039 (N_27039,N_26861,N_26819);
or U27040 (N_27040,N_26994,N_26890);
and U27041 (N_27041,N_26801,N_26957);
xor U27042 (N_27042,N_26882,N_26958);
or U27043 (N_27043,N_26873,N_26841);
nand U27044 (N_27044,N_26843,N_26818);
or U27045 (N_27045,N_26928,N_26807);
nand U27046 (N_27046,N_26899,N_26838);
or U27047 (N_27047,N_26936,N_26846);
xor U27048 (N_27048,N_26943,N_26999);
nor U27049 (N_27049,N_26963,N_26964);
nor U27050 (N_27050,N_26837,N_26950);
and U27051 (N_27051,N_26863,N_26990);
or U27052 (N_27052,N_26885,N_26855);
and U27053 (N_27053,N_26869,N_26978);
xor U27054 (N_27054,N_26896,N_26876);
nand U27055 (N_27055,N_26875,N_26893);
or U27056 (N_27056,N_26814,N_26836);
nor U27057 (N_27057,N_26824,N_26830);
nor U27058 (N_27058,N_26880,N_26911);
nand U27059 (N_27059,N_26805,N_26887);
nor U27060 (N_27060,N_26891,N_26954);
or U27061 (N_27061,N_26992,N_26806);
and U27062 (N_27062,N_26914,N_26961);
nor U27063 (N_27063,N_26867,N_26927);
nand U27064 (N_27064,N_26991,N_26864);
xnor U27065 (N_27065,N_26832,N_26998);
nor U27066 (N_27066,N_26850,N_26881);
or U27067 (N_27067,N_26937,N_26829);
xnor U27068 (N_27068,N_26878,N_26898);
nor U27069 (N_27069,N_26921,N_26949);
nor U27070 (N_27070,N_26944,N_26989);
nor U27071 (N_27071,N_26808,N_26960);
xnor U27072 (N_27072,N_26967,N_26997);
nand U27073 (N_27073,N_26844,N_26906);
xor U27074 (N_27074,N_26945,N_26834);
xnor U27075 (N_27075,N_26804,N_26856);
xnor U27076 (N_27076,N_26845,N_26835);
nor U27077 (N_27077,N_26933,N_26904);
nand U27078 (N_27078,N_26905,N_26912);
or U27079 (N_27079,N_26827,N_26947);
nand U27080 (N_27080,N_26951,N_26879);
nor U27081 (N_27081,N_26925,N_26825);
xnor U27082 (N_27082,N_26888,N_26853);
nor U27083 (N_27083,N_26942,N_26985);
nor U27084 (N_27084,N_26919,N_26883);
nor U27085 (N_27085,N_26988,N_26860);
nand U27086 (N_27086,N_26993,N_26833);
nand U27087 (N_27087,N_26970,N_26894);
nor U27088 (N_27088,N_26987,N_26956);
xor U27089 (N_27089,N_26931,N_26892);
nand U27090 (N_27090,N_26909,N_26870);
nand U27091 (N_27091,N_26966,N_26810);
nor U27092 (N_27092,N_26831,N_26922);
nor U27093 (N_27093,N_26842,N_26962);
and U27094 (N_27094,N_26979,N_26910);
xnor U27095 (N_27095,N_26981,N_26815);
and U27096 (N_27096,N_26974,N_26913);
nand U27097 (N_27097,N_26976,N_26941);
nor U27098 (N_27098,N_26858,N_26828);
xor U27099 (N_27099,N_26930,N_26809);
xnor U27100 (N_27100,N_26815,N_26881);
and U27101 (N_27101,N_26979,N_26805);
and U27102 (N_27102,N_26851,N_26983);
and U27103 (N_27103,N_26890,N_26820);
xor U27104 (N_27104,N_26906,N_26867);
nand U27105 (N_27105,N_26896,N_26915);
xnor U27106 (N_27106,N_26833,N_26810);
and U27107 (N_27107,N_26966,N_26954);
nor U27108 (N_27108,N_26862,N_26866);
xnor U27109 (N_27109,N_26845,N_26970);
and U27110 (N_27110,N_26871,N_26998);
and U27111 (N_27111,N_26926,N_26883);
nor U27112 (N_27112,N_26810,N_26977);
or U27113 (N_27113,N_26988,N_26867);
nor U27114 (N_27114,N_26921,N_26826);
xor U27115 (N_27115,N_26941,N_26849);
nor U27116 (N_27116,N_26894,N_26857);
xor U27117 (N_27117,N_26842,N_26938);
nand U27118 (N_27118,N_26988,N_26876);
nand U27119 (N_27119,N_26960,N_26893);
nand U27120 (N_27120,N_26923,N_26974);
and U27121 (N_27121,N_26869,N_26938);
nor U27122 (N_27122,N_26949,N_26837);
nor U27123 (N_27123,N_26998,N_26924);
and U27124 (N_27124,N_26816,N_26808);
or U27125 (N_27125,N_26844,N_26924);
nand U27126 (N_27126,N_26904,N_26870);
and U27127 (N_27127,N_26929,N_26953);
nor U27128 (N_27128,N_26836,N_26801);
nor U27129 (N_27129,N_26866,N_26947);
and U27130 (N_27130,N_26875,N_26890);
nand U27131 (N_27131,N_26880,N_26863);
and U27132 (N_27132,N_26999,N_26885);
nor U27133 (N_27133,N_26920,N_26837);
nand U27134 (N_27134,N_26841,N_26944);
and U27135 (N_27135,N_26944,N_26894);
nand U27136 (N_27136,N_26877,N_26945);
nor U27137 (N_27137,N_26833,N_26965);
xor U27138 (N_27138,N_26973,N_26906);
nor U27139 (N_27139,N_26871,N_26891);
and U27140 (N_27140,N_26802,N_26903);
nor U27141 (N_27141,N_26846,N_26969);
xnor U27142 (N_27142,N_26856,N_26848);
xnor U27143 (N_27143,N_26890,N_26872);
and U27144 (N_27144,N_26835,N_26979);
or U27145 (N_27145,N_26922,N_26930);
xnor U27146 (N_27146,N_26817,N_26836);
and U27147 (N_27147,N_26831,N_26891);
xor U27148 (N_27148,N_26860,N_26809);
xnor U27149 (N_27149,N_26845,N_26884);
nor U27150 (N_27150,N_26807,N_26809);
xnor U27151 (N_27151,N_26985,N_26913);
xor U27152 (N_27152,N_26912,N_26814);
nand U27153 (N_27153,N_26831,N_26954);
nand U27154 (N_27154,N_26850,N_26989);
nand U27155 (N_27155,N_26903,N_26996);
and U27156 (N_27156,N_26994,N_26882);
and U27157 (N_27157,N_26864,N_26921);
nor U27158 (N_27158,N_26815,N_26911);
nand U27159 (N_27159,N_26997,N_26800);
nand U27160 (N_27160,N_26963,N_26959);
and U27161 (N_27161,N_26958,N_26828);
xor U27162 (N_27162,N_26919,N_26903);
and U27163 (N_27163,N_26958,N_26836);
nand U27164 (N_27164,N_26863,N_26925);
and U27165 (N_27165,N_26803,N_26947);
nand U27166 (N_27166,N_26830,N_26973);
nor U27167 (N_27167,N_26963,N_26836);
xnor U27168 (N_27168,N_26976,N_26905);
nand U27169 (N_27169,N_26985,N_26823);
nor U27170 (N_27170,N_26912,N_26931);
nand U27171 (N_27171,N_26801,N_26993);
xnor U27172 (N_27172,N_26953,N_26911);
and U27173 (N_27173,N_26964,N_26918);
xor U27174 (N_27174,N_26847,N_26815);
nor U27175 (N_27175,N_26823,N_26861);
xor U27176 (N_27176,N_26892,N_26842);
xnor U27177 (N_27177,N_26932,N_26979);
xor U27178 (N_27178,N_26980,N_26855);
nor U27179 (N_27179,N_26965,N_26828);
nor U27180 (N_27180,N_26901,N_26984);
nor U27181 (N_27181,N_26960,N_26901);
and U27182 (N_27182,N_26849,N_26842);
or U27183 (N_27183,N_26927,N_26805);
nand U27184 (N_27184,N_26917,N_26825);
or U27185 (N_27185,N_26868,N_26963);
nor U27186 (N_27186,N_26917,N_26935);
and U27187 (N_27187,N_26952,N_26982);
xnor U27188 (N_27188,N_26842,N_26826);
xor U27189 (N_27189,N_26938,N_26890);
nor U27190 (N_27190,N_26979,N_26885);
or U27191 (N_27191,N_26914,N_26811);
or U27192 (N_27192,N_26880,N_26852);
nor U27193 (N_27193,N_26932,N_26878);
nand U27194 (N_27194,N_26957,N_26914);
or U27195 (N_27195,N_26953,N_26862);
or U27196 (N_27196,N_26955,N_26926);
and U27197 (N_27197,N_26851,N_26947);
nand U27198 (N_27198,N_26847,N_26977);
and U27199 (N_27199,N_26961,N_26991);
nor U27200 (N_27200,N_27022,N_27128);
nor U27201 (N_27201,N_27151,N_27092);
nor U27202 (N_27202,N_27167,N_27169);
xor U27203 (N_27203,N_27061,N_27197);
or U27204 (N_27204,N_27107,N_27080);
or U27205 (N_27205,N_27194,N_27133);
or U27206 (N_27206,N_27196,N_27135);
xnor U27207 (N_27207,N_27104,N_27020);
xnor U27208 (N_27208,N_27030,N_27038);
or U27209 (N_27209,N_27003,N_27053);
or U27210 (N_27210,N_27097,N_27012);
xnor U27211 (N_27211,N_27102,N_27117);
or U27212 (N_27212,N_27199,N_27016);
nand U27213 (N_27213,N_27142,N_27183);
nor U27214 (N_27214,N_27024,N_27172);
nand U27215 (N_27215,N_27126,N_27192);
or U27216 (N_27216,N_27051,N_27068);
nor U27217 (N_27217,N_27120,N_27028);
nor U27218 (N_27218,N_27087,N_27059);
and U27219 (N_27219,N_27094,N_27138);
xnor U27220 (N_27220,N_27180,N_27041);
xnor U27221 (N_27221,N_27074,N_27177);
and U27222 (N_27222,N_27039,N_27116);
nor U27223 (N_27223,N_27156,N_27014);
nand U27224 (N_27224,N_27084,N_27069);
xnor U27225 (N_27225,N_27027,N_27054);
nor U27226 (N_27226,N_27029,N_27137);
nand U27227 (N_27227,N_27155,N_27079);
nor U27228 (N_27228,N_27110,N_27179);
or U27229 (N_27229,N_27032,N_27103);
nand U27230 (N_27230,N_27000,N_27129);
xnor U27231 (N_27231,N_27066,N_27047);
xor U27232 (N_27232,N_27122,N_27037);
nand U27233 (N_27233,N_27021,N_27001);
or U27234 (N_27234,N_27096,N_27191);
nor U27235 (N_27235,N_27072,N_27046);
xor U27236 (N_27236,N_27174,N_27050);
nand U27237 (N_27237,N_27176,N_27064);
and U27238 (N_27238,N_27056,N_27026);
or U27239 (N_27239,N_27140,N_27111);
nand U27240 (N_27240,N_27168,N_27090);
nor U27241 (N_27241,N_27034,N_27067);
nor U27242 (N_27242,N_27171,N_27076);
and U27243 (N_27243,N_27058,N_27152);
nor U27244 (N_27244,N_27143,N_27006);
or U27245 (N_27245,N_27189,N_27081);
nor U27246 (N_27246,N_27109,N_27184);
and U27247 (N_27247,N_27091,N_27100);
nor U27248 (N_27248,N_27086,N_27164);
nand U27249 (N_27249,N_27132,N_27009);
xnor U27250 (N_27250,N_27130,N_27190);
nor U27251 (N_27251,N_27042,N_27139);
nor U27252 (N_27252,N_27101,N_27013);
nor U27253 (N_27253,N_27134,N_27125);
xnor U27254 (N_27254,N_27002,N_27017);
nand U27255 (N_27255,N_27075,N_27188);
xnor U27256 (N_27256,N_27055,N_27088);
or U27257 (N_27257,N_27112,N_27023);
or U27258 (N_27258,N_27173,N_27153);
nor U27259 (N_27259,N_27011,N_27186);
or U27260 (N_27260,N_27078,N_27162);
xnor U27261 (N_27261,N_27052,N_27063);
nand U27262 (N_27262,N_27070,N_27115);
and U27263 (N_27263,N_27114,N_27145);
and U27264 (N_27264,N_27044,N_27165);
xnor U27265 (N_27265,N_27118,N_27040);
and U27266 (N_27266,N_27144,N_27163);
and U27267 (N_27267,N_27045,N_27121);
or U27268 (N_27268,N_27105,N_27010);
and U27269 (N_27269,N_27182,N_27060);
or U27270 (N_27270,N_27178,N_27095);
nor U27271 (N_27271,N_27057,N_27147);
or U27272 (N_27272,N_27043,N_27181);
and U27273 (N_27273,N_27099,N_27158);
or U27274 (N_27274,N_27015,N_27157);
or U27275 (N_27275,N_27004,N_27089);
xnor U27276 (N_27276,N_27035,N_27093);
nor U27277 (N_27277,N_27085,N_27019);
nor U27278 (N_27278,N_27036,N_27166);
nor U27279 (N_27279,N_27175,N_27187);
nor U27280 (N_27280,N_27170,N_27154);
and U27281 (N_27281,N_27033,N_27025);
or U27282 (N_27282,N_27127,N_27106);
nor U27283 (N_27283,N_27031,N_27071);
and U27284 (N_27284,N_27005,N_27098);
and U27285 (N_27285,N_27065,N_27161);
nand U27286 (N_27286,N_27150,N_27124);
nand U27287 (N_27287,N_27073,N_27008);
nor U27288 (N_27288,N_27062,N_27148);
nor U27289 (N_27289,N_27149,N_27131);
or U27290 (N_27290,N_27193,N_27185);
and U27291 (N_27291,N_27146,N_27141);
and U27292 (N_27292,N_27113,N_27159);
or U27293 (N_27293,N_27119,N_27136);
or U27294 (N_27294,N_27108,N_27123);
xor U27295 (N_27295,N_27018,N_27083);
xor U27296 (N_27296,N_27160,N_27049);
nand U27297 (N_27297,N_27198,N_27077);
xor U27298 (N_27298,N_27048,N_27195);
nand U27299 (N_27299,N_27082,N_27007);
xnor U27300 (N_27300,N_27141,N_27001);
nand U27301 (N_27301,N_27165,N_27069);
and U27302 (N_27302,N_27166,N_27136);
and U27303 (N_27303,N_27122,N_27008);
nand U27304 (N_27304,N_27086,N_27120);
or U27305 (N_27305,N_27196,N_27091);
nand U27306 (N_27306,N_27069,N_27009);
xor U27307 (N_27307,N_27079,N_27151);
nand U27308 (N_27308,N_27189,N_27050);
and U27309 (N_27309,N_27072,N_27097);
or U27310 (N_27310,N_27071,N_27157);
and U27311 (N_27311,N_27198,N_27048);
or U27312 (N_27312,N_27029,N_27000);
nor U27313 (N_27313,N_27039,N_27127);
nand U27314 (N_27314,N_27159,N_27154);
or U27315 (N_27315,N_27022,N_27017);
or U27316 (N_27316,N_27053,N_27022);
nor U27317 (N_27317,N_27180,N_27141);
xnor U27318 (N_27318,N_27191,N_27082);
xor U27319 (N_27319,N_27070,N_27028);
and U27320 (N_27320,N_27086,N_27146);
or U27321 (N_27321,N_27107,N_27198);
nor U27322 (N_27322,N_27023,N_27026);
and U27323 (N_27323,N_27118,N_27137);
nand U27324 (N_27324,N_27005,N_27022);
and U27325 (N_27325,N_27038,N_27059);
and U27326 (N_27326,N_27018,N_27161);
nand U27327 (N_27327,N_27164,N_27144);
and U27328 (N_27328,N_27092,N_27112);
and U27329 (N_27329,N_27030,N_27173);
or U27330 (N_27330,N_27020,N_27184);
xor U27331 (N_27331,N_27157,N_27167);
and U27332 (N_27332,N_27059,N_27179);
xnor U27333 (N_27333,N_27079,N_27017);
and U27334 (N_27334,N_27120,N_27169);
and U27335 (N_27335,N_27035,N_27004);
nand U27336 (N_27336,N_27077,N_27134);
and U27337 (N_27337,N_27057,N_27042);
nand U27338 (N_27338,N_27188,N_27074);
xnor U27339 (N_27339,N_27161,N_27035);
nor U27340 (N_27340,N_27006,N_27044);
and U27341 (N_27341,N_27008,N_27059);
xnor U27342 (N_27342,N_27121,N_27017);
nand U27343 (N_27343,N_27195,N_27102);
xor U27344 (N_27344,N_27073,N_27117);
or U27345 (N_27345,N_27067,N_27065);
nor U27346 (N_27346,N_27043,N_27158);
and U27347 (N_27347,N_27002,N_27013);
nor U27348 (N_27348,N_27141,N_27078);
and U27349 (N_27349,N_27159,N_27186);
or U27350 (N_27350,N_27169,N_27139);
xnor U27351 (N_27351,N_27091,N_27006);
xor U27352 (N_27352,N_27064,N_27011);
and U27353 (N_27353,N_27135,N_27187);
or U27354 (N_27354,N_27101,N_27128);
or U27355 (N_27355,N_27137,N_27183);
and U27356 (N_27356,N_27124,N_27079);
nand U27357 (N_27357,N_27090,N_27156);
and U27358 (N_27358,N_27015,N_27082);
or U27359 (N_27359,N_27180,N_27039);
or U27360 (N_27360,N_27121,N_27006);
xnor U27361 (N_27361,N_27173,N_27062);
xor U27362 (N_27362,N_27032,N_27078);
nor U27363 (N_27363,N_27032,N_27147);
and U27364 (N_27364,N_27148,N_27023);
or U27365 (N_27365,N_27003,N_27034);
nor U27366 (N_27366,N_27023,N_27047);
or U27367 (N_27367,N_27127,N_27176);
nand U27368 (N_27368,N_27138,N_27028);
nor U27369 (N_27369,N_27127,N_27167);
xnor U27370 (N_27370,N_27131,N_27094);
nor U27371 (N_27371,N_27010,N_27071);
and U27372 (N_27372,N_27091,N_27020);
nand U27373 (N_27373,N_27180,N_27059);
nand U27374 (N_27374,N_27082,N_27127);
and U27375 (N_27375,N_27060,N_27123);
or U27376 (N_27376,N_27117,N_27190);
or U27377 (N_27377,N_27139,N_27125);
or U27378 (N_27378,N_27105,N_27159);
nor U27379 (N_27379,N_27139,N_27003);
xor U27380 (N_27380,N_27145,N_27146);
nand U27381 (N_27381,N_27086,N_27123);
xnor U27382 (N_27382,N_27002,N_27056);
xor U27383 (N_27383,N_27122,N_27004);
nand U27384 (N_27384,N_27144,N_27107);
nand U27385 (N_27385,N_27060,N_27002);
nor U27386 (N_27386,N_27131,N_27044);
nor U27387 (N_27387,N_27008,N_27141);
nand U27388 (N_27388,N_27073,N_27063);
nand U27389 (N_27389,N_27074,N_27009);
or U27390 (N_27390,N_27091,N_27176);
or U27391 (N_27391,N_27109,N_27046);
and U27392 (N_27392,N_27084,N_27159);
nand U27393 (N_27393,N_27126,N_27173);
xnor U27394 (N_27394,N_27109,N_27089);
nor U27395 (N_27395,N_27067,N_27195);
and U27396 (N_27396,N_27156,N_27020);
nor U27397 (N_27397,N_27094,N_27179);
xnor U27398 (N_27398,N_27010,N_27129);
nor U27399 (N_27399,N_27199,N_27157);
or U27400 (N_27400,N_27248,N_27285);
xnor U27401 (N_27401,N_27364,N_27326);
xnor U27402 (N_27402,N_27276,N_27322);
xnor U27403 (N_27403,N_27339,N_27396);
or U27404 (N_27404,N_27218,N_27342);
or U27405 (N_27405,N_27266,N_27347);
nand U27406 (N_27406,N_27205,N_27201);
nor U27407 (N_27407,N_27354,N_27331);
or U27408 (N_27408,N_27295,N_27301);
xnor U27409 (N_27409,N_27319,N_27255);
nor U27410 (N_27410,N_27258,N_27320);
or U27411 (N_27411,N_27346,N_27333);
and U27412 (N_27412,N_27225,N_27351);
or U27413 (N_27413,N_27374,N_27361);
or U27414 (N_27414,N_27227,N_27239);
and U27415 (N_27415,N_27274,N_27304);
or U27416 (N_27416,N_27352,N_27307);
xnor U27417 (N_27417,N_27337,N_27233);
xnor U27418 (N_27418,N_27311,N_27338);
nor U27419 (N_27419,N_27355,N_27244);
xor U27420 (N_27420,N_27300,N_27267);
or U27421 (N_27421,N_27395,N_27213);
and U27422 (N_27422,N_27341,N_27343);
nor U27423 (N_27423,N_27393,N_27321);
or U27424 (N_27424,N_27348,N_27232);
nor U27425 (N_27425,N_27282,N_27387);
or U27426 (N_27426,N_27256,N_27373);
or U27427 (N_27427,N_27357,N_27297);
nand U27428 (N_27428,N_27356,N_27215);
and U27429 (N_27429,N_27280,N_27249);
and U27430 (N_27430,N_27221,N_27236);
nand U27431 (N_27431,N_27240,N_27262);
and U27432 (N_27432,N_27241,N_27340);
or U27433 (N_27433,N_27305,N_27330);
xnor U27434 (N_27434,N_27214,N_27345);
or U27435 (N_27435,N_27389,N_27370);
nand U27436 (N_27436,N_27223,N_27367);
or U27437 (N_27437,N_27378,N_27308);
xnor U27438 (N_27438,N_27278,N_27335);
and U27439 (N_27439,N_27230,N_27277);
and U27440 (N_27440,N_27380,N_27224);
xnor U27441 (N_27441,N_27220,N_27287);
nor U27442 (N_27442,N_27344,N_27360);
and U27443 (N_27443,N_27273,N_27349);
nor U27444 (N_27444,N_27254,N_27327);
and U27445 (N_27445,N_27366,N_27303);
or U27446 (N_27446,N_27288,N_27313);
xnor U27447 (N_27447,N_27328,N_27394);
xnor U27448 (N_27448,N_27231,N_27271);
nand U27449 (N_27449,N_27290,N_27376);
and U27450 (N_27450,N_27245,N_27226);
nor U27451 (N_27451,N_27358,N_27250);
or U27452 (N_27452,N_27203,N_27207);
nand U27453 (N_27453,N_27261,N_27210);
nand U27454 (N_27454,N_27264,N_27242);
or U27455 (N_27455,N_27329,N_27291);
xnor U27456 (N_27456,N_27292,N_27238);
nor U27457 (N_27457,N_27353,N_27257);
and U27458 (N_27458,N_27222,N_27229);
xor U27459 (N_27459,N_27211,N_27212);
nor U27460 (N_27460,N_27279,N_27252);
and U27461 (N_27461,N_27316,N_27293);
xor U27462 (N_27462,N_27296,N_27369);
and U27463 (N_27463,N_27235,N_27315);
nand U27464 (N_27464,N_27383,N_27391);
nand U27465 (N_27465,N_27397,N_27314);
and U27466 (N_27466,N_27398,N_27318);
or U27467 (N_27467,N_27390,N_27332);
and U27468 (N_27468,N_27251,N_27372);
nor U27469 (N_27469,N_27382,N_27268);
or U27470 (N_27470,N_27200,N_27334);
nor U27471 (N_27471,N_27260,N_27371);
nand U27472 (N_27472,N_27272,N_27263);
nand U27473 (N_27473,N_27265,N_27312);
xor U27474 (N_27474,N_27325,N_27298);
and U27475 (N_27475,N_27243,N_27234);
and U27476 (N_27476,N_27377,N_27247);
or U27477 (N_27477,N_27310,N_27359);
or U27478 (N_27478,N_27237,N_27379);
nand U27479 (N_27479,N_27368,N_27317);
nand U27480 (N_27480,N_27365,N_27362);
nand U27481 (N_27481,N_27309,N_27208);
nand U27482 (N_27482,N_27375,N_27219);
and U27483 (N_27483,N_27270,N_27385);
nor U27484 (N_27484,N_27284,N_27209);
and U27485 (N_27485,N_27399,N_27283);
or U27486 (N_27486,N_27294,N_27386);
or U27487 (N_27487,N_27202,N_27281);
or U27488 (N_27488,N_27206,N_27381);
and U27489 (N_27489,N_27269,N_27350);
and U27490 (N_27490,N_27286,N_27204);
xor U27491 (N_27491,N_27306,N_27363);
xnor U27492 (N_27492,N_27302,N_27289);
or U27493 (N_27493,N_27275,N_27392);
and U27494 (N_27494,N_27384,N_27246);
and U27495 (N_27495,N_27299,N_27324);
nor U27496 (N_27496,N_27216,N_27253);
xnor U27497 (N_27497,N_27228,N_27217);
nand U27498 (N_27498,N_27388,N_27259);
and U27499 (N_27499,N_27336,N_27323);
and U27500 (N_27500,N_27272,N_27274);
xor U27501 (N_27501,N_27269,N_27218);
and U27502 (N_27502,N_27322,N_27254);
nand U27503 (N_27503,N_27353,N_27232);
nand U27504 (N_27504,N_27366,N_27358);
xor U27505 (N_27505,N_27326,N_27323);
nand U27506 (N_27506,N_27220,N_27214);
or U27507 (N_27507,N_27348,N_27316);
and U27508 (N_27508,N_27223,N_27369);
xor U27509 (N_27509,N_27280,N_27370);
or U27510 (N_27510,N_27281,N_27209);
and U27511 (N_27511,N_27394,N_27370);
nor U27512 (N_27512,N_27399,N_27239);
nand U27513 (N_27513,N_27397,N_27293);
or U27514 (N_27514,N_27337,N_27323);
nor U27515 (N_27515,N_27394,N_27288);
xnor U27516 (N_27516,N_27244,N_27256);
nand U27517 (N_27517,N_27355,N_27347);
nor U27518 (N_27518,N_27300,N_27256);
or U27519 (N_27519,N_27398,N_27284);
nor U27520 (N_27520,N_27358,N_27293);
nor U27521 (N_27521,N_27255,N_27398);
nor U27522 (N_27522,N_27216,N_27213);
nand U27523 (N_27523,N_27299,N_27230);
nor U27524 (N_27524,N_27272,N_27365);
nor U27525 (N_27525,N_27360,N_27365);
nand U27526 (N_27526,N_27276,N_27311);
nand U27527 (N_27527,N_27295,N_27338);
nand U27528 (N_27528,N_27226,N_27301);
and U27529 (N_27529,N_27211,N_27392);
or U27530 (N_27530,N_27261,N_27355);
and U27531 (N_27531,N_27324,N_27218);
nand U27532 (N_27532,N_27379,N_27291);
and U27533 (N_27533,N_27306,N_27320);
nand U27534 (N_27534,N_27346,N_27293);
nand U27535 (N_27535,N_27250,N_27285);
or U27536 (N_27536,N_27335,N_27399);
nor U27537 (N_27537,N_27261,N_27378);
or U27538 (N_27538,N_27230,N_27375);
xnor U27539 (N_27539,N_27202,N_27359);
xnor U27540 (N_27540,N_27292,N_27291);
and U27541 (N_27541,N_27270,N_27368);
or U27542 (N_27542,N_27226,N_27326);
xor U27543 (N_27543,N_27321,N_27303);
nand U27544 (N_27544,N_27335,N_27223);
xnor U27545 (N_27545,N_27236,N_27377);
nor U27546 (N_27546,N_27237,N_27271);
and U27547 (N_27547,N_27235,N_27273);
nor U27548 (N_27548,N_27333,N_27362);
xnor U27549 (N_27549,N_27216,N_27281);
nand U27550 (N_27550,N_27341,N_27317);
or U27551 (N_27551,N_27306,N_27315);
or U27552 (N_27552,N_27295,N_27312);
xnor U27553 (N_27553,N_27343,N_27377);
nor U27554 (N_27554,N_27269,N_27259);
or U27555 (N_27555,N_27340,N_27234);
nor U27556 (N_27556,N_27268,N_27248);
or U27557 (N_27557,N_27361,N_27363);
and U27558 (N_27558,N_27383,N_27366);
and U27559 (N_27559,N_27273,N_27293);
xor U27560 (N_27560,N_27336,N_27260);
nand U27561 (N_27561,N_27292,N_27398);
and U27562 (N_27562,N_27203,N_27232);
xor U27563 (N_27563,N_27378,N_27223);
nor U27564 (N_27564,N_27245,N_27319);
xor U27565 (N_27565,N_27326,N_27390);
or U27566 (N_27566,N_27359,N_27305);
or U27567 (N_27567,N_27208,N_27294);
nor U27568 (N_27568,N_27368,N_27369);
or U27569 (N_27569,N_27271,N_27225);
or U27570 (N_27570,N_27317,N_27320);
nor U27571 (N_27571,N_27255,N_27301);
xor U27572 (N_27572,N_27350,N_27323);
nor U27573 (N_27573,N_27398,N_27231);
nand U27574 (N_27574,N_27237,N_27376);
or U27575 (N_27575,N_27226,N_27224);
and U27576 (N_27576,N_27224,N_27373);
and U27577 (N_27577,N_27386,N_27205);
nor U27578 (N_27578,N_27278,N_27230);
and U27579 (N_27579,N_27362,N_27320);
and U27580 (N_27580,N_27308,N_27223);
xnor U27581 (N_27581,N_27304,N_27212);
nand U27582 (N_27582,N_27208,N_27269);
nand U27583 (N_27583,N_27330,N_27341);
nor U27584 (N_27584,N_27220,N_27325);
nand U27585 (N_27585,N_27321,N_27345);
and U27586 (N_27586,N_27224,N_27269);
nand U27587 (N_27587,N_27357,N_27347);
nor U27588 (N_27588,N_27312,N_27228);
or U27589 (N_27589,N_27283,N_27346);
xnor U27590 (N_27590,N_27358,N_27261);
xnor U27591 (N_27591,N_27361,N_27367);
nand U27592 (N_27592,N_27297,N_27343);
nand U27593 (N_27593,N_27261,N_27335);
and U27594 (N_27594,N_27259,N_27283);
nor U27595 (N_27595,N_27209,N_27237);
or U27596 (N_27596,N_27354,N_27219);
or U27597 (N_27597,N_27348,N_27388);
nand U27598 (N_27598,N_27360,N_27315);
nand U27599 (N_27599,N_27224,N_27352);
and U27600 (N_27600,N_27410,N_27579);
nand U27601 (N_27601,N_27571,N_27439);
nand U27602 (N_27602,N_27400,N_27426);
xor U27603 (N_27603,N_27429,N_27585);
nor U27604 (N_27604,N_27447,N_27436);
nor U27605 (N_27605,N_27463,N_27591);
nand U27606 (N_27606,N_27493,N_27432);
nor U27607 (N_27607,N_27531,N_27525);
nor U27608 (N_27608,N_27510,N_27547);
or U27609 (N_27609,N_27478,N_27402);
or U27610 (N_27610,N_27504,N_27552);
or U27611 (N_27611,N_27580,N_27454);
and U27612 (N_27612,N_27409,N_27536);
xnor U27613 (N_27613,N_27405,N_27545);
nor U27614 (N_27614,N_27456,N_27496);
xor U27615 (N_27615,N_27475,N_27526);
nand U27616 (N_27616,N_27584,N_27520);
nand U27617 (N_27617,N_27502,N_27407);
and U27618 (N_27618,N_27430,N_27530);
xnor U27619 (N_27619,N_27557,N_27467);
nand U27620 (N_27620,N_27458,N_27418);
nand U27621 (N_27621,N_27550,N_27509);
or U27622 (N_27622,N_27434,N_27574);
nor U27623 (N_27623,N_27566,N_27414);
or U27624 (N_27624,N_27421,N_27570);
nor U27625 (N_27625,N_27578,N_27543);
xor U27626 (N_27626,N_27482,N_27450);
or U27627 (N_27627,N_27512,N_27551);
xor U27628 (N_27628,N_27565,N_27464);
xor U27629 (N_27629,N_27466,N_27457);
nand U27630 (N_27630,N_27495,N_27440);
and U27631 (N_27631,N_27535,N_27537);
nor U27632 (N_27632,N_27597,N_27437);
or U27633 (N_27633,N_27592,N_27511);
xor U27634 (N_27634,N_27553,N_27415);
or U27635 (N_27635,N_27499,N_27517);
nand U27636 (N_27636,N_27522,N_27538);
nand U27637 (N_27637,N_27427,N_27423);
nand U27638 (N_27638,N_27455,N_27523);
nand U27639 (N_27639,N_27483,N_27404);
and U27640 (N_27640,N_27424,N_27575);
and U27641 (N_27641,N_27472,N_27459);
or U27642 (N_27642,N_27542,N_27486);
nor U27643 (N_27643,N_27559,N_27420);
xor U27644 (N_27644,N_27446,N_27441);
nand U27645 (N_27645,N_27480,N_27546);
xnor U27646 (N_27646,N_27471,N_27507);
xor U27647 (N_27647,N_27521,N_27503);
and U27648 (N_27648,N_27411,N_27481);
nand U27649 (N_27649,N_27563,N_27422);
nor U27650 (N_27650,N_27595,N_27473);
nor U27651 (N_27651,N_27470,N_27445);
xnor U27652 (N_27652,N_27583,N_27569);
xor U27653 (N_27653,N_27449,N_27462);
xor U27654 (N_27654,N_27492,N_27577);
nand U27655 (N_27655,N_27528,N_27489);
nor U27656 (N_27656,N_27541,N_27479);
nand U27657 (N_27657,N_27556,N_27460);
or U27658 (N_27658,N_27514,N_27469);
nand U27659 (N_27659,N_27539,N_27431);
nor U27660 (N_27660,N_27555,N_27527);
and U27661 (N_27661,N_27506,N_27451);
or U27662 (N_27662,N_27501,N_27582);
nand U27663 (N_27663,N_27533,N_27477);
and U27664 (N_27664,N_27453,N_27428);
and U27665 (N_27665,N_27588,N_27476);
nand U27666 (N_27666,N_27433,N_27573);
and U27667 (N_27667,N_27488,N_27491);
and U27668 (N_27668,N_27474,N_27549);
nand U27669 (N_27669,N_27544,N_27465);
nor U27670 (N_27670,N_27419,N_27442);
and U27671 (N_27671,N_27508,N_27438);
or U27672 (N_27672,N_27417,N_27505);
xor U27673 (N_27673,N_27534,N_27576);
nand U27674 (N_27674,N_27452,N_27529);
xor U27675 (N_27675,N_27598,N_27444);
xor U27676 (N_27676,N_27562,N_27401);
xor U27677 (N_27677,N_27443,N_27567);
or U27678 (N_27678,N_27558,N_27518);
or U27679 (N_27679,N_27524,N_27435);
xor U27680 (N_27680,N_27568,N_27516);
nand U27681 (N_27681,N_27572,N_27515);
nor U27682 (N_27682,N_27416,N_27412);
nand U27683 (N_27683,N_27406,N_27425);
xor U27684 (N_27684,N_27468,N_27513);
nor U27685 (N_27685,N_27590,N_27448);
and U27686 (N_27686,N_27581,N_27519);
or U27687 (N_27687,N_27490,N_27403);
and U27688 (N_27688,N_27564,N_27599);
or U27689 (N_27689,N_27594,N_27498);
and U27690 (N_27690,N_27593,N_27540);
and U27691 (N_27691,N_27408,N_27494);
xnor U27692 (N_27692,N_27500,N_27484);
and U27693 (N_27693,N_27586,N_27532);
nand U27694 (N_27694,N_27560,N_27487);
nor U27695 (N_27695,N_27485,N_27589);
xor U27696 (N_27696,N_27561,N_27413);
nor U27697 (N_27697,N_27461,N_27587);
and U27698 (N_27698,N_27554,N_27497);
xnor U27699 (N_27699,N_27548,N_27596);
xor U27700 (N_27700,N_27562,N_27415);
nor U27701 (N_27701,N_27438,N_27549);
nand U27702 (N_27702,N_27586,N_27496);
nand U27703 (N_27703,N_27478,N_27445);
xor U27704 (N_27704,N_27595,N_27452);
nor U27705 (N_27705,N_27469,N_27458);
nand U27706 (N_27706,N_27584,N_27589);
and U27707 (N_27707,N_27478,N_27589);
nand U27708 (N_27708,N_27548,N_27493);
nand U27709 (N_27709,N_27497,N_27527);
xor U27710 (N_27710,N_27488,N_27503);
or U27711 (N_27711,N_27471,N_27416);
nor U27712 (N_27712,N_27423,N_27463);
xor U27713 (N_27713,N_27536,N_27588);
nand U27714 (N_27714,N_27514,N_27429);
nand U27715 (N_27715,N_27501,N_27524);
and U27716 (N_27716,N_27459,N_27537);
and U27717 (N_27717,N_27505,N_27559);
or U27718 (N_27718,N_27463,N_27458);
nand U27719 (N_27719,N_27455,N_27529);
xor U27720 (N_27720,N_27434,N_27452);
nand U27721 (N_27721,N_27476,N_27545);
nor U27722 (N_27722,N_27407,N_27488);
nor U27723 (N_27723,N_27413,N_27518);
nand U27724 (N_27724,N_27460,N_27437);
xnor U27725 (N_27725,N_27432,N_27504);
nor U27726 (N_27726,N_27577,N_27459);
or U27727 (N_27727,N_27430,N_27477);
nor U27728 (N_27728,N_27565,N_27538);
xnor U27729 (N_27729,N_27463,N_27502);
and U27730 (N_27730,N_27402,N_27570);
xor U27731 (N_27731,N_27400,N_27542);
and U27732 (N_27732,N_27405,N_27547);
or U27733 (N_27733,N_27493,N_27507);
nand U27734 (N_27734,N_27516,N_27558);
nor U27735 (N_27735,N_27502,N_27417);
nand U27736 (N_27736,N_27402,N_27431);
xor U27737 (N_27737,N_27412,N_27560);
nor U27738 (N_27738,N_27580,N_27541);
nand U27739 (N_27739,N_27478,N_27578);
or U27740 (N_27740,N_27523,N_27518);
or U27741 (N_27741,N_27416,N_27581);
nor U27742 (N_27742,N_27536,N_27471);
and U27743 (N_27743,N_27540,N_27433);
nand U27744 (N_27744,N_27402,N_27429);
xor U27745 (N_27745,N_27524,N_27467);
nor U27746 (N_27746,N_27571,N_27529);
nor U27747 (N_27747,N_27582,N_27575);
and U27748 (N_27748,N_27495,N_27417);
or U27749 (N_27749,N_27508,N_27540);
xor U27750 (N_27750,N_27505,N_27419);
nor U27751 (N_27751,N_27520,N_27547);
and U27752 (N_27752,N_27545,N_27442);
and U27753 (N_27753,N_27407,N_27529);
nor U27754 (N_27754,N_27540,N_27405);
and U27755 (N_27755,N_27475,N_27503);
or U27756 (N_27756,N_27430,N_27584);
nor U27757 (N_27757,N_27447,N_27480);
nor U27758 (N_27758,N_27419,N_27489);
nand U27759 (N_27759,N_27447,N_27586);
nand U27760 (N_27760,N_27586,N_27564);
xnor U27761 (N_27761,N_27481,N_27561);
xor U27762 (N_27762,N_27526,N_27471);
or U27763 (N_27763,N_27578,N_27459);
nand U27764 (N_27764,N_27414,N_27492);
xor U27765 (N_27765,N_27553,N_27518);
nand U27766 (N_27766,N_27567,N_27581);
or U27767 (N_27767,N_27456,N_27448);
or U27768 (N_27768,N_27579,N_27498);
xnor U27769 (N_27769,N_27444,N_27455);
or U27770 (N_27770,N_27592,N_27490);
and U27771 (N_27771,N_27452,N_27542);
xnor U27772 (N_27772,N_27413,N_27431);
or U27773 (N_27773,N_27576,N_27535);
nor U27774 (N_27774,N_27449,N_27558);
nor U27775 (N_27775,N_27477,N_27577);
nor U27776 (N_27776,N_27407,N_27562);
nand U27777 (N_27777,N_27577,N_27420);
nand U27778 (N_27778,N_27480,N_27534);
or U27779 (N_27779,N_27504,N_27498);
nor U27780 (N_27780,N_27591,N_27482);
or U27781 (N_27781,N_27527,N_27523);
xor U27782 (N_27782,N_27462,N_27558);
nor U27783 (N_27783,N_27478,N_27598);
nand U27784 (N_27784,N_27482,N_27445);
xor U27785 (N_27785,N_27517,N_27425);
nand U27786 (N_27786,N_27511,N_27571);
or U27787 (N_27787,N_27520,N_27522);
xnor U27788 (N_27788,N_27593,N_27591);
nand U27789 (N_27789,N_27567,N_27570);
nand U27790 (N_27790,N_27423,N_27547);
nand U27791 (N_27791,N_27566,N_27489);
or U27792 (N_27792,N_27447,N_27544);
nor U27793 (N_27793,N_27546,N_27440);
or U27794 (N_27794,N_27481,N_27555);
and U27795 (N_27795,N_27585,N_27496);
and U27796 (N_27796,N_27408,N_27448);
nor U27797 (N_27797,N_27477,N_27479);
nor U27798 (N_27798,N_27473,N_27421);
or U27799 (N_27799,N_27555,N_27485);
nand U27800 (N_27800,N_27606,N_27705);
nand U27801 (N_27801,N_27666,N_27657);
nand U27802 (N_27802,N_27625,N_27683);
nor U27803 (N_27803,N_27677,N_27698);
xnor U27804 (N_27804,N_27739,N_27624);
nor U27805 (N_27805,N_27729,N_27785);
xnor U27806 (N_27806,N_27675,N_27740);
nand U27807 (N_27807,N_27619,N_27717);
nor U27808 (N_27808,N_27798,N_27608);
nor U27809 (N_27809,N_27688,N_27747);
xnor U27810 (N_27810,N_27644,N_27661);
or U27811 (N_27811,N_27707,N_27646);
xor U27812 (N_27812,N_27792,N_27744);
and U27813 (N_27813,N_27713,N_27794);
xor U27814 (N_27814,N_27746,N_27687);
nand U27815 (N_27815,N_27647,N_27730);
nand U27816 (N_27816,N_27708,N_27775);
xor U27817 (N_27817,N_27702,N_27658);
xor U27818 (N_27818,N_27632,N_27762);
xor U27819 (N_27819,N_27628,N_27635);
or U27820 (N_27820,N_27768,N_27736);
or U27821 (N_27821,N_27641,N_27604);
xnor U27822 (N_27822,N_27672,N_27694);
nor U27823 (N_27823,N_27753,N_27784);
nor U27824 (N_27824,N_27665,N_27638);
and U27825 (N_27825,N_27699,N_27640);
and U27826 (N_27826,N_27718,N_27710);
and U27827 (N_27827,N_27685,N_27626);
or U27828 (N_27828,N_27701,N_27787);
or U27829 (N_27829,N_27793,N_27652);
nand U27830 (N_27830,N_27720,N_27735);
nand U27831 (N_27831,N_27791,N_27680);
and U27832 (N_27832,N_27689,N_27603);
nor U27833 (N_27833,N_27732,N_27622);
nand U27834 (N_27834,N_27748,N_27754);
and U27835 (N_27835,N_27654,N_27734);
nand U27836 (N_27836,N_27769,N_27673);
nand U27837 (N_27837,N_27613,N_27648);
and U27838 (N_27838,N_27656,N_27786);
or U27839 (N_27839,N_27712,N_27767);
xnor U27840 (N_27840,N_27738,N_27618);
nor U27841 (N_27841,N_27684,N_27715);
nand U27842 (N_27842,N_27636,N_27779);
or U27843 (N_27843,N_27758,N_27686);
and U27844 (N_27844,N_27716,N_27772);
nand U27845 (N_27845,N_27771,N_27700);
and U27846 (N_27846,N_27601,N_27679);
or U27847 (N_27847,N_27759,N_27782);
or U27848 (N_27848,N_27722,N_27653);
nand U27849 (N_27849,N_27755,N_27721);
xnor U27850 (N_27850,N_27728,N_27778);
nand U27851 (N_27851,N_27690,N_27693);
and U27852 (N_27852,N_27612,N_27692);
xor U27853 (N_27853,N_27627,N_27639);
nand U27854 (N_27854,N_27725,N_27674);
and U27855 (N_27855,N_27695,N_27663);
or U27856 (N_27856,N_27760,N_27678);
and U27857 (N_27857,N_27602,N_27799);
or U27858 (N_27858,N_27671,N_27696);
or U27859 (N_27859,N_27670,N_27697);
and U27860 (N_27860,N_27764,N_27777);
nor U27861 (N_27861,N_27743,N_27714);
and U27862 (N_27862,N_27774,N_27751);
or U27863 (N_27863,N_27643,N_27709);
nand U27864 (N_27864,N_27669,N_27691);
nand U27865 (N_27865,N_27719,N_27745);
and U27866 (N_27866,N_27733,N_27763);
nand U27867 (N_27867,N_27617,N_27660);
and U27868 (N_27868,N_27650,N_27757);
nor U27869 (N_27869,N_27620,N_27655);
and U27870 (N_27870,N_27727,N_27780);
nand U27871 (N_27871,N_27607,N_27731);
xor U27872 (N_27872,N_27796,N_27776);
nor U27873 (N_27873,N_27797,N_27706);
xnor U27874 (N_27874,N_27667,N_27681);
or U27875 (N_27875,N_27614,N_27605);
nand U27876 (N_27876,N_27723,N_27742);
xor U27877 (N_27877,N_27789,N_27703);
or U27878 (N_27878,N_27621,N_27741);
nand U27879 (N_27879,N_27756,N_27682);
or U27880 (N_27880,N_27750,N_27600);
and U27881 (N_27881,N_27752,N_27761);
nor U27882 (N_27882,N_27737,N_27711);
and U27883 (N_27883,N_27795,N_27634);
xnor U27884 (N_27884,N_27664,N_27609);
or U27885 (N_27885,N_27724,N_27704);
or U27886 (N_27886,N_27637,N_27676);
and U27887 (N_27887,N_27629,N_27668);
or U27888 (N_27888,N_27659,N_27790);
nand U27889 (N_27889,N_27630,N_27766);
or U27890 (N_27890,N_27631,N_27749);
or U27891 (N_27891,N_27633,N_27783);
and U27892 (N_27892,N_27781,N_27645);
nor U27893 (N_27893,N_27773,N_27623);
or U27894 (N_27894,N_27662,N_27642);
nand U27895 (N_27895,N_27615,N_27770);
and U27896 (N_27896,N_27616,N_27788);
or U27897 (N_27897,N_27651,N_27726);
or U27898 (N_27898,N_27765,N_27610);
and U27899 (N_27899,N_27611,N_27649);
xnor U27900 (N_27900,N_27728,N_27769);
nor U27901 (N_27901,N_27690,N_27608);
or U27902 (N_27902,N_27607,N_27679);
nor U27903 (N_27903,N_27753,N_27781);
nand U27904 (N_27904,N_27759,N_27704);
and U27905 (N_27905,N_27735,N_27672);
or U27906 (N_27906,N_27627,N_27772);
and U27907 (N_27907,N_27773,N_27632);
or U27908 (N_27908,N_27628,N_27717);
and U27909 (N_27909,N_27602,N_27744);
xor U27910 (N_27910,N_27722,N_27773);
and U27911 (N_27911,N_27680,N_27679);
xnor U27912 (N_27912,N_27624,N_27727);
nand U27913 (N_27913,N_27765,N_27708);
xor U27914 (N_27914,N_27632,N_27684);
xor U27915 (N_27915,N_27659,N_27617);
xor U27916 (N_27916,N_27751,N_27740);
nand U27917 (N_27917,N_27651,N_27600);
nand U27918 (N_27918,N_27625,N_27719);
or U27919 (N_27919,N_27784,N_27700);
nand U27920 (N_27920,N_27799,N_27683);
and U27921 (N_27921,N_27742,N_27758);
nand U27922 (N_27922,N_27701,N_27628);
and U27923 (N_27923,N_27660,N_27635);
or U27924 (N_27924,N_27751,N_27667);
nand U27925 (N_27925,N_27792,N_27714);
nand U27926 (N_27926,N_27770,N_27656);
or U27927 (N_27927,N_27632,N_27627);
nand U27928 (N_27928,N_27674,N_27710);
nand U27929 (N_27929,N_27705,N_27728);
nand U27930 (N_27930,N_27727,N_27796);
xor U27931 (N_27931,N_27790,N_27665);
nand U27932 (N_27932,N_27772,N_27661);
nor U27933 (N_27933,N_27740,N_27716);
nor U27934 (N_27934,N_27730,N_27600);
xor U27935 (N_27935,N_27779,N_27604);
or U27936 (N_27936,N_27606,N_27624);
nand U27937 (N_27937,N_27786,N_27751);
nand U27938 (N_27938,N_27656,N_27732);
nor U27939 (N_27939,N_27683,N_27605);
nand U27940 (N_27940,N_27690,N_27767);
nand U27941 (N_27941,N_27675,N_27786);
and U27942 (N_27942,N_27740,N_27747);
or U27943 (N_27943,N_27656,N_27600);
and U27944 (N_27944,N_27763,N_27727);
nand U27945 (N_27945,N_27768,N_27737);
or U27946 (N_27946,N_27730,N_27637);
and U27947 (N_27947,N_27676,N_27770);
nor U27948 (N_27948,N_27612,N_27731);
and U27949 (N_27949,N_27773,N_27635);
nor U27950 (N_27950,N_27618,N_27737);
xnor U27951 (N_27951,N_27769,N_27626);
and U27952 (N_27952,N_27770,N_27661);
nand U27953 (N_27953,N_27758,N_27702);
and U27954 (N_27954,N_27748,N_27779);
nor U27955 (N_27955,N_27777,N_27720);
and U27956 (N_27956,N_27718,N_27627);
and U27957 (N_27957,N_27677,N_27611);
nor U27958 (N_27958,N_27731,N_27756);
or U27959 (N_27959,N_27758,N_27792);
nand U27960 (N_27960,N_27790,N_27620);
nor U27961 (N_27961,N_27658,N_27604);
nor U27962 (N_27962,N_27667,N_27743);
nand U27963 (N_27963,N_27719,N_27640);
nor U27964 (N_27964,N_27704,N_27647);
nand U27965 (N_27965,N_27725,N_27741);
and U27966 (N_27966,N_27698,N_27632);
and U27967 (N_27967,N_27660,N_27753);
nand U27968 (N_27968,N_27710,N_27626);
nor U27969 (N_27969,N_27656,N_27624);
and U27970 (N_27970,N_27713,N_27660);
nor U27971 (N_27971,N_27656,N_27617);
nand U27972 (N_27972,N_27767,N_27773);
xor U27973 (N_27973,N_27678,N_27699);
and U27974 (N_27974,N_27711,N_27729);
xor U27975 (N_27975,N_27673,N_27654);
or U27976 (N_27976,N_27754,N_27652);
or U27977 (N_27977,N_27742,N_27777);
xor U27978 (N_27978,N_27770,N_27634);
xor U27979 (N_27979,N_27795,N_27689);
xnor U27980 (N_27980,N_27765,N_27728);
and U27981 (N_27981,N_27780,N_27731);
xnor U27982 (N_27982,N_27636,N_27709);
or U27983 (N_27983,N_27653,N_27752);
or U27984 (N_27984,N_27710,N_27610);
xnor U27985 (N_27985,N_27702,N_27786);
nand U27986 (N_27986,N_27611,N_27748);
xnor U27987 (N_27987,N_27627,N_27762);
xor U27988 (N_27988,N_27651,N_27760);
nand U27989 (N_27989,N_27748,N_27733);
and U27990 (N_27990,N_27723,N_27632);
nor U27991 (N_27991,N_27630,N_27707);
nor U27992 (N_27992,N_27707,N_27681);
xor U27993 (N_27993,N_27792,N_27746);
and U27994 (N_27994,N_27648,N_27644);
xnor U27995 (N_27995,N_27705,N_27712);
xnor U27996 (N_27996,N_27784,N_27655);
nor U27997 (N_27997,N_27723,N_27662);
xor U27998 (N_27998,N_27717,N_27655);
xnor U27999 (N_27999,N_27601,N_27681);
xnor U28000 (N_28000,N_27990,N_27902);
xnor U28001 (N_28001,N_27802,N_27836);
xnor U28002 (N_28002,N_27983,N_27847);
nor U28003 (N_28003,N_27935,N_27813);
nand U28004 (N_28004,N_27807,N_27894);
xor U28005 (N_28005,N_27900,N_27861);
nand U28006 (N_28006,N_27995,N_27823);
or U28007 (N_28007,N_27930,N_27924);
nand U28008 (N_28008,N_27821,N_27824);
and U28009 (N_28009,N_27942,N_27875);
xnor U28010 (N_28010,N_27944,N_27825);
or U28011 (N_28011,N_27876,N_27830);
nand U28012 (N_28012,N_27801,N_27997);
nor U28013 (N_28013,N_27984,N_27870);
nand U28014 (N_28014,N_27957,N_27895);
and U28015 (N_28015,N_27916,N_27989);
xor U28016 (N_28016,N_27881,N_27993);
and U28017 (N_28017,N_27908,N_27933);
nor U28018 (N_28018,N_27804,N_27854);
xnor U28019 (N_28019,N_27873,N_27891);
or U28020 (N_28020,N_27858,N_27954);
nor U28021 (N_28021,N_27831,N_27976);
nand U28022 (N_28022,N_27960,N_27961);
and U28023 (N_28023,N_27835,N_27827);
nor U28024 (N_28024,N_27864,N_27969);
nand U28025 (N_28025,N_27965,N_27917);
xnor U28026 (N_28026,N_27975,N_27842);
nand U28027 (N_28027,N_27951,N_27867);
nor U28028 (N_28028,N_27885,N_27849);
nor U28029 (N_28029,N_27928,N_27991);
nand U28030 (N_28030,N_27994,N_27898);
or U28031 (N_28031,N_27906,N_27946);
nand U28032 (N_28032,N_27803,N_27953);
nor U28033 (N_28033,N_27886,N_27815);
xnor U28034 (N_28034,N_27818,N_27879);
or U28035 (N_28035,N_27940,N_27808);
xor U28036 (N_28036,N_27986,N_27926);
xor U28037 (N_28037,N_27959,N_27950);
xnor U28038 (N_28038,N_27880,N_27923);
or U28039 (N_28039,N_27812,N_27988);
xor U28040 (N_28040,N_27914,N_27982);
nand U28041 (N_28041,N_27996,N_27871);
xnor U28042 (N_28042,N_27862,N_27838);
and U28043 (N_28043,N_27806,N_27826);
and U28044 (N_28044,N_27841,N_27979);
nor U28045 (N_28045,N_27853,N_27850);
xor U28046 (N_28046,N_27839,N_27913);
and U28047 (N_28047,N_27922,N_27868);
xnor U28048 (N_28048,N_27855,N_27943);
and U28049 (N_28049,N_27848,N_27890);
and U28050 (N_28050,N_27910,N_27819);
nand U28051 (N_28051,N_27893,N_27929);
or U28052 (N_28052,N_27896,N_27927);
nand U28053 (N_28053,N_27810,N_27919);
nor U28054 (N_28054,N_27814,N_27901);
xnor U28055 (N_28055,N_27963,N_27816);
nand U28056 (N_28056,N_27846,N_27905);
xor U28057 (N_28057,N_27955,N_27973);
nand U28058 (N_28058,N_27949,N_27903);
or U28059 (N_28059,N_27947,N_27852);
or U28060 (N_28060,N_27833,N_27840);
nor U28061 (N_28061,N_27844,N_27811);
and U28062 (N_28062,N_27941,N_27921);
and U28063 (N_28063,N_27837,N_27859);
or U28064 (N_28064,N_27998,N_27809);
nor U28065 (N_28065,N_27909,N_27931);
xnor U28066 (N_28066,N_27860,N_27925);
nand U28067 (N_28067,N_27851,N_27987);
and U28068 (N_28068,N_27932,N_27966);
and U28069 (N_28069,N_27805,N_27834);
nand U28070 (N_28070,N_27968,N_27883);
and U28071 (N_28071,N_27897,N_27934);
nor U28072 (N_28072,N_27939,N_27937);
and U28073 (N_28073,N_27978,N_27962);
and U28074 (N_28074,N_27822,N_27820);
or U28075 (N_28075,N_27887,N_27918);
xor U28076 (N_28076,N_27872,N_27828);
xnor U28077 (N_28077,N_27977,N_27936);
and U28078 (N_28078,N_27938,N_27845);
and U28079 (N_28079,N_27843,N_27958);
xor U28080 (N_28080,N_27948,N_27964);
or U28081 (N_28081,N_27863,N_27865);
nor U28082 (N_28082,N_27911,N_27952);
nand U28083 (N_28083,N_27912,N_27920);
and U28084 (N_28084,N_27945,N_27889);
or U28085 (N_28085,N_27980,N_27832);
nand U28086 (N_28086,N_27800,N_27857);
xor U28087 (N_28087,N_27882,N_27869);
nor U28088 (N_28088,N_27899,N_27970);
nand U28089 (N_28089,N_27856,N_27884);
xnor U28090 (N_28090,N_27878,N_27866);
nor U28091 (N_28091,N_27907,N_27915);
or U28092 (N_28092,N_27992,N_27974);
and U28093 (N_28093,N_27985,N_27967);
and U28094 (N_28094,N_27817,N_27904);
and U28095 (N_28095,N_27972,N_27956);
xnor U28096 (N_28096,N_27971,N_27981);
nor U28097 (N_28097,N_27874,N_27877);
or U28098 (N_28098,N_27888,N_27999);
xnor U28099 (N_28099,N_27829,N_27892);
xor U28100 (N_28100,N_27879,N_27979);
and U28101 (N_28101,N_27871,N_27957);
or U28102 (N_28102,N_27961,N_27955);
xor U28103 (N_28103,N_27972,N_27872);
xor U28104 (N_28104,N_27848,N_27841);
nand U28105 (N_28105,N_27840,N_27938);
or U28106 (N_28106,N_27859,N_27953);
and U28107 (N_28107,N_27816,N_27945);
xnor U28108 (N_28108,N_27988,N_27823);
nand U28109 (N_28109,N_27849,N_27974);
and U28110 (N_28110,N_27829,N_27961);
or U28111 (N_28111,N_27813,N_27809);
nor U28112 (N_28112,N_27901,N_27884);
nor U28113 (N_28113,N_27913,N_27942);
and U28114 (N_28114,N_27958,N_27971);
nor U28115 (N_28115,N_27951,N_27846);
nor U28116 (N_28116,N_27901,N_27911);
nor U28117 (N_28117,N_27944,N_27869);
nand U28118 (N_28118,N_27962,N_27844);
and U28119 (N_28119,N_27884,N_27921);
nand U28120 (N_28120,N_27994,N_27830);
xnor U28121 (N_28121,N_27980,N_27921);
or U28122 (N_28122,N_27967,N_27876);
nor U28123 (N_28123,N_27921,N_27903);
and U28124 (N_28124,N_27948,N_27999);
or U28125 (N_28125,N_27997,N_27882);
xor U28126 (N_28126,N_27998,N_27829);
xnor U28127 (N_28127,N_27964,N_27892);
xor U28128 (N_28128,N_27993,N_27832);
and U28129 (N_28129,N_27889,N_27946);
or U28130 (N_28130,N_27836,N_27835);
nor U28131 (N_28131,N_27922,N_27812);
xnor U28132 (N_28132,N_27938,N_27854);
nand U28133 (N_28133,N_27950,N_27867);
nor U28134 (N_28134,N_27849,N_27846);
nand U28135 (N_28135,N_27846,N_27947);
or U28136 (N_28136,N_27814,N_27902);
or U28137 (N_28137,N_27997,N_27902);
nand U28138 (N_28138,N_27945,N_27941);
nor U28139 (N_28139,N_27809,N_27988);
or U28140 (N_28140,N_27830,N_27877);
nand U28141 (N_28141,N_27928,N_27911);
or U28142 (N_28142,N_27995,N_27845);
and U28143 (N_28143,N_27867,N_27998);
and U28144 (N_28144,N_27890,N_27819);
nor U28145 (N_28145,N_27820,N_27913);
nand U28146 (N_28146,N_27969,N_27894);
and U28147 (N_28147,N_27857,N_27836);
or U28148 (N_28148,N_27980,N_27920);
nor U28149 (N_28149,N_27915,N_27989);
or U28150 (N_28150,N_27823,N_27847);
and U28151 (N_28151,N_27962,N_27996);
xor U28152 (N_28152,N_27873,N_27859);
xor U28153 (N_28153,N_27899,N_27845);
or U28154 (N_28154,N_27933,N_27841);
and U28155 (N_28155,N_27856,N_27946);
nor U28156 (N_28156,N_27911,N_27881);
nor U28157 (N_28157,N_27968,N_27953);
and U28158 (N_28158,N_27878,N_27940);
or U28159 (N_28159,N_27977,N_27911);
or U28160 (N_28160,N_27892,N_27849);
nand U28161 (N_28161,N_27957,N_27969);
nand U28162 (N_28162,N_27855,N_27871);
xnor U28163 (N_28163,N_27934,N_27917);
nor U28164 (N_28164,N_27993,N_27807);
nand U28165 (N_28165,N_27937,N_27823);
or U28166 (N_28166,N_27897,N_27945);
xnor U28167 (N_28167,N_27956,N_27806);
nand U28168 (N_28168,N_27946,N_27959);
nand U28169 (N_28169,N_27897,N_27816);
or U28170 (N_28170,N_27940,N_27817);
or U28171 (N_28171,N_27820,N_27975);
nor U28172 (N_28172,N_27858,N_27966);
xnor U28173 (N_28173,N_27934,N_27960);
or U28174 (N_28174,N_27866,N_27927);
xor U28175 (N_28175,N_27899,N_27810);
nor U28176 (N_28176,N_27808,N_27990);
and U28177 (N_28177,N_27976,N_27824);
nand U28178 (N_28178,N_27892,N_27946);
and U28179 (N_28179,N_27876,N_27944);
xor U28180 (N_28180,N_27907,N_27844);
nor U28181 (N_28181,N_27960,N_27824);
and U28182 (N_28182,N_27921,N_27871);
and U28183 (N_28183,N_27932,N_27955);
nand U28184 (N_28184,N_27938,N_27841);
and U28185 (N_28185,N_27960,N_27914);
or U28186 (N_28186,N_27899,N_27922);
or U28187 (N_28187,N_27901,N_27968);
or U28188 (N_28188,N_27861,N_27936);
and U28189 (N_28189,N_27904,N_27873);
and U28190 (N_28190,N_27983,N_27897);
nor U28191 (N_28191,N_27933,N_27984);
nand U28192 (N_28192,N_27955,N_27927);
xnor U28193 (N_28193,N_27808,N_27836);
and U28194 (N_28194,N_27912,N_27900);
xor U28195 (N_28195,N_27916,N_27941);
or U28196 (N_28196,N_27950,N_27825);
or U28197 (N_28197,N_27867,N_27841);
nand U28198 (N_28198,N_27899,N_27997);
nor U28199 (N_28199,N_27905,N_27855);
nand U28200 (N_28200,N_28039,N_28126);
nor U28201 (N_28201,N_28100,N_28078);
nand U28202 (N_28202,N_28085,N_28043);
xor U28203 (N_28203,N_28006,N_28068);
and U28204 (N_28204,N_28000,N_28155);
nand U28205 (N_28205,N_28028,N_28011);
xnor U28206 (N_28206,N_28056,N_28088);
and U28207 (N_28207,N_28076,N_28116);
nand U28208 (N_28208,N_28159,N_28025);
and U28209 (N_28209,N_28045,N_28102);
nand U28210 (N_28210,N_28103,N_28147);
xnor U28211 (N_28211,N_28125,N_28049);
xnor U28212 (N_28212,N_28086,N_28097);
xnor U28213 (N_28213,N_28072,N_28142);
or U28214 (N_28214,N_28041,N_28164);
nand U28215 (N_28215,N_28062,N_28090);
nand U28216 (N_28216,N_28027,N_28128);
or U28217 (N_28217,N_28193,N_28141);
nor U28218 (N_28218,N_28196,N_28077);
and U28219 (N_28219,N_28019,N_28163);
or U28220 (N_28220,N_28152,N_28190);
nor U28221 (N_28221,N_28178,N_28013);
nor U28222 (N_28222,N_28122,N_28038);
xnor U28223 (N_28223,N_28124,N_28053);
or U28224 (N_28224,N_28160,N_28092);
xor U28225 (N_28225,N_28114,N_28172);
nor U28226 (N_28226,N_28071,N_28018);
and U28227 (N_28227,N_28179,N_28131);
xnor U28228 (N_28228,N_28058,N_28166);
and U28229 (N_28229,N_28067,N_28066);
nand U28230 (N_28230,N_28079,N_28009);
xor U28231 (N_28231,N_28199,N_28171);
xor U28232 (N_28232,N_28096,N_28177);
or U28233 (N_28233,N_28005,N_28063);
nor U28234 (N_28234,N_28134,N_28111);
nor U28235 (N_28235,N_28051,N_28149);
nand U28236 (N_28236,N_28161,N_28098);
or U28237 (N_28237,N_28115,N_28198);
nand U28238 (N_28238,N_28113,N_28118);
nor U28239 (N_28239,N_28082,N_28004);
and U28240 (N_28240,N_28055,N_28065);
nor U28241 (N_28241,N_28094,N_28099);
or U28242 (N_28242,N_28117,N_28061);
xnor U28243 (N_28243,N_28133,N_28074);
or U28244 (N_28244,N_28144,N_28042);
nand U28245 (N_28245,N_28120,N_28022);
nand U28246 (N_28246,N_28154,N_28129);
and U28247 (N_28247,N_28084,N_28162);
xnor U28248 (N_28248,N_28057,N_28060);
xnor U28249 (N_28249,N_28010,N_28180);
nand U28250 (N_28250,N_28073,N_28137);
xnor U28251 (N_28251,N_28015,N_28087);
and U28252 (N_28252,N_28101,N_28192);
xnor U28253 (N_28253,N_28020,N_28023);
nand U28254 (N_28254,N_28044,N_28031);
nand U28255 (N_28255,N_28003,N_28059);
xnor U28256 (N_28256,N_28104,N_28143);
nor U28257 (N_28257,N_28151,N_28140);
and U28258 (N_28258,N_28046,N_28127);
and U28259 (N_28259,N_28109,N_28107);
or U28260 (N_28260,N_28052,N_28170);
xor U28261 (N_28261,N_28167,N_28145);
and U28262 (N_28262,N_28093,N_28070);
xnor U28263 (N_28263,N_28110,N_28157);
xnor U28264 (N_28264,N_28139,N_28001);
nand U28265 (N_28265,N_28105,N_28150);
and U28266 (N_28266,N_28012,N_28138);
or U28267 (N_28267,N_28069,N_28081);
or U28268 (N_28268,N_28030,N_28156);
or U28269 (N_28269,N_28007,N_28123);
and U28270 (N_28270,N_28106,N_28002);
nor U28271 (N_28271,N_28064,N_28029);
or U28272 (N_28272,N_28026,N_28014);
nand U28273 (N_28273,N_28054,N_28047);
xor U28274 (N_28274,N_28095,N_28165);
and U28275 (N_28275,N_28189,N_28040);
and U28276 (N_28276,N_28173,N_28032);
xnor U28277 (N_28277,N_28181,N_28037);
or U28278 (N_28278,N_28036,N_28083);
or U28279 (N_28279,N_28175,N_28197);
xor U28280 (N_28280,N_28194,N_28187);
xnor U28281 (N_28281,N_28130,N_28158);
or U28282 (N_28282,N_28091,N_28136);
nand U28283 (N_28283,N_28182,N_28017);
or U28284 (N_28284,N_28168,N_28184);
nor U28285 (N_28285,N_28024,N_28121);
and U28286 (N_28286,N_28148,N_28112);
nand U28287 (N_28287,N_28119,N_28185);
or U28288 (N_28288,N_28186,N_28075);
or U28289 (N_28289,N_28169,N_28188);
nor U28290 (N_28290,N_28108,N_28195);
xor U28291 (N_28291,N_28191,N_28034);
nor U28292 (N_28292,N_28016,N_28050);
nor U28293 (N_28293,N_28135,N_28132);
and U28294 (N_28294,N_28080,N_28008);
xor U28295 (N_28295,N_28048,N_28174);
xnor U28296 (N_28296,N_28176,N_28021);
or U28297 (N_28297,N_28089,N_28035);
or U28298 (N_28298,N_28153,N_28183);
xor U28299 (N_28299,N_28146,N_28033);
nor U28300 (N_28300,N_28093,N_28109);
nand U28301 (N_28301,N_28121,N_28147);
and U28302 (N_28302,N_28181,N_28026);
nand U28303 (N_28303,N_28173,N_28013);
or U28304 (N_28304,N_28049,N_28022);
nand U28305 (N_28305,N_28196,N_28179);
nor U28306 (N_28306,N_28165,N_28030);
nand U28307 (N_28307,N_28035,N_28087);
nand U28308 (N_28308,N_28003,N_28180);
nand U28309 (N_28309,N_28052,N_28171);
nor U28310 (N_28310,N_28044,N_28098);
and U28311 (N_28311,N_28114,N_28092);
and U28312 (N_28312,N_28108,N_28199);
and U28313 (N_28313,N_28198,N_28125);
nand U28314 (N_28314,N_28081,N_28139);
nand U28315 (N_28315,N_28092,N_28139);
and U28316 (N_28316,N_28062,N_28098);
and U28317 (N_28317,N_28198,N_28122);
and U28318 (N_28318,N_28056,N_28010);
nand U28319 (N_28319,N_28145,N_28029);
and U28320 (N_28320,N_28182,N_28054);
nand U28321 (N_28321,N_28158,N_28015);
and U28322 (N_28322,N_28128,N_28087);
xor U28323 (N_28323,N_28081,N_28072);
and U28324 (N_28324,N_28099,N_28165);
nor U28325 (N_28325,N_28165,N_28004);
or U28326 (N_28326,N_28134,N_28193);
or U28327 (N_28327,N_28182,N_28105);
nor U28328 (N_28328,N_28163,N_28184);
nand U28329 (N_28329,N_28138,N_28104);
nor U28330 (N_28330,N_28144,N_28028);
and U28331 (N_28331,N_28181,N_28077);
nor U28332 (N_28332,N_28120,N_28159);
xor U28333 (N_28333,N_28130,N_28079);
and U28334 (N_28334,N_28198,N_28064);
xor U28335 (N_28335,N_28001,N_28044);
nand U28336 (N_28336,N_28020,N_28111);
or U28337 (N_28337,N_28008,N_28034);
xnor U28338 (N_28338,N_28089,N_28011);
and U28339 (N_28339,N_28173,N_28199);
and U28340 (N_28340,N_28039,N_28085);
or U28341 (N_28341,N_28147,N_28146);
or U28342 (N_28342,N_28185,N_28145);
nor U28343 (N_28343,N_28182,N_28131);
or U28344 (N_28344,N_28078,N_28013);
nand U28345 (N_28345,N_28142,N_28081);
xor U28346 (N_28346,N_28139,N_28184);
and U28347 (N_28347,N_28104,N_28177);
nand U28348 (N_28348,N_28143,N_28000);
xor U28349 (N_28349,N_28015,N_28164);
and U28350 (N_28350,N_28185,N_28148);
and U28351 (N_28351,N_28170,N_28097);
nor U28352 (N_28352,N_28171,N_28091);
or U28353 (N_28353,N_28184,N_28092);
nor U28354 (N_28354,N_28038,N_28089);
and U28355 (N_28355,N_28168,N_28124);
nand U28356 (N_28356,N_28014,N_28020);
nand U28357 (N_28357,N_28079,N_28135);
and U28358 (N_28358,N_28160,N_28086);
or U28359 (N_28359,N_28003,N_28131);
nand U28360 (N_28360,N_28066,N_28166);
nand U28361 (N_28361,N_28057,N_28095);
or U28362 (N_28362,N_28179,N_28103);
nand U28363 (N_28363,N_28024,N_28140);
nor U28364 (N_28364,N_28044,N_28005);
nand U28365 (N_28365,N_28099,N_28044);
nor U28366 (N_28366,N_28130,N_28173);
nand U28367 (N_28367,N_28145,N_28055);
xnor U28368 (N_28368,N_28035,N_28021);
nand U28369 (N_28369,N_28038,N_28136);
and U28370 (N_28370,N_28008,N_28049);
nand U28371 (N_28371,N_28129,N_28131);
nand U28372 (N_28372,N_28144,N_28153);
or U28373 (N_28373,N_28013,N_28184);
or U28374 (N_28374,N_28085,N_28075);
nand U28375 (N_28375,N_28172,N_28085);
and U28376 (N_28376,N_28073,N_28143);
and U28377 (N_28377,N_28010,N_28074);
or U28378 (N_28378,N_28059,N_28151);
or U28379 (N_28379,N_28045,N_28024);
and U28380 (N_28380,N_28084,N_28119);
or U28381 (N_28381,N_28135,N_28087);
xnor U28382 (N_28382,N_28071,N_28046);
nand U28383 (N_28383,N_28123,N_28001);
and U28384 (N_28384,N_28014,N_28168);
nor U28385 (N_28385,N_28152,N_28173);
xnor U28386 (N_28386,N_28155,N_28008);
nand U28387 (N_28387,N_28116,N_28068);
nor U28388 (N_28388,N_28119,N_28150);
xor U28389 (N_28389,N_28023,N_28086);
and U28390 (N_28390,N_28020,N_28120);
nand U28391 (N_28391,N_28171,N_28191);
nand U28392 (N_28392,N_28053,N_28035);
or U28393 (N_28393,N_28065,N_28109);
xor U28394 (N_28394,N_28082,N_28167);
nor U28395 (N_28395,N_28151,N_28097);
nor U28396 (N_28396,N_28190,N_28073);
and U28397 (N_28397,N_28022,N_28117);
xor U28398 (N_28398,N_28098,N_28085);
or U28399 (N_28399,N_28175,N_28154);
xnor U28400 (N_28400,N_28272,N_28278);
xor U28401 (N_28401,N_28369,N_28239);
xor U28402 (N_28402,N_28286,N_28379);
or U28403 (N_28403,N_28360,N_28389);
nand U28404 (N_28404,N_28245,N_28335);
nand U28405 (N_28405,N_28364,N_28208);
and U28406 (N_28406,N_28355,N_28248);
or U28407 (N_28407,N_28229,N_28366);
or U28408 (N_28408,N_28331,N_28304);
and U28409 (N_28409,N_28361,N_28319);
and U28410 (N_28410,N_28214,N_28223);
nor U28411 (N_28411,N_28289,N_28235);
xnor U28412 (N_28412,N_28377,N_28329);
xor U28413 (N_28413,N_28232,N_28336);
and U28414 (N_28414,N_28343,N_28399);
or U28415 (N_28415,N_28337,N_28397);
xnor U28416 (N_28416,N_28376,N_28370);
xor U28417 (N_28417,N_28259,N_28238);
and U28418 (N_28418,N_28398,N_28263);
nor U28419 (N_28419,N_28274,N_28270);
nor U28420 (N_28420,N_28385,N_28316);
or U28421 (N_28421,N_28254,N_28326);
and U28422 (N_28422,N_28260,N_28344);
and U28423 (N_28423,N_28320,N_28382);
nor U28424 (N_28424,N_28368,N_28293);
and U28425 (N_28425,N_28313,N_28381);
nor U28426 (N_28426,N_28384,N_28297);
or U28427 (N_28427,N_28202,N_28394);
nand U28428 (N_28428,N_28213,N_28252);
nor U28429 (N_28429,N_28255,N_28277);
nor U28430 (N_28430,N_28328,N_28350);
or U28431 (N_28431,N_28296,N_28221);
nor U28432 (N_28432,N_28318,N_28287);
nor U28433 (N_28433,N_28317,N_28386);
or U28434 (N_28434,N_28325,N_28338);
nor U28435 (N_28435,N_28341,N_28210);
nand U28436 (N_28436,N_28392,N_28268);
or U28437 (N_28437,N_28351,N_28378);
nor U28438 (N_28438,N_28256,N_28310);
and U28439 (N_28439,N_28375,N_28315);
or U28440 (N_28440,N_28393,N_28371);
and U28441 (N_28441,N_28215,N_28227);
or U28442 (N_28442,N_28226,N_28345);
nand U28443 (N_28443,N_28373,N_28200);
or U28444 (N_28444,N_28363,N_28233);
and U28445 (N_28445,N_28251,N_28246);
nand U28446 (N_28446,N_28295,N_28311);
xor U28447 (N_28447,N_28240,N_28241);
nor U28448 (N_28448,N_28307,N_28211);
and U28449 (N_28449,N_28222,N_28249);
nor U28450 (N_28450,N_28264,N_28282);
and U28451 (N_28451,N_28340,N_28281);
and U28452 (N_28452,N_28288,N_28275);
xor U28453 (N_28453,N_28216,N_28262);
and U28454 (N_28454,N_28280,N_28327);
and U28455 (N_28455,N_28243,N_28266);
nand U28456 (N_28456,N_28261,N_28242);
or U28457 (N_28457,N_28212,N_28285);
xor U28458 (N_28458,N_28205,N_28383);
xnor U28459 (N_28459,N_28395,N_28225);
and U28460 (N_28460,N_28312,N_28306);
nand U28461 (N_28461,N_28358,N_28390);
or U28462 (N_28462,N_28324,N_28333);
nand U28463 (N_28463,N_28298,N_28244);
nand U28464 (N_28464,N_28291,N_28339);
nand U28465 (N_28465,N_28203,N_28299);
nand U28466 (N_28466,N_28354,N_28365);
nand U28467 (N_28467,N_28357,N_28367);
xor U28468 (N_28468,N_28234,N_28359);
xor U28469 (N_28469,N_28250,N_28330);
nor U28470 (N_28470,N_28253,N_28353);
xor U28471 (N_28471,N_28257,N_28219);
or U28472 (N_28472,N_28224,N_28396);
nand U28473 (N_28473,N_28207,N_28391);
xor U28474 (N_28474,N_28332,N_28321);
xor U28475 (N_28475,N_28267,N_28269);
xnor U28476 (N_28476,N_28294,N_28362);
nor U28477 (N_28477,N_28220,N_28292);
xnor U28478 (N_28478,N_28273,N_28301);
and U28479 (N_28479,N_28303,N_28276);
or U28480 (N_28480,N_28305,N_28322);
nand U28481 (N_28481,N_28380,N_28209);
and U28482 (N_28482,N_28346,N_28247);
and U28483 (N_28483,N_28283,N_28204);
or U28484 (N_28484,N_28279,N_28342);
nand U28485 (N_28485,N_28265,N_28228);
and U28486 (N_28486,N_28206,N_28308);
nor U28487 (N_28487,N_28334,N_28372);
or U28488 (N_28488,N_28314,N_28352);
nor U28489 (N_28489,N_28218,N_28348);
nand U28490 (N_28490,N_28388,N_28300);
nand U28491 (N_28491,N_28356,N_28258);
xor U28492 (N_28492,N_28231,N_28323);
and U28493 (N_28493,N_28349,N_28290);
nand U28494 (N_28494,N_28347,N_28284);
nand U28495 (N_28495,N_28236,N_28271);
or U28496 (N_28496,N_28217,N_28309);
xnor U28497 (N_28497,N_28237,N_28387);
nor U28498 (N_28498,N_28374,N_28302);
or U28499 (N_28499,N_28230,N_28201);
nor U28500 (N_28500,N_28227,N_28359);
and U28501 (N_28501,N_28376,N_28241);
or U28502 (N_28502,N_28250,N_28396);
or U28503 (N_28503,N_28263,N_28350);
nand U28504 (N_28504,N_28360,N_28319);
nor U28505 (N_28505,N_28332,N_28254);
nand U28506 (N_28506,N_28206,N_28393);
nand U28507 (N_28507,N_28215,N_28303);
or U28508 (N_28508,N_28282,N_28288);
or U28509 (N_28509,N_28242,N_28294);
xor U28510 (N_28510,N_28307,N_28222);
and U28511 (N_28511,N_28329,N_28335);
and U28512 (N_28512,N_28252,N_28394);
or U28513 (N_28513,N_28238,N_28221);
or U28514 (N_28514,N_28379,N_28363);
nand U28515 (N_28515,N_28328,N_28292);
nor U28516 (N_28516,N_28383,N_28366);
and U28517 (N_28517,N_28218,N_28298);
nor U28518 (N_28518,N_28332,N_28339);
and U28519 (N_28519,N_28367,N_28244);
or U28520 (N_28520,N_28302,N_28288);
or U28521 (N_28521,N_28274,N_28279);
and U28522 (N_28522,N_28343,N_28333);
nor U28523 (N_28523,N_28393,N_28389);
nand U28524 (N_28524,N_28254,N_28379);
and U28525 (N_28525,N_28293,N_28321);
nor U28526 (N_28526,N_28274,N_28225);
xnor U28527 (N_28527,N_28317,N_28243);
xnor U28528 (N_28528,N_28393,N_28314);
and U28529 (N_28529,N_28233,N_28356);
and U28530 (N_28530,N_28372,N_28374);
nor U28531 (N_28531,N_28206,N_28262);
or U28532 (N_28532,N_28239,N_28203);
xor U28533 (N_28533,N_28231,N_28347);
and U28534 (N_28534,N_28317,N_28309);
nand U28535 (N_28535,N_28277,N_28373);
or U28536 (N_28536,N_28351,N_28278);
nor U28537 (N_28537,N_28353,N_28224);
nor U28538 (N_28538,N_28217,N_28322);
xnor U28539 (N_28539,N_28237,N_28232);
nor U28540 (N_28540,N_28230,N_28386);
nand U28541 (N_28541,N_28348,N_28335);
and U28542 (N_28542,N_28388,N_28284);
xnor U28543 (N_28543,N_28335,N_28320);
or U28544 (N_28544,N_28201,N_28232);
xor U28545 (N_28545,N_28216,N_28368);
nor U28546 (N_28546,N_28346,N_28291);
or U28547 (N_28547,N_28246,N_28370);
nor U28548 (N_28548,N_28245,N_28200);
nand U28549 (N_28549,N_28221,N_28209);
nor U28550 (N_28550,N_28347,N_28253);
or U28551 (N_28551,N_28307,N_28206);
nand U28552 (N_28552,N_28271,N_28388);
and U28553 (N_28553,N_28206,N_28382);
xor U28554 (N_28554,N_28244,N_28289);
or U28555 (N_28555,N_28289,N_28374);
nand U28556 (N_28556,N_28383,N_28364);
nor U28557 (N_28557,N_28369,N_28212);
or U28558 (N_28558,N_28398,N_28308);
or U28559 (N_28559,N_28388,N_28353);
xnor U28560 (N_28560,N_28284,N_28386);
nand U28561 (N_28561,N_28331,N_28282);
nand U28562 (N_28562,N_28240,N_28272);
xor U28563 (N_28563,N_28248,N_28374);
or U28564 (N_28564,N_28234,N_28279);
and U28565 (N_28565,N_28252,N_28301);
nand U28566 (N_28566,N_28261,N_28336);
xnor U28567 (N_28567,N_28386,N_28240);
and U28568 (N_28568,N_28297,N_28264);
xor U28569 (N_28569,N_28399,N_28331);
and U28570 (N_28570,N_28201,N_28221);
nor U28571 (N_28571,N_28278,N_28237);
xor U28572 (N_28572,N_28386,N_28343);
nor U28573 (N_28573,N_28325,N_28256);
nand U28574 (N_28574,N_28237,N_28368);
xnor U28575 (N_28575,N_28362,N_28296);
or U28576 (N_28576,N_28329,N_28281);
and U28577 (N_28577,N_28229,N_28224);
nand U28578 (N_28578,N_28283,N_28248);
nor U28579 (N_28579,N_28371,N_28211);
xor U28580 (N_28580,N_28334,N_28204);
xnor U28581 (N_28581,N_28286,N_28359);
or U28582 (N_28582,N_28282,N_28350);
nand U28583 (N_28583,N_28251,N_28314);
nand U28584 (N_28584,N_28324,N_28204);
nand U28585 (N_28585,N_28277,N_28355);
or U28586 (N_28586,N_28308,N_28399);
or U28587 (N_28587,N_28237,N_28357);
and U28588 (N_28588,N_28203,N_28356);
nor U28589 (N_28589,N_28261,N_28347);
or U28590 (N_28590,N_28375,N_28247);
and U28591 (N_28591,N_28363,N_28315);
nor U28592 (N_28592,N_28254,N_28391);
xor U28593 (N_28593,N_28248,N_28261);
nor U28594 (N_28594,N_28215,N_28264);
or U28595 (N_28595,N_28390,N_28391);
and U28596 (N_28596,N_28270,N_28297);
nand U28597 (N_28597,N_28305,N_28255);
xnor U28598 (N_28598,N_28361,N_28328);
or U28599 (N_28599,N_28298,N_28266);
nor U28600 (N_28600,N_28575,N_28441);
xor U28601 (N_28601,N_28409,N_28506);
or U28602 (N_28602,N_28527,N_28455);
nand U28603 (N_28603,N_28595,N_28522);
nand U28604 (N_28604,N_28531,N_28478);
nor U28605 (N_28605,N_28592,N_28507);
and U28606 (N_28606,N_28412,N_28508);
nor U28607 (N_28607,N_28538,N_28540);
and U28608 (N_28608,N_28563,N_28517);
or U28609 (N_28609,N_28535,N_28405);
nand U28610 (N_28610,N_28464,N_28461);
or U28611 (N_28611,N_28480,N_28417);
nand U28612 (N_28612,N_28568,N_28536);
nand U28613 (N_28613,N_28463,N_28411);
or U28614 (N_28614,N_28526,N_28550);
xor U28615 (N_28615,N_28452,N_28499);
and U28616 (N_28616,N_28477,N_28494);
or U28617 (N_28617,N_28487,N_28559);
xor U28618 (N_28618,N_28496,N_28509);
or U28619 (N_28619,N_28533,N_28403);
nand U28620 (N_28620,N_28485,N_28497);
nand U28621 (N_28621,N_28484,N_28593);
nor U28622 (N_28622,N_28591,N_28489);
nand U28623 (N_28623,N_28493,N_28436);
nand U28624 (N_28624,N_28547,N_28472);
xor U28625 (N_28625,N_28425,N_28513);
nor U28626 (N_28626,N_28459,N_28467);
nor U28627 (N_28627,N_28514,N_28569);
xor U28628 (N_28628,N_28416,N_28537);
or U28629 (N_28629,N_28521,N_28561);
nand U28630 (N_28630,N_28528,N_28439);
xnor U28631 (N_28631,N_28468,N_28515);
xnor U28632 (N_28632,N_28437,N_28519);
or U28633 (N_28633,N_28510,N_28566);
and U28634 (N_28634,N_28486,N_28544);
or U28635 (N_28635,N_28539,N_28431);
nand U28636 (N_28636,N_28542,N_28580);
or U28637 (N_28637,N_28476,N_28564);
and U28638 (N_28638,N_28562,N_28512);
nand U28639 (N_28639,N_28483,N_28599);
or U28640 (N_28640,N_28490,N_28549);
nor U28641 (N_28641,N_28546,N_28402);
nor U28642 (N_28642,N_28554,N_28498);
xnor U28643 (N_28643,N_28598,N_28415);
nor U28644 (N_28644,N_28462,N_28430);
xnor U28645 (N_28645,N_28551,N_28432);
xor U28646 (N_28646,N_28534,N_28543);
nand U28647 (N_28647,N_28434,N_28438);
xnor U28648 (N_28648,N_28421,N_28488);
or U28649 (N_28649,N_28502,N_28520);
nand U28650 (N_28650,N_28456,N_28453);
nand U28651 (N_28651,N_28524,N_28571);
nor U28652 (N_28652,N_28423,N_28572);
and U28653 (N_28653,N_28470,N_28586);
nand U28654 (N_28654,N_28530,N_28473);
nor U28655 (N_28655,N_28597,N_28541);
or U28656 (N_28656,N_28511,N_28451);
nand U28657 (N_28657,N_28408,N_28492);
and U28658 (N_28658,N_28573,N_28577);
or U28659 (N_28659,N_28504,N_28525);
xnor U28660 (N_28660,N_28454,N_28435);
nor U28661 (N_28661,N_28594,N_28406);
nor U28662 (N_28662,N_28448,N_28558);
nand U28663 (N_28663,N_28555,N_28529);
nor U28664 (N_28664,N_28419,N_28427);
and U28665 (N_28665,N_28589,N_28420);
nor U28666 (N_28666,N_28576,N_28505);
and U28667 (N_28667,N_28545,N_28449);
or U28668 (N_28668,N_28422,N_28458);
nor U28669 (N_28669,N_28578,N_28560);
nor U28670 (N_28670,N_28479,N_28447);
nand U28671 (N_28671,N_28410,N_28474);
nor U28672 (N_28672,N_28428,N_28401);
xnor U28673 (N_28673,N_28582,N_28475);
nor U28674 (N_28674,N_28481,N_28596);
xnor U28675 (N_28675,N_28482,N_28585);
nand U28676 (N_28676,N_28501,N_28418);
xor U28677 (N_28677,N_28556,N_28495);
and U28678 (N_28678,N_28553,N_28518);
xor U28679 (N_28679,N_28523,N_28446);
nor U28680 (N_28680,N_28457,N_28413);
and U28681 (N_28681,N_28579,N_28584);
nor U28682 (N_28682,N_28570,N_28450);
nand U28683 (N_28683,N_28583,N_28590);
and U28684 (N_28684,N_28407,N_28426);
and U28685 (N_28685,N_28444,N_28491);
or U28686 (N_28686,N_28429,N_28565);
xor U28687 (N_28687,N_28465,N_28574);
and U28688 (N_28688,N_28588,N_28442);
or U28689 (N_28689,N_28532,N_28433);
and U28690 (N_28690,N_28460,N_28552);
xor U28691 (N_28691,N_28503,N_28548);
xnor U28692 (N_28692,N_28445,N_28500);
xor U28693 (N_28693,N_28567,N_28404);
or U28694 (N_28694,N_28557,N_28414);
and U28695 (N_28695,N_28466,N_28424);
and U28696 (N_28696,N_28471,N_28400);
xnor U28697 (N_28697,N_28469,N_28581);
or U28698 (N_28698,N_28587,N_28516);
nand U28699 (N_28699,N_28443,N_28440);
xnor U28700 (N_28700,N_28583,N_28507);
and U28701 (N_28701,N_28506,N_28431);
and U28702 (N_28702,N_28482,N_28533);
or U28703 (N_28703,N_28409,N_28477);
nor U28704 (N_28704,N_28490,N_28534);
nor U28705 (N_28705,N_28577,N_28492);
xnor U28706 (N_28706,N_28565,N_28553);
xnor U28707 (N_28707,N_28520,N_28416);
nor U28708 (N_28708,N_28543,N_28538);
nand U28709 (N_28709,N_28569,N_28451);
or U28710 (N_28710,N_28455,N_28469);
or U28711 (N_28711,N_28436,N_28599);
xor U28712 (N_28712,N_28403,N_28422);
nor U28713 (N_28713,N_28501,N_28455);
xor U28714 (N_28714,N_28592,N_28437);
and U28715 (N_28715,N_28490,N_28464);
nand U28716 (N_28716,N_28543,N_28552);
or U28717 (N_28717,N_28562,N_28559);
and U28718 (N_28718,N_28466,N_28465);
nor U28719 (N_28719,N_28516,N_28442);
or U28720 (N_28720,N_28558,N_28556);
xnor U28721 (N_28721,N_28576,N_28411);
and U28722 (N_28722,N_28541,N_28503);
nand U28723 (N_28723,N_28487,N_28568);
or U28724 (N_28724,N_28561,N_28441);
xnor U28725 (N_28725,N_28477,N_28411);
nand U28726 (N_28726,N_28484,N_28514);
or U28727 (N_28727,N_28502,N_28499);
and U28728 (N_28728,N_28484,N_28430);
or U28729 (N_28729,N_28412,N_28500);
xor U28730 (N_28730,N_28580,N_28559);
and U28731 (N_28731,N_28429,N_28538);
nand U28732 (N_28732,N_28485,N_28548);
or U28733 (N_28733,N_28500,N_28571);
nor U28734 (N_28734,N_28462,N_28517);
and U28735 (N_28735,N_28463,N_28487);
and U28736 (N_28736,N_28405,N_28479);
xnor U28737 (N_28737,N_28497,N_28433);
xor U28738 (N_28738,N_28505,N_28550);
nor U28739 (N_28739,N_28494,N_28469);
xor U28740 (N_28740,N_28527,N_28529);
xor U28741 (N_28741,N_28578,N_28428);
nand U28742 (N_28742,N_28486,N_28431);
nor U28743 (N_28743,N_28493,N_28509);
or U28744 (N_28744,N_28546,N_28429);
nand U28745 (N_28745,N_28532,N_28557);
nand U28746 (N_28746,N_28566,N_28434);
xor U28747 (N_28747,N_28561,N_28477);
xor U28748 (N_28748,N_28531,N_28406);
or U28749 (N_28749,N_28483,N_28450);
or U28750 (N_28750,N_28583,N_28511);
nor U28751 (N_28751,N_28424,N_28480);
xor U28752 (N_28752,N_28530,N_28523);
nor U28753 (N_28753,N_28489,N_28461);
nor U28754 (N_28754,N_28437,N_28483);
nand U28755 (N_28755,N_28422,N_28594);
xor U28756 (N_28756,N_28401,N_28507);
or U28757 (N_28757,N_28452,N_28519);
or U28758 (N_28758,N_28598,N_28490);
nand U28759 (N_28759,N_28400,N_28512);
and U28760 (N_28760,N_28402,N_28589);
nor U28761 (N_28761,N_28469,N_28449);
or U28762 (N_28762,N_28512,N_28556);
nor U28763 (N_28763,N_28598,N_28431);
or U28764 (N_28764,N_28525,N_28559);
or U28765 (N_28765,N_28580,N_28419);
and U28766 (N_28766,N_28435,N_28443);
nand U28767 (N_28767,N_28498,N_28447);
and U28768 (N_28768,N_28420,N_28580);
nor U28769 (N_28769,N_28478,N_28484);
nor U28770 (N_28770,N_28579,N_28432);
or U28771 (N_28771,N_28572,N_28414);
nor U28772 (N_28772,N_28463,N_28529);
nand U28773 (N_28773,N_28445,N_28546);
nand U28774 (N_28774,N_28460,N_28458);
or U28775 (N_28775,N_28571,N_28441);
nor U28776 (N_28776,N_28515,N_28417);
nand U28777 (N_28777,N_28557,N_28415);
or U28778 (N_28778,N_28561,N_28440);
xor U28779 (N_28779,N_28508,N_28498);
nand U28780 (N_28780,N_28414,N_28549);
nand U28781 (N_28781,N_28428,N_28570);
xnor U28782 (N_28782,N_28476,N_28596);
nor U28783 (N_28783,N_28498,N_28558);
xor U28784 (N_28784,N_28438,N_28563);
or U28785 (N_28785,N_28502,N_28507);
and U28786 (N_28786,N_28559,N_28546);
xnor U28787 (N_28787,N_28547,N_28586);
or U28788 (N_28788,N_28558,N_28555);
and U28789 (N_28789,N_28403,N_28545);
and U28790 (N_28790,N_28458,N_28551);
xnor U28791 (N_28791,N_28467,N_28494);
nand U28792 (N_28792,N_28587,N_28418);
and U28793 (N_28793,N_28435,N_28429);
or U28794 (N_28794,N_28573,N_28451);
xor U28795 (N_28795,N_28474,N_28470);
nand U28796 (N_28796,N_28545,N_28440);
nand U28797 (N_28797,N_28572,N_28549);
or U28798 (N_28798,N_28524,N_28563);
nor U28799 (N_28799,N_28442,N_28522);
and U28800 (N_28800,N_28610,N_28630);
and U28801 (N_28801,N_28623,N_28782);
or U28802 (N_28802,N_28673,N_28735);
nor U28803 (N_28803,N_28702,N_28769);
nand U28804 (N_28804,N_28786,N_28747);
and U28805 (N_28805,N_28723,N_28622);
xor U28806 (N_28806,N_28665,N_28671);
nor U28807 (N_28807,N_28685,N_28729);
nand U28808 (N_28808,N_28749,N_28701);
or U28809 (N_28809,N_28770,N_28645);
xor U28810 (N_28810,N_28664,N_28619);
xnor U28811 (N_28811,N_28670,N_28601);
or U28812 (N_28812,N_28710,N_28632);
xor U28813 (N_28813,N_28794,N_28773);
xnor U28814 (N_28814,N_28621,N_28774);
xnor U28815 (N_28815,N_28733,N_28765);
and U28816 (N_28816,N_28618,N_28654);
nand U28817 (N_28817,N_28694,N_28681);
xor U28818 (N_28818,N_28688,N_28675);
nand U28819 (N_28819,N_28649,N_28740);
or U28820 (N_28820,N_28613,N_28745);
nor U28821 (N_28821,N_28792,N_28793);
nand U28822 (N_28822,N_28795,N_28689);
nor U28823 (N_28823,N_28785,N_28627);
xor U28824 (N_28824,N_28600,N_28668);
nor U28825 (N_28825,N_28693,N_28763);
nor U28826 (N_28826,N_28755,N_28642);
and U28827 (N_28827,N_28636,N_28663);
nand U28828 (N_28828,N_28635,N_28698);
and U28829 (N_28829,N_28738,N_28638);
and U28830 (N_28830,N_28692,N_28691);
xor U28831 (N_28831,N_28617,N_28787);
xnor U28832 (N_28832,N_28620,N_28760);
nand U28833 (N_28833,N_28797,N_28661);
or U28834 (N_28834,N_28752,N_28759);
and U28835 (N_28835,N_28736,N_28644);
or U28836 (N_28836,N_28737,N_28669);
nand U28837 (N_28837,N_28777,N_28624);
and U28838 (N_28838,N_28742,N_28750);
and U28839 (N_28839,N_28775,N_28614);
nand U28840 (N_28840,N_28626,N_28656);
nor U28841 (N_28841,N_28608,N_28612);
nand U28842 (N_28842,N_28732,N_28653);
nand U28843 (N_28843,N_28726,N_28660);
or U28844 (N_28844,N_28764,N_28696);
nand U28845 (N_28845,N_28659,N_28607);
xnor U28846 (N_28846,N_28799,N_28634);
nand U28847 (N_28847,N_28643,N_28754);
nand U28848 (N_28848,N_28672,N_28666);
or U28849 (N_28849,N_28639,N_28730);
nor U28850 (N_28850,N_28652,N_28717);
nand U28851 (N_28851,N_28628,N_28791);
and U28852 (N_28852,N_28758,N_28728);
or U28853 (N_28853,N_28798,N_28684);
nand U28854 (N_28854,N_28743,N_28768);
and U28855 (N_28855,N_28678,N_28767);
or U28856 (N_28856,N_28780,N_28748);
xnor U28857 (N_28857,N_28676,N_28746);
nor U28858 (N_28858,N_28625,N_28631);
xnor U28859 (N_28859,N_28706,N_28646);
xnor U28860 (N_28860,N_28603,N_28658);
or U28861 (N_28861,N_28602,N_28761);
nor U28862 (N_28862,N_28680,N_28705);
xnor U28863 (N_28863,N_28699,N_28637);
and U28864 (N_28864,N_28725,N_28762);
or U28865 (N_28865,N_28779,N_28715);
xor U28866 (N_28866,N_28790,N_28741);
and U28867 (N_28867,N_28709,N_28690);
and U28868 (N_28868,N_28667,N_28718);
nor U28869 (N_28869,N_28766,N_28674);
and U28870 (N_28870,N_28784,N_28713);
or U28871 (N_28871,N_28605,N_28616);
and U28872 (N_28872,N_28778,N_28606);
and U28873 (N_28873,N_28716,N_28739);
xnor U28874 (N_28874,N_28640,N_28783);
and U28875 (N_28875,N_28744,N_28756);
and U28876 (N_28876,N_28700,N_28662);
nand U28877 (N_28877,N_28714,N_28703);
and U28878 (N_28878,N_28731,N_28751);
nand U28879 (N_28879,N_28734,N_28776);
nor U28880 (N_28880,N_28651,N_28772);
and U28881 (N_28881,N_28720,N_28704);
and U28882 (N_28882,N_28712,N_28722);
nor U28883 (N_28883,N_28641,N_28707);
nand U28884 (N_28884,N_28629,N_28708);
xor U28885 (N_28885,N_28604,N_28695);
nand U28886 (N_28886,N_28615,N_28655);
xor U28887 (N_28887,N_28683,N_28788);
xor U28888 (N_28888,N_28724,N_28648);
nand U28889 (N_28889,N_28796,N_28611);
nand U28890 (N_28890,N_28727,N_28757);
or U28891 (N_28891,N_28633,N_28771);
nand U28892 (N_28892,N_28682,N_28686);
nand U28893 (N_28893,N_28697,N_28789);
or U28894 (N_28894,N_28650,N_28679);
or U28895 (N_28895,N_28677,N_28657);
nand U28896 (N_28896,N_28753,N_28711);
nor U28897 (N_28897,N_28687,N_28609);
or U28898 (N_28898,N_28781,N_28719);
and U28899 (N_28899,N_28721,N_28647);
or U28900 (N_28900,N_28770,N_28745);
or U28901 (N_28901,N_28764,N_28617);
and U28902 (N_28902,N_28753,N_28736);
nor U28903 (N_28903,N_28774,N_28604);
or U28904 (N_28904,N_28724,N_28677);
nor U28905 (N_28905,N_28776,N_28689);
and U28906 (N_28906,N_28696,N_28734);
or U28907 (N_28907,N_28742,N_28684);
xor U28908 (N_28908,N_28754,N_28697);
nand U28909 (N_28909,N_28675,N_28702);
xnor U28910 (N_28910,N_28664,N_28610);
nor U28911 (N_28911,N_28618,N_28686);
and U28912 (N_28912,N_28733,N_28685);
nor U28913 (N_28913,N_28753,N_28793);
or U28914 (N_28914,N_28627,N_28770);
nand U28915 (N_28915,N_28608,N_28675);
or U28916 (N_28916,N_28622,N_28741);
xor U28917 (N_28917,N_28609,N_28741);
and U28918 (N_28918,N_28786,N_28717);
nor U28919 (N_28919,N_28631,N_28600);
nand U28920 (N_28920,N_28658,N_28790);
and U28921 (N_28921,N_28787,N_28614);
or U28922 (N_28922,N_28647,N_28638);
xnor U28923 (N_28923,N_28797,N_28722);
nor U28924 (N_28924,N_28631,N_28784);
nand U28925 (N_28925,N_28688,N_28737);
or U28926 (N_28926,N_28688,N_28625);
and U28927 (N_28927,N_28739,N_28681);
and U28928 (N_28928,N_28773,N_28692);
nor U28929 (N_28929,N_28769,N_28766);
nor U28930 (N_28930,N_28665,N_28674);
or U28931 (N_28931,N_28733,N_28663);
nand U28932 (N_28932,N_28762,N_28729);
nand U28933 (N_28933,N_28792,N_28605);
and U28934 (N_28934,N_28722,N_28720);
and U28935 (N_28935,N_28655,N_28660);
or U28936 (N_28936,N_28607,N_28634);
or U28937 (N_28937,N_28783,N_28760);
or U28938 (N_28938,N_28787,N_28733);
or U28939 (N_28939,N_28791,N_28775);
or U28940 (N_28940,N_28668,N_28770);
xnor U28941 (N_28941,N_28689,N_28697);
nor U28942 (N_28942,N_28612,N_28700);
nor U28943 (N_28943,N_28753,N_28737);
or U28944 (N_28944,N_28695,N_28660);
or U28945 (N_28945,N_28619,N_28655);
nor U28946 (N_28946,N_28782,N_28626);
xor U28947 (N_28947,N_28735,N_28728);
and U28948 (N_28948,N_28696,N_28677);
nor U28949 (N_28949,N_28778,N_28726);
and U28950 (N_28950,N_28609,N_28709);
nor U28951 (N_28951,N_28650,N_28794);
or U28952 (N_28952,N_28678,N_28700);
and U28953 (N_28953,N_28715,N_28645);
xor U28954 (N_28954,N_28730,N_28753);
nand U28955 (N_28955,N_28601,N_28645);
nor U28956 (N_28956,N_28614,N_28729);
xor U28957 (N_28957,N_28600,N_28782);
and U28958 (N_28958,N_28661,N_28779);
or U28959 (N_28959,N_28736,N_28646);
nor U28960 (N_28960,N_28740,N_28614);
nand U28961 (N_28961,N_28601,N_28755);
or U28962 (N_28962,N_28603,N_28782);
and U28963 (N_28963,N_28715,N_28778);
nor U28964 (N_28964,N_28713,N_28624);
and U28965 (N_28965,N_28662,N_28726);
or U28966 (N_28966,N_28789,N_28756);
nand U28967 (N_28967,N_28753,N_28624);
and U28968 (N_28968,N_28753,N_28689);
xor U28969 (N_28969,N_28670,N_28799);
and U28970 (N_28970,N_28787,N_28773);
xnor U28971 (N_28971,N_28703,N_28757);
xnor U28972 (N_28972,N_28746,N_28703);
and U28973 (N_28973,N_28765,N_28698);
nor U28974 (N_28974,N_28780,N_28724);
or U28975 (N_28975,N_28665,N_28703);
nand U28976 (N_28976,N_28624,N_28718);
or U28977 (N_28977,N_28636,N_28696);
nand U28978 (N_28978,N_28793,N_28705);
xor U28979 (N_28979,N_28786,N_28691);
and U28980 (N_28980,N_28644,N_28673);
or U28981 (N_28981,N_28607,N_28621);
and U28982 (N_28982,N_28716,N_28675);
or U28983 (N_28983,N_28743,N_28651);
xnor U28984 (N_28984,N_28672,N_28620);
nor U28985 (N_28985,N_28724,N_28628);
nor U28986 (N_28986,N_28752,N_28601);
or U28987 (N_28987,N_28739,N_28637);
nand U28988 (N_28988,N_28707,N_28788);
and U28989 (N_28989,N_28754,N_28765);
nor U28990 (N_28990,N_28650,N_28701);
nor U28991 (N_28991,N_28705,N_28792);
or U28992 (N_28992,N_28798,N_28766);
nor U28993 (N_28993,N_28674,N_28692);
nand U28994 (N_28994,N_28766,N_28729);
and U28995 (N_28995,N_28682,N_28740);
or U28996 (N_28996,N_28743,N_28631);
nand U28997 (N_28997,N_28674,N_28757);
nand U28998 (N_28998,N_28641,N_28741);
or U28999 (N_28999,N_28768,N_28780);
xnor U29000 (N_29000,N_28818,N_28857);
or U29001 (N_29001,N_28983,N_28896);
nor U29002 (N_29002,N_28942,N_28986);
or U29003 (N_29003,N_28807,N_28899);
or U29004 (N_29004,N_28909,N_28877);
or U29005 (N_29005,N_28805,N_28953);
xor U29006 (N_29006,N_28940,N_28936);
nand U29007 (N_29007,N_28801,N_28961);
and U29008 (N_29008,N_28887,N_28907);
or U29009 (N_29009,N_28965,N_28883);
or U29010 (N_29010,N_28931,N_28834);
and U29011 (N_29011,N_28910,N_28826);
xor U29012 (N_29012,N_28958,N_28941);
or U29013 (N_29013,N_28841,N_28959);
xnor U29014 (N_29014,N_28812,N_28995);
or U29015 (N_29015,N_28911,N_28985);
and U29016 (N_29016,N_28922,N_28919);
nor U29017 (N_29017,N_28978,N_28992);
and U29018 (N_29018,N_28854,N_28855);
and U29019 (N_29019,N_28902,N_28938);
xnor U29020 (N_29020,N_28871,N_28939);
nor U29021 (N_29021,N_28847,N_28886);
xor U29022 (N_29022,N_28976,N_28969);
nand U29023 (N_29023,N_28957,N_28858);
nand U29024 (N_29024,N_28815,N_28878);
and U29025 (N_29025,N_28913,N_28945);
nand U29026 (N_29026,N_28845,N_28989);
and U29027 (N_29027,N_28993,N_28814);
nor U29028 (N_29028,N_28954,N_28817);
xor U29029 (N_29029,N_28905,N_28808);
nand U29030 (N_29030,N_28920,N_28926);
xnor U29031 (N_29031,N_28864,N_28991);
and U29032 (N_29032,N_28984,N_28839);
or U29033 (N_29033,N_28891,N_28937);
nor U29034 (N_29034,N_28876,N_28832);
or U29035 (N_29035,N_28830,N_28868);
xor U29036 (N_29036,N_28990,N_28974);
nor U29037 (N_29037,N_28835,N_28924);
or U29038 (N_29038,N_28856,N_28944);
or U29039 (N_29039,N_28947,N_28897);
nand U29040 (N_29040,N_28943,N_28867);
or U29041 (N_29041,N_28934,N_28904);
nand U29042 (N_29042,N_28803,N_28853);
xnor U29043 (N_29043,N_28888,N_28823);
nor U29044 (N_29044,N_28873,N_28975);
or U29045 (N_29045,N_28800,N_28999);
nor U29046 (N_29046,N_28962,N_28972);
and U29047 (N_29047,N_28849,N_28948);
xor U29048 (N_29048,N_28949,N_28960);
and U29049 (N_29049,N_28932,N_28863);
nor U29050 (N_29050,N_28874,N_28982);
or U29051 (N_29051,N_28851,N_28901);
nor U29052 (N_29052,N_28816,N_28895);
nand U29053 (N_29053,N_28956,N_28935);
nor U29054 (N_29054,N_28870,N_28912);
nor U29055 (N_29055,N_28997,N_28894);
nand U29056 (N_29056,N_28981,N_28987);
nor U29057 (N_29057,N_28881,N_28806);
nand U29058 (N_29058,N_28963,N_28890);
and U29059 (N_29059,N_28859,N_28929);
or U29060 (N_29060,N_28980,N_28852);
xnor U29061 (N_29061,N_28875,N_28880);
or U29062 (N_29062,N_28996,N_28914);
nand U29063 (N_29063,N_28906,N_28872);
nand U29064 (N_29064,N_28885,N_28862);
xnor U29065 (N_29065,N_28952,N_28955);
nor U29066 (N_29066,N_28824,N_28933);
and U29067 (N_29067,N_28903,N_28898);
nor U29068 (N_29068,N_28916,N_28820);
nor U29069 (N_29069,N_28810,N_28811);
or U29070 (N_29070,N_28804,N_28950);
xnor U29071 (N_29071,N_28893,N_28973);
and U29072 (N_29072,N_28840,N_28848);
xnor U29073 (N_29073,N_28838,N_28918);
or U29074 (N_29074,N_28844,N_28998);
nand U29075 (N_29075,N_28821,N_28843);
nand U29076 (N_29076,N_28846,N_28928);
xor U29077 (N_29077,N_28979,N_28977);
nand U29078 (N_29078,N_28842,N_28825);
nor U29079 (N_29079,N_28946,N_28860);
or U29080 (N_29080,N_28861,N_28831);
nand U29081 (N_29081,N_28813,N_28966);
and U29082 (N_29082,N_28869,N_28829);
or U29083 (N_29083,N_28951,N_28967);
or U29084 (N_29084,N_28964,N_28994);
nand U29085 (N_29085,N_28915,N_28802);
xnor U29086 (N_29086,N_28819,N_28970);
nand U29087 (N_29087,N_28971,N_28827);
xnor U29088 (N_29088,N_28968,N_28865);
and U29089 (N_29089,N_28822,N_28917);
xor U29090 (N_29090,N_28927,N_28879);
or U29091 (N_29091,N_28900,N_28836);
and U29092 (N_29092,N_28837,N_28930);
nor U29093 (N_29093,N_28882,N_28828);
or U29094 (N_29094,N_28889,N_28892);
or U29095 (N_29095,N_28850,N_28809);
or U29096 (N_29096,N_28925,N_28988);
or U29097 (N_29097,N_28866,N_28908);
or U29098 (N_29098,N_28921,N_28884);
nand U29099 (N_29099,N_28833,N_28923);
nand U29100 (N_29100,N_28817,N_28868);
and U29101 (N_29101,N_28886,N_28987);
xor U29102 (N_29102,N_28950,N_28843);
or U29103 (N_29103,N_28870,N_28985);
nor U29104 (N_29104,N_28993,N_28855);
nor U29105 (N_29105,N_28908,N_28811);
or U29106 (N_29106,N_28812,N_28985);
and U29107 (N_29107,N_28926,N_28806);
and U29108 (N_29108,N_28869,N_28966);
and U29109 (N_29109,N_28971,N_28805);
nand U29110 (N_29110,N_28993,N_28813);
nand U29111 (N_29111,N_28936,N_28911);
and U29112 (N_29112,N_28861,N_28854);
xnor U29113 (N_29113,N_28872,N_28817);
or U29114 (N_29114,N_28824,N_28862);
nand U29115 (N_29115,N_28809,N_28912);
nand U29116 (N_29116,N_28849,N_28825);
nand U29117 (N_29117,N_28974,N_28873);
nand U29118 (N_29118,N_28880,N_28950);
xnor U29119 (N_29119,N_28883,N_28957);
xnor U29120 (N_29120,N_28876,N_28885);
nand U29121 (N_29121,N_28912,N_28994);
and U29122 (N_29122,N_28887,N_28805);
xnor U29123 (N_29123,N_28846,N_28961);
and U29124 (N_29124,N_28907,N_28919);
nor U29125 (N_29125,N_28822,N_28932);
or U29126 (N_29126,N_28873,N_28803);
or U29127 (N_29127,N_28844,N_28944);
xnor U29128 (N_29128,N_28873,N_28813);
nor U29129 (N_29129,N_28983,N_28866);
nand U29130 (N_29130,N_28831,N_28990);
or U29131 (N_29131,N_28999,N_28962);
nor U29132 (N_29132,N_28912,N_28814);
and U29133 (N_29133,N_28898,N_28951);
nand U29134 (N_29134,N_28897,N_28993);
nor U29135 (N_29135,N_28909,N_28853);
xor U29136 (N_29136,N_28955,N_28899);
nor U29137 (N_29137,N_28881,N_28925);
or U29138 (N_29138,N_28985,N_28950);
or U29139 (N_29139,N_28852,N_28848);
or U29140 (N_29140,N_28856,N_28937);
or U29141 (N_29141,N_28871,N_28949);
xnor U29142 (N_29142,N_28862,N_28900);
and U29143 (N_29143,N_28944,N_28910);
nand U29144 (N_29144,N_28894,N_28803);
nand U29145 (N_29145,N_28897,N_28976);
xor U29146 (N_29146,N_28815,N_28969);
and U29147 (N_29147,N_28824,N_28931);
nor U29148 (N_29148,N_28858,N_28806);
nand U29149 (N_29149,N_28900,N_28944);
nand U29150 (N_29150,N_28991,N_28911);
xnor U29151 (N_29151,N_28932,N_28979);
nand U29152 (N_29152,N_28957,N_28891);
nor U29153 (N_29153,N_28802,N_28898);
xnor U29154 (N_29154,N_28808,N_28950);
and U29155 (N_29155,N_28808,N_28813);
xnor U29156 (N_29156,N_28948,N_28899);
nor U29157 (N_29157,N_28811,N_28844);
nand U29158 (N_29158,N_28981,N_28808);
nand U29159 (N_29159,N_28852,N_28926);
or U29160 (N_29160,N_28929,N_28842);
xnor U29161 (N_29161,N_28858,N_28872);
or U29162 (N_29162,N_28983,N_28827);
nand U29163 (N_29163,N_28996,N_28990);
nand U29164 (N_29164,N_28981,N_28982);
xor U29165 (N_29165,N_28902,N_28819);
xor U29166 (N_29166,N_28942,N_28889);
nand U29167 (N_29167,N_28811,N_28854);
nand U29168 (N_29168,N_28871,N_28815);
or U29169 (N_29169,N_28803,N_28948);
nand U29170 (N_29170,N_28980,N_28900);
nand U29171 (N_29171,N_28960,N_28822);
or U29172 (N_29172,N_28873,N_28889);
and U29173 (N_29173,N_28888,N_28851);
or U29174 (N_29174,N_28999,N_28895);
nand U29175 (N_29175,N_28850,N_28910);
and U29176 (N_29176,N_28955,N_28821);
or U29177 (N_29177,N_28953,N_28974);
and U29178 (N_29178,N_28994,N_28990);
nand U29179 (N_29179,N_28902,N_28975);
nand U29180 (N_29180,N_28918,N_28870);
xor U29181 (N_29181,N_28922,N_28856);
or U29182 (N_29182,N_28890,N_28960);
nor U29183 (N_29183,N_28958,N_28806);
nand U29184 (N_29184,N_28950,N_28915);
and U29185 (N_29185,N_28986,N_28902);
and U29186 (N_29186,N_28819,N_28822);
nand U29187 (N_29187,N_28804,N_28946);
or U29188 (N_29188,N_28892,N_28921);
or U29189 (N_29189,N_28816,N_28818);
and U29190 (N_29190,N_28806,N_28874);
xor U29191 (N_29191,N_28946,N_28887);
nor U29192 (N_29192,N_28812,N_28948);
xor U29193 (N_29193,N_28832,N_28922);
xnor U29194 (N_29194,N_28986,N_28867);
nand U29195 (N_29195,N_28869,N_28981);
nand U29196 (N_29196,N_28847,N_28819);
nand U29197 (N_29197,N_28813,N_28835);
or U29198 (N_29198,N_28906,N_28958);
or U29199 (N_29199,N_28981,N_28888);
or U29200 (N_29200,N_29073,N_29050);
and U29201 (N_29201,N_29088,N_29119);
xor U29202 (N_29202,N_29036,N_29165);
or U29203 (N_29203,N_29125,N_29030);
nand U29204 (N_29204,N_29103,N_29011);
nor U29205 (N_29205,N_29173,N_29010);
nor U29206 (N_29206,N_29100,N_29107);
nand U29207 (N_29207,N_29059,N_29002);
nor U29208 (N_29208,N_29185,N_29066);
nor U29209 (N_29209,N_29101,N_29195);
and U29210 (N_29210,N_29074,N_29120);
and U29211 (N_29211,N_29003,N_29131);
and U29212 (N_29212,N_29175,N_29182);
xnor U29213 (N_29213,N_29089,N_29017);
nor U29214 (N_29214,N_29190,N_29106);
xnor U29215 (N_29215,N_29147,N_29031);
xnor U29216 (N_29216,N_29150,N_29012);
nor U29217 (N_29217,N_29133,N_29080);
xor U29218 (N_29218,N_29186,N_29157);
nand U29219 (N_29219,N_29057,N_29128);
nor U29220 (N_29220,N_29027,N_29086);
nand U29221 (N_29221,N_29054,N_29159);
or U29222 (N_29222,N_29124,N_29007);
nor U29223 (N_29223,N_29081,N_29016);
or U29224 (N_29224,N_29166,N_29009);
or U29225 (N_29225,N_29055,N_29155);
nor U29226 (N_29226,N_29047,N_29114);
nand U29227 (N_29227,N_29065,N_29113);
and U29228 (N_29228,N_29192,N_29033);
nor U29229 (N_29229,N_29077,N_29079);
nor U29230 (N_29230,N_29104,N_29044);
nor U29231 (N_29231,N_29025,N_29177);
xnor U29232 (N_29232,N_29041,N_29092);
or U29233 (N_29233,N_29162,N_29142);
nand U29234 (N_29234,N_29085,N_29035);
or U29235 (N_29235,N_29004,N_29102);
nor U29236 (N_29236,N_29134,N_29170);
nand U29237 (N_29237,N_29115,N_29069);
and U29238 (N_29238,N_29038,N_29161);
nor U29239 (N_29239,N_29014,N_29176);
and U29240 (N_29240,N_29046,N_29148);
or U29241 (N_29241,N_29156,N_29168);
nand U29242 (N_29242,N_29169,N_29179);
xor U29243 (N_29243,N_29060,N_29058);
xnor U29244 (N_29244,N_29049,N_29024);
nor U29245 (N_29245,N_29068,N_29196);
and U29246 (N_29246,N_29109,N_29015);
and U29247 (N_29247,N_29139,N_29132);
xnor U29248 (N_29248,N_29043,N_29140);
nor U29249 (N_29249,N_29199,N_29037);
nor U29250 (N_29250,N_29181,N_29076);
nand U29251 (N_29251,N_29137,N_29141);
nor U29252 (N_29252,N_29153,N_29056);
nand U29253 (N_29253,N_29075,N_29136);
and U29254 (N_29254,N_29138,N_29091);
nand U29255 (N_29255,N_29112,N_29197);
or U29256 (N_29256,N_29116,N_29152);
and U29257 (N_29257,N_29122,N_29174);
nand U29258 (N_29258,N_29172,N_29040);
and U29259 (N_29259,N_29063,N_29082);
and U29260 (N_29260,N_29039,N_29129);
nor U29261 (N_29261,N_29094,N_29064);
or U29262 (N_29262,N_29078,N_29093);
or U29263 (N_29263,N_29117,N_29163);
xor U29264 (N_29264,N_29105,N_29097);
xnor U29265 (N_29265,N_29029,N_29019);
xnor U29266 (N_29266,N_29171,N_29053);
or U29267 (N_29267,N_29087,N_29111);
or U29268 (N_29268,N_29130,N_29028);
and U29269 (N_29269,N_29167,N_29121);
or U29270 (N_29270,N_29052,N_29000);
nand U29271 (N_29271,N_29084,N_29126);
or U29272 (N_29272,N_29178,N_29083);
nor U29273 (N_29273,N_29021,N_29098);
nor U29274 (N_29274,N_29020,N_29135);
nand U29275 (N_29275,N_29072,N_29071);
nand U29276 (N_29276,N_29051,N_29045);
nand U29277 (N_29277,N_29149,N_29183);
xnor U29278 (N_29278,N_29006,N_29160);
xor U29279 (N_29279,N_29187,N_29118);
or U29280 (N_29280,N_29188,N_29090);
nor U29281 (N_29281,N_29032,N_29062);
and U29282 (N_29282,N_29198,N_29018);
and U29283 (N_29283,N_29026,N_29145);
nor U29284 (N_29284,N_29189,N_29061);
xor U29285 (N_29285,N_29193,N_29013);
or U29286 (N_29286,N_29008,N_29127);
nand U29287 (N_29287,N_29095,N_29096);
xnor U29288 (N_29288,N_29180,N_29110);
xor U29289 (N_29289,N_29022,N_29146);
nand U29290 (N_29290,N_29070,N_29184);
nand U29291 (N_29291,N_29143,N_29023);
nor U29292 (N_29292,N_29108,N_29144);
nor U29293 (N_29293,N_29005,N_29164);
or U29294 (N_29294,N_29048,N_29191);
or U29295 (N_29295,N_29123,N_29158);
or U29296 (N_29296,N_29099,N_29034);
nor U29297 (N_29297,N_29001,N_29154);
and U29298 (N_29298,N_29042,N_29194);
nor U29299 (N_29299,N_29067,N_29151);
nand U29300 (N_29300,N_29012,N_29121);
xor U29301 (N_29301,N_29031,N_29088);
and U29302 (N_29302,N_29053,N_29155);
xnor U29303 (N_29303,N_29066,N_29106);
or U29304 (N_29304,N_29094,N_29115);
and U29305 (N_29305,N_29075,N_29108);
nor U29306 (N_29306,N_29177,N_29062);
or U29307 (N_29307,N_29060,N_29118);
and U29308 (N_29308,N_29128,N_29111);
xnor U29309 (N_29309,N_29144,N_29050);
nor U29310 (N_29310,N_29122,N_29021);
nor U29311 (N_29311,N_29121,N_29109);
or U29312 (N_29312,N_29014,N_29179);
and U29313 (N_29313,N_29159,N_29098);
or U29314 (N_29314,N_29052,N_29033);
nand U29315 (N_29315,N_29130,N_29023);
or U29316 (N_29316,N_29080,N_29168);
nor U29317 (N_29317,N_29080,N_29035);
and U29318 (N_29318,N_29018,N_29088);
nand U29319 (N_29319,N_29124,N_29027);
nand U29320 (N_29320,N_29141,N_29071);
or U29321 (N_29321,N_29143,N_29183);
xnor U29322 (N_29322,N_29072,N_29084);
and U29323 (N_29323,N_29192,N_29104);
xnor U29324 (N_29324,N_29173,N_29141);
nor U29325 (N_29325,N_29114,N_29042);
nand U29326 (N_29326,N_29197,N_29196);
xor U29327 (N_29327,N_29105,N_29159);
nand U29328 (N_29328,N_29097,N_29191);
xnor U29329 (N_29329,N_29087,N_29098);
xnor U29330 (N_29330,N_29014,N_29148);
or U29331 (N_29331,N_29134,N_29178);
and U29332 (N_29332,N_29115,N_29018);
or U29333 (N_29333,N_29105,N_29009);
and U29334 (N_29334,N_29134,N_29168);
and U29335 (N_29335,N_29114,N_29054);
nor U29336 (N_29336,N_29129,N_29044);
nand U29337 (N_29337,N_29076,N_29023);
and U29338 (N_29338,N_29189,N_29114);
and U29339 (N_29339,N_29138,N_29058);
nand U29340 (N_29340,N_29179,N_29042);
and U29341 (N_29341,N_29117,N_29094);
nand U29342 (N_29342,N_29020,N_29000);
xor U29343 (N_29343,N_29195,N_29159);
nand U29344 (N_29344,N_29047,N_29120);
and U29345 (N_29345,N_29075,N_29148);
xnor U29346 (N_29346,N_29097,N_29107);
nor U29347 (N_29347,N_29188,N_29098);
and U29348 (N_29348,N_29064,N_29102);
or U29349 (N_29349,N_29060,N_29187);
xnor U29350 (N_29350,N_29178,N_29137);
or U29351 (N_29351,N_29106,N_29094);
nor U29352 (N_29352,N_29089,N_29044);
or U29353 (N_29353,N_29142,N_29063);
nand U29354 (N_29354,N_29000,N_29156);
xor U29355 (N_29355,N_29096,N_29113);
nor U29356 (N_29356,N_29102,N_29048);
and U29357 (N_29357,N_29004,N_29169);
or U29358 (N_29358,N_29162,N_29125);
xnor U29359 (N_29359,N_29039,N_29168);
nand U29360 (N_29360,N_29107,N_29021);
xnor U29361 (N_29361,N_29111,N_29060);
nand U29362 (N_29362,N_29045,N_29196);
nor U29363 (N_29363,N_29091,N_29179);
nor U29364 (N_29364,N_29100,N_29173);
xor U29365 (N_29365,N_29035,N_29000);
xor U29366 (N_29366,N_29059,N_29199);
nor U29367 (N_29367,N_29184,N_29100);
nor U29368 (N_29368,N_29077,N_29010);
or U29369 (N_29369,N_29019,N_29136);
nand U29370 (N_29370,N_29030,N_29013);
and U29371 (N_29371,N_29050,N_29148);
nand U29372 (N_29372,N_29126,N_29086);
xnor U29373 (N_29373,N_29172,N_29136);
nand U29374 (N_29374,N_29178,N_29194);
nand U29375 (N_29375,N_29073,N_29162);
and U29376 (N_29376,N_29040,N_29036);
nand U29377 (N_29377,N_29052,N_29030);
nand U29378 (N_29378,N_29001,N_29045);
or U29379 (N_29379,N_29081,N_29077);
nand U29380 (N_29380,N_29177,N_29090);
and U29381 (N_29381,N_29085,N_29170);
xor U29382 (N_29382,N_29116,N_29066);
or U29383 (N_29383,N_29072,N_29128);
nand U29384 (N_29384,N_29185,N_29195);
nand U29385 (N_29385,N_29151,N_29113);
xnor U29386 (N_29386,N_29039,N_29113);
nor U29387 (N_29387,N_29114,N_29086);
or U29388 (N_29388,N_29000,N_29111);
xor U29389 (N_29389,N_29099,N_29146);
or U29390 (N_29390,N_29093,N_29006);
nor U29391 (N_29391,N_29178,N_29177);
and U29392 (N_29392,N_29159,N_29129);
or U29393 (N_29393,N_29135,N_29186);
nor U29394 (N_29394,N_29039,N_29189);
or U29395 (N_29395,N_29043,N_29023);
or U29396 (N_29396,N_29057,N_29082);
or U29397 (N_29397,N_29190,N_29068);
xor U29398 (N_29398,N_29174,N_29140);
xor U29399 (N_29399,N_29194,N_29182);
and U29400 (N_29400,N_29234,N_29226);
nor U29401 (N_29401,N_29214,N_29329);
or U29402 (N_29402,N_29351,N_29233);
or U29403 (N_29403,N_29304,N_29279);
and U29404 (N_29404,N_29339,N_29349);
xnor U29405 (N_29405,N_29338,N_29385);
nand U29406 (N_29406,N_29227,N_29383);
nand U29407 (N_29407,N_29298,N_29330);
nor U29408 (N_29408,N_29312,N_29332);
xnor U29409 (N_29409,N_29259,N_29372);
nor U29410 (N_29410,N_29201,N_29391);
nor U29411 (N_29411,N_29296,N_29240);
and U29412 (N_29412,N_29366,N_29369);
nor U29413 (N_29413,N_29202,N_29311);
or U29414 (N_29414,N_29295,N_29356);
and U29415 (N_29415,N_29216,N_29337);
xnor U29416 (N_29416,N_29348,N_29245);
and U29417 (N_29417,N_29275,N_29260);
or U29418 (N_29418,N_29324,N_29255);
nand U29419 (N_29419,N_29297,N_29209);
and U29420 (N_29420,N_29381,N_29250);
xnor U29421 (N_29421,N_29359,N_29398);
and U29422 (N_29422,N_29328,N_29397);
nand U29423 (N_29423,N_29343,N_29310);
nand U29424 (N_29424,N_29253,N_29238);
nand U29425 (N_29425,N_29344,N_29283);
and U29426 (N_29426,N_29387,N_29321);
xor U29427 (N_29427,N_29284,N_29322);
and U29428 (N_29428,N_29352,N_29241);
xnor U29429 (N_29429,N_29292,N_29270);
nor U29430 (N_29430,N_29323,N_29257);
xor U29431 (N_29431,N_29247,N_29221);
nor U29432 (N_29432,N_29236,N_29293);
nor U29433 (N_29433,N_29389,N_29220);
or U29434 (N_29434,N_29217,N_29224);
nand U29435 (N_29435,N_29336,N_29318);
xnor U29436 (N_29436,N_29291,N_29365);
nand U29437 (N_29437,N_29347,N_29264);
nor U29438 (N_29438,N_29363,N_29263);
xnor U29439 (N_29439,N_29206,N_29205);
nand U29440 (N_29440,N_29314,N_29285);
nand U29441 (N_29441,N_29288,N_29392);
xor U29442 (N_29442,N_29305,N_29353);
or U29443 (N_29443,N_29340,N_29300);
and U29444 (N_29444,N_29213,N_29244);
nor U29445 (N_29445,N_29371,N_29273);
and U29446 (N_29446,N_29393,N_29327);
or U29447 (N_29447,N_29289,N_29341);
nand U29448 (N_29448,N_29333,N_29254);
xnor U29449 (N_29449,N_29281,N_29223);
nor U29450 (N_29450,N_29320,N_29361);
nand U29451 (N_29451,N_29390,N_29331);
and U29452 (N_29452,N_29350,N_29301);
xor U29453 (N_29453,N_29242,N_29265);
nor U29454 (N_29454,N_29267,N_29225);
nor U29455 (N_29455,N_29274,N_29294);
or U29456 (N_29456,N_29252,N_29222);
nand U29457 (N_29457,N_29268,N_29200);
nor U29458 (N_29458,N_29269,N_29290);
xor U29459 (N_29459,N_29382,N_29230);
and U29460 (N_29460,N_29282,N_29251);
nand U29461 (N_29461,N_29280,N_29218);
nor U29462 (N_29462,N_29335,N_29319);
nor U29463 (N_29463,N_29309,N_29307);
and U29464 (N_29464,N_29286,N_29326);
or U29465 (N_29465,N_29258,N_29266);
and U29466 (N_29466,N_29243,N_29278);
and U29467 (N_29467,N_29231,N_29203);
or U29468 (N_29468,N_29376,N_29210);
and U29469 (N_29469,N_29377,N_29364);
or U29470 (N_29470,N_29208,N_29207);
and U29471 (N_29471,N_29237,N_29211);
or U29472 (N_29472,N_29248,N_29261);
xor U29473 (N_29473,N_29373,N_29358);
xor U29474 (N_29474,N_29316,N_29362);
xnor U29475 (N_29475,N_29256,N_29396);
and U29476 (N_29476,N_29394,N_29239);
nor U29477 (N_29477,N_29215,N_29303);
nor U29478 (N_29478,N_29246,N_29379);
nand U29479 (N_29479,N_29346,N_29212);
and U29480 (N_29480,N_29308,N_29219);
or U29481 (N_29481,N_29262,N_29317);
or U29482 (N_29482,N_29287,N_29375);
nand U29483 (N_29483,N_29277,N_29342);
nor U29484 (N_29484,N_29374,N_29325);
and U29485 (N_29485,N_29315,N_29368);
xor U29486 (N_29486,N_29380,N_29235);
nor U29487 (N_29487,N_29272,N_29271);
or U29488 (N_29488,N_29384,N_29204);
nand U29489 (N_29489,N_29388,N_29299);
and U29490 (N_29490,N_29370,N_29229);
xnor U29491 (N_29491,N_29378,N_29355);
nand U29492 (N_29492,N_29395,N_29360);
or U29493 (N_29493,N_29232,N_29249);
or U29494 (N_29494,N_29354,N_29357);
xnor U29495 (N_29495,N_29367,N_29276);
xor U29496 (N_29496,N_29313,N_29228);
and U29497 (N_29497,N_29386,N_29399);
or U29498 (N_29498,N_29334,N_29306);
nand U29499 (N_29499,N_29345,N_29302);
xnor U29500 (N_29500,N_29204,N_29348);
nand U29501 (N_29501,N_29394,N_29206);
xnor U29502 (N_29502,N_29306,N_29305);
and U29503 (N_29503,N_29399,N_29301);
nor U29504 (N_29504,N_29240,N_29321);
nand U29505 (N_29505,N_29319,N_29302);
nor U29506 (N_29506,N_29371,N_29353);
and U29507 (N_29507,N_29279,N_29286);
nand U29508 (N_29508,N_29378,N_29220);
nor U29509 (N_29509,N_29375,N_29388);
or U29510 (N_29510,N_29231,N_29254);
nor U29511 (N_29511,N_29328,N_29364);
or U29512 (N_29512,N_29321,N_29262);
and U29513 (N_29513,N_29247,N_29389);
or U29514 (N_29514,N_29217,N_29243);
xor U29515 (N_29515,N_29268,N_29351);
xor U29516 (N_29516,N_29313,N_29223);
and U29517 (N_29517,N_29330,N_29365);
nand U29518 (N_29518,N_29235,N_29392);
nor U29519 (N_29519,N_29249,N_29239);
xor U29520 (N_29520,N_29360,N_29270);
or U29521 (N_29521,N_29325,N_29383);
nand U29522 (N_29522,N_29390,N_29357);
or U29523 (N_29523,N_29290,N_29297);
or U29524 (N_29524,N_29362,N_29306);
and U29525 (N_29525,N_29219,N_29329);
xor U29526 (N_29526,N_29322,N_29333);
xor U29527 (N_29527,N_29310,N_29391);
xor U29528 (N_29528,N_29280,N_29331);
nand U29529 (N_29529,N_29346,N_29318);
xnor U29530 (N_29530,N_29342,N_29359);
nand U29531 (N_29531,N_29215,N_29369);
xnor U29532 (N_29532,N_29335,N_29266);
or U29533 (N_29533,N_29329,N_29250);
or U29534 (N_29534,N_29217,N_29236);
nand U29535 (N_29535,N_29388,N_29255);
xnor U29536 (N_29536,N_29385,N_29282);
and U29537 (N_29537,N_29286,N_29261);
nor U29538 (N_29538,N_29246,N_29245);
and U29539 (N_29539,N_29249,N_29203);
nor U29540 (N_29540,N_29208,N_29379);
xor U29541 (N_29541,N_29292,N_29229);
nand U29542 (N_29542,N_29293,N_29210);
and U29543 (N_29543,N_29325,N_29321);
or U29544 (N_29544,N_29289,N_29252);
or U29545 (N_29545,N_29214,N_29270);
or U29546 (N_29546,N_29268,N_29253);
or U29547 (N_29547,N_29368,N_29310);
xor U29548 (N_29548,N_29305,N_29243);
nand U29549 (N_29549,N_29256,N_29348);
or U29550 (N_29550,N_29284,N_29358);
xnor U29551 (N_29551,N_29307,N_29323);
or U29552 (N_29552,N_29206,N_29264);
nor U29553 (N_29553,N_29288,N_29334);
or U29554 (N_29554,N_29235,N_29296);
or U29555 (N_29555,N_29274,N_29226);
xor U29556 (N_29556,N_29337,N_29237);
xor U29557 (N_29557,N_29354,N_29358);
nand U29558 (N_29558,N_29314,N_29301);
and U29559 (N_29559,N_29295,N_29303);
xnor U29560 (N_29560,N_29219,N_29330);
nand U29561 (N_29561,N_29353,N_29301);
or U29562 (N_29562,N_29322,N_29231);
or U29563 (N_29563,N_29372,N_29393);
and U29564 (N_29564,N_29252,N_29393);
xor U29565 (N_29565,N_29259,N_29285);
and U29566 (N_29566,N_29289,N_29306);
nor U29567 (N_29567,N_29387,N_29379);
nor U29568 (N_29568,N_29205,N_29343);
nand U29569 (N_29569,N_29226,N_29383);
nand U29570 (N_29570,N_29252,N_29314);
and U29571 (N_29571,N_29342,N_29357);
xnor U29572 (N_29572,N_29228,N_29338);
and U29573 (N_29573,N_29219,N_29298);
nand U29574 (N_29574,N_29298,N_29323);
xor U29575 (N_29575,N_29203,N_29258);
and U29576 (N_29576,N_29371,N_29305);
xor U29577 (N_29577,N_29250,N_29219);
nand U29578 (N_29578,N_29278,N_29318);
nand U29579 (N_29579,N_29349,N_29321);
and U29580 (N_29580,N_29282,N_29299);
nand U29581 (N_29581,N_29240,N_29204);
and U29582 (N_29582,N_29255,N_29244);
or U29583 (N_29583,N_29256,N_29389);
nand U29584 (N_29584,N_29200,N_29384);
nand U29585 (N_29585,N_29298,N_29204);
or U29586 (N_29586,N_29308,N_29256);
xor U29587 (N_29587,N_29234,N_29257);
xnor U29588 (N_29588,N_29253,N_29208);
nor U29589 (N_29589,N_29313,N_29330);
nor U29590 (N_29590,N_29368,N_29276);
xnor U29591 (N_29591,N_29215,N_29397);
and U29592 (N_29592,N_29306,N_29394);
or U29593 (N_29593,N_29312,N_29292);
and U29594 (N_29594,N_29251,N_29298);
nand U29595 (N_29595,N_29230,N_29397);
xnor U29596 (N_29596,N_29278,N_29331);
and U29597 (N_29597,N_29285,N_29358);
nand U29598 (N_29598,N_29339,N_29265);
and U29599 (N_29599,N_29248,N_29275);
or U29600 (N_29600,N_29529,N_29579);
or U29601 (N_29601,N_29571,N_29532);
and U29602 (N_29602,N_29415,N_29435);
or U29603 (N_29603,N_29487,N_29482);
or U29604 (N_29604,N_29462,N_29500);
nand U29605 (N_29605,N_29537,N_29510);
nor U29606 (N_29606,N_29596,N_29432);
xnor U29607 (N_29607,N_29502,N_29599);
or U29608 (N_29608,N_29468,N_29454);
nor U29609 (N_29609,N_29551,N_29485);
or U29610 (N_29610,N_29550,N_29452);
and U29611 (N_29611,N_29536,N_29554);
nand U29612 (N_29612,N_29507,N_29541);
xnor U29613 (N_29613,N_29408,N_29506);
and U29614 (N_29614,N_29475,N_29509);
and U29615 (N_29615,N_29456,N_29401);
nor U29616 (N_29616,N_29497,N_29520);
nand U29617 (N_29617,N_29548,N_29543);
xnor U29618 (N_29618,N_29593,N_29442);
nand U29619 (N_29619,N_29441,N_29413);
nand U29620 (N_29620,N_29400,N_29528);
xor U29621 (N_29621,N_29463,N_29453);
nor U29622 (N_29622,N_29518,N_29527);
nor U29623 (N_29623,N_29498,N_29483);
xor U29624 (N_29624,N_29444,N_29531);
nand U29625 (N_29625,N_29594,N_29587);
nor U29626 (N_29626,N_29577,N_29557);
nor U29627 (N_29627,N_29414,N_29486);
nor U29628 (N_29628,N_29501,N_29575);
or U29629 (N_29629,N_29583,N_29553);
or U29630 (N_29630,N_29458,N_29445);
and U29631 (N_29631,N_29515,N_29581);
or U29632 (N_29632,N_29512,N_29546);
nand U29633 (N_29633,N_29410,N_29514);
nor U29634 (N_29634,N_29547,N_29451);
nand U29635 (N_29635,N_29565,N_29523);
xnor U29636 (N_29636,N_29406,N_29504);
xnor U29637 (N_29637,N_29484,N_29521);
or U29638 (N_29638,N_29404,N_29568);
xnor U29639 (N_29639,N_29459,N_29429);
nand U29640 (N_29640,N_29479,N_29480);
xnor U29641 (N_29641,N_29467,N_29461);
or U29642 (N_29642,N_29533,N_29574);
nand U29643 (N_29643,N_29490,N_29446);
xor U29644 (N_29644,N_29590,N_29427);
xnor U29645 (N_29645,N_29416,N_29465);
and U29646 (N_29646,N_29503,N_29505);
nor U29647 (N_29647,N_29477,N_29492);
and U29648 (N_29648,N_29496,N_29539);
xnor U29649 (N_29649,N_29585,N_29576);
nor U29650 (N_29650,N_29561,N_29582);
nor U29651 (N_29651,N_29438,N_29426);
and U29652 (N_29652,N_29597,N_29471);
or U29653 (N_29653,N_29567,N_29522);
xor U29654 (N_29654,N_29476,N_29556);
xor U29655 (N_29655,N_29455,N_29535);
nor U29656 (N_29656,N_29469,N_29544);
nor U29657 (N_29657,N_29472,N_29562);
or U29658 (N_29658,N_29508,N_29499);
and U29659 (N_29659,N_29434,N_29598);
xnor U29660 (N_29660,N_29552,N_29428);
or U29661 (N_29661,N_29489,N_29517);
nand U29662 (N_29662,N_29572,N_29491);
xnor U29663 (N_29663,N_29569,N_29560);
and U29664 (N_29664,N_29588,N_29423);
or U29665 (N_29665,N_29566,N_29589);
nand U29666 (N_29666,N_29481,N_29412);
xor U29667 (N_29667,N_29563,N_29542);
or U29668 (N_29668,N_29430,N_29433);
or U29669 (N_29669,N_29519,N_29586);
nand U29670 (N_29670,N_29470,N_29540);
nand U29671 (N_29671,N_29460,N_29447);
or U29672 (N_29672,N_29407,N_29448);
nand U29673 (N_29673,N_29573,N_29564);
nand U29674 (N_29674,N_29559,N_29403);
or U29675 (N_29675,N_29513,N_29534);
nor U29676 (N_29676,N_29443,N_29431);
nor U29677 (N_29677,N_29495,N_29402);
or U29678 (N_29678,N_29449,N_29516);
nor U29679 (N_29679,N_29419,N_29584);
nand U29680 (N_29680,N_29592,N_29545);
xnor U29681 (N_29681,N_29439,N_29420);
or U29682 (N_29682,N_29549,N_29457);
nor U29683 (N_29683,N_29422,N_29425);
nand U29684 (N_29684,N_29555,N_29450);
and U29685 (N_29685,N_29511,N_29409);
nand U29686 (N_29686,N_29421,N_29417);
xnor U29687 (N_29687,N_29524,N_29464);
and U29688 (N_29688,N_29526,N_29473);
xnor U29689 (N_29689,N_29440,N_29493);
nand U29690 (N_29690,N_29591,N_29578);
nor U29691 (N_29691,N_29525,N_29558);
xor U29692 (N_29692,N_29538,N_29405);
nor U29693 (N_29693,N_29494,N_29474);
or U29694 (N_29694,N_29530,N_29570);
xor U29695 (N_29695,N_29466,N_29411);
nor U29696 (N_29696,N_29424,N_29478);
nor U29697 (N_29697,N_29488,N_29595);
and U29698 (N_29698,N_29418,N_29580);
nor U29699 (N_29699,N_29437,N_29436);
xnor U29700 (N_29700,N_29472,N_29430);
nor U29701 (N_29701,N_29584,N_29527);
xnor U29702 (N_29702,N_29590,N_29461);
and U29703 (N_29703,N_29456,N_29437);
nor U29704 (N_29704,N_29413,N_29585);
or U29705 (N_29705,N_29414,N_29526);
nand U29706 (N_29706,N_29532,N_29463);
nor U29707 (N_29707,N_29489,N_29515);
xnor U29708 (N_29708,N_29590,N_29554);
and U29709 (N_29709,N_29437,N_29517);
nor U29710 (N_29710,N_29559,N_29448);
nand U29711 (N_29711,N_29532,N_29462);
nor U29712 (N_29712,N_29543,N_29587);
nand U29713 (N_29713,N_29401,N_29509);
xnor U29714 (N_29714,N_29503,N_29461);
or U29715 (N_29715,N_29492,N_29415);
xnor U29716 (N_29716,N_29468,N_29540);
xnor U29717 (N_29717,N_29538,N_29569);
xnor U29718 (N_29718,N_29505,N_29470);
nor U29719 (N_29719,N_29453,N_29550);
and U29720 (N_29720,N_29468,N_29559);
and U29721 (N_29721,N_29551,N_29523);
or U29722 (N_29722,N_29505,N_29558);
nand U29723 (N_29723,N_29500,N_29429);
nor U29724 (N_29724,N_29444,N_29448);
nor U29725 (N_29725,N_29542,N_29521);
and U29726 (N_29726,N_29438,N_29575);
nand U29727 (N_29727,N_29579,N_29590);
and U29728 (N_29728,N_29582,N_29539);
nand U29729 (N_29729,N_29579,N_29482);
xor U29730 (N_29730,N_29511,N_29498);
xor U29731 (N_29731,N_29482,N_29425);
nor U29732 (N_29732,N_29502,N_29504);
or U29733 (N_29733,N_29466,N_29587);
and U29734 (N_29734,N_29469,N_29464);
xor U29735 (N_29735,N_29581,N_29417);
xor U29736 (N_29736,N_29483,N_29568);
nand U29737 (N_29737,N_29400,N_29424);
xor U29738 (N_29738,N_29465,N_29594);
and U29739 (N_29739,N_29552,N_29599);
or U29740 (N_29740,N_29496,N_29404);
and U29741 (N_29741,N_29432,N_29486);
nand U29742 (N_29742,N_29597,N_29428);
xor U29743 (N_29743,N_29446,N_29439);
nor U29744 (N_29744,N_29569,N_29517);
nand U29745 (N_29745,N_29461,N_29505);
and U29746 (N_29746,N_29471,N_29409);
nand U29747 (N_29747,N_29402,N_29430);
nor U29748 (N_29748,N_29400,N_29436);
xnor U29749 (N_29749,N_29549,N_29445);
or U29750 (N_29750,N_29534,N_29483);
or U29751 (N_29751,N_29434,N_29588);
nand U29752 (N_29752,N_29507,N_29471);
or U29753 (N_29753,N_29573,N_29576);
xor U29754 (N_29754,N_29524,N_29402);
nand U29755 (N_29755,N_29466,N_29580);
and U29756 (N_29756,N_29517,N_29465);
or U29757 (N_29757,N_29431,N_29545);
and U29758 (N_29758,N_29418,N_29534);
or U29759 (N_29759,N_29404,N_29462);
or U29760 (N_29760,N_29566,N_29531);
or U29761 (N_29761,N_29408,N_29491);
nand U29762 (N_29762,N_29521,N_29446);
nor U29763 (N_29763,N_29482,N_29594);
xor U29764 (N_29764,N_29520,N_29504);
xnor U29765 (N_29765,N_29416,N_29586);
nor U29766 (N_29766,N_29526,N_29429);
nand U29767 (N_29767,N_29444,N_29451);
and U29768 (N_29768,N_29560,N_29483);
and U29769 (N_29769,N_29429,N_29440);
or U29770 (N_29770,N_29462,N_29489);
nor U29771 (N_29771,N_29532,N_29511);
xor U29772 (N_29772,N_29483,N_29422);
and U29773 (N_29773,N_29412,N_29560);
or U29774 (N_29774,N_29512,N_29408);
nor U29775 (N_29775,N_29418,N_29425);
or U29776 (N_29776,N_29527,N_29553);
and U29777 (N_29777,N_29462,N_29407);
or U29778 (N_29778,N_29525,N_29507);
or U29779 (N_29779,N_29411,N_29561);
nor U29780 (N_29780,N_29461,N_29511);
nor U29781 (N_29781,N_29449,N_29495);
nand U29782 (N_29782,N_29544,N_29405);
and U29783 (N_29783,N_29594,N_29596);
and U29784 (N_29784,N_29444,N_29453);
or U29785 (N_29785,N_29593,N_29482);
or U29786 (N_29786,N_29590,N_29485);
nor U29787 (N_29787,N_29498,N_29484);
xor U29788 (N_29788,N_29510,N_29435);
nor U29789 (N_29789,N_29474,N_29486);
and U29790 (N_29790,N_29530,N_29481);
and U29791 (N_29791,N_29498,N_29411);
xnor U29792 (N_29792,N_29420,N_29452);
nand U29793 (N_29793,N_29411,N_29456);
or U29794 (N_29794,N_29431,N_29435);
xnor U29795 (N_29795,N_29468,N_29424);
or U29796 (N_29796,N_29400,N_29506);
or U29797 (N_29797,N_29594,N_29534);
nor U29798 (N_29798,N_29412,N_29441);
or U29799 (N_29799,N_29516,N_29430);
or U29800 (N_29800,N_29762,N_29609);
xor U29801 (N_29801,N_29705,N_29698);
or U29802 (N_29802,N_29777,N_29786);
nor U29803 (N_29803,N_29793,N_29730);
nor U29804 (N_29804,N_29729,N_29714);
or U29805 (N_29805,N_29772,N_29709);
or U29806 (N_29806,N_29690,N_29677);
or U29807 (N_29807,N_29618,N_29656);
or U29808 (N_29808,N_29683,N_29684);
xnor U29809 (N_29809,N_29655,N_29608);
or U29810 (N_29810,N_29769,N_29695);
and U29811 (N_29811,N_29616,N_29724);
nand U29812 (N_29812,N_29667,N_29676);
and U29813 (N_29813,N_29693,N_29703);
nor U29814 (N_29814,N_29704,N_29672);
nand U29815 (N_29815,N_29715,N_29623);
and U29816 (N_29816,N_29645,N_29648);
xnor U29817 (N_29817,N_29750,N_29621);
nor U29818 (N_29818,N_29707,N_29642);
and U29819 (N_29819,N_29612,N_29658);
and U29820 (N_29820,N_29792,N_29706);
or U29821 (N_29821,N_29619,N_29652);
or U29822 (N_29822,N_29785,N_29751);
nor U29823 (N_29823,N_29637,N_29668);
nand U29824 (N_29824,N_29726,N_29691);
and U29825 (N_29825,N_29613,N_29789);
and U29826 (N_29826,N_29747,N_29727);
nand U29827 (N_29827,N_29687,N_29685);
nor U29828 (N_29828,N_29711,N_29630);
nor U29829 (N_29829,N_29610,N_29669);
or U29830 (N_29830,N_29733,N_29660);
or U29831 (N_29831,N_29788,N_29659);
xor U29832 (N_29832,N_29752,N_29775);
xnor U29833 (N_29833,N_29702,N_29761);
xor U29834 (N_29834,N_29634,N_29743);
nor U29835 (N_29835,N_29646,N_29620);
and U29836 (N_29836,N_29745,N_29746);
nor U29837 (N_29837,N_29717,N_29723);
nand U29838 (N_29838,N_29719,N_29631);
and U29839 (N_29839,N_29689,N_29649);
xnor U29840 (N_29840,N_29755,N_29657);
nand U29841 (N_29841,N_29661,N_29638);
xor U29842 (N_29842,N_29674,N_29765);
or U29843 (N_29843,N_29787,N_29712);
or U29844 (N_29844,N_29644,N_29688);
xor U29845 (N_29845,N_29636,N_29664);
nand U29846 (N_29846,N_29641,N_29611);
xor U29847 (N_29847,N_29678,N_29696);
nand U29848 (N_29848,N_29640,N_29754);
nor U29849 (N_29849,N_29662,N_29757);
xor U29850 (N_29850,N_29756,N_29605);
or U29851 (N_29851,N_29736,N_29795);
nand U29852 (N_29852,N_29758,N_29673);
nand U29853 (N_29853,N_29694,N_29654);
or U29854 (N_29854,N_29763,N_29679);
or U29855 (N_29855,N_29759,N_29783);
nand U29856 (N_29856,N_29774,N_29603);
xnor U29857 (N_29857,N_29606,N_29771);
nand U29858 (N_29858,N_29764,N_29778);
or U29859 (N_29859,N_29749,N_29602);
xnor U29860 (N_29860,N_29639,N_29735);
nor U29861 (N_29861,N_29713,N_29665);
and U29862 (N_29862,N_29737,N_29716);
and U29863 (N_29863,N_29692,N_29760);
nor U29864 (N_29864,N_29615,N_29797);
nand U29865 (N_29865,N_29701,N_29627);
or U29866 (N_29866,N_29790,N_29643);
nand U29867 (N_29867,N_29651,N_29770);
and U29868 (N_29868,N_29728,N_29784);
or U29869 (N_29869,N_29748,N_29614);
nor U29870 (N_29870,N_29731,N_29742);
nand U29871 (N_29871,N_29617,N_29607);
and U29872 (N_29872,N_29782,N_29601);
or U29873 (N_29873,N_29740,N_29779);
xnor U29874 (N_29874,N_29626,N_29734);
nor U29875 (N_29875,N_29738,N_29768);
nand U29876 (N_29876,N_29721,N_29624);
and U29877 (N_29877,N_29708,N_29650);
xnor U29878 (N_29878,N_29799,N_29622);
and U29879 (N_29879,N_29675,N_29633);
and U29880 (N_29880,N_29700,N_29710);
nor U29881 (N_29881,N_29681,N_29632);
xor U29882 (N_29882,N_29796,N_29604);
or U29883 (N_29883,N_29744,N_29718);
and U29884 (N_29884,N_29647,N_29722);
nor U29885 (N_29885,N_29725,N_29699);
nand U29886 (N_29886,N_29666,N_29628);
nand U29887 (N_29887,N_29780,N_29781);
nand U29888 (N_29888,N_29682,N_29670);
nor U29889 (N_29889,N_29720,N_29773);
nand U29890 (N_29890,N_29741,N_29794);
or U29891 (N_29891,N_29686,N_29776);
xor U29892 (N_29892,N_29732,N_29791);
or U29893 (N_29893,N_29767,N_29663);
nand U29894 (N_29894,N_29635,N_29680);
and U29895 (N_29895,N_29625,N_29653);
nand U29896 (N_29896,N_29697,N_29671);
or U29897 (N_29897,N_29798,N_29766);
and U29898 (N_29898,N_29629,N_29600);
nor U29899 (N_29899,N_29739,N_29753);
or U29900 (N_29900,N_29735,N_29614);
xor U29901 (N_29901,N_29723,N_29776);
xnor U29902 (N_29902,N_29717,N_29601);
nand U29903 (N_29903,N_29749,N_29786);
nand U29904 (N_29904,N_29754,N_29627);
nand U29905 (N_29905,N_29614,N_29701);
and U29906 (N_29906,N_29717,N_29790);
nor U29907 (N_29907,N_29786,N_29741);
xor U29908 (N_29908,N_29647,N_29798);
nand U29909 (N_29909,N_29745,N_29715);
nand U29910 (N_29910,N_29789,N_29609);
xor U29911 (N_29911,N_29613,N_29728);
nand U29912 (N_29912,N_29737,N_29778);
nand U29913 (N_29913,N_29757,N_29755);
xnor U29914 (N_29914,N_29644,N_29787);
or U29915 (N_29915,N_29757,N_29726);
nor U29916 (N_29916,N_29755,N_29651);
xor U29917 (N_29917,N_29650,N_29787);
nor U29918 (N_29918,N_29656,N_29707);
nor U29919 (N_29919,N_29738,N_29640);
and U29920 (N_29920,N_29723,N_29663);
and U29921 (N_29921,N_29644,N_29648);
nand U29922 (N_29922,N_29742,N_29639);
xor U29923 (N_29923,N_29678,N_29647);
nand U29924 (N_29924,N_29734,N_29680);
or U29925 (N_29925,N_29782,N_29609);
and U29926 (N_29926,N_29704,N_29608);
or U29927 (N_29927,N_29642,N_29792);
xnor U29928 (N_29928,N_29721,N_29608);
xnor U29929 (N_29929,N_29728,N_29748);
nand U29930 (N_29930,N_29731,N_29609);
and U29931 (N_29931,N_29770,N_29650);
xor U29932 (N_29932,N_29732,N_29653);
nor U29933 (N_29933,N_29659,N_29670);
or U29934 (N_29934,N_29775,N_29777);
nand U29935 (N_29935,N_29726,N_29778);
or U29936 (N_29936,N_29606,N_29603);
or U29937 (N_29937,N_29638,N_29740);
nor U29938 (N_29938,N_29724,N_29663);
or U29939 (N_29939,N_29679,N_29618);
or U29940 (N_29940,N_29608,N_29601);
or U29941 (N_29941,N_29690,N_29643);
and U29942 (N_29942,N_29788,N_29638);
and U29943 (N_29943,N_29609,N_29707);
and U29944 (N_29944,N_29683,N_29789);
nand U29945 (N_29945,N_29604,N_29788);
nor U29946 (N_29946,N_29612,N_29648);
nand U29947 (N_29947,N_29753,N_29686);
and U29948 (N_29948,N_29624,N_29729);
nor U29949 (N_29949,N_29721,N_29644);
nor U29950 (N_29950,N_29794,N_29633);
nand U29951 (N_29951,N_29711,N_29791);
nand U29952 (N_29952,N_29683,N_29608);
or U29953 (N_29953,N_29688,N_29775);
nor U29954 (N_29954,N_29643,N_29659);
and U29955 (N_29955,N_29725,N_29708);
xnor U29956 (N_29956,N_29678,N_29618);
or U29957 (N_29957,N_29703,N_29666);
and U29958 (N_29958,N_29643,N_29623);
and U29959 (N_29959,N_29732,N_29610);
nor U29960 (N_29960,N_29629,N_29756);
nor U29961 (N_29961,N_29789,N_29769);
and U29962 (N_29962,N_29777,N_29718);
and U29963 (N_29963,N_29668,N_29638);
and U29964 (N_29964,N_29639,N_29730);
and U29965 (N_29965,N_29753,N_29736);
xnor U29966 (N_29966,N_29666,N_29689);
nor U29967 (N_29967,N_29726,N_29697);
or U29968 (N_29968,N_29660,N_29669);
and U29969 (N_29969,N_29646,N_29723);
xnor U29970 (N_29970,N_29607,N_29713);
nand U29971 (N_29971,N_29686,N_29761);
nand U29972 (N_29972,N_29635,N_29637);
and U29973 (N_29973,N_29775,N_29702);
or U29974 (N_29974,N_29726,N_29705);
nor U29975 (N_29975,N_29644,N_29614);
xnor U29976 (N_29976,N_29737,N_29671);
nor U29977 (N_29977,N_29614,N_29771);
nand U29978 (N_29978,N_29693,N_29686);
and U29979 (N_29979,N_29620,N_29722);
nor U29980 (N_29980,N_29746,N_29611);
or U29981 (N_29981,N_29715,N_29792);
xor U29982 (N_29982,N_29675,N_29724);
nand U29983 (N_29983,N_29751,N_29734);
or U29984 (N_29984,N_29756,N_29667);
or U29985 (N_29985,N_29604,N_29666);
nand U29986 (N_29986,N_29782,N_29773);
or U29987 (N_29987,N_29685,N_29666);
nand U29988 (N_29988,N_29759,N_29764);
xor U29989 (N_29989,N_29641,N_29637);
and U29990 (N_29990,N_29786,N_29778);
nor U29991 (N_29991,N_29749,N_29765);
and U29992 (N_29992,N_29758,N_29672);
or U29993 (N_29993,N_29781,N_29793);
nand U29994 (N_29994,N_29721,N_29716);
nor U29995 (N_29995,N_29633,N_29605);
nand U29996 (N_29996,N_29763,N_29744);
and U29997 (N_29997,N_29608,N_29706);
nand U29998 (N_29998,N_29763,N_29701);
xor U29999 (N_29999,N_29765,N_29626);
nor UO_0 (O_0,N_29919,N_29833);
nor UO_1 (O_1,N_29868,N_29858);
nor UO_2 (O_2,N_29977,N_29986);
and UO_3 (O_3,N_29872,N_29918);
or UO_4 (O_4,N_29997,N_29839);
xor UO_5 (O_5,N_29812,N_29963);
xnor UO_6 (O_6,N_29821,N_29865);
xnor UO_7 (O_7,N_29826,N_29827);
xor UO_8 (O_8,N_29804,N_29916);
or UO_9 (O_9,N_29859,N_29990);
or UO_10 (O_10,N_29863,N_29896);
and UO_11 (O_11,N_29964,N_29874);
xnor UO_12 (O_12,N_29803,N_29862);
xor UO_13 (O_13,N_29974,N_29835);
nor UO_14 (O_14,N_29973,N_29851);
or UO_15 (O_15,N_29917,N_29840);
nor UO_16 (O_16,N_29985,N_29817);
xnor UO_17 (O_17,N_29956,N_29807);
nor UO_18 (O_18,N_29908,N_29824);
and UO_19 (O_19,N_29879,N_29932);
nand UO_20 (O_20,N_29888,N_29993);
and UO_21 (O_21,N_29836,N_29837);
nor UO_22 (O_22,N_29884,N_29909);
nand UO_23 (O_23,N_29819,N_29971);
nand UO_24 (O_24,N_29999,N_29900);
and UO_25 (O_25,N_29844,N_29915);
and UO_26 (O_26,N_29968,N_29950);
nor UO_27 (O_27,N_29843,N_29982);
nor UO_28 (O_28,N_29972,N_29853);
and UO_29 (O_29,N_29922,N_29887);
xor UO_30 (O_30,N_29806,N_29924);
nor UO_31 (O_31,N_29962,N_29861);
and UO_32 (O_32,N_29912,N_29944);
and UO_33 (O_33,N_29866,N_29903);
xnor UO_34 (O_34,N_29953,N_29805);
or UO_35 (O_35,N_29829,N_29845);
or UO_36 (O_36,N_29847,N_29966);
nand UO_37 (O_37,N_29869,N_29931);
nand UO_38 (O_38,N_29808,N_29907);
nor UO_39 (O_39,N_29855,N_29846);
nand UO_40 (O_40,N_29929,N_29957);
nor UO_41 (O_41,N_29942,N_29969);
xor UO_42 (O_42,N_29961,N_29889);
nand UO_43 (O_43,N_29975,N_29838);
xnor UO_44 (O_44,N_29867,N_29935);
nor UO_45 (O_45,N_29832,N_29885);
xnor UO_46 (O_46,N_29981,N_29893);
and UO_47 (O_47,N_29938,N_29979);
and UO_48 (O_48,N_29860,N_29923);
and UO_49 (O_49,N_29927,N_29864);
and UO_50 (O_50,N_29989,N_29800);
and UO_51 (O_51,N_29914,N_29801);
or UO_52 (O_52,N_29959,N_29877);
or UO_53 (O_53,N_29992,N_29820);
nand UO_54 (O_54,N_29823,N_29928);
or UO_55 (O_55,N_29876,N_29899);
nand UO_56 (O_56,N_29849,N_29978);
nor UO_57 (O_57,N_29960,N_29842);
xnor UO_58 (O_58,N_29822,N_29983);
nand UO_59 (O_59,N_29892,N_29949);
nand UO_60 (O_60,N_29848,N_29911);
xnor UO_61 (O_61,N_29818,N_29873);
nor UO_62 (O_62,N_29815,N_29967);
and UO_63 (O_63,N_29948,N_29926);
or UO_64 (O_64,N_29882,N_29905);
and UO_65 (O_65,N_29886,N_29947);
xor UO_66 (O_66,N_29991,N_29952);
xor UO_67 (O_67,N_29883,N_29902);
nor UO_68 (O_68,N_29878,N_29894);
xor UO_69 (O_69,N_29813,N_29897);
and UO_70 (O_70,N_29870,N_29910);
or UO_71 (O_71,N_29834,N_29841);
nor UO_72 (O_72,N_29831,N_29939);
or UO_73 (O_73,N_29987,N_29994);
or UO_74 (O_74,N_29891,N_29921);
or UO_75 (O_75,N_29925,N_29995);
nand UO_76 (O_76,N_29998,N_29936);
xnor UO_77 (O_77,N_29828,N_29970);
xnor UO_78 (O_78,N_29830,N_29996);
xor UO_79 (O_79,N_29898,N_29920);
nor UO_80 (O_80,N_29940,N_29941);
or UO_81 (O_81,N_29954,N_29854);
xor UO_82 (O_82,N_29930,N_29856);
or UO_83 (O_83,N_29937,N_29814);
and UO_84 (O_84,N_29875,N_29880);
and UO_85 (O_85,N_29895,N_29825);
or UO_86 (O_86,N_29871,N_29946);
or UO_87 (O_87,N_29976,N_29852);
nor UO_88 (O_88,N_29984,N_29901);
or UO_89 (O_89,N_29810,N_29958);
nand UO_90 (O_90,N_29850,N_29934);
nand UO_91 (O_91,N_29955,N_29943);
or UO_92 (O_92,N_29980,N_29913);
xnor UO_93 (O_93,N_29857,N_29816);
and UO_94 (O_94,N_29890,N_29988);
nor UO_95 (O_95,N_29881,N_29811);
nand UO_96 (O_96,N_29802,N_29906);
or UO_97 (O_97,N_29951,N_29809);
nand UO_98 (O_98,N_29933,N_29904);
nor UO_99 (O_99,N_29945,N_29965);
nor UO_100 (O_100,N_29850,N_29941);
nor UO_101 (O_101,N_29806,N_29963);
or UO_102 (O_102,N_29820,N_29999);
nor UO_103 (O_103,N_29998,N_29953);
and UO_104 (O_104,N_29828,N_29853);
nor UO_105 (O_105,N_29865,N_29822);
and UO_106 (O_106,N_29880,N_29889);
xnor UO_107 (O_107,N_29944,N_29801);
nand UO_108 (O_108,N_29929,N_29888);
or UO_109 (O_109,N_29849,N_29922);
or UO_110 (O_110,N_29850,N_29936);
nand UO_111 (O_111,N_29891,N_29812);
or UO_112 (O_112,N_29953,N_29845);
and UO_113 (O_113,N_29948,N_29913);
and UO_114 (O_114,N_29815,N_29982);
and UO_115 (O_115,N_29919,N_29890);
xnor UO_116 (O_116,N_29957,N_29890);
xnor UO_117 (O_117,N_29879,N_29937);
or UO_118 (O_118,N_29882,N_29868);
or UO_119 (O_119,N_29878,N_29879);
and UO_120 (O_120,N_29908,N_29927);
xnor UO_121 (O_121,N_29805,N_29916);
or UO_122 (O_122,N_29835,N_29946);
xor UO_123 (O_123,N_29892,N_29916);
or UO_124 (O_124,N_29879,N_29890);
and UO_125 (O_125,N_29906,N_29854);
nand UO_126 (O_126,N_29985,N_29806);
or UO_127 (O_127,N_29842,N_29899);
and UO_128 (O_128,N_29878,N_29986);
xor UO_129 (O_129,N_29970,N_29904);
nand UO_130 (O_130,N_29822,N_29834);
nand UO_131 (O_131,N_29866,N_29958);
nand UO_132 (O_132,N_29941,N_29820);
and UO_133 (O_133,N_29964,N_29911);
or UO_134 (O_134,N_29974,N_29908);
nand UO_135 (O_135,N_29900,N_29997);
or UO_136 (O_136,N_29948,N_29819);
nand UO_137 (O_137,N_29877,N_29833);
nor UO_138 (O_138,N_29811,N_29847);
nor UO_139 (O_139,N_29921,N_29936);
nand UO_140 (O_140,N_29939,N_29849);
nor UO_141 (O_141,N_29886,N_29985);
or UO_142 (O_142,N_29879,N_29917);
or UO_143 (O_143,N_29954,N_29908);
and UO_144 (O_144,N_29917,N_29825);
nand UO_145 (O_145,N_29913,N_29869);
and UO_146 (O_146,N_29908,N_29940);
xor UO_147 (O_147,N_29915,N_29806);
and UO_148 (O_148,N_29837,N_29887);
or UO_149 (O_149,N_29807,N_29868);
nand UO_150 (O_150,N_29964,N_29991);
nand UO_151 (O_151,N_29853,N_29821);
nor UO_152 (O_152,N_29901,N_29970);
or UO_153 (O_153,N_29905,N_29959);
and UO_154 (O_154,N_29861,N_29834);
and UO_155 (O_155,N_29917,N_29990);
and UO_156 (O_156,N_29825,N_29887);
nor UO_157 (O_157,N_29989,N_29883);
nand UO_158 (O_158,N_29817,N_29967);
xnor UO_159 (O_159,N_29991,N_29926);
xor UO_160 (O_160,N_29937,N_29980);
xnor UO_161 (O_161,N_29923,N_29984);
or UO_162 (O_162,N_29859,N_29942);
or UO_163 (O_163,N_29978,N_29861);
nor UO_164 (O_164,N_29995,N_29938);
xor UO_165 (O_165,N_29922,N_29933);
xnor UO_166 (O_166,N_29918,N_29902);
or UO_167 (O_167,N_29973,N_29831);
and UO_168 (O_168,N_29857,N_29921);
xnor UO_169 (O_169,N_29917,N_29937);
or UO_170 (O_170,N_29928,N_29801);
xor UO_171 (O_171,N_29935,N_29975);
and UO_172 (O_172,N_29805,N_29946);
nor UO_173 (O_173,N_29896,N_29968);
xor UO_174 (O_174,N_29918,N_29840);
xor UO_175 (O_175,N_29808,N_29955);
xnor UO_176 (O_176,N_29999,N_29963);
xor UO_177 (O_177,N_29896,N_29819);
and UO_178 (O_178,N_29836,N_29933);
and UO_179 (O_179,N_29800,N_29812);
nand UO_180 (O_180,N_29890,N_29972);
xor UO_181 (O_181,N_29932,N_29923);
nor UO_182 (O_182,N_29896,N_29841);
nor UO_183 (O_183,N_29895,N_29995);
nand UO_184 (O_184,N_29850,N_29826);
xor UO_185 (O_185,N_29998,N_29900);
or UO_186 (O_186,N_29800,N_29903);
and UO_187 (O_187,N_29887,N_29976);
and UO_188 (O_188,N_29851,N_29908);
nand UO_189 (O_189,N_29996,N_29962);
xor UO_190 (O_190,N_29871,N_29901);
or UO_191 (O_191,N_29999,N_29961);
xnor UO_192 (O_192,N_29975,N_29978);
or UO_193 (O_193,N_29948,N_29866);
nor UO_194 (O_194,N_29960,N_29879);
xnor UO_195 (O_195,N_29977,N_29905);
nor UO_196 (O_196,N_29821,N_29881);
xor UO_197 (O_197,N_29969,N_29885);
and UO_198 (O_198,N_29919,N_29914);
nand UO_199 (O_199,N_29830,N_29975);
and UO_200 (O_200,N_29848,N_29939);
nor UO_201 (O_201,N_29854,N_29812);
nand UO_202 (O_202,N_29926,N_29993);
xor UO_203 (O_203,N_29967,N_29968);
nand UO_204 (O_204,N_29964,N_29834);
nor UO_205 (O_205,N_29827,N_29840);
and UO_206 (O_206,N_29926,N_29902);
xnor UO_207 (O_207,N_29964,N_29902);
xor UO_208 (O_208,N_29990,N_29983);
or UO_209 (O_209,N_29927,N_29858);
nand UO_210 (O_210,N_29942,N_29847);
nand UO_211 (O_211,N_29830,N_29898);
nor UO_212 (O_212,N_29812,N_29840);
and UO_213 (O_213,N_29918,N_29906);
or UO_214 (O_214,N_29959,N_29906);
or UO_215 (O_215,N_29868,N_29910);
or UO_216 (O_216,N_29874,N_29938);
or UO_217 (O_217,N_29908,N_29800);
xor UO_218 (O_218,N_29995,N_29813);
nor UO_219 (O_219,N_29965,N_29930);
or UO_220 (O_220,N_29806,N_29811);
and UO_221 (O_221,N_29928,N_29937);
and UO_222 (O_222,N_29992,N_29972);
and UO_223 (O_223,N_29918,N_29834);
or UO_224 (O_224,N_29878,N_29848);
or UO_225 (O_225,N_29873,N_29970);
nand UO_226 (O_226,N_29918,N_29919);
nor UO_227 (O_227,N_29812,N_29873);
or UO_228 (O_228,N_29905,N_29851);
and UO_229 (O_229,N_29914,N_29964);
or UO_230 (O_230,N_29832,N_29884);
nand UO_231 (O_231,N_29979,N_29929);
xnor UO_232 (O_232,N_29916,N_29954);
and UO_233 (O_233,N_29851,N_29871);
nand UO_234 (O_234,N_29927,N_29926);
nand UO_235 (O_235,N_29940,N_29999);
xnor UO_236 (O_236,N_29869,N_29919);
nand UO_237 (O_237,N_29907,N_29980);
nor UO_238 (O_238,N_29811,N_29920);
and UO_239 (O_239,N_29851,N_29916);
nor UO_240 (O_240,N_29895,N_29954);
nand UO_241 (O_241,N_29822,N_29909);
nor UO_242 (O_242,N_29893,N_29904);
or UO_243 (O_243,N_29914,N_29957);
xnor UO_244 (O_244,N_29978,N_29973);
xnor UO_245 (O_245,N_29834,N_29917);
nor UO_246 (O_246,N_29917,N_29827);
nand UO_247 (O_247,N_29861,N_29851);
nand UO_248 (O_248,N_29832,N_29829);
or UO_249 (O_249,N_29840,N_29922);
or UO_250 (O_250,N_29973,N_29999);
or UO_251 (O_251,N_29955,N_29825);
or UO_252 (O_252,N_29829,N_29945);
and UO_253 (O_253,N_29868,N_29812);
nand UO_254 (O_254,N_29963,N_29905);
nand UO_255 (O_255,N_29935,N_29854);
nand UO_256 (O_256,N_29919,N_29924);
nand UO_257 (O_257,N_29895,N_29951);
nor UO_258 (O_258,N_29883,N_29884);
nor UO_259 (O_259,N_29896,N_29852);
or UO_260 (O_260,N_29961,N_29946);
or UO_261 (O_261,N_29888,N_29957);
and UO_262 (O_262,N_29883,N_29821);
nor UO_263 (O_263,N_29898,N_29919);
or UO_264 (O_264,N_29831,N_29985);
and UO_265 (O_265,N_29983,N_29805);
and UO_266 (O_266,N_29907,N_29922);
or UO_267 (O_267,N_29939,N_29979);
and UO_268 (O_268,N_29945,N_29825);
nor UO_269 (O_269,N_29896,N_29950);
xnor UO_270 (O_270,N_29970,N_29858);
or UO_271 (O_271,N_29892,N_29812);
nor UO_272 (O_272,N_29986,N_29804);
nand UO_273 (O_273,N_29956,N_29952);
nand UO_274 (O_274,N_29815,N_29858);
xnor UO_275 (O_275,N_29971,N_29889);
and UO_276 (O_276,N_29933,N_29886);
and UO_277 (O_277,N_29947,N_29989);
xor UO_278 (O_278,N_29801,N_29883);
or UO_279 (O_279,N_29836,N_29826);
and UO_280 (O_280,N_29949,N_29868);
nand UO_281 (O_281,N_29882,N_29864);
nand UO_282 (O_282,N_29977,N_29899);
nand UO_283 (O_283,N_29874,N_29888);
nand UO_284 (O_284,N_29933,N_29998);
nor UO_285 (O_285,N_29999,N_29833);
nand UO_286 (O_286,N_29934,N_29800);
or UO_287 (O_287,N_29872,N_29983);
and UO_288 (O_288,N_29921,N_29925);
nor UO_289 (O_289,N_29911,N_29937);
xnor UO_290 (O_290,N_29852,N_29802);
xor UO_291 (O_291,N_29854,N_29805);
xor UO_292 (O_292,N_29817,N_29959);
xor UO_293 (O_293,N_29850,N_29981);
and UO_294 (O_294,N_29954,N_29975);
xor UO_295 (O_295,N_29898,N_29996);
nor UO_296 (O_296,N_29853,N_29995);
and UO_297 (O_297,N_29862,N_29902);
xnor UO_298 (O_298,N_29867,N_29886);
nor UO_299 (O_299,N_29827,N_29965);
nand UO_300 (O_300,N_29851,N_29829);
nor UO_301 (O_301,N_29831,N_29930);
nand UO_302 (O_302,N_29856,N_29956);
nand UO_303 (O_303,N_29897,N_29891);
nor UO_304 (O_304,N_29941,N_29881);
or UO_305 (O_305,N_29971,N_29904);
nand UO_306 (O_306,N_29874,N_29919);
nand UO_307 (O_307,N_29842,N_29945);
nor UO_308 (O_308,N_29852,N_29850);
nor UO_309 (O_309,N_29852,N_29876);
xor UO_310 (O_310,N_29846,N_29913);
nand UO_311 (O_311,N_29879,N_29979);
xor UO_312 (O_312,N_29915,N_29841);
or UO_313 (O_313,N_29921,N_29875);
xnor UO_314 (O_314,N_29806,N_29908);
xnor UO_315 (O_315,N_29835,N_29823);
nor UO_316 (O_316,N_29902,N_29936);
or UO_317 (O_317,N_29800,N_29888);
xnor UO_318 (O_318,N_29879,N_29812);
nand UO_319 (O_319,N_29837,N_29999);
nand UO_320 (O_320,N_29803,N_29972);
nor UO_321 (O_321,N_29814,N_29982);
xor UO_322 (O_322,N_29892,N_29826);
and UO_323 (O_323,N_29915,N_29962);
nor UO_324 (O_324,N_29866,N_29957);
xnor UO_325 (O_325,N_29851,N_29800);
xor UO_326 (O_326,N_29907,N_29852);
nand UO_327 (O_327,N_29992,N_29940);
nor UO_328 (O_328,N_29960,N_29853);
xor UO_329 (O_329,N_29882,N_29941);
and UO_330 (O_330,N_29931,N_29936);
nand UO_331 (O_331,N_29991,N_29815);
nor UO_332 (O_332,N_29821,N_29886);
nor UO_333 (O_333,N_29803,N_29898);
or UO_334 (O_334,N_29965,N_29889);
nor UO_335 (O_335,N_29939,N_29821);
nand UO_336 (O_336,N_29868,N_29863);
and UO_337 (O_337,N_29848,N_29970);
nand UO_338 (O_338,N_29826,N_29977);
and UO_339 (O_339,N_29889,N_29898);
and UO_340 (O_340,N_29927,N_29896);
nand UO_341 (O_341,N_29848,N_29917);
nor UO_342 (O_342,N_29851,N_29913);
or UO_343 (O_343,N_29807,N_29947);
or UO_344 (O_344,N_29915,N_29830);
and UO_345 (O_345,N_29941,N_29883);
nand UO_346 (O_346,N_29872,N_29942);
and UO_347 (O_347,N_29980,N_29867);
and UO_348 (O_348,N_29934,N_29919);
nor UO_349 (O_349,N_29850,N_29957);
nand UO_350 (O_350,N_29979,N_29875);
nand UO_351 (O_351,N_29898,N_29870);
and UO_352 (O_352,N_29816,N_29962);
xor UO_353 (O_353,N_29992,N_29981);
nand UO_354 (O_354,N_29955,N_29906);
xor UO_355 (O_355,N_29853,N_29926);
and UO_356 (O_356,N_29803,N_29920);
and UO_357 (O_357,N_29941,N_29833);
or UO_358 (O_358,N_29879,N_29805);
nand UO_359 (O_359,N_29937,N_29939);
nor UO_360 (O_360,N_29804,N_29919);
xnor UO_361 (O_361,N_29987,N_29906);
and UO_362 (O_362,N_29967,N_29923);
or UO_363 (O_363,N_29860,N_29854);
nor UO_364 (O_364,N_29973,N_29845);
xor UO_365 (O_365,N_29913,N_29888);
nand UO_366 (O_366,N_29829,N_29984);
nand UO_367 (O_367,N_29875,N_29897);
and UO_368 (O_368,N_29863,N_29812);
nor UO_369 (O_369,N_29959,N_29937);
or UO_370 (O_370,N_29939,N_29971);
xor UO_371 (O_371,N_29898,N_29875);
nor UO_372 (O_372,N_29894,N_29980);
nand UO_373 (O_373,N_29864,N_29966);
nand UO_374 (O_374,N_29841,N_29851);
and UO_375 (O_375,N_29873,N_29822);
and UO_376 (O_376,N_29829,N_29815);
and UO_377 (O_377,N_29987,N_29867);
xnor UO_378 (O_378,N_29949,N_29843);
nand UO_379 (O_379,N_29964,N_29891);
nor UO_380 (O_380,N_29936,N_29811);
xor UO_381 (O_381,N_29876,N_29900);
and UO_382 (O_382,N_29900,N_29813);
or UO_383 (O_383,N_29830,N_29952);
nand UO_384 (O_384,N_29908,N_29837);
nor UO_385 (O_385,N_29917,N_29841);
or UO_386 (O_386,N_29871,N_29958);
or UO_387 (O_387,N_29955,N_29853);
xor UO_388 (O_388,N_29882,N_29946);
nand UO_389 (O_389,N_29907,N_29961);
and UO_390 (O_390,N_29833,N_29952);
and UO_391 (O_391,N_29977,N_29908);
or UO_392 (O_392,N_29805,N_29943);
xnor UO_393 (O_393,N_29822,N_29963);
or UO_394 (O_394,N_29971,N_29991);
and UO_395 (O_395,N_29947,N_29801);
or UO_396 (O_396,N_29905,N_29844);
xnor UO_397 (O_397,N_29988,N_29820);
and UO_398 (O_398,N_29849,N_29942);
nand UO_399 (O_399,N_29892,N_29894);
and UO_400 (O_400,N_29934,N_29993);
nand UO_401 (O_401,N_29957,N_29810);
or UO_402 (O_402,N_29923,N_29995);
nor UO_403 (O_403,N_29824,N_29811);
xnor UO_404 (O_404,N_29992,N_29970);
nor UO_405 (O_405,N_29951,N_29947);
nor UO_406 (O_406,N_29986,N_29964);
and UO_407 (O_407,N_29997,N_29802);
and UO_408 (O_408,N_29830,N_29859);
nand UO_409 (O_409,N_29950,N_29921);
nor UO_410 (O_410,N_29940,N_29961);
or UO_411 (O_411,N_29869,N_29871);
nand UO_412 (O_412,N_29857,N_29990);
or UO_413 (O_413,N_29885,N_29821);
and UO_414 (O_414,N_29957,N_29804);
nor UO_415 (O_415,N_29889,N_29829);
nand UO_416 (O_416,N_29949,N_29836);
and UO_417 (O_417,N_29884,N_29941);
and UO_418 (O_418,N_29867,N_29849);
xor UO_419 (O_419,N_29831,N_29853);
xor UO_420 (O_420,N_29861,N_29864);
nand UO_421 (O_421,N_29937,N_29925);
or UO_422 (O_422,N_29851,N_29890);
nor UO_423 (O_423,N_29826,N_29854);
nand UO_424 (O_424,N_29814,N_29831);
xor UO_425 (O_425,N_29934,N_29848);
xnor UO_426 (O_426,N_29912,N_29922);
and UO_427 (O_427,N_29934,N_29925);
and UO_428 (O_428,N_29836,N_29891);
and UO_429 (O_429,N_29969,N_29815);
nor UO_430 (O_430,N_29902,N_29943);
and UO_431 (O_431,N_29898,N_29945);
nand UO_432 (O_432,N_29815,N_29837);
or UO_433 (O_433,N_29809,N_29802);
nor UO_434 (O_434,N_29816,N_29873);
nand UO_435 (O_435,N_29954,N_29900);
xor UO_436 (O_436,N_29872,N_29830);
nor UO_437 (O_437,N_29880,N_29838);
nand UO_438 (O_438,N_29821,N_29986);
or UO_439 (O_439,N_29914,N_29988);
and UO_440 (O_440,N_29907,N_29885);
xor UO_441 (O_441,N_29929,N_29995);
and UO_442 (O_442,N_29806,N_29880);
or UO_443 (O_443,N_29924,N_29890);
nand UO_444 (O_444,N_29992,N_29921);
and UO_445 (O_445,N_29946,N_29887);
xor UO_446 (O_446,N_29894,N_29974);
or UO_447 (O_447,N_29889,N_29943);
or UO_448 (O_448,N_29838,N_29908);
xnor UO_449 (O_449,N_29893,N_29978);
nor UO_450 (O_450,N_29810,N_29864);
nor UO_451 (O_451,N_29850,N_29854);
nor UO_452 (O_452,N_29802,N_29844);
nor UO_453 (O_453,N_29934,N_29834);
and UO_454 (O_454,N_29961,N_29971);
or UO_455 (O_455,N_29882,N_29896);
and UO_456 (O_456,N_29945,N_29812);
and UO_457 (O_457,N_29994,N_29859);
nand UO_458 (O_458,N_29920,N_29886);
and UO_459 (O_459,N_29834,N_29837);
nand UO_460 (O_460,N_29903,N_29978);
nand UO_461 (O_461,N_29932,N_29815);
nor UO_462 (O_462,N_29893,N_29840);
xor UO_463 (O_463,N_29819,N_29962);
xor UO_464 (O_464,N_29824,N_29900);
xnor UO_465 (O_465,N_29966,N_29976);
and UO_466 (O_466,N_29972,N_29979);
and UO_467 (O_467,N_29926,N_29987);
and UO_468 (O_468,N_29909,N_29814);
or UO_469 (O_469,N_29921,N_29837);
and UO_470 (O_470,N_29979,N_29989);
or UO_471 (O_471,N_29905,N_29862);
or UO_472 (O_472,N_29947,N_29908);
and UO_473 (O_473,N_29909,N_29992);
nor UO_474 (O_474,N_29839,N_29835);
xnor UO_475 (O_475,N_29882,N_29955);
or UO_476 (O_476,N_29923,N_29904);
xor UO_477 (O_477,N_29968,N_29972);
and UO_478 (O_478,N_29874,N_29863);
nand UO_479 (O_479,N_29838,N_29857);
xnor UO_480 (O_480,N_29907,N_29860);
and UO_481 (O_481,N_29861,N_29941);
and UO_482 (O_482,N_29911,N_29953);
or UO_483 (O_483,N_29986,N_29887);
xor UO_484 (O_484,N_29854,N_29835);
or UO_485 (O_485,N_29877,N_29818);
nand UO_486 (O_486,N_29845,N_29954);
and UO_487 (O_487,N_29813,N_29825);
or UO_488 (O_488,N_29878,N_29824);
and UO_489 (O_489,N_29857,N_29946);
nor UO_490 (O_490,N_29933,N_29999);
or UO_491 (O_491,N_29975,N_29940);
or UO_492 (O_492,N_29870,N_29922);
nor UO_493 (O_493,N_29885,N_29941);
or UO_494 (O_494,N_29828,N_29979);
and UO_495 (O_495,N_29803,N_29941);
nor UO_496 (O_496,N_29883,N_29828);
and UO_497 (O_497,N_29813,N_29914);
xnor UO_498 (O_498,N_29914,N_29909);
or UO_499 (O_499,N_29864,N_29904);
and UO_500 (O_500,N_29991,N_29902);
xor UO_501 (O_501,N_29884,N_29802);
xor UO_502 (O_502,N_29846,N_29862);
nand UO_503 (O_503,N_29819,N_29891);
or UO_504 (O_504,N_29865,N_29929);
or UO_505 (O_505,N_29864,N_29867);
nand UO_506 (O_506,N_29984,N_29909);
nand UO_507 (O_507,N_29818,N_29808);
nand UO_508 (O_508,N_29900,N_29962);
nand UO_509 (O_509,N_29825,N_29828);
and UO_510 (O_510,N_29879,N_29970);
xor UO_511 (O_511,N_29926,N_29888);
xor UO_512 (O_512,N_29910,N_29985);
or UO_513 (O_513,N_29977,N_29913);
xor UO_514 (O_514,N_29971,N_29852);
and UO_515 (O_515,N_29985,N_29984);
nor UO_516 (O_516,N_29835,N_29955);
nand UO_517 (O_517,N_29979,N_29984);
and UO_518 (O_518,N_29923,N_29826);
or UO_519 (O_519,N_29992,N_29923);
nand UO_520 (O_520,N_29876,N_29828);
nand UO_521 (O_521,N_29819,N_29909);
and UO_522 (O_522,N_29870,N_29846);
xnor UO_523 (O_523,N_29897,N_29882);
nand UO_524 (O_524,N_29937,N_29895);
xnor UO_525 (O_525,N_29830,N_29909);
xnor UO_526 (O_526,N_29858,N_29867);
nor UO_527 (O_527,N_29832,N_29820);
and UO_528 (O_528,N_29833,N_29940);
or UO_529 (O_529,N_29904,N_29813);
nor UO_530 (O_530,N_29923,N_29875);
or UO_531 (O_531,N_29958,N_29944);
nand UO_532 (O_532,N_29952,N_29992);
nand UO_533 (O_533,N_29900,N_29888);
nand UO_534 (O_534,N_29972,N_29807);
or UO_535 (O_535,N_29820,N_29858);
xor UO_536 (O_536,N_29860,N_29992);
xnor UO_537 (O_537,N_29961,N_29899);
xor UO_538 (O_538,N_29922,N_29950);
or UO_539 (O_539,N_29838,N_29832);
xor UO_540 (O_540,N_29934,N_29990);
nand UO_541 (O_541,N_29904,N_29937);
and UO_542 (O_542,N_29966,N_29865);
and UO_543 (O_543,N_29908,N_29867);
nor UO_544 (O_544,N_29904,N_29982);
or UO_545 (O_545,N_29824,N_29997);
nand UO_546 (O_546,N_29955,N_29830);
and UO_547 (O_547,N_29957,N_29988);
or UO_548 (O_548,N_29851,N_29835);
nand UO_549 (O_549,N_29903,N_29981);
nand UO_550 (O_550,N_29933,N_29926);
nor UO_551 (O_551,N_29864,N_29832);
xnor UO_552 (O_552,N_29822,N_29928);
xor UO_553 (O_553,N_29828,N_29965);
xor UO_554 (O_554,N_29921,N_29896);
nand UO_555 (O_555,N_29927,N_29840);
and UO_556 (O_556,N_29927,N_29938);
nand UO_557 (O_557,N_29858,N_29807);
or UO_558 (O_558,N_29818,N_29804);
xor UO_559 (O_559,N_29988,N_29909);
or UO_560 (O_560,N_29916,N_29870);
and UO_561 (O_561,N_29997,N_29831);
xor UO_562 (O_562,N_29923,N_29823);
nor UO_563 (O_563,N_29915,N_29803);
and UO_564 (O_564,N_29913,N_29840);
and UO_565 (O_565,N_29961,N_29882);
and UO_566 (O_566,N_29897,N_29923);
nand UO_567 (O_567,N_29818,N_29915);
or UO_568 (O_568,N_29833,N_29826);
and UO_569 (O_569,N_29978,N_29904);
or UO_570 (O_570,N_29833,N_29869);
or UO_571 (O_571,N_29892,N_29936);
nor UO_572 (O_572,N_29917,N_29821);
or UO_573 (O_573,N_29821,N_29859);
xor UO_574 (O_574,N_29932,N_29968);
or UO_575 (O_575,N_29985,N_29918);
and UO_576 (O_576,N_29819,N_29992);
and UO_577 (O_577,N_29828,N_29856);
xnor UO_578 (O_578,N_29871,N_29863);
nand UO_579 (O_579,N_29954,N_29949);
nand UO_580 (O_580,N_29913,N_29979);
nor UO_581 (O_581,N_29986,N_29976);
or UO_582 (O_582,N_29957,N_29851);
and UO_583 (O_583,N_29873,N_29831);
and UO_584 (O_584,N_29974,N_29810);
nor UO_585 (O_585,N_29806,N_29883);
or UO_586 (O_586,N_29896,N_29907);
xor UO_587 (O_587,N_29808,N_29947);
and UO_588 (O_588,N_29868,N_29835);
or UO_589 (O_589,N_29918,N_29959);
or UO_590 (O_590,N_29823,N_29855);
xor UO_591 (O_591,N_29825,N_29938);
and UO_592 (O_592,N_29909,N_29857);
xnor UO_593 (O_593,N_29867,N_29883);
nand UO_594 (O_594,N_29834,N_29859);
xor UO_595 (O_595,N_29932,N_29937);
nand UO_596 (O_596,N_29865,N_29998);
nor UO_597 (O_597,N_29894,N_29924);
nand UO_598 (O_598,N_29960,N_29984);
xor UO_599 (O_599,N_29974,N_29985);
or UO_600 (O_600,N_29821,N_29987);
nand UO_601 (O_601,N_29909,N_29974);
and UO_602 (O_602,N_29958,N_29884);
and UO_603 (O_603,N_29846,N_29977);
nand UO_604 (O_604,N_29964,N_29869);
nor UO_605 (O_605,N_29948,N_29816);
xnor UO_606 (O_606,N_29874,N_29900);
nand UO_607 (O_607,N_29811,N_29923);
and UO_608 (O_608,N_29805,N_29891);
nand UO_609 (O_609,N_29906,N_29840);
nand UO_610 (O_610,N_29910,N_29842);
and UO_611 (O_611,N_29975,N_29981);
nand UO_612 (O_612,N_29932,N_29870);
xor UO_613 (O_613,N_29963,N_29850);
nor UO_614 (O_614,N_29860,N_29931);
nand UO_615 (O_615,N_29963,N_29939);
and UO_616 (O_616,N_29942,N_29970);
xnor UO_617 (O_617,N_29924,N_29989);
xor UO_618 (O_618,N_29834,N_29997);
or UO_619 (O_619,N_29874,N_29969);
xor UO_620 (O_620,N_29903,N_29855);
nand UO_621 (O_621,N_29822,N_29969);
nor UO_622 (O_622,N_29830,N_29956);
or UO_623 (O_623,N_29846,N_29886);
nand UO_624 (O_624,N_29970,N_29969);
xor UO_625 (O_625,N_29808,N_29805);
xnor UO_626 (O_626,N_29825,N_29919);
or UO_627 (O_627,N_29870,N_29896);
or UO_628 (O_628,N_29996,N_29959);
nand UO_629 (O_629,N_29857,N_29947);
and UO_630 (O_630,N_29907,N_29877);
nor UO_631 (O_631,N_29858,N_29877);
nor UO_632 (O_632,N_29852,N_29829);
xnor UO_633 (O_633,N_29850,N_29894);
nor UO_634 (O_634,N_29977,N_29837);
or UO_635 (O_635,N_29975,N_29957);
nand UO_636 (O_636,N_29846,N_29984);
nand UO_637 (O_637,N_29916,N_29947);
nor UO_638 (O_638,N_29999,N_29871);
nand UO_639 (O_639,N_29924,N_29864);
or UO_640 (O_640,N_29940,N_29876);
xor UO_641 (O_641,N_29855,N_29816);
and UO_642 (O_642,N_29965,N_29873);
nand UO_643 (O_643,N_29982,N_29921);
and UO_644 (O_644,N_29943,N_29988);
and UO_645 (O_645,N_29966,N_29859);
and UO_646 (O_646,N_29824,N_29958);
xnor UO_647 (O_647,N_29909,N_29844);
nor UO_648 (O_648,N_29873,N_29937);
nor UO_649 (O_649,N_29983,N_29949);
nor UO_650 (O_650,N_29870,N_29967);
and UO_651 (O_651,N_29858,N_29906);
xor UO_652 (O_652,N_29969,N_29893);
and UO_653 (O_653,N_29978,N_29968);
nor UO_654 (O_654,N_29926,N_29838);
nand UO_655 (O_655,N_29852,N_29822);
nand UO_656 (O_656,N_29857,N_29934);
or UO_657 (O_657,N_29952,N_29940);
nand UO_658 (O_658,N_29882,N_29924);
nand UO_659 (O_659,N_29871,N_29840);
and UO_660 (O_660,N_29847,N_29957);
nand UO_661 (O_661,N_29818,N_29813);
nor UO_662 (O_662,N_29864,N_29945);
and UO_663 (O_663,N_29897,N_29880);
nand UO_664 (O_664,N_29830,N_29862);
nor UO_665 (O_665,N_29853,N_29943);
and UO_666 (O_666,N_29928,N_29941);
xor UO_667 (O_667,N_29818,N_29987);
nand UO_668 (O_668,N_29847,N_29947);
nor UO_669 (O_669,N_29894,N_29807);
nor UO_670 (O_670,N_29875,N_29819);
or UO_671 (O_671,N_29878,N_29829);
xor UO_672 (O_672,N_29820,N_29944);
xor UO_673 (O_673,N_29952,N_29960);
nor UO_674 (O_674,N_29949,N_29834);
nor UO_675 (O_675,N_29969,N_29827);
nand UO_676 (O_676,N_29874,N_29839);
nand UO_677 (O_677,N_29841,N_29975);
and UO_678 (O_678,N_29836,N_29931);
nor UO_679 (O_679,N_29825,N_29801);
nand UO_680 (O_680,N_29883,N_29948);
and UO_681 (O_681,N_29857,N_29996);
nand UO_682 (O_682,N_29928,N_29991);
and UO_683 (O_683,N_29851,N_29966);
and UO_684 (O_684,N_29934,N_29873);
nor UO_685 (O_685,N_29885,N_29888);
or UO_686 (O_686,N_29954,N_29938);
nor UO_687 (O_687,N_29941,N_29961);
and UO_688 (O_688,N_29964,N_29997);
or UO_689 (O_689,N_29856,N_29841);
xor UO_690 (O_690,N_29858,N_29918);
or UO_691 (O_691,N_29841,N_29883);
and UO_692 (O_692,N_29876,N_29845);
nand UO_693 (O_693,N_29969,N_29847);
and UO_694 (O_694,N_29956,N_29979);
and UO_695 (O_695,N_29900,N_29977);
and UO_696 (O_696,N_29819,N_29955);
xnor UO_697 (O_697,N_29930,N_29809);
and UO_698 (O_698,N_29891,N_29971);
nor UO_699 (O_699,N_29901,N_29982);
nor UO_700 (O_700,N_29846,N_29919);
and UO_701 (O_701,N_29999,N_29867);
or UO_702 (O_702,N_29999,N_29937);
nand UO_703 (O_703,N_29965,N_29915);
nor UO_704 (O_704,N_29832,N_29841);
nand UO_705 (O_705,N_29953,N_29924);
nor UO_706 (O_706,N_29907,N_29999);
or UO_707 (O_707,N_29902,N_29954);
nor UO_708 (O_708,N_29812,N_29836);
nor UO_709 (O_709,N_29913,N_29908);
nor UO_710 (O_710,N_29858,N_29893);
nor UO_711 (O_711,N_29810,N_29913);
or UO_712 (O_712,N_29973,N_29926);
nand UO_713 (O_713,N_29827,N_29813);
and UO_714 (O_714,N_29864,N_29990);
or UO_715 (O_715,N_29854,N_29823);
and UO_716 (O_716,N_29846,N_29986);
nor UO_717 (O_717,N_29902,N_29957);
xnor UO_718 (O_718,N_29817,N_29944);
and UO_719 (O_719,N_29807,N_29935);
nor UO_720 (O_720,N_29984,N_29952);
nor UO_721 (O_721,N_29840,N_29894);
and UO_722 (O_722,N_29983,N_29811);
nor UO_723 (O_723,N_29903,N_29909);
nor UO_724 (O_724,N_29804,N_29901);
and UO_725 (O_725,N_29940,N_29939);
nand UO_726 (O_726,N_29926,N_29813);
nand UO_727 (O_727,N_29874,N_29861);
nor UO_728 (O_728,N_29802,N_29988);
and UO_729 (O_729,N_29836,N_29970);
xor UO_730 (O_730,N_29975,N_29941);
nor UO_731 (O_731,N_29966,N_29989);
nand UO_732 (O_732,N_29861,N_29946);
xor UO_733 (O_733,N_29872,N_29804);
and UO_734 (O_734,N_29832,N_29972);
nand UO_735 (O_735,N_29801,N_29929);
or UO_736 (O_736,N_29823,N_29880);
nand UO_737 (O_737,N_29813,N_29996);
nand UO_738 (O_738,N_29920,N_29967);
nand UO_739 (O_739,N_29839,N_29953);
xor UO_740 (O_740,N_29952,N_29924);
xor UO_741 (O_741,N_29939,N_29861);
xnor UO_742 (O_742,N_29887,N_29991);
xnor UO_743 (O_743,N_29888,N_29886);
xor UO_744 (O_744,N_29813,N_29812);
nor UO_745 (O_745,N_29818,N_29930);
or UO_746 (O_746,N_29851,N_29986);
nor UO_747 (O_747,N_29814,N_29880);
or UO_748 (O_748,N_29801,N_29941);
nor UO_749 (O_749,N_29974,N_29818);
xor UO_750 (O_750,N_29911,N_29912);
nor UO_751 (O_751,N_29833,N_29907);
nor UO_752 (O_752,N_29892,N_29813);
and UO_753 (O_753,N_29950,N_29811);
xnor UO_754 (O_754,N_29874,N_29860);
or UO_755 (O_755,N_29933,N_29807);
nor UO_756 (O_756,N_29805,N_29874);
nor UO_757 (O_757,N_29820,N_29910);
or UO_758 (O_758,N_29997,N_29885);
and UO_759 (O_759,N_29871,N_29954);
nand UO_760 (O_760,N_29965,N_29901);
xnor UO_761 (O_761,N_29910,N_29837);
or UO_762 (O_762,N_29831,N_29890);
nand UO_763 (O_763,N_29818,N_29947);
or UO_764 (O_764,N_29935,N_29982);
xnor UO_765 (O_765,N_29827,N_29890);
or UO_766 (O_766,N_29885,N_29938);
and UO_767 (O_767,N_29888,N_29927);
nor UO_768 (O_768,N_29943,N_29976);
and UO_769 (O_769,N_29946,N_29972);
xor UO_770 (O_770,N_29957,N_29939);
xnor UO_771 (O_771,N_29853,N_29947);
xor UO_772 (O_772,N_29959,N_29892);
and UO_773 (O_773,N_29908,N_29903);
nand UO_774 (O_774,N_29819,N_29817);
nor UO_775 (O_775,N_29829,N_29934);
xnor UO_776 (O_776,N_29853,N_29933);
nor UO_777 (O_777,N_29891,N_29910);
xnor UO_778 (O_778,N_29976,N_29971);
and UO_779 (O_779,N_29866,N_29821);
xor UO_780 (O_780,N_29996,N_29852);
nor UO_781 (O_781,N_29851,N_29920);
xnor UO_782 (O_782,N_29830,N_29908);
or UO_783 (O_783,N_29871,N_29825);
or UO_784 (O_784,N_29950,N_29962);
or UO_785 (O_785,N_29925,N_29920);
or UO_786 (O_786,N_29830,N_29865);
xor UO_787 (O_787,N_29972,N_29867);
or UO_788 (O_788,N_29966,N_29973);
xnor UO_789 (O_789,N_29973,N_29991);
xnor UO_790 (O_790,N_29955,N_29814);
and UO_791 (O_791,N_29841,N_29858);
xnor UO_792 (O_792,N_29839,N_29990);
and UO_793 (O_793,N_29933,N_29846);
or UO_794 (O_794,N_29838,N_29883);
xnor UO_795 (O_795,N_29973,N_29957);
and UO_796 (O_796,N_29845,N_29859);
and UO_797 (O_797,N_29886,N_29876);
or UO_798 (O_798,N_29816,N_29901);
or UO_799 (O_799,N_29812,N_29988);
or UO_800 (O_800,N_29903,N_29968);
or UO_801 (O_801,N_29840,N_29949);
and UO_802 (O_802,N_29848,N_29829);
xnor UO_803 (O_803,N_29895,N_29814);
xnor UO_804 (O_804,N_29845,N_29941);
nand UO_805 (O_805,N_29967,N_29931);
or UO_806 (O_806,N_29831,N_29803);
and UO_807 (O_807,N_29968,N_29957);
nor UO_808 (O_808,N_29838,N_29847);
nor UO_809 (O_809,N_29878,N_29976);
nor UO_810 (O_810,N_29827,N_29904);
nor UO_811 (O_811,N_29899,N_29955);
xor UO_812 (O_812,N_29836,N_29832);
nand UO_813 (O_813,N_29821,N_29925);
nor UO_814 (O_814,N_29893,N_29825);
xnor UO_815 (O_815,N_29828,N_29967);
xnor UO_816 (O_816,N_29899,N_29834);
nand UO_817 (O_817,N_29844,N_29877);
and UO_818 (O_818,N_29849,N_29850);
xor UO_819 (O_819,N_29934,N_29862);
or UO_820 (O_820,N_29849,N_29879);
xnor UO_821 (O_821,N_29819,N_29833);
and UO_822 (O_822,N_29957,N_29800);
nand UO_823 (O_823,N_29877,N_29865);
nand UO_824 (O_824,N_29967,N_29946);
or UO_825 (O_825,N_29987,N_29997);
nor UO_826 (O_826,N_29973,N_29816);
xor UO_827 (O_827,N_29945,N_29822);
and UO_828 (O_828,N_29947,N_29919);
or UO_829 (O_829,N_29940,N_29808);
and UO_830 (O_830,N_29800,N_29932);
nand UO_831 (O_831,N_29818,N_29992);
nor UO_832 (O_832,N_29981,N_29888);
and UO_833 (O_833,N_29967,N_29917);
nor UO_834 (O_834,N_29897,N_29810);
nor UO_835 (O_835,N_29814,N_29851);
and UO_836 (O_836,N_29849,N_29946);
and UO_837 (O_837,N_29830,N_29838);
or UO_838 (O_838,N_29956,N_29829);
and UO_839 (O_839,N_29952,N_29931);
xnor UO_840 (O_840,N_29887,N_29912);
nor UO_841 (O_841,N_29818,N_29856);
nand UO_842 (O_842,N_29806,N_29855);
or UO_843 (O_843,N_29921,N_29983);
xnor UO_844 (O_844,N_29983,N_29916);
nand UO_845 (O_845,N_29900,N_29949);
xnor UO_846 (O_846,N_29828,N_29925);
or UO_847 (O_847,N_29833,N_29959);
nor UO_848 (O_848,N_29848,N_29918);
and UO_849 (O_849,N_29957,N_29846);
nand UO_850 (O_850,N_29816,N_29992);
nor UO_851 (O_851,N_29925,N_29894);
and UO_852 (O_852,N_29865,N_29871);
and UO_853 (O_853,N_29810,N_29945);
nor UO_854 (O_854,N_29997,N_29812);
nor UO_855 (O_855,N_29902,N_29821);
and UO_856 (O_856,N_29846,N_29804);
nor UO_857 (O_857,N_29961,N_29831);
nor UO_858 (O_858,N_29897,N_29975);
xor UO_859 (O_859,N_29991,N_29896);
and UO_860 (O_860,N_29895,N_29935);
xor UO_861 (O_861,N_29850,N_29838);
nand UO_862 (O_862,N_29871,N_29952);
nor UO_863 (O_863,N_29845,N_29862);
nor UO_864 (O_864,N_29828,N_29807);
or UO_865 (O_865,N_29973,N_29817);
nand UO_866 (O_866,N_29906,N_29878);
nor UO_867 (O_867,N_29827,N_29824);
nand UO_868 (O_868,N_29973,N_29850);
nand UO_869 (O_869,N_29800,N_29865);
nand UO_870 (O_870,N_29908,N_29855);
nand UO_871 (O_871,N_29990,N_29974);
and UO_872 (O_872,N_29994,N_29846);
xor UO_873 (O_873,N_29841,N_29882);
xnor UO_874 (O_874,N_29992,N_29880);
nand UO_875 (O_875,N_29994,N_29972);
xnor UO_876 (O_876,N_29806,N_29889);
or UO_877 (O_877,N_29901,N_29957);
nor UO_878 (O_878,N_29997,N_29844);
or UO_879 (O_879,N_29975,N_29843);
nor UO_880 (O_880,N_29849,N_29958);
xor UO_881 (O_881,N_29919,N_29977);
nand UO_882 (O_882,N_29904,N_29844);
and UO_883 (O_883,N_29813,N_29943);
and UO_884 (O_884,N_29823,N_29843);
or UO_885 (O_885,N_29938,N_29981);
xnor UO_886 (O_886,N_29897,N_29979);
xnor UO_887 (O_887,N_29827,N_29971);
and UO_888 (O_888,N_29979,N_29815);
and UO_889 (O_889,N_29891,N_29825);
xnor UO_890 (O_890,N_29956,N_29811);
xnor UO_891 (O_891,N_29938,N_29903);
nor UO_892 (O_892,N_29815,N_29809);
and UO_893 (O_893,N_29946,N_29942);
or UO_894 (O_894,N_29973,N_29825);
nor UO_895 (O_895,N_29843,N_29881);
nand UO_896 (O_896,N_29973,N_29933);
or UO_897 (O_897,N_29870,N_29878);
nor UO_898 (O_898,N_29992,N_29984);
nand UO_899 (O_899,N_29811,N_29969);
xor UO_900 (O_900,N_29892,N_29822);
nand UO_901 (O_901,N_29812,N_29804);
xnor UO_902 (O_902,N_29927,N_29992);
nand UO_903 (O_903,N_29827,N_29900);
nand UO_904 (O_904,N_29898,N_29956);
or UO_905 (O_905,N_29878,N_29819);
nor UO_906 (O_906,N_29818,N_29942);
or UO_907 (O_907,N_29916,N_29904);
nand UO_908 (O_908,N_29810,N_29955);
and UO_909 (O_909,N_29918,N_29842);
xnor UO_910 (O_910,N_29863,N_29950);
or UO_911 (O_911,N_29858,N_29899);
nand UO_912 (O_912,N_29894,N_29971);
nor UO_913 (O_913,N_29945,N_29983);
and UO_914 (O_914,N_29861,N_29957);
xor UO_915 (O_915,N_29872,N_29990);
and UO_916 (O_916,N_29818,N_29853);
nand UO_917 (O_917,N_29841,N_29959);
nor UO_918 (O_918,N_29855,N_29976);
nor UO_919 (O_919,N_29919,N_29932);
xnor UO_920 (O_920,N_29850,N_29952);
nand UO_921 (O_921,N_29851,N_29832);
or UO_922 (O_922,N_29881,N_29924);
xor UO_923 (O_923,N_29817,N_29989);
or UO_924 (O_924,N_29934,N_29833);
nand UO_925 (O_925,N_29897,N_29890);
or UO_926 (O_926,N_29930,N_29823);
nor UO_927 (O_927,N_29943,N_29809);
nand UO_928 (O_928,N_29856,N_29976);
nand UO_929 (O_929,N_29901,N_29810);
and UO_930 (O_930,N_29875,N_29975);
or UO_931 (O_931,N_29930,N_29828);
nand UO_932 (O_932,N_29900,N_29873);
xnor UO_933 (O_933,N_29828,N_29997);
or UO_934 (O_934,N_29913,N_29806);
or UO_935 (O_935,N_29826,N_29965);
xor UO_936 (O_936,N_29943,N_29939);
xnor UO_937 (O_937,N_29950,N_29873);
xnor UO_938 (O_938,N_29889,N_29929);
and UO_939 (O_939,N_29904,N_29920);
nor UO_940 (O_940,N_29935,N_29848);
xor UO_941 (O_941,N_29888,N_29805);
and UO_942 (O_942,N_29992,N_29872);
nor UO_943 (O_943,N_29875,N_29988);
xor UO_944 (O_944,N_29880,N_29893);
or UO_945 (O_945,N_29829,N_29915);
nor UO_946 (O_946,N_29922,N_29846);
nand UO_947 (O_947,N_29830,N_29882);
nor UO_948 (O_948,N_29916,N_29961);
or UO_949 (O_949,N_29905,N_29951);
and UO_950 (O_950,N_29824,N_29898);
xnor UO_951 (O_951,N_29956,N_29821);
and UO_952 (O_952,N_29909,N_29824);
nor UO_953 (O_953,N_29822,N_29861);
xor UO_954 (O_954,N_29883,N_29844);
and UO_955 (O_955,N_29819,N_29890);
and UO_956 (O_956,N_29997,N_29805);
nor UO_957 (O_957,N_29988,N_29898);
nor UO_958 (O_958,N_29876,N_29812);
or UO_959 (O_959,N_29957,N_29977);
or UO_960 (O_960,N_29914,N_29905);
or UO_961 (O_961,N_29953,N_29946);
xnor UO_962 (O_962,N_29988,N_29805);
or UO_963 (O_963,N_29928,N_29855);
nand UO_964 (O_964,N_29937,N_29998);
nor UO_965 (O_965,N_29966,N_29825);
xnor UO_966 (O_966,N_29965,N_29905);
and UO_967 (O_967,N_29871,N_29864);
nand UO_968 (O_968,N_29819,N_29864);
or UO_969 (O_969,N_29901,N_29841);
and UO_970 (O_970,N_29977,N_29865);
or UO_971 (O_971,N_29883,N_29885);
nand UO_972 (O_972,N_29805,N_29952);
nand UO_973 (O_973,N_29808,N_29894);
nand UO_974 (O_974,N_29875,N_29866);
nor UO_975 (O_975,N_29949,N_29826);
xnor UO_976 (O_976,N_29986,N_29825);
nand UO_977 (O_977,N_29984,N_29930);
and UO_978 (O_978,N_29915,N_29997);
and UO_979 (O_979,N_29818,N_29887);
nor UO_980 (O_980,N_29964,N_29903);
or UO_981 (O_981,N_29854,N_29875);
or UO_982 (O_982,N_29955,N_29987);
nor UO_983 (O_983,N_29906,N_29985);
xor UO_984 (O_984,N_29805,N_29910);
and UO_985 (O_985,N_29949,N_29975);
or UO_986 (O_986,N_29800,N_29853);
or UO_987 (O_987,N_29973,N_29871);
nand UO_988 (O_988,N_29872,N_29949);
nor UO_989 (O_989,N_29989,N_29885);
xor UO_990 (O_990,N_29838,N_29903);
nor UO_991 (O_991,N_29972,N_29925);
and UO_992 (O_992,N_29855,N_29895);
or UO_993 (O_993,N_29850,N_29985);
nand UO_994 (O_994,N_29824,N_29992);
xor UO_995 (O_995,N_29909,N_29949);
xor UO_996 (O_996,N_29936,N_29887);
nor UO_997 (O_997,N_29969,N_29830);
or UO_998 (O_998,N_29917,N_29874);
nand UO_999 (O_999,N_29858,N_29926);
nand UO_1000 (O_1000,N_29999,N_29868);
and UO_1001 (O_1001,N_29889,N_29850);
nand UO_1002 (O_1002,N_29803,N_29946);
nand UO_1003 (O_1003,N_29935,N_29808);
or UO_1004 (O_1004,N_29951,N_29896);
and UO_1005 (O_1005,N_29923,N_29854);
and UO_1006 (O_1006,N_29930,N_29959);
xor UO_1007 (O_1007,N_29838,N_29937);
nor UO_1008 (O_1008,N_29828,N_29869);
nor UO_1009 (O_1009,N_29969,N_29932);
nand UO_1010 (O_1010,N_29858,N_29869);
nand UO_1011 (O_1011,N_29943,N_29870);
nand UO_1012 (O_1012,N_29881,N_29842);
and UO_1013 (O_1013,N_29896,N_29928);
and UO_1014 (O_1014,N_29938,N_29906);
and UO_1015 (O_1015,N_29897,N_29924);
nand UO_1016 (O_1016,N_29988,N_29999);
and UO_1017 (O_1017,N_29999,N_29950);
xnor UO_1018 (O_1018,N_29900,N_29995);
xor UO_1019 (O_1019,N_29962,N_29939);
xnor UO_1020 (O_1020,N_29955,N_29822);
nand UO_1021 (O_1021,N_29960,N_29989);
or UO_1022 (O_1022,N_29992,N_29802);
and UO_1023 (O_1023,N_29862,N_29881);
and UO_1024 (O_1024,N_29880,N_29936);
or UO_1025 (O_1025,N_29928,N_29964);
or UO_1026 (O_1026,N_29898,N_29954);
nand UO_1027 (O_1027,N_29903,N_29853);
xor UO_1028 (O_1028,N_29979,N_29908);
nand UO_1029 (O_1029,N_29809,N_29882);
and UO_1030 (O_1030,N_29993,N_29914);
nor UO_1031 (O_1031,N_29939,N_29857);
nor UO_1032 (O_1032,N_29899,N_29869);
or UO_1033 (O_1033,N_29885,N_29879);
nor UO_1034 (O_1034,N_29960,N_29980);
nor UO_1035 (O_1035,N_29894,N_29896);
nor UO_1036 (O_1036,N_29997,N_29982);
nand UO_1037 (O_1037,N_29898,N_29986);
nand UO_1038 (O_1038,N_29836,N_29843);
nor UO_1039 (O_1039,N_29927,N_29834);
nor UO_1040 (O_1040,N_29928,N_29909);
or UO_1041 (O_1041,N_29912,N_29832);
xor UO_1042 (O_1042,N_29820,N_29879);
and UO_1043 (O_1043,N_29853,N_29849);
and UO_1044 (O_1044,N_29845,N_29957);
xnor UO_1045 (O_1045,N_29926,N_29817);
nand UO_1046 (O_1046,N_29945,N_29892);
or UO_1047 (O_1047,N_29930,N_29919);
and UO_1048 (O_1048,N_29843,N_29855);
or UO_1049 (O_1049,N_29865,N_29873);
and UO_1050 (O_1050,N_29987,N_29803);
nand UO_1051 (O_1051,N_29901,N_29873);
xnor UO_1052 (O_1052,N_29916,N_29984);
and UO_1053 (O_1053,N_29953,N_29978);
xnor UO_1054 (O_1054,N_29826,N_29928);
nand UO_1055 (O_1055,N_29963,N_29880);
nand UO_1056 (O_1056,N_29948,N_29831);
nor UO_1057 (O_1057,N_29876,N_29887);
and UO_1058 (O_1058,N_29870,N_29982);
nand UO_1059 (O_1059,N_29869,N_29808);
xnor UO_1060 (O_1060,N_29862,N_29843);
nand UO_1061 (O_1061,N_29850,N_29965);
xor UO_1062 (O_1062,N_29912,N_29932);
nand UO_1063 (O_1063,N_29950,N_29849);
and UO_1064 (O_1064,N_29860,N_29885);
nand UO_1065 (O_1065,N_29844,N_29888);
xnor UO_1066 (O_1066,N_29846,N_29920);
and UO_1067 (O_1067,N_29909,N_29977);
or UO_1068 (O_1068,N_29904,N_29899);
xor UO_1069 (O_1069,N_29815,N_29900);
nand UO_1070 (O_1070,N_29975,N_29845);
nor UO_1071 (O_1071,N_29960,N_29978);
or UO_1072 (O_1072,N_29946,N_29990);
xor UO_1073 (O_1073,N_29968,N_29994);
nor UO_1074 (O_1074,N_29908,N_29876);
nor UO_1075 (O_1075,N_29804,N_29931);
and UO_1076 (O_1076,N_29805,N_29870);
and UO_1077 (O_1077,N_29892,N_29935);
nor UO_1078 (O_1078,N_29987,N_29963);
or UO_1079 (O_1079,N_29845,N_29833);
and UO_1080 (O_1080,N_29852,N_29968);
or UO_1081 (O_1081,N_29843,N_29846);
nand UO_1082 (O_1082,N_29977,N_29872);
nand UO_1083 (O_1083,N_29928,N_29864);
or UO_1084 (O_1084,N_29973,N_29937);
and UO_1085 (O_1085,N_29868,N_29898);
nor UO_1086 (O_1086,N_29895,N_29874);
or UO_1087 (O_1087,N_29914,N_29920);
nor UO_1088 (O_1088,N_29921,N_29820);
or UO_1089 (O_1089,N_29924,N_29867);
xnor UO_1090 (O_1090,N_29864,N_29994);
nand UO_1091 (O_1091,N_29929,N_29816);
nor UO_1092 (O_1092,N_29871,N_29968);
or UO_1093 (O_1093,N_29883,N_29953);
nor UO_1094 (O_1094,N_29846,N_29830);
or UO_1095 (O_1095,N_29901,N_29968);
nand UO_1096 (O_1096,N_29984,N_29904);
and UO_1097 (O_1097,N_29938,N_29942);
and UO_1098 (O_1098,N_29870,N_29988);
or UO_1099 (O_1099,N_29944,N_29847);
nor UO_1100 (O_1100,N_29995,N_29844);
nand UO_1101 (O_1101,N_29852,N_29949);
or UO_1102 (O_1102,N_29955,N_29944);
nor UO_1103 (O_1103,N_29861,N_29889);
nor UO_1104 (O_1104,N_29905,N_29950);
nor UO_1105 (O_1105,N_29861,N_29981);
and UO_1106 (O_1106,N_29922,N_29815);
nand UO_1107 (O_1107,N_29843,N_29815);
nand UO_1108 (O_1108,N_29818,N_29815);
nor UO_1109 (O_1109,N_29805,N_29927);
xor UO_1110 (O_1110,N_29857,N_29852);
nor UO_1111 (O_1111,N_29890,N_29875);
or UO_1112 (O_1112,N_29873,N_29817);
nand UO_1113 (O_1113,N_29850,N_29879);
nor UO_1114 (O_1114,N_29973,N_29952);
xor UO_1115 (O_1115,N_29833,N_29821);
nand UO_1116 (O_1116,N_29861,N_29924);
xor UO_1117 (O_1117,N_29828,N_29993);
nand UO_1118 (O_1118,N_29925,N_29895);
nand UO_1119 (O_1119,N_29829,N_29982);
nand UO_1120 (O_1120,N_29952,N_29923);
xnor UO_1121 (O_1121,N_29955,N_29828);
xnor UO_1122 (O_1122,N_29992,N_29948);
or UO_1123 (O_1123,N_29830,N_29979);
nor UO_1124 (O_1124,N_29972,N_29938);
nor UO_1125 (O_1125,N_29809,N_29931);
and UO_1126 (O_1126,N_29896,N_29818);
nand UO_1127 (O_1127,N_29943,N_29839);
and UO_1128 (O_1128,N_29842,N_29984);
nand UO_1129 (O_1129,N_29854,N_29926);
nand UO_1130 (O_1130,N_29806,N_29803);
nor UO_1131 (O_1131,N_29992,N_29832);
and UO_1132 (O_1132,N_29913,N_29978);
xor UO_1133 (O_1133,N_29885,N_29929);
nand UO_1134 (O_1134,N_29825,N_29918);
xor UO_1135 (O_1135,N_29939,N_29915);
nand UO_1136 (O_1136,N_29972,N_29993);
xor UO_1137 (O_1137,N_29924,N_29801);
or UO_1138 (O_1138,N_29943,N_29949);
nand UO_1139 (O_1139,N_29820,N_29823);
and UO_1140 (O_1140,N_29834,N_29931);
xor UO_1141 (O_1141,N_29854,N_29991);
nand UO_1142 (O_1142,N_29811,N_29839);
and UO_1143 (O_1143,N_29846,N_29965);
xnor UO_1144 (O_1144,N_29836,N_29977);
and UO_1145 (O_1145,N_29839,N_29971);
nand UO_1146 (O_1146,N_29967,N_29860);
and UO_1147 (O_1147,N_29858,N_29992);
nand UO_1148 (O_1148,N_29922,N_29981);
or UO_1149 (O_1149,N_29905,N_29984);
and UO_1150 (O_1150,N_29827,N_29819);
or UO_1151 (O_1151,N_29841,N_29918);
nor UO_1152 (O_1152,N_29822,N_29804);
xor UO_1153 (O_1153,N_29930,N_29918);
nand UO_1154 (O_1154,N_29867,N_29976);
xor UO_1155 (O_1155,N_29973,N_29818);
xor UO_1156 (O_1156,N_29892,N_29837);
nand UO_1157 (O_1157,N_29872,N_29897);
xor UO_1158 (O_1158,N_29941,N_29947);
nand UO_1159 (O_1159,N_29954,N_29840);
xor UO_1160 (O_1160,N_29879,N_29965);
or UO_1161 (O_1161,N_29842,N_29800);
nand UO_1162 (O_1162,N_29969,N_29976);
nand UO_1163 (O_1163,N_29916,N_29853);
and UO_1164 (O_1164,N_29991,N_29905);
xnor UO_1165 (O_1165,N_29979,N_29918);
or UO_1166 (O_1166,N_29852,N_29868);
nand UO_1167 (O_1167,N_29978,N_29824);
xnor UO_1168 (O_1168,N_29830,N_29819);
xnor UO_1169 (O_1169,N_29887,N_29983);
xnor UO_1170 (O_1170,N_29853,N_29837);
nor UO_1171 (O_1171,N_29894,N_29936);
nor UO_1172 (O_1172,N_29979,N_29882);
xor UO_1173 (O_1173,N_29943,N_29963);
or UO_1174 (O_1174,N_29850,N_29898);
or UO_1175 (O_1175,N_29893,N_29900);
or UO_1176 (O_1176,N_29868,N_29953);
nand UO_1177 (O_1177,N_29831,N_29964);
nor UO_1178 (O_1178,N_29948,N_29811);
nand UO_1179 (O_1179,N_29959,N_29834);
nand UO_1180 (O_1180,N_29842,N_29840);
or UO_1181 (O_1181,N_29820,N_29942);
xor UO_1182 (O_1182,N_29997,N_29949);
nor UO_1183 (O_1183,N_29969,N_29935);
or UO_1184 (O_1184,N_29938,N_29880);
or UO_1185 (O_1185,N_29976,N_29939);
xnor UO_1186 (O_1186,N_29976,N_29822);
nor UO_1187 (O_1187,N_29818,N_29912);
xor UO_1188 (O_1188,N_29845,N_29988);
nor UO_1189 (O_1189,N_29909,N_29854);
nor UO_1190 (O_1190,N_29869,N_29888);
and UO_1191 (O_1191,N_29800,N_29816);
and UO_1192 (O_1192,N_29935,N_29907);
xnor UO_1193 (O_1193,N_29814,N_29827);
nand UO_1194 (O_1194,N_29965,N_29993);
nand UO_1195 (O_1195,N_29879,N_29999);
and UO_1196 (O_1196,N_29943,N_29819);
or UO_1197 (O_1197,N_29931,N_29982);
nor UO_1198 (O_1198,N_29864,N_29984);
or UO_1199 (O_1199,N_29807,N_29967);
xnor UO_1200 (O_1200,N_29986,N_29983);
or UO_1201 (O_1201,N_29934,N_29831);
xor UO_1202 (O_1202,N_29859,N_29833);
nor UO_1203 (O_1203,N_29946,N_29952);
or UO_1204 (O_1204,N_29958,N_29939);
xor UO_1205 (O_1205,N_29929,N_29959);
xor UO_1206 (O_1206,N_29950,N_29943);
or UO_1207 (O_1207,N_29897,N_29982);
and UO_1208 (O_1208,N_29924,N_29937);
and UO_1209 (O_1209,N_29865,N_29979);
xor UO_1210 (O_1210,N_29857,N_29847);
nand UO_1211 (O_1211,N_29987,N_29998);
and UO_1212 (O_1212,N_29978,N_29819);
nand UO_1213 (O_1213,N_29910,N_29955);
nor UO_1214 (O_1214,N_29857,N_29936);
and UO_1215 (O_1215,N_29933,N_29802);
nand UO_1216 (O_1216,N_29891,N_29953);
nand UO_1217 (O_1217,N_29891,N_29877);
and UO_1218 (O_1218,N_29953,N_29995);
xor UO_1219 (O_1219,N_29836,N_29905);
nor UO_1220 (O_1220,N_29917,N_29898);
nand UO_1221 (O_1221,N_29867,N_29913);
or UO_1222 (O_1222,N_29895,N_29861);
nand UO_1223 (O_1223,N_29972,N_29939);
xnor UO_1224 (O_1224,N_29839,N_29854);
nand UO_1225 (O_1225,N_29912,N_29925);
and UO_1226 (O_1226,N_29836,N_29916);
nand UO_1227 (O_1227,N_29850,N_29903);
nor UO_1228 (O_1228,N_29936,N_29843);
or UO_1229 (O_1229,N_29860,N_29870);
or UO_1230 (O_1230,N_29890,N_29951);
or UO_1231 (O_1231,N_29887,N_29870);
nor UO_1232 (O_1232,N_29993,N_29944);
xnor UO_1233 (O_1233,N_29878,N_29943);
and UO_1234 (O_1234,N_29860,N_29966);
nand UO_1235 (O_1235,N_29922,N_29914);
or UO_1236 (O_1236,N_29976,N_29884);
or UO_1237 (O_1237,N_29902,N_29976);
xnor UO_1238 (O_1238,N_29823,N_29979);
nor UO_1239 (O_1239,N_29898,N_29873);
or UO_1240 (O_1240,N_29916,N_29900);
or UO_1241 (O_1241,N_29864,N_29883);
nor UO_1242 (O_1242,N_29873,N_29929);
nor UO_1243 (O_1243,N_29972,N_29969);
xor UO_1244 (O_1244,N_29893,N_29889);
nand UO_1245 (O_1245,N_29832,N_29901);
xnor UO_1246 (O_1246,N_29942,N_29994);
nor UO_1247 (O_1247,N_29860,N_29897);
or UO_1248 (O_1248,N_29918,N_29856);
and UO_1249 (O_1249,N_29958,N_29874);
nand UO_1250 (O_1250,N_29880,N_29877);
nor UO_1251 (O_1251,N_29821,N_29827);
and UO_1252 (O_1252,N_29809,N_29973);
xnor UO_1253 (O_1253,N_29818,N_29983);
and UO_1254 (O_1254,N_29896,N_29966);
xor UO_1255 (O_1255,N_29880,N_29939);
xnor UO_1256 (O_1256,N_29919,N_29913);
or UO_1257 (O_1257,N_29929,N_29948);
nor UO_1258 (O_1258,N_29953,N_29821);
and UO_1259 (O_1259,N_29995,N_29926);
or UO_1260 (O_1260,N_29871,N_29913);
xnor UO_1261 (O_1261,N_29889,N_29957);
nand UO_1262 (O_1262,N_29832,N_29971);
nor UO_1263 (O_1263,N_29863,N_29925);
nand UO_1264 (O_1264,N_29830,N_29950);
and UO_1265 (O_1265,N_29871,N_29839);
and UO_1266 (O_1266,N_29824,N_29934);
and UO_1267 (O_1267,N_29871,N_29894);
nor UO_1268 (O_1268,N_29813,N_29958);
nor UO_1269 (O_1269,N_29953,N_29802);
nand UO_1270 (O_1270,N_29813,N_29816);
nand UO_1271 (O_1271,N_29829,N_29914);
or UO_1272 (O_1272,N_29831,N_29855);
and UO_1273 (O_1273,N_29837,N_29878);
nand UO_1274 (O_1274,N_29987,N_29988);
and UO_1275 (O_1275,N_29878,N_29917);
and UO_1276 (O_1276,N_29821,N_29872);
xnor UO_1277 (O_1277,N_29919,N_29838);
nor UO_1278 (O_1278,N_29880,N_29885);
xnor UO_1279 (O_1279,N_29876,N_29802);
nor UO_1280 (O_1280,N_29803,N_29992);
or UO_1281 (O_1281,N_29886,N_29907);
nor UO_1282 (O_1282,N_29892,N_29975);
nor UO_1283 (O_1283,N_29818,N_29846);
and UO_1284 (O_1284,N_29889,N_29844);
nor UO_1285 (O_1285,N_29910,N_29831);
nand UO_1286 (O_1286,N_29846,N_29954);
nand UO_1287 (O_1287,N_29908,N_29892);
or UO_1288 (O_1288,N_29841,N_29853);
or UO_1289 (O_1289,N_29869,N_29872);
and UO_1290 (O_1290,N_29957,N_29820);
nor UO_1291 (O_1291,N_29935,N_29938);
nand UO_1292 (O_1292,N_29966,N_29975);
and UO_1293 (O_1293,N_29950,N_29856);
and UO_1294 (O_1294,N_29841,N_29839);
or UO_1295 (O_1295,N_29998,N_29813);
and UO_1296 (O_1296,N_29851,N_29967);
xnor UO_1297 (O_1297,N_29879,N_29918);
xnor UO_1298 (O_1298,N_29888,N_29903);
or UO_1299 (O_1299,N_29934,N_29860);
or UO_1300 (O_1300,N_29958,N_29881);
nand UO_1301 (O_1301,N_29838,N_29873);
xor UO_1302 (O_1302,N_29880,N_29969);
or UO_1303 (O_1303,N_29903,N_29868);
nor UO_1304 (O_1304,N_29924,N_29985);
or UO_1305 (O_1305,N_29990,N_29970);
nand UO_1306 (O_1306,N_29950,N_29945);
or UO_1307 (O_1307,N_29873,N_29839);
xnor UO_1308 (O_1308,N_29921,N_29852);
xnor UO_1309 (O_1309,N_29982,N_29968);
and UO_1310 (O_1310,N_29810,N_29857);
or UO_1311 (O_1311,N_29934,N_29802);
and UO_1312 (O_1312,N_29884,N_29918);
and UO_1313 (O_1313,N_29858,N_29931);
xor UO_1314 (O_1314,N_29858,N_29960);
and UO_1315 (O_1315,N_29814,N_29894);
xor UO_1316 (O_1316,N_29801,N_29839);
xor UO_1317 (O_1317,N_29923,N_29869);
nor UO_1318 (O_1318,N_29890,N_29964);
nand UO_1319 (O_1319,N_29949,N_29908);
nand UO_1320 (O_1320,N_29957,N_29887);
nand UO_1321 (O_1321,N_29805,N_29923);
and UO_1322 (O_1322,N_29803,N_29934);
or UO_1323 (O_1323,N_29832,N_29809);
and UO_1324 (O_1324,N_29927,N_29851);
xnor UO_1325 (O_1325,N_29961,N_29864);
and UO_1326 (O_1326,N_29991,N_29908);
xnor UO_1327 (O_1327,N_29889,N_29952);
xnor UO_1328 (O_1328,N_29906,N_29892);
or UO_1329 (O_1329,N_29948,N_29923);
and UO_1330 (O_1330,N_29837,N_29903);
nor UO_1331 (O_1331,N_29902,N_29837);
or UO_1332 (O_1332,N_29975,N_29911);
or UO_1333 (O_1333,N_29935,N_29899);
nand UO_1334 (O_1334,N_29810,N_29952);
nand UO_1335 (O_1335,N_29837,N_29949);
xnor UO_1336 (O_1336,N_29893,N_29879);
and UO_1337 (O_1337,N_29924,N_29850);
or UO_1338 (O_1338,N_29900,N_29976);
and UO_1339 (O_1339,N_29885,N_29924);
and UO_1340 (O_1340,N_29963,N_29838);
nor UO_1341 (O_1341,N_29839,N_29947);
or UO_1342 (O_1342,N_29895,N_29893);
xor UO_1343 (O_1343,N_29815,N_29807);
nor UO_1344 (O_1344,N_29870,N_29806);
or UO_1345 (O_1345,N_29931,N_29832);
and UO_1346 (O_1346,N_29866,N_29825);
or UO_1347 (O_1347,N_29943,N_29938);
xor UO_1348 (O_1348,N_29894,N_29873);
nor UO_1349 (O_1349,N_29963,N_29805);
nand UO_1350 (O_1350,N_29821,N_29903);
or UO_1351 (O_1351,N_29805,N_29931);
nor UO_1352 (O_1352,N_29878,N_29888);
or UO_1353 (O_1353,N_29878,N_29987);
or UO_1354 (O_1354,N_29861,N_29919);
xor UO_1355 (O_1355,N_29936,N_29874);
xnor UO_1356 (O_1356,N_29946,N_29907);
nand UO_1357 (O_1357,N_29900,N_29938);
nor UO_1358 (O_1358,N_29999,N_29864);
and UO_1359 (O_1359,N_29865,N_29863);
nor UO_1360 (O_1360,N_29819,N_29857);
or UO_1361 (O_1361,N_29940,N_29965);
or UO_1362 (O_1362,N_29885,N_29800);
nor UO_1363 (O_1363,N_29994,N_29888);
and UO_1364 (O_1364,N_29918,N_29889);
or UO_1365 (O_1365,N_29976,N_29996);
and UO_1366 (O_1366,N_29999,N_29832);
xor UO_1367 (O_1367,N_29808,N_29874);
nand UO_1368 (O_1368,N_29937,N_29851);
nand UO_1369 (O_1369,N_29812,N_29834);
or UO_1370 (O_1370,N_29956,N_29971);
nor UO_1371 (O_1371,N_29913,N_29819);
and UO_1372 (O_1372,N_29838,N_29948);
nand UO_1373 (O_1373,N_29903,N_29883);
nor UO_1374 (O_1374,N_29831,N_29801);
nor UO_1375 (O_1375,N_29955,N_29879);
or UO_1376 (O_1376,N_29826,N_29807);
or UO_1377 (O_1377,N_29972,N_29836);
xnor UO_1378 (O_1378,N_29957,N_29829);
and UO_1379 (O_1379,N_29818,N_29889);
xnor UO_1380 (O_1380,N_29946,N_29913);
or UO_1381 (O_1381,N_29933,N_29839);
or UO_1382 (O_1382,N_29896,N_29909);
and UO_1383 (O_1383,N_29855,N_29901);
nand UO_1384 (O_1384,N_29905,N_29990);
or UO_1385 (O_1385,N_29993,N_29977);
xnor UO_1386 (O_1386,N_29907,N_29827);
and UO_1387 (O_1387,N_29970,N_29973);
and UO_1388 (O_1388,N_29904,N_29889);
and UO_1389 (O_1389,N_29875,N_29808);
nor UO_1390 (O_1390,N_29999,N_29968);
or UO_1391 (O_1391,N_29987,N_29822);
and UO_1392 (O_1392,N_29906,N_29805);
nand UO_1393 (O_1393,N_29884,N_29824);
nor UO_1394 (O_1394,N_29963,N_29967);
nand UO_1395 (O_1395,N_29983,N_29984);
and UO_1396 (O_1396,N_29950,N_29882);
nand UO_1397 (O_1397,N_29869,N_29998);
or UO_1398 (O_1398,N_29823,N_29940);
nand UO_1399 (O_1399,N_29849,N_29800);
or UO_1400 (O_1400,N_29968,N_29909);
nor UO_1401 (O_1401,N_29803,N_29965);
and UO_1402 (O_1402,N_29847,N_29851);
xor UO_1403 (O_1403,N_29941,N_29873);
nand UO_1404 (O_1404,N_29843,N_29827);
and UO_1405 (O_1405,N_29919,N_29851);
xor UO_1406 (O_1406,N_29838,N_29951);
and UO_1407 (O_1407,N_29849,N_29855);
nor UO_1408 (O_1408,N_29883,N_29805);
nor UO_1409 (O_1409,N_29846,N_29831);
or UO_1410 (O_1410,N_29810,N_29907);
xnor UO_1411 (O_1411,N_29944,N_29800);
xor UO_1412 (O_1412,N_29961,N_29879);
nor UO_1413 (O_1413,N_29901,N_29976);
xor UO_1414 (O_1414,N_29823,N_29985);
nand UO_1415 (O_1415,N_29846,N_29947);
nor UO_1416 (O_1416,N_29892,N_29885);
xor UO_1417 (O_1417,N_29906,N_29948);
and UO_1418 (O_1418,N_29931,N_29932);
nand UO_1419 (O_1419,N_29868,N_29801);
nor UO_1420 (O_1420,N_29821,N_29999);
or UO_1421 (O_1421,N_29962,N_29945);
or UO_1422 (O_1422,N_29911,N_29843);
xnor UO_1423 (O_1423,N_29935,N_29995);
xnor UO_1424 (O_1424,N_29899,N_29978);
nand UO_1425 (O_1425,N_29814,N_29970);
and UO_1426 (O_1426,N_29940,N_29887);
and UO_1427 (O_1427,N_29868,N_29809);
nand UO_1428 (O_1428,N_29996,N_29824);
or UO_1429 (O_1429,N_29947,N_29892);
xnor UO_1430 (O_1430,N_29884,N_29872);
and UO_1431 (O_1431,N_29821,N_29815);
and UO_1432 (O_1432,N_29816,N_29987);
xnor UO_1433 (O_1433,N_29918,N_29838);
xnor UO_1434 (O_1434,N_29859,N_29923);
or UO_1435 (O_1435,N_29905,N_29925);
or UO_1436 (O_1436,N_29885,N_29995);
or UO_1437 (O_1437,N_29998,N_29816);
xnor UO_1438 (O_1438,N_29948,N_29995);
nor UO_1439 (O_1439,N_29996,N_29998);
or UO_1440 (O_1440,N_29823,N_29978);
and UO_1441 (O_1441,N_29913,N_29958);
nor UO_1442 (O_1442,N_29985,N_29965);
and UO_1443 (O_1443,N_29851,N_29939);
or UO_1444 (O_1444,N_29818,N_29835);
and UO_1445 (O_1445,N_29945,N_29933);
or UO_1446 (O_1446,N_29980,N_29912);
nand UO_1447 (O_1447,N_29942,N_29981);
or UO_1448 (O_1448,N_29957,N_29982);
xnor UO_1449 (O_1449,N_29927,N_29986);
xnor UO_1450 (O_1450,N_29867,N_29929);
nor UO_1451 (O_1451,N_29996,N_29940);
xnor UO_1452 (O_1452,N_29816,N_29847);
and UO_1453 (O_1453,N_29914,N_29917);
nor UO_1454 (O_1454,N_29850,N_29886);
xor UO_1455 (O_1455,N_29929,N_29804);
or UO_1456 (O_1456,N_29945,N_29800);
nand UO_1457 (O_1457,N_29809,N_29976);
nand UO_1458 (O_1458,N_29942,N_29901);
or UO_1459 (O_1459,N_29818,N_29834);
or UO_1460 (O_1460,N_29912,N_29964);
nor UO_1461 (O_1461,N_29864,N_29846);
nand UO_1462 (O_1462,N_29961,N_29902);
nor UO_1463 (O_1463,N_29869,N_29946);
nor UO_1464 (O_1464,N_29911,N_29982);
nor UO_1465 (O_1465,N_29880,N_29829);
or UO_1466 (O_1466,N_29984,N_29990);
or UO_1467 (O_1467,N_29861,N_29983);
or UO_1468 (O_1468,N_29957,N_29841);
nor UO_1469 (O_1469,N_29974,N_29868);
and UO_1470 (O_1470,N_29946,N_29816);
nand UO_1471 (O_1471,N_29853,N_29938);
and UO_1472 (O_1472,N_29867,N_29958);
nand UO_1473 (O_1473,N_29883,N_29977);
nor UO_1474 (O_1474,N_29988,N_29867);
nand UO_1475 (O_1475,N_29894,N_29913);
nor UO_1476 (O_1476,N_29806,N_29917);
and UO_1477 (O_1477,N_29897,N_29931);
or UO_1478 (O_1478,N_29992,N_29951);
and UO_1479 (O_1479,N_29920,N_29930);
or UO_1480 (O_1480,N_29929,N_29926);
nor UO_1481 (O_1481,N_29811,N_29915);
nor UO_1482 (O_1482,N_29822,N_29838);
nand UO_1483 (O_1483,N_29947,N_29845);
nand UO_1484 (O_1484,N_29812,N_29845);
nand UO_1485 (O_1485,N_29863,N_29920);
or UO_1486 (O_1486,N_29987,N_29836);
nand UO_1487 (O_1487,N_29814,N_29967);
nand UO_1488 (O_1488,N_29911,N_29929);
and UO_1489 (O_1489,N_29879,N_29906);
nor UO_1490 (O_1490,N_29943,N_29970);
or UO_1491 (O_1491,N_29955,N_29837);
nand UO_1492 (O_1492,N_29804,N_29956);
xnor UO_1493 (O_1493,N_29829,N_29943);
or UO_1494 (O_1494,N_29838,N_29871);
and UO_1495 (O_1495,N_29993,N_29874);
nand UO_1496 (O_1496,N_29882,N_29971);
nor UO_1497 (O_1497,N_29909,N_29954);
nand UO_1498 (O_1498,N_29804,N_29970);
xor UO_1499 (O_1499,N_29927,N_29833);
or UO_1500 (O_1500,N_29931,N_29864);
nor UO_1501 (O_1501,N_29971,N_29895);
and UO_1502 (O_1502,N_29867,N_29970);
xnor UO_1503 (O_1503,N_29868,N_29969);
and UO_1504 (O_1504,N_29890,N_29882);
nand UO_1505 (O_1505,N_29979,N_29868);
or UO_1506 (O_1506,N_29844,N_29971);
nand UO_1507 (O_1507,N_29911,N_29910);
and UO_1508 (O_1508,N_29847,N_29894);
nor UO_1509 (O_1509,N_29903,N_29852);
and UO_1510 (O_1510,N_29884,N_29840);
xor UO_1511 (O_1511,N_29993,N_29833);
nor UO_1512 (O_1512,N_29833,N_29812);
or UO_1513 (O_1513,N_29861,N_29859);
nor UO_1514 (O_1514,N_29905,N_29910);
xor UO_1515 (O_1515,N_29802,N_29801);
or UO_1516 (O_1516,N_29999,N_29810);
or UO_1517 (O_1517,N_29833,N_29903);
and UO_1518 (O_1518,N_29906,N_29946);
and UO_1519 (O_1519,N_29937,N_29913);
nor UO_1520 (O_1520,N_29859,N_29880);
xnor UO_1521 (O_1521,N_29924,N_29992);
nand UO_1522 (O_1522,N_29938,N_29975);
and UO_1523 (O_1523,N_29888,N_29959);
nor UO_1524 (O_1524,N_29998,N_29824);
and UO_1525 (O_1525,N_29870,N_29850);
and UO_1526 (O_1526,N_29995,N_29964);
xnor UO_1527 (O_1527,N_29894,N_29819);
or UO_1528 (O_1528,N_29869,N_29926);
or UO_1529 (O_1529,N_29937,N_29878);
nor UO_1530 (O_1530,N_29957,N_29923);
xor UO_1531 (O_1531,N_29956,N_29845);
and UO_1532 (O_1532,N_29917,N_29957);
xnor UO_1533 (O_1533,N_29850,N_29958);
nand UO_1534 (O_1534,N_29915,N_29927);
nand UO_1535 (O_1535,N_29994,N_29806);
nor UO_1536 (O_1536,N_29866,N_29990);
and UO_1537 (O_1537,N_29995,N_29913);
nor UO_1538 (O_1538,N_29903,N_29925);
or UO_1539 (O_1539,N_29838,N_29959);
nor UO_1540 (O_1540,N_29827,N_29973);
nor UO_1541 (O_1541,N_29810,N_29882);
nand UO_1542 (O_1542,N_29860,N_29861);
xor UO_1543 (O_1543,N_29808,N_29995);
or UO_1544 (O_1544,N_29910,N_29841);
xnor UO_1545 (O_1545,N_29917,N_29812);
nor UO_1546 (O_1546,N_29844,N_29902);
and UO_1547 (O_1547,N_29811,N_29982);
nand UO_1548 (O_1548,N_29857,N_29884);
xor UO_1549 (O_1549,N_29953,N_29842);
and UO_1550 (O_1550,N_29863,N_29843);
and UO_1551 (O_1551,N_29978,N_29984);
nand UO_1552 (O_1552,N_29903,N_29912);
or UO_1553 (O_1553,N_29996,N_29958);
or UO_1554 (O_1554,N_29981,N_29802);
and UO_1555 (O_1555,N_29836,N_29935);
nand UO_1556 (O_1556,N_29876,N_29893);
nand UO_1557 (O_1557,N_29967,N_29864);
or UO_1558 (O_1558,N_29859,N_29976);
nor UO_1559 (O_1559,N_29951,N_29999);
nand UO_1560 (O_1560,N_29912,N_29858);
or UO_1561 (O_1561,N_29974,N_29960);
and UO_1562 (O_1562,N_29968,N_29951);
nand UO_1563 (O_1563,N_29993,N_29842);
and UO_1564 (O_1564,N_29844,N_29947);
nand UO_1565 (O_1565,N_29836,N_29994);
nand UO_1566 (O_1566,N_29890,N_29966);
and UO_1567 (O_1567,N_29978,N_29894);
or UO_1568 (O_1568,N_29994,N_29869);
nor UO_1569 (O_1569,N_29852,N_29878);
nor UO_1570 (O_1570,N_29978,N_29808);
nand UO_1571 (O_1571,N_29858,N_29850);
xnor UO_1572 (O_1572,N_29865,N_29801);
nor UO_1573 (O_1573,N_29946,N_29993);
nor UO_1574 (O_1574,N_29808,N_29845);
nand UO_1575 (O_1575,N_29919,N_29892);
nand UO_1576 (O_1576,N_29980,N_29961);
or UO_1577 (O_1577,N_29811,N_29984);
or UO_1578 (O_1578,N_29976,N_29962);
and UO_1579 (O_1579,N_29808,N_29826);
nor UO_1580 (O_1580,N_29983,N_29839);
nand UO_1581 (O_1581,N_29804,N_29918);
and UO_1582 (O_1582,N_29908,N_29960);
or UO_1583 (O_1583,N_29977,N_29823);
or UO_1584 (O_1584,N_29862,N_29817);
or UO_1585 (O_1585,N_29846,N_29860);
nand UO_1586 (O_1586,N_29844,N_29899);
nor UO_1587 (O_1587,N_29833,N_29880);
or UO_1588 (O_1588,N_29859,N_29979);
nand UO_1589 (O_1589,N_29913,N_29989);
xnor UO_1590 (O_1590,N_29879,N_29998);
and UO_1591 (O_1591,N_29905,N_29904);
xor UO_1592 (O_1592,N_29934,N_29945);
and UO_1593 (O_1593,N_29907,N_29890);
nand UO_1594 (O_1594,N_29843,N_29931);
nand UO_1595 (O_1595,N_29941,N_29822);
nand UO_1596 (O_1596,N_29800,N_29920);
nand UO_1597 (O_1597,N_29931,N_29866);
and UO_1598 (O_1598,N_29904,N_29939);
and UO_1599 (O_1599,N_29935,N_29916);
nor UO_1600 (O_1600,N_29937,N_29986);
and UO_1601 (O_1601,N_29995,N_29868);
nor UO_1602 (O_1602,N_29952,N_29942);
nor UO_1603 (O_1603,N_29862,N_29812);
nand UO_1604 (O_1604,N_29968,N_29926);
nand UO_1605 (O_1605,N_29887,N_29871);
nand UO_1606 (O_1606,N_29901,N_29920);
nor UO_1607 (O_1607,N_29822,N_29840);
and UO_1608 (O_1608,N_29812,N_29924);
nand UO_1609 (O_1609,N_29827,N_29956);
nor UO_1610 (O_1610,N_29833,N_29831);
nor UO_1611 (O_1611,N_29999,N_29971);
or UO_1612 (O_1612,N_29954,N_29944);
or UO_1613 (O_1613,N_29813,N_29957);
nor UO_1614 (O_1614,N_29897,N_29854);
or UO_1615 (O_1615,N_29971,N_29970);
nor UO_1616 (O_1616,N_29894,N_29889);
nand UO_1617 (O_1617,N_29991,N_29999);
xor UO_1618 (O_1618,N_29812,N_29926);
nor UO_1619 (O_1619,N_29801,N_29864);
nor UO_1620 (O_1620,N_29910,N_29977);
or UO_1621 (O_1621,N_29953,N_29851);
xor UO_1622 (O_1622,N_29863,N_29971);
and UO_1623 (O_1623,N_29836,N_29803);
xor UO_1624 (O_1624,N_29855,N_29960);
nor UO_1625 (O_1625,N_29801,N_29809);
xnor UO_1626 (O_1626,N_29858,N_29979);
nand UO_1627 (O_1627,N_29904,N_29825);
or UO_1628 (O_1628,N_29936,N_29970);
and UO_1629 (O_1629,N_29822,N_29985);
nor UO_1630 (O_1630,N_29984,N_29936);
and UO_1631 (O_1631,N_29881,N_29850);
xnor UO_1632 (O_1632,N_29819,N_29834);
nand UO_1633 (O_1633,N_29916,N_29971);
nand UO_1634 (O_1634,N_29896,N_29918);
xnor UO_1635 (O_1635,N_29933,N_29913);
or UO_1636 (O_1636,N_29954,N_29800);
nor UO_1637 (O_1637,N_29895,N_29818);
or UO_1638 (O_1638,N_29963,N_29928);
xnor UO_1639 (O_1639,N_29894,N_29976);
and UO_1640 (O_1640,N_29844,N_29890);
or UO_1641 (O_1641,N_29898,N_29897);
nor UO_1642 (O_1642,N_29865,N_29839);
xnor UO_1643 (O_1643,N_29801,N_29903);
xnor UO_1644 (O_1644,N_29986,N_29854);
xor UO_1645 (O_1645,N_29805,N_29921);
and UO_1646 (O_1646,N_29880,N_29891);
and UO_1647 (O_1647,N_29823,N_29976);
or UO_1648 (O_1648,N_29974,N_29998);
nor UO_1649 (O_1649,N_29986,N_29910);
and UO_1650 (O_1650,N_29972,N_29841);
nor UO_1651 (O_1651,N_29988,N_29968);
or UO_1652 (O_1652,N_29887,N_29963);
xnor UO_1653 (O_1653,N_29913,N_29872);
nor UO_1654 (O_1654,N_29829,N_29894);
and UO_1655 (O_1655,N_29935,N_29981);
xor UO_1656 (O_1656,N_29882,N_29995);
nor UO_1657 (O_1657,N_29932,N_29840);
or UO_1658 (O_1658,N_29884,N_29907);
nand UO_1659 (O_1659,N_29897,N_29950);
nand UO_1660 (O_1660,N_29916,N_29958);
nor UO_1661 (O_1661,N_29870,N_29869);
or UO_1662 (O_1662,N_29993,N_29974);
xor UO_1663 (O_1663,N_29986,N_29808);
or UO_1664 (O_1664,N_29916,N_29869);
or UO_1665 (O_1665,N_29983,N_29959);
xor UO_1666 (O_1666,N_29963,N_29858);
and UO_1667 (O_1667,N_29814,N_29856);
nor UO_1668 (O_1668,N_29827,N_29948);
xnor UO_1669 (O_1669,N_29824,N_29970);
nor UO_1670 (O_1670,N_29816,N_29907);
nand UO_1671 (O_1671,N_29897,N_29940);
nand UO_1672 (O_1672,N_29899,N_29968);
or UO_1673 (O_1673,N_29994,N_29899);
and UO_1674 (O_1674,N_29847,N_29993);
and UO_1675 (O_1675,N_29883,N_29911);
and UO_1676 (O_1676,N_29913,N_29922);
nor UO_1677 (O_1677,N_29989,N_29873);
or UO_1678 (O_1678,N_29933,N_29868);
nand UO_1679 (O_1679,N_29888,N_29966);
nand UO_1680 (O_1680,N_29875,N_29837);
or UO_1681 (O_1681,N_29934,N_29935);
nand UO_1682 (O_1682,N_29980,N_29979);
xor UO_1683 (O_1683,N_29801,N_29855);
and UO_1684 (O_1684,N_29877,N_29927);
nor UO_1685 (O_1685,N_29872,N_29979);
xnor UO_1686 (O_1686,N_29806,N_29974);
xnor UO_1687 (O_1687,N_29924,N_29884);
nor UO_1688 (O_1688,N_29972,N_29999);
nand UO_1689 (O_1689,N_29908,N_29905);
nor UO_1690 (O_1690,N_29958,N_29897);
nand UO_1691 (O_1691,N_29964,N_29867);
or UO_1692 (O_1692,N_29805,N_29842);
and UO_1693 (O_1693,N_29954,N_29803);
xnor UO_1694 (O_1694,N_29965,N_29960);
nor UO_1695 (O_1695,N_29804,N_29875);
and UO_1696 (O_1696,N_29912,N_29828);
and UO_1697 (O_1697,N_29950,N_29942);
xnor UO_1698 (O_1698,N_29836,N_29860);
xnor UO_1699 (O_1699,N_29954,N_29940);
nand UO_1700 (O_1700,N_29857,N_29926);
nor UO_1701 (O_1701,N_29937,N_29880);
and UO_1702 (O_1702,N_29879,N_29947);
or UO_1703 (O_1703,N_29853,N_29859);
xor UO_1704 (O_1704,N_29802,N_29828);
or UO_1705 (O_1705,N_29968,N_29935);
nand UO_1706 (O_1706,N_29910,N_29872);
nand UO_1707 (O_1707,N_29835,N_29954);
nor UO_1708 (O_1708,N_29944,N_29874);
xor UO_1709 (O_1709,N_29892,N_29922);
and UO_1710 (O_1710,N_29868,N_29884);
nor UO_1711 (O_1711,N_29831,N_29937);
or UO_1712 (O_1712,N_29960,N_29849);
or UO_1713 (O_1713,N_29839,N_29877);
and UO_1714 (O_1714,N_29891,N_29823);
nor UO_1715 (O_1715,N_29842,N_29938);
or UO_1716 (O_1716,N_29889,N_29933);
and UO_1717 (O_1717,N_29839,N_29916);
nor UO_1718 (O_1718,N_29981,N_29842);
or UO_1719 (O_1719,N_29809,N_29851);
nand UO_1720 (O_1720,N_29941,N_29807);
and UO_1721 (O_1721,N_29826,N_29868);
or UO_1722 (O_1722,N_29814,N_29876);
nor UO_1723 (O_1723,N_29972,N_29879);
and UO_1724 (O_1724,N_29895,N_29898);
xnor UO_1725 (O_1725,N_29846,N_29893);
xor UO_1726 (O_1726,N_29832,N_29888);
nand UO_1727 (O_1727,N_29843,N_29941);
nand UO_1728 (O_1728,N_29940,N_29828);
and UO_1729 (O_1729,N_29918,N_29992);
nor UO_1730 (O_1730,N_29804,N_29937);
and UO_1731 (O_1731,N_29842,N_29835);
nor UO_1732 (O_1732,N_29803,N_29813);
nor UO_1733 (O_1733,N_29843,N_29804);
or UO_1734 (O_1734,N_29908,N_29887);
nand UO_1735 (O_1735,N_29988,N_29803);
or UO_1736 (O_1736,N_29922,N_29837);
and UO_1737 (O_1737,N_29998,N_29854);
nand UO_1738 (O_1738,N_29971,N_29967);
nand UO_1739 (O_1739,N_29881,N_29930);
xnor UO_1740 (O_1740,N_29838,N_29885);
nand UO_1741 (O_1741,N_29905,N_29923);
or UO_1742 (O_1742,N_29802,N_29860);
and UO_1743 (O_1743,N_29903,N_29818);
or UO_1744 (O_1744,N_29909,N_29852);
or UO_1745 (O_1745,N_29885,N_29927);
nor UO_1746 (O_1746,N_29934,N_29926);
nor UO_1747 (O_1747,N_29911,N_29966);
nand UO_1748 (O_1748,N_29976,N_29801);
xnor UO_1749 (O_1749,N_29937,N_29837);
nand UO_1750 (O_1750,N_29983,N_29923);
or UO_1751 (O_1751,N_29806,N_29818);
xor UO_1752 (O_1752,N_29909,N_29860);
nor UO_1753 (O_1753,N_29875,N_29874);
nand UO_1754 (O_1754,N_29810,N_29865);
and UO_1755 (O_1755,N_29924,N_29933);
and UO_1756 (O_1756,N_29964,N_29927);
and UO_1757 (O_1757,N_29917,N_29900);
and UO_1758 (O_1758,N_29820,N_29951);
xor UO_1759 (O_1759,N_29908,N_29963);
xnor UO_1760 (O_1760,N_29824,N_29844);
xor UO_1761 (O_1761,N_29930,N_29934);
nor UO_1762 (O_1762,N_29805,N_29903);
nand UO_1763 (O_1763,N_29924,N_29930);
nand UO_1764 (O_1764,N_29913,N_29844);
and UO_1765 (O_1765,N_29828,N_29909);
or UO_1766 (O_1766,N_29824,N_29886);
nor UO_1767 (O_1767,N_29942,N_29882);
and UO_1768 (O_1768,N_29819,N_29859);
or UO_1769 (O_1769,N_29917,N_29890);
and UO_1770 (O_1770,N_29828,N_29960);
or UO_1771 (O_1771,N_29988,N_29899);
and UO_1772 (O_1772,N_29841,N_29989);
nor UO_1773 (O_1773,N_29995,N_29894);
nand UO_1774 (O_1774,N_29908,N_29864);
nor UO_1775 (O_1775,N_29926,N_29930);
nand UO_1776 (O_1776,N_29949,N_29979);
nand UO_1777 (O_1777,N_29906,N_29800);
nor UO_1778 (O_1778,N_29946,N_29820);
and UO_1779 (O_1779,N_29842,N_29964);
or UO_1780 (O_1780,N_29834,N_29809);
and UO_1781 (O_1781,N_29971,N_29840);
or UO_1782 (O_1782,N_29801,N_29920);
or UO_1783 (O_1783,N_29857,N_29997);
and UO_1784 (O_1784,N_29977,N_29880);
and UO_1785 (O_1785,N_29879,N_29927);
or UO_1786 (O_1786,N_29985,N_29879);
xor UO_1787 (O_1787,N_29819,N_29886);
or UO_1788 (O_1788,N_29906,N_29899);
nand UO_1789 (O_1789,N_29836,N_29801);
xnor UO_1790 (O_1790,N_29848,N_29861);
or UO_1791 (O_1791,N_29996,N_29880);
nor UO_1792 (O_1792,N_29826,N_29958);
nand UO_1793 (O_1793,N_29826,N_29803);
xnor UO_1794 (O_1794,N_29989,N_29872);
nor UO_1795 (O_1795,N_29940,N_29849);
nor UO_1796 (O_1796,N_29900,N_29961);
or UO_1797 (O_1797,N_29969,N_29860);
and UO_1798 (O_1798,N_29995,N_29972);
xnor UO_1799 (O_1799,N_29974,N_29982);
and UO_1800 (O_1800,N_29812,N_29817);
and UO_1801 (O_1801,N_29996,N_29802);
and UO_1802 (O_1802,N_29902,N_29827);
nor UO_1803 (O_1803,N_29894,N_29845);
xnor UO_1804 (O_1804,N_29985,N_29876);
and UO_1805 (O_1805,N_29905,N_29992);
or UO_1806 (O_1806,N_29953,N_29960);
nor UO_1807 (O_1807,N_29868,N_29836);
nand UO_1808 (O_1808,N_29809,N_29954);
or UO_1809 (O_1809,N_29995,N_29968);
xnor UO_1810 (O_1810,N_29929,N_29819);
nand UO_1811 (O_1811,N_29969,N_29939);
or UO_1812 (O_1812,N_29989,N_29978);
or UO_1813 (O_1813,N_29868,N_29966);
xor UO_1814 (O_1814,N_29887,N_29820);
nor UO_1815 (O_1815,N_29937,N_29991);
xor UO_1816 (O_1816,N_29926,N_29821);
xor UO_1817 (O_1817,N_29849,N_29803);
nand UO_1818 (O_1818,N_29872,N_29972);
nand UO_1819 (O_1819,N_29990,N_29899);
and UO_1820 (O_1820,N_29970,N_29812);
xor UO_1821 (O_1821,N_29951,N_29955);
nor UO_1822 (O_1822,N_29820,N_29888);
and UO_1823 (O_1823,N_29802,N_29823);
xnor UO_1824 (O_1824,N_29861,N_29842);
xor UO_1825 (O_1825,N_29977,N_29848);
xnor UO_1826 (O_1826,N_29831,N_29996);
xor UO_1827 (O_1827,N_29955,N_29992);
and UO_1828 (O_1828,N_29892,N_29817);
or UO_1829 (O_1829,N_29950,N_29935);
nand UO_1830 (O_1830,N_29916,N_29933);
nor UO_1831 (O_1831,N_29930,N_29980);
nand UO_1832 (O_1832,N_29920,N_29900);
or UO_1833 (O_1833,N_29894,N_29879);
xor UO_1834 (O_1834,N_29969,N_29856);
and UO_1835 (O_1835,N_29861,N_29839);
or UO_1836 (O_1836,N_29974,N_29999);
nand UO_1837 (O_1837,N_29989,N_29818);
or UO_1838 (O_1838,N_29954,N_29896);
and UO_1839 (O_1839,N_29800,N_29987);
nand UO_1840 (O_1840,N_29855,N_29957);
xnor UO_1841 (O_1841,N_29854,N_29908);
xor UO_1842 (O_1842,N_29860,N_29948);
nor UO_1843 (O_1843,N_29963,N_29922);
nand UO_1844 (O_1844,N_29884,N_29895);
or UO_1845 (O_1845,N_29909,N_29943);
nor UO_1846 (O_1846,N_29870,N_29826);
or UO_1847 (O_1847,N_29875,N_29946);
and UO_1848 (O_1848,N_29833,N_29815);
xnor UO_1849 (O_1849,N_29975,N_29800);
and UO_1850 (O_1850,N_29837,N_29829);
xor UO_1851 (O_1851,N_29841,N_29979);
nand UO_1852 (O_1852,N_29836,N_29914);
xor UO_1853 (O_1853,N_29983,N_29976);
or UO_1854 (O_1854,N_29865,N_29941);
xnor UO_1855 (O_1855,N_29893,N_29826);
or UO_1856 (O_1856,N_29804,N_29941);
nor UO_1857 (O_1857,N_29939,N_29872);
nor UO_1858 (O_1858,N_29806,N_29948);
or UO_1859 (O_1859,N_29906,N_29811);
nor UO_1860 (O_1860,N_29938,N_29990);
or UO_1861 (O_1861,N_29972,N_29873);
xnor UO_1862 (O_1862,N_29858,N_29994);
nor UO_1863 (O_1863,N_29901,N_29886);
and UO_1864 (O_1864,N_29947,N_29960);
or UO_1865 (O_1865,N_29975,N_29952);
nor UO_1866 (O_1866,N_29824,N_29901);
or UO_1867 (O_1867,N_29849,N_29866);
nor UO_1868 (O_1868,N_29827,N_29908);
or UO_1869 (O_1869,N_29929,N_29949);
nand UO_1870 (O_1870,N_29860,N_29882);
nand UO_1871 (O_1871,N_29951,N_29855);
xnor UO_1872 (O_1872,N_29886,N_29899);
nor UO_1873 (O_1873,N_29990,N_29957);
and UO_1874 (O_1874,N_29937,N_29828);
or UO_1875 (O_1875,N_29864,N_29888);
xnor UO_1876 (O_1876,N_29918,N_29833);
nand UO_1877 (O_1877,N_29925,N_29976);
or UO_1878 (O_1878,N_29982,N_29915);
or UO_1879 (O_1879,N_29818,N_29939);
xnor UO_1880 (O_1880,N_29881,N_29913);
and UO_1881 (O_1881,N_29827,N_29802);
or UO_1882 (O_1882,N_29961,N_29964);
nor UO_1883 (O_1883,N_29954,N_29992);
or UO_1884 (O_1884,N_29849,N_29959);
nand UO_1885 (O_1885,N_29910,N_29936);
nor UO_1886 (O_1886,N_29818,N_29964);
nor UO_1887 (O_1887,N_29986,N_29914);
and UO_1888 (O_1888,N_29898,N_29802);
or UO_1889 (O_1889,N_29810,N_29869);
and UO_1890 (O_1890,N_29975,N_29823);
and UO_1891 (O_1891,N_29991,N_29976);
xnor UO_1892 (O_1892,N_29985,N_29935);
nand UO_1893 (O_1893,N_29992,N_29852);
or UO_1894 (O_1894,N_29829,N_29857);
or UO_1895 (O_1895,N_29853,N_29835);
or UO_1896 (O_1896,N_29839,N_29853);
or UO_1897 (O_1897,N_29905,N_29873);
xnor UO_1898 (O_1898,N_29897,N_29942);
and UO_1899 (O_1899,N_29805,N_29956);
nor UO_1900 (O_1900,N_29923,N_29993);
nand UO_1901 (O_1901,N_29896,N_29890);
or UO_1902 (O_1902,N_29816,N_29932);
nand UO_1903 (O_1903,N_29985,N_29930);
or UO_1904 (O_1904,N_29819,N_29906);
and UO_1905 (O_1905,N_29874,N_29974);
nand UO_1906 (O_1906,N_29844,N_29952);
xor UO_1907 (O_1907,N_29860,N_29983);
and UO_1908 (O_1908,N_29862,N_29811);
nand UO_1909 (O_1909,N_29976,N_29827);
and UO_1910 (O_1910,N_29947,N_29973);
xnor UO_1911 (O_1911,N_29900,N_29880);
nor UO_1912 (O_1912,N_29971,N_29960);
and UO_1913 (O_1913,N_29908,N_29945);
nor UO_1914 (O_1914,N_29872,N_29998);
and UO_1915 (O_1915,N_29804,N_29857);
and UO_1916 (O_1916,N_29967,N_29981);
or UO_1917 (O_1917,N_29853,N_29911);
nor UO_1918 (O_1918,N_29987,N_29938);
nand UO_1919 (O_1919,N_29980,N_29808);
nand UO_1920 (O_1920,N_29869,N_29902);
nor UO_1921 (O_1921,N_29906,N_29983);
and UO_1922 (O_1922,N_29980,N_29959);
nor UO_1923 (O_1923,N_29948,N_29884);
xnor UO_1924 (O_1924,N_29924,N_29857);
or UO_1925 (O_1925,N_29823,N_29961);
nand UO_1926 (O_1926,N_29864,N_29841);
xnor UO_1927 (O_1927,N_29889,N_29930);
xor UO_1928 (O_1928,N_29896,N_29945);
nand UO_1929 (O_1929,N_29925,N_29877);
xor UO_1930 (O_1930,N_29851,N_29985);
nor UO_1931 (O_1931,N_29967,N_29813);
or UO_1932 (O_1932,N_29967,N_29891);
nand UO_1933 (O_1933,N_29902,N_29931);
xnor UO_1934 (O_1934,N_29921,N_29975);
nor UO_1935 (O_1935,N_29991,N_29837);
and UO_1936 (O_1936,N_29994,N_29978);
xnor UO_1937 (O_1937,N_29812,N_29937);
nand UO_1938 (O_1938,N_29874,N_29814);
xor UO_1939 (O_1939,N_29934,N_29978);
or UO_1940 (O_1940,N_29860,N_29927);
or UO_1941 (O_1941,N_29851,N_29948);
nand UO_1942 (O_1942,N_29857,N_29968);
nor UO_1943 (O_1943,N_29917,N_29933);
or UO_1944 (O_1944,N_29984,N_29910);
nand UO_1945 (O_1945,N_29886,N_29994);
nor UO_1946 (O_1946,N_29945,N_29932);
or UO_1947 (O_1947,N_29867,N_29888);
xor UO_1948 (O_1948,N_29821,N_29974);
and UO_1949 (O_1949,N_29821,N_29802);
nor UO_1950 (O_1950,N_29910,N_29951);
or UO_1951 (O_1951,N_29883,N_29898);
xnor UO_1952 (O_1952,N_29966,N_29853);
or UO_1953 (O_1953,N_29867,N_29950);
nand UO_1954 (O_1954,N_29923,N_29891);
nor UO_1955 (O_1955,N_29986,N_29826);
nand UO_1956 (O_1956,N_29937,N_29883);
xor UO_1957 (O_1957,N_29844,N_29853);
and UO_1958 (O_1958,N_29925,N_29985);
and UO_1959 (O_1959,N_29920,N_29994);
and UO_1960 (O_1960,N_29918,N_29887);
or UO_1961 (O_1961,N_29824,N_29956);
and UO_1962 (O_1962,N_29979,N_29874);
nand UO_1963 (O_1963,N_29998,N_29956);
and UO_1964 (O_1964,N_29856,N_29948);
nor UO_1965 (O_1965,N_29826,N_29996);
and UO_1966 (O_1966,N_29988,N_29956);
and UO_1967 (O_1967,N_29938,N_29831);
nand UO_1968 (O_1968,N_29915,N_29966);
and UO_1969 (O_1969,N_29906,N_29956);
xor UO_1970 (O_1970,N_29930,N_29902);
nand UO_1971 (O_1971,N_29844,N_29895);
nor UO_1972 (O_1972,N_29850,N_29869);
and UO_1973 (O_1973,N_29850,N_29926);
or UO_1974 (O_1974,N_29934,N_29975);
and UO_1975 (O_1975,N_29836,N_29942);
and UO_1976 (O_1976,N_29835,N_29988);
nand UO_1977 (O_1977,N_29973,N_29931);
nor UO_1978 (O_1978,N_29981,N_29882);
or UO_1979 (O_1979,N_29903,N_29944);
or UO_1980 (O_1980,N_29969,N_29821);
nand UO_1981 (O_1981,N_29830,N_29988);
and UO_1982 (O_1982,N_29816,N_29933);
xnor UO_1983 (O_1983,N_29877,N_29873);
or UO_1984 (O_1984,N_29995,N_29825);
xor UO_1985 (O_1985,N_29949,N_29915);
xor UO_1986 (O_1986,N_29825,N_29851);
and UO_1987 (O_1987,N_29835,N_29808);
or UO_1988 (O_1988,N_29878,N_29970);
or UO_1989 (O_1989,N_29868,N_29943);
nor UO_1990 (O_1990,N_29998,N_29860);
nand UO_1991 (O_1991,N_29942,N_29837);
and UO_1992 (O_1992,N_29991,N_29954);
nor UO_1993 (O_1993,N_29973,N_29864);
or UO_1994 (O_1994,N_29898,N_29900);
or UO_1995 (O_1995,N_29899,N_29943);
nand UO_1996 (O_1996,N_29828,N_29820);
nor UO_1997 (O_1997,N_29913,N_29952);
and UO_1998 (O_1998,N_29923,N_29982);
and UO_1999 (O_1999,N_29806,N_29937);
and UO_2000 (O_2000,N_29876,N_29956);
and UO_2001 (O_2001,N_29822,N_29870);
nand UO_2002 (O_2002,N_29906,N_29873);
and UO_2003 (O_2003,N_29843,N_29919);
and UO_2004 (O_2004,N_29823,N_29800);
nor UO_2005 (O_2005,N_29931,N_29994);
or UO_2006 (O_2006,N_29812,N_29906);
nor UO_2007 (O_2007,N_29900,N_29941);
nand UO_2008 (O_2008,N_29837,N_29958);
nor UO_2009 (O_2009,N_29862,N_29887);
or UO_2010 (O_2010,N_29990,N_29925);
nor UO_2011 (O_2011,N_29808,N_29932);
nor UO_2012 (O_2012,N_29914,N_29877);
nor UO_2013 (O_2013,N_29972,N_29953);
and UO_2014 (O_2014,N_29876,N_29868);
xor UO_2015 (O_2015,N_29830,N_29923);
or UO_2016 (O_2016,N_29930,N_29812);
and UO_2017 (O_2017,N_29966,N_29909);
nor UO_2018 (O_2018,N_29898,N_29817);
and UO_2019 (O_2019,N_29991,N_29871);
nor UO_2020 (O_2020,N_29965,N_29820);
xor UO_2021 (O_2021,N_29824,N_29902);
nor UO_2022 (O_2022,N_29987,N_29805);
and UO_2023 (O_2023,N_29820,N_29863);
nand UO_2024 (O_2024,N_29811,N_29981);
xnor UO_2025 (O_2025,N_29945,N_29968);
xor UO_2026 (O_2026,N_29870,N_29848);
nand UO_2027 (O_2027,N_29875,N_29832);
nand UO_2028 (O_2028,N_29862,N_29899);
or UO_2029 (O_2029,N_29938,N_29936);
xnor UO_2030 (O_2030,N_29998,N_29930);
or UO_2031 (O_2031,N_29986,N_29869);
or UO_2032 (O_2032,N_29933,N_29804);
nor UO_2033 (O_2033,N_29984,N_29913);
and UO_2034 (O_2034,N_29983,N_29928);
nand UO_2035 (O_2035,N_29889,N_29869);
nor UO_2036 (O_2036,N_29880,N_29947);
xnor UO_2037 (O_2037,N_29865,N_29957);
or UO_2038 (O_2038,N_29995,N_29824);
or UO_2039 (O_2039,N_29949,N_29965);
nand UO_2040 (O_2040,N_29818,N_29990);
and UO_2041 (O_2041,N_29822,N_29931);
and UO_2042 (O_2042,N_29901,N_29845);
nand UO_2043 (O_2043,N_29817,N_29923);
xor UO_2044 (O_2044,N_29984,N_29926);
or UO_2045 (O_2045,N_29959,N_29823);
and UO_2046 (O_2046,N_29810,N_29860);
and UO_2047 (O_2047,N_29815,N_29862);
nand UO_2048 (O_2048,N_29955,N_29813);
xor UO_2049 (O_2049,N_29971,N_29868);
nand UO_2050 (O_2050,N_29878,N_29856);
nand UO_2051 (O_2051,N_29816,N_29879);
nand UO_2052 (O_2052,N_29953,N_29881);
or UO_2053 (O_2053,N_29930,N_29803);
nor UO_2054 (O_2054,N_29938,N_29826);
xnor UO_2055 (O_2055,N_29964,N_29948);
nor UO_2056 (O_2056,N_29801,N_29968);
nand UO_2057 (O_2057,N_29808,N_29988);
nor UO_2058 (O_2058,N_29925,N_29953);
nand UO_2059 (O_2059,N_29996,N_29864);
and UO_2060 (O_2060,N_29973,N_29868);
or UO_2061 (O_2061,N_29963,N_29977);
xor UO_2062 (O_2062,N_29903,N_29856);
or UO_2063 (O_2063,N_29994,N_29983);
or UO_2064 (O_2064,N_29924,N_29957);
xor UO_2065 (O_2065,N_29876,N_29822);
xor UO_2066 (O_2066,N_29947,N_29987);
and UO_2067 (O_2067,N_29804,N_29971);
and UO_2068 (O_2068,N_29975,N_29854);
nor UO_2069 (O_2069,N_29976,N_29885);
xor UO_2070 (O_2070,N_29864,N_29902);
xor UO_2071 (O_2071,N_29972,N_29974);
nor UO_2072 (O_2072,N_29958,N_29946);
nand UO_2073 (O_2073,N_29942,N_29848);
nor UO_2074 (O_2074,N_29894,N_29979);
nor UO_2075 (O_2075,N_29912,N_29916);
nand UO_2076 (O_2076,N_29843,N_29898);
and UO_2077 (O_2077,N_29914,N_29923);
nor UO_2078 (O_2078,N_29989,N_29929);
and UO_2079 (O_2079,N_29960,N_29895);
and UO_2080 (O_2080,N_29969,N_29914);
nor UO_2081 (O_2081,N_29958,N_29921);
xnor UO_2082 (O_2082,N_29874,N_29803);
or UO_2083 (O_2083,N_29925,N_29938);
xor UO_2084 (O_2084,N_29870,N_29843);
nand UO_2085 (O_2085,N_29835,N_29952);
nand UO_2086 (O_2086,N_29937,N_29898);
xnor UO_2087 (O_2087,N_29863,N_29937);
or UO_2088 (O_2088,N_29842,N_29987);
and UO_2089 (O_2089,N_29956,N_29873);
nand UO_2090 (O_2090,N_29884,N_29839);
nand UO_2091 (O_2091,N_29814,N_29885);
nand UO_2092 (O_2092,N_29996,N_29917);
and UO_2093 (O_2093,N_29957,N_29984);
nor UO_2094 (O_2094,N_29960,N_29976);
nor UO_2095 (O_2095,N_29810,N_29972);
nor UO_2096 (O_2096,N_29844,N_29801);
xnor UO_2097 (O_2097,N_29852,N_29813);
and UO_2098 (O_2098,N_29892,N_29855);
and UO_2099 (O_2099,N_29835,N_29925);
nor UO_2100 (O_2100,N_29887,N_29974);
nor UO_2101 (O_2101,N_29862,N_29894);
nand UO_2102 (O_2102,N_29899,N_29805);
xor UO_2103 (O_2103,N_29878,N_29883);
nand UO_2104 (O_2104,N_29845,N_29998);
xnor UO_2105 (O_2105,N_29923,N_29862);
and UO_2106 (O_2106,N_29927,N_29996);
or UO_2107 (O_2107,N_29950,N_29964);
nand UO_2108 (O_2108,N_29968,N_29985);
nand UO_2109 (O_2109,N_29892,N_29909);
nor UO_2110 (O_2110,N_29911,N_29828);
nand UO_2111 (O_2111,N_29899,N_29881);
or UO_2112 (O_2112,N_29919,N_29880);
xnor UO_2113 (O_2113,N_29842,N_29817);
nand UO_2114 (O_2114,N_29941,N_29944);
xnor UO_2115 (O_2115,N_29973,N_29990);
nor UO_2116 (O_2116,N_29910,N_29877);
nand UO_2117 (O_2117,N_29872,N_29828);
xor UO_2118 (O_2118,N_29873,N_29993);
nand UO_2119 (O_2119,N_29867,N_29898);
nor UO_2120 (O_2120,N_29952,N_29989);
and UO_2121 (O_2121,N_29822,N_29889);
nand UO_2122 (O_2122,N_29970,N_29884);
xor UO_2123 (O_2123,N_29940,N_29900);
xnor UO_2124 (O_2124,N_29906,N_29814);
xnor UO_2125 (O_2125,N_29982,N_29929);
or UO_2126 (O_2126,N_29856,N_29967);
and UO_2127 (O_2127,N_29884,N_29902);
xnor UO_2128 (O_2128,N_29825,N_29926);
and UO_2129 (O_2129,N_29954,N_29823);
and UO_2130 (O_2130,N_29873,N_29939);
or UO_2131 (O_2131,N_29920,N_29978);
nor UO_2132 (O_2132,N_29884,N_29806);
nand UO_2133 (O_2133,N_29918,N_29829);
nand UO_2134 (O_2134,N_29999,N_29905);
or UO_2135 (O_2135,N_29800,N_29834);
nor UO_2136 (O_2136,N_29909,N_29893);
nor UO_2137 (O_2137,N_29912,N_29906);
or UO_2138 (O_2138,N_29915,N_29943);
nor UO_2139 (O_2139,N_29955,N_29918);
and UO_2140 (O_2140,N_29898,N_29935);
and UO_2141 (O_2141,N_29884,N_29844);
and UO_2142 (O_2142,N_29901,N_29847);
nand UO_2143 (O_2143,N_29811,N_29807);
nor UO_2144 (O_2144,N_29824,N_29890);
nand UO_2145 (O_2145,N_29876,N_29962);
or UO_2146 (O_2146,N_29899,N_29828);
xnor UO_2147 (O_2147,N_29906,N_29866);
nand UO_2148 (O_2148,N_29858,N_29853);
and UO_2149 (O_2149,N_29826,N_29841);
or UO_2150 (O_2150,N_29925,N_29999);
xor UO_2151 (O_2151,N_29871,N_29817);
or UO_2152 (O_2152,N_29905,N_29930);
nand UO_2153 (O_2153,N_29846,N_29937);
and UO_2154 (O_2154,N_29873,N_29986);
nor UO_2155 (O_2155,N_29975,N_29997);
and UO_2156 (O_2156,N_29928,N_29976);
xnor UO_2157 (O_2157,N_29946,N_29994);
and UO_2158 (O_2158,N_29882,N_29910);
or UO_2159 (O_2159,N_29821,N_29963);
or UO_2160 (O_2160,N_29875,N_29959);
and UO_2161 (O_2161,N_29885,N_29922);
nor UO_2162 (O_2162,N_29833,N_29813);
and UO_2163 (O_2163,N_29964,N_29863);
or UO_2164 (O_2164,N_29933,N_29934);
or UO_2165 (O_2165,N_29892,N_29954);
and UO_2166 (O_2166,N_29910,N_29941);
nor UO_2167 (O_2167,N_29810,N_29904);
and UO_2168 (O_2168,N_29818,N_29838);
and UO_2169 (O_2169,N_29810,N_29951);
or UO_2170 (O_2170,N_29803,N_29885);
and UO_2171 (O_2171,N_29915,N_29828);
nor UO_2172 (O_2172,N_29876,N_29949);
nor UO_2173 (O_2173,N_29988,N_29813);
or UO_2174 (O_2174,N_29904,N_29814);
and UO_2175 (O_2175,N_29817,N_29820);
nor UO_2176 (O_2176,N_29830,N_29945);
or UO_2177 (O_2177,N_29943,N_29953);
nor UO_2178 (O_2178,N_29826,N_29985);
xnor UO_2179 (O_2179,N_29963,N_29825);
nand UO_2180 (O_2180,N_29885,N_29851);
or UO_2181 (O_2181,N_29900,N_29980);
nand UO_2182 (O_2182,N_29920,N_29979);
and UO_2183 (O_2183,N_29885,N_29967);
or UO_2184 (O_2184,N_29809,N_29975);
nand UO_2185 (O_2185,N_29861,N_29897);
nor UO_2186 (O_2186,N_29928,N_29905);
xnor UO_2187 (O_2187,N_29915,N_29901);
nor UO_2188 (O_2188,N_29940,N_29831);
nor UO_2189 (O_2189,N_29948,N_29989);
and UO_2190 (O_2190,N_29893,N_29836);
and UO_2191 (O_2191,N_29882,N_29820);
and UO_2192 (O_2192,N_29854,N_29890);
nor UO_2193 (O_2193,N_29824,N_29954);
nand UO_2194 (O_2194,N_29954,N_29875);
nor UO_2195 (O_2195,N_29924,N_29852);
nor UO_2196 (O_2196,N_29971,N_29979);
or UO_2197 (O_2197,N_29834,N_29970);
and UO_2198 (O_2198,N_29890,N_29909);
and UO_2199 (O_2199,N_29948,N_29889);
and UO_2200 (O_2200,N_29966,N_29872);
or UO_2201 (O_2201,N_29836,N_29968);
and UO_2202 (O_2202,N_29808,N_29975);
and UO_2203 (O_2203,N_29921,N_29854);
or UO_2204 (O_2204,N_29932,N_29939);
nor UO_2205 (O_2205,N_29915,N_29919);
xor UO_2206 (O_2206,N_29990,N_29977);
and UO_2207 (O_2207,N_29999,N_29854);
and UO_2208 (O_2208,N_29928,N_29852);
or UO_2209 (O_2209,N_29864,N_29969);
nand UO_2210 (O_2210,N_29914,N_29935);
xor UO_2211 (O_2211,N_29893,N_29851);
nand UO_2212 (O_2212,N_29903,N_29811);
nor UO_2213 (O_2213,N_29836,N_29867);
xnor UO_2214 (O_2214,N_29888,N_29881);
or UO_2215 (O_2215,N_29863,N_29910);
and UO_2216 (O_2216,N_29979,N_29812);
or UO_2217 (O_2217,N_29930,N_29887);
and UO_2218 (O_2218,N_29895,N_29813);
nand UO_2219 (O_2219,N_29969,N_29853);
xor UO_2220 (O_2220,N_29945,N_29967);
and UO_2221 (O_2221,N_29925,N_29964);
and UO_2222 (O_2222,N_29928,N_29907);
and UO_2223 (O_2223,N_29903,N_29906);
and UO_2224 (O_2224,N_29985,N_29802);
or UO_2225 (O_2225,N_29958,N_29903);
and UO_2226 (O_2226,N_29835,N_29814);
or UO_2227 (O_2227,N_29963,N_29936);
nor UO_2228 (O_2228,N_29852,N_29994);
xnor UO_2229 (O_2229,N_29981,N_29829);
nor UO_2230 (O_2230,N_29917,N_29983);
and UO_2231 (O_2231,N_29973,N_29857);
nor UO_2232 (O_2232,N_29933,N_29844);
xor UO_2233 (O_2233,N_29920,N_29889);
xnor UO_2234 (O_2234,N_29862,N_29962);
xnor UO_2235 (O_2235,N_29879,N_29943);
nor UO_2236 (O_2236,N_29939,N_29858);
xor UO_2237 (O_2237,N_29871,N_29844);
nor UO_2238 (O_2238,N_29970,N_29979);
or UO_2239 (O_2239,N_29889,N_29913);
xor UO_2240 (O_2240,N_29838,N_29852);
xnor UO_2241 (O_2241,N_29860,N_29905);
or UO_2242 (O_2242,N_29820,N_29961);
xor UO_2243 (O_2243,N_29866,N_29949);
nor UO_2244 (O_2244,N_29995,N_29819);
nor UO_2245 (O_2245,N_29976,N_29906);
and UO_2246 (O_2246,N_29909,N_29821);
nor UO_2247 (O_2247,N_29856,N_29808);
and UO_2248 (O_2248,N_29819,N_29888);
and UO_2249 (O_2249,N_29994,N_29981);
and UO_2250 (O_2250,N_29801,N_29872);
and UO_2251 (O_2251,N_29832,N_29951);
and UO_2252 (O_2252,N_29850,N_29843);
nor UO_2253 (O_2253,N_29802,N_29958);
nor UO_2254 (O_2254,N_29967,N_29986);
nor UO_2255 (O_2255,N_29927,N_29983);
nor UO_2256 (O_2256,N_29850,N_29966);
xor UO_2257 (O_2257,N_29850,N_29914);
or UO_2258 (O_2258,N_29853,N_29942);
and UO_2259 (O_2259,N_29886,N_29976);
and UO_2260 (O_2260,N_29874,N_29832);
or UO_2261 (O_2261,N_29996,N_29982);
nor UO_2262 (O_2262,N_29993,N_29970);
and UO_2263 (O_2263,N_29936,N_29856);
nand UO_2264 (O_2264,N_29907,N_29968);
or UO_2265 (O_2265,N_29864,N_29885);
or UO_2266 (O_2266,N_29921,N_29816);
and UO_2267 (O_2267,N_29870,N_29867);
nand UO_2268 (O_2268,N_29906,N_29941);
or UO_2269 (O_2269,N_29884,N_29891);
nor UO_2270 (O_2270,N_29974,N_29826);
or UO_2271 (O_2271,N_29860,N_29982);
or UO_2272 (O_2272,N_29976,N_29959);
nand UO_2273 (O_2273,N_29898,N_29946);
nand UO_2274 (O_2274,N_29992,N_29941);
nand UO_2275 (O_2275,N_29983,N_29919);
xor UO_2276 (O_2276,N_29822,N_29959);
xnor UO_2277 (O_2277,N_29943,N_29947);
nor UO_2278 (O_2278,N_29806,N_29843);
or UO_2279 (O_2279,N_29979,N_29992);
nand UO_2280 (O_2280,N_29961,N_29922);
or UO_2281 (O_2281,N_29808,N_29886);
nor UO_2282 (O_2282,N_29992,N_29807);
nor UO_2283 (O_2283,N_29902,N_29818);
nor UO_2284 (O_2284,N_29914,N_29975);
nand UO_2285 (O_2285,N_29802,N_29825);
and UO_2286 (O_2286,N_29816,N_29862);
xor UO_2287 (O_2287,N_29845,N_29949);
or UO_2288 (O_2288,N_29805,N_29837);
xor UO_2289 (O_2289,N_29940,N_29943);
or UO_2290 (O_2290,N_29902,N_29811);
nor UO_2291 (O_2291,N_29805,N_29851);
nor UO_2292 (O_2292,N_29951,N_29938);
or UO_2293 (O_2293,N_29920,N_29916);
nor UO_2294 (O_2294,N_29915,N_29847);
nand UO_2295 (O_2295,N_29857,N_29970);
and UO_2296 (O_2296,N_29991,N_29870);
nor UO_2297 (O_2297,N_29924,N_29941);
and UO_2298 (O_2298,N_29828,N_29847);
or UO_2299 (O_2299,N_29809,N_29910);
or UO_2300 (O_2300,N_29809,N_29959);
nor UO_2301 (O_2301,N_29973,N_29813);
and UO_2302 (O_2302,N_29982,N_29984);
and UO_2303 (O_2303,N_29848,N_29880);
and UO_2304 (O_2304,N_29863,N_29967);
and UO_2305 (O_2305,N_29875,N_29939);
nor UO_2306 (O_2306,N_29997,N_29961);
nand UO_2307 (O_2307,N_29947,N_29867);
xor UO_2308 (O_2308,N_29844,N_29970);
and UO_2309 (O_2309,N_29893,N_29821);
nor UO_2310 (O_2310,N_29911,N_29838);
nand UO_2311 (O_2311,N_29960,N_29827);
nand UO_2312 (O_2312,N_29809,N_29871);
nand UO_2313 (O_2313,N_29982,N_29899);
nor UO_2314 (O_2314,N_29949,N_29851);
xor UO_2315 (O_2315,N_29927,N_29857);
or UO_2316 (O_2316,N_29948,N_29934);
xor UO_2317 (O_2317,N_29914,N_29867);
xnor UO_2318 (O_2318,N_29977,N_29821);
nand UO_2319 (O_2319,N_29882,N_29915);
nor UO_2320 (O_2320,N_29966,N_29830);
nor UO_2321 (O_2321,N_29887,N_29811);
xor UO_2322 (O_2322,N_29910,N_29862);
nand UO_2323 (O_2323,N_29877,N_29980);
nand UO_2324 (O_2324,N_29994,N_29990);
nor UO_2325 (O_2325,N_29861,N_29863);
xnor UO_2326 (O_2326,N_29864,N_29926);
xnor UO_2327 (O_2327,N_29877,N_29983);
xnor UO_2328 (O_2328,N_29871,N_29812);
or UO_2329 (O_2329,N_29874,N_29890);
and UO_2330 (O_2330,N_29828,N_29976);
xnor UO_2331 (O_2331,N_29960,N_29874);
xnor UO_2332 (O_2332,N_29989,N_29918);
xor UO_2333 (O_2333,N_29893,N_29874);
and UO_2334 (O_2334,N_29973,N_29891);
xor UO_2335 (O_2335,N_29871,N_29967);
or UO_2336 (O_2336,N_29894,N_29803);
nand UO_2337 (O_2337,N_29995,N_29850);
and UO_2338 (O_2338,N_29852,N_29845);
nand UO_2339 (O_2339,N_29878,N_29910);
xor UO_2340 (O_2340,N_29982,N_29991);
and UO_2341 (O_2341,N_29856,N_29839);
and UO_2342 (O_2342,N_29808,N_29878);
and UO_2343 (O_2343,N_29897,N_29948);
xnor UO_2344 (O_2344,N_29825,N_29864);
nor UO_2345 (O_2345,N_29839,N_29909);
nand UO_2346 (O_2346,N_29872,N_29816);
nand UO_2347 (O_2347,N_29853,N_29843);
or UO_2348 (O_2348,N_29889,N_29854);
and UO_2349 (O_2349,N_29845,N_29880);
nor UO_2350 (O_2350,N_29900,N_29910);
nand UO_2351 (O_2351,N_29831,N_29824);
or UO_2352 (O_2352,N_29868,N_29991);
nor UO_2353 (O_2353,N_29885,N_29942);
xnor UO_2354 (O_2354,N_29997,N_29927);
xor UO_2355 (O_2355,N_29814,N_29849);
nor UO_2356 (O_2356,N_29854,N_29904);
xnor UO_2357 (O_2357,N_29862,N_29819);
nand UO_2358 (O_2358,N_29962,N_29919);
and UO_2359 (O_2359,N_29952,N_29823);
xnor UO_2360 (O_2360,N_29996,N_29936);
nand UO_2361 (O_2361,N_29856,N_29953);
nor UO_2362 (O_2362,N_29838,N_29961);
and UO_2363 (O_2363,N_29959,N_29842);
xnor UO_2364 (O_2364,N_29861,N_29905);
xor UO_2365 (O_2365,N_29890,N_29846);
nand UO_2366 (O_2366,N_29978,N_29858);
nor UO_2367 (O_2367,N_29997,N_29813);
nand UO_2368 (O_2368,N_29920,N_29879);
nand UO_2369 (O_2369,N_29855,N_29848);
xor UO_2370 (O_2370,N_29978,N_29969);
and UO_2371 (O_2371,N_29835,N_29869);
or UO_2372 (O_2372,N_29885,N_29940);
and UO_2373 (O_2373,N_29929,N_29859);
xor UO_2374 (O_2374,N_29923,N_29990);
or UO_2375 (O_2375,N_29831,N_29933);
and UO_2376 (O_2376,N_29898,N_29995);
nand UO_2377 (O_2377,N_29809,N_29919);
and UO_2378 (O_2378,N_29936,N_29822);
nand UO_2379 (O_2379,N_29951,N_29913);
xor UO_2380 (O_2380,N_29886,N_29917);
xnor UO_2381 (O_2381,N_29887,N_29903);
xor UO_2382 (O_2382,N_29881,N_29934);
or UO_2383 (O_2383,N_29936,N_29847);
or UO_2384 (O_2384,N_29938,N_29899);
or UO_2385 (O_2385,N_29938,N_29971);
and UO_2386 (O_2386,N_29855,N_29931);
nand UO_2387 (O_2387,N_29868,N_29934);
nand UO_2388 (O_2388,N_29968,N_29959);
or UO_2389 (O_2389,N_29800,N_29847);
nor UO_2390 (O_2390,N_29815,N_29963);
and UO_2391 (O_2391,N_29925,N_29940);
nand UO_2392 (O_2392,N_29987,N_29917);
or UO_2393 (O_2393,N_29876,N_29914);
nor UO_2394 (O_2394,N_29903,N_29953);
and UO_2395 (O_2395,N_29974,N_29861);
xnor UO_2396 (O_2396,N_29874,N_29845);
xnor UO_2397 (O_2397,N_29980,N_29840);
and UO_2398 (O_2398,N_29907,N_29972);
and UO_2399 (O_2399,N_29872,N_29958);
and UO_2400 (O_2400,N_29869,N_29948);
nand UO_2401 (O_2401,N_29865,N_29951);
nand UO_2402 (O_2402,N_29839,N_29867);
xnor UO_2403 (O_2403,N_29849,N_29840);
xor UO_2404 (O_2404,N_29998,N_29982);
nand UO_2405 (O_2405,N_29927,N_29970);
nor UO_2406 (O_2406,N_29997,N_29938);
nor UO_2407 (O_2407,N_29873,N_29860);
and UO_2408 (O_2408,N_29893,N_29899);
or UO_2409 (O_2409,N_29977,N_29894);
and UO_2410 (O_2410,N_29951,N_29843);
and UO_2411 (O_2411,N_29874,N_29813);
nor UO_2412 (O_2412,N_29919,N_29927);
nor UO_2413 (O_2413,N_29974,N_29978);
nor UO_2414 (O_2414,N_29813,N_29928);
or UO_2415 (O_2415,N_29992,N_29857);
or UO_2416 (O_2416,N_29838,N_29906);
nand UO_2417 (O_2417,N_29882,N_29944);
xnor UO_2418 (O_2418,N_29864,N_29954);
xnor UO_2419 (O_2419,N_29937,N_29861);
nand UO_2420 (O_2420,N_29904,N_29908);
xor UO_2421 (O_2421,N_29805,N_29893);
or UO_2422 (O_2422,N_29957,N_29965);
or UO_2423 (O_2423,N_29999,N_29979);
or UO_2424 (O_2424,N_29913,N_29934);
nor UO_2425 (O_2425,N_29809,N_29807);
nor UO_2426 (O_2426,N_29944,N_29823);
and UO_2427 (O_2427,N_29958,N_29985);
or UO_2428 (O_2428,N_29986,N_29843);
xnor UO_2429 (O_2429,N_29987,N_29886);
or UO_2430 (O_2430,N_29852,N_29853);
nand UO_2431 (O_2431,N_29971,N_29859);
xor UO_2432 (O_2432,N_29908,N_29874);
nor UO_2433 (O_2433,N_29863,N_29807);
or UO_2434 (O_2434,N_29956,N_29912);
nor UO_2435 (O_2435,N_29987,N_29916);
xor UO_2436 (O_2436,N_29803,N_29845);
and UO_2437 (O_2437,N_29804,N_29848);
and UO_2438 (O_2438,N_29882,N_29900);
xnor UO_2439 (O_2439,N_29881,N_29918);
xnor UO_2440 (O_2440,N_29975,N_29833);
and UO_2441 (O_2441,N_29876,N_29950);
nor UO_2442 (O_2442,N_29939,N_29801);
and UO_2443 (O_2443,N_29994,N_29862);
or UO_2444 (O_2444,N_29919,N_29837);
xor UO_2445 (O_2445,N_29864,N_29964);
nand UO_2446 (O_2446,N_29879,N_29986);
or UO_2447 (O_2447,N_29885,N_29901);
nand UO_2448 (O_2448,N_29818,N_29816);
and UO_2449 (O_2449,N_29995,N_29851);
nand UO_2450 (O_2450,N_29926,N_29985);
or UO_2451 (O_2451,N_29938,N_29884);
nand UO_2452 (O_2452,N_29934,N_29946);
or UO_2453 (O_2453,N_29837,N_29862);
xor UO_2454 (O_2454,N_29895,N_29997);
nand UO_2455 (O_2455,N_29940,N_29945);
nor UO_2456 (O_2456,N_29863,N_29875);
and UO_2457 (O_2457,N_29991,N_29929);
xor UO_2458 (O_2458,N_29873,N_29868);
nand UO_2459 (O_2459,N_29889,N_29941);
nor UO_2460 (O_2460,N_29809,N_29957);
or UO_2461 (O_2461,N_29847,N_29806);
nor UO_2462 (O_2462,N_29852,N_29916);
and UO_2463 (O_2463,N_29834,N_29922);
nand UO_2464 (O_2464,N_29823,N_29935);
xor UO_2465 (O_2465,N_29931,N_29953);
and UO_2466 (O_2466,N_29923,N_29842);
nand UO_2467 (O_2467,N_29830,N_29929);
nand UO_2468 (O_2468,N_29808,N_29895);
nand UO_2469 (O_2469,N_29998,N_29920);
nand UO_2470 (O_2470,N_29924,N_29950);
nor UO_2471 (O_2471,N_29951,N_29874);
xnor UO_2472 (O_2472,N_29980,N_29874);
and UO_2473 (O_2473,N_29878,N_29909);
nor UO_2474 (O_2474,N_29955,N_29902);
nand UO_2475 (O_2475,N_29808,N_29804);
and UO_2476 (O_2476,N_29943,N_29855);
and UO_2477 (O_2477,N_29880,N_29935);
nand UO_2478 (O_2478,N_29829,N_29898);
nand UO_2479 (O_2479,N_29932,N_29948);
and UO_2480 (O_2480,N_29908,N_29870);
nand UO_2481 (O_2481,N_29993,N_29992);
xnor UO_2482 (O_2482,N_29963,N_29944);
nand UO_2483 (O_2483,N_29930,N_29829);
xnor UO_2484 (O_2484,N_29865,N_29846);
nor UO_2485 (O_2485,N_29937,N_29990);
and UO_2486 (O_2486,N_29853,N_29857);
or UO_2487 (O_2487,N_29993,N_29801);
or UO_2488 (O_2488,N_29847,N_29865);
nor UO_2489 (O_2489,N_29920,N_29982);
nor UO_2490 (O_2490,N_29922,N_29854);
xor UO_2491 (O_2491,N_29832,N_29943);
nand UO_2492 (O_2492,N_29983,N_29871);
nor UO_2493 (O_2493,N_29951,N_29877);
and UO_2494 (O_2494,N_29859,N_29803);
nor UO_2495 (O_2495,N_29809,N_29912);
nor UO_2496 (O_2496,N_29921,N_29815);
nand UO_2497 (O_2497,N_29993,N_29860);
and UO_2498 (O_2498,N_29810,N_29839);
and UO_2499 (O_2499,N_29986,N_29810);
nor UO_2500 (O_2500,N_29957,N_29926);
xnor UO_2501 (O_2501,N_29921,N_29915);
xor UO_2502 (O_2502,N_29809,N_29945);
nand UO_2503 (O_2503,N_29923,N_29848);
xor UO_2504 (O_2504,N_29897,N_29959);
xor UO_2505 (O_2505,N_29961,N_29825);
or UO_2506 (O_2506,N_29922,N_29803);
xnor UO_2507 (O_2507,N_29998,N_29941);
nand UO_2508 (O_2508,N_29935,N_29903);
and UO_2509 (O_2509,N_29821,N_29887);
nand UO_2510 (O_2510,N_29806,N_29968);
xnor UO_2511 (O_2511,N_29881,N_29835);
or UO_2512 (O_2512,N_29926,N_29830);
or UO_2513 (O_2513,N_29801,N_29862);
xor UO_2514 (O_2514,N_29968,N_29931);
nor UO_2515 (O_2515,N_29895,N_29833);
nor UO_2516 (O_2516,N_29883,N_29901);
xor UO_2517 (O_2517,N_29967,N_29821);
and UO_2518 (O_2518,N_29909,N_29997);
nand UO_2519 (O_2519,N_29977,N_29812);
or UO_2520 (O_2520,N_29938,N_29941);
and UO_2521 (O_2521,N_29909,N_29849);
and UO_2522 (O_2522,N_29987,N_29953);
xnor UO_2523 (O_2523,N_29903,N_29945);
nand UO_2524 (O_2524,N_29931,N_29896);
or UO_2525 (O_2525,N_29815,N_29990);
or UO_2526 (O_2526,N_29856,N_29827);
nand UO_2527 (O_2527,N_29903,N_29990);
and UO_2528 (O_2528,N_29817,N_29802);
nor UO_2529 (O_2529,N_29981,N_29902);
nand UO_2530 (O_2530,N_29849,N_29893);
xnor UO_2531 (O_2531,N_29968,N_29890);
nor UO_2532 (O_2532,N_29823,N_29826);
nand UO_2533 (O_2533,N_29968,N_29906);
xor UO_2534 (O_2534,N_29963,N_29864);
and UO_2535 (O_2535,N_29945,N_29931);
and UO_2536 (O_2536,N_29876,N_29860);
nand UO_2537 (O_2537,N_29897,N_29863);
or UO_2538 (O_2538,N_29814,N_29866);
nor UO_2539 (O_2539,N_29808,N_29815);
and UO_2540 (O_2540,N_29938,N_29980);
or UO_2541 (O_2541,N_29998,N_29802);
and UO_2542 (O_2542,N_29836,N_29918);
and UO_2543 (O_2543,N_29939,N_29840);
xor UO_2544 (O_2544,N_29949,N_29944);
xor UO_2545 (O_2545,N_29811,N_29856);
or UO_2546 (O_2546,N_29810,N_29803);
and UO_2547 (O_2547,N_29973,N_29988);
nor UO_2548 (O_2548,N_29852,N_29929);
or UO_2549 (O_2549,N_29910,N_29990);
nor UO_2550 (O_2550,N_29827,N_29990);
nor UO_2551 (O_2551,N_29852,N_29953);
nor UO_2552 (O_2552,N_29851,N_29853);
nand UO_2553 (O_2553,N_29973,N_29873);
and UO_2554 (O_2554,N_29984,N_29939);
or UO_2555 (O_2555,N_29805,N_29896);
nor UO_2556 (O_2556,N_29965,N_29894);
and UO_2557 (O_2557,N_29856,N_29891);
and UO_2558 (O_2558,N_29905,N_29957);
xnor UO_2559 (O_2559,N_29957,N_29951);
and UO_2560 (O_2560,N_29978,N_29882);
nor UO_2561 (O_2561,N_29951,N_29830);
and UO_2562 (O_2562,N_29887,N_29980);
nand UO_2563 (O_2563,N_29938,N_29896);
nor UO_2564 (O_2564,N_29828,N_29945);
xor UO_2565 (O_2565,N_29804,N_29888);
nor UO_2566 (O_2566,N_29887,N_29848);
xor UO_2567 (O_2567,N_29956,N_29911);
nor UO_2568 (O_2568,N_29865,N_29967);
or UO_2569 (O_2569,N_29880,N_29978);
nand UO_2570 (O_2570,N_29832,N_29944);
nor UO_2571 (O_2571,N_29896,N_29860);
nand UO_2572 (O_2572,N_29808,N_29870);
or UO_2573 (O_2573,N_29852,N_29869);
xnor UO_2574 (O_2574,N_29889,N_29896);
xor UO_2575 (O_2575,N_29842,N_29950);
and UO_2576 (O_2576,N_29913,N_29994);
or UO_2577 (O_2577,N_29932,N_29838);
xor UO_2578 (O_2578,N_29827,N_29817);
or UO_2579 (O_2579,N_29824,N_29973);
nand UO_2580 (O_2580,N_29923,N_29824);
or UO_2581 (O_2581,N_29988,N_29952);
xor UO_2582 (O_2582,N_29864,N_29890);
and UO_2583 (O_2583,N_29832,N_29911);
and UO_2584 (O_2584,N_29871,N_29853);
nor UO_2585 (O_2585,N_29842,N_29995);
nand UO_2586 (O_2586,N_29952,N_29972);
nor UO_2587 (O_2587,N_29866,N_29804);
and UO_2588 (O_2588,N_29827,N_29873);
nor UO_2589 (O_2589,N_29890,N_29937);
or UO_2590 (O_2590,N_29966,N_29874);
and UO_2591 (O_2591,N_29989,N_29838);
xnor UO_2592 (O_2592,N_29979,N_29808);
and UO_2593 (O_2593,N_29908,N_29919);
or UO_2594 (O_2594,N_29930,N_29871);
or UO_2595 (O_2595,N_29949,N_29878);
xnor UO_2596 (O_2596,N_29958,N_29978);
nand UO_2597 (O_2597,N_29800,N_29845);
xor UO_2598 (O_2598,N_29823,N_29929);
nor UO_2599 (O_2599,N_29986,N_29866);
nand UO_2600 (O_2600,N_29807,N_29819);
nor UO_2601 (O_2601,N_29995,N_29871);
or UO_2602 (O_2602,N_29878,N_29980);
xnor UO_2603 (O_2603,N_29877,N_29948);
or UO_2604 (O_2604,N_29861,N_29831);
or UO_2605 (O_2605,N_29958,N_29927);
xor UO_2606 (O_2606,N_29977,N_29817);
xor UO_2607 (O_2607,N_29963,N_29801);
nand UO_2608 (O_2608,N_29870,N_29973);
nand UO_2609 (O_2609,N_29816,N_29958);
nand UO_2610 (O_2610,N_29905,N_29943);
or UO_2611 (O_2611,N_29954,N_29878);
nor UO_2612 (O_2612,N_29992,N_29914);
xor UO_2613 (O_2613,N_29945,N_29946);
nand UO_2614 (O_2614,N_29981,N_29828);
xnor UO_2615 (O_2615,N_29967,N_29869);
xnor UO_2616 (O_2616,N_29890,N_29861);
xor UO_2617 (O_2617,N_29946,N_29888);
nand UO_2618 (O_2618,N_29941,N_29988);
xnor UO_2619 (O_2619,N_29967,N_29903);
or UO_2620 (O_2620,N_29887,N_29934);
nor UO_2621 (O_2621,N_29935,N_29924);
and UO_2622 (O_2622,N_29991,N_29835);
and UO_2623 (O_2623,N_29810,N_29856);
nand UO_2624 (O_2624,N_29916,N_29951);
xor UO_2625 (O_2625,N_29845,N_29834);
xnor UO_2626 (O_2626,N_29948,N_29867);
nand UO_2627 (O_2627,N_29879,N_29974);
or UO_2628 (O_2628,N_29897,N_29822);
and UO_2629 (O_2629,N_29910,N_29945);
xnor UO_2630 (O_2630,N_29844,N_29803);
and UO_2631 (O_2631,N_29978,N_29817);
xnor UO_2632 (O_2632,N_29980,N_29921);
nand UO_2633 (O_2633,N_29891,N_29986);
nand UO_2634 (O_2634,N_29869,N_29894);
nand UO_2635 (O_2635,N_29817,N_29868);
nor UO_2636 (O_2636,N_29984,N_29969);
and UO_2637 (O_2637,N_29877,N_29884);
and UO_2638 (O_2638,N_29802,N_29808);
or UO_2639 (O_2639,N_29836,N_29965);
nand UO_2640 (O_2640,N_29946,N_29826);
xnor UO_2641 (O_2641,N_29977,N_29827);
xnor UO_2642 (O_2642,N_29840,N_29802);
nor UO_2643 (O_2643,N_29832,N_29966);
nand UO_2644 (O_2644,N_29937,N_29943);
nand UO_2645 (O_2645,N_29869,N_29863);
xnor UO_2646 (O_2646,N_29849,N_29830);
and UO_2647 (O_2647,N_29988,N_29865);
xor UO_2648 (O_2648,N_29852,N_29875);
nand UO_2649 (O_2649,N_29862,N_29935);
and UO_2650 (O_2650,N_29926,N_29999);
or UO_2651 (O_2651,N_29937,N_29824);
xor UO_2652 (O_2652,N_29836,N_29818);
nand UO_2653 (O_2653,N_29931,N_29962);
xor UO_2654 (O_2654,N_29800,N_29946);
or UO_2655 (O_2655,N_29860,N_29891);
xor UO_2656 (O_2656,N_29841,N_29944);
or UO_2657 (O_2657,N_29907,N_29804);
xor UO_2658 (O_2658,N_29838,N_29958);
nor UO_2659 (O_2659,N_29801,N_29934);
and UO_2660 (O_2660,N_29996,N_29869);
or UO_2661 (O_2661,N_29864,N_29823);
and UO_2662 (O_2662,N_29872,N_29955);
nand UO_2663 (O_2663,N_29851,N_29868);
xnor UO_2664 (O_2664,N_29936,N_29968);
or UO_2665 (O_2665,N_29801,N_29820);
nand UO_2666 (O_2666,N_29865,N_29999);
nor UO_2667 (O_2667,N_29806,N_29905);
xnor UO_2668 (O_2668,N_29886,N_29980);
xnor UO_2669 (O_2669,N_29811,N_29980);
nor UO_2670 (O_2670,N_29810,N_29815);
or UO_2671 (O_2671,N_29834,N_29824);
xnor UO_2672 (O_2672,N_29972,N_29831);
or UO_2673 (O_2673,N_29862,N_29929);
nand UO_2674 (O_2674,N_29889,N_29921);
or UO_2675 (O_2675,N_29835,N_29999);
xnor UO_2676 (O_2676,N_29871,N_29807);
or UO_2677 (O_2677,N_29914,N_29999);
xnor UO_2678 (O_2678,N_29889,N_29942);
or UO_2679 (O_2679,N_29867,N_29887);
or UO_2680 (O_2680,N_29828,N_29863);
xor UO_2681 (O_2681,N_29808,N_29844);
or UO_2682 (O_2682,N_29903,N_29983);
and UO_2683 (O_2683,N_29903,N_29863);
xor UO_2684 (O_2684,N_29830,N_29939);
nand UO_2685 (O_2685,N_29996,N_29866);
nor UO_2686 (O_2686,N_29948,N_29890);
nor UO_2687 (O_2687,N_29815,N_29845);
xnor UO_2688 (O_2688,N_29843,N_29942);
or UO_2689 (O_2689,N_29861,N_29844);
and UO_2690 (O_2690,N_29837,N_29930);
or UO_2691 (O_2691,N_29966,N_29866);
xor UO_2692 (O_2692,N_29888,N_29955);
nand UO_2693 (O_2693,N_29965,N_29998);
xor UO_2694 (O_2694,N_29977,N_29969);
xor UO_2695 (O_2695,N_29964,N_29988);
nor UO_2696 (O_2696,N_29805,N_29920);
and UO_2697 (O_2697,N_29950,N_29837);
or UO_2698 (O_2698,N_29839,N_29852);
xor UO_2699 (O_2699,N_29873,N_29996);
nand UO_2700 (O_2700,N_29860,N_29807);
nand UO_2701 (O_2701,N_29996,N_29832);
nor UO_2702 (O_2702,N_29826,N_29815);
xor UO_2703 (O_2703,N_29890,N_29908);
or UO_2704 (O_2704,N_29852,N_29898);
nor UO_2705 (O_2705,N_29904,N_29924);
nand UO_2706 (O_2706,N_29973,N_29828);
nor UO_2707 (O_2707,N_29935,N_29891);
nor UO_2708 (O_2708,N_29939,N_29888);
xnor UO_2709 (O_2709,N_29885,N_29870);
nor UO_2710 (O_2710,N_29968,N_29834);
nor UO_2711 (O_2711,N_29849,N_29887);
nor UO_2712 (O_2712,N_29913,N_29830);
nand UO_2713 (O_2713,N_29848,N_29844);
and UO_2714 (O_2714,N_29851,N_29903);
or UO_2715 (O_2715,N_29924,N_29874);
and UO_2716 (O_2716,N_29915,N_29987);
and UO_2717 (O_2717,N_29998,N_29970);
xnor UO_2718 (O_2718,N_29997,N_29957);
xor UO_2719 (O_2719,N_29984,N_29941);
or UO_2720 (O_2720,N_29913,N_29877);
nand UO_2721 (O_2721,N_29847,N_29819);
or UO_2722 (O_2722,N_29962,N_29888);
and UO_2723 (O_2723,N_29844,N_29964);
xnor UO_2724 (O_2724,N_29976,N_29875);
nand UO_2725 (O_2725,N_29899,N_29907);
or UO_2726 (O_2726,N_29829,N_29952);
or UO_2727 (O_2727,N_29944,N_29964);
or UO_2728 (O_2728,N_29965,N_29947);
nand UO_2729 (O_2729,N_29811,N_29957);
and UO_2730 (O_2730,N_29888,N_29973);
nor UO_2731 (O_2731,N_29966,N_29936);
nand UO_2732 (O_2732,N_29994,N_29948);
nand UO_2733 (O_2733,N_29887,N_29860);
and UO_2734 (O_2734,N_29956,N_29861);
or UO_2735 (O_2735,N_29999,N_29981);
nand UO_2736 (O_2736,N_29819,N_29996);
nor UO_2737 (O_2737,N_29871,N_29848);
nor UO_2738 (O_2738,N_29880,N_29962);
and UO_2739 (O_2739,N_29922,N_29904);
xor UO_2740 (O_2740,N_29820,N_29839);
nor UO_2741 (O_2741,N_29882,N_29919);
and UO_2742 (O_2742,N_29869,N_29971);
nor UO_2743 (O_2743,N_29948,N_29950);
and UO_2744 (O_2744,N_29819,N_29848);
nor UO_2745 (O_2745,N_29821,N_29981);
and UO_2746 (O_2746,N_29922,N_29897);
nor UO_2747 (O_2747,N_29826,N_29857);
or UO_2748 (O_2748,N_29841,N_29836);
and UO_2749 (O_2749,N_29984,N_29844);
nand UO_2750 (O_2750,N_29993,N_29963);
nand UO_2751 (O_2751,N_29854,N_29825);
nand UO_2752 (O_2752,N_29887,N_29994);
nor UO_2753 (O_2753,N_29803,N_29938);
or UO_2754 (O_2754,N_29913,N_29932);
and UO_2755 (O_2755,N_29815,N_29835);
and UO_2756 (O_2756,N_29909,N_29937);
nand UO_2757 (O_2757,N_29829,N_29859);
xor UO_2758 (O_2758,N_29918,N_29973);
nor UO_2759 (O_2759,N_29943,N_29914);
xor UO_2760 (O_2760,N_29969,N_29890);
or UO_2761 (O_2761,N_29906,N_29884);
and UO_2762 (O_2762,N_29880,N_29968);
nand UO_2763 (O_2763,N_29912,N_29945);
or UO_2764 (O_2764,N_29837,N_29984);
or UO_2765 (O_2765,N_29879,N_29977);
and UO_2766 (O_2766,N_29921,N_29898);
or UO_2767 (O_2767,N_29868,N_29888);
or UO_2768 (O_2768,N_29987,N_29812);
nor UO_2769 (O_2769,N_29868,N_29856);
nand UO_2770 (O_2770,N_29973,N_29841);
or UO_2771 (O_2771,N_29918,N_29956);
nor UO_2772 (O_2772,N_29809,N_29853);
nor UO_2773 (O_2773,N_29830,N_29935);
and UO_2774 (O_2774,N_29996,N_29999);
or UO_2775 (O_2775,N_29934,N_29949);
nor UO_2776 (O_2776,N_29925,N_29823);
xor UO_2777 (O_2777,N_29907,N_29930);
or UO_2778 (O_2778,N_29814,N_29842);
xor UO_2779 (O_2779,N_29954,N_29859);
nor UO_2780 (O_2780,N_29856,N_29965);
nand UO_2781 (O_2781,N_29953,N_29940);
or UO_2782 (O_2782,N_29802,N_29804);
and UO_2783 (O_2783,N_29886,N_29982);
xor UO_2784 (O_2784,N_29942,N_29974);
nand UO_2785 (O_2785,N_29810,N_29954);
or UO_2786 (O_2786,N_29859,N_29974);
and UO_2787 (O_2787,N_29948,N_29861);
xnor UO_2788 (O_2788,N_29977,N_29932);
xnor UO_2789 (O_2789,N_29965,N_29870);
nand UO_2790 (O_2790,N_29851,N_29943);
nand UO_2791 (O_2791,N_29964,N_29850);
or UO_2792 (O_2792,N_29851,N_29821);
nand UO_2793 (O_2793,N_29953,N_29901);
nand UO_2794 (O_2794,N_29853,N_29847);
nand UO_2795 (O_2795,N_29824,N_29813);
xor UO_2796 (O_2796,N_29853,N_29965);
and UO_2797 (O_2797,N_29917,N_29985);
nor UO_2798 (O_2798,N_29898,N_29966);
xnor UO_2799 (O_2799,N_29930,N_29903);
nor UO_2800 (O_2800,N_29963,N_29957);
nand UO_2801 (O_2801,N_29953,N_29907);
nand UO_2802 (O_2802,N_29901,N_29909);
xnor UO_2803 (O_2803,N_29908,N_29970);
nand UO_2804 (O_2804,N_29804,N_29895);
nand UO_2805 (O_2805,N_29946,N_29921);
nor UO_2806 (O_2806,N_29823,N_29953);
or UO_2807 (O_2807,N_29906,N_29867);
and UO_2808 (O_2808,N_29933,N_29893);
nor UO_2809 (O_2809,N_29864,N_29881);
and UO_2810 (O_2810,N_29945,N_29813);
nor UO_2811 (O_2811,N_29989,N_29827);
and UO_2812 (O_2812,N_29872,N_29838);
xor UO_2813 (O_2813,N_29995,N_29817);
nor UO_2814 (O_2814,N_29850,N_29841);
and UO_2815 (O_2815,N_29845,N_29925);
nor UO_2816 (O_2816,N_29865,N_29824);
nand UO_2817 (O_2817,N_29956,N_29820);
nand UO_2818 (O_2818,N_29846,N_29849);
nand UO_2819 (O_2819,N_29835,N_29894);
and UO_2820 (O_2820,N_29922,N_29902);
xor UO_2821 (O_2821,N_29912,N_29863);
nand UO_2822 (O_2822,N_29999,N_29909);
nor UO_2823 (O_2823,N_29803,N_29914);
nor UO_2824 (O_2824,N_29843,N_29972);
nor UO_2825 (O_2825,N_29832,N_29872);
nand UO_2826 (O_2826,N_29985,N_29872);
nor UO_2827 (O_2827,N_29896,N_29871);
nor UO_2828 (O_2828,N_29965,N_29811);
xnor UO_2829 (O_2829,N_29866,N_29879);
and UO_2830 (O_2830,N_29983,N_29814);
nor UO_2831 (O_2831,N_29810,N_29899);
nand UO_2832 (O_2832,N_29998,N_29981);
or UO_2833 (O_2833,N_29808,N_29814);
nand UO_2834 (O_2834,N_29893,N_29925);
nor UO_2835 (O_2835,N_29937,N_29941);
xor UO_2836 (O_2836,N_29904,N_29882);
or UO_2837 (O_2837,N_29924,N_29833);
xnor UO_2838 (O_2838,N_29917,N_29849);
nand UO_2839 (O_2839,N_29874,N_29865);
and UO_2840 (O_2840,N_29877,N_29881);
or UO_2841 (O_2841,N_29899,N_29985);
and UO_2842 (O_2842,N_29942,N_29927);
nor UO_2843 (O_2843,N_29824,N_29947);
nand UO_2844 (O_2844,N_29892,N_29923);
xor UO_2845 (O_2845,N_29841,N_29862);
and UO_2846 (O_2846,N_29854,N_29804);
or UO_2847 (O_2847,N_29966,N_29858);
and UO_2848 (O_2848,N_29866,N_29907);
or UO_2849 (O_2849,N_29810,N_29990);
and UO_2850 (O_2850,N_29913,N_29801);
nand UO_2851 (O_2851,N_29960,N_29917);
nand UO_2852 (O_2852,N_29917,N_29943);
or UO_2853 (O_2853,N_29886,N_29968);
or UO_2854 (O_2854,N_29886,N_29877);
xor UO_2855 (O_2855,N_29939,N_29876);
or UO_2856 (O_2856,N_29861,N_29824);
or UO_2857 (O_2857,N_29931,N_29963);
and UO_2858 (O_2858,N_29973,N_29881);
nor UO_2859 (O_2859,N_29974,N_29986);
and UO_2860 (O_2860,N_29898,N_29960);
nand UO_2861 (O_2861,N_29815,N_29998);
nand UO_2862 (O_2862,N_29850,N_29949);
or UO_2863 (O_2863,N_29825,N_29844);
xor UO_2864 (O_2864,N_29816,N_29832);
xnor UO_2865 (O_2865,N_29900,N_29832);
or UO_2866 (O_2866,N_29895,N_29879);
or UO_2867 (O_2867,N_29958,N_29975);
or UO_2868 (O_2868,N_29889,N_29999);
or UO_2869 (O_2869,N_29903,N_29917);
nand UO_2870 (O_2870,N_29982,N_29825);
nand UO_2871 (O_2871,N_29920,N_29873);
or UO_2872 (O_2872,N_29810,N_29964);
xnor UO_2873 (O_2873,N_29919,N_29902);
and UO_2874 (O_2874,N_29948,N_29859);
nand UO_2875 (O_2875,N_29868,N_29828);
xnor UO_2876 (O_2876,N_29872,N_29982);
xor UO_2877 (O_2877,N_29921,N_29866);
nand UO_2878 (O_2878,N_29999,N_29982);
and UO_2879 (O_2879,N_29929,N_29992);
nor UO_2880 (O_2880,N_29869,N_29938);
nor UO_2881 (O_2881,N_29872,N_29975);
nand UO_2882 (O_2882,N_29957,N_29852);
xnor UO_2883 (O_2883,N_29939,N_29917);
nor UO_2884 (O_2884,N_29908,N_29942);
xnor UO_2885 (O_2885,N_29837,N_29944);
or UO_2886 (O_2886,N_29987,N_29944);
and UO_2887 (O_2887,N_29891,N_29872);
nor UO_2888 (O_2888,N_29860,N_29930);
and UO_2889 (O_2889,N_29911,N_29920);
nor UO_2890 (O_2890,N_29955,N_29801);
and UO_2891 (O_2891,N_29989,N_29829);
nor UO_2892 (O_2892,N_29947,N_29992);
and UO_2893 (O_2893,N_29903,N_29926);
nand UO_2894 (O_2894,N_29807,N_29822);
xnor UO_2895 (O_2895,N_29925,N_29827);
nand UO_2896 (O_2896,N_29953,N_29854);
nor UO_2897 (O_2897,N_29812,N_29808);
nand UO_2898 (O_2898,N_29995,N_29934);
xnor UO_2899 (O_2899,N_29906,N_29977);
xnor UO_2900 (O_2900,N_29834,N_29835);
nor UO_2901 (O_2901,N_29835,N_29848);
and UO_2902 (O_2902,N_29999,N_29899);
or UO_2903 (O_2903,N_29868,N_29860);
or UO_2904 (O_2904,N_29941,N_29954);
and UO_2905 (O_2905,N_29927,N_29837);
or UO_2906 (O_2906,N_29911,N_29962);
or UO_2907 (O_2907,N_29923,N_29821);
nand UO_2908 (O_2908,N_29912,N_29983);
xnor UO_2909 (O_2909,N_29987,N_29885);
and UO_2910 (O_2910,N_29837,N_29824);
or UO_2911 (O_2911,N_29909,N_29970);
xor UO_2912 (O_2912,N_29878,N_29972);
nor UO_2913 (O_2913,N_29847,N_29883);
and UO_2914 (O_2914,N_29828,N_29849);
and UO_2915 (O_2915,N_29845,N_29966);
xor UO_2916 (O_2916,N_29911,N_29836);
or UO_2917 (O_2917,N_29920,N_29858);
and UO_2918 (O_2918,N_29968,N_29939);
nor UO_2919 (O_2919,N_29832,N_29987);
and UO_2920 (O_2920,N_29971,N_29905);
xnor UO_2921 (O_2921,N_29906,N_29928);
xor UO_2922 (O_2922,N_29920,N_29809);
nand UO_2923 (O_2923,N_29845,N_29905);
nand UO_2924 (O_2924,N_29851,N_29940);
nor UO_2925 (O_2925,N_29985,N_29860);
nor UO_2926 (O_2926,N_29916,N_29934);
or UO_2927 (O_2927,N_29867,N_29851);
nor UO_2928 (O_2928,N_29854,N_29883);
xor UO_2929 (O_2929,N_29910,N_29824);
and UO_2930 (O_2930,N_29924,N_29896);
nand UO_2931 (O_2931,N_29879,N_29912);
and UO_2932 (O_2932,N_29924,N_29829);
and UO_2933 (O_2933,N_29850,N_29867);
and UO_2934 (O_2934,N_29969,N_29863);
nor UO_2935 (O_2935,N_29864,N_29837);
or UO_2936 (O_2936,N_29810,N_29936);
or UO_2937 (O_2937,N_29892,N_29895);
xor UO_2938 (O_2938,N_29869,N_29903);
nor UO_2939 (O_2939,N_29819,N_29808);
xnor UO_2940 (O_2940,N_29894,N_29926);
or UO_2941 (O_2941,N_29806,N_29991);
xnor UO_2942 (O_2942,N_29833,N_29962);
xnor UO_2943 (O_2943,N_29919,N_29982);
and UO_2944 (O_2944,N_29806,N_29842);
or UO_2945 (O_2945,N_29886,N_29988);
xor UO_2946 (O_2946,N_29805,N_29816);
nand UO_2947 (O_2947,N_29827,N_29931);
nor UO_2948 (O_2948,N_29943,N_29831);
xor UO_2949 (O_2949,N_29918,N_29826);
nor UO_2950 (O_2950,N_29956,N_29962);
or UO_2951 (O_2951,N_29843,N_29839);
nand UO_2952 (O_2952,N_29836,N_29944);
nor UO_2953 (O_2953,N_29873,N_29921);
xor UO_2954 (O_2954,N_29802,N_29816);
nor UO_2955 (O_2955,N_29863,N_29955);
nor UO_2956 (O_2956,N_29892,N_29910);
and UO_2957 (O_2957,N_29977,N_29938);
or UO_2958 (O_2958,N_29949,N_29856);
xor UO_2959 (O_2959,N_29803,N_29912);
or UO_2960 (O_2960,N_29828,N_29890);
or UO_2961 (O_2961,N_29863,N_29838);
and UO_2962 (O_2962,N_29883,N_29809);
and UO_2963 (O_2963,N_29984,N_29873);
nand UO_2964 (O_2964,N_29918,N_29835);
or UO_2965 (O_2965,N_29891,N_29950);
or UO_2966 (O_2966,N_29826,N_29956);
nor UO_2967 (O_2967,N_29883,N_29866);
xor UO_2968 (O_2968,N_29944,N_29994);
xor UO_2969 (O_2969,N_29983,N_29849);
nor UO_2970 (O_2970,N_29849,N_29836);
xnor UO_2971 (O_2971,N_29803,N_29974);
nor UO_2972 (O_2972,N_29895,N_29831);
xnor UO_2973 (O_2973,N_29954,N_29884);
nand UO_2974 (O_2974,N_29842,N_29858);
or UO_2975 (O_2975,N_29948,N_29805);
nor UO_2976 (O_2976,N_29911,N_29863);
and UO_2977 (O_2977,N_29975,N_29816);
or UO_2978 (O_2978,N_29920,N_29947);
nand UO_2979 (O_2979,N_29945,N_29878);
nor UO_2980 (O_2980,N_29994,N_29853);
xor UO_2981 (O_2981,N_29997,N_29866);
or UO_2982 (O_2982,N_29959,N_29819);
nand UO_2983 (O_2983,N_29895,N_29940);
nand UO_2984 (O_2984,N_29854,N_29844);
and UO_2985 (O_2985,N_29881,N_29807);
nor UO_2986 (O_2986,N_29937,N_29931);
and UO_2987 (O_2987,N_29865,N_29848);
or UO_2988 (O_2988,N_29966,N_29987);
nor UO_2989 (O_2989,N_29922,N_29921);
and UO_2990 (O_2990,N_29992,N_29846);
xnor UO_2991 (O_2991,N_29813,N_29936);
or UO_2992 (O_2992,N_29842,N_29811);
and UO_2993 (O_2993,N_29940,N_29942);
xor UO_2994 (O_2994,N_29805,N_29813);
nand UO_2995 (O_2995,N_29837,N_29917);
xnor UO_2996 (O_2996,N_29895,N_29920);
or UO_2997 (O_2997,N_29943,N_29883);
or UO_2998 (O_2998,N_29929,N_29829);
nand UO_2999 (O_2999,N_29945,N_29876);
nand UO_3000 (O_3000,N_29934,N_29997);
xor UO_3001 (O_3001,N_29838,N_29816);
nand UO_3002 (O_3002,N_29893,N_29856);
and UO_3003 (O_3003,N_29965,N_29955);
or UO_3004 (O_3004,N_29990,N_29895);
nor UO_3005 (O_3005,N_29975,N_29915);
or UO_3006 (O_3006,N_29882,N_29854);
nand UO_3007 (O_3007,N_29845,N_29999);
xnor UO_3008 (O_3008,N_29919,N_29888);
nor UO_3009 (O_3009,N_29925,N_29910);
xor UO_3010 (O_3010,N_29975,N_29848);
nand UO_3011 (O_3011,N_29896,N_29804);
or UO_3012 (O_3012,N_29900,N_29825);
and UO_3013 (O_3013,N_29879,N_29857);
nor UO_3014 (O_3014,N_29997,N_29858);
nor UO_3015 (O_3015,N_29852,N_29890);
nand UO_3016 (O_3016,N_29888,N_29935);
and UO_3017 (O_3017,N_29807,N_29916);
nand UO_3018 (O_3018,N_29890,N_29926);
xor UO_3019 (O_3019,N_29985,N_29885);
xnor UO_3020 (O_3020,N_29909,N_29805);
xor UO_3021 (O_3021,N_29893,N_29906);
and UO_3022 (O_3022,N_29825,N_29826);
xor UO_3023 (O_3023,N_29984,N_29922);
xnor UO_3024 (O_3024,N_29856,N_29843);
xor UO_3025 (O_3025,N_29881,N_29936);
or UO_3026 (O_3026,N_29940,N_29877);
xnor UO_3027 (O_3027,N_29878,N_29800);
nand UO_3028 (O_3028,N_29910,N_29821);
nor UO_3029 (O_3029,N_29800,N_29864);
or UO_3030 (O_3030,N_29898,N_29975);
and UO_3031 (O_3031,N_29895,N_29869);
nor UO_3032 (O_3032,N_29961,N_29979);
or UO_3033 (O_3033,N_29818,N_29922);
xor UO_3034 (O_3034,N_29806,N_29829);
or UO_3035 (O_3035,N_29893,N_29831);
and UO_3036 (O_3036,N_29927,N_29847);
xor UO_3037 (O_3037,N_29852,N_29888);
nor UO_3038 (O_3038,N_29911,N_29985);
nand UO_3039 (O_3039,N_29881,N_29834);
xor UO_3040 (O_3040,N_29859,N_29951);
xnor UO_3041 (O_3041,N_29991,N_29892);
or UO_3042 (O_3042,N_29802,N_29874);
or UO_3043 (O_3043,N_29853,N_29964);
nand UO_3044 (O_3044,N_29914,N_29851);
or UO_3045 (O_3045,N_29828,N_29946);
or UO_3046 (O_3046,N_29805,N_29966);
and UO_3047 (O_3047,N_29979,N_29832);
or UO_3048 (O_3048,N_29903,N_29890);
nor UO_3049 (O_3049,N_29852,N_29864);
or UO_3050 (O_3050,N_29801,N_29961);
nand UO_3051 (O_3051,N_29959,N_29947);
nand UO_3052 (O_3052,N_29989,N_29877);
and UO_3053 (O_3053,N_29988,N_29913);
nand UO_3054 (O_3054,N_29807,N_29872);
nor UO_3055 (O_3055,N_29867,N_29823);
xnor UO_3056 (O_3056,N_29976,N_29956);
or UO_3057 (O_3057,N_29966,N_29836);
or UO_3058 (O_3058,N_29847,N_29924);
nor UO_3059 (O_3059,N_29927,N_29843);
nor UO_3060 (O_3060,N_29924,N_29811);
and UO_3061 (O_3061,N_29950,N_29926);
nand UO_3062 (O_3062,N_29901,N_29857);
xnor UO_3063 (O_3063,N_29859,N_29980);
xor UO_3064 (O_3064,N_29828,N_29891);
or UO_3065 (O_3065,N_29978,N_29860);
or UO_3066 (O_3066,N_29811,N_29964);
xor UO_3067 (O_3067,N_29992,N_29967);
nand UO_3068 (O_3068,N_29805,N_29818);
nand UO_3069 (O_3069,N_29966,N_29844);
xor UO_3070 (O_3070,N_29936,N_29866);
or UO_3071 (O_3071,N_29956,N_29953);
or UO_3072 (O_3072,N_29835,N_29960);
nor UO_3073 (O_3073,N_29881,N_29962);
nor UO_3074 (O_3074,N_29868,N_29837);
or UO_3075 (O_3075,N_29888,N_29916);
nand UO_3076 (O_3076,N_29850,N_29868);
nor UO_3077 (O_3077,N_29960,N_29843);
xor UO_3078 (O_3078,N_29820,N_29960);
and UO_3079 (O_3079,N_29916,N_29988);
or UO_3080 (O_3080,N_29899,N_29967);
xnor UO_3081 (O_3081,N_29888,N_29861);
or UO_3082 (O_3082,N_29971,N_29871);
and UO_3083 (O_3083,N_29958,N_29902);
nand UO_3084 (O_3084,N_29807,N_29830);
nand UO_3085 (O_3085,N_29905,N_29897);
and UO_3086 (O_3086,N_29988,N_29872);
or UO_3087 (O_3087,N_29874,N_29848);
nand UO_3088 (O_3088,N_29987,N_29939);
or UO_3089 (O_3089,N_29970,N_29949);
xnor UO_3090 (O_3090,N_29819,N_29916);
nand UO_3091 (O_3091,N_29984,N_29949);
nand UO_3092 (O_3092,N_29999,N_29850);
nand UO_3093 (O_3093,N_29853,N_29913);
nor UO_3094 (O_3094,N_29948,N_29810);
xnor UO_3095 (O_3095,N_29950,N_29909);
and UO_3096 (O_3096,N_29994,N_29979);
xnor UO_3097 (O_3097,N_29907,N_29843);
nor UO_3098 (O_3098,N_29847,N_29807);
xnor UO_3099 (O_3099,N_29896,N_29892);
nand UO_3100 (O_3100,N_29963,N_29890);
nand UO_3101 (O_3101,N_29906,N_29944);
and UO_3102 (O_3102,N_29994,N_29832);
xor UO_3103 (O_3103,N_29852,N_29926);
xor UO_3104 (O_3104,N_29896,N_29972);
xor UO_3105 (O_3105,N_29964,N_29846);
nor UO_3106 (O_3106,N_29866,N_29933);
or UO_3107 (O_3107,N_29831,N_29953);
nor UO_3108 (O_3108,N_29839,N_29950);
nand UO_3109 (O_3109,N_29940,N_29863);
xor UO_3110 (O_3110,N_29986,N_29885);
or UO_3111 (O_3111,N_29889,N_29954);
nand UO_3112 (O_3112,N_29886,N_29826);
xnor UO_3113 (O_3113,N_29801,N_29978);
or UO_3114 (O_3114,N_29838,N_29915);
nor UO_3115 (O_3115,N_29838,N_29934);
nor UO_3116 (O_3116,N_29835,N_29992);
nand UO_3117 (O_3117,N_29950,N_29916);
nor UO_3118 (O_3118,N_29992,N_29810);
nor UO_3119 (O_3119,N_29865,N_29939);
or UO_3120 (O_3120,N_29943,N_29962);
or UO_3121 (O_3121,N_29895,N_29981);
xnor UO_3122 (O_3122,N_29857,N_29980);
nand UO_3123 (O_3123,N_29863,N_29848);
nor UO_3124 (O_3124,N_29937,N_29910);
and UO_3125 (O_3125,N_29953,N_29934);
nand UO_3126 (O_3126,N_29952,N_29840);
nand UO_3127 (O_3127,N_29843,N_29956);
nor UO_3128 (O_3128,N_29815,N_29989);
and UO_3129 (O_3129,N_29984,N_29882);
xnor UO_3130 (O_3130,N_29833,N_29979);
and UO_3131 (O_3131,N_29853,N_29813);
nor UO_3132 (O_3132,N_29954,N_29894);
xor UO_3133 (O_3133,N_29884,N_29927);
nor UO_3134 (O_3134,N_29873,N_29842);
nor UO_3135 (O_3135,N_29931,N_29859);
nor UO_3136 (O_3136,N_29917,N_29949);
and UO_3137 (O_3137,N_29960,N_29808);
or UO_3138 (O_3138,N_29857,N_29889);
nor UO_3139 (O_3139,N_29925,N_29849);
and UO_3140 (O_3140,N_29820,N_29806);
nand UO_3141 (O_3141,N_29967,N_29974);
xnor UO_3142 (O_3142,N_29947,N_29896);
and UO_3143 (O_3143,N_29965,N_29802);
nor UO_3144 (O_3144,N_29810,N_29827);
nor UO_3145 (O_3145,N_29868,N_29946);
xor UO_3146 (O_3146,N_29944,N_29957);
xnor UO_3147 (O_3147,N_29849,N_29897);
and UO_3148 (O_3148,N_29933,N_29882);
nand UO_3149 (O_3149,N_29807,N_29926);
nor UO_3150 (O_3150,N_29902,N_29890);
nand UO_3151 (O_3151,N_29953,N_29886);
or UO_3152 (O_3152,N_29882,N_29969);
nor UO_3153 (O_3153,N_29806,N_29899);
xor UO_3154 (O_3154,N_29821,N_29965);
and UO_3155 (O_3155,N_29902,N_29809);
xnor UO_3156 (O_3156,N_29926,N_29901);
nor UO_3157 (O_3157,N_29930,N_29805);
and UO_3158 (O_3158,N_29918,N_29849);
and UO_3159 (O_3159,N_29947,N_29971);
and UO_3160 (O_3160,N_29916,N_29810);
or UO_3161 (O_3161,N_29995,N_29974);
nand UO_3162 (O_3162,N_29881,N_29865);
or UO_3163 (O_3163,N_29821,N_29838);
xor UO_3164 (O_3164,N_29802,N_29830);
or UO_3165 (O_3165,N_29804,N_29883);
nand UO_3166 (O_3166,N_29989,N_29935);
nor UO_3167 (O_3167,N_29869,N_29988);
and UO_3168 (O_3168,N_29861,N_29901);
nor UO_3169 (O_3169,N_29802,N_29926);
or UO_3170 (O_3170,N_29909,N_29911);
and UO_3171 (O_3171,N_29869,N_29890);
nor UO_3172 (O_3172,N_29826,N_29914);
or UO_3173 (O_3173,N_29827,N_29874);
nand UO_3174 (O_3174,N_29814,N_29875);
nor UO_3175 (O_3175,N_29802,N_29850);
xnor UO_3176 (O_3176,N_29812,N_29921);
nand UO_3177 (O_3177,N_29912,N_29806);
and UO_3178 (O_3178,N_29909,N_29836);
xnor UO_3179 (O_3179,N_29999,N_29922);
or UO_3180 (O_3180,N_29881,N_29984);
nor UO_3181 (O_3181,N_29863,N_29894);
xor UO_3182 (O_3182,N_29806,N_29955);
nand UO_3183 (O_3183,N_29881,N_29989);
or UO_3184 (O_3184,N_29804,N_29973);
xor UO_3185 (O_3185,N_29838,N_29802);
and UO_3186 (O_3186,N_29935,N_29837);
nand UO_3187 (O_3187,N_29963,N_29974);
or UO_3188 (O_3188,N_29854,N_29879);
and UO_3189 (O_3189,N_29929,N_29831);
nand UO_3190 (O_3190,N_29892,N_29830);
or UO_3191 (O_3191,N_29907,N_29942);
or UO_3192 (O_3192,N_29992,N_29829);
nor UO_3193 (O_3193,N_29878,N_29866);
xnor UO_3194 (O_3194,N_29998,N_29877);
or UO_3195 (O_3195,N_29908,N_29883);
nand UO_3196 (O_3196,N_29849,N_29941);
nand UO_3197 (O_3197,N_29824,N_29961);
xor UO_3198 (O_3198,N_29957,N_29844);
and UO_3199 (O_3199,N_29837,N_29816);
and UO_3200 (O_3200,N_29937,N_29844);
nand UO_3201 (O_3201,N_29846,N_29841);
nand UO_3202 (O_3202,N_29875,N_29951);
xor UO_3203 (O_3203,N_29904,N_29872);
nand UO_3204 (O_3204,N_29953,N_29859);
nor UO_3205 (O_3205,N_29997,N_29908);
or UO_3206 (O_3206,N_29877,N_29805);
nor UO_3207 (O_3207,N_29856,N_29906);
nand UO_3208 (O_3208,N_29951,N_29940);
nor UO_3209 (O_3209,N_29918,N_29999);
nand UO_3210 (O_3210,N_29922,N_29816);
or UO_3211 (O_3211,N_29883,N_29826);
or UO_3212 (O_3212,N_29982,N_29951);
or UO_3213 (O_3213,N_29821,N_29948);
nand UO_3214 (O_3214,N_29933,N_29829);
or UO_3215 (O_3215,N_29975,N_29972);
nor UO_3216 (O_3216,N_29995,N_29904);
xnor UO_3217 (O_3217,N_29882,N_29914);
xnor UO_3218 (O_3218,N_29980,N_29914);
xor UO_3219 (O_3219,N_29899,N_29923);
xor UO_3220 (O_3220,N_29866,N_29985);
or UO_3221 (O_3221,N_29965,N_29805);
nor UO_3222 (O_3222,N_29811,N_29938);
xor UO_3223 (O_3223,N_29861,N_29892);
and UO_3224 (O_3224,N_29937,N_29994);
or UO_3225 (O_3225,N_29822,N_29944);
or UO_3226 (O_3226,N_29993,N_29959);
or UO_3227 (O_3227,N_29814,N_29826);
nand UO_3228 (O_3228,N_29971,N_29873);
nor UO_3229 (O_3229,N_29892,N_29815);
and UO_3230 (O_3230,N_29853,N_29953);
and UO_3231 (O_3231,N_29946,N_29832);
and UO_3232 (O_3232,N_29944,N_29833);
nand UO_3233 (O_3233,N_29864,N_29993);
nand UO_3234 (O_3234,N_29901,N_29966);
and UO_3235 (O_3235,N_29884,N_29870);
xor UO_3236 (O_3236,N_29807,N_29902);
nand UO_3237 (O_3237,N_29845,N_29871);
or UO_3238 (O_3238,N_29851,N_29999);
and UO_3239 (O_3239,N_29946,N_29983);
nand UO_3240 (O_3240,N_29805,N_29859);
nand UO_3241 (O_3241,N_29894,N_29864);
nand UO_3242 (O_3242,N_29884,N_29837);
nor UO_3243 (O_3243,N_29819,N_29953);
or UO_3244 (O_3244,N_29901,N_29828);
nor UO_3245 (O_3245,N_29864,N_29829);
and UO_3246 (O_3246,N_29908,N_29805);
nor UO_3247 (O_3247,N_29996,N_29811);
or UO_3248 (O_3248,N_29827,N_29928);
xor UO_3249 (O_3249,N_29998,N_29977);
nor UO_3250 (O_3250,N_29839,N_29882);
xor UO_3251 (O_3251,N_29953,N_29945);
nand UO_3252 (O_3252,N_29866,N_29981);
and UO_3253 (O_3253,N_29865,N_29953);
xor UO_3254 (O_3254,N_29843,N_29913);
and UO_3255 (O_3255,N_29875,N_29844);
nor UO_3256 (O_3256,N_29891,N_29985);
nor UO_3257 (O_3257,N_29954,N_29870);
xor UO_3258 (O_3258,N_29871,N_29846);
or UO_3259 (O_3259,N_29857,N_29855);
nor UO_3260 (O_3260,N_29861,N_29908);
or UO_3261 (O_3261,N_29925,N_29864);
nand UO_3262 (O_3262,N_29922,N_29804);
nand UO_3263 (O_3263,N_29990,N_29826);
xor UO_3264 (O_3264,N_29826,N_29929);
nor UO_3265 (O_3265,N_29958,N_29846);
xor UO_3266 (O_3266,N_29874,N_29838);
and UO_3267 (O_3267,N_29912,N_29875);
or UO_3268 (O_3268,N_29927,N_29959);
and UO_3269 (O_3269,N_29891,N_29944);
nor UO_3270 (O_3270,N_29909,N_29964);
nor UO_3271 (O_3271,N_29853,N_29905);
nor UO_3272 (O_3272,N_29887,N_29889);
and UO_3273 (O_3273,N_29874,N_29851);
xor UO_3274 (O_3274,N_29904,N_29913);
nor UO_3275 (O_3275,N_29894,N_29875);
or UO_3276 (O_3276,N_29804,N_29892);
xnor UO_3277 (O_3277,N_29839,N_29951);
nand UO_3278 (O_3278,N_29862,N_29818);
xnor UO_3279 (O_3279,N_29949,N_29807);
nand UO_3280 (O_3280,N_29945,N_29951);
or UO_3281 (O_3281,N_29867,N_29982);
or UO_3282 (O_3282,N_29810,N_29938);
nor UO_3283 (O_3283,N_29866,N_29836);
nand UO_3284 (O_3284,N_29947,N_29873);
and UO_3285 (O_3285,N_29845,N_29979);
nor UO_3286 (O_3286,N_29937,N_29809);
and UO_3287 (O_3287,N_29890,N_29833);
and UO_3288 (O_3288,N_29819,N_29805);
xor UO_3289 (O_3289,N_29973,N_29898);
nor UO_3290 (O_3290,N_29846,N_29906);
and UO_3291 (O_3291,N_29877,N_29946);
and UO_3292 (O_3292,N_29890,N_29856);
xnor UO_3293 (O_3293,N_29853,N_29919);
nand UO_3294 (O_3294,N_29808,N_29951);
xnor UO_3295 (O_3295,N_29870,N_29983);
xor UO_3296 (O_3296,N_29985,N_29887);
nand UO_3297 (O_3297,N_29985,N_29883);
or UO_3298 (O_3298,N_29884,N_29882);
nand UO_3299 (O_3299,N_29825,N_29846);
nor UO_3300 (O_3300,N_29983,N_29947);
and UO_3301 (O_3301,N_29992,N_29957);
nor UO_3302 (O_3302,N_29875,N_29829);
or UO_3303 (O_3303,N_29861,N_29985);
xor UO_3304 (O_3304,N_29902,N_29956);
and UO_3305 (O_3305,N_29838,N_29920);
or UO_3306 (O_3306,N_29912,N_29881);
or UO_3307 (O_3307,N_29925,N_29914);
nor UO_3308 (O_3308,N_29873,N_29862);
nand UO_3309 (O_3309,N_29943,N_29820);
or UO_3310 (O_3310,N_29843,N_29867);
nand UO_3311 (O_3311,N_29931,N_29819);
nor UO_3312 (O_3312,N_29871,N_29979);
or UO_3313 (O_3313,N_29998,N_29864);
nand UO_3314 (O_3314,N_29857,N_29802);
nor UO_3315 (O_3315,N_29839,N_29806);
or UO_3316 (O_3316,N_29880,N_29914);
nor UO_3317 (O_3317,N_29882,N_29965);
or UO_3318 (O_3318,N_29957,N_29818);
or UO_3319 (O_3319,N_29818,N_29819);
or UO_3320 (O_3320,N_29816,N_29884);
xnor UO_3321 (O_3321,N_29856,N_29864);
nor UO_3322 (O_3322,N_29802,N_29902);
or UO_3323 (O_3323,N_29805,N_29958);
and UO_3324 (O_3324,N_29895,N_29918);
nand UO_3325 (O_3325,N_29930,N_29991);
nor UO_3326 (O_3326,N_29979,N_29878);
xor UO_3327 (O_3327,N_29955,N_29919);
or UO_3328 (O_3328,N_29801,N_29958);
or UO_3329 (O_3329,N_29911,N_29817);
and UO_3330 (O_3330,N_29992,N_29861);
or UO_3331 (O_3331,N_29977,N_29907);
nor UO_3332 (O_3332,N_29952,N_29885);
xor UO_3333 (O_3333,N_29805,N_29949);
nand UO_3334 (O_3334,N_29904,N_29842);
nor UO_3335 (O_3335,N_29906,N_29934);
nor UO_3336 (O_3336,N_29977,N_29946);
and UO_3337 (O_3337,N_29901,N_29934);
nor UO_3338 (O_3338,N_29859,N_29828);
and UO_3339 (O_3339,N_29886,N_29881);
and UO_3340 (O_3340,N_29987,N_29868);
nor UO_3341 (O_3341,N_29874,N_29844);
or UO_3342 (O_3342,N_29935,N_29859);
or UO_3343 (O_3343,N_29934,N_29836);
nor UO_3344 (O_3344,N_29957,N_29919);
nor UO_3345 (O_3345,N_29885,N_29854);
nand UO_3346 (O_3346,N_29855,N_29900);
and UO_3347 (O_3347,N_29868,N_29918);
and UO_3348 (O_3348,N_29951,N_29831);
nand UO_3349 (O_3349,N_29909,N_29868);
or UO_3350 (O_3350,N_29929,N_29988);
xnor UO_3351 (O_3351,N_29814,N_29942);
xor UO_3352 (O_3352,N_29970,N_29988);
nor UO_3353 (O_3353,N_29942,N_29865);
and UO_3354 (O_3354,N_29922,N_29865);
xnor UO_3355 (O_3355,N_29861,N_29936);
xnor UO_3356 (O_3356,N_29803,N_29936);
nand UO_3357 (O_3357,N_29994,N_29837);
or UO_3358 (O_3358,N_29863,N_29811);
and UO_3359 (O_3359,N_29813,N_29948);
xnor UO_3360 (O_3360,N_29936,N_29933);
nand UO_3361 (O_3361,N_29836,N_29846);
nor UO_3362 (O_3362,N_29990,N_29892);
nand UO_3363 (O_3363,N_29808,N_29906);
or UO_3364 (O_3364,N_29839,N_29993);
and UO_3365 (O_3365,N_29895,N_29837);
and UO_3366 (O_3366,N_29984,N_29836);
nor UO_3367 (O_3367,N_29971,N_29959);
or UO_3368 (O_3368,N_29921,N_29909);
xnor UO_3369 (O_3369,N_29990,N_29877);
nand UO_3370 (O_3370,N_29831,N_29925);
nand UO_3371 (O_3371,N_29855,N_29926);
nor UO_3372 (O_3372,N_29958,N_29925);
or UO_3373 (O_3373,N_29931,N_29813);
nor UO_3374 (O_3374,N_29953,N_29847);
or UO_3375 (O_3375,N_29892,N_29869);
xor UO_3376 (O_3376,N_29918,N_29808);
xor UO_3377 (O_3377,N_29914,N_29938);
nand UO_3378 (O_3378,N_29910,N_29981);
xor UO_3379 (O_3379,N_29941,N_29836);
nand UO_3380 (O_3380,N_29841,N_29949);
nand UO_3381 (O_3381,N_29891,N_29833);
or UO_3382 (O_3382,N_29811,N_29928);
and UO_3383 (O_3383,N_29980,N_29801);
or UO_3384 (O_3384,N_29802,N_29862);
and UO_3385 (O_3385,N_29801,N_29887);
nor UO_3386 (O_3386,N_29922,N_29923);
nand UO_3387 (O_3387,N_29875,N_29984);
xor UO_3388 (O_3388,N_29898,N_29813);
nor UO_3389 (O_3389,N_29932,N_29873);
nor UO_3390 (O_3390,N_29902,N_29939);
nand UO_3391 (O_3391,N_29804,N_29899);
nand UO_3392 (O_3392,N_29925,N_29991);
nand UO_3393 (O_3393,N_29898,N_29861);
or UO_3394 (O_3394,N_29849,N_29987);
nor UO_3395 (O_3395,N_29888,N_29848);
and UO_3396 (O_3396,N_29863,N_29939);
and UO_3397 (O_3397,N_29969,N_29836);
and UO_3398 (O_3398,N_29885,N_29853);
xor UO_3399 (O_3399,N_29958,N_29869);
and UO_3400 (O_3400,N_29958,N_29984);
or UO_3401 (O_3401,N_29840,N_29926);
nand UO_3402 (O_3402,N_29805,N_29810);
and UO_3403 (O_3403,N_29968,N_29990);
nand UO_3404 (O_3404,N_29858,N_29903);
nand UO_3405 (O_3405,N_29916,N_29905);
or UO_3406 (O_3406,N_29802,N_29858);
xnor UO_3407 (O_3407,N_29932,N_29911);
nor UO_3408 (O_3408,N_29829,N_29976);
nand UO_3409 (O_3409,N_29883,N_29802);
and UO_3410 (O_3410,N_29847,N_29948);
xor UO_3411 (O_3411,N_29821,N_29892);
nand UO_3412 (O_3412,N_29900,N_29833);
nand UO_3413 (O_3413,N_29832,N_29825);
nor UO_3414 (O_3414,N_29841,N_29902);
or UO_3415 (O_3415,N_29965,N_29875);
xnor UO_3416 (O_3416,N_29983,N_29863);
nand UO_3417 (O_3417,N_29867,N_29853);
or UO_3418 (O_3418,N_29801,N_29964);
and UO_3419 (O_3419,N_29892,N_29956);
or UO_3420 (O_3420,N_29861,N_29912);
or UO_3421 (O_3421,N_29945,N_29897);
or UO_3422 (O_3422,N_29807,N_29991);
nor UO_3423 (O_3423,N_29889,N_29801);
or UO_3424 (O_3424,N_29912,N_29976);
xnor UO_3425 (O_3425,N_29937,N_29919);
nor UO_3426 (O_3426,N_29877,N_29970);
nand UO_3427 (O_3427,N_29901,N_29967);
or UO_3428 (O_3428,N_29895,N_29922);
nor UO_3429 (O_3429,N_29952,N_29891);
nand UO_3430 (O_3430,N_29939,N_29966);
xnor UO_3431 (O_3431,N_29848,N_29847);
xor UO_3432 (O_3432,N_29823,N_29840);
xnor UO_3433 (O_3433,N_29890,N_29802);
xor UO_3434 (O_3434,N_29819,N_29905);
and UO_3435 (O_3435,N_29969,N_29966);
xnor UO_3436 (O_3436,N_29958,N_29951);
nand UO_3437 (O_3437,N_29878,N_29818);
nor UO_3438 (O_3438,N_29809,N_29826);
nor UO_3439 (O_3439,N_29900,N_29957);
and UO_3440 (O_3440,N_29983,N_29894);
xnor UO_3441 (O_3441,N_29873,N_29836);
nor UO_3442 (O_3442,N_29997,N_29825);
xnor UO_3443 (O_3443,N_29841,N_29998);
nand UO_3444 (O_3444,N_29867,N_29952);
and UO_3445 (O_3445,N_29951,N_29897);
and UO_3446 (O_3446,N_29856,N_29970);
xnor UO_3447 (O_3447,N_29907,N_29955);
and UO_3448 (O_3448,N_29889,N_29814);
and UO_3449 (O_3449,N_29911,N_29839);
or UO_3450 (O_3450,N_29900,N_29828);
nor UO_3451 (O_3451,N_29833,N_29998);
nand UO_3452 (O_3452,N_29984,N_29859);
and UO_3453 (O_3453,N_29814,N_29888);
or UO_3454 (O_3454,N_29966,N_29827);
or UO_3455 (O_3455,N_29902,N_29871);
or UO_3456 (O_3456,N_29870,N_29835);
or UO_3457 (O_3457,N_29938,N_29872);
nand UO_3458 (O_3458,N_29983,N_29853);
nor UO_3459 (O_3459,N_29888,N_29889);
nand UO_3460 (O_3460,N_29825,N_29856);
nand UO_3461 (O_3461,N_29979,N_29804);
and UO_3462 (O_3462,N_29928,N_29858);
nand UO_3463 (O_3463,N_29990,N_29900);
nor UO_3464 (O_3464,N_29998,N_29989);
nor UO_3465 (O_3465,N_29820,N_29805);
or UO_3466 (O_3466,N_29869,N_29918);
xnor UO_3467 (O_3467,N_29816,N_29989);
or UO_3468 (O_3468,N_29931,N_29806);
and UO_3469 (O_3469,N_29958,N_29833);
nor UO_3470 (O_3470,N_29952,N_29846);
or UO_3471 (O_3471,N_29864,N_29866);
xor UO_3472 (O_3472,N_29822,N_29888);
or UO_3473 (O_3473,N_29856,N_29888);
nor UO_3474 (O_3474,N_29995,N_29896);
nand UO_3475 (O_3475,N_29850,N_29902);
and UO_3476 (O_3476,N_29945,N_29999);
xor UO_3477 (O_3477,N_29800,N_29951);
nor UO_3478 (O_3478,N_29818,N_29801);
or UO_3479 (O_3479,N_29810,N_29914);
xnor UO_3480 (O_3480,N_29928,N_29865);
and UO_3481 (O_3481,N_29959,N_29870);
xor UO_3482 (O_3482,N_29922,N_29893);
nor UO_3483 (O_3483,N_29886,N_29855);
xnor UO_3484 (O_3484,N_29817,N_29864);
nand UO_3485 (O_3485,N_29873,N_29931);
and UO_3486 (O_3486,N_29899,N_29926);
nand UO_3487 (O_3487,N_29965,N_29937);
and UO_3488 (O_3488,N_29894,N_29944);
xnor UO_3489 (O_3489,N_29848,N_29969);
or UO_3490 (O_3490,N_29819,N_29946);
nand UO_3491 (O_3491,N_29994,N_29934);
xnor UO_3492 (O_3492,N_29974,N_29916);
nand UO_3493 (O_3493,N_29958,N_29963);
or UO_3494 (O_3494,N_29975,N_29917);
or UO_3495 (O_3495,N_29977,N_29955);
nand UO_3496 (O_3496,N_29871,N_29868);
nand UO_3497 (O_3497,N_29881,N_29838);
or UO_3498 (O_3498,N_29990,N_29908);
xor UO_3499 (O_3499,N_29910,N_29858);
endmodule