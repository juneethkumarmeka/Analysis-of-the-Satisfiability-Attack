module basic_1500_15000_2000_10_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_297,In_1009);
and U1 (N_1,In_460,In_14);
nor U2 (N_2,In_794,In_18);
nand U3 (N_3,In_286,In_23);
nor U4 (N_4,In_731,In_912);
nand U5 (N_5,In_84,In_696);
nand U6 (N_6,In_643,In_1247);
nand U7 (N_7,In_1464,In_152);
nor U8 (N_8,In_228,In_1208);
and U9 (N_9,In_87,In_24);
nor U10 (N_10,In_3,In_1287);
nand U11 (N_11,In_1115,In_32);
xor U12 (N_12,In_1405,In_19);
and U13 (N_13,In_311,In_1063);
nand U14 (N_14,In_190,In_498);
nor U15 (N_15,In_887,In_1141);
nor U16 (N_16,In_560,In_1304);
and U17 (N_17,In_43,In_7);
xor U18 (N_18,In_544,In_1463);
nand U19 (N_19,In_1457,In_475);
nand U20 (N_20,In_334,In_295);
and U21 (N_21,In_419,In_770);
nor U22 (N_22,In_568,In_871);
nand U23 (N_23,In_403,In_1467);
nor U24 (N_24,In_1184,In_1205);
nor U25 (N_25,In_216,In_741);
and U26 (N_26,In_1368,In_446);
nand U27 (N_27,In_955,In_478);
and U28 (N_28,In_561,In_1163);
or U29 (N_29,In_550,In_719);
or U30 (N_30,In_1165,In_1278);
or U31 (N_31,In_652,In_1377);
nor U32 (N_32,In_786,In_232);
nor U33 (N_33,In_1474,In_125);
nor U34 (N_34,In_844,In_1284);
or U35 (N_35,In_407,In_66);
nor U36 (N_36,In_171,In_793);
or U37 (N_37,In_114,In_1495);
nor U38 (N_38,In_848,In_1309);
nand U39 (N_39,In_957,In_335);
and U40 (N_40,In_679,In_1466);
and U41 (N_41,In_875,In_1478);
nand U42 (N_42,In_624,In_722);
nand U43 (N_43,In_733,In_527);
nor U44 (N_44,In_950,In_395);
nor U45 (N_45,In_942,In_1359);
nand U46 (N_46,In_867,In_674);
and U47 (N_47,In_422,In_1370);
or U48 (N_48,In_1088,In_281);
nor U49 (N_49,In_1401,In_933);
xor U50 (N_50,In_149,In_1151);
or U51 (N_51,In_103,In_52);
xor U52 (N_52,In_646,In_1119);
and U53 (N_53,In_943,In_655);
nand U54 (N_54,In_264,In_1122);
and U55 (N_55,In_1067,In_850);
or U56 (N_56,In_807,In_501);
xnor U57 (N_57,In_657,In_362);
and U58 (N_58,In_805,In_1048);
nand U59 (N_59,In_296,In_1186);
nor U60 (N_60,In_869,In_1485);
nand U61 (N_61,In_1499,In_1159);
and U62 (N_62,In_810,In_1385);
or U63 (N_63,In_927,In_278);
or U64 (N_64,In_914,In_504);
nand U65 (N_65,In_174,In_1130);
nor U66 (N_66,In_67,In_481);
or U67 (N_67,In_440,In_1396);
and U68 (N_68,In_255,In_874);
nand U69 (N_69,In_1496,In_1053);
nor U70 (N_70,In_393,In_95);
nand U71 (N_71,In_203,In_354);
nand U72 (N_72,In_75,In_99);
or U73 (N_73,In_359,In_737);
nor U74 (N_74,In_1353,In_378);
nand U75 (N_75,In_136,In_1337);
or U76 (N_76,In_329,In_1367);
xor U77 (N_77,In_890,In_345);
and U78 (N_78,In_179,In_252);
and U79 (N_79,In_298,In_828);
or U80 (N_80,In_779,In_1104);
nand U81 (N_81,In_505,In_797);
nand U82 (N_82,In_1095,In_396);
and U83 (N_83,In_1065,In_1289);
and U84 (N_84,In_206,In_186);
and U85 (N_85,In_804,In_249);
nand U86 (N_86,In_109,In_305);
or U87 (N_87,In_1218,In_146);
and U88 (N_88,In_928,In_932);
and U89 (N_89,In_865,In_938);
nand U90 (N_90,In_840,In_1308);
nand U91 (N_91,In_668,In_1384);
and U92 (N_92,In_65,In_1021);
nor U93 (N_93,In_1280,In_1275);
nor U94 (N_94,In_925,In_832);
nor U95 (N_95,In_1259,In_158);
nor U96 (N_96,In_113,In_1258);
or U97 (N_97,In_257,In_1213);
nand U98 (N_98,In_1041,In_852);
nand U99 (N_99,In_870,In_219);
or U100 (N_100,In_1271,In_433);
nor U101 (N_101,In_1288,In_740);
or U102 (N_102,In_897,In_1164);
nor U103 (N_103,In_1200,In_1197);
and U104 (N_104,In_616,In_953);
xnor U105 (N_105,In_511,In_8);
nand U106 (N_106,In_1383,In_626);
nor U107 (N_107,In_439,In_833);
and U108 (N_108,In_1248,In_682);
nand U109 (N_109,In_96,In_473);
or U110 (N_110,In_566,In_165);
and U111 (N_111,In_1492,In_1029);
nand U112 (N_112,In_525,In_1406);
or U113 (N_113,In_1303,In_303);
or U114 (N_114,In_792,In_1030);
and U115 (N_115,In_201,In_892);
or U116 (N_116,In_226,In_670);
xnor U117 (N_117,In_1068,In_1253);
or U118 (N_118,In_61,In_1292);
or U119 (N_119,In_160,In_391);
nand U120 (N_120,In_313,In_1486);
or U121 (N_121,In_796,In_1042);
xor U122 (N_122,In_1071,In_428);
nor U123 (N_123,In_614,In_1223);
and U124 (N_124,In_126,In_776);
or U125 (N_125,In_649,In_635);
or U126 (N_126,In_751,In_542);
nor U127 (N_127,In_367,In_1416);
or U128 (N_128,In_1187,In_1059);
xnor U129 (N_129,In_1290,In_1402);
or U130 (N_130,In_1108,In_110);
nor U131 (N_131,In_1376,In_1142);
nor U132 (N_132,In_548,In_1243);
nand U133 (N_133,In_464,In_389);
or U134 (N_134,In_1459,In_1144);
and U135 (N_135,In_347,In_929);
nand U136 (N_136,In_51,In_157);
or U137 (N_137,In_268,In_651);
xor U138 (N_138,In_233,In_767);
nor U139 (N_139,In_429,In_918);
nor U140 (N_140,In_1056,In_284);
nor U141 (N_141,In_491,In_181);
nor U142 (N_142,In_220,In_1375);
or U143 (N_143,In_762,In_137);
or U144 (N_144,In_1132,In_312);
nand U145 (N_145,In_130,In_16);
and U146 (N_146,In_1234,In_374);
nand U147 (N_147,In_808,In_769);
nor U148 (N_148,In_1023,In_860);
nor U149 (N_149,In_60,In_813);
nand U150 (N_150,In_325,In_1039);
and U151 (N_151,In_846,In_836);
xnor U152 (N_152,In_331,In_1311);
or U153 (N_153,In_894,In_678);
or U154 (N_154,In_58,In_1414);
and U155 (N_155,In_547,In_431);
and U156 (N_156,In_1343,In_1211);
nor U157 (N_157,In_739,In_975);
and U158 (N_158,In_405,In_915);
nor U159 (N_159,In_798,In_764);
nor U160 (N_160,In_1236,In_91);
nor U161 (N_161,In_386,In_726);
and U162 (N_162,In_666,In_585);
nand U163 (N_163,In_1319,In_1279);
xor U164 (N_164,In_490,In_586);
and U165 (N_165,In_1484,In_885);
xor U166 (N_166,In_178,In_17);
and U167 (N_167,In_127,In_237);
nand U168 (N_168,In_1404,In_36);
and U169 (N_169,In_350,In_549);
nand U170 (N_170,In_310,In_992);
or U171 (N_171,In_1116,In_1323);
nor U172 (N_172,In_115,In_111);
nand U173 (N_173,In_366,In_71);
nor U174 (N_174,In_1450,In_673);
nor U175 (N_175,In_1462,In_77);
nor U176 (N_176,In_57,In_990);
and U177 (N_177,In_148,In_30);
and U178 (N_178,In_1036,In_292);
and U179 (N_179,In_514,In_876);
or U180 (N_180,In_97,In_1326);
or U181 (N_181,In_754,In_935);
nor U182 (N_182,In_177,In_699);
or U183 (N_183,In_261,In_664);
nor U184 (N_184,In_214,In_820);
and U185 (N_185,In_629,In_708);
and U186 (N_186,In_289,In_841);
or U187 (N_187,In_135,In_1183);
nor U188 (N_188,In_200,In_1155);
nor U189 (N_189,In_94,In_517);
or U190 (N_190,In_1101,In_720);
and U191 (N_191,In_946,In_905);
or U192 (N_192,In_1334,In_742);
xnor U193 (N_193,In_316,In_1246);
and U194 (N_194,In_0,In_326);
or U195 (N_195,In_1300,In_818);
xnor U196 (N_196,In_1096,In_904);
nand U197 (N_197,In_1113,In_202);
or U198 (N_198,In_1228,In_623);
xnor U199 (N_199,In_477,In_659);
nor U200 (N_200,In_732,In_1427);
or U201 (N_201,In_138,In_1476);
or U202 (N_202,In_50,In_901);
xor U203 (N_203,In_22,In_599);
nor U204 (N_204,In_82,In_132);
and U205 (N_205,In_1410,In_1245);
and U206 (N_206,In_829,In_817);
nand U207 (N_207,In_315,In_610);
and U208 (N_208,In_958,In_1381);
or U209 (N_209,In_1294,In_107);
nand U210 (N_210,In_1254,In_1328);
and U211 (N_211,In_633,In_27);
and U212 (N_212,In_520,In_1480);
and U213 (N_213,In_1324,In_499);
or U214 (N_214,In_883,In_410);
and U215 (N_215,In_479,In_360);
nand U216 (N_216,In_815,In_744);
and U217 (N_217,In_920,In_1097);
xor U218 (N_218,In_620,In_1120);
nor U219 (N_219,In_265,In_377);
nor U220 (N_220,In_385,In_1192);
nand U221 (N_221,In_523,In_748);
nor U222 (N_222,In_1188,In_824);
nand U223 (N_223,In_400,In_1161);
or U224 (N_224,In_645,In_642);
nand U225 (N_225,In_618,In_986);
and U226 (N_226,In_1051,In_902);
xnor U227 (N_227,In_38,In_516);
nor U228 (N_228,In_13,In_809);
or U229 (N_229,In_746,In_859);
or U230 (N_230,In_729,In_1090);
nand U231 (N_231,In_736,In_1412);
nor U232 (N_232,In_1318,In_830);
or U233 (N_233,In_591,In_583);
nand U234 (N_234,In_1317,In_1293);
nor U235 (N_235,In_145,In_691);
nand U236 (N_236,In_1106,In_1100);
or U237 (N_237,In_1085,In_1157);
xnor U238 (N_238,In_1389,In_789);
and U239 (N_239,In_1014,In_1491);
and U240 (N_240,In_924,In_254);
nor U241 (N_241,In_880,In_529);
nor U242 (N_242,In_323,In_1267);
or U243 (N_243,In_761,In_217);
or U244 (N_244,In_1475,In_680);
or U245 (N_245,In_543,In_967);
and U246 (N_246,In_37,In_535);
nor U247 (N_247,In_1212,In_166);
nand U248 (N_248,In_294,In_1227);
nand U249 (N_249,In_1229,In_1215);
nor U250 (N_250,In_1235,In_944);
or U251 (N_251,In_1173,In_35);
nor U252 (N_252,In_1291,In_161);
xnor U253 (N_253,In_879,In_1007);
nor U254 (N_254,In_572,In_994);
nand U255 (N_255,In_811,In_392);
and U256 (N_256,In_884,In_1452);
xor U257 (N_257,In_845,In_697);
nand U258 (N_258,In_1449,In_688);
or U259 (N_259,In_106,In_379);
nand U260 (N_260,In_101,In_44);
and U261 (N_261,In_907,In_351);
and U262 (N_262,In_939,In_1341);
and U263 (N_263,In_675,In_1241);
nor U264 (N_264,In_959,In_483);
and U265 (N_265,In_877,In_898);
or U266 (N_266,In_416,In_1268);
or U267 (N_267,In_1182,In_319);
nand U268 (N_268,In_1369,In_1340);
and U269 (N_269,In_459,In_600);
or U270 (N_270,In_253,In_401);
xnor U271 (N_271,In_105,In_622);
and U272 (N_272,In_187,In_556);
or U273 (N_273,In_1072,In_337);
nor U274 (N_274,In_12,In_1336);
nand U275 (N_275,In_1066,In_1176);
and U276 (N_276,In_1430,In_74);
nand U277 (N_277,In_215,In_128);
and U278 (N_278,In_1004,In_795);
xnor U279 (N_279,In_172,In_262);
or U280 (N_280,In_1454,In_1167);
or U281 (N_281,In_133,In_300);
xnor U282 (N_282,In_54,In_948);
nand U283 (N_283,In_1320,In_438);
nand U284 (N_284,In_271,In_248);
and U285 (N_285,In_1202,In_25);
nand U286 (N_286,In_234,In_225);
or U287 (N_287,In_162,In_1128);
nand U288 (N_288,In_1017,In_458);
or U289 (N_289,In_1198,In_1307);
nor U290 (N_290,In_601,In_540);
and U291 (N_291,In_508,In_1458);
nor U292 (N_292,In_408,In_1332);
and U293 (N_293,In_49,In_63);
nand U294 (N_294,In_686,In_1087);
nor U295 (N_295,In_308,In_246);
or U296 (N_296,In_369,In_839);
nand U297 (N_297,In_1082,In_1361);
and U298 (N_298,In_453,In_814);
xor U299 (N_299,In_383,In_198);
nor U300 (N_300,In_590,In_1049);
or U301 (N_301,In_1135,In_1084);
nor U302 (N_302,In_412,In_352);
or U303 (N_303,In_290,In_92);
or U304 (N_304,In_1424,In_1225);
or U305 (N_305,In_409,In_578);
nor U306 (N_306,In_580,In_983);
xnor U307 (N_307,In_628,In_671);
and U308 (N_308,In_218,In_978);
or U309 (N_309,In_1070,In_1360);
nor U310 (N_310,In_661,In_1026);
and U311 (N_311,In_906,In_900);
or U312 (N_312,In_33,In_449);
or U313 (N_313,In_280,In_1121);
xor U314 (N_314,In_102,In_608);
xor U315 (N_315,In_538,In_317);
nor U316 (N_316,In_812,In_1362);
and U317 (N_317,In_765,In_421);
nand U318 (N_318,In_987,In_68);
nor U319 (N_319,In_539,In_42);
and U320 (N_320,In_1020,In_124);
nor U321 (N_321,In_1455,In_1002);
nor U322 (N_322,In_1170,In_768);
nor U323 (N_323,In_1327,In_1177);
nor U324 (N_324,In_653,In_909);
nor U325 (N_325,In_903,In_1216);
xor U326 (N_326,In_1044,In_1180);
or U327 (N_327,In_169,In_480);
and U328 (N_328,In_1387,In_1315);
xnor U329 (N_329,In_328,In_1018);
nand U330 (N_330,In_1199,In_1147);
or U331 (N_331,In_1277,In_1005);
nor U332 (N_332,In_1411,In_1333);
nor U333 (N_333,In_940,In_1335);
nand U334 (N_334,In_90,In_753);
and U335 (N_335,In_507,In_258);
nor U336 (N_336,In_916,In_364);
nand U337 (N_337,In_562,In_864);
nor U338 (N_338,In_781,In_447);
nand U339 (N_339,In_727,In_175);
nor U340 (N_340,In_999,In_1055);
nand U341 (N_341,In_10,In_1482);
xor U342 (N_342,In_183,In_752);
nand U343 (N_343,In_1162,In_579);
or U344 (N_344,In_150,In_151);
and U345 (N_345,In_1440,In_384);
xor U346 (N_346,In_1103,In_207);
nand U347 (N_347,In_1125,In_1060);
or U348 (N_348,In_274,In_755);
xnor U349 (N_349,In_1078,In_1425);
xor U350 (N_350,In_123,In_573);
nor U351 (N_351,In_1388,In_1352);
and U352 (N_352,In_9,In_773);
nor U353 (N_353,In_1305,In_656);
nand U354 (N_354,In_921,In_698);
or U355 (N_355,In_427,In_108);
nor U356 (N_356,In_822,In_275);
nor U357 (N_357,In_725,In_260);
nand U358 (N_358,In_868,In_502);
nor U359 (N_359,In_1262,In_1407);
nand U360 (N_360,In_80,In_567);
nand U361 (N_361,In_1081,In_602);
xor U362 (N_362,In_293,In_782);
or U363 (N_363,In_79,In_1016);
and U364 (N_364,In_291,In_470);
or U365 (N_365,In_1062,In_436);
and U366 (N_366,In_182,In_154);
and U367 (N_367,In_684,In_155);
and U368 (N_368,In_1456,In_1477);
and U369 (N_369,In_783,In_163);
xor U370 (N_370,In_1110,In_1347);
nand U371 (N_371,In_716,In_521);
nand U372 (N_372,In_1260,In_1460);
nor U373 (N_373,In_861,In_518);
nand U374 (N_374,In_1083,In_59);
or U375 (N_375,In_760,In_1446);
xnor U376 (N_376,In_1421,In_277);
nor U377 (N_377,In_996,In_1179);
and U378 (N_378,In_1150,In_660);
and U379 (N_379,In_48,In_631);
nor U380 (N_380,In_411,In_714);
or U381 (N_381,In_320,In_306);
and U382 (N_382,In_596,In_1439);
nor U383 (N_383,In_64,In_546);
nor U384 (N_384,In_122,In_144);
and U385 (N_385,In_1222,In_509);
and U386 (N_386,In_692,In_1175);
or U387 (N_387,In_168,In_1057);
nor U388 (N_388,In_609,In_639);
and U389 (N_389,In_777,In_1312);
nand U390 (N_390,In_1330,In_1217);
xnor U391 (N_391,In_823,In_448);
nor U392 (N_392,In_39,In_1143);
nand U393 (N_393,In_526,In_488);
xor U394 (N_394,In_1261,In_891);
and U395 (N_395,In_474,In_1252);
or U396 (N_396,In_247,In_53);
or U397 (N_397,In_1392,In_1178);
or U398 (N_398,In_667,In_503);
and U399 (N_399,In_658,In_766);
nor U400 (N_400,In_1408,In_457);
nand U401 (N_401,In_778,In_1283);
nor U402 (N_402,In_531,In_1274);
and U403 (N_403,In_993,In_47);
xnor U404 (N_404,In_1047,In_1358);
or U405 (N_405,In_1089,In_309);
or U406 (N_406,In_279,In_513);
and U407 (N_407,In_250,In_98);
nor U408 (N_408,In_563,In_984);
nand U409 (N_409,In_1093,In_595);
or U410 (N_410,In_493,In_238);
and U411 (N_411,In_966,In_119);
nor U412 (N_412,In_486,In_1302);
nor U413 (N_413,In_73,In_299);
nor U414 (N_414,In_497,In_1210);
nand U415 (N_415,In_1498,In_1378);
and U416 (N_416,In_1298,In_571);
xor U417 (N_417,In_598,In_533);
nand U418 (N_418,In_46,In_689);
nor U419 (N_419,In_1465,In_1365);
nand U420 (N_420,In_28,In_1043);
xor U421 (N_421,In_156,In_1270);
xor U422 (N_422,In_711,In_785);
nor U423 (N_423,In_683,In_707);
and U424 (N_424,In_6,In_387);
nor U425 (N_425,In_34,In_1196);
or U426 (N_426,In_1429,In_842);
nand U427 (N_427,In_1420,In_1058);
nand U428 (N_428,In_1181,In_467);
nand U429 (N_429,In_519,In_569);
nand U430 (N_430,In_715,In_878);
nand U431 (N_431,In_534,In_758);
nor U432 (N_432,In_1437,In_1444);
or U433 (N_433,In_1203,In_873);
nor U434 (N_434,In_1117,In_1397);
nand U435 (N_435,In_330,In_1349);
or U436 (N_436,In_376,In_397);
xnor U437 (N_437,In_496,In_1092);
or U438 (N_438,In_788,In_441);
nor U439 (N_439,In_1154,In_704);
or U440 (N_440,In_952,In_338);
nor U441 (N_441,In_1189,In_1028);
nor U442 (N_442,In_973,In_1338);
and U443 (N_443,In_390,In_1138);
and U444 (N_444,In_1105,In_693);
xnor U445 (N_445,In_314,In_370);
nand U446 (N_446,In_372,In_1490);
xnor U447 (N_447,In_703,In_989);
or U448 (N_448,In_584,In_239);
nand U449 (N_449,In_922,In_327);
or U450 (N_450,In_834,In_545);
and U451 (N_451,In_1357,In_1479);
and U452 (N_452,In_554,In_5);
or U453 (N_453,In_500,In_476);
or U454 (N_454,In_418,In_694);
nor U455 (N_455,In_750,In_709);
nor U456 (N_456,In_734,In_1145);
nor U457 (N_457,In_321,In_965);
nand U458 (N_458,In_197,In_801);
or U459 (N_459,In_995,In_1069);
nor U460 (N_460,In_650,In_1201);
nor U461 (N_461,In_357,In_211);
or U462 (N_462,In_230,In_613);
nand U463 (N_463,In_961,In_343);
nand U464 (N_464,In_1011,In_1386);
nand U465 (N_465,In_1107,In_229);
nor U466 (N_466,In_1239,In_302);
nand U467 (N_467,In_1426,In_1226);
or U468 (N_468,In_581,In_1322);
and U469 (N_469,In_988,In_1140);
and U470 (N_470,In_1481,In_837);
xnor U471 (N_471,In_611,In_373);
nor U472 (N_472,In_241,In_1443);
nor U473 (N_473,In_721,In_997);
nor U474 (N_474,In_1191,In_129);
and U475 (N_475,In_341,In_324);
xor U476 (N_476,In_245,In_594);
nand U477 (N_477,In_283,In_461);
nand U478 (N_478,In_826,In_20);
and U479 (N_479,In_242,In_466);
and U480 (N_480,In_866,In_1314);
nor U481 (N_481,In_456,In_1149);
and U482 (N_482,In_167,In_1024);
nand U483 (N_483,In_700,In_1432);
nand U484 (N_484,In_936,In_388);
nand U485 (N_485,In_333,In_1372);
nand U486 (N_486,In_559,In_76);
nor U487 (N_487,In_799,In_1313);
or U488 (N_488,In_450,In_827);
or U489 (N_489,In_1255,In_1214);
xor U490 (N_490,In_1185,In_552);
or U491 (N_491,In_1109,In_862);
nand U492 (N_492,In_577,In_1356);
or U493 (N_493,In_1346,In_349);
nor U494 (N_494,In_749,In_1025);
and U495 (N_495,In_886,In_1310);
nand U496 (N_496,In_1301,In_1129);
nor U497 (N_497,In_194,In_318);
nand U498 (N_498,In_1127,In_849);
nand U499 (N_499,In_638,In_164);
or U500 (N_500,In_724,In_831);
or U501 (N_501,In_1472,In_872);
nand U502 (N_502,In_971,In_471);
nor U503 (N_503,In_597,In_1264);
nor U504 (N_504,In_224,In_951);
nand U505 (N_505,In_1395,In_485);
and U506 (N_506,In_821,In_816);
or U507 (N_507,In_1428,In_557);
nor U508 (N_508,In_147,In_941);
or U509 (N_509,In_348,In_882);
or U510 (N_510,In_1094,In_1249);
or U511 (N_511,In_487,In_1445);
nor U512 (N_512,In_1393,In_1399);
or U513 (N_513,In_863,In_506);
or U514 (N_514,In_512,In_236);
nand U515 (N_515,In_1281,In_1156);
and U516 (N_516,In_1469,In_1231);
or U517 (N_517,In_340,In_1015);
xor U518 (N_518,In_1204,In_1345);
and U519 (N_519,In_70,In_510);
nand U520 (N_520,In_256,In_888);
xor U521 (N_521,In_763,In_1342);
or U522 (N_522,In_1061,In_911);
nor U523 (N_523,In_747,In_399);
and U524 (N_524,In_919,In_717);
nor U525 (N_525,In_847,In_1403);
nor U526 (N_526,In_1035,In_435);
nand U527 (N_527,In_803,In_88);
xor U528 (N_528,In_430,In_1263);
or U529 (N_529,In_434,In_273);
and U530 (N_530,In_701,In_630);
nand U531 (N_531,In_1232,In_1046);
xor U532 (N_532,In_553,In_462);
or U533 (N_533,In_802,In_1297);
or U534 (N_534,In_1038,In_632);
or U535 (N_535,In_153,In_695);
or U536 (N_536,In_1012,In_931);
and U537 (N_537,In_235,In_677);
or U538 (N_538,In_210,In_825);
and U539 (N_539,In_143,In_1052);
or U540 (N_540,In_1073,In_322);
nand U541 (N_541,In_368,In_1098);
nand U542 (N_542,In_536,In_1398);
or U543 (N_543,In_979,In_593);
and U544 (N_544,In_117,In_575);
xnor U545 (N_545,In_468,In_784);
and U546 (N_546,In_1000,In_227);
nor U547 (N_547,In_881,In_1219);
nor U548 (N_548,In_1033,In_853);
and U549 (N_549,In_282,In_1137);
nand U550 (N_550,In_209,In_1240);
or U551 (N_551,In_445,In_1453);
and U552 (N_552,In_221,In_908);
and U553 (N_553,In_1409,In_1483);
xnor U554 (N_554,In_1224,In_647);
xor U555 (N_555,In_414,In_196);
nand U556 (N_556,In_41,In_1447);
or U557 (N_557,In_240,In_855);
xnor U558 (N_558,In_743,In_270);
nand U559 (N_559,In_31,In_1473);
nor U560 (N_560,In_1153,In_1497);
nand U561 (N_561,In_1001,In_492);
and U562 (N_562,In_259,In_991);
and U563 (N_563,In_1244,In_759);
nand U564 (N_564,In_665,In_1433);
nor U565 (N_565,In_1152,In_1400);
nor U566 (N_566,In_970,In_524);
or U567 (N_567,In_1086,In_1037);
xnor U568 (N_568,In_15,In_772);
nor U569 (N_569,In_1374,In_4);
or U570 (N_570,In_757,In_960);
or U571 (N_571,In_705,In_288);
and U572 (N_572,In_968,In_285);
and U573 (N_573,In_1350,In_1276);
nand U574 (N_574,In_851,In_204);
nor U575 (N_575,In_56,In_1139);
or U576 (N_576,In_565,In_454);
nand U577 (N_577,In_582,In_452);
nand U578 (N_578,In_1131,In_118);
or U579 (N_579,In_1050,In_1299);
nand U580 (N_580,In_1494,In_1134);
or U581 (N_581,In_712,In_587);
and U582 (N_582,In_1080,In_89);
or U583 (N_583,In_528,In_1451);
and U584 (N_584,In_1114,In_1471);
or U585 (N_585,In_1285,In_251);
and U586 (N_586,In_184,In_947);
xnor U587 (N_587,In_272,In_856);
or U588 (N_588,In_365,In_199);
xor U589 (N_589,In_62,In_465);
xor U590 (N_590,In_706,In_361);
or U591 (N_591,In_854,In_1436);
and U592 (N_592,In_615,In_787);
xor U593 (N_593,In_735,In_1112);
nand U594 (N_594,In_417,In_188);
nor U595 (N_595,In_1373,In_1079);
nor U596 (N_596,In_1256,In_1431);
and U597 (N_597,In_998,In_1064);
and U598 (N_598,In_899,In_1250);
and U599 (N_599,In_934,In_402);
nor U600 (N_600,In_1221,In_78);
nor U601 (N_601,In_923,In_304);
nand U602 (N_602,In_404,In_432);
nor U603 (N_603,In_672,In_603);
or U604 (N_604,In_205,In_1423);
or U605 (N_605,In_141,In_558);
nand U606 (N_606,In_969,In_926);
and U607 (N_607,In_85,In_1027);
xor U608 (N_608,In_243,In_1032);
nor U609 (N_609,In_104,In_344);
nand U610 (N_610,In_917,In_140);
and U611 (N_611,In_790,In_985);
nand U612 (N_612,In_681,In_1099);
and U613 (N_613,In_120,In_627);
and U614 (N_614,In_223,In_1054);
or U615 (N_615,In_1209,In_895);
nor U616 (N_616,In_116,In_606);
and U617 (N_617,In_482,In_26);
or U618 (N_618,In_604,In_956);
nand U619 (N_619,In_442,In_81);
nand U620 (N_620,In_974,In_1194);
or U621 (N_621,In_185,In_949);
or U622 (N_622,In_208,In_644);
or U623 (N_623,In_121,In_634);
and U624 (N_624,In_222,In_687);
nor U625 (N_625,In_267,In_592);
nand U626 (N_626,In_972,In_937);
and U627 (N_627,In_1448,In_1045);
and U628 (N_628,In_1331,In_588);
xor U629 (N_629,In_522,In_771);
nand U630 (N_630,In_738,In_195);
and U631 (N_631,In_662,In_469);
or U632 (N_632,In_637,In_685);
or U633 (N_633,In_358,In_718);
nor U634 (N_634,In_730,In_1379);
or U635 (N_635,In_495,In_702);
nor U636 (N_636,In_515,In_382);
or U637 (N_637,In_806,In_857);
or U638 (N_638,In_1380,In_858);
nand U639 (N_639,In_1074,In_1418);
and U640 (N_640,In_287,In_1329);
nor U641 (N_641,In_1273,In_193);
and U642 (N_642,In_1136,In_1371);
nand U643 (N_643,In_1206,In_1470);
nor U644 (N_644,In_530,In_1195);
nor U645 (N_645,In_1158,In_1111);
and U646 (N_646,In_1091,In_619);
and U647 (N_647,In_394,In_444);
and U648 (N_648,In_1415,In_641);
nand U649 (N_649,In_1230,In_1488);
nor U650 (N_650,In_1487,In_244);
nand U651 (N_651,In_1193,In_489);
nor U652 (N_652,In_72,In_1251);
nor U653 (N_653,In_1123,In_131);
or U654 (N_654,In_676,In_494);
and U655 (N_655,In_380,In_1171);
and U656 (N_656,In_11,In_756);
or U657 (N_657,In_1075,In_663);
nor U658 (N_658,In_45,In_589);
xor U659 (N_659,In_93,In_29);
and U660 (N_660,In_532,In_266);
and U661 (N_661,In_191,In_332);
and U662 (N_662,In_963,In_1172);
nand U663 (N_663,In_455,In_424);
or U664 (N_664,In_112,In_69);
nand U665 (N_665,In_1238,In_1006);
and U666 (N_666,In_774,In_1394);
nor U667 (N_667,In_1133,In_1417);
nor U668 (N_668,In_1422,In_893);
nand U669 (N_669,In_139,In_86);
or U670 (N_670,In_1242,In_1220);
xor U671 (N_671,In_723,In_40);
and U672 (N_672,In_896,In_1282);
nand U673 (N_673,In_170,In_100);
and U674 (N_674,In_1435,In_213);
nor U675 (N_675,In_1169,In_910);
and U676 (N_676,In_1355,In_1390);
nand U677 (N_677,In_964,In_371);
nor U678 (N_678,In_981,In_713);
and U679 (N_679,In_1442,In_1022);
and U680 (N_680,In_640,In_913);
or U681 (N_681,In_353,In_363);
and U682 (N_682,In_356,In_819);
nor U683 (N_683,In_21,In_1321);
or U684 (N_684,In_212,In_537);
nor U685 (N_685,In_1441,In_1102);
xor U686 (N_686,In_621,In_1339);
nor U687 (N_687,In_1031,In_1207);
or U688 (N_688,In_1,In_1166);
nor U689 (N_689,In_484,In_1348);
nor U690 (N_690,In_339,In_1272);
or U691 (N_691,In_1316,In_1366);
nor U692 (N_692,In_1419,In_1146);
and U693 (N_693,In_1019,In_55);
and U694 (N_694,In_1003,In_1382);
nor U695 (N_695,In_346,In_1160);
nor U696 (N_696,In_1010,In_301);
or U697 (N_697,In_1286,In_2);
nor U698 (N_698,In_617,In_745);
nand U699 (N_699,In_1351,In_415);
nand U700 (N_700,In_838,In_1148);
and U701 (N_701,In_189,In_463);
and U702 (N_702,In_1364,In_945);
nand U703 (N_703,In_1076,In_355);
or U704 (N_704,In_1190,In_982);
nor U705 (N_705,In_1391,In_1325);
and U706 (N_706,In_192,In_443);
or U707 (N_707,In_231,In_648);
nor U708 (N_708,In_1266,In_1126);
or U709 (N_709,In_977,In_843);
xor U710 (N_710,In_1168,In_269);
nand U711 (N_711,In_962,In_1077);
nor U712 (N_712,In_1008,In_800);
or U713 (N_713,In_690,In_1034);
xnor U714 (N_714,In_472,In_176);
or U715 (N_715,In_423,In_605);
or U716 (N_716,In_1013,In_1295);
nor U717 (N_717,In_1237,In_1461);
and U718 (N_718,In_551,In_980);
and U719 (N_719,In_425,In_1344);
and U720 (N_720,In_710,In_420);
nand U721 (N_721,In_83,In_954);
xor U722 (N_722,In_1434,In_654);
nand U723 (N_723,In_173,In_574);
and U724 (N_724,In_307,In_142);
and U725 (N_725,In_780,In_1269);
nand U726 (N_726,In_1468,In_342);
and U727 (N_727,In_791,In_636);
xor U728 (N_728,In_134,In_1040);
or U729 (N_729,In_775,In_1233);
nand U730 (N_730,In_612,In_1306);
and U731 (N_731,In_1493,In_541);
or U732 (N_732,In_1296,In_1118);
or U733 (N_733,In_1363,In_1489);
and U734 (N_734,In_1413,In_1354);
nor U735 (N_735,In_406,In_835);
and U736 (N_736,In_180,In_889);
nor U737 (N_737,In_576,In_375);
and U738 (N_738,In_1265,In_555);
or U739 (N_739,In_276,In_381);
or U740 (N_740,In_625,In_159);
or U741 (N_741,In_930,In_570);
or U742 (N_742,In_1124,In_564);
and U743 (N_743,In_426,In_728);
and U744 (N_744,In_1257,In_669);
nor U745 (N_745,In_336,In_607);
nand U746 (N_746,In_976,In_413);
nor U747 (N_747,In_1438,In_398);
or U748 (N_748,In_451,In_263);
nor U749 (N_749,In_1174,In_437);
and U750 (N_750,In_983,In_578);
nand U751 (N_751,In_392,In_826);
or U752 (N_752,In_1133,In_1292);
or U753 (N_753,In_1148,In_256);
or U754 (N_754,In_131,In_305);
or U755 (N_755,In_754,In_183);
xnor U756 (N_756,In_870,In_1366);
nand U757 (N_757,In_147,In_1306);
nand U758 (N_758,In_1223,In_1490);
nand U759 (N_759,In_1484,In_1138);
nor U760 (N_760,In_1491,In_345);
or U761 (N_761,In_800,In_1418);
or U762 (N_762,In_1416,In_59);
nand U763 (N_763,In_1321,In_212);
nand U764 (N_764,In_1496,In_1458);
and U765 (N_765,In_752,In_93);
and U766 (N_766,In_277,In_1307);
or U767 (N_767,In_651,In_276);
xor U768 (N_768,In_1278,In_468);
nor U769 (N_769,In_349,In_1294);
nor U770 (N_770,In_217,In_331);
or U771 (N_771,In_1293,In_1022);
nand U772 (N_772,In_1058,In_789);
nor U773 (N_773,In_1175,In_1313);
nand U774 (N_774,In_1193,In_269);
xnor U775 (N_775,In_947,In_973);
or U776 (N_776,In_210,In_1212);
nand U777 (N_777,In_630,In_1246);
and U778 (N_778,In_746,In_430);
nor U779 (N_779,In_1141,In_294);
or U780 (N_780,In_1458,In_1202);
xor U781 (N_781,In_1402,In_1308);
nand U782 (N_782,In_420,In_19);
nand U783 (N_783,In_871,In_634);
nor U784 (N_784,In_1402,In_1240);
and U785 (N_785,In_542,In_164);
nor U786 (N_786,In_1170,In_450);
or U787 (N_787,In_572,In_1167);
or U788 (N_788,In_9,In_1478);
nand U789 (N_789,In_902,In_185);
nor U790 (N_790,In_391,In_554);
nand U791 (N_791,In_214,In_46);
and U792 (N_792,In_884,In_16);
nor U793 (N_793,In_1041,In_212);
or U794 (N_794,In_1283,In_71);
nor U795 (N_795,In_768,In_155);
or U796 (N_796,In_1370,In_139);
and U797 (N_797,In_0,In_235);
and U798 (N_798,In_1122,In_840);
or U799 (N_799,In_1102,In_0);
nand U800 (N_800,In_671,In_1225);
and U801 (N_801,In_1288,In_234);
nand U802 (N_802,In_419,In_984);
and U803 (N_803,In_76,In_828);
nor U804 (N_804,In_83,In_339);
xnor U805 (N_805,In_348,In_1119);
nor U806 (N_806,In_1418,In_665);
nand U807 (N_807,In_635,In_911);
and U808 (N_808,In_690,In_679);
and U809 (N_809,In_1153,In_359);
or U810 (N_810,In_118,In_1251);
nand U811 (N_811,In_361,In_948);
xor U812 (N_812,In_538,In_1405);
nor U813 (N_813,In_792,In_1113);
and U814 (N_814,In_460,In_1084);
nand U815 (N_815,In_814,In_487);
nand U816 (N_816,In_1323,In_1400);
or U817 (N_817,In_1074,In_1359);
and U818 (N_818,In_53,In_486);
nor U819 (N_819,In_855,In_615);
nor U820 (N_820,In_775,In_1375);
or U821 (N_821,In_1267,In_687);
nor U822 (N_822,In_1079,In_1068);
nor U823 (N_823,In_332,In_987);
or U824 (N_824,In_966,In_1438);
nand U825 (N_825,In_558,In_125);
and U826 (N_826,In_1133,In_544);
xor U827 (N_827,In_1111,In_344);
nor U828 (N_828,In_117,In_927);
or U829 (N_829,In_1286,In_1460);
or U830 (N_830,In_1248,In_714);
nand U831 (N_831,In_238,In_1151);
xnor U832 (N_832,In_896,In_274);
nand U833 (N_833,In_755,In_69);
nand U834 (N_834,In_253,In_394);
nand U835 (N_835,In_821,In_304);
xnor U836 (N_836,In_1173,In_1220);
or U837 (N_837,In_1067,In_1263);
or U838 (N_838,In_1273,In_801);
nand U839 (N_839,In_971,In_853);
xnor U840 (N_840,In_144,In_242);
or U841 (N_841,In_657,In_1062);
and U842 (N_842,In_0,In_399);
or U843 (N_843,In_227,In_804);
or U844 (N_844,In_711,In_1463);
nand U845 (N_845,In_460,In_18);
nand U846 (N_846,In_163,In_661);
nor U847 (N_847,In_190,In_129);
and U848 (N_848,In_1427,In_921);
nand U849 (N_849,In_520,In_688);
xor U850 (N_850,In_768,In_6);
nor U851 (N_851,In_177,In_1158);
nand U852 (N_852,In_971,In_946);
nand U853 (N_853,In_800,In_1346);
nor U854 (N_854,In_305,In_1216);
and U855 (N_855,In_929,In_1100);
nor U856 (N_856,In_1379,In_50);
nor U857 (N_857,In_630,In_473);
nand U858 (N_858,In_1025,In_439);
nand U859 (N_859,In_641,In_180);
nand U860 (N_860,In_469,In_1295);
and U861 (N_861,In_1492,In_1342);
and U862 (N_862,In_376,In_153);
nor U863 (N_863,In_1378,In_501);
and U864 (N_864,In_1166,In_981);
xor U865 (N_865,In_143,In_1487);
nor U866 (N_866,In_1171,In_735);
nand U867 (N_867,In_1497,In_895);
or U868 (N_868,In_1102,In_986);
nand U869 (N_869,In_1241,In_649);
nand U870 (N_870,In_1443,In_531);
nand U871 (N_871,In_688,In_55);
and U872 (N_872,In_1401,In_150);
or U873 (N_873,In_394,In_492);
nand U874 (N_874,In_167,In_563);
nor U875 (N_875,In_886,In_770);
and U876 (N_876,In_1055,In_351);
or U877 (N_877,In_557,In_433);
and U878 (N_878,In_494,In_539);
or U879 (N_879,In_391,In_516);
nand U880 (N_880,In_786,In_1490);
nor U881 (N_881,In_1234,In_119);
nor U882 (N_882,In_928,In_582);
or U883 (N_883,In_1074,In_1195);
xor U884 (N_884,In_1116,In_1142);
nor U885 (N_885,In_441,In_1378);
and U886 (N_886,In_724,In_1163);
nand U887 (N_887,In_1425,In_1308);
or U888 (N_888,In_794,In_806);
and U889 (N_889,In_741,In_74);
nand U890 (N_890,In_1368,In_1458);
nor U891 (N_891,In_385,In_433);
or U892 (N_892,In_913,In_26);
and U893 (N_893,In_136,In_348);
or U894 (N_894,In_1109,In_67);
xnor U895 (N_895,In_650,In_560);
xnor U896 (N_896,In_25,In_144);
nor U897 (N_897,In_212,In_63);
nor U898 (N_898,In_970,In_1135);
and U899 (N_899,In_681,In_696);
or U900 (N_900,In_1184,In_918);
nor U901 (N_901,In_985,In_458);
nand U902 (N_902,In_397,In_1446);
nor U903 (N_903,In_828,In_1091);
or U904 (N_904,In_65,In_464);
nand U905 (N_905,In_1336,In_274);
xnor U906 (N_906,In_1126,In_849);
nor U907 (N_907,In_250,In_439);
and U908 (N_908,In_1212,In_954);
nor U909 (N_909,In_939,In_1363);
and U910 (N_910,In_916,In_931);
or U911 (N_911,In_188,In_1024);
or U912 (N_912,In_179,In_1076);
nor U913 (N_913,In_668,In_336);
nor U914 (N_914,In_29,In_1288);
and U915 (N_915,In_520,In_997);
nand U916 (N_916,In_814,In_1246);
nand U917 (N_917,In_1496,In_395);
and U918 (N_918,In_495,In_328);
and U919 (N_919,In_1258,In_728);
and U920 (N_920,In_1035,In_18);
nand U921 (N_921,In_632,In_1285);
or U922 (N_922,In_1482,In_791);
xor U923 (N_923,In_1363,In_10);
and U924 (N_924,In_439,In_374);
nor U925 (N_925,In_270,In_130);
nor U926 (N_926,In_645,In_604);
nand U927 (N_927,In_706,In_716);
or U928 (N_928,In_489,In_657);
xnor U929 (N_929,In_731,In_1454);
or U930 (N_930,In_164,In_786);
and U931 (N_931,In_429,In_334);
xor U932 (N_932,In_203,In_715);
or U933 (N_933,In_776,In_217);
nor U934 (N_934,In_329,In_227);
or U935 (N_935,In_1031,In_1234);
or U936 (N_936,In_1408,In_1158);
nor U937 (N_937,In_210,In_209);
nand U938 (N_938,In_594,In_595);
nor U939 (N_939,In_956,In_644);
or U940 (N_940,In_263,In_1034);
nand U941 (N_941,In_388,In_640);
and U942 (N_942,In_760,In_26);
and U943 (N_943,In_24,In_503);
xor U944 (N_944,In_803,In_902);
or U945 (N_945,In_209,In_750);
and U946 (N_946,In_553,In_575);
and U947 (N_947,In_992,In_833);
nor U948 (N_948,In_1178,In_1393);
nor U949 (N_949,In_534,In_206);
and U950 (N_950,In_163,In_1204);
nand U951 (N_951,In_1299,In_1400);
nor U952 (N_952,In_1046,In_1020);
nor U953 (N_953,In_656,In_728);
or U954 (N_954,In_783,In_491);
or U955 (N_955,In_416,In_825);
nor U956 (N_956,In_711,In_1269);
and U957 (N_957,In_272,In_615);
and U958 (N_958,In_738,In_363);
nand U959 (N_959,In_510,In_349);
nand U960 (N_960,In_2,In_1130);
and U961 (N_961,In_1343,In_839);
or U962 (N_962,In_873,In_1396);
xor U963 (N_963,In_1338,In_586);
or U964 (N_964,In_84,In_568);
nor U965 (N_965,In_1330,In_408);
and U966 (N_966,In_8,In_1032);
or U967 (N_967,In_739,In_240);
or U968 (N_968,In_657,In_182);
and U969 (N_969,In_193,In_1123);
xor U970 (N_970,In_728,In_465);
nand U971 (N_971,In_1480,In_565);
nand U972 (N_972,In_1400,In_1282);
xor U973 (N_973,In_519,In_292);
nand U974 (N_974,In_664,In_612);
or U975 (N_975,In_1214,In_1107);
nand U976 (N_976,In_725,In_749);
nand U977 (N_977,In_566,In_385);
and U978 (N_978,In_1285,In_1114);
and U979 (N_979,In_684,In_504);
nor U980 (N_980,In_275,In_283);
or U981 (N_981,In_1461,In_698);
or U982 (N_982,In_439,In_1024);
nand U983 (N_983,In_161,In_1339);
nand U984 (N_984,In_1123,In_214);
and U985 (N_985,In_326,In_520);
nor U986 (N_986,In_451,In_157);
nor U987 (N_987,In_593,In_1248);
and U988 (N_988,In_1122,In_972);
or U989 (N_989,In_319,In_821);
nor U990 (N_990,In_790,In_1340);
nor U991 (N_991,In_1496,In_674);
xor U992 (N_992,In_279,In_868);
nand U993 (N_993,In_1034,In_1262);
and U994 (N_994,In_441,In_1247);
and U995 (N_995,In_1487,In_1454);
nand U996 (N_996,In_261,In_934);
nand U997 (N_997,In_1469,In_200);
or U998 (N_998,In_1363,In_893);
and U999 (N_999,In_523,In_350);
or U1000 (N_1000,In_10,In_1220);
nand U1001 (N_1001,In_107,In_900);
nor U1002 (N_1002,In_428,In_1055);
nand U1003 (N_1003,In_201,In_577);
nand U1004 (N_1004,In_1289,In_1131);
nor U1005 (N_1005,In_516,In_598);
and U1006 (N_1006,In_489,In_611);
xnor U1007 (N_1007,In_626,In_1118);
or U1008 (N_1008,In_853,In_904);
xor U1009 (N_1009,In_135,In_690);
or U1010 (N_1010,In_602,In_1032);
or U1011 (N_1011,In_568,In_1233);
nand U1012 (N_1012,In_731,In_566);
nor U1013 (N_1013,In_1129,In_268);
nor U1014 (N_1014,In_1361,In_388);
nand U1015 (N_1015,In_1401,In_844);
nor U1016 (N_1016,In_1256,In_950);
nand U1017 (N_1017,In_298,In_1297);
and U1018 (N_1018,In_1303,In_861);
or U1019 (N_1019,In_1160,In_793);
and U1020 (N_1020,In_1152,In_454);
and U1021 (N_1021,In_1286,In_631);
and U1022 (N_1022,In_1077,In_1301);
nand U1023 (N_1023,In_1413,In_165);
xor U1024 (N_1024,In_228,In_1387);
nor U1025 (N_1025,In_100,In_673);
or U1026 (N_1026,In_1163,In_1476);
nand U1027 (N_1027,In_777,In_103);
nand U1028 (N_1028,In_808,In_411);
nor U1029 (N_1029,In_209,In_736);
or U1030 (N_1030,In_913,In_1146);
nor U1031 (N_1031,In_1081,In_1075);
nand U1032 (N_1032,In_1116,In_333);
xor U1033 (N_1033,In_927,In_633);
nand U1034 (N_1034,In_1447,In_1306);
and U1035 (N_1035,In_402,In_1317);
or U1036 (N_1036,In_974,In_367);
or U1037 (N_1037,In_523,In_334);
xor U1038 (N_1038,In_205,In_831);
nor U1039 (N_1039,In_496,In_499);
or U1040 (N_1040,In_767,In_1455);
and U1041 (N_1041,In_232,In_723);
xnor U1042 (N_1042,In_267,In_634);
nand U1043 (N_1043,In_369,In_637);
nor U1044 (N_1044,In_1164,In_748);
and U1045 (N_1045,In_658,In_1127);
nor U1046 (N_1046,In_1143,In_355);
and U1047 (N_1047,In_726,In_1497);
nor U1048 (N_1048,In_1428,In_134);
or U1049 (N_1049,In_1160,In_1494);
nor U1050 (N_1050,In_404,In_834);
nor U1051 (N_1051,In_950,In_463);
or U1052 (N_1052,In_233,In_264);
xor U1053 (N_1053,In_283,In_1231);
nor U1054 (N_1054,In_513,In_559);
nand U1055 (N_1055,In_1491,In_1198);
and U1056 (N_1056,In_1085,In_16);
or U1057 (N_1057,In_922,In_425);
nand U1058 (N_1058,In_394,In_340);
nand U1059 (N_1059,In_530,In_1318);
nor U1060 (N_1060,In_156,In_1377);
and U1061 (N_1061,In_688,In_739);
xnor U1062 (N_1062,In_1394,In_1425);
and U1063 (N_1063,In_1123,In_845);
and U1064 (N_1064,In_750,In_378);
nor U1065 (N_1065,In_1228,In_1410);
nor U1066 (N_1066,In_957,In_1024);
nor U1067 (N_1067,In_451,In_318);
nand U1068 (N_1068,In_1000,In_1332);
nand U1069 (N_1069,In_1065,In_1348);
xor U1070 (N_1070,In_880,In_449);
or U1071 (N_1071,In_1331,In_344);
nand U1072 (N_1072,In_1066,In_653);
nor U1073 (N_1073,In_937,In_678);
or U1074 (N_1074,In_1024,In_255);
and U1075 (N_1075,In_248,In_1051);
nor U1076 (N_1076,In_356,In_716);
or U1077 (N_1077,In_1168,In_210);
nand U1078 (N_1078,In_227,In_506);
and U1079 (N_1079,In_883,In_946);
xor U1080 (N_1080,In_1284,In_1296);
or U1081 (N_1081,In_145,In_677);
or U1082 (N_1082,In_1274,In_942);
nand U1083 (N_1083,In_1158,In_1315);
nand U1084 (N_1084,In_640,In_1477);
or U1085 (N_1085,In_538,In_63);
and U1086 (N_1086,In_64,In_839);
or U1087 (N_1087,In_1259,In_406);
or U1088 (N_1088,In_1002,In_1189);
xnor U1089 (N_1089,In_886,In_917);
and U1090 (N_1090,In_810,In_1224);
nand U1091 (N_1091,In_875,In_644);
nor U1092 (N_1092,In_1279,In_939);
or U1093 (N_1093,In_795,In_268);
nand U1094 (N_1094,In_1360,In_1497);
nor U1095 (N_1095,In_1322,In_572);
and U1096 (N_1096,In_1444,In_928);
nand U1097 (N_1097,In_433,In_769);
and U1098 (N_1098,In_1463,In_1469);
or U1099 (N_1099,In_837,In_1047);
xnor U1100 (N_1100,In_1036,In_1068);
xnor U1101 (N_1101,In_662,In_324);
nand U1102 (N_1102,In_740,In_564);
or U1103 (N_1103,In_683,In_341);
nand U1104 (N_1104,In_371,In_558);
and U1105 (N_1105,In_1309,In_925);
xor U1106 (N_1106,In_314,In_385);
nor U1107 (N_1107,In_913,In_23);
or U1108 (N_1108,In_239,In_611);
or U1109 (N_1109,In_122,In_1127);
or U1110 (N_1110,In_199,In_1032);
or U1111 (N_1111,In_937,In_100);
nand U1112 (N_1112,In_1486,In_721);
nor U1113 (N_1113,In_1290,In_872);
and U1114 (N_1114,In_898,In_1445);
nand U1115 (N_1115,In_1325,In_65);
xor U1116 (N_1116,In_1212,In_900);
and U1117 (N_1117,In_145,In_952);
and U1118 (N_1118,In_1383,In_384);
and U1119 (N_1119,In_1093,In_433);
nor U1120 (N_1120,In_699,In_805);
or U1121 (N_1121,In_454,In_1063);
or U1122 (N_1122,In_1412,In_1154);
and U1123 (N_1123,In_994,In_1195);
nand U1124 (N_1124,In_985,In_689);
or U1125 (N_1125,In_562,In_1124);
nand U1126 (N_1126,In_1463,In_1244);
xor U1127 (N_1127,In_1034,In_211);
or U1128 (N_1128,In_186,In_1361);
xnor U1129 (N_1129,In_775,In_847);
nor U1130 (N_1130,In_629,In_124);
or U1131 (N_1131,In_391,In_119);
and U1132 (N_1132,In_22,In_1467);
and U1133 (N_1133,In_1376,In_667);
xor U1134 (N_1134,In_637,In_641);
nand U1135 (N_1135,In_1083,In_943);
or U1136 (N_1136,In_1245,In_632);
or U1137 (N_1137,In_920,In_1350);
and U1138 (N_1138,In_894,In_177);
and U1139 (N_1139,In_321,In_1205);
nand U1140 (N_1140,In_121,In_1444);
nand U1141 (N_1141,In_1007,In_139);
or U1142 (N_1142,In_71,In_635);
nor U1143 (N_1143,In_220,In_186);
xor U1144 (N_1144,In_801,In_1478);
or U1145 (N_1145,In_484,In_1008);
nor U1146 (N_1146,In_275,In_385);
or U1147 (N_1147,In_1226,In_1441);
nand U1148 (N_1148,In_336,In_20);
nor U1149 (N_1149,In_604,In_97);
or U1150 (N_1150,In_312,In_1292);
nor U1151 (N_1151,In_276,In_1155);
nor U1152 (N_1152,In_787,In_1170);
or U1153 (N_1153,In_685,In_464);
xor U1154 (N_1154,In_1418,In_407);
nor U1155 (N_1155,In_53,In_1231);
xor U1156 (N_1156,In_877,In_454);
nand U1157 (N_1157,In_672,In_1111);
or U1158 (N_1158,In_387,In_167);
and U1159 (N_1159,In_1443,In_1195);
nand U1160 (N_1160,In_60,In_199);
nand U1161 (N_1161,In_57,In_533);
xnor U1162 (N_1162,In_257,In_1171);
or U1163 (N_1163,In_854,In_635);
nor U1164 (N_1164,In_969,In_1327);
nor U1165 (N_1165,In_656,In_1046);
or U1166 (N_1166,In_431,In_715);
nand U1167 (N_1167,In_923,In_1490);
nor U1168 (N_1168,In_1320,In_160);
nand U1169 (N_1169,In_849,In_1190);
nand U1170 (N_1170,In_1141,In_958);
and U1171 (N_1171,In_344,In_777);
nand U1172 (N_1172,In_1005,In_178);
nand U1173 (N_1173,In_434,In_967);
and U1174 (N_1174,In_341,In_1123);
or U1175 (N_1175,In_286,In_256);
nor U1176 (N_1176,In_165,In_1248);
nor U1177 (N_1177,In_5,In_762);
or U1178 (N_1178,In_129,In_707);
and U1179 (N_1179,In_1166,In_1381);
nor U1180 (N_1180,In_250,In_1285);
and U1181 (N_1181,In_1402,In_879);
or U1182 (N_1182,In_855,In_1094);
nor U1183 (N_1183,In_917,In_738);
and U1184 (N_1184,In_1273,In_760);
nand U1185 (N_1185,In_603,In_478);
xor U1186 (N_1186,In_773,In_776);
nand U1187 (N_1187,In_239,In_452);
nor U1188 (N_1188,In_467,In_97);
or U1189 (N_1189,In_173,In_841);
nor U1190 (N_1190,In_1494,In_57);
nor U1191 (N_1191,In_789,In_912);
xnor U1192 (N_1192,In_131,In_199);
nor U1193 (N_1193,In_783,In_607);
or U1194 (N_1194,In_1198,In_1103);
nor U1195 (N_1195,In_511,In_297);
xor U1196 (N_1196,In_585,In_42);
or U1197 (N_1197,In_477,In_715);
nand U1198 (N_1198,In_304,In_806);
nor U1199 (N_1199,In_703,In_1048);
or U1200 (N_1200,In_1264,In_349);
or U1201 (N_1201,In_1283,In_1073);
nor U1202 (N_1202,In_436,In_1167);
xnor U1203 (N_1203,In_1134,In_1159);
and U1204 (N_1204,In_46,In_880);
or U1205 (N_1205,In_1204,In_434);
nor U1206 (N_1206,In_791,In_1301);
nor U1207 (N_1207,In_1482,In_1018);
and U1208 (N_1208,In_1306,In_346);
nand U1209 (N_1209,In_822,In_1358);
or U1210 (N_1210,In_281,In_24);
nand U1211 (N_1211,In_1113,In_819);
or U1212 (N_1212,In_304,In_1008);
and U1213 (N_1213,In_162,In_1154);
xor U1214 (N_1214,In_474,In_1413);
or U1215 (N_1215,In_362,In_597);
and U1216 (N_1216,In_226,In_599);
nor U1217 (N_1217,In_609,In_619);
xnor U1218 (N_1218,In_319,In_797);
or U1219 (N_1219,In_728,In_471);
or U1220 (N_1220,In_326,In_523);
or U1221 (N_1221,In_967,In_493);
or U1222 (N_1222,In_507,In_352);
and U1223 (N_1223,In_948,In_417);
nor U1224 (N_1224,In_824,In_921);
or U1225 (N_1225,In_1497,In_936);
or U1226 (N_1226,In_111,In_1135);
or U1227 (N_1227,In_568,In_1091);
and U1228 (N_1228,In_961,In_610);
nor U1229 (N_1229,In_15,In_1100);
and U1230 (N_1230,In_484,In_436);
nand U1231 (N_1231,In_1099,In_578);
nor U1232 (N_1232,In_742,In_173);
and U1233 (N_1233,In_383,In_613);
nand U1234 (N_1234,In_532,In_763);
and U1235 (N_1235,In_435,In_1496);
and U1236 (N_1236,In_1416,In_1114);
xor U1237 (N_1237,In_1056,In_285);
or U1238 (N_1238,In_1227,In_192);
or U1239 (N_1239,In_946,In_1284);
and U1240 (N_1240,In_227,In_936);
nor U1241 (N_1241,In_314,In_890);
nor U1242 (N_1242,In_1199,In_1260);
nand U1243 (N_1243,In_1355,In_200);
or U1244 (N_1244,In_1374,In_784);
xnor U1245 (N_1245,In_1038,In_278);
nor U1246 (N_1246,In_381,In_1105);
or U1247 (N_1247,In_942,In_972);
and U1248 (N_1248,In_50,In_44);
and U1249 (N_1249,In_1023,In_22);
nand U1250 (N_1250,In_875,In_1069);
nor U1251 (N_1251,In_1314,In_613);
nor U1252 (N_1252,In_1270,In_656);
or U1253 (N_1253,In_911,In_816);
and U1254 (N_1254,In_1368,In_881);
or U1255 (N_1255,In_1290,In_114);
and U1256 (N_1256,In_136,In_1490);
or U1257 (N_1257,In_998,In_17);
or U1258 (N_1258,In_1302,In_52);
and U1259 (N_1259,In_1282,In_882);
xnor U1260 (N_1260,In_940,In_671);
nor U1261 (N_1261,In_13,In_343);
and U1262 (N_1262,In_435,In_774);
or U1263 (N_1263,In_288,In_1277);
nand U1264 (N_1264,In_1275,In_772);
nor U1265 (N_1265,In_393,In_1242);
or U1266 (N_1266,In_394,In_956);
xor U1267 (N_1267,In_3,In_477);
or U1268 (N_1268,In_1444,In_336);
and U1269 (N_1269,In_1477,In_1401);
xnor U1270 (N_1270,In_3,In_473);
or U1271 (N_1271,In_867,In_414);
xor U1272 (N_1272,In_739,In_396);
nor U1273 (N_1273,In_872,In_678);
nand U1274 (N_1274,In_43,In_54);
or U1275 (N_1275,In_871,In_179);
and U1276 (N_1276,In_760,In_369);
nor U1277 (N_1277,In_1222,In_730);
or U1278 (N_1278,In_24,In_813);
and U1279 (N_1279,In_743,In_1460);
and U1280 (N_1280,In_499,In_638);
or U1281 (N_1281,In_1193,In_610);
nor U1282 (N_1282,In_162,In_814);
nor U1283 (N_1283,In_275,In_913);
nor U1284 (N_1284,In_1190,In_1472);
or U1285 (N_1285,In_839,In_751);
and U1286 (N_1286,In_492,In_1487);
nor U1287 (N_1287,In_970,In_330);
nor U1288 (N_1288,In_1274,In_1305);
nand U1289 (N_1289,In_315,In_1195);
or U1290 (N_1290,In_693,In_156);
nor U1291 (N_1291,In_1227,In_141);
or U1292 (N_1292,In_699,In_410);
and U1293 (N_1293,In_486,In_386);
xnor U1294 (N_1294,In_730,In_285);
nor U1295 (N_1295,In_555,In_1311);
nor U1296 (N_1296,In_296,In_230);
nor U1297 (N_1297,In_685,In_145);
or U1298 (N_1298,In_410,In_590);
nor U1299 (N_1299,In_1085,In_385);
nor U1300 (N_1300,In_243,In_116);
nand U1301 (N_1301,In_253,In_710);
nand U1302 (N_1302,In_2,In_906);
or U1303 (N_1303,In_1383,In_380);
or U1304 (N_1304,In_245,In_850);
and U1305 (N_1305,In_1258,In_1004);
or U1306 (N_1306,In_437,In_1489);
nor U1307 (N_1307,In_819,In_1095);
and U1308 (N_1308,In_229,In_867);
xor U1309 (N_1309,In_783,In_1274);
or U1310 (N_1310,In_311,In_169);
nand U1311 (N_1311,In_1232,In_222);
xor U1312 (N_1312,In_530,In_1012);
nand U1313 (N_1313,In_631,In_620);
or U1314 (N_1314,In_924,In_217);
nand U1315 (N_1315,In_1357,In_114);
nor U1316 (N_1316,In_713,In_782);
or U1317 (N_1317,In_88,In_251);
or U1318 (N_1318,In_130,In_1197);
nor U1319 (N_1319,In_729,In_1447);
and U1320 (N_1320,In_1377,In_638);
or U1321 (N_1321,In_547,In_186);
nor U1322 (N_1322,In_1476,In_266);
or U1323 (N_1323,In_463,In_1243);
nand U1324 (N_1324,In_991,In_74);
nand U1325 (N_1325,In_387,In_1045);
nor U1326 (N_1326,In_271,In_1156);
or U1327 (N_1327,In_156,In_1331);
nand U1328 (N_1328,In_220,In_540);
or U1329 (N_1329,In_233,In_49);
and U1330 (N_1330,In_524,In_409);
nor U1331 (N_1331,In_760,In_1033);
xnor U1332 (N_1332,In_1107,In_544);
nor U1333 (N_1333,In_1033,In_377);
or U1334 (N_1334,In_519,In_92);
or U1335 (N_1335,In_249,In_304);
nand U1336 (N_1336,In_243,In_1416);
and U1337 (N_1337,In_1303,In_1238);
or U1338 (N_1338,In_1177,In_1157);
and U1339 (N_1339,In_632,In_1484);
nand U1340 (N_1340,In_1408,In_1184);
nand U1341 (N_1341,In_415,In_318);
nor U1342 (N_1342,In_1165,In_1006);
and U1343 (N_1343,In_1147,In_593);
and U1344 (N_1344,In_489,In_622);
xor U1345 (N_1345,In_26,In_1239);
xnor U1346 (N_1346,In_669,In_1273);
or U1347 (N_1347,In_56,In_1459);
and U1348 (N_1348,In_202,In_223);
xor U1349 (N_1349,In_380,In_1205);
nand U1350 (N_1350,In_364,In_743);
or U1351 (N_1351,In_1434,In_608);
or U1352 (N_1352,In_1177,In_285);
nand U1353 (N_1353,In_1155,In_974);
nor U1354 (N_1354,In_1433,In_67);
and U1355 (N_1355,In_119,In_252);
or U1356 (N_1356,In_330,In_681);
and U1357 (N_1357,In_574,In_1366);
nand U1358 (N_1358,In_89,In_392);
nand U1359 (N_1359,In_1065,In_560);
nor U1360 (N_1360,In_413,In_435);
or U1361 (N_1361,In_649,In_1211);
nand U1362 (N_1362,In_140,In_159);
or U1363 (N_1363,In_250,In_807);
and U1364 (N_1364,In_493,In_1204);
nor U1365 (N_1365,In_550,In_563);
xnor U1366 (N_1366,In_1319,In_414);
nand U1367 (N_1367,In_589,In_707);
nand U1368 (N_1368,In_740,In_27);
or U1369 (N_1369,In_961,In_327);
nor U1370 (N_1370,In_94,In_186);
or U1371 (N_1371,In_666,In_663);
and U1372 (N_1372,In_964,In_967);
and U1373 (N_1373,In_1012,In_472);
or U1374 (N_1374,In_1156,In_291);
and U1375 (N_1375,In_946,In_658);
nor U1376 (N_1376,In_384,In_1488);
nor U1377 (N_1377,In_1410,In_456);
xor U1378 (N_1378,In_770,In_207);
nor U1379 (N_1379,In_1490,In_1446);
or U1380 (N_1380,In_419,In_50);
and U1381 (N_1381,In_159,In_1252);
and U1382 (N_1382,In_1084,In_1188);
and U1383 (N_1383,In_139,In_1097);
or U1384 (N_1384,In_1063,In_733);
or U1385 (N_1385,In_409,In_808);
nand U1386 (N_1386,In_964,In_22);
xor U1387 (N_1387,In_1192,In_247);
or U1388 (N_1388,In_1378,In_253);
nor U1389 (N_1389,In_1096,In_801);
nand U1390 (N_1390,In_1234,In_672);
nor U1391 (N_1391,In_111,In_726);
nand U1392 (N_1392,In_679,In_446);
and U1393 (N_1393,In_5,In_818);
nor U1394 (N_1394,In_1104,In_925);
or U1395 (N_1395,In_485,In_581);
nand U1396 (N_1396,In_1482,In_1366);
nand U1397 (N_1397,In_1204,In_456);
nor U1398 (N_1398,In_824,In_1070);
nor U1399 (N_1399,In_191,In_308);
nand U1400 (N_1400,In_280,In_836);
nor U1401 (N_1401,In_695,In_268);
and U1402 (N_1402,In_512,In_999);
and U1403 (N_1403,In_424,In_1073);
nor U1404 (N_1404,In_705,In_1077);
nand U1405 (N_1405,In_941,In_1263);
and U1406 (N_1406,In_1302,In_1330);
nor U1407 (N_1407,In_92,In_1489);
or U1408 (N_1408,In_1301,In_20);
xnor U1409 (N_1409,In_1122,In_37);
nand U1410 (N_1410,In_484,In_673);
xor U1411 (N_1411,In_887,In_520);
nor U1412 (N_1412,In_894,In_172);
nor U1413 (N_1413,In_1309,In_1115);
and U1414 (N_1414,In_1010,In_1404);
and U1415 (N_1415,In_493,In_873);
and U1416 (N_1416,In_153,In_1143);
xnor U1417 (N_1417,In_95,In_1177);
nor U1418 (N_1418,In_1036,In_1428);
nand U1419 (N_1419,In_1045,In_1105);
or U1420 (N_1420,In_1431,In_583);
nor U1421 (N_1421,In_794,In_660);
nor U1422 (N_1422,In_560,In_1059);
and U1423 (N_1423,In_372,In_440);
nand U1424 (N_1424,In_1207,In_551);
xnor U1425 (N_1425,In_552,In_124);
or U1426 (N_1426,In_1003,In_723);
nand U1427 (N_1427,In_812,In_1423);
or U1428 (N_1428,In_308,In_728);
nand U1429 (N_1429,In_309,In_133);
nand U1430 (N_1430,In_1433,In_951);
or U1431 (N_1431,In_16,In_74);
and U1432 (N_1432,In_126,In_1371);
and U1433 (N_1433,In_1085,In_1042);
nor U1434 (N_1434,In_369,In_183);
nand U1435 (N_1435,In_1331,In_645);
nand U1436 (N_1436,In_789,In_1131);
and U1437 (N_1437,In_568,In_1434);
and U1438 (N_1438,In_817,In_1480);
nor U1439 (N_1439,In_1124,In_213);
nor U1440 (N_1440,In_911,In_686);
nor U1441 (N_1441,In_1004,In_179);
and U1442 (N_1442,In_1334,In_467);
and U1443 (N_1443,In_590,In_248);
or U1444 (N_1444,In_1137,In_1467);
nand U1445 (N_1445,In_1323,In_845);
and U1446 (N_1446,In_1192,In_1296);
xnor U1447 (N_1447,In_1399,In_785);
nor U1448 (N_1448,In_939,In_570);
and U1449 (N_1449,In_1175,In_715);
nor U1450 (N_1450,In_1101,In_1404);
nand U1451 (N_1451,In_1233,In_1449);
nor U1452 (N_1452,In_806,In_944);
and U1453 (N_1453,In_531,In_663);
nand U1454 (N_1454,In_671,In_1466);
and U1455 (N_1455,In_981,In_676);
nor U1456 (N_1456,In_931,In_349);
nand U1457 (N_1457,In_657,In_1323);
nand U1458 (N_1458,In_1210,In_1152);
and U1459 (N_1459,In_1286,In_37);
nor U1460 (N_1460,In_623,In_1021);
and U1461 (N_1461,In_1020,In_1323);
nor U1462 (N_1462,In_915,In_44);
nand U1463 (N_1463,In_757,In_1017);
nand U1464 (N_1464,In_10,In_248);
nand U1465 (N_1465,In_557,In_1427);
or U1466 (N_1466,In_387,In_856);
and U1467 (N_1467,In_1408,In_1483);
nor U1468 (N_1468,In_916,In_778);
nand U1469 (N_1469,In_1282,In_1216);
nand U1470 (N_1470,In_287,In_1428);
or U1471 (N_1471,In_1383,In_931);
nand U1472 (N_1472,In_1117,In_664);
and U1473 (N_1473,In_1047,In_476);
or U1474 (N_1474,In_1489,In_253);
nand U1475 (N_1475,In_682,In_195);
or U1476 (N_1476,In_513,In_1274);
nor U1477 (N_1477,In_225,In_424);
nor U1478 (N_1478,In_646,In_1085);
and U1479 (N_1479,In_1485,In_62);
and U1480 (N_1480,In_79,In_209);
and U1481 (N_1481,In_1042,In_399);
nand U1482 (N_1482,In_180,In_374);
xnor U1483 (N_1483,In_1203,In_1053);
and U1484 (N_1484,In_21,In_982);
nand U1485 (N_1485,In_539,In_979);
nor U1486 (N_1486,In_1265,In_1135);
and U1487 (N_1487,In_1062,In_910);
nand U1488 (N_1488,In_200,In_904);
nand U1489 (N_1489,In_1035,In_1157);
or U1490 (N_1490,In_1089,In_1392);
nor U1491 (N_1491,In_1022,In_1361);
xnor U1492 (N_1492,In_137,In_1306);
nor U1493 (N_1493,In_800,In_815);
xnor U1494 (N_1494,In_765,In_526);
or U1495 (N_1495,In_1487,In_795);
and U1496 (N_1496,In_875,In_868);
or U1497 (N_1497,In_226,In_791);
and U1498 (N_1498,In_1091,In_712);
nor U1499 (N_1499,In_1011,In_790);
nand U1500 (N_1500,N_218,N_1477);
nand U1501 (N_1501,N_827,N_166);
nor U1502 (N_1502,N_114,N_377);
nand U1503 (N_1503,N_519,N_388);
and U1504 (N_1504,N_376,N_515);
and U1505 (N_1505,N_821,N_652);
nand U1506 (N_1506,N_1225,N_1167);
nand U1507 (N_1507,N_776,N_1107);
or U1508 (N_1508,N_862,N_1012);
nor U1509 (N_1509,N_354,N_900);
and U1510 (N_1510,N_493,N_834);
xnor U1511 (N_1511,N_846,N_241);
and U1512 (N_1512,N_471,N_344);
and U1513 (N_1513,N_1111,N_614);
nand U1514 (N_1514,N_1089,N_1437);
or U1515 (N_1515,N_1323,N_1258);
and U1516 (N_1516,N_1356,N_486);
xor U1517 (N_1517,N_1267,N_587);
nor U1518 (N_1518,N_865,N_758);
or U1519 (N_1519,N_929,N_221);
and U1520 (N_1520,N_504,N_501);
nor U1521 (N_1521,N_1337,N_603);
or U1522 (N_1522,N_193,N_563);
or U1523 (N_1523,N_693,N_357);
nor U1524 (N_1524,N_1009,N_11);
or U1525 (N_1525,N_1142,N_1499);
or U1526 (N_1526,N_1412,N_286);
nand U1527 (N_1527,N_1261,N_764);
or U1528 (N_1528,N_582,N_932);
or U1529 (N_1529,N_491,N_120);
or U1530 (N_1530,N_886,N_371);
or U1531 (N_1531,N_709,N_295);
nor U1532 (N_1532,N_627,N_1112);
or U1533 (N_1533,N_480,N_439);
nand U1534 (N_1534,N_367,N_1372);
and U1535 (N_1535,N_1404,N_1057);
nor U1536 (N_1536,N_1393,N_1446);
and U1537 (N_1537,N_250,N_421);
xnor U1538 (N_1538,N_847,N_879);
or U1539 (N_1539,N_628,N_269);
or U1540 (N_1540,N_451,N_970);
nor U1541 (N_1541,N_1357,N_204);
nand U1542 (N_1542,N_671,N_1378);
or U1543 (N_1543,N_229,N_601);
or U1544 (N_1544,N_1185,N_490);
nor U1545 (N_1545,N_1215,N_980);
or U1546 (N_1546,N_925,N_706);
and U1547 (N_1547,N_561,N_19);
or U1548 (N_1548,N_1491,N_931);
or U1549 (N_1549,N_972,N_1166);
or U1550 (N_1550,N_502,N_658);
nor U1551 (N_1551,N_757,N_24);
and U1552 (N_1552,N_968,N_347);
nand U1553 (N_1553,N_898,N_498);
nand U1554 (N_1554,N_517,N_1450);
and U1555 (N_1555,N_1483,N_16);
and U1556 (N_1556,N_395,N_368);
nand U1557 (N_1557,N_613,N_456);
nand U1558 (N_1558,N_861,N_130);
nor U1559 (N_1559,N_339,N_753);
and U1560 (N_1560,N_335,N_213);
nand U1561 (N_1561,N_1333,N_997);
xor U1562 (N_1562,N_346,N_1328);
or U1563 (N_1563,N_806,N_280);
xor U1564 (N_1564,N_169,N_650);
or U1565 (N_1565,N_1350,N_1298);
nor U1566 (N_1566,N_1135,N_577);
nand U1567 (N_1567,N_528,N_707);
nor U1568 (N_1568,N_773,N_1196);
or U1569 (N_1569,N_1113,N_793);
nor U1570 (N_1570,N_410,N_768);
nor U1571 (N_1571,N_946,N_1061);
or U1572 (N_1572,N_791,N_180);
nand U1573 (N_1573,N_1115,N_1233);
and U1574 (N_1574,N_1385,N_230);
nand U1575 (N_1575,N_387,N_242);
nor U1576 (N_1576,N_1486,N_722);
nor U1577 (N_1577,N_589,N_217);
nor U1578 (N_1578,N_181,N_850);
nand U1579 (N_1579,N_749,N_401);
nor U1580 (N_1580,N_1432,N_562);
and U1581 (N_1581,N_22,N_303);
and U1582 (N_1582,N_1489,N_141);
or U1583 (N_1583,N_1237,N_1044);
or U1584 (N_1584,N_625,N_161);
xor U1585 (N_1585,N_1133,N_822);
nand U1586 (N_1586,N_164,N_1119);
or U1587 (N_1587,N_632,N_285);
and U1588 (N_1588,N_1152,N_231);
and U1589 (N_1589,N_1314,N_1321);
nor U1590 (N_1590,N_422,N_1076);
and U1591 (N_1591,N_1433,N_730);
nor U1592 (N_1592,N_794,N_802);
and U1593 (N_1593,N_581,N_1081);
and U1594 (N_1594,N_311,N_1439);
nand U1595 (N_1595,N_152,N_187);
nor U1596 (N_1596,N_290,N_369);
xor U1597 (N_1597,N_174,N_678);
or U1598 (N_1598,N_672,N_856);
nor U1599 (N_1599,N_1036,N_267);
nor U1600 (N_1600,N_453,N_1202);
and U1601 (N_1601,N_792,N_873);
nand U1602 (N_1602,N_44,N_389);
nand U1603 (N_1603,N_10,N_1210);
nand U1604 (N_1604,N_1100,N_333);
xor U1605 (N_1605,N_1330,N_844);
and U1606 (N_1606,N_547,N_194);
or U1607 (N_1607,N_179,N_740);
or U1608 (N_1608,N_1183,N_1426);
nand U1609 (N_1609,N_4,N_291);
nand U1610 (N_1610,N_1259,N_49);
or U1611 (N_1611,N_765,N_699);
nand U1612 (N_1612,N_1071,N_511);
or U1613 (N_1613,N_636,N_789);
nor U1614 (N_1614,N_153,N_97);
nand U1615 (N_1615,N_780,N_915);
nand U1616 (N_1616,N_67,N_397);
or U1617 (N_1617,N_405,N_1224);
nand U1618 (N_1618,N_183,N_1286);
nor U1619 (N_1619,N_1200,N_1014);
or U1620 (N_1620,N_341,N_365);
nor U1621 (N_1621,N_969,N_1216);
nand U1622 (N_1622,N_447,N_340);
nor U1623 (N_1623,N_345,N_543);
and U1624 (N_1624,N_40,N_586);
xnor U1625 (N_1625,N_1053,N_415);
nor U1626 (N_1626,N_1129,N_718);
nand U1627 (N_1627,N_1205,N_994);
or U1628 (N_1628,N_1223,N_560);
nor U1629 (N_1629,N_556,N_131);
xor U1630 (N_1630,N_380,N_1230);
or U1631 (N_1631,N_1460,N_1000);
nor U1632 (N_1632,N_1042,N_445);
nand U1633 (N_1633,N_1363,N_665);
nand U1634 (N_1634,N_597,N_1464);
nor U1635 (N_1635,N_739,N_378);
nor U1636 (N_1636,N_403,N_939);
nand U1637 (N_1637,N_619,N_1040);
or U1638 (N_1638,N_147,N_1151);
and U1639 (N_1639,N_578,N_1322);
or U1640 (N_1640,N_647,N_266);
nand U1641 (N_1641,N_1377,N_452);
nand U1642 (N_1642,N_914,N_440);
or U1643 (N_1643,N_808,N_190);
or U1644 (N_1644,N_795,N_866);
and U1645 (N_1645,N_458,N_1257);
nor U1646 (N_1646,N_1279,N_1410);
or U1647 (N_1647,N_362,N_656);
nor U1648 (N_1648,N_721,N_165);
xor U1649 (N_1649,N_653,N_256);
or U1650 (N_1650,N_1045,N_930);
or U1651 (N_1651,N_951,N_503);
and U1652 (N_1652,N_759,N_897);
or U1653 (N_1653,N_558,N_940);
xor U1654 (N_1654,N_818,N_1120);
nor U1655 (N_1655,N_573,N_938);
or U1656 (N_1656,N_1059,N_463);
nor U1657 (N_1657,N_436,N_1398);
and U1658 (N_1658,N_966,N_1461);
and U1659 (N_1659,N_1272,N_1428);
nor U1660 (N_1660,N_1329,N_1271);
or U1661 (N_1661,N_1282,N_959);
or U1662 (N_1662,N_198,N_427);
and U1663 (N_1663,N_323,N_1062);
or U1664 (N_1664,N_513,N_492);
nand U1665 (N_1665,N_983,N_325);
nand U1666 (N_1666,N_418,N_936);
or U1667 (N_1667,N_819,N_37);
and U1668 (N_1668,N_8,N_253);
and U1669 (N_1669,N_1317,N_159);
nor U1670 (N_1670,N_13,N_279);
nor U1671 (N_1671,N_813,N_1452);
nand U1672 (N_1672,N_139,N_684);
nor U1673 (N_1673,N_1043,N_449);
nand U1674 (N_1674,N_352,N_584);
and U1675 (N_1675,N_167,N_1488);
or U1676 (N_1676,N_814,N_408);
and U1677 (N_1677,N_225,N_785);
nand U1678 (N_1678,N_23,N_1197);
or U1679 (N_1679,N_58,N_893);
nor U1680 (N_1680,N_904,N_1025);
or U1681 (N_1681,N_1096,N_76);
and U1682 (N_1682,N_880,N_216);
and U1683 (N_1683,N_934,N_985);
or U1684 (N_1684,N_1281,N_640);
nor U1685 (N_1685,N_510,N_738);
nor U1686 (N_1686,N_145,N_605);
nand U1687 (N_1687,N_289,N_1245);
and U1688 (N_1688,N_1029,N_1239);
xor U1689 (N_1689,N_1265,N_1073);
and U1690 (N_1690,N_843,N_948);
nor U1691 (N_1691,N_824,N_746);
nand U1692 (N_1692,N_276,N_1274);
nor U1693 (N_1693,N_396,N_1019);
or U1694 (N_1694,N_499,N_639);
nand U1695 (N_1695,N_943,N_461);
and U1696 (N_1696,N_129,N_441);
and U1697 (N_1697,N_544,N_1131);
nand U1698 (N_1698,N_1163,N_1332);
nand U1699 (N_1699,N_1026,N_545);
or U1700 (N_1700,N_710,N_1015);
nand U1701 (N_1701,N_1427,N_784);
nor U1702 (N_1702,N_975,N_384);
or U1703 (N_1703,N_783,N_1095);
and U1704 (N_1704,N_1307,N_361);
and U1705 (N_1705,N_782,N_271);
or U1706 (N_1706,N_134,N_111);
nand U1707 (N_1707,N_1132,N_1207);
or U1708 (N_1708,N_48,N_398);
xor U1709 (N_1709,N_1481,N_1003);
nor U1710 (N_1710,N_686,N_1291);
nor U1711 (N_1711,N_328,N_43);
nor U1712 (N_1712,N_1312,N_1208);
and U1713 (N_1713,N_65,N_863);
nor U1714 (N_1714,N_1448,N_1227);
nand U1715 (N_1715,N_1134,N_1313);
nand U1716 (N_1716,N_1300,N_79);
or U1717 (N_1717,N_1381,N_1238);
or U1718 (N_1718,N_443,N_1380);
nor U1719 (N_1719,N_529,N_790);
nor U1720 (N_1720,N_992,N_338);
or U1721 (N_1721,N_105,N_482);
nand U1722 (N_1722,N_1161,N_1295);
and U1723 (N_1723,N_1066,N_976);
or U1724 (N_1724,N_332,N_1214);
xnor U1725 (N_1725,N_595,N_151);
or U1726 (N_1726,N_777,N_84);
nand U1727 (N_1727,N_1054,N_296);
nand U1728 (N_1728,N_500,N_1422);
nor U1729 (N_1729,N_702,N_1386);
nand U1730 (N_1730,N_54,N_786);
and U1731 (N_1731,N_263,N_733);
nor U1732 (N_1732,N_284,N_1174);
nand U1733 (N_1733,N_958,N_68);
or U1734 (N_1734,N_1405,N_487);
nor U1735 (N_1735,N_1253,N_1110);
nor U1736 (N_1736,N_1269,N_17);
and U1737 (N_1737,N_1114,N_826);
and U1738 (N_1738,N_322,N_428);
nor U1739 (N_1739,N_1474,N_3);
xor U1740 (N_1740,N_1084,N_743);
nand U1741 (N_1741,N_1479,N_1434);
nor U1742 (N_1742,N_287,N_26);
or U1743 (N_1743,N_1440,N_849);
and U1744 (N_1744,N_60,N_591);
or U1745 (N_1745,N_1088,N_747);
nor U1746 (N_1746,N_809,N_497);
xor U1747 (N_1747,N_767,N_1423);
nor U1748 (N_1748,N_27,N_1374);
nor U1749 (N_1749,N_1429,N_805);
nor U1750 (N_1750,N_524,N_756);
nor U1751 (N_1751,N_126,N_891);
and U1752 (N_1752,N_655,N_1229);
xnor U1753 (N_1753,N_1010,N_425);
or U1754 (N_1754,N_1361,N_1090);
nor U1755 (N_1755,N_1204,N_402);
and U1756 (N_1756,N_184,N_884);
or U1757 (N_1757,N_1348,N_246);
nand U1758 (N_1758,N_189,N_1123);
or U1759 (N_1759,N_797,N_356);
or U1760 (N_1760,N_192,N_803);
nand U1761 (N_1761,N_919,N_771);
nor U1762 (N_1762,N_1168,N_888);
nor U1763 (N_1763,N_927,N_80);
nor U1764 (N_1764,N_600,N_518);
nor U1765 (N_1765,N_608,N_1487);
or U1766 (N_1766,N_649,N_996);
or U1767 (N_1767,N_400,N_1341);
and U1768 (N_1768,N_31,N_761);
and U1769 (N_1769,N_588,N_66);
and U1770 (N_1770,N_644,N_546);
or U1771 (N_1771,N_375,N_760);
or U1772 (N_1772,N_478,N_56);
xor U1773 (N_1773,N_788,N_472);
nor U1774 (N_1774,N_481,N_485);
nand U1775 (N_1775,N_676,N_53);
nand U1776 (N_1776,N_1454,N_697);
nor U1777 (N_1777,N_1158,N_1050);
and U1778 (N_1778,N_1343,N_583);
nand U1779 (N_1779,N_1376,N_137);
xnor U1780 (N_1780,N_751,N_540);
nand U1781 (N_1781,N_52,N_232);
and U1782 (N_1782,N_1340,N_1251);
and U1783 (N_1783,N_1222,N_1453);
and U1784 (N_1784,N_615,N_1401);
and U1785 (N_1785,N_1389,N_1425);
or U1786 (N_1786,N_1463,N_57);
nand U1787 (N_1787,N_298,N_538);
nand U1788 (N_1788,N_342,N_437);
and U1789 (N_1789,N_1455,N_720);
nand U1790 (N_1790,N_1156,N_567);
nand U1791 (N_1791,N_306,N_299);
xor U1792 (N_1792,N_1247,N_728);
and U1793 (N_1793,N_1149,N_1130);
and U1794 (N_1794,N_651,N_799);
xnor U1795 (N_1795,N_146,N_313);
and U1796 (N_1796,N_909,N_574);
xnor U1797 (N_1797,N_737,N_370);
or U1798 (N_1798,N_406,N_1028);
xor U1799 (N_1799,N_248,N_667);
nor U1800 (N_1800,N_1234,N_1480);
and U1801 (N_1801,N_1419,N_477);
nor U1802 (N_1802,N_81,N_177);
nand U1803 (N_1803,N_811,N_1209);
and U1804 (N_1804,N_7,N_2);
nor U1805 (N_1805,N_358,N_373);
and U1806 (N_1806,N_235,N_1470);
xor U1807 (N_1807,N_366,N_264);
and U1808 (N_1808,N_1417,N_305);
and U1809 (N_1809,N_1153,N_1394);
xor U1810 (N_1810,N_536,N_292);
xnor U1811 (N_1811,N_315,N_386);
xnor U1812 (N_1812,N_300,N_916);
nand U1813 (N_1813,N_454,N_233);
nand U1814 (N_1814,N_407,N_727);
nand U1815 (N_1815,N_662,N_205);
and U1816 (N_1816,N_1495,N_801);
nand U1817 (N_1817,N_896,N_1033);
nand U1818 (N_1818,N_1139,N_95);
or U1819 (N_1819,N_281,N_864);
or U1820 (N_1820,N_1218,N_330);
and U1821 (N_1821,N_1327,N_1415);
nor U1822 (N_1822,N_1387,N_45);
nor U1823 (N_1823,N_839,N_1442);
nand U1824 (N_1824,N_355,N_476);
nor U1825 (N_1825,N_1031,N_1018);
nand U1826 (N_1826,N_918,N_1353);
or U1827 (N_1827,N_572,N_956);
and U1828 (N_1828,N_1497,N_611);
nand U1829 (N_1829,N_838,N_91);
or U1830 (N_1830,N_566,N_1263);
xnor U1831 (N_1831,N_155,N_555);
nor U1832 (N_1832,N_118,N_201);
xnor U1833 (N_1833,N_138,N_1369);
and U1834 (N_1834,N_175,N_1324);
nor U1835 (N_1835,N_942,N_537);
nand U1836 (N_1836,N_668,N_553);
and U1837 (N_1837,N_1346,N_55);
or U1838 (N_1838,N_73,N_1436);
nor U1839 (N_1839,N_1005,N_430);
nor U1840 (N_1840,N_475,N_1485);
nand U1841 (N_1841,N_1254,N_987);
xnor U1842 (N_1842,N_157,N_535);
xor U1843 (N_1843,N_239,N_1297);
nor U1844 (N_1844,N_1288,N_1220);
nor U1845 (N_1845,N_1368,N_1217);
xor U1846 (N_1846,N_1468,N_324);
or U1847 (N_1847,N_735,N_435);
and U1848 (N_1848,N_1030,N_754);
nor U1849 (N_1849,N_92,N_673);
or U1850 (N_1850,N_715,N_1391);
xnor U1851 (N_1851,N_1087,N_1256);
nand U1852 (N_1852,N_1373,N_913);
nand U1853 (N_1853,N_908,N_1235);
nor U1854 (N_1854,N_964,N_331);
nand U1855 (N_1855,N_820,N_307);
nand U1856 (N_1856,N_734,N_1124);
or U1857 (N_1857,N_921,N_1409);
nand U1858 (N_1858,N_197,N_549);
or U1859 (N_1859,N_237,N_320);
nor U1860 (N_1860,N_1072,N_390);
or U1861 (N_1861,N_1178,N_1459);
xnor U1862 (N_1862,N_209,N_351);
nor U1863 (N_1863,N_411,N_579);
and U1864 (N_1864,N_1413,N_714);
and U1865 (N_1865,N_1165,N_265);
nand U1866 (N_1866,N_663,N_182);
nand U1867 (N_1867,N_986,N_116);
and U1868 (N_1868,N_1125,N_698);
and U1869 (N_1869,N_1482,N_832);
nor U1870 (N_1870,N_829,N_1325);
nor U1871 (N_1871,N_890,N_115);
and U1872 (N_1872,N_853,N_30);
or U1873 (N_1873,N_1308,N_12);
nor U1874 (N_1874,N_688,N_25);
xor U1875 (N_1875,N_1462,N_643);
or U1876 (N_1876,N_399,N_314);
or U1877 (N_1877,N_319,N_282);
xnor U1878 (N_1878,N_383,N_701);
xor U1879 (N_1879,N_828,N_1347);
nor U1880 (N_1880,N_1024,N_1086);
nand U1881 (N_1881,N_1358,N_318);
and U1882 (N_1882,N_554,N_874);
or U1883 (N_1883,N_1342,N_70);
and U1884 (N_1884,N_1335,N_755);
xnor U1885 (N_1885,N_1206,N_110);
or U1886 (N_1886,N_1293,N_1458);
and U1887 (N_1887,N_766,N_1083);
or U1888 (N_1888,N_160,N_1336);
xor U1889 (N_1889,N_855,N_128);
nand U1890 (N_1890,N_618,N_188);
xnor U1891 (N_1891,N_1157,N_1211);
xor U1892 (N_1892,N_816,N_1078);
xnor U1893 (N_1893,N_675,N_1475);
nand U1894 (N_1894,N_877,N_1188);
and U1895 (N_1895,N_532,N_831);
and U1896 (N_1896,N_283,N_542);
nand U1897 (N_1897,N_1023,N_1296);
nand U1898 (N_1898,N_962,N_1243);
nand U1899 (N_1899,N_1219,N_920);
nor U1900 (N_1900,N_132,N_531);
and U1901 (N_1901,N_876,N_1289);
or U1902 (N_1902,N_1035,N_228);
or U1903 (N_1903,N_88,N_859);
nor U1904 (N_1904,N_657,N_779);
and U1905 (N_1905,N_541,N_316);
nor U1906 (N_1906,N_1292,N_1456);
nor U1907 (N_1907,N_1077,N_123);
or U1908 (N_1908,N_158,N_262);
nand U1909 (N_1909,N_1406,N_273);
and U1910 (N_1910,N_1118,N_1193);
and U1911 (N_1911,N_1349,N_1146);
nor U1912 (N_1912,N_593,N_691);
nand U1913 (N_1913,N_769,N_1365);
nand U1914 (N_1914,N_108,N_1169);
and U1915 (N_1915,N_885,N_385);
or U1916 (N_1916,N_329,N_1424);
nand U1917 (N_1917,N_1266,N_965);
nand U1918 (N_1918,N_364,N_326);
nand U1919 (N_1919,N_878,N_270);
and U1920 (N_1920,N_669,N_1469);
nand U1921 (N_1921,N_261,N_381);
nand U1922 (N_1922,N_121,N_1299);
nor U1923 (N_1923,N_1354,N_1320);
or U1924 (N_1924,N_752,N_349);
and U1925 (N_1925,N_1304,N_508);
and U1926 (N_1926,N_1260,N_744);
nor U1927 (N_1927,N_1067,N_170);
nand U1928 (N_1928,N_641,N_87);
nand U1929 (N_1929,N_33,N_494);
nor U1930 (N_1930,N_1284,N_1060);
and U1931 (N_1931,N_729,N_419);
nor U1932 (N_1932,N_1172,N_633);
and U1933 (N_1933,N_473,N_244);
nand U1934 (N_1934,N_1148,N_1283);
nor U1935 (N_1935,N_176,N_1303);
nand U1936 (N_1936,N_124,N_882);
or U1937 (N_1937,N_798,N_787);
nand U1938 (N_1938,N_220,N_840);
nor U1939 (N_1939,N_215,N_1476);
nor U1940 (N_1940,N_417,N_414);
nor U1941 (N_1941,N_1127,N_89);
or U1942 (N_1942,N_1242,N_1136);
and U1943 (N_1943,N_903,N_631);
and U1944 (N_1944,N_1221,N_569);
or U1945 (N_1945,N_995,N_372);
xnor U1946 (N_1946,N_570,N_450);
and U1947 (N_1947,N_1290,N_29);
or U1948 (N_1948,N_599,N_858);
nand U1949 (N_1949,N_1140,N_150);
or U1950 (N_1950,N_214,N_1075);
and U1951 (N_1951,N_967,N_1103);
xnor U1952 (N_1952,N_199,N_868);
and U1953 (N_1953,N_1408,N_690);
and U1954 (N_1954,N_99,N_719);
nor U1955 (N_1955,N_695,N_680);
nor U1956 (N_1956,N_78,N_38);
and U1957 (N_1957,N_1435,N_867);
or U1958 (N_1958,N_464,N_35);
and U1959 (N_1959,N_148,N_963);
or U1960 (N_1960,N_781,N_240);
or U1961 (N_1961,N_774,N_1232);
nand U1962 (N_1962,N_252,N_947);
and U1963 (N_1963,N_926,N_1117);
nand U1964 (N_1964,N_1187,N_1264);
and U1965 (N_1965,N_924,N_526);
or U1966 (N_1966,N_1164,N_149);
and U1967 (N_1967,N_571,N_1109);
nand U1968 (N_1968,N_724,N_807);
nand U1969 (N_1969,N_1085,N_61);
nor U1970 (N_1970,N_1301,N_106);
nor U1971 (N_1971,N_1318,N_18);
and U1972 (N_1972,N_991,N_534);
or U1973 (N_1973,N_1038,N_899);
nor U1974 (N_1974,N_413,N_1101);
nor U1975 (N_1975,N_21,N_14);
nand U1976 (N_1976,N_1375,N_96);
or U1977 (N_1977,N_1315,N_604);
nor U1978 (N_1978,N_1370,N_1143);
or U1979 (N_1979,N_207,N_1447);
nand U1980 (N_1980,N_64,N_870);
nand U1981 (N_1981,N_664,N_1244);
nand U1982 (N_1982,N_171,N_634);
nand U1983 (N_1983,N_654,N_800);
nor U1984 (N_1984,N_509,N_1277);
or U1985 (N_1985,N_1063,N_1102);
or U1986 (N_1986,N_630,N_1198);
xnor U1987 (N_1987,N_382,N_848);
nor U1988 (N_1988,N_564,N_750);
xor U1989 (N_1989,N_258,N_810);
xor U1990 (N_1990,N_103,N_304);
nor U1991 (N_1991,N_1493,N_394);
nand U1992 (N_1992,N_1180,N_135);
and U1993 (N_1993,N_682,N_39);
nor U1994 (N_1994,N_1116,N_1013);
nand U1995 (N_1995,N_426,N_15);
and U1996 (N_1996,N_1457,N_516);
nor U1997 (N_1997,N_1065,N_446);
xnor U1998 (N_1998,N_119,N_923);
or U1999 (N_1999,N_6,N_359);
and U2000 (N_2000,N_666,N_71);
or U2001 (N_2001,N_895,N_1016);
xnor U2002 (N_2002,N_700,N_1175);
nand U2003 (N_2003,N_69,N_211);
nand U2004 (N_2004,N_1122,N_1021);
nand U2005 (N_2005,N_1362,N_1184);
nand U2006 (N_2006,N_1310,N_72);
nor U2007 (N_2007,N_857,N_548);
xnor U2008 (N_2008,N_1159,N_255);
or U2009 (N_2009,N_905,N_527);
nor U2010 (N_2010,N_195,N_716);
and U2011 (N_2011,N_635,N_1046);
xnor U2012 (N_2012,N_140,N_1186);
or U2013 (N_2013,N_465,N_1388);
and U2014 (N_2014,N_902,N_1181);
nand U2015 (N_2015,N_467,N_694);
nand U2016 (N_2016,N_741,N_42);
nor U2017 (N_2017,N_83,N_208);
nor U2018 (N_2018,N_901,N_815);
and U2019 (N_2019,N_1002,N_978);
nand U2020 (N_2020,N_954,N_1064);
xnor U2021 (N_2021,N_871,N_957);
or U2022 (N_2022,N_1212,N_28);
and U2023 (N_2023,N_565,N_685);
nand U2024 (N_2024,N_429,N_1311);
nor U2025 (N_2025,N_881,N_1007);
nand U2026 (N_2026,N_1392,N_460);
and U2027 (N_2027,N_622,N_825);
nor U2028 (N_2028,N_278,N_1141);
xnor U2029 (N_2029,N_1270,N_112);
nor U2030 (N_2030,N_607,N_185);
nand U2031 (N_2031,N_745,N_1097);
and U2032 (N_2032,N_254,N_277);
and U2033 (N_2033,N_122,N_945);
nor U2034 (N_2034,N_1400,N_889);
xor U2035 (N_2035,N_136,N_955);
nor U2036 (N_2036,N_661,N_869);
and U2037 (N_2037,N_1231,N_1001);
nand U2038 (N_2038,N_196,N_683);
or U2039 (N_2039,N_1199,N_1438);
nand U2040 (N_2040,N_260,N_1176);
xor U2041 (N_2041,N_1047,N_1445);
and U2042 (N_2042,N_1294,N_448);
xnor U2043 (N_2043,N_598,N_696);
and U2044 (N_2044,N_842,N_1416);
or U2045 (N_2045,N_444,N_872);
and U2046 (N_2046,N_712,N_272);
and U2047 (N_2047,N_725,N_717);
and U2048 (N_2048,N_557,N_1384);
or U2049 (N_2049,N_41,N_226);
or U2050 (N_2050,N_883,N_1);
xor U2051 (N_2051,N_93,N_294);
xnor U2052 (N_2052,N_1248,N_1331);
or U2053 (N_2053,N_982,N_539);
nand U2054 (N_2054,N_1498,N_496);
nand U2055 (N_2055,N_186,N_830);
and U2056 (N_2056,N_1367,N_1352);
nand U2057 (N_2057,N_257,N_1171);
nor U2058 (N_2058,N_961,N_1364);
and U2059 (N_2059,N_455,N_1451);
xnor U2060 (N_2060,N_1213,N_1032);
xor U2061 (N_2061,N_736,N_732);
nor U2062 (N_2062,N_90,N_142);
and U2063 (N_2063,N_1179,N_952);
nand U2064 (N_2064,N_552,N_979);
or U2065 (N_2065,N_949,N_156);
nor U2066 (N_2066,N_1020,N_894);
and U2067 (N_2067,N_1195,N_687);
or U2068 (N_2068,N_1011,N_268);
or U2069 (N_2069,N_47,N_1444);
and U2070 (N_2070,N_297,N_1048);
or U2071 (N_2071,N_59,N_1170);
nand U2072 (N_2072,N_117,N_993);
nor U2073 (N_2073,N_404,N_293);
and U2074 (N_2074,N_202,N_1051);
nand U2075 (N_2075,N_833,N_9);
nor U2076 (N_2076,N_416,N_505);
or U2077 (N_2077,N_1431,N_1371);
nand U2078 (N_2078,N_506,N_34);
nor U2079 (N_2079,N_409,N_1056);
nor U2080 (N_2080,N_484,N_32);
nand U2081 (N_2081,N_1236,N_275);
or U2082 (N_2082,N_742,N_778);
and U2083 (N_2083,N_1402,N_576);
and U2084 (N_2084,N_1121,N_1004);
xor U2085 (N_2085,N_343,N_1411);
nand U2086 (N_2086,N_999,N_1275);
or U2087 (N_2087,N_520,N_337);
xor U2088 (N_2088,N_679,N_1467);
nand U2089 (N_2089,N_845,N_1108);
nor U2090 (N_2090,N_935,N_852);
xnor U2091 (N_2091,N_726,N_1147);
nand U2092 (N_2092,N_1360,N_1074);
xnor U2093 (N_2093,N_243,N_507);
nand U2094 (N_2094,N_1414,N_1104);
nand U2095 (N_2095,N_1226,N_775);
or U2096 (N_2096,N_1144,N_36);
xor U2097 (N_2097,N_353,N_1273);
nand U2098 (N_2098,N_236,N_629);
or U2099 (N_2099,N_1278,N_249);
or U2100 (N_2100,N_1055,N_907);
or U2101 (N_2101,N_1407,N_247);
or U2102 (N_2102,N_227,N_770);
nor U2103 (N_2103,N_162,N_1150);
or U2104 (N_2104,N_1162,N_1092);
or U2105 (N_2105,N_1490,N_432);
nand U2106 (N_2106,N_708,N_575);
xor U2107 (N_2107,N_163,N_1079);
xor U2108 (N_2108,N_602,N_200);
nand U2109 (N_2109,N_1155,N_626);
nand U2110 (N_2110,N_168,N_1098);
and U2111 (N_2111,N_1177,N_1154);
nand U2112 (N_2112,N_1246,N_1344);
xor U2113 (N_2113,N_1355,N_474);
nand U2114 (N_2114,N_100,N_1441);
and U2115 (N_2115,N_144,N_420);
or U2116 (N_2116,N_74,N_1397);
nor U2117 (N_2117,N_1099,N_178);
or U2118 (N_2118,N_1203,N_470);
nor U2119 (N_2119,N_887,N_998);
nand U2120 (N_2120,N_521,N_1145);
or U2121 (N_2121,N_1396,N_391);
or U2122 (N_2122,N_606,N_841);
or U2123 (N_2123,N_1189,N_875);
or U2124 (N_2124,N_812,N_312);
nand U2125 (N_2125,N_1466,N_512);
or U2126 (N_2126,N_1262,N_1250);
nor U2127 (N_2127,N_1137,N_1082);
nor U2128 (N_2128,N_203,N_1091);
nand U2129 (N_2129,N_219,N_748);
nand U2130 (N_2130,N_988,N_525);
nor U2131 (N_2131,N_836,N_1228);
and U2132 (N_2132,N_1041,N_1068);
or U2133 (N_2133,N_483,N_94);
nand U2134 (N_2134,N_568,N_1070);
or U2135 (N_2135,N_392,N_1390);
nand U2136 (N_2136,N_660,N_172);
or U2137 (N_2137,N_1338,N_1473);
or U2138 (N_2138,N_837,N_514);
or U2139 (N_2139,N_703,N_670);
nand U2140 (N_2140,N_125,N_645);
nor U2141 (N_2141,N_224,N_86);
or U2142 (N_2142,N_1190,N_620);
or U2143 (N_2143,N_1191,N_309);
or U2144 (N_2144,N_288,N_251);
and U2145 (N_2145,N_704,N_533);
nand U2146 (N_2146,N_46,N_933);
and U2147 (N_2147,N_911,N_977);
and U2148 (N_2148,N_692,N_1182);
and U2149 (N_2149,N_206,N_723);
nand U2150 (N_2150,N_638,N_1496);
xor U2151 (N_2151,N_336,N_1022);
xor U2152 (N_2152,N_610,N_1403);
nand U2153 (N_2153,N_1008,N_468);
xnor U2154 (N_2154,N_0,N_621);
nand U2155 (N_2155,N_523,N_941);
nand U2156 (N_2156,N_950,N_1094);
or U2157 (N_2157,N_51,N_590);
nand U2158 (N_2158,N_469,N_5);
or U2159 (N_2159,N_62,N_1049);
or U2160 (N_2160,N_559,N_1334);
and U2161 (N_2161,N_1249,N_522);
nand U2162 (N_2162,N_711,N_981);
or U2163 (N_2163,N_127,N_1285);
xnor U2164 (N_2164,N_772,N_1449);
nand U2165 (N_2165,N_1430,N_1255);
xnor U2166 (N_2166,N_960,N_133);
or U2167 (N_2167,N_310,N_1106);
nor U2168 (N_2168,N_1126,N_609);
or U2169 (N_2169,N_212,N_245);
or U2170 (N_2170,N_301,N_1339);
nand U2171 (N_2171,N_642,N_191);
and U2172 (N_2172,N_360,N_143);
or U2173 (N_2173,N_1494,N_624);
or U2174 (N_2174,N_442,N_763);
nand U2175 (N_2175,N_85,N_350);
nand U2176 (N_2176,N_1037,N_580);
nand U2177 (N_2177,N_101,N_1276);
or U2178 (N_2178,N_804,N_989);
and U2179 (N_2179,N_796,N_851);
and U2180 (N_2180,N_912,N_823);
xnor U2181 (N_2181,N_434,N_689);
and U2182 (N_2182,N_1201,N_393);
nand U2183 (N_2183,N_1302,N_713);
or U2184 (N_2184,N_107,N_1359);
nor U2185 (N_2185,N_1418,N_596);
or U2186 (N_2186,N_1173,N_222);
and U2187 (N_2187,N_860,N_705);
or U2188 (N_2188,N_922,N_1316);
or U2189 (N_2189,N_1484,N_82);
nand U2190 (N_2190,N_104,N_1395);
or U2191 (N_2191,N_50,N_77);
nand U2192 (N_2192,N_835,N_731);
xnor U2193 (N_2193,N_308,N_1309);
nand U2194 (N_2194,N_1240,N_928);
nand U2195 (N_2195,N_892,N_1241);
nor U2196 (N_2196,N_612,N_1027);
or U2197 (N_2197,N_334,N_1471);
and U2198 (N_2198,N_906,N_1034);
and U2199 (N_2199,N_412,N_585);
nor U2200 (N_2200,N_1138,N_223);
or U2201 (N_2201,N_990,N_1160);
and U2202 (N_2202,N_637,N_154);
or U2203 (N_2203,N_937,N_1492);
nand U2204 (N_2204,N_327,N_1287);
nor U2205 (N_2205,N_495,N_1420);
or U2206 (N_2206,N_423,N_466);
nor U2207 (N_2207,N_98,N_1268);
nor U2208 (N_2208,N_113,N_530);
or U2209 (N_2209,N_1069,N_462);
nor U2210 (N_2210,N_321,N_374);
and U2211 (N_2211,N_944,N_1280);
and U2212 (N_2212,N_63,N_363);
nor U2213 (N_2213,N_1006,N_1326);
nor U2214 (N_2214,N_102,N_1379);
and U2215 (N_2215,N_1192,N_424);
or U2216 (N_2216,N_1382,N_75);
xnor U2217 (N_2217,N_1052,N_910);
or U2218 (N_2218,N_1306,N_1465);
or U2219 (N_2219,N_762,N_917);
nor U2220 (N_2220,N_274,N_1319);
nor U2221 (N_2221,N_550,N_210);
and U2222 (N_2222,N_1478,N_302);
or U2223 (N_2223,N_317,N_1105);
nand U2224 (N_2224,N_1039,N_1351);
nand U2225 (N_2225,N_971,N_20);
nor U2226 (N_2226,N_677,N_1399);
nor U2227 (N_2227,N_1252,N_973);
or U2228 (N_2228,N_1366,N_488);
nor U2229 (N_2229,N_1472,N_974);
nand U2230 (N_2230,N_459,N_623);
nor U2231 (N_2231,N_551,N_489);
and U2232 (N_2232,N_348,N_1305);
xor U2233 (N_2233,N_1345,N_431);
and U2234 (N_2234,N_1093,N_1421);
xor U2235 (N_2235,N_173,N_438);
or U2236 (N_2236,N_109,N_433);
or U2237 (N_2237,N_648,N_681);
nand U2238 (N_2238,N_953,N_659);
and U2239 (N_2239,N_457,N_238);
nand U2240 (N_2240,N_479,N_234);
or U2241 (N_2241,N_817,N_379);
nand U2242 (N_2242,N_259,N_1128);
and U2243 (N_2243,N_1058,N_1194);
nand U2244 (N_2244,N_617,N_616);
and U2245 (N_2245,N_854,N_594);
and U2246 (N_2246,N_674,N_984);
nand U2247 (N_2247,N_1017,N_1443);
nor U2248 (N_2248,N_592,N_646);
nand U2249 (N_2249,N_1383,N_1080);
nor U2250 (N_2250,N_678,N_363);
nand U2251 (N_2251,N_1212,N_96);
xor U2252 (N_2252,N_1097,N_937);
nor U2253 (N_2253,N_423,N_909);
xnor U2254 (N_2254,N_1381,N_229);
nand U2255 (N_2255,N_40,N_279);
nand U2256 (N_2256,N_704,N_1032);
nand U2257 (N_2257,N_1313,N_1304);
nand U2258 (N_2258,N_664,N_64);
and U2259 (N_2259,N_791,N_1258);
nor U2260 (N_2260,N_10,N_32);
nand U2261 (N_2261,N_383,N_417);
nor U2262 (N_2262,N_357,N_1068);
xor U2263 (N_2263,N_508,N_502);
nor U2264 (N_2264,N_508,N_821);
and U2265 (N_2265,N_1400,N_1263);
xnor U2266 (N_2266,N_881,N_857);
and U2267 (N_2267,N_1029,N_865);
or U2268 (N_2268,N_969,N_446);
nor U2269 (N_2269,N_1114,N_537);
nand U2270 (N_2270,N_989,N_770);
nor U2271 (N_2271,N_555,N_672);
nor U2272 (N_2272,N_873,N_657);
nor U2273 (N_2273,N_430,N_433);
and U2274 (N_2274,N_400,N_1265);
or U2275 (N_2275,N_386,N_550);
nand U2276 (N_2276,N_797,N_754);
nor U2277 (N_2277,N_370,N_25);
or U2278 (N_2278,N_1359,N_398);
nand U2279 (N_2279,N_1252,N_1497);
or U2280 (N_2280,N_355,N_34);
and U2281 (N_2281,N_896,N_707);
nand U2282 (N_2282,N_14,N_867);
nor U2283 (N_2283,N_1201,N_1377);
nor U2284 (N_2284,N_213,N_1252);
nor U2285 (N_2285,N_180,N_1455);
xnor U2286 (N_2286,N_265,N_291);
nor U2287 (N_2287,N_3,N_1235);
nand U2288 (N_2288,N_1030,N_923);
nor U2289 (N_2289,N_984,N_1458);
nor U2290 (N_2290,N_1308,N_799);
or U2291 (N_2291,N_325,N_766);
or U2292 (N_2292,N_753,N_700);
nand U2293 (N_2293,N_169,N_768);
and U2294 (N_2294,N_1476,N_941);
or U2295 (N_2295,N_941,N_256);
and U2296 (N_2296,N_898,N_632);
or U2297 (N_2297,N_58,N_1086);
or U2298 (N_2298,N_232,N_938);
nor U2299 (N_2299,N_214,N_353);
nor U2300 (N_2300,N_1145,N_1498);
and U2301 (N_2301,N_748,N_862);
and U2302 (N_2302,N_931,N_950);
nor U2303 (N_2303,N_1181,N_1477);
or U2304 (N_2304,N_23,N_635);
or U2305 (N_2305,N_979,N_275);
and U2306 (N_2306,N_170,N_1235);
and U2307 (N_2307,N_654,N_453);
or U2308 (N_2308,N_375,N_1470);
or U2309 (N_2309,N_426,N_609);
xor U2310 (N_2310,N_472,N_1484);
nor U2311 (N_2311,N_1140,N_1136);
or U2312 (N_2312,N_1290,N_922);
nor U2313 (N_2313,N_1324,N_437);
and U2314 (N_2314,N_1384,N_1356);
nor U2315 (N_2315,N_1082,N_25);
or U2316 (N_2316,N_975,N_959);
or U2317 (N_2317,N_189,N_1221);
nor U2318 (N_2318,N_1359,N_1393);
and U2319 (N_2319,N_1486,N_1359);
nand U2320 (N_2320,N_1228,N_308);
xor U2321 (N_2321,N_1390,N_379);
or U2322 (N_2322,N_1495,N_235);
and U2323 (N_2323,N_1127,N_116);
nand U2324 (N_2324,N_1087,N_451);
nor U2325 (N_2325,N_903,N_431);
or U2326 (N_2326,N_1199,N_424);
xnor U2327 (N_2327,N_15,N_1413);
nand U2328 (N_2328,N_324,N_1195);
nand U2329 (N_2329,N_972,N_785);
or U2330 (N_2330,N_652,N_127);
or U2331 (N_2331,N_1361,N_444);
nor U2332 (N_2332,N_88,N_499);
nand U2333 (N_2333,N_1216,N_334);
nor U2334 (N_2334,N_366,N_1443);
xor U2335 (N_2335,N_3,N_952);
nor U2336 (N_2336,N_78,N_1282);
nor U2337 (N_2337,N_1143,N_91);
nand U2338 (N_2338,N_145,N_140);
or U2339 (N_2339,N_1169,N_1235);
xor U2340 (N_2340,N_239,N_315);
nand U2341 (N_2341,N_488,N_43);
nor U2342 (N_2342,N_1278,N_669);
nor U2343 (N_2343,N_1266,N_1214);
nor U2344 (N_2344,N_181,N_1096);
or U2345 (N_2345,N_1244,N_460);
and U2346 (N_2346,N_1168,N_928);
nand U2347 (N_2347,N_545,N_1316);
nand U2348 (N_2348,N_748,N_896);
and U2349 (N_2349,N_113,N_467);
xnor U2350 (N_2350,N_1019,N_1079);
xnor U2351 (N_2351,N_199,N_979);
and U2352 (N_2352,N_655,N_749);
xnor U2353 (N_2353,N_168,N_1326);
nor U2354 (N_2354,N_188,N_1265);
xor U2355 (N_2355,N_461,N_260);
nor U2356 (N_2356,N_139,N_1453);
nand U2357 (N_2357,N_270,N_1025);
and U2358 (N_2358,N_473,N_422);
nor U2359 (N_2359,N_517,N_452);
nand U2360 (N_2360,N_1091,N_318);
or U2361 (N_2361,N_477,N_213);
nor U2362 (N_2362,N_1279,N_993);
and U2363 (N_2363,N_142,N_992);
nand U2364 (N_2364,N_1026,N_747);
nand U2365 (N_2365,N_192,N_538);
nor U2366 (N_2366,N_1187,N_863);
or U2367 (N_2367,N_1313,N_1432);
and U2368 (N_2368,N_876,N_93);
nor U2369 (N_2369,N_1172,N_274);
or U2370 (N_2370,N_68,N_232);
and U2371 (N_2371,N_954,N_457);
or U2372 (N_2372,N_171,N_1190);
nand U2373 (N_2373,N_972,N_586);
or U2374 (N_2374,N_943,N_713);
and U2375 (N_2375,N_427,N_1272);
xnor U2376 (N_2376,N_676,N_736);
or U2377 (N_2377,N_1358,N_1108);
and U2378 (N_2378,N_1368,N_48);
nor U2379 (N_2379,N_720,N_257);
and U2380 (N_2380,N_1294,N_1366);
or U2381 (N_2381,N_1089,N_44);
nand U2382 (N_2382,N_1202,N_162);
and U2383 (N_2383,N_1062,N_890);
nand U2384 (N_2384,N_639,N_1410);
nor U2385 (N_2385,N_1418,N_1212);
nand U2386 (N_2386,N_361,N_535);
nor U2387 (N_2387,N_1464,N_890);
nor U2388 (N_2388,N_1246,N_823);
nand U2389 (N_2389,N_219,N_1022);
and U2390 (N_2390,N_409,N_281);
and U2391 (N_2391,N_857,N_555);
nor U2392 (N_2392,N_658,N_1380);
or U2393 (N_2393,N_383,N_545);
nor U2394 (N_2394,N_1150,N_582);
and U2395 (N_2395,N_120,N_472);
nor U2396 (N_2396,N_1452,N_739);
or U2397 (N_2397,N_660,N_830);
or U2398 (N_2398,N_869,N_778);
nor U2399 (N_2399,N_1161,N_599);
and U2400 (N_2400,N_1248,N_221);
nor U2401 (N_2401,N_1087,N_843);
or U2402 (N_2402,N_1345,N_811);
nand U2403 (N_2403,N_624,N_1055);
nand U2404 (N_2404,N_401,N_920);
nand U2405 (N_2405,N_293,N_1303);
or U2406 (N_2406,N_371,N_713);
nand U2407 (N_2407,N_218,N_1476);
and U2408 (N_2408,N_927,N_25);
nor U2409 (N_2409,N_180,N_1014);
and U2410 (N_2410,N_362,N_544);
nor U2411 (N_2411,N_514,N_29);
and U2412 (N_2412,N_1329,N_787);
nor U2413 (N_2413,N_208,N_1136);
nand U2414 (N_2414,N_1362,N_1427);
xor U2415 (N_2415,N_689,N_367);
nor U2416 (N_2416,N_1345,N_1229);
or U2417 (N_2417,N_473,N_166);
and U2418 (N_2418,N_898,N_720);
nor U2419 (N_2419,N_211,N_934);
nor U2420 (N_2420,N_1330,N_1310);
and U2421 (N_2421,N_1156,N_957);
nand U2422 (N_2422,N_901,N_467);
or U2423 (N_2423,N_1389,N_1326);
nand U2424 (N_2424,N_1039,N_1035);
nor U2425 (N_2425,N_1439,N_776);
or U2426 (N_2426,N_940,N_821);
nor U2427 (N_2427,N_972,N_1145);
nand U2428 (N_2428,N_650,N_53);
nand U2429 (N_2429,N_287,N_126);
xnor U2430 (N_2430,N_653,N_1049);
xor U2431 (N_2431,N_1034,N_1173);
or U2432 (N_2432,N_1099,N_1426);
nand U2433 (N_2433,N_388,N_1269);
xnor U2434 (N_2434,N_481,N_895);
nand U2435 (N_2435,N_41,N_679);
nor U2436 (N_2436,N_906,N_1009);
or U2437 (N_2437,N_478,N_1139);
or U2438 (N_2438,N_58,N_1184);
nor U2439 (N_2439,N_101,N_599);
nand U2440 (N_2440,N_1282,N_228);
nand U2441 (N_2441,N_1284,N_535);
nand U2442 (N_2442,N_78,N_1273);
nor U2443 (N_2443,N_382,N_949);
xnor U2444 (N_2444,N_901,N_566);
and U2445 (N_2445,N_890,N_682);
and U2446 (N_2446,N_221,N_375);
nand U2447 (N_2447,N_143,N_708);
nand U2448 (N_2448,N_1401,N_1472);
and U2449 (N_2449,N_866,N_156);
and U2450 (N_2450,N_1286,N_1499);
and U2451 (N_2451,N_926,N_783);
xnor U2452 (N_2452,N_69,N_1158);
or U2453 (N_2453,N_1306,N_1429);
nor U2454 (N_2454,N_624,N_969);
nor U2455 (N_2455,N_591,N_959);
nor U2456 (N_2456,N_1490,N_31);
nor U2457 (N_2457,N_1147,N_331);
nor U2458 (N_2458,N_238,N_454);
nor U2459 (N_2459,N_688,N_198);
nand U2460 (N_2460,N_1320,N_634);
and U2461 (N_2461,N_125,N_0);
or U2462 (N_2462,N_186,N_121);
and U2463 (N_2463,N_1305,N_995);
nand U2464 (N_2464,N_386,N_1042);
nand U2465 (N_2465,N_821,N_1282);
or U2466 (N_2466,N_255,N_1009);
xor U2467 (N_2467,N_763,N_121);
nand U2468 (N_2468,N_580,N_186);
and U2469 (N_2469,N_151,N_869);
xor U2470 (N_2470,N_157,N_1364);
and U2471 (N_2471,N_561,N_386);
xnor U2472 (N_2472,N_815,N_1095);
and U2473 (N_2473,N_1347,N_882);
xnor U2474 (N_2474,N_10,N_865);
nand U2475 (N_2475,N_683,N_432);
nor U2476 (N_2476,N_948,N_132);
and U2477 (N_2477,N_480,N_626);
nand U2478 (N_2478,N_888,N_1322);
nand U2479 (N_2479,N_1263,N_894);
and U2480 (N_2480,N_679,N_1236);
nand U2481 (N_2481,N_645,N_595);
nand U2482 (N_2482,N_917,N_1294);
nor U2483 (N_2483,N_1454,N_844);
and U2484 (N_2484,N_836,N_972);
nor U2485 (N_2485,N_1030,N_628);
nand U2486 (N_2486,N_574,N_772);
nand U2487 (N_2487,N_648,N_1377);
nor U2488 (N_2488,N_167,N_1078);
nor U2489 (N_2489,N_1217,N_290);
xor U2490 (N_2490,N_1437,N_1198);
nand U2491 (N_2491,N_1403,N_880);
and U2492 (N_2492,N_892,N_864);
or U2493 (N_2493,N_376,N_405);
and U2494 (N_2494,N_1294,N_1359);
and U2495 (N_2495,N_222,N_731);
nor U2496 (N_2496,N_1368,N_1383);
nand U2497 (N_2497,N_643,N_19);
and U2498 (N_2498,N_210,N_661);
xor U2499 (N_2499,N_519,N_910);
nor U2500 (N_2500,N_607,N_1302);
nor U2501 (N_2501,N_164,N_70);
or U2502 (N_2502,N_385,N_131);
nor U2503 (N_2503,N_1325,N_338);
xor U2504 (N_2504,N_937,N_228);
nor U2505 (N_2505,N_1223,N_951);
and U2506 (N_2506,N_632,N_1304);
nor U2507 (N_2507,N_706,N_1123);
and U2508 (N_2508,N_342,N_1045);
or U2509 (N_2509,N_1265,N_770);
and U2510 (N_2510,N_352,N_748);
and U2511 (N_2511,N_550,N_1207);
or U2512 (N_2512,N_1187,N_1020);
nor U2513 (N_2513,N_839,N_197);
nand U2514 (N_2514,N_585,N_1102);
or U2515 (N_2515,N_1322,N_897);
nor U2516 (N_2516,N_356,N_1270);
nand U2517 (N_2517,N_557,N_611);
nand U2518 (N_2518,N_784,N_1122);
and U2519 (N_2519,N_311,N_898);
or U2520 (N_2520,N_3,N_530);
nor U2521 (N_2521,N_1488,N_765);
nor U2522 (N_2522,N_150,N_262);
xnor U2523 (N_2523,N_6,N_1312);
xor U2524 (N_2524,N_600,N_958);
xnor U2525 (N_2525,N_1028,N_867);
and U2526 (N_2526,N_106,N_397);
nor U2527 (N_2527,N_390,N_257);
nor U2528 (N_2528,N_533,N_979);
xnor U2529 (N_2529,N_1067,N_1224);
or U2530 (N_2530,N_1120,N_597);
nand U2531 (N_2531,N_559,N_882);
or U2532 (N_2532,N_967,N_717);
and U2533 (N_2533,N_25,N_785);
and U2534 (N_2534,N_1412,N_244);
nand U2535 (N_2535,N_931,N_638);
xor U2536 (N_2536,N_921,N_1031);
nand U2537 (N_2537,N_611,N_16);
or U2538 (N_2538,N_1271,N_743);
xor U2539 (N_2539,N_1349,N_449);
and U2540 (N_2540,N_597,N_562);
nand U2541 (N_2541,N_1017,N_958);
nor U2542 (N_2542,N_1334,N_764);
or U2543 (N_2543,N_417,N_1174);
nor U2544 (N_2544,N_249,N_1357);
or U2545 (N_2545,N_461,N_1293);
xor U2546 (N_2546,N_91,N_346);
nand U2547 (N_2547,N_1313,N_278);
and U2548 (N_2548,N_684,N_107);
xnor U2549 (N_2549,N_1296,N_545);
nand U2550 (N_2550,N_266,N_962);
nor U2551 (N_2551,N_1128,N_347);
or U2552 (N_2552,N_1301,N_884);
or U2553 (N_2553,N_1104,N_114);
or U2554 (N_2554,N_1457,N_191);
xor U2555 (N_2555,N_425,N_595);
nor U2556 (N_2556,N_1025,N_935);
nand U2557 (N_2557,N_610,N_1063);
or U2558 (N_2558,N_603,N_1034);
nor U2559 (N_2559,N_1128,N_195);
nand U2560 (N_2560,N_571,N_395);
and U2561 (N_2561,N_663,N_525);
and U2562 (N_2562,N_1415,N_181);
or U2563 (N_2563,N_619,N_1282);
nor U2564 (N_2564,N_27,N_1361);
or U2565 (N_2565,N_397,N_434);
nand U2566 (N_2566,N_68,N_1337);
nor U2567 (N_2567,N_614,N_5);
nor U2568 (N_2568,N_880,N_149);
nor U2569 (N_2569,N_964,N_961);
and U2570 (N_2570,N_1407,N_1121);
or U2571 (N_2571,N_955,N_1229);
or U2572 (N_2572,N_1217,N_519);
nor U2573 (N_2573,N_906,N_188);
or U2574 (N_2574,N_1119,N_1065);
nor U2575 (N_2575,N_1359,N_571);
or U2576 (N_2576,N_963,N_675);
or U2577 (N_2577,N_810,N_149);
or U2578 (N_2578,N_281,N_1111);
nor U2579 (N_2579,N_1221,N_655);
and U2580 (N_2580,N_365,N_715);
and U2581 (N_2581,N_215,N_1117);
or U2582 (N_2582,N_1250,N_318);
and U2583 (N_2583,N_1224,N_1099);
and U2584 (N_2584,N_1149,N_518);
nand U2585 (N_2585,N_1392,N_1480);
nand U2586 (N_2586,N_949,N_1109);
or U2587 (N_2587,N_830,N_1101);
or U2588 (N_2588,N_379,N_218);
nor U2589 (N_2589,N_182,N_220);
or U2590 (N_2590,N_1021,N_544);
or U2591 (N_2591,N_899,N_1414);
nand U2592 (N_2592,N_1107,N_901);
or U2593 (N_2593,N_83,N_616);
nand U2594 (N_2594,N_1124,N_912);
nor U2595 (N_2595,N_778,N_269);
nand U2596 (N_2596,N_350,N_222);
nand U2597 (N_2597,N_937,N_399);
nand U2598 (N_2598,N_804,N_56);
nor U2599 (N_2599,N_627,N_588);
and U2600 (N_2600,N_403,N_673);
and U2601 (N_2601,N_1074,N_237);
and U2602 (N_2602,N_92,N_173);
xnor U2603 (N_2603,N_1083,N_972);
and U2604 (N_2604,N_1215,N_237);
or U2605 (N_2605,N_49,N_248);
nand U2606 (N_2606,N_350,N_972);
xnor U2607 (N_2607,N_1445,N_50);
and U2608 (N_2608,N_1014,N_1148);
xnor U2609 (N_2609,N_191,N_1036);
and U2610 (N_2610,N_10,N_839);
and U2611 (N_2611,N_405,N_1089);
nor U2612 (N_2612,N_992,N_429);
or U2613 (N_2613,N_75,N_1125);
or U2614 (N_2614,N_196,N_296);
or U2615 (N_2615,N_418,N_1371);
and U2616 (N_2616,N_391,N_1197);
nand U2617 (N_2617,N_691,N_1165);
and U2618 (N_2618,N_1417,N_652);
and U2619 (N_2619,N_644,N_982);
nand U2620 (N_2620,N_488,N_500);
or U2621 (N_2621,N_131,N_687);
or U2622 (N_2622,N_1470,N_1188);
nor U2623 (N_2623,N_325,N_191);
nor U2624 (N_2624,N_721,N_915);
nor U2625 (N_2625,N_361,N_969);
and U2626 (N_2626,N_626,N_695);
xnor U2627 (N_2627,N_1209,N_240);
nor U2628 (N_2628,N_830,N_1293);
or U2629 (N_2629,N_201,N_1249);
or U2630 (N_2630,N_239,N_299);
xnor U2631 (N_2631,N_633,N_1296);
and U2632 (N_2632,N_1180,N_23);
and U2633 (N_2633,N_381,N_630);
or U2634 (N_2634,N_540,N_1365);
and U2635 (N_2635,N_59,N_285);
nand U2636 (N_2636,N_102,N_228);
and U2637 (N_2637,N_670,N_334);
nand U2638 (N_2638,N_647,N_307);
or U2639 (N_2639,N_840,N_839);
xor U2640 (N_2640,N_805,N_332);
nor U2641 (N_2641,N_1137,N_944);
and U2642 (N_2642,N_544,N_152);
or U2643 (N_2643,N_205,N_833);
nand U2644 (N_2644,N_635,N_265);
nor U2645 (N_2645,N_356,N_1222);
and U2646 (N_2646,N_434,N_933);
nand U2647 (N_2647,N_365,N_1298);
nor U2648 (N_2648,N_921,N_289);
or U2649 (N_2649,N_1388,N_452);
nor U2650 (N_2650,N_1026,N_582);
nor U2651 (N_2651,N_974,N_283);
xor U2652 (N_2652,N_1465,N_1302);
nor U2653 (N_2653,N_1421,N_829);
and U2654 (N_2654,N_619,N_1175);
and U2655 (N_2655,N_1068,N_324);
nand U2656 (N_2656,N_501,N_650);
or U2657 (N_2657,N_509,N_716);
nor U2658 (N_2658,N_750,N_379);
or U2659 (N_2659,N_26,N_902);
nor U2660 (N_2660,N_967,N_292);
or U2661 (N_2661,N_589,N_395);
or U2662 (N_2662,N_1219,N_479);
or U2663 (N_2663,N_459,N_939);
nor U2664 (N_2664,N_612,N_233);
or U2665 (N_2665,N_283,N_142);
and U2666 (N_2666,N_1153,N_1264);
xnor U2667 (N_2667,N_214,N_561);
nor U2668 (N_2668,N_142,N_191);
xor U2669 (N_2669,N_854,N_1283);
or U2670 (N_2670,N_1211,N_1303);
and U2671 (N_2671,N_1344,N_371);
nand U2672 (N_2672,N_1126,N_173);
xnor U2673 (N_2673,N_1102,N_400);
xnor U2674 (N_2674,N_1236,N_364);
and U2675 (N_2675,N_39,N_1462);
and U2676 (N_2676,N_437,N_508);
and U2677 (N_2677,N_1320,N_778);
or U2678 (N_2678,N_724,N_1355);
xor U2679 (N_2679,N_85,N_767);
nand U2680 (N_2680,N_211,N_662);
and U2681 (N_2681,N_926,N_104);
or U2682 (N_2682,N_1352,N_879);
nand U2683 (N_2683,N_461,N_52);
and U2684 (N_2684,N_553,N_775);
and U2685 (N_2685,N_739,N_543);
xor U2686 (N_2686,N_894,N_253);
nor U2687 (N_2687,N_735,N_1120);
nand U2688 (N_2688,N_12,N_1091);
nand U2689 (N_2689,N_816,N_1398);
nor U2690 (N_2690,N_369,N_124);
nor U2691 (N_2691,N_80,N_489);
xor U2692 (N_2692,N_226,N_847);
nor U2693 (N_2693,N_136,N_400);
nor U2694 (N_2694,N_107,N_1009);
and U2695 (N_2695,N_1363,N_1040);
nand U2696 (N_2696,N_100,N_875);
or U2697 (N_2697,N_1116,N_345);
nor U2698 (N_2698,N_232,N_804);
nand U2699 (N_2699,N_610,N_297);
xnor U2700 (N_2700,N_1020,N_1052);
and U2701 (N_2701,N_1448,N_713);
or U2702 (N_2702,N_118,N_861);
and U2703 (N_2703,N_1048,N_152);
and U2704 (N_2704,N_137,N_1);
xor U2705 (N_2705,N_714,N_779);
xor U2706 (N_2706,N_380,N_1411);
or U2707 (N_2707,N_1093,N_1077);
nand U2708 (N_2708,N_1318,N_77);
and U2709 (N_2709,N_50,N_41);
xnor U2710 (N_2710,N_571,N_931);
nor U2711 (N_2711,N_1172,N_654);
nand U2712 (N_2712,N_1042,N_225);
and U2713 (N_2713,N_167,N_1148);
or U2714 (N_2714,N_693,N_237);
nand U2715 (N_2715,N_97,N_1187);
and U2716 (N_2716,N_317,N_589);
xor U2717 (N_2717,N_1159,N_1003);
or U2718 (N_2718,N_998,N_137);
or U2719 (N_2719,N_1024,N_713);
or U2720 (N_2720,N_385,N_1133);
xnor U2721 (N_2721,N_749,N_432);
nor U2722 (N_2722,N_1429,N_349);
nor U2723 (N_2723,N_426,N_227);
or U2724 (N_2724,N_94,N_408);
nor U2725 (N_2725,N_1376,N_1390);
and U2726 (N_2726,N_903,N_36);
nor U2727 (N_2727,N_365,N_944);
nand U2728 (N_2728,N_1166,N_1352);
nor U2729 (N_2729,N_1024,N_916);
and U2730 (N_2730,N_494,N_602);
and U2731 (N_2731,N_230,N_1449);
nor U2732 (N_2732,N_1333,N_447);
and U2733 (N_2733,N_1039,N_1311);
or U2734 (N_2734,N_525,N_41);
and U2735 (N_2735,N_1115,N_353);
nor U2736 (N_2736,N_855,N_853);
nor U2737 (N_2737,N_1431,N_1451);
or U2738 (N_2738,N_382,N_1004);
nor U2739 (N_2739,N_399,N_640);
nand U2740 (N_2740,N_1103,N_802);
and U2741 (N_2741,N_163,N_625);
or U2742 (N_2742,N_153,N_1036);
and U2743 (N_2743,N_603,N_1033);
xnor U2744 (N_2744,N_837,N_178);
nand U2745 (N_2745,N_1350,N_636);
nand U2746 (N_2746,N_226,N_355);
nand U2747 (N_2747,N_989,N_696);
or U2748 (N_2748,N_252,N_737);
nor U2749 (N_2749,N_288,N_444);
or U2750 (N_2750,N_50,N_970);
nand U2751 (N_2751,N_184,N_701);
nor U2752 (N_2752,N_86,N_642);
xor U2753 (N_2753,N_949,N_252);
or U2754 (N_2754,N_143,N_1289);
nor U2755 (N_2755,N_577,N_1022);
xor U2756 (N_2756,N_406,N_510);
nand U2757 (N_2757,N_1299,N_917);
or U2758 (N_2758,N_1385,N_443);
or U2759 (N_2759,N_1420,N_723);
nand U2760 (N_2760,N_508,N_184);
xor U2761 (N_2761,N_1379,N_656);
and U2762 (N_2762,N_380,N_389);
nand U2763 (N_2763,N_795,N_1082);
or U2764 (N_2764,N_700,N_1046);
nand U2765 (N_2765,N_1314,N_264);
nand U2766 (N_2766,N_146,N_1170);
nand U2767 (N_2767,N_572,N_525);
nand U2768 (N_2768,N_403,N_590);
or U2769 (N_2769,N_214,N_571);
xnor U2770 (N_2770,N_1206,N_364);
or U2771 (N_2771,N_184,N_709);
nor U2772 (N_2772,N_23,N_1255);
and U2773 (N_2773,N_471,N_1441);
nor U2774 (N_2774,N_154,N_437);
xnor U2775 (N_2775,N_145,N_1231);
nor U2776 (N_2776,N_1289,N_1166);
nand U2777 (N_2777,N_799,N_712);
nor U2778 (N_2778,N_28,N_770);
nor U2779 (N_2779,N_1057,N_235);
nor U2780 (N_2780,N_983,N_1212);
and U2781 (N_2781,N_803,N_522);
and U2782 (N_2782,N_864,N_510);
and U2783 (N_2783,N_161,N_1053);
nor U2784 (N_2784,N_42,N_1401);
or U2785 (N_2785,N_989,N_1336);
nand U2786 (N_2786,N_273,N_917);
nand U2787 (N_2787,N_658,N_747);
and U2788 (N_2788,N_1299,N_1346);
and U2789 (N_2789,N_818,N_852);
and U2790 (N_2790,N_1480,N_1180);
and U2791 (N_2791,N_17,N_1046);
nor U2792 (N_2792,N_969,N_620);
or U2793 (N_2793,N_1294,N_454);
nor U2794 (N_2794,N_1463,N_375);
nor U2795 (N_2795,N_1421,N_1396);
nand U2796 (N_2796,N_93,N_1249);
nand U2797 (N_2797,N_542,N_50);
and U2798 (N_2798,N_1119,N_986);
or U2799 (N_2799,N_41,N_744);
or U2800 (N_2800,N_1076,N_1063);
nand U2801 (N_2801,N_1069,N_1165);
xor U2802 (N_2802,N_419,N_616);
nor U2803 (N_2803,N_45,N_483);
or U2804 (N_2804,N_248,N_93);
xnor U2805 (N_2805,N_167,N_1261);
and U2806 (N_2806,N_54,N_850);
nand U2807 (N_2807,N_411,N_992);
xnor U2808 (N_2808,N_85,N_1296);
nor U2809 (N_2809,N_774,N_1212);
nor U2810 (N_2810,N_1367,N_142);
and U2811 (N_2811,N_1124,N_439);
and U2812 (N_2812,N_46,N_748);
nand U2813 (N_2813,N_1038,N_361);
or U2814 (N_2814,N_1442,N_1135);
nand U2815 (N_2815,N_674,N_907);
nor U2816 (N_2816,N_781,N_1284);
or U2817 (N_2817,N_28,N_1400);
and U2818 (N_2818,N_1389,N_775);
nor U2819 (N_2819,N_1256,N_880);
and U2820 (N_2820,N_1091,N_1423);
xnor U2821 (N_2821,N_1291,N_761);
and U2822 (N_2822,N_1086,N_418);
or U2823 (N_2823,N_471,N_117);
nand U2824 (N_2824,N_823,N_1393);
xor U2825 (N_2825,N_645,N_1476);
nand U2826 (N_2826,N_1291,N_823);
nand U2827 (N_2827,N_369,N_94);
nor U2828 (N_2828,N_983,N_474);
xnor U2829 (N_2829,N_1048,N_18);
and U2830 (N_2830,N_1069,N_706);
nand U2831 (N_2831,N_227,N_794);
xor U2832 (N_2832,N_980,N_1293);
and U2833 (N_2833,N_427,N_70);
nor U2834 (N_2834,N_140,N_360);
nand U2835 (N_2835,N_211,N_11);
nor U2836 (N_2836,N_901,N_140);
nor U2837 (N_2837,N_1075,N_1322);
and U2838 (N_2838,N_1236,N_395);
nor U2839 (N_2839,N_718,N_1287);
nand U2840 (N_2840,N_1464,N_1357);
or U2841 (N_2841,N_801,N_1068);
nand U2842 (N_2842,N_731,N_439);
nand U2843 (N_2843,N_13,N_1465);
nand U2844 (N_2844,N_462,N_504);
nor U2845 (N_2845,N_1311,N_396);
or U2846 (N_2846,N_862,N_1320);
nand U2847 (N_2847,N_685,N_229);
nand U2848 (N_2848,N_785,N_1284);
nor U2849 (N_2849,N_1014,N_963);
nand U2850 (N_2850,N_113,N_354);
and U2851 (N_2851,N_1017,N_303);
or U2852 (N_2852,N_909,N_1400);
and U2853 (N_2853,N_1077,N_512);
and U2854 (N_2854,N_1279,N_1168);
or U2855 (N_2855,N_104,N_435);
and U2856 (N_2856,N_815,N_1417);
and U2857 (N_2857,N_800,N_1286);
and U2858 (N_2858,N_107,N_1101);
or U2859 (N_2859,N_1418,N_816);
nand U2860 (N_2860,N_1216,N_1067);
nor U2861 (N_2861,N_622,N_714);
xor U2862 (N_2862,N_1341,N_758);
nand U2863 (N_2863,N_525,N_77);
and U2864 (N_2864,N_671,N_155);
nand U2865 (N_2865,N_1168,N_855);
nand U2866 (N_2866,N_335,N_163);
nand U2867 (N_2867,N_1120,N_426);
or U2868 (N_2868,N_636,N_823);
or U2869 (N_2869,N_1326,N_1247);
nand U2870 (N_2870,N_469,N_798);
or U2871 (N_2871,N_1005,N_57);
or U2872 (N_2872,N_1104,N_453);
nor U2873 (N_2873,N_881,N_597);
nor U2874 (N_2874,N_315,N_128);
nor U2875 (N_2875,N_413,N_1340);
or U2876 (N_2876,N_1434,N_1134);
nand U2877 (N_2877,N_1043,N_1490);
nand U2878 (N_2878,N_913,N_1193);
nor U2879 (N_2879,N_983,N_976);
or U2880 (N_2880,N_1185,N_1120);
nand U2881 (N_2881,N_1211,N_51);
nand U2882 (N_2882,N_1408,N_704);
nor U2883 (N_2883,N_1014,N_36);
nand U2884 (N_2884,N_948,N_319);
nand U2885 (N_2885,N_976,N_675);
nand U2886 (N_2886,N_980,N_265);
or U2887 (N_2887,N_900,N_789);
or U2888 (N_2888,N_184,N_98);
nor U2889 (N_2889,N_858,N_795);
nand U2890 (N_2890,N_1421,N_777);
nor U2891 (N_2891,N_734,N_1471);
nor U2892 (N_2892,N_1259,N_1060);
and U2893 (N_2893,N_929,N_1422);
xor U2894 (N_2894,N_787,N_24);
or U2895 (N_2895,N_782,N_370);
xor U2896 (N_2896,N_736,N_1239);
nor U2897 (N_2897,N_634,N_318);
xor U2898 (N_2898,N_1299,N_419);
nand U2899 (N_2899,N_593,N_332);
nor U2900 (N_2900,N_560,N_365);
nor U2901 (N_2901,N_605,N_4);
or U2902 (N_2902,N_1383,N_1336);
nor U2903 (N_2903,N_172,N_430);
nand U2904 (N_2904,N_999,N_118);
or U2905 (N_2905,N_927,N_1045);
or U2906 (N_2906,N_1324,N_1117);
and U2907 (N_2907,N_662,N_271);
nand U2908 (N_2908,N_73,N_153);
and U2909 (N_2909,N_362,N_189);
nor U2910 (N_2910,N_822,N_1127);
nor U2911 (N_2911,N_1307,N_381);
xnor U2912 (N_2912,N_810,N_890);
xnor U2913 (N_2913,N_1194,N_238);
nor U2914 (N_2914,N_989,N_595);
nor U2915 (N_2915,N_52,N_81);
or U2916 (N_2916,N_1314,N_371);
xnor U2917 (N_2917,N_1426,N_842);
and U2918 (N_2918,N_1113,N_383);
and U2919 (N_2919,N_1138,N_1207);
nand U2920 (N_2920,N_65,N_732);
nand U2921 (N_2921,N_628,N_1076);
and U2922 (N_2922,N_1156,N_1432);
xnor U2923 (N_2923,N_1226,N_153);
nor U2924 (N_2924,N_1208,N_495);
and U2925 (N_2925,N_1361,N_494);
or U2926 (N_2926,N_341,N_748);
nor U2927 (N_2927,N_236,N_271);
nand U2928 (N_2928,N_1310,N_962);
nor U2929 (N_2929,N_1333,N_1181);
nand U2930 (N_2930,N_1358,N_141);
or U2931 (N_2931,N_1128,N_752);
and U2932 (N_2932,N_222,N_408);
or U2933 (N_2933,N_1061,N_834);
or U2934 (N_2934,N_254,N_722);
or U2935 (N_2935,N_291,N_680);
nand U2936 (N_2936,N_789,N_1310);
nor U2937 (N_2937,N_1376,N_489);
or U2938 (N_2938,N_114,N_527);
and U2939 (N_2939,N_826,N_945);
and U2940 (N_2940,N_1391,N_1380);
nor U2941 (N_2941,N_474,N_358);
and U2942 (N_2942,N_188,N_552);
nand U2943 (N_2943,N_1290,N_1267);
and U2944 (N_2944,N_1193,N_1089);
or U2945 (N_2945,N_128,N_426);
nand U2946 (N_2946,N_353,N_1279);
or U2947 (N_2947,N_283,N_234);
nor U2948 (N_2948,N_1019,N_763);
or U2949 (N_2949,N_523,N_558);
and U2950 (N_2950,N_690,N_25);
and U2951 (N_2951,N_341,N_917);
or U2952 (N_2952,N_1016,N_443);
or U2953 (N_2953,N_479,N_1163);
or U2954 (N_2954,N_1219,N_1121);
or U2955 (N_2955,N_34,N_660);
nor U2956 (N_2956,N_1010,N_73);
and U2957 (N_2957,N_279,N_841);
nor U2958 (N_2958,N_863,N_53);
or U2959 (N_2959,N_1488,N_565);
nand U2960 (N_2960,N_1381,N_1158);
and U2961 (N_2961,N_1467,N_162);
xor U2962 (N_2962,N_1031,N_948);
nor U2963 (N_2963,N_332,N_939);
nor U2964 (N_2964,N_1345,N_696);
or U2965 (N_2965,N_1151,N_1219);
xor U2966 (N_2966,N_935,N_479);
or U2967 (N_2967,N_1426,N_838);
nand U2968 (N_2968,N_780,N_311);
nor U2969 (N_2969,N_1056,N_1040);
nand U2970 (N_2970,N_124,N_986);
nand U2971 (N_2971,N_654,N_952);
xor U2972 (N_2972,N_550,N_143);
nor U2973 (N_2973,N_541,N_833);
or U2974 (N_2974,N_1064,N_114);
xnor U2975 (N_2975,N_345,N_1436);
and U2976 (N_2976,N_697,N_217);
nand U2977 (N_2977,N_728,N_152);
nand U2978 (N_2978,N_594,N_266);
and U2979 (N_2979,N_1318,N_708);
and U2980 (N_2980,N_828,N_159);
xor U2981 (N_2981,N_733,N_353);
nor U2982 (N_2982,N_1197,N_1486);
nor U2983 (N_2983,N_516,N_549);
or U2984 (N_2984,N_657,N_93);
and U2985 (N_2985,N_755,N_312);
nand U2986 (N_2986,N_1040,N_246);
or U2987 (N_2987,N_1378,N_1445);
or U2988 (N_2988,N_54,N_72);
and U2989 (N_2989,N_62,N_682);
nand U2990 (N_2990,N_1317,N_1150);
and U2991 (N_2991,N_849,N_1181);
and U2992 (N_2992,N_202,N_1079);
nand U2993 (N_2993,N_390,N_898);
nand U2994 (N_2994,N_1073,N_128);
xor U2995 (N_2995,N_1046,N_759);
nand U2996 (N_2996,N_1480,N_1449);
and U2997 (N_2997,N_50,N_385);
and U2998 (N_2998,N_763,N_378);
nor U2999 (N_2999,N_296,N_584);
or U3000 (N_3000,N_1618,N_2270);
or U3001 (N_3001,N_2367,N_2194);
nor U3002 (N_3002,N_1927,N_2856);
xnor U3003 (N_3003,N_1870,N_2731);
and U3004 (N_3004,N_2206,N_2983);
nand U3005 (N_3005,N_2891,N_2583);
or U3006 (N_3006,N_2309,N_1982);
and U3007 (N_3007,N_2578,N_1955);
nand U3008 (N_3008,N_1680,N_1771);
nand U3009 (N_3009,N_1911,N_1905);
or U3010 (N_3010,N_1980,N_2709);
or U3011 (N_3011,N_1501,N_2223);
and U3012 (N_3012,N_2786,N_1882);
nor U3013 (N_3013,N_2712,N_1790);
and U3014 (N_3014,N_2002,N_1749);
or U3015 (N_3015,N_2326,N_2279);
nor U3016 (N_3016,N_2886,N_2796);
nor U3017 (N_3017,N_2657,N_1957);
nand U3018 (N_3018,N_1694,N_2242);
and U3019 (N_3019,N_1736,N_2869);
nor U3020 (N_3020,N_1699,N_2970);
nand U3021 (N_3021,N_2400,N_2409);
nor U3022 (N_3022,N_2445,N_2331);
or U3023 (N_3023,N_1880,N_2962);
and U3024 (N_3024,N_2902,N_2256);
or U3025 (N_3025,N_2939,N_1944);
and U3026 (N_3026,N_2757,N_2384);
nor U3027 (N_3027,N_2129,N_2503);
and U3028 (N_3028,N_2428,N_2297);
or U3029 (N_3029,N_2147,N_1634);
or U3030 (N_3030,N_2555,N_2673);
nor U3031 (N_3031,N_1938,N_1710);
xnor U3032 (N_3032,N_2986,N_1825);
and U3033 (N_3033,N_2062,N_2130);
or U3034 (N_3034,N_1846,N_2966);
and U3035 (N_3035,N_1620,N_2004);
nand U3036 (N_3036,N_2009,N_2292);
nand U3037 (N_3037,N_2680,N_1670);
and U3038 (N_3038,N_2416,N_2581);
xnor U3039 (N_3039,N_2879,N_2821);
nand U3040 (N_3040,N_1777,N_2267);
and U3041 (N_3041,N_1948,N_2815);
nand U3042 (N_3042,N_2105,N_2855);
nor U3043 (N_3043,N_2411,N_2064);
and U3044 (N_3044,N_2713,N_2807);
and U3045 (N_3045,N_1525,N_2412);
xnor U3046 (N_3046,N_2317,N_2823);
nand U3047 (N_3047,N_2133,N_2199);
and U3048 (N_3048,N_1586,N_1742);
nand U3049 (N_3049,N_1812,N_1807);
or U3050 (N_3050,N_2521,N_2429);
and U3051 (N_3051,N_2020,N_1619);
or U3052 (N_3052,N_2638,N_2539);
and U3053 (N_3053,N_2566,N_2554);
or U3054 (N_3054,N_2028,N_2979);
xnor U3055 (N_3055,N_1719,N_2775);
or U3056 (N_3056,N_1928,N_2865);
or U3057 (N_3057,N_2330,N_2904);
and U3058 (N_3058,N_2667,N_1843);
and U3059 (N_3059,N_2625,N_1998);
or U3060 (N_3060,N_2664,N_1939);
nand U3061 (N_3061,N_1861,N_2487);
nor U3062 (N_3062,N_2585,N_2965);
or U3063 (N_3063,N_1971,N_2284);
and U3064 (N_3064,N_2635,N_2361);
nand U3065 (N_3065,N_2588,N_1675);
or U3066 (N_3066,N_2721,N_2946);
or U3067 (N_3067,N_2640,N_1811);
nor U3068 (N_3068,N_2257,N_2321);
nor U3069 (N_3069,N_1916,N_2380);
nor U3070 (N_3070,N_2327,N_1612);
or U3071 (N_3071,N_2570,N_1746);
and U3072 (N_3072,N_1862,N_2463);
or U3073 (N_3073,N_2829,N_1655);
nand U3074 (N_3074,N_2055,N_1667);
and U3075 (N_3075,N_1588,N_1885);
and U3076 (N_3076,N_2510,N_2379);
xnor U3077 (N_3077,N_2508,N_1889);
nand U3078 (N_3078,N_2278,N_2870);
xnor U3079 (N_3079,N_1900,N_2750);
and U3080 (N_3080,N_1554,N_2915);
xor U3081 (N_3081,N_1651,N_2526);
xor U3082 (N_3082,N_2280,N_2112);
and U3083 (N_3083,N_2111,N_2711);
xnor U3084 (N_3084,N_2971,N_2740);
and U3085 (N_3085,N_2191,N_1839);
and U3086 (N_3086,N_2603,N_2652);
nand U3087 (N_3087,N_2698,N_2401);
and U3088 (N_3088,N_2138,N_2695);
nand U3089 (N_3089,N_2003,N_2747);
nand U3090 (N_3090,N_2114,N_1599);
and U3091 (N_3091,N_2837,N_1570);
nand U3092 (N_3092,N_2077,N_2476);
and U3093 (N_3093,N_2994,N_1520);
nor U3094 (N_3094,N_2039,N_2726);
or U3095 (N_3095,N_1813,N_2955);
or U3096 (N_3096,N_1726,N_2110);
or U3097 (N_3097,N_2972,N_1738);
or U3098 (N_3098,N_2057,N_2499);
nor U3099 (N_3099,N_2844,N_2387);
or U3100 (N_3100,N_2593,N_1737);
nor U3101 (N_3101,N_1616,N_1997);
nor U3102 (N_3102,N_2549,N_1921);
xnor U3103 (N_3103,N_1818,N_2885);
nor U3104 (N_3104,N_2440,N_2291);
nor U3105 (N_3105,N_2420,N_2614);
or U3106 (N_3106,N_1510,N_2218);
xor U3107 (N_3107,N_1578,N_1535);
and U3108 (N_3108,N_1996,N_2377);
or U3109 (N_3109,N_1933,N_1696);
or U3110 (N_3110,N_2683,N_2316);
nand U3111 (N_3111,N_2315,N_1931);
and U3112 (N_3112,N_1635,N_1942);
xnor U3113 (N_3113,N_2023,N_2107);
and U3114 (N_3114,N_1574,N_1781);
nor U3115 (N_3115,N_2090,N_1962);
nor U3116 (N_3116,N_2001,N_2532);
nor U3117 (N_3117,N_2505,N_2515);
nor U3118 (N_3118,N_1898,N_2557);
nand U3119 (N_3119,N_2442,N_1633);
and U3120 (N_3120,N_2386,N_2069);
nand U3121 (N_3121,N_2758,N_1621);
nand U3122 (N_3122,N_2804,N_2550);
or U3123 (N_3123,N_1592,N_2459);
nor U3124 (N_3124,N_2332,N_2745);
nor U3125 (N_3125,N_2137,N_2254);
nor U3126 (N_3126,N_2343,N_2708);
or U3127 (N_3127,N_1598,N_2392);
or U3128 (N_3128,N_2932,N_2417);
nor U3129 (N_3129,N_2150,N_2000);
and U3130 (N_3130,N_2849,N_2956);
and U3131 (N_3131,N_2875,N_2053);
or U3132 (N_3132,N_2688,N_2789);
or U3133 (N_3133,N_2471,N_1848);
and U3134 (N_3134,N_2957,N_2738);
or U3135 (N_3135,N_2120,N_2236);
nand U3136 (N_3136,N_1645,N_2960);
or U3137 (N_3137,N_1565,N_2093);
nor U3138 (N_3138,N_1557,N_2501);
or U3139 (N_3139,N_1528,N_1664);
xor U3140 (N_3140,N_1668,N_2220);
nand U3141 (N_3141,N_2852,N_1687);
nand U3142 (N_3142,N_1689,N_2959);
nand U3143 (N_3143,N_2743,N_1760);
xnor U3144 (N_3144,N_2142,N_2636);
or U3145 (N_3145,N_1561,N_2108);
and U3146 (N_3146,N_2214,N_2877);
or U3147 (N_3147,N_2397,N_1802);
xor U3148 (N_3148,N_1819,N_1963);
or U3149 (N_3149,N_1833,N_1556);
nand U3150 (N_3150,N_2669,N_2597);
or U3151 (N_3151,N_1759,N_1513);
and U3152 (N_3152,N_1608,N_2671);
nor U3153 (N_3153,N_2928,N_2851);
nand U3154 (N_3154,N_2990,N_2127);
or U3155 (N_3155,N_1748,N_2181);
nand U3156 (N_3156,N_1704,N_2826);
nor U3157 (N_3157,N_1823,N_2937);
and U3158 (N_3158,N_2500,N_2168);
nand U3159 (N_3159,N_1568,N_2564);
or U3160 (N_3160,N_2847,N_2352);
or U3161 (N_3161,N_2567,N_2224);
and U3162 (N_3162,N_1888,N_1897);
xnor U3163 (N_3163,N_2022,N_1653);
and U3164 (N_3164,N_1829,N_1896);
or U3165 (N_3165,N_1571,N_2616);
nand U3166 (N_3166,N_1991,N_1935);
xor U3167 (N_3167,N_2014,N_1787);
xnor U3168 (N_3168,N_2540,N_2774);
xnor U3169 (N_3169,N_2228,N_2430);
or U3170 (N_3170,N_2484,N_2854);
nand U3171 (N_3171,N_2996,N_2729);
and U3172 (N_3172,N_1851,N_1547);
nor U3173 (N_3173,N_2706,N_2453);
xnor U3174 (N_3174,N_1577,N_2702);
and U3175 (N_3175,N_2486,N_1709);
or U3176 (N_3176,N_2963,N_2272);
nor U3177 (N_3177,N_2897,N_2241);
or U3178 (N_3178,N_2227,N_1828);
or U3179 (N_3179,N_1590,N_1626);
nor U3180 (N_3180,N_2162,N_2719);
and U3181 (N_3181,N_2243,N_2630);
and U3182 (N_3182,N_2820,N_1611);
nor U3183 (N_3183,N_2303,N_2040);
and U3184 (N_3184,N_2883,N_2867);
or U3185 (N_3185,N_2180,N_1920);
nor U3186 (N_3186,N_1775,N_2917);
and U3187 (N_3187,N_2152,N_2969);
nor U3188 (N_3188,N_2030,N_1832);
nand U3189 (N_3189,N_1569,N_1683);
nor U3190 (N_3190,N_1863,N_1815);
nor U3191 (N_3191,N_2158,N_2460);
nand U3192 (N_3192,N_2761,N_2329);
xor U3193 (N_3193,N_2911,N_1617);
xnor U3194 (N_3194,N_1817,N_1659);
nor U3195 (N_3195,N_2368,N_2164);
or U3196 (N_3196,N_2863,N_2705);
nand U3197 (N_3197,N_2200,N_2827);
nor U3198 (N_3198,N_1529,N_2478);
nor U3199 (N_3199,N_2466,N_1684);
nand U3200 (N_3200,N_1702,N_1548);
nor U3201 (N_3201,N_2447,N_2776);
and U3202 (N_3202,N_1596,N_2251);
nor U3203 (N_3203,N_2798,N_2535);
or U3204 (N_3204,N_2506,N_2978);
and U3205 (N_3205,N_2454,N_1542);
xor U3206 (N_3206,N_1932,N_1890);
or U3207 (N_3207,N_1835,N_2682);
xnor U3208 (N_3208,N_1627,N_2339);
nand U3209 (N_3209,N_2139,N_2882);
nor U3210 (N_3210,N_1875,N_2300);
nand U3211 (N_3211,N_2922,N_2382);
nor U3212 (N_3212,N_2018,N_1808);
nand U3213 (N_3213,N_2259,N_2950);
nand U3214 (N_3214,N_2071,N_1572);
xnor U3215 (N_3215,N_2029,N_1720);
nand U3216 (N_3216,N_2253,N_2099);
or U3217 (N_3217,N_2514,N_1895);
and U3218 (N_3218,N_2903,N_1663);
nor U3219 (N_3219,N_2656,N_1614);
xnor U3220 (N_3220,N_1891,N_2086);
and U3221 (N_3221,N_2271,N_1526);
and U3222 (N_3222,N_1682,N_1541);
nor U3223 (N_3223,N_2073,N_2318);
nor U3224 (N_3224,N_2639,N_2311);
nand U3225 (N_3225,N_2948,N_1629);
and U3226 (N_3226,N_2225,N_2252);
and U3227 (N_3227,N_1551,N_1671);
nor U3228 (N_3228,N_1794,N_2104);
and U3229 (N_3229,N_2791,N_1773);
and U3230 (N_3230,N_1806,N_1822);
nor U3231 (N_3231,N_1532,N_1714);
or U3232 (N_3232,N_2308,N_2010);
or U3233 (N_3233,N_1909,N_2733);
nand U3234 (N_3234,N_2623,N_2208);
nor U3235 (N_3235,N_2952,N_1864);
nor U3236 (N_3236,N_2910,N_1638);
nor U3237 (N_3237,N_2624,N_1950);
nor U3238 (N_3238,N_1915,N_2350);
nand U3239 (N_3239,N_2295,N_2131);
xor U3240 (N_3240,N_2480,N_2860);
or U3241 (N_3241,N_2780,N_2488);
nand U3242 (N_3242,N_2103,N_2998);
and U3243 (N_3243,N_2472,N_1881);
nand U3244 (N_3244,N_1508,N_1757);
nand U3245 (N_3245,N_1706,N_2646);
nor U3246 (N_3246,N_2078,N_2779);
nand U3247 (N_3247,N_2600,N_2833);
and U3248 (N_3248,N_2470,N_2919);
nand U3249 (N_3249,N_2146,N_2545);
and U3250 (N_3250,N_2958,N_1867);
or U3251 (N_3251,N_1566,N_2007);
nor U3252 (N_3252,N_2404,N_1511);
or U3253 (N_3253,N_2628,N_1856);
nor U3254 (N_3254,N_2684,N_2128);
and U3255 (N_3255,N_2770,N_1560);
or U3256 (N_3256,N_2511,N_1770);
and U3257 (N_3257,N_2512,N_2362);
nor U3258 (N_3258,N_2677,N_1695);
or U3259 (N_3259,N_2642,N_2755);
and U3260 (N_3260,N_2670,N_2301);
xnor U3261 (N_3261,N_2398,N_2230);
or U3262 (N_3262,N_2405,N_2687);
nor U3263 (N_3263,N_2898,N_2661);
nand U3264 (N_3264,N_1879,N_2734);
and U3265 (N_3265,N_1868,N_1892);
nand U3266 (N_3266,N_1647,N_2756);
nor U3267 (N_3267,N_2519,N_1562);
and U3268 (N_3268,N_2644,N_2172);
or U3269 (N_3269,N_2634,N_2226);
nor U3270 (N_3270,N_2161,N_1966);
nor U3271 (N_3271,N_2772,N_2801);
nand U3272 (N_3272,N_2452,N_2042);
nand U3273 (N_3273,N_2536,N_2675);
and U3274 (N_3274,N_1721,N_1857);
xor U3275 (N_3275,N_2619,N_1594);
or U3276 (N_3276,N_1643,N_2313);
nand U3277 (N_3277,N_2989,N_1923);
nand U3278 (N_3278,N_2370,N_1537);
xnor U3279 (N_3279,N_2446,N_1953);
and U3280 (N_3280,N_2117,N_2806);
nor U3281 (N_3281,N_1949,N_2373);
nand U3282 (N_3282,N_1826,N_2560);
or U3283 (N_3283,N_2151,N_2249);
xnor U3284 (N_3284,N_1536,N_1874);
nor U3285 (N_3285,N_2627,N_1549);
nor U3286 (N_3286,N_2631,N_2461);
nand U3287 (N_3287,N_2838,N_2097);
nor U3288 (N_3288,N_2534,N_1965);
and U3289 (N_3289,N_2795,N_2113);
or U3290 (N_3290,N_2074,N_2765);
and U3291 (N_3291,N_1740,N_2144);
and U3292 (N_3292,N_1673,N_2169);
and U3293 (N_3293,N_1576,N_1834);
xor U3294 (N_3294,N_2509,N_1941);
nand U3295 (N_3295,N_2633,N_1649);
or U3296 (N_3296,N_2759,N_1984);
xnor U3297 (N_3297,N_2424,N_2828);
or U3298 (N_3298,N_1713,N_2265);
xor U3299 (N_3299,N_2234,N_2914);
or U3300 (N_3300,N_2418,N_2155);
and U3301 (N_3301,N_2122,N_1735);
and U3302 (N_3302,N_1968,N_1503);
or U3303 (N_3303,N_1934,N_1956);
nor U3304 (N_3304,N_2075,N_2217);
or U3305 (N_3305,N_2027,N_1518);
and U3306 (N_3306,N_1601,N_1550);
nor U3307 (N_3307,N_2887,N_1575);
xor U3308 (N_3308,N_2654,N_2021);
nand U3309 (N_3309,N_1899,N_1539);
and U3310 (N_3310,N_2703,N_2982);
or U3311 (N_3311,N_1609,N_1803);
nor U3312 (N_3312,N_2612,N_2929);
nand U3313 (N_3313,N_2666,N_1747);
and U3314 (N_3314,N_2338,N_2035);
xnor U3315 (N_3315,N_2717,N_2561);
nor U3316 (N_3316,N_2866,N_2668);
nand U3317 (N_3317,N_2413,N_2651);
nor U3318 (N_3318,N_1733,N_1852);
nand U3319 (N_3319,N_1821,N_1715);
nand U3320 (N_3320,N_2571,N_1782);
nand U3321 (N_3321,N_1688,N_2337);
or U3322 (N_3322,N_1869,N_1585);
nor U3323 (N_3323,N_2354,N_1724);
and U3324 (N_3324,N_2991,N_2741);
nor U3325 (N_3325,N_1778,N_2813);
and U3326 (N_3326,N_2809,N_2876);
or U3327 (N_3327,N_2601,N_2394);
nand U3328 (N_3328,N_1661,N_1691);
nand U3329 (N_3329,N_1504,N_1700);
nand U3330 (N_3330,N_1761,N_1669);
or U3331 (N_3331,N_2559,N_1660);
and U3332 (N_3332,N_2543,N_1768);
xor U3333 (N_3333,N_1959,N_1693);
or U3334 (N_3334,N_2448,N_2115);
nand U3335 (N_3335,N_2662,N_2558);
or U3336 (N_3336,N_2482,N_2552);
nand U3337 (N_3337,N_2930,N_2961);
and U3338 (N_3338,N_1774,N_2212);
xor U3339 (N_3339,N_2530,N_2419);
or U3340 (N_3340,N_2988,N_1951);
and U3341 (N_3341,N_2525,N_1628);
nand U3342 (N_3342,N_2153,N_2762);
nor U3343 (N_3343,N_2195,N_2921);
xor U3344 (N_3344,N_2736,N_1922);
and U3345 (N_3345,N_1679,N_1564);
and U3346 (N_3346,N_1717,N_1583);
and U3347 (N_3347,N_2551,N_2784);
nor U3348 (N_3348,N_1810,N_1917);
and U3349 (N_3349,N_2553,N_2371);
or U3350 (N_3350,N_2589,N_1772);
or U3351 (N_3351,N_1908,N_2310);
nand U3352 (N_3352,N_2328,N_2546);
nand U3353 (N_3353,N_2766,N_1697);
and U3354 (N_3354,N_2451,N_2993);
or U3355 (N_3355,N_2443,N_1506);
nor U3356 (N_3356,N_2365,N_2647);
or U3357 (N_3357,N_2274,N_1716);
nor U3358 (N_3358,N_2095,N_2954);
and U3359 (N_3359,N_2210,N_2247);
nand U3360 (N_3360,N_1558,N_1622);
and U3361 (N_3361,N_1707,N_2598);
nor U3362 (N_3362,N_1745,N_2066);
nand U3363 (N_3363,N_2154,N_2385);
or U3364 (N_3364,N_2528,N_2781);
nor U3365 (N_3365,N_2285,N_1866);
and U3366 (N_3366,N_1589,N_1855);
nand U3367 (N_3367,N_2043,N_2892);
and U3368 (N_3368,N_2562,N_1906);
or U3369 (N_3369,N_2728,N_2531);
xor U3370 (N_3370,N_2319,N_2984);
nand U3371 (N_3371,N_1854,N_2611);
xnor U3372 (N_3372,N_2678,N_1860);
nor U3373 (N_3373,N_2016,N_2768);
xor U3374 (N_3374,N_2699,N_2473);
and U3375 (N_3375,N_1902,N_1553);
or U3376 (N_3376,N_2685,N_1952);
or U3377 (N_3377,N_2034,N_2606);
or U3378 (N_3378,N_2302,N_1958);
nand U3379 (N_3379,N_1545,N_1750);
and U3380 (N_3380,N_1995,N_1657);
nand U3381 (N_3381,N_2835,N_2977);
xnor U3382 (N_3382,N_2579,N_2931);
nand U3383 (N_3383,N_2193,N_1850);
nand U3384 (N_3384,N_2026,N_1989);
and U3385 (N_3385,N_1582,N_1840);
or U3386 (N_3386,N_1783,N_2934);
nor U3387 (N_3387,N_2175,N_1692);
xor U3388 (N_3388,N_2692,N_1799);
nor U3389 (N_3389,N_2165,N_2818);
nor U3390 (N_3390,N_2156,N_2832);
nand U3391 (N_3391,N_2576,N_2788);
xnor U3392 (N_3392,N_1637,N_2502);
and U3393 (N_3393,N_1701,N_2622);
nor U3394 (N_3394,N_1816,N_2602);
nor U3395 (N_3395,N_2490,N_2314);
nand U3396 (N_3396,N_2215,N_1983);
and U3397 (N_3397,N_2495,N_2198);
and U3398 (N_3398,N_2785,N_2858);
and U3399 (N_3399,N_2477,N_2693);
nor U3400 (N_3400,N_2873,N_2229);
and U3401 (N_3401,N_1780,N_1521);
nor U3402 (N_3402,N_2083,N_2202);
and U3403 (N_3403,N_1784,N_2565);
nand U3404 (N_3404,N_2645,N_2469);
and U3405 (N_3405,N_2237,N_2933);
or U3406 (N_3406,N_1753,N_1625);
or U3407 (N_3407,N_2938,N_2032);
nor U3408 (N_3408,N_2076,N_1978);
and U3409 (N_3409,N_2596,N_1741);
or U3410 (N_3410,N_2305,N_2658);
nand U3411 (N_3411,N_2805,N_2935);
nand U3412 (N_3412,N_1903,N_1992);
or U3413 (N_3413,N_1672,N_1734);
nand U3414 (N_3414,N_2947,N_2081);
nand U3415 (N_3415,N_2100,N_1804);
or U3416 (N_3416,N_2132,N_2749);
xor U3417 (N_3417,N_1930,N_1827);
nand U3418 (N_3418,N_2594,N_1678);
or U3419 (N_3419,N_2307,N_1555);
and U3420 (N_3420,N_1936,N_2348);
xnor U3421 (N_3421,N_2790,N_2171);
xnor U3422 (N_3422,N_2383,N_2008);
nand U3423 (N_3423,N_2894,N_1722);
nor U3424 (N_3424,N_2590,N_2290);
nand U3425 (N_3425,N_1987,N_2219);
or U3426 (N_3426,N_2462,N_2696);
nor U3427 (N_3427,N_2408,N_1584);
nor U3428 (N_3428,N_2414,N_1544);
and U3429 (N_3429,N_1615,N_1876);
nand U3430 (N_3430,N_1604,N_2455);
nand U3431 (N_3431,N_2556,N_2334);
and U3432 (N_3432,N_2769,N_1509);
or U3433 (N_3433,N_2068,N_2739);
and U3434 (N_3434,N_2389,N_1972);
or U3435 (N_3435,N_1849,N_2817);
nor U3436 (N_3436,N_1837,N_1805);
nand U3437 (N_3437,N_1648,N_1602);
xnor U3438 (N_3438,N_1919,N_2893);
xnor U3439 (N_3439,N_1865,N_2239);
or U3440 (N_3440,N_2190,N_2494);
and U3441 (N_3441,N_1797,N_2822);
or U3442 (N_3442,N_1563,N_2800);
nor U3443 (N_3443,N_2116,N_2691);
and U3444 (N_3444,N_2799,N_2906);
nor U3445 (N_3445,N_1641,N_2676);
nor U3446 (N_3446,N_1642,N_2126);
nand U3447 (N_3447,N_2613,N_2672);
or U3448 (N_3448,N_1725,N_2197);
nor U3449 (N_3449,N_2096,N_2572);
xor U3450 (N_3450,N_2087,N_1603);
nor U3451 (N_3451,N_1779,N_2140);
xnor U3452 (N_3452,N_2773,N_2450);
xnor U3453 (N_3453,N_1727,N_1765);
nor U3454 (N_3454,N_1674,N_1698);
nor U3455 (N_3455,N_1685,N_2192);
or U3456 (N_3456,N_2433,N_1690);
nor U3457 (N_3457,N_2841,N_1636);
or U3458 (N_3458,N_2595,N_2909);
nand U3459 (N_3459,N_2046,N_2372);
or U3460 (N_3460,N_2293,N_2632);
nand U3461 (N_3461,N_1976,N_1606);
nor U3462 (N_3462,N_2746,N_2872);
xnor U3463 (N_3463,N_2880,N_2378);
nor U3464 (N_3464,N_2432,N_2084);
nand U3465 (N_3465,N_1907,N_1686);
nand U3466 (N_3466,N_2723,N_2563);
nand U3467 (N_3467,N_2124,N_2533);
and U3468 (N_3468,N_2347,N_2045);
nor U3469 (N_3469,N_2051,N_1795);
nand U3470 (N_3470,N_1587,N_2707);
and U3471 (N_3471,N_1666,N_2504);
and U3472 (N_3472,N_2255,N_2065);
or U3473 (N_3473,N_2067,N_1792);
and U3474 (N_3474,N_2541,N_2831);
or U3475 (N_3475,N_2012,N_2336);
and U3476 (N_3476,N_1994,N_2346);
nor U3477 (N_3477,N_1912,N_2846);
nor U3478 (N_3478,N_2052,N_2054);
and U3479 (N_3479,N_2771,N_2975);
nand U3480 (N_3480,N_2125,N_2744);
nor U3481 (N_3481,N_2943,N_2735);
nor U3482 (N_3482,N_2592,N_2643);
nand U3483 (N_3483,N_2088,N_2423);
xor U3484 (N_3484,N_2686,N_1801);
or U3485 (N_3485,N_2918,N_2940);
and U3486 (N_3486,N_2663,N_1744);
nand U3487 (N_3487,N_2390,N_2655);
nand U3488 (N_3488,N_2752,N_1524);
nand U3489 (N_3489,N_1538,N_2748);
and U3490 (N_3490,N_1961,N_2174);
nor U3491 (N_3491,N_2196,N_2182);
and U3492 (N_3492,N_2610,N_1877);
or U3493 (N_3493,N_1523,N_2778);
and U3494 (N_3494,N_2276,N_2092);
and U3495 (N_3495,N_2340,N_1986);
or U3496 (N_3496,N_1591,N_1540);
nor U3497 (N_3497,N_1798,N_2923);
and U3498 (N_3498,N_1945,N_2840);
xnor U3499 (N_3499,N_2522,N_1796);
nand U3500 (N_3500,N_2186,N_2288);
and U3501 (N_3501,N_2715,N_2575);
nand U3502 (N_3502,N_2080,N_2015);
and U3503 (N_3503,N_2577,N_2964);
nor U3504 (N_3504,N_2421,N_2238);
or U3505 (N_3505,N_1677,N_2005);
and U3506 (N_3506,N_2465,N_1527);
nand U3507 (N_3507,N_1559,N_1530);
nand U3508 (N_3508,N_2282,N_2987);
nor U3509 (N_3509,N_2437,N_2233);
nor U3510 (N_3510,N_2263,N_1516);
nand U3511 (N_3511,N_2159,N_2245);
and U3512 (N_3512,N_2679,N_1739);
and U3513 (N_3513,N_2407,N_2584);
nand U3514 (N_3514,N_2369,N_2542);
nand U3515 (N_3515,N_2942,N_1990);
or U3516 (N_3516,N_2425,N_1999);
and U3517 (N_3517,N_1593,N_2358);
nand U3518 (N_3518,N_2041,N_1533);
and U3519 (N_3519,N_1820,N_2608);
nor U3520 (N_3520,N_2845,N_2905);
nand U3521 (N_3521,N_1567,N_2901);
xnor U3522 (N_3522,N_1831,N_1718);
nor U3523 (N_3523,N_2363,N_2250);
nand U3524 (N_3524,N_2615,N_2261);
or U3525 (N_3525,N_2763,N_1988);
xor U3526 (N_3526,N_2205,N_2006);
and U3527 (N_3527,N_2091,N_2836);
and U3528 (N_3528,N_2518,N_1873);
nand U3529 (N_3529,N_2058,N_2496);
or U3530 (N_3530,N_2374,N_1979);
nor U3531 (N_3531,N_2173,N_1607);
xnor U3532 (N_3532,N_2925,N_1964);
nor U3533 (N_3533,N_2900,N_2388);
and U3534 (N_3534,N_1600,N_1893);
nor U3535 (N_3535,N_2294,N_1573);
nand U3536 (N_3536,N_1977,N_1512);
nand U3537 (N_3537,N_2277,N_2121);
or U3538 (N_3538,N_2185,N_2949);
nand U3539 (N_3539,N_2232,N_2497);
nor U3540 (N_3540,N_1845,N_2751);
nor U3541 (N_3541,N_1762,N_2483);
nor U3542 (N_3542,N_1729,N_2629);
or U3543 (N_3543,N_1776,N_1764);
nor U3544 (N_3544,N_2427,N_2710);
or U3545 (N_3545,N_2816,N_2246);
or U3546 (N_3546,N_2941,N_2649);
or U3547 (N_3547,N_2620,N_2356);
or U3548 (N_3548,N_2722,N_1894);
or U3549 (N_3549,N_2357,N_2697);
and U3550 (N_3550,N_1711,N_2479);
or U3551 (N_3551,N_2997,N_2410);
nand U3552 (N_3552,N_2529,N_2730);
or U3553 (N_3553,N_1904,N_2013);
or U3554 (N_3554,N_2268,N_2980);
and U3555 (N_3555,N_1640,N_2626);
or U3556 (N_3556,N_1960,N_2402);
and U3557 (N_3557,N_2258,N_2936);
and U3558 (N_3558,N_1858,N_2689);
nand U3559 (N_3559,N_2782,N_2767);
nand U3560 (N_3560,N_2580,N_2393);
nor U3561 (N_3561,N_2777,N_1519);
nand U3562 (N_3562,N_2913,N_1853);
and U3563 (N_3563,N_2351,N_1723);
nor U3564 (N_3564,N_2884,N_1924);
nor U3565 (N_3565,N_2439,N_1836);
or U3566 (N_3566,N_2375,N_2260);
and U3567 (N_3567,N_1652,N_2825);
nor U3568 (N_3568,N_2742,N_2641);
nor U3569 (N_3569,N_2498,N_2916);
xnor U3570 (N_3570,N_2468,N_2797);
nor U3571 (N_3571,N_2353,N_2814);
and U3572 (N_3572,N_2718,N_2184);
nand U3573 (N_3573,N_2912,N_2716);
nor U3574 (N_3574,N_2537,N_2783);
nor U3575 (N_3575,N_2431,N_2527);
nand U3576 (N_3576,N_1755,N_2187);
or U3577 (N_3577,N_2240,N_2135);
xnor U3578 (N_3578,N_1767,N_1656);
nor U3579 (N_3579,N_2467,N_2060);
xnor U3580 (N_3580,N_2434,N_1597);
xnor U3581 (N_3581,N_2166,N_1517);
or U3582 (N_3582,N_2170,N_2209);
nor U3583 (N_3583,N_2896,N_2281);
and U3584 (N_3584,N_2102,N_1728);
and U3585 (N_3585,N_2048,N_2059);
nand U3586 (N_3586,N_2216,N_1754);
and U3587 (N_3587,N_2618,N_1993);
xnor U3588 (N_3588,N_2038,N_1859);
or U3589 (N_3589,N_1844,N_2148);
or U3590 (N_3590,N_2458,N_1841);
or U3591 (N_3591,N_2399,N_2296);
or U3592 (N_3592,N_2793,N_1732);
nand U3593 (N_3593,N_2136,N_2507);
nand U3594 (N_3594,N_2160,N_2544);
or U3595 (N_3595,N_2167,N_2235);
nand U3596 (N_3596,N_2422,N_1743);
nor U3597 (N_3597,N_1676,N_2665);
and U3598 (N_3598,N_1763,N_2701);
nand U3599 (N_3599,N_2704,N_2681);
nand U3600 (N_3600,N_2079,N_2438);
or U3601 (N_3601,N_2953,N_1624);
xor U3602 (N_3602,N_1824,N_1981);
nand U3603 (N_3603,N_1901,N_1946);
or U3604 (N_3604,N_2920,N_2406);
or U3605 (N_3605,N_2044,N_2819);
nor U3606 (N_3606,N_2737,N_2538);
nor U3607 (N_3607,N_2441,N_2927);
and U3608 (N_3608,N_2492,N_2082);
nor U3609 (N_3609,N_2868,N_2725);
or U3610 (N_3610,N_2275,N_2548);
nand U3611 (N_3611,N_2201,N_1552);
nor U3612 (N_3612,N_1646,N_2951);
nand U3613 (N_3613,N_1752,N_1886);
or U3614 (N_3614,N_1631,N_1947);
xnor U3615 (N_3615,N_2335,N_2207);
nor U3616 (N_3616,N_2436,N_1758);
xor U3617 (N_3617,N_2811,N_2907);
or U3618 (N_3618,N_1662,N_2485);
and U3619 (N_3619,N_1500,N_2178);
nor U3620 (N_3620,N_2475,N_1883);
or U3621 (N_3621,N_2049,N_2266);
nand U3622 (N_3622,N_2342,N_1788);
nor U3623 (N_3623,N_1929,N_1665);
nand U3624 (N_3624,N_2037,N_2724);
xnor U3625 (N_3625,N_2320,N_1632);
and U3626 (N_3626,N_2690,N_2322);
and U3627 (N_3627,N_2714,N_1630);
or U3628 (N_3628,N_2569,N_2070);
and U3629 (N_3629,N_2853,N_2349);
or U3630 (N_3630,N_1531,N_2824);
xnor U3631 (N_3631,N_2609,N_2449);
or U3632 (N_3632,N_2481,N_2637);
nand U3633 (N_3633,N_1878,N_2648);
nor U3634 (N_3634,N_2244,N_1580);
xnor U3635 (N_3635,N_2025,N_1605);
xnor U3636 (N_3636,N_1708,N_1830);
nand U3637 (N_3637,N_2426,N_2812);
or U3638 (N_3638,N_1967,N_2992);
and U3639 (N_3639,N_2842,N_1793);
nor U3640 (N_3640,N_2574,N_2848);
nand U3641 (N_3641,N_1943,N_2926);
nand U3642 (N_3642,N_2444,N_1756);
nor U3643 (N_3643,N_2976,N_2061);
nand U3644 (N_3644,N_2547,N_2861);
nand U3645 (N_3645,N_1639,N_2345);
and U3646 (N_3646,N_2360,N_2456);
nand U3647 (N_3647,N_2188,N_2211);
xnor U3648 (N_3648,N_1751,N_1515);
nor U3649 (N_3649,N_2094,N_2333);
xnor U3650 (N_3650,N_2273,N_2999);
or U3651 (N_3651,N_1789,N_1791);
nor U3652 (N_3652,N_2366,N_2944);
nand U3653 (N_3653,N_2024,N_2464);
xor U3654 (N_3654,N_2810,N_2085);
or U3655 (N_3655,N_2568,N_2031);
nor U3656 (N_3656,N_2888,N_1623);
nor U3657 (N_3657,N_1914,N_1872);
nand U3658 (N_3658,N_2491,N_1613);
nor U3659 (N_3659,N_2204,N_1884);
and U3660 (N_3660,N_2019,N_2203);
nand U3661 (N_3661,N_2050,N_2968);
and U3662 (N_3662,N_2700,N_2262);
nor U3663 (N_3663,N_1766,N_2299);
nand U3664 (N_3664,N_2889,N_1507);
or U3665 (N_3665,N_2857,N_2324);
nand U3666 (N_3666,N_2047,N_2248);
nand U3667 (N_3667,N_2298,N_2304);
nor U3668 (N_3668,N_2231,N_2808);
or U3669 (N_3669,N_2359,N_2839);
nor U3670 (N_3670,N_1918,N_2415);
nand U3671 (N_3671,N_2862,N_1681);
nand U3672 (N_3672,N_2489,N_2607);
and U3673 (N_3673,N_2653,N_1658);
nor U3674 (N_3674,N_2118,N_2396);
and U3675 (N_3675,N_2787,N_1534);
nand U3676 (N_3676,N_1937,N_1730);
or U3677 (N_3677,N_2179,N_1975);
nor U3678 (N_3678,N_1809,N_2843);
nand U3679 (N_3679,N_2222,N_2134);
and U3680 (N_3680,N_2011,N_2995);
nor U3681 (N_3681,N_1926,N_2283);
nor U3682 (N_3682,N_2376,N_2355);
nand U3683 (N_3683,N_2605,N_2794);
nor U3684 (N_3684,N_1814,N_2106);
and U3685 (N_3685,N_1973,N_2881);
and U3686 (N_3686,N_2694,N_2157);
and U3687 (N_3687,N_1940,N_2650);
and U3688 (N_3688,N_2753,N_1925);
or U3689 (N_3689,N_2973,N_2899);
and U3690 (N_3690,N_1974,N_2189);
and U3691 (N_3691,N_1650,N_2063);
nor U3692 (N_3692,N_2878,N_1800);
or U3693 (N_3693,N_2764,N_2306);
xor U3694 (N_3694,N_1514,N_2591);
nor U3695 (N_3695,N_1546,N_1785);
or U3696 (N_3696,N_2732,N_2802);
nor U3697 (N_3697,N_2513,N_2727);
nand U3698 (N_3698,N_1954,N_2072);
and U3699 (N_3699,N_2754,N_2341);
xor U3700 (N_3700,N_2524,N_2163);
or U3701 (N_3701,N_2177,N_1581);
or U3702 (N_3702,N_1910,N_1543);
nor U3703 (N_3703,N_2874,N_1610);
nor U3704 (N_3704,N_1502,N_2098);
nor U3705 (N_3705,N_1969,N_2517);
xnor U3706 (N_3706,N_2967,N_1842);
nor U3707 (N_3707,N_1731,N_2573);
and U3708 (N_3708,N_2523,N_2325);
nand U3709 (N_3709,N_2149,N_2109);
nor U3710 (N_3710,N_2850,N_2289);
or U3711 (N_3711,N_2056,N_2760);
nand U3712 (N_3712,N_2660,N_2143);
and U3713 (N_3713,N_2435,N_1505);
or U3714 (N_3714,N_2895,N_2803);
or U3715 (N_3715,N_2312,N_2017);
or U3716 (N_3716,N_2621,N_1654);
nor U3717 (N_3717,N_2792,N_2145);
or U3718 (N_3718,N_2286,N_2587);
nand U3719 (N_3719,N_2582,N_2493);
and U3720 (N_3720,N_1595,N_2981);
nor U3721 (N_3721,N_1913,N_1522);
and U3722 (N_3722,N_1887,N_2036);
and U3723 (N_3723,N_2344,N_2586);
nand U3724 (N_3724,N_2221,N_2381);
or U3725 (N_3725,N_2974,N_2864);
nor U3726 (N_3726,N_2659,N_2520);
nor U3727 (N_3727,N_1712,N_1644);
xor U3728 (N_3728,N_2457,N_2033);
nand U3729 (N_3729,N_2985,N_2830);
or U3730 (N_3730,N_2924,N_2123);
nor U3731 (N_3731,N_2395,N_2364);
or U3732 (N_3732,N_2720,N_1970);
nand U3733 (N_3733,N_2141,N_2264);
or U3734 (N_3734,N_2516,N_2119);
nand U3735 (N_3735,N_2183,N_1705);
xor U3736 (N_3736,N_1871,N_2474);
nand U3737 (N_3737,N_2599,N_2269);
nor U3738 (N_3738,N_2859,N_2908);
nor U3739 (N_3739,N_2403,N_2287);
xor U3740 (N_3740,N_2213,N_1838);
nor U3741 (N_3741,N_2871,N_1786);
nand U3742 (N_3742,N_1985,N_1703);
nor U3743 (N_3743,N_2617,N_1579);
xor U3744 (N_3744,N_2834,N_1847);
nand U3745 (N_3745,N_2674,N_2945);
and U3746 (N_3746,N_2176,N_2890);
nand U3747 (N_3747,N_2604,N_2089);
and U3748 (N_3748,N_1769,N_2101);
nor U3749 (N_3749,N_2323,N_2391);
xor U3750 (N_3750,N_2794,N_2830);
nand U3751 (N_3751,N_2847,N_2706);
nand U3752 (N_3752,N_2180,N_2909);
nand U3753 (N_3753,N_2938,N_1788);
or U3754 (N_3754,N_1643,N_2683);
or U3755 (N_3755,N_2202,N_2912);
and U3756 (N_3756,N_2161,N_2827);
or U3757 (N_3757,N_2037,N_2486);
or U3758 (N_3758,N_2165,N_2864);
nand U3759 (N_3759,N_2734,N_2939);
nand U3760 (N_3760,N_2748,N_1992);
or U3761 (N_3761,N_1873,N_2626);
xnor U3762 (N_3762,N_2233,N_1827);
nor U3763 (N_3763,N_1784,N_2316);
and U3764 (N_3764,N_1982,N_2154);
or U3765 (N_3765,N_2451,N_2567);
nor U3766 (N_3766,N_2088,N_2534);
nand U3767 (N_3767,N_2555,N_1521);
nor U3768 (N_3768,N_1745,N_1869);
and U3769 (N_3769,N_2698,N_2907);
nor U3770 (N_3770,N_2787,N_2864);
nand U3771 (N_3771,N_1771,N_2637);
and U3772 (N_3772,N_1905,N_2700);
and U3773 (N_3773,N_1557,N_2702);
and U3774 (N_3774,N_2185,N_1951);
nor U3775 (N_3775,N_1595,N_2304);
or U3776 (N_3776,N_2913,N_1885);
or U3777 (N_3777,N_2524,N_1995);
nor U3778 (N_3778,N_2758,N_1558);
nand U3779 (N_3779,N_2032,N_1758);
nand U3780 (N_3780,N_2847,N_1596);
and U3781 (N_3781,N_2517,N_2471);
and U3782 (N_3782,N_2428,N_2339);
nand U3783 (N_3783,N_1927,N_2955);
nor U3784 (N_3784,N_2549,N_1859);
nor U3785 (N_3785,N_2420,N_1722);
xor U3786 (N_3786,N_2158,N_2559);
nand U3787 (N_3787,N_2371,N_2082);
or U3788 (N_3788,N_1538,N_2353);
nand U3789 (N_3789,N_2642,N_2232);
nor U3790 (N_3790,N_1919,N_1738);
and U3791 (N_3791,N_2990,N_2001);
nand U3792 (N_3792,N_1635,N_1979);
nand U3793 (N_3793,N_2021,N_2369);
or U3794 (N_3794,N_2704,N_2903);
nand U3795 (N_3795,N_2344,N_2395);
xor U3796 (N_3796,N_2717,N_2111);
and U3797 (N_3797,N_2198,N_2500);
nand U3798 (N_3798,N_1520,N_2443);
nand U3799 (N_3799,N_1990,N_2144);
nand U3800 (N_3800,N_2876,N_1653);
xor U3801 (N_3801,N_1983,N_2755);
nand U3802 (N_3802,N_2431,N_2408);
nand U3803 (N_3803,N_2939,N_2995);
nor U3804 (N_3804,N_1720,N_1840);
nand U3805 (N_3805,N_2535,N_2208);
nor U3806 (N_3806,N_2061,N_2562);
and U3807 (N_3807,N_2702,N_2650);
nor U3808 (N_3808,N_2707,N_1807);
and U3809 (N_3809,N_2047,N_1581);
nand U3810 (N_3810,N_1542,N_2195);
or U3811 (N_3811,N_2276,N_2857);
nand U3812 (N_3812,N_2398,N_1650);
nand U3813 (N_3813,N_2949,N_1718);
nand U3814 (N_3814,N_2897,N_2239);
xnor U3815 (N_3815,N_2178,N_1929);
nand U3816 (N_3816,N_1704,N_2409);
or U3817 (N_3817,N_2128,N_2446);
and U3818 (N_3818,N_2600,N_1759);
and U3819 (N_3819,N_1992,N_1773);
and U3820 (N_3820,N_2001,N_1539);
xor U3821 (N_3821,N_2245,N_2874);
nor U3822 (N_3822,N_2831,N_2648);
or U3823 (N_3823,N_1942,N_1965);
nor U3824 (N_3824,N_2683,N_2381);
and U3825 (N_3825,N_2544,N_2442);
or U3826 (N_3826,N_2352,N_2295);
nand U3827 (N_3827,N_2352,N_2966);
nor U3828 (N_3828,N_2665,N_2410);
nand U3829 (N_3829,N_2639,N_2270);
nor U3830 (N_3830,N_2491,N_1676);
and U3831 (N_3831,N_2888,N_2856);
nand U3832 (N_3832,N_2098,N_2659);
nor U3833 (N_3833,N_1866,N_1649);
nand U3834 (N_3834,N_1528,N_1583);
nor U3835 (N_3835,N_2886,N_2531);
or U3836 (N_3836,N_2012,N_2145);
nor U3837 (N_3837,N_2782,N_2257);
or U3838 (N_3838,N_1999,N_2706);
nor U3839 (N_3839,N_2578,N_2236);
nand U3840 (N_3840,N_1892,N_1910);
nand U3841 (N_3841,N_1823,N_2403);
nor U3842 (N_3842,N_1925,N_2524);
or U3843 (N_3843,N_1790,N_2677);
nand U3844 (N_3844,N_2693,N_2465);
nand U3845 (N_3845,N_2352,N_2357);
nand U3846 (N_3846,N_1654,N_1988);
or U3847 (N_3847,N_2781,N_2676);
nor U3848 (N_3848,N_2210,N_1726);
nand U3849 (N_3849,N_1603,N_2002);
nand U3850 (N_3850,N_2944,N_2656);
and U3851 (N_3851,N_2535,N_2147);
or U3852 (N_3852,N_2292,N_1635);
nand U3853 (N_3853,N_2399,N_2962);
nand U3854 (N_3854,N_1731,N_2225);
nor U3855 (N_3855,N_2544,N_1987);
or U3856 (N_3856,N_2100,N_1882);
nor U3857 (N_3857,N_1946,N_2447);
and U3858 (N_3858,N_1507,N_1664);
nand U3859 (N_3859,N_1538,N_1696);
or U3860 (N_3860,N_2011,N_1891);
or U3861 (N_3861,N_2906,N_1982);
nor U3862 (N_3862,N_2001,N_1773);
xnor U3863 (N_3863,N_2090,N_2913);
nand U3864 (N_3864,N_2949,N_1534);
or U3865 (N_3865,N_2476,N_2373);
xor U3866 (N_3866,N_2953,N_2456);
nor U3867 (N_3867,N_2357,N_2422);
nand U3868 (N_3868,N_1761,N_2234);
or U3869 (N_3869,N_2224,N_1755);
and U3870 (N_3870,N_1955,N_2654);
nor U3871 (N_3871,N_2493,N_2734);
nor U3872 (N_3872,N_2204,N_1789);
and U3873 (N_3873,N_1762,N_1943);
or U3874 (N_3874,N_1901,N_2565);
or U3875 (N_3875,N_2355,N_2186);
or U3876 (N_3876,N_2144,N_2646);
and U3877 (N_3877,N_2897,N_2801);
nand U3878 (N_3878,N_2846,N_2094);
nand U3879 (N_3879,N_2638,N_2108);
nor U3880 (N_3880,N_2524,N_2723);
and U3881 (N_3881,N_2606,N_1539);
and U3882 (N_3882,N_1688,N_1789);
or U3883 (N_3883,N_2921,N_1967);
or U3884 (N_3884,N_1889,N_2732);
and U3885 (N_3885,N_2064,N_1972);
nor U3886 (N_3886,N_2336,N_2597);
and U3887 (N_3887,N_2799,N_2682);
nand U3888 (N_3888,N_2715,N_1564);
nor U3889 (N_3889,N_2142,N_2159);
nor U3890 (N_3890,N_2300,N_1755);
nor U3891 (N_3891,N_2450,N_2683);
or U3892 (N_3892,N_1603,N_2316);
or U3893 (N_3893,N_2251,N_1711);
xnor U3894 (N_3894,N_2023,N_1633);
or U3895 (N_3895,N_2083,N_2479);
nand U3896 (N_3896,N_1982,N_2615);
and U3897 (N_3897,N_2571,N_2450);
and U3898 (N_3898,N_1949,N_2360);
nor U3899 (N_3899,N_2155,N_1911);
or U3900 (N_3900,N_2334,N_1667);
nand U3901 (N_3901,N_1694,N_2468);
nand U3902 (N_3902,N_2321,N_2821);
xor U3903 (N_3903,N_2441,N_2899);
nor U3904 (N_3904,N_2083,N_2418);
nand U3905 (N_3905,N_2199,N_2745);
nand U3906 (N_3906,N_1646,N_2279);
or U3907 (N_3907,N_2992,N_2103);
xnor U3908 (N_3908,N_2553,N_1574);
xnor U3909 (N_3909,N_2326,N_2232);
nor U3910 (N_3910,N_2060,N_2817);
nor U3911 (N_3911,N_2534,N_1751);
nand U3912 (N_3912,N_1919,N_2915);
and U3913 (N_3913,N_2953,N_2850);
and U3914 (N_3914,N_1549,N_2186);
nor U3915 (N_3915,N_2275,N_2915);
and U3916 (N_3916,N_2154,N_2295);
xnor U3917 (N_3917,N_2412,N_1657);
or U3918 (N_3918,N_2799,N_1536);
nand U3919 (N_3919,N_1965,N_2589);
and U3920 (N_3920,N_1694,N_2043);
nor U3921 (N_3921,N_2284,N_2312);
nor U3922 (N_3922,N_2023,N_2353);
and U3923 (N_3923,N_2986,N_2258);
or U3924 (N_3924,N_2190,N_2147);
xor U3925 (N_3925,N_2789,N_1569);
and U3926 (N_3926,N_2853,N_2279);
and U3927 (N_3927,N_2120,N_2685);
nor U3928 (N_3928,N_2552,N_2627);
and U3929 (N_3929,N_2883,N_2416);
nor U3930 (N_3930,N_1923,N_1638);
xor U3931 (N_3931,N_1770,N_2110);
and U3932 (N_3932,N_2855,N_1753);
and U3933 (N_3933,N_2010,N_1959);
or U3934 (N_3934,N_2805,N_2216);
nand U3935 (N_3935,N_2701,N_2904);
or U3936 (N_3936,N_2950,N_2459);
or U3937 (N_3937,N_2074,N_1872);
nor U3938 (N_3938,N_2372,N_1947);
nor U3939 (N_3939,N_2487,N_1902);
nand U3940 (N_3940,N_2546,N_2120);
and U3941 (N_3941,N_2308,N_2603);
and U3942 (N_3942,N_2857,N_2199);
and U3943 (N_3943,N_1546,N_2197);
nand U3944 (N_3944,N_2306,N_1706);
nor U3945 (N_3945,N_2373,N_2197);
nor U3946 (N_3946,N_2844,N_2680);
or U3947 (N_3947,N_2562,N_1977);
nand U3948 (N_3948,N_1797,N_2881);
xor U3949 (N_3949,N_1520,N_1952);
nor U3950 (N_3950,N_2422,N_1797);
and U3951 (N_3951,N_2070,N_2369);
or U3952 (N_3952,N_2306,N_2507);
and U3953 (N_3953,N_1777,N_2764);
and U3954 (N_3954,N_2151,N_1948);
nand U3955 (N_3955,N_2887,N_2781);
nor U3956 (N_3956,N_2851,N_1791);
nand U3957 (N_3957,N_2791,N_2064);
nand U3958 (N_3958,N_1959,N_2551);
nor U3959 (N_3959,N_2508,N_2475);
nor U3960 (N_3960,N_2465,N_2933);
nor U3961 (N_3961,N_2926,N_2633);
xnor U3962 (N_3962,N_2785,N_2926);
or U3963 (N_3963,N_2488,N_1814);
and U3964 (N_3964,N_2083,N_1664);
nor U3965 (N_3965,N_1797,N_2014);
or U3966 (N_3966,N_2260,N_2822);
xnor U3967 (N_3967,N_1917,N_1558);
nand U3968 (N_3968,N_2288,N_2702);
nand U3969 (N_3969,N_2521,N_2010);
nand U3970 (N_3970,N_2207,N_1542);
and U3971 (N_3971,N_1743,N_2580);
nand U3972 (N_3972,N_1856,N_2831);
nor U3973 (N_3973,N_2222,N_1864);
xnor U3974 (N_3974,N_1960,N_1957);
or U3975 (N_3975,N_1881,N_2738);
nor U3976 (N_3976,N_2802,N_2501);
or U3977 (N_3977,N_2886,N_2272);
nor U3978 (N_3978,N_2630,N_1916);
nand U3979 (N_3979,N_2930,N_2287);
nand U3980 (N_3980,N_2308,N_2024);
xor U3981 (N_3981,N_2366,N_2651);
xor U3982 (N_3982,N_2462,N_2362);
and U3983 (N_3983,N_1800,N_1688);
xor U3984 (N_3984,N_2759,N_1900);
or U3985 (N_3985,N_2650,N_2240);
nor U3986 (N_3986,N_2314,N_1848);
xor U3987 (N_3987,N_1505,N_2921);
nand U3988 (N_3988,N_2936,N_2397);
or U3989 (N_3989,N_2159,N_2586);
nand U3990 (N_3990,N_1783,N_2270);
nand U3991 (N_3991,N_1833,N_2361);
nor U3992 (N_3992,N_2785,N_2208);
nand U3993 (N_3993,N_2304,N_1531);
nor U3994 (N_3994,N_1588,N_2080);
and U3995 (N_3995,N_2228,N_2124);
nand U3996 (N_3996,N_2983,N_2674);
and U3997 (N_3997,N_1598,N_2339);
or U3998 (N_3998,N_2819,N_1920);
nand U3999 (N_3999,N_1941,N_2668);
nand U4000 (N_4000,N_2506,N_2541);
nand U4001 (N_4001,N_2600,N_2063);
or U4002 (N_4002,N_2601,N_1576);
nor U4003 (N_4003,N_2359,N_2935);
xor U4004 (N_4004,N_1530,N_1767);
nor U4005 (N_4005,N_2911,N_1503);
and U4006 (N_4006,N_2255,N_1595);
nand U4007 (N_4007,N_2880,N_1608);
and U4008 (N_4008,N_1716,N_2768);
and U4009 (N_4009,N_1992,N_2199);
and U4010 (N_4010,N_2994,N_2893);
or U4011 (N_4011,N_2189,N_2069);
nor U4012 (N_4012,N_1767,N_1821);
nand U4013 (N_4013,N_2456,N_1564);
xor U4014 (N_4014,N_2738,N_1999);
or U4015 (N_4015,N_2384,N_2313);
and U4016 (N_4016,N_2001,N_2513);
nand U4017 (N_4017,N_2378,N_2548);
and U4018 (N_4018,N_1835,N_2453);
or U4019 (N_4019,N_2818,N_2617);
and U4020 (N_4020,N_2018,N_1626);
nand U4021 (N_4021,N_2362,N_1538);
nor U4022 (N_4022,N_2794,N_2304);
or U4023 (N_4023,N_1921,N_1998);
xor U4024 (N_4024,N_2263,N_1992);
nand U4025 (N_4025,N_2154,N_1530);
nand U4026 (N_4026,N_2346,N_2286);
or U4027 (N_4027,N_1875,N_2299);
nor U4028 (N_4028,N_1808,N_1605);
nor U4029 (N_4029,N_2247,N_1672);
nor U4030 (N_4030,N_2005,N_1861);
or U4031 (N_4031,N_2716,N_2097);
nor U4032 (N_4032,N_2820,N_2439);
nand U4033 (N_4033,N_2132,N_1776);
nand U4034 (N_4034,N_2765,N_2920);
nand U4035 (N_4035,N_1691,N_2954);
xnor U4036 (N_4036,N_2408,N_2513);
nor U4037 (N_4037,N_2210,N_2354);
nand U4038 (N_4038,N_1654,N_1597);
nand U4039 (N_4039,N_1952,N_2733);
nor U4040 (N_4040,N_2638,N_1675);
nor U4041 (N_4041,N_2888,N_1652);
or U4042 (N_4042,N_2799,N_1705);
or U4043 (N_4043,N_1817,N_2731);
or U4044 (N_4044,N_2538,N_1968);
nor U4045 (N_4045,N_1761,N_1573);
nor U4046 (N_4046,N_2571,N_2262);
or U4047 (N_4047,N_1805,N_1940);
nor U4048 (N_4048,N_1524,N_2824);
and U4049 (N_4049,N_2575,N_1685);
nor U4050 (N_4050,N_1803,N_2508);
nand U4051 (N_4051,N_2234,N_2210);
xor U4052 (N_4052,N_1879,N_2136);
nand U4053 (N_4053,N_2993,N_2923);
and U4054 (N_4054,N_1503,N_1553);
or U4055 (N_4055,N_1546,N_2226);
or U4056 (N_4056,N_2865,N_2013);
or U4057 (N_4057,N_2742,N_2134);
xor U4058 (N_4058,N_1530,N_2202);
and U4059 (N_4059,N_2431,N_2351);
nor U4060 (N_4060,N_2672,N_1801);
nand U4061 (N_4061,N_2017,N_2276);
and U4062 (N_4062,N_1592,N_2439);
nor U4063 (N_4063,N_1556,N_2645);
nand U4064 (N_4064,N_1597,N_2216);
or U4065 (N_4065,N_2961,N_2982);
nand U4066 (N_4066,N_2227,N_2437);
nor U4067 (N_4067,N_2336,N_2092);
nand U4068 (N_4068,N_2687,N_1969);
and U4069 (N_4069,N_1827,N_2094);
xnor U4070 (N_4070,N_2892,N_1689);
nor U4071 (N_4071,N_1514,N_2869);
xnor U4072 (N_4072,N_2188,N_2912);
and U4073 (N_4073,N_2421,N_2506);
and U4074 (N_4074,N_2026,N_2463);
nand U4075 (N_4075,N_1530,N_2819);
nand U4076 (N_4076,N_2051,N_2392);
nand U4077 (N_4077,N_1765,N_2420);
and U4078 (N_4078,N_2328,N_2786);
and U4079 (N_4079,N_2790,N_1735);
nor U4080 (N_4080,N_2226,N_1653);
nand U4081 (N_4081,N_2660,N_2652);
nor U4082 (N_4082,N_2385,N_1582);
nor U4083 (N_4083,N_1918,N_2039);
nand U4084 (N_4084,N_2689,N_2485);
or U4085 (N_4085,N_2424,N_1571);
nand U4086 (N_4086,N_2329,N_1761);
and U4087 (N_4087,N_1861,N_2188);
or U4088 (N_4088,N_2268,N_2304);
nor U4089 (N_4089,N_2695,N_2306);
nand U4090 (N_4090,N_2273,N_1624);
or U4091 (N_4091,N_2539,N_1817);
nand U4092 (N_4092,N_1992,N_2881);
nor U4093 (N_4093,N_1519,N_2464);
nand U4094 (N_4094,N_2870,N_1592);
nor U4095 (N_4095,N_1873,N_1508);
nor U4096 (N_4096,N_1756,N_1822);
nand U4097 (N_4097,N_2173,N_2166);
or U4098 (N_4098,N_1652,N_2510);
or U4099 (N_4099,N_2388,N_2432);
xor U4100 (N_4100,N_1516,N_1791);
xnor U4101 (N_4101,N_1893,N_1978);
and U4102 (N_4102,N_1818,N_2910);
nor U4103 (N_4103,N_2471,N_2714);
or U4104 (N_4104,N_2130,N_2286);
nand U4105 (N_4105,N_2365,N_2392);
and U4106 (N_4106,N_2660,N_2071);
or U4107 (N_4107,N_1760,N_1927);
or U4108 (N_4108,N_2249,N_1693);
and U4109 (N_4109,N_1751,N_1509);
or U4110 (N_4110,N_1926,N_2278);
or U4111 (N_4111,N_2478,N_1874);
nand U4112 (N_4112,N_2265,N_2111);
nor U4113 (N_4113,N_1913,N_2088);
nand U4114 (N_4114,N_1805,N_2569);
nand U4115 (N_4115,N_2970,N_1965);
nor U4116 (N_4116,N_2496,N_2244);
nor U4117 (N_4117,N_2755,N_2136);
xor U4118 (N_4118,N_2103,N_2273);
nor U4119 (N_4119,N_2739,N_2849);
and U4120 (N_4120,N_1807,N_1775);
and U4121 (N_4121,N_2076,N_1643);
or U4122 (N_4122,N_1737,N_2256);
nand U4123 (N_4123,N_2324,N_1868);
and U4124 (N_4124,N_2377,N_1545);
nand U4125 (N_4125,N_2492,N_1956);
nand U4126 (N_4126,N_2070,N_2524);
xor U4127 (N_4127,N_1757,N_2727);
or U4128 (N_4128,N_1538,N_1787);
or U4129 (N_4129,N_2537,N_2483);
and U4130 (N_4130,N_2819,N_2937);
xor U4131 (N_4131,N_2955,N_2567);
and U4132 (N_4132,N_2472,N_1660);
nand U4133 (N_4133,N_1907,N_2989);
or U4134 (N_4134,N_2738,N_2378);
nor U4135 (N_4135,N_2172,N_2035);
nand U4136 (N_4136,N_2379,N_2299);
and U4137 (N_4137,N_1576,N_2218);
xor U4138 (N_4138,N_2321,N_2018);
or U4139 (N_4139,N_2119,N_2890);
nand U4140 (N_4140,N_2781,N_2652);
nand U4141 (N_4141,N_1658,N_1584);
nor U4142 (N_4142,N_2803,N_2861);
or U4143 (N_4143,N_2835,N_2819);
and U4144 (N_4144,N_2749,N_2681);
nand U4145 (N_4145,N_1897,N_2639);
xnor U4146 (N_4146,N_2840,N_2263);
nor U4147 (N_4147,N_2938,N_2016);
or U4148 (N_4148,N_2432,N_1687);
or U4149 (N_4149,N_2798,N_1954);
nor U4150 (N_4150,N_2516,N_1637);
or U4151 (N_4151,N_2409,N_2976);
xnor U4152 (N_4152,N_2235,N_2592);
nand U4153 (N_4153,N_2398,N_2858);
nand U4154 (N_4154,N_1963,N_2485);
and U4155 (N_4155,N_2542,N_2943);
or U4156 (N_4156,N_2183,N_1671);
nor U4157 (N_4157,N_2206,N_1774);
or U4158 (N_4158,N_1735,N_2414);
nor U4159 (N_4159,N_2313,N_2864);
or U4160 (N_4160,N_2098,N_1961);
nand U4161 (N_4161,N_2393,N_2169);
nand U4162 (N_4162,N_2379,N_2459);
nor U4163 (N_4163,N_1812,N_2703);
nor U4164 (N_4164,N_2217,N_2626);
nor U4165 (N_4165,N_2071,N_1774);
or U4166 (N_4166,N_2483,N_2784);
nand U4167 (N_4167,N_1804,N_2973);
nor U4168 (N_4168,N_1661,N_2058);
and U4169 (N_4169,N_1609,N_2618);
or U4170 (N_4170,N_2885,N_1820);
and U4171 (N_4171,N_2976,N_2794);
xor U4172 (N_4172,N_1595,N_2270);
nor U4173 (N_4173,N_2812,N_2792);
xor U4174 (N_4174,N_1751,N_2212);
and U4175 (N_4175,N_2839,N_2116);
or U4176 (N_4176,N_2982,N_1657);
nand U4177 (N_4177,N_2957,N_1830);
and U4178 (N_4178,N_1984,N_2033);
nand U4179 (N_4179,N_2579,N_1876);
nand U4180 (N_4180,N_2301,N_1575);
xor U4181 (N_4181,N_2837,N_2341);
or U4182 (N_4182,N_2081,N_2511);
or U4183 (N_4183,N_2956,N_2091);
nor U4184 (N_4184,N_1918,N_2711);
or U4185 (N_4185,N_2000,N_2606);
nand U4186 (N_4186,N_2952,N_2426);
or U4187 (N_4187,N_1583,N_2706);
or U4188 (N_4188,N_2306,N_1695);
nor U4189 (N_4189,N_1969,N_2648);
or U4190 (N_4190,N_2156,N_2890);
and U4191 (N_4191,N_1897,N_2444);
or U4192 (N_4192,N_2897,N_2867);
or U4193 (N_4193,N_2415,N_2308);
xor U4194 (N_4194,N_1991,N_2137);
or U4195 (N_4195,N_2163,N_1768);
and U4196 (N_4196,N_2633,N_2235);
nor U4197 (N_4197,N_2244,N_2396);
nor U4198 (N_4198,N_2887,N_2079);
nand U4199 (N_4199,N_2882,N_1703);
and U4200 (N_4200,N_2533,N_1772);
or U4201 (N_4201,N_2201,N_1968);
or U4202 (N_4202,N_2559,N_1866);
and U4203 (N_4203,N_2889,N_2602);
and U4204 (N_4204,N_2172,N_2947);
or U4205 (N_4205,N_2784,N_2152);
nor U4206 (N_4206,N_2374,N_2765);
and U4207 (N_4207,N_2189,N_1795);
and U4208 (N_4208,N_1754,N_2553);
or U4209 (N_4209,N_2589,N_1606);
xnor U4210 (N_4210,N_1782,N_2334);
nor U4211 (N_4211,N_2628,N_2603);
nand U4212 (N_4212,N_2816,N_2629);
and U4213 (N_4213,N_2807,N_2559);
and U4214 (N_4214,N_2129,N_2957);
xnor U4215 (N_4215,N_1903,N_1821);
nand U4216 (N_4216,N_2593,N_1775);
nand U4217 (N_4217,N_1567,N_1726);
nand U4218 (N_4218,N_2937,N_2820);
or U4219 (N_4219,N_2441,N_2385);
and U4220 (N_4220,N_2088,N_2628);
nor U4221 (N_4221,N_2323,N_2250);
nand U4222 (N_4222,N_1806,N_1610);
and U4223 (N_4223,N_2901,N_2548);
nand U4224 (N_4224,N_1842,N_2929);
or U4225 (N_4225,N_1554,N_2290);
and U4226 (N_4226,N_1671,N_1632);
nand U4227 (N_4227,N_1697,N_1906);
and U4228 (N_4228,N_1978,N_2949);
and U4229 (N_4229,N_1883,N_1833);
nand U4230 (N_4230,N_1771,N_2765);
and U4231 (N_4231,N_2284,N_2575);
or U4232 (N_4232,N_2452,N_2765);
xor U4233 (N_4233,N_2936,N_1675);
nor U4234 (N_4234,N_2224,N_2963);
nor U4235 (N_4235,N_2560,N_2926);
or U4236 (N_4236,N_1694,N_2849);
or U4237 (N_4237,N_2283,N_2132);
nor U4238 (N_4238,N_2041,N_1764);
and U4239 (N_4239,N_1559,N_1862);
or U4240 (N_4240,N_1605,N_2585);
and U4241 (N_4241,N_2105,N_2225);
nand U4242 (N_4242,N_2745,N_2774);
nor U4243 (N_4243,N_2345,N_2111);
or U4244 (N_4244,N_2973,N_1826);
nand U4245 (N_4245,N_2215,N_1598);
and U4246 (N_4246,N_1567,N_2435);
xnor U4247 (N_4247,N_1978,N_1584);
and U4248 (N_4248,N_2876,N_2060);
or U4249 (N_4249,N_2646,N_2136);
or U4250 (N_4250,N_2692,N_2821);
or U4251 (N_4251,N_2912,N_1755);
or U4252 (N_4252,N_1667,N_1712);
and U4253 (N_4253,N_2901,N_2453);
nor U4254 (N_4254,N_2491,N_2969);
nand U4255 (N_4255,N_2633,N_1547);
and U4256 (N_4256,N_1877,N_1510);
or U4257 (N_4257,N_1732,N_2871);
and U4258 (N_4258,N_2489,N_2566);
nand U4259 (N_4259,N_2360,N_2784);
nand U4260 (N_4260,N_2448,N_2400);
or U4261 (N_4261,N_2352,N_2427);
or U4262 (N_4262,N_2359,N_2229);
nand U4263 (N_4263,N_1981,N_2268);
nor U4264 (N_4264,N_2043,N_1634);
xnor U4265 (N_4265,N_2509,N_2997);
nor U4266 (N_4266,N_2152,N_2463);
xnor U4267 (N_4267,N_2092,N_2921);
nor U4268 (N_4268,N_2807,N_2389);
and U4269 (N_4269,N_1509,N_2796);
xor U4270 (N_4270,N_2651,N_1865);
nand U4271 (N_4271,N_1662,N_2001);
or U4272 (N_4272,N_2981,N_2572);
or U4273 (N_4273,N_2948,N_1720);
or U4274 (N_4274,N_1999,N_2959);
or U4275 (N_4275,N_2188,N_2590);
and U4276 (N_4276,N_2329,N_2728);
nand U4277 (N_4277,N_2084,N_2351);
nand U4278 (N_4278,N_2178,N_2596);
nand U4279 (N_4279,N_2454,N_2887);
nor U4280 (N_4280,N_2746,N_2104);
and U4281 (N_4281,N_2934,N_2484);
nand U4282 (N_4282,N_2142,N_1517);
xnor U4283 (N_4283,N_2319,N_1850);
nand U4284 (N_4284,N_2621,N_1570);
xnor U4285 (N_4285,N_2049,N_2802);
nor U4286 (N_4286,N_2272,N_2372);
nor U4287 (N_4287,N_2549,N_2822);
or U4288 (N_4288,N_2257,N_2726);
or U4289 (N_4289,N_2874,N_2573);
nand U4290 (N_4290,N_2836,N_2246);
xor U4291 (N_4291,N_2104,N_1828);
and U4292 (N_4292,N_2158,N_1858);
nand U4293 (N_4293,N_2012,N_2808);
nand U4294 (N_4294,N_1724,N_2533);
xnor U4295 (N_4295,N_2254,N_2470);
and U4296 (N_4296,N_1809,N_1967);
nand U4297 (N_4297,N_2851,N_2482);
or U4298 (N_4298,N_1624,N_2418);
nand U4299 (N_4299,N_1858,N_2802);
and U4300 (N_4300,N_2371,N_2514);
nor U4301 (N_4301,N_2298,N_2955);
xor U4302 (N_4302,N_2085,N_2657);
xor U4303 (N_4303,N_1793,N_1897);
and U4304 (N_4304,N_2342,N_2476);
or U4305 (N_4305,N_2452,N_1976);
nor U4306 (N_4306,N_2248,N_2346);
or U4307 (N_4307,N_1696,N_1748);
nand U4308 (N_4308,N_2026,N_2273);
or U4309 (N_4309,N_2407,N_1583);
nand U4310 (N_4310,N_1585,N_2701);
xor U4311 (N_4311,N_2179,N_2503);
nor U4312 (N_4312,N_1555,N_2509);
and U4313 (N_4313,N_2472,N_2380);
nor U4314 (N_4314,N_1907,N_1983);
xnor U4315 (N_4315,N_1960,N_1779);
and U4316 (N_4316,N_2674,N_2222);
nand U4317 (N_4317,N_1917,N_2811);
or U4318 (N_4318,N_2362,N_2030);
and U4319 (N_4319,N_1537,N_2239);
or U4320 (N_4320,N_2908,N_2466);
and U4321 (N_4321,N_2660,N_1973);
nor U4322 (N_4322,N_1500,N_2648);
nand U4323 (N_4323,N_1601,N_2505);
or U4324 (N_4324,N_2141,N_2903);
or U4325 (N_4325,N_2802,N_1758);
nand U4326 (N_4326,N_2272,N_2716);
or U4327 (N_4327,N_2806,N_2859);
and U4328 (N_4328,N_2119,N_2782);
xor U4329 (N_4329,N_1624,N_1577);
xor U4330 (N_4330,N_1807,N_2071);
nand U4331 (N_4331,N_1785,N_2733);
or U4332 (N_4332,N_2133,N_2271);
nand U4333 (N_4333,N_2105,N_2962);
nand U4334 (N_4334,N_2714,N_2664);
and U4335 (N_4335,N_1594,N_2729);
xnor U4336 (N_4336,N_2037,N_1586);
and U4337 (N_4337,N_2067,N_1712);
nor U4338 (N_4338,N_2304,N_1788);
nor U4339 (N_4339,N_2824,N_2240);
and U4340 (N_4340,N_1868,N_2573);
xor U4341 (N_4341,N_2083,N_2401);
nor U4342 (N_4342,N_2728,N_1895);
and U4343 (N_4343,N_2043,N_2731);
or U4344 (N_4344,N_2770,N_1668);
nor U4345 (N_4345,N_1792,N_2142);
or U4346 (N_4346,N_1650,N_1936);
or U4347 (N_4347,N_2377,N_2416);
nor U4348 (N_4348,N_2217,N_2782);
nand U4349 (N_4349,N_2836,N_1521);
nand U4350 (N_4350,N_2648,N_1771);
nand U4351 (N_4351,N_2057,N_2533);
and U4352 (N_4352,N_2144,N_1879);
or U4353 (N_4353,N_2472,N_2116);
or U4354 (N_4354,N_1782,N_2355);
and U4355 (N_4355,N_2191,N_1989);
nor U4356 (N_4356,N_1872,N_2621);
and U4357 (N_4357,N_1676,N_2004);
nor U4358 (N_4358,N_2627,N_2428);
or U4359 (N_4359,N_1944,N_2253);
nand U4360 (N_4360,N_2461,N_2951);
and U4361 (N_4361,N_1751,N_2022);
nor U4362 (N_4362,N_2836,N_2718);
and U4363 (N_4363,N_1896,N_2049);
or U4364 (N_4364,N_1742,N_2199);
and U4365 (N_4365,N_2459,N_2841);
and U4366 (N_4366,N_1762,N_1835);
or U4367 (N_4367,N_1750,N_2999);
and U4368 (N_4368,N_1625,N_2151);
and U4369 (N_4369,N_2690,N_2890);
nand U4370 (N_4370,N_2403,N_1998);
nand U4371 (N_4371,N_1932,N_2248);
nor U4372 (N_4372,N_2670,N_2168);
xnor U4373 (N_4373,N_2766,N_1677);
xnor U4374 (N_4374,N_1549,N_2773);
or U4375 (N_4375,N_2756,N_2805);
and U4376 (N_4376,N_2799,N_2329);
nor U4377 (N_4377,N_1872,N_2775);
xor U4378 (N_4378,N_2365,N_2682);
xnor U4379 (N_4379,N_1726,N_1608);
and U4380 (N_4380,N_2626,N_1614);
nor U4381 (N_4381,N_1580,N_1574);
and U4382 (N_4382,N_2811,N_2401);
or U4383 (N_4383,N_1929,N_1924);
nor U4384 (N_4384,N_2101,N_2531);
nand U4385 (N_4385,N_2016,N_2037);
and U4386 (N_4386,N_2483,N_2464);
and U4387 (N_4387,N_2462,N_2843);
nor U4388 (N_4388,N_1807,N_1818);
nor U4389 (N_4389,N_2008,N_2979);
or U4390 (N_4390,N_1820,N_2141);
nand U4391 (N_4391,N_2363,N_2249);
nor U4392 (N_4392,N_2035,N_2657);
nand U4393 (N_4393,N_1706,N_2565);
and U4394 (N_4394,N_1808,N_1589);
and U4395 (N_4395,N_1986,N_2505);
and U4396 (N_4396,N_1946,N_2616);
or U4397 (N_4397,N_2648,N_1599);
and U4398 (N_4398,N_1898,N_2092);
or U4399 (N_4399,N_2182,N_2120);
and U4400 (N_4400,N_2337,N_2235);
and U4401 (N_4401,N_1641,N_1647);
nand U4402 (N_4402,N_2485,N_2244);
nand U4403 (N_4403,N_1793,N_2153);
or U4404 (N_4404,N_2856,N_2737);
nor U4405 (N_4405,N_2730,N_2412);
or U4406 (N_4406,N_2275,N_2567);
or U4407 (N_4407,N_2542,N_2567);
or U4408 (N_4408,N_2663,N_2673);
and U4409 (N_4409,N_1796,N_2576);
and U4410 (N_4410,N_1926,N_2518);
nor U4411 (N_4411,N_2661,N_2716);
or U4412 (N_4412,N_1641,N_2217);
or U4413 (N_4413,N_2617,N_2886);
and U4414 (N_4414,N_2304,N_1924);
or U4415 (N_4415,N_2282,N_2529);
nand U4416 (N_4416,N_2388,N_1916);
xnor U4417 (N_4417,N_2181,N_1549);
or U4418 (N_4418,N_1740,N_2197);
and U4419 (N_4419,N_2746,N_1548);
and U4420 (N_4420,N_2372,N_2576);
or U4421 (N_4421,N_1714,N_2702);
nor U4422 (N_4422,N_2796,N_1630);
nand U4423 (N_4423,N_2562,N_1720);
nor U4424 (N_4424,N_2911,N_2082);
nor U4425 (N_4425,N_2076,N_1703);
and U4426 (N_4426,N_2458,N_1873);
nor U4427 (N_4427,N_1941,N_2273);
nand U4428 (N_4428,N_2631,N_1737);
nand U4429 (N_4429,N_2649,N_2335);
nand U4430 (N_4430,N_2835,N_1577);
and U4431 (N_4431,N_2303,N_2842);
nor U4432 (N_4432,N_2675,N_2817);
and U4433 (N_4433,N_2617,N_1628);
nor U4434 (N_4434,N_2925,N_2714);
and U4435 (N_4435,N_2407,N_2374);
or U4436 (N_4436,N_2284,N_2572);
xor U4437 (N_4437,N_1662,N_2162);
xor U4438 (N_4438,N_2012,N_2534);
or U4439 (N_4439,N_2789,N_2817);
nor U4440 (N_4440,N_2208,N_2313);
nand U4441 (N_4441,N_2873,N_2182);
or U4442 (N_4442,N_1629,N_2345);
and U4443 (N_4443,N_1774,N_1687);
nand U4444 (N_4444,N_2640,N_2177);
nor U4445 (N_4445,N_1742,N_1636);
nand U4446 (N_4446,N_1625,N_2320);
or U4447 (N_4447,N_1651,N_2351);
nand U4448 (N_4448,N_1746,N_2400);
xor U4449 (N_4449,N_1719,N_2625);
nand U4450 (N_4450,N_2233,N_1596);
or U4451 (N_4451,N_2516,N_1931);
nand U4452 (N_4452,N_1951,N_2318);
nor U4453 (N_4453,N_2829,N_1522);
nor U4454 (N_4454,N_1862,N_2511);
xnor U4455 (N_4455,N_2301,N_2624);
and U4456 (N_4456,N_1672,N_1775);
or U4457 (N_4457,N_2659,N_2094);
nor U4458 (N_4458,N_2837,N_2031);
nand U4459 (N_4459,N_2871,N_1969);
and U4460 (N_4460,N_1608,N_1873);
or U4461 (N_4461,N_2430,N_2579);
or U4462 (N_4462,N_2208,N_2711);
nand U4463 (N_4463,N_1939,N_2856);
and U4464 (N_4464,N_1777,N_1605);
xor U4465 (N_4465,N_1902,N_1726);
xor U4466 (N_4466,N_2557,N_2990);
or U4467 (N_4467,N_2907,N_2445);
nand U4468 (N_4468,N_2642,N_1564);
or U4469 (N_4469,N_2516,N_1817);
nand U4470 (N_4470,N_1683,N_1592);
nor U4471 (N_4471,N_1800,N_1518);
or U4472 (N_4472,N_1812,N_2704);
nor U4473 (N_4473,N_2834,N_2601);
nor U4474 (N_4474,N_2563,N_2502);
nand U4475 (N_4475,N_2737,N_2489);
or U4476 (N_4476,N_1649,N_1755);
or U4477 (N_4477,N_1879,N_2523);
nand U4478 (N_4478,N_2314,N_2013);
or U4479 (N_4479,N_2667,N_2157);
nor U4480 (N_4480,N_2584,N_1889);
or U4481 (N_4481,N_1980,N_1748);
or U4482 (N_4482,N_1632,N_2910);
nand U4483 (N_4483,N_2053,N_1818);
nor U4484 (N_4484,N_2577,N_2410);
xor U4485 (N_4485,N_2255,N_2772);
xor U4486 (N_4486,N_2017,N_2910);
or U4487 (N_4487,N_2866,N_1705);
or U4488 (N_4488,N_2857,N_1715);
nor U4489 (N_4489,N_1545,N_2727);
nand U4490 (N_4490,N_1538,N_2402);
or U4491 (N_4491,N_2748,N_2985);
or U4492 (N_4492,N_2124,N_1770);
and U4493 (N_4493,N_2271,N_1947);
nor U4494 (N_4494,N_1935,N_1843);
and U4495 (N_4495,N_1607,N_2660);
nor U4496 (N_4496,N_2005,N_2846);
and U4497 (N_4497,N_1873,N_2067);
or U4498 (N_4498,N_2131,N_2664);
and U4499 (N_4499,N_2461,N_1905);
nor U4500 (N_4500,N_3362,N_4266);
nand U4501 (N_4501,N_3925,N_4249);
and U4502 (N_4502,N_3759,N_4165);
nand U4503 (N_4503,N_4365,N_3817);
or U4504 (N_4504,N_3417,N_3806);
and U4505 (N_4505,N_3116,N_3299);
or U4506 (N_4506,N_4236,N_4119);
and U4507 (N_4507,N_3536,N_3283);
nand U4508 (N_4508,N_4333,N_4486);
or U4509 (N_4509,N_3413,N_3408);
and U4510 (N_4510,N_3240,N_3168);
nor U4511 (N_4511,N_3169,N_4086);
nor U4512 (N_4512,N_3361,N_4116);
xor U4513 (N_4513,N_3162,N_3991);
and U4514 (N_4514,N_3881,N_3357);
and U4515 (N_4515,N_3173,N_3515);
or U4516 (N_4516,N_3183,N_3669);
or U4517 (N_4517,N_3238,N_3314);
nor U4518 (N_4518,N_3657,N_3172);
nor U4519 (N_4519,N_4408,N_3031);
or U4520 (N_4520,N_3223,N_3092);
nand U4521 (N_4521,N_3834,N_3527);
and U4522 (N_4522,N_4391,N_4207);
nor U4523 (N_4523,N_3562,N_3350);
and U4524 (N_4524,N_3139,N_3454);
nand U4525 (N_4525,N_3504,N_3973);
or U4526 (N_4526,N_4407,N_3672);
nor U4527 (N_4527,N_3255,N_3488);
and U4528 (N_4528,N_4025,N_3443);
or U4529 (N_4529,N_4421,N_3127);
nor U4530 (N_4530,N_3550,N_3206);
nor U4531 (N_4531,N_4048,N_3793);
nand U4532 (N_4532,N_3658,N_3323);
nand U4533 (N_4533,N_4477,N_4087);
nand U4534 (N_4534,N_3298,N_4103);
nor U4535 (N_4535,N_3105,N_3847);
nor U4536 (N_4536,N_3122,N_4109);
xor U4537 (N_4537,N_3479,N_4436);
or U4538 (N_4538,N_3341,N_3349);
nor U4539 (N_4539,N_3107,N_4425);
and U4540 (N_4540,N_3640,N_4275);
nor U4541 (N_4541,N_4305,N_3854);
or U4542 (N_4542,N_3900,N_3216);
and U4543 (N_4543,N_3386,N_3970);
nand U4544 (N_4544,N_3044,N_3701);
xor U4545 (N_4545,N_3019,N_3387);
nor U4546 (N_4546,N_3380,N_4495);
nor U4547 (N_4547,N_3346,N_3251);
nand U4548 (N_4548,N_4221,N_4016);
or U4549 (N_4549,N_3750,N_3020);
and U4550 (N_4550,N_3115,N_3785);
or U4551 (N_4551,N_4121,N_4398);
nor U4552 (N_4552,N_4198,N_3078);
nand U4553 (N_4553,N_4279,N_3871);
nor U4554 (N_4554,N_4232,N_3137);
nor U4555 (N_4555,N_3998,N_3334);
and U4556 (N_4556,N_4280,N_3911);
and U4557 (N_4557,N_3419,N_3682);
nor U4558 (N_4558,N_3581,N_4335);
nor U4559 (N_4559,N_3770,N_4475);
nand U4560 (N_4560,N_3502,N_3542);
nand U4561 (N_4561,N_4277,N_4471);
and U4562 (N_4562,N_3561,N_3426);
or U4563 (N_4563,N_4110,N_4388);
xnor U4564 (N_4564,N_4215,N_3538);
nor U4565 (N_4565,N_3858,N_3850);
nand U4566 (N_4566,N_4002,N_3807);
and U4567 (N_4567,N_3204,N_3874);
or U4568 (N_4568,N_4019,N_3933);
xor U4569 (N_4569,N_4273,N_3400);
nand U4570 (N_4570,N_3348,N_4132);
nand U4571 (N_4571,N_3754,N_4341);
or U4572 (N_4572,N_3668,N_3614);
xor U4573 (N_4573,N_4428,N_4252);
nor U4574 (N_4574,N_3663,N_3302);
or U4575 (N_4575,N_3574,N_3601);
or U4576 (N_4576,N_3758,N_4043);
or U4577 (N_4577,N_3069,N_3823);
xnor U4578 (N_4578,N_3352,N_3313);
or U4579 (N_4579,N_3276,N_4039);
nor U4580 (N_4580,N_4395,N_3587);
xnor U4581 (N_4581,N_3976,N_4061);
nand U4582 (N_4582,N_4464,N_3713);
and U4583 (N_4583,N_3372,N_3332);
nor U4584 (N_4584,N_3039,N_4022);
xnor U4585 (N_4585,N_3779,N_3154);
nand U4586 (N_4586,N_4248,N_3336);
or U4587 (N_4587,N_3471,N_3133);
nor U4588 (N_4588,N_3493,N_4312);
and U4589 (N_4589,N_4005,N_4447);
nor U4590 (N_4590,N_3395,N_4065);
and U4591 (N_4591,N_4090,N_3214);
and U4592 (N_4592,N_3860,N_3450);
and U4593 (N_4593,N_4091,N_4327);
and U4594 (N_4594,N_3163,N_4489);
nand U4595 (N_4595,N_3123,N_3664);
xnor U4596 (N_4596,N_3370,N_3083);
or U4597 (N_4597,N_3947,N_3492);
nor U4598 (N_4598,N_3821,N_3851);
and U4599 (N_4599,N_3178,N_4401);
and U4600 (N_4600,N_4367,N_3780);
or U4601 (N_4601,N_3665,N_3928);
nand U4602 (N_4602,N_4353,N_3813);
nor U4603 (N_4603,N_4179,N_4308);
or U4604 (N_4604,N_3108,N_3942);
and U4605 (N_4605,N_4290,N_4117);
and U4606 (N_4606,N_4182,N_3433);
or U4607 (N_4607,N_3559,N_3756);
nand U4608 (N_4608,N_3247,N_3193);
and U4609 (N_4609,N_3610,N_3205);
or U4610 (N_4610,N_3902,N_3161);
or U4611 (N_4611,N_4427,N_3316);
or U4612 (N_4612,N_3279,N_3189);
and U4613 (N_4613,N_3062,N_3795);
and U4614 (N_4614,N_3853,N_3571);
nand U4615 (N_4615,N_3697,N_4097);
nand U4616 (N_4616,N_3551,N_3744);
nor U4617 (N_4617,N_3838,N_4054);
nand U4618 (N_4618,N_4219,N_3937);
nand U4619 (N_4619,N_3993,N_3704);
or U4620 (N_4620,N_3028,N_3954);
and U4621 (N_4621,N_4493,N_3337);
nand U4622 (N_4622,N_4191,N_4386);
or U4623 (N_4623,N_3125,N_3434);
and U4624 (N_4624,N_4155,N_3960);
or U4625 (N_4625,N_3643,N_3102);
and U4626 (N_4626,N_3285,N_4498);
and U4627 (N_4627,N_4139,N_4224);
or U4628 (N_4628,N_3344,N_3495);
nand U4629 (N_4629,N_3311,N_4185);
and U4630 (N_4630,N_3849,N_4411);
or U4631 (N_4631,N_3535,N_3702);
or U4632 (N_4632,N_3401,N_3877);
nand U4633 (N_4633,N_3962,N_3604);
xor U4634 (N_4634,N_4067,N_3570);
nor U4635 (N_4635,N_3320,N_4373);
xor U4636 (N_4636,N_3243,N_4034);
and U4637 (N_4637,N_3649,N_3233);
xor U4638 (N_4638,N_3670,N_3384);
and U4639 (N_4639,N_3152,N_3376);
nand U4640 (N_4640,N_3995,N_4233);
nor U4641 (N_4641,N_3715,N_3235);
or U4642 (N_4642,N_3690,N_3718);
or U4643 (N_4643,N_4080,N_3526);
and U4644 (N_4644,N_3470,N_3733);
nand U4645 (N_4645,N_3174,N_4461);
xor U4646 (N_4646,N_4038,N_4337);
or U4647 (N_4647,N_3772,N_3883);
nor U4648 (N_4648,N_4378,N_3143);
or U4649 (N_4649,N_4431,N_4063);
nor U4650 (N_4650,N_3671,N_4009);
and U4651 (N_4651,N_3931,N_3816);
nand U4652 (N_4652,N_4285,N_3113);
or U4653 (N_4653,N_3468,N_4326);
or U4654 (N_4654,N_3138,N_3425);
nor U4655 (N_4655,N_4348,N_3398);
or U4656 (N_4656,N_3792,N_4200);
nor U4657 (N_4657,N_4451,N_4301);
xor U4658 (N_4658,N_4294,N_3256);
or U4659 (N_4659,N_4357,N_4469);
nor U4660 (N_4660,N_3404,N_4089);
nor U4661 (N_4661,N_4223,N_4206);
or U4662 (N_4662,N_3148,N_4050);
and U4663 (N_4663,N_4258,N_4217);
nand U4664 (N_4664,N_4209,N_4346);
nand U4665 (N_4665,N_3119,N_4030);
and U4666 (N_4666,N_3629,N_3885);
nor U4667 (N_4667,N_4330,N_3677);
nor U4668 (N_4668,N_3236,N_4351);
nor U4669 (N_4669,N_3711,N_4146);
nand U4670 (N_4670,N_3104,N_3363);
or U4671 (N_4671,N_3819,N_4000);
nand U4672 (N_4672,N_3814,N_3192);
or U4673 (N_4673,N_3534,N_3429);
or U4674 (N_4674,N_3703,N_3953);
nand U4675 (N_4675,N_4366,N_4203);
or U4676 (N_4676,N_3552,N_3165);
xor U4677 (N_4677,N_3167,N_3655);
or U4678 (N_4678,N_4186,N_3449);
nor U4679 (N_4679,N_3719,N_4216);
nor U4680 (N_4680,N_3209,N_3354);
or U4681 (N_4681,N_4068,N_4083);
and U4682 (N_4682,N_3340,N_3013);
and U4683 (N_4683,N_3257,N_3961);
or U4684 (N_4684,N_3179,N_3540);
nor U4685 (N_4685,N_4144,N_3940);
or U4686 (N_4686,N_3339,N_4251);
and U4687 (N_4687,N_4066,N_3430);
or U4688 (N_4688,N_3654,N_3010);
and U4689 (N_4689,N_3373,N_4482);
and U4690 (N_4690,N_3788,N_3290);
and U4691 (N_4691,N_3547,N_3842);
nor U4692 (N_4692,N_3259,N_3465);
xor U4693 (N_4693,N_3140,N_3996);
nand U4694 (N_4694,N_3674,N_3843);
or U4695 (N_4695,N_4446,N_4164);
or U4696 (N_4696,N_3225,N_3331);
and U4697 (N_4697,N_3406,N_4350);
or U4698 (N_4698,N_3781,N_4332);
and U4699 (N_4699,N_3639,N_3926);
and U4700 (N_4700,N_3500,N_3729);
nand U4701 (N_4701,N_3676,N_4361);
and U4702 (N_4702,N_3695,N_3367);
or U4703 (N_4703,N_4174,N_4283);
xnor U4704 (N_4704,N_4118,N_3660);
nand U4705 (N_4705,N_3506,N_3051);
nor U4706 (N_4706,N_3560,N_3597);
and U4707 (N_4707,N_3907,N_3002);
nand U4708 (N_4708,N_3895,N_4169);
nor U4709 (N_4709,N_3977,N_3723);
or U4710 (N_4710,N_3833,N_3136);
nor U4711 (N_4711,N_3324,N_4007);
nand U4712 (N_4712,N_4081,N_4385);
nor U4713 (N_4713,N_4392,N_3056);
or U4714 (N_4714,N_3009,N_3612);
nand U4715 (N_4715,N_3472,N_4454);
and U4716 (N_4716,N_4276,N_3837);
and U4717 (N_4717,N_3171,N_3799);
nand U4718 (N_4718,N_3399,N_3959);
or U4719 (N_4719,N_3351,N_4499);
and U4720 (N_4720,N_3983,N_3721);
nand U4721 (N_4721,N_4329,N_3090);
and U4722 (N_4722,N_4404,N_3846);
and U4723 (N_4723,N_3096,N_4100);
and U4724 (N_4724,N_3045,N_3826);
and U4725 (N_4725,N_4462,N_4101);
or U4726 (N_4726,N_3200,N_4137);
nand U4727 (N_4727,N_3705,N_3130);
and U4728 (N_4728,N_4450,N_3912);
nor U4729 (N_4729,N_3360,N_3884);
or U4730 (N_4730,N_3445,N_3517);
nor U4731 (N_4731,N_3353,N_4126);
nand U4732 (N_4732,N_3730,N_3371);
nor U4733 (N_4733,N_3185,N_3249);
xnor U4734 (N_4734,N_4419,N_3789);
nand U4735 (N_4735,N_3613,N_4228);
xnor U4736 (N_4736,N_4140,N_3263);
and U4737 (N_4737,N_3924,N_3291);
xor U4738 (N_4738,N_3295,N_4439);
or U4739 (N_4739,N_3575,N_4311);
and U4740 (N_4740,N_4458,N_3057);
and U4741 (N_4741,N_3865,N_3067);
or U4742 (N_4742,N_3753,N_3231);
and U4743 (N_4743,N_3927,N_3461);
nand U4744 (N_4744,N_4355,N_3876);
and U4745 (N_4745,N_3024,N_4304);
or U4746 (N_4746,N_4014,N_3510);
or U4747 (N_4747,N_4173,N_4470);
nand U4748 (N_4748,N_4271,N_4284);
or U4749 (N_4749,N_3751,N_3687);
or U4750 (N_4750,N_4115,N_4131);
nand U4751 (N_4751,N_4405,N_4375);
and U4752 (N_4752,N_3988,N_3685);
and U4753 (N_4753,N_3981,N_4166);
xor U4754 (N_4754,N_3978,N_3388);
nand U4755 (N_4755,N_3935,N_4295);
or U4756 (N_4756,N_3309,N_3945);
nor U4757 (N_4757,N_3511,N_3153);
nor U4758 (N_4758,N_4124,N_3519);
nand U4759 (N_4759,N_4085,N_4261);
and U4760 (N_4760,N_4128,N_3058);
or U4761 (N_4761,N_4457,N_4210);
and U4762 (N_4762,N_3661,N_4278);
or U4763 (N_4763,N_3573,N_4364);
and U4764 (N_4764,N_3539,N_4269);
or U4765 (N_4765,N_3757,N_4363);
nand U4766 (N_4766,N_3748,N_3805);
nand U4767 (N_4767,N_4288,N_4073);
or U4768 (N_4768,N_3916,N_3512);
nand U4769 (N_4769,N_3260,N_3422);
and U4770 (N_4770,N_3393,N_3673);
nor U4771 (N_4771,N_3164,N_3446);
nor U4772 (N_4772,N_3097,N_3158);
and U4773 (N_4773,N_4352,N_3227);
nand U4774 (N_4774,N_3415,N_3159);
and U4775 (N_4775,N_3142,N_3287);
or U4776 (N_4776,N_3878,N_4231);
nand U4777 (N_4777,N_3347,N_4374);
xor U4778 (N_4778,N_4018,N_4322);
xor U4779 (N_4779,N_3368,N_3889);
nand U4780 (N_4780,N_3693,N_3600);
nand U4781 (N_4781,N_4317,N_4157);
nor U4782 (N_4782,N_4176,N_3210);
xnor U4783 (N_4783,N_4306,N_3557);
nor U4784 (N_4784,N_4340,N_4243);
nand U4785 (N_4785,N_4412,N_3199);
nand U4786 (N_4786,N_3830,N_3755);
and U4787 (N_4787,N_3622,N_3856);
and U4788 (N_4788,N_4430,N_3330);
xnor U4789 (N_4789,N_3088,N_3220);
nor U4790 (N_4790,N_4456,N_4397);
nand U4791 (N_4791,N_3118,N_3879);
and U4792 (N_4792,N_4298,N_4441);
or U4793 (N_4793,N_3463,N_4102);
xnor U4794 (N_4794,N_4187,N_3607);
or U4795 (N_4795,N_4370,N_3036);
and U4796 (N_4796,N_4171,N_3859);
nand U4797 (N_4797,N_3207,N_4256);
nor U4798 (N_4798,N_3052,N_4349);
or U4799 (N_4799,N_3228,N_3892);
or U4800 (N_4800,N_4247,N_4193);
xor U4801 (N_4801,N_3768,N_4422);
nand U4802 (N_4802,N_4133,N_3694);
nor U4803 (N_4803,N_3619,N_4196);
xor U4804 (N_4804,N_4282,N_3197);
nand U4805 (N_4805,N_3620,N_4088);
or U4806 (N_4806,N_3577,N_3219);
nor U4807 (N_4807,N_3369,N_3265);
xor U4808 (N_4808,N_3952,N_3794);
or U4809 (N_4809,N_3893,N_4094);
nand U4810 (N_4810,N_3188,N_4082);
or U4811 (N_4811,N_3822,N_3868);
or U4812 (N_4812,N_4180,N_3741);
nand U4813 (N_4813,N_3385,N_4234);
nand U4814 (N_4814,N_3021,N_3128);
nand U4815 (N_4815,N_3499,N_3835);
or U4816 (N_4816,N_3091,N_3094);
xor U4817 (N_4817,N_3477,N_3017);
xnor U4818 (N_4818,N_3064,N_3201);
nand U4819 (N_4819,N_3432,N_4031);
nand U4820 (N_4820,N_4310,N_4172);
and U4821 (N_4821,N_4112,N_4199);
and U4822 (N_4822,N_3531,N_4476);
nor U4823 (N_4823,N_4024,N_3637);
and U4824 (N_4824,N_3431,N_4409);
nand U4825 (N_4825,N_3599,N_4181);
or U4826 (N_4826,N_3319,N_4315);
xnor U4827 (N_4827,N_3111,N_3921);
nor U4828 (N_4828,N_3899,N_3913);
nand U4829 (N_4829,N_4064,N_3034);
and U4830 (N_4830,N_3955,N_4154);
or U4831 (N_4831,N_4455,N_4041);
and U4832 (N_4832,N_4313,N_4339);
xnor U4833 (N_4833,N_3621,N_3880);
xor U4834 (N_4834,N_3990,N_4059);
nand U4835 (N_4835,N_4225,N_4170);
nor U4836 (N_4836,N_3727,N_3603);
or U4837 (N_4837,N_3356,N_3558);
nand U4838 (N_4838,N_4437,N_3213);
and U4839 (N_4839,N_4342,N_3686);
or U4840 (N_4840,N_3605,N_3743);
xnor U4841 (N_4841,N_3901,N_4260);
xnor U4842 (N_4842,N_3079,N_4163);
nor U4843 (N_4843,N_3784,N_3641);
and U4844 (N_4844,N_3864,N_3266);
nor U4845 (N_4845,N_4449,N_4344);
xor U4846 (N_4846,N_4316,N_4426);
or U4847 (N_4847,N_3076,N_4138);
nor U4848 (N_4848,N_3170,N_3335);
xor U4849 (N_4849,N_4293,N_3292);
nor U4850 (N_4850,N_3563,N_3882);
and U4851 (N_4851,N_3326,N_3724);
nor U4852 (N_4852,N_3897,N_3439);
or U4853 (N_4853,N_3989,N_3866);
xnor U4854 (N_4854,N_4197,N_4062);
nor U4855 (N_4855,N_3254,N_4074);
or U4856 (N_4856,N_4204,N_4220);
or U4857 (N_4857,N_3483,N_3273);
xnor U4858 (N_4858,N_3274,N_4497);
xnor U4859 (N_4859,N_3720,N_4020);
nand U4860 (N_4860,N_3414,N_3548);
and U4861 (N_4861,N_3410,N_3475);
xnor U4862 (N_4862,N_3777,N_3012);
nor U4863 (N_4863,N_3590,N_4387);
xnor U4864 (N_4864,N_4253,N_3046);
nor U4865 (N_4865,N_3364,N_4432);
or U4866 (N_4866,N_4488,N_3824);
nor U4867 (N_4867,N_3825,N_3409);
nand U4868 (N_4868,N_4177,N_4297);
and U4869 (N_4869,N_3459,N_4072);
nor U4870 (N_4870,N_3271,N_4208);
and U4871 (N_4871,N_4268,N_4319);
or U4872 (N_4872,N_4026,N_4056);
xnor U4873 (N_4873,N_4382,N_3121);
nand U4874 (N_4874,N_4255,N_4053);
or U4875 (N_4875,N_4104,N_3109);
and U4876 (N_4876,N_4372,N_3229);
or U4877 (N_4877,N_3016,N_3239);
xnor U4878 (N_4878,N_3957,N_3131);
xnor U4879 (N_4879,N_4257,N_3150);
xor U4880 (N_4880,N_3948,N_3919);
or U4881 (N_4881,N_4281,N_3891);
and U4882 (N_4882,N_4093,N_4202);
nor U4883 (N_4883,N_3195,N_4226);
nand U4884 (N_4884,N_3038,N_4438);
nor U4885 (N_4885,N_3049,N_4148);
nand U4886 (N_4886,N_3725,N_4338);
nand U4887 (N_4887,N_4047,N_4472);
or U4888 (N_4888,N_4046,N_3489);
and U4889 (N_4889,N_3532,N_3582);
nor U4890 (N_4890,N_3774,N_4213);
or U4891 (N_4891,N_3848,N_3533);
or U4892 (N_4892,N_3037,N_3716);
and U4893 (N_4893,N_3505,N_3861);
or U4894 (N_4894,N_3345,N_3938);
nor U4895 (N_4895,N_4235,N_4040);
nand U4896 (N_4896,N_4334,N_3307);
and U4897 (N_4897,N_4152,N_3760);
nand U4898 (N_4898,N_3606,N_3073);
nor U4899 (N_4899,N_3635,N_3412);
nor U4900 (N_4900,N_3827,N_4192);
nand U4901 (N_4901,N_3869,N_3761);
nand U4902 (N_4902,N_3775,N_3253);
nand U4903 (N_4903,N_3802,N_3653);
or U4904 (N_4904,N_4106,N_4218);
xor U4905 (N_4905,N_4211,N_3980);
or U4906 (N_4906,N_4205,N_3797);
or U4907 (N_4907,N_3969,N_4122);
xnor U4908 (N_4908,N_3250,N_3035);
or U4909 (N_4909,N_4023,N_4347);
nand U4910 (N_4910,N_3004,N_3804);
and U4911 (N_4911,N_3764,N_3544);
and U4912 (N_4912,N_3282,N_3958);
nand U4913 (N_4913,N_3625,N_3246);
nor U4914 (N_4914,N_4071,N_4123);
and U4915 (N_4915,N_3992,N_3390);
nor U4916 (N_4916,N_3041,N_4423);
or U4917 (N_4917,N_3281,N_4027);
and U4918 (N_4918,N_4245,N_3456);
and U4919 (N_4919,N_3029,N_3732);
or U4920 (N_4920,N_4270,N_3615);
xor U4921 (N_4921,N_3196,N_3217);
and U4922 (N_4922,N_3554,N_3224);
nor U4923 (N_4923,N_3636,N_4049);
nor U4924 (N_4924,N_3646,N_4162);
or U4925 (N_4925,N_3114,N_3528);
xor U4926 (N_4926,N_3106,N_3343);
nand U4927 (N_4927,N_3166,N_3609);
and U4928 (N_4928,N_4079,N_3521);
nor U4929 (N_4929,N_3160,N_3394);
or U4930 (N_4930,N_4429,N_3923);
and U4931 (N_4931,N_3712,N_4325);
nand U4932 (N_4932,N_3135,N_3054);
or U4933 (N_4933,N_3579,N_4473);
or U4934 (N_4934,N_3645,N_3678);
and U4935 (N_4935,N_3707,N_3809);
nor U4936 (N_4936,N_3242,N_4479);
nand U4937 (N_4937,N_3918,N_4175);
or U4938 (N_4938,N_3999,N_4036);
and U4939 (N_4939,N_4003,N_3187);
nor U4940 (N_4940,N_3863,N_3626);
nand U4941 (N_4941,N_3182,N_3726);
and U4942 (N_4942,N_4459,N_4291);
xor U4943 (N_4943,N_4096,N_4384);
nand U4944 (N_4944,N_3585,N_3829);
and U4945 (N_4945,N_4195,N_4055);
or U4946 (N_4946,N_3151,N_4077);
nor U4947 (N_4947,N_3181,N_4360);
nor U4948 (N_4948,N_3714,N_3120);
or U4949 (N_4949,N_3277,N_3416);
and U4950 (N_4950,N_3244,N_4336);
or U4951 (N_4951,N_3939,N_3627);
and U4952 (N_4952,N_3175,N_3382);
nand U4953 (N_4953,N_4309,N_3936);
nor U4954 (N_4954,N_3767,N_4390);
or U4955 (N_4955,N_3011,N_3460);
nor U4956 (N_4956,N_3487,N_4136);
xnor U4957 (N_4957,N_3070,N_3194);
nand U4958 (N_4958,N_3950,N_3867);
nor U4959 (N_4959,N_3498,N_4448);
and U4960 (N_4960,N_3061,N_3374);
xor U4961 (N_4961,N_4267,N_3101);
and U4962 (N_4962,N_3221,N_3684);
or U4963 (N_4963,N_3667,N_4099);
and U4964 (N_4964,N_4286,N_3852);
nand U4965 (N_4965,N_3303,N_3841);
or U4966 (N_4966,N_4159,N_3644);
nand U4967 (N_4967,N_3769,N_3222);
nand U4968 (N_4968,N_3033,N_3252);
or U4969 (N_4969,N_4444,N_3642);
and U4970 (N_4970,N_4010,N_3457);
and U4971 (N_4971,N_3782,N_3699);
nand U4972 (N_4972,N_3358,N_3008);
xnor U4973 (N_4973,N_3972,N_4318);
nor U4974 (N_4974,N_4440,N_3328);
and U4975 (N_4975,N_3839,N_3503);
xnor U4976 (N_4976,N_4402,N_3566);
and U4977 (N_4977,N_4396,N_4017);
nor U4978 (N_4978,N_3383,N_4107);
and U4979 (N_4979,N_3624,N_3740);
xnor U4980 (N_4980,N_3578,N_4480);
and U4981 (N_4981,N_3000,N_3176);
and U4982 (N_4982,N_4452,N_3875);
nand U4983 (N_4983,N_3530,N_4274);
nor U4984 (N_4984,N_4150,N_3402);
and U4985 (N_4985,N_4381,N_3553);
nor U4986 (N_4986,N_4414,N_3706);
and U4987 (N_4987,N_3831,N_3453);
xnor U4988 (N_4988,N_3043,N_3071);
nand U4989 (N_4989,N_3126,N_3411);
and U4990 (N_4990,N_3084,N_4021);
nand U4991 (N_4991,N_3177,N_3006);
or U4992 (N_4992,N_3100,N_3280);
or U4993 (N_4993,N_4359,N_4149);
and U4994 (N_4994,N_3906,N_4035);
nor U4995 (N_4995,N_4075,N_3381);
or U4996 (N_4996,N_3509,N_3647);
nor U4997 (N_4997,N_3342,N_3746);
xor U4998 (N_4998,N_3300,N_3284);
nand U4999 (N_4999,N_3914,N_3700);
or U5000 (N_5000,N_3656,N_3820);
or U5001 (N_5001,N_3979,N_3628);
or U5002 (N_5002,N_4345,N_3596);
xnor U5003 (N_5003,N_3968,N_3355);
nand U5004 (N_5004,N_3230,N_4418);
or U5005 (N_5005,N_3815,N_3591);
xnor U5006 (N_5006,N_3366,N_3237);
and U5007 (N_5007,N_3787,N_3301);
xor U5008 (N_5008,N_3068,N_3778);
nor U5009 (N_5009,N_4001,N_3447);
or U5010 (N_5010,N_3966,N_3812);
and U5011 (N_5011,N_3808,N_3147);
and U5012 (N_5012,N_3870,N_3692);
or U5013 (N_5013,N_3507,N_4037);
and U5014 (N_5014,N_3844,N_3329);
or U5015 (N_5015,N_3728,N_4433);
nand U5016 (N_5016,N_4416,N_4368);
nand U5017 (N_5017,N_3588,N_4135);
and U5018 (N_5018,N_3681,N_4393);
or U5019 (N_5019,N_3666,N_3598);
xor U5020 (N_5020,N_3190,N_4328);
nand U5021 (N_5021,N_3086,N_3541);
nor U5022 (N_5022,N_3435,N_4012);
nor U5023 (N_5023,N_3943,N_3180);
or U5024 (N_5024,N_4141,N_4424);
nand U5025 (N_5025,N_3310,N_3005);
or U5026 (N_5026,N_3987,N_4227);
or U5027 (N_5027,N_3896,N_3496);
and U5028 (N_5028,N_4442,N_3407);
and U5029 (N_5029,N_3080,N_3632);
or U5030 (N_5030,N_4029,N_3576);
xor U5031 (N_5031,N_3971,N_3248);
xor U5032 (N_5032,N_3872,N_3389);
nand U5033 (N_5033,N_3322,N_3623);
or U5034 (N_5034,N_3391,N_3075);
nand U5035 (N_5035,N_4406,N_3066);
and U5036 (N_5036,N_3857,N_3484);
nor U5037 (N_5037,N_4445,N_3065);
and U5038 (N_5038,N_3146,N_3543);
and U5039 (N_5039,N_3377,N_3286);
nor U5040 (N_5040,N_3275,N_3473);
and U5041 (N_5041,N_3630,N_4161);
or U5042 (N_5042,N_3611,N_4264);
nand U5043 (N_5043,N_3003,N_3072);
or U5044 (N_5044,N_3513,N_3261);
nor U5045 (N_5045,N_4057,N_3735);
nor U5046 (N_5046,N_3564,N_3032);
and U5047 (N_5047,N_3556,N_3691);
nor U5048 (N_5048,N_3589,N_3099);
nor U5049 (N_5049,N_3651,N_3469);
nor U5050 (N_5050,N_3652,N_3234);
nand U5051 (N_5051,N_4467,N_3796);
nor U5052 (N_5052,N_3186,N_3482);
nand U5053 (N_5053,N_4052,N_3327);
nor U5054 (N_5054,N_3932,N_3731);
nor U5055 (N_5055,N_3688,N_4147);
nand U5056 (N_5056,N_3396,N_3680);
nand U5057 (N_5057,N_3436,N_4142);
and U5058 (N_5058,N_4466,N_3949);
nand U5059 (N_5059,N_3631,N_3765);
nand U5060 (N_5060,N_3508,N_3616);
or U5061 (N_5061,N_3903,N_3001);
nor U5062 (N_5062,N_3964,N_4435);
nor U5063 (N_5063,N_3752,N_4028);
nand U5064 (N_5064,N_4343,N_3862);
nor U5065 (N_5065,N_4379,N_4143);
nor U5066 (N_5066,N_3698,N_3832);
nor U5067 (N_5067,N_3110,N_4060);
and U5068 (N_5068,N_3594,N_3894);
nand U5069 (N_5069,N_4491,N_3828);
and U5070 (N_5070,N_3497,N_4465);
and U5071 (N_5071,N_4380,N_3144);
or U5072 (N_5072,N_3129,N_4400);
nand U5073 (N_5073,N_3984,N_3022);
xnor U5074 (N_5074,N_3659,N_3569);
xnor U5075 (N_5075,N_3710,N_3887);
or U5076 (N_5076,N_4399,N_3040);
nor U5077 (N_5077,N_3749,N_4362);
nor U5078 (N_5078,N_4032,N_3397);
and U5079 (N_5079,N_4212,N_3059);
or U5080 (N_5080,N_3689,N_3458);
or U5081 (N_5081,N_3648,N_3023);
nor U5082 (N_5082,N_3568,N_3845);
or U5083 (N_5083,N_3294,N_3904);
and U5084 (N_5084,N_3956,N_3215);
and U5085 (N_5085,N_4113,N_3790);
and U5086 (N_5086,N_3909,N_4383);
or U5087 (N_5087,N_4168,N_3027);
xnor U5088 (N_5088,N_3523,N_3803);
and U5089 (N_5089,N_3420,N_4006);
nand U5090 (N_5090,N_3709,N_4259);
nor U5091 (N_5091,N_4324,N_3696);
and U5092 (N_5092,N_3438,N_3915);
nor U5093 (N_5093,N_3184,N_3567);
nand U5094 (N_5094,N_3963,N_3424);
xor U5095 (N_5095,N_3905,N_4484);
and U5096 (N_5096,N_4004,N_4108);
or U5097 (N_5097,N_3773,N_4468);
nor U5098 (N_5098,N_4420,N_3095);
nand U5099 (N_5099,N_3318,N_3325);
nand U5100 (N_5100,N_3268,N_3791);
xor U5101 (N_5101,N_3975,N_4413);
nand U5102 (N_5102,N_4237,N_4410);
or U5103 (N_5103,N_3055,N_3077);
nor U5104 (N_5104,N_3592,N_3258);
and U5105 (N_5105,N_3451,N_3516);
nand U5106 (N_5106,N_4229,N_3304);
and U5107 (N_5107,N_4190,N_4222);
nor U5108 (N_5108,N_3306,N_3742);
or U5109 (N_5109,N_3514,N_4167);
or U5110 (N_5110,N_4496,N_3305);
nor U5111 (N_5111,N_4292,N_3490);
nor U5112 (N_5112,N_4463,N_4214);
and U5113 (N_5113,N_3771,N_3047);
nor U5114 (N_5114,N_4434,N_4300);
nor U5115 (N_5115,N_3974,N_3308);
xnor U5116 (N_5116,N_3801,N_3317);
xor U5117 (N_5117,N_4453,N_3873);
nor U5118 (N_5118,N_3633,N_4241);
nand U5119 (N_5119,N_3634,N_4323);
nand U5120 (N_5120,N_3737,N_4058);
and U5121 (N_5121,N_4262,N_3437);
or U5122 (N_5122,N_3103,N_4417);
or U5123 (N_5123,N_4250,N_3087);
or U5124 (N_5124,N_4371,N_4051);
and U5125 (N_5125,N_3478,N_4490);
or U5126 (N_5126,N_3074,N_4403);
nand U5127 (N_5127,N_3650,N_4084);
nand U5128 (N_5128,N_3297,N_3427);
or U5129 (N_5129,N_4008,N_3026);
and U5130 (N_5130,N_3085,N_3211);
and U5131 (N_5131,N_4240,N_3783);
nand U5132 (N_5132,N_3917,N_3134);
nand U5133 (N_5133,N_3485,N_3117);
nor U5134 (N_5134,N_3155,N_3662);
nand U5135 (N_5135,N_4069,N_3602);
nand U5136 (N_5136,N_3333,N_3467);
xnor U5137 (N_5137,N_3638,N_3440);
nor U5138 (N_5138,N_3191,N_3442);
nand U5139 (N_5139,N_3312,N_3994);
nand U5140 (N_5140,N_3157,N_4153);
nor U5141 (N_5141,N_3572,N_4242);
or U5142 (N_5142,N_4320,N_3455);
nand U5143 (N_5143,N_4045,N_3141);
nand U5144 (N_5144,N_3930,N_4158);
or U5145 (N_5145,N_4289,N_4354);
or U5146 (N_5146,N_3048,N_3745);
or U5147 (N_5147,N_3908,N_4389);
or U5148 (N_5148,N_3403,N_4302);
or U5149 (N_5149,N_4263,N_4194);
or U5150 (N_5150,N_3811,N_3722);
and U5151 (N_5151,N_3739,N_4474);
nand U5152 (N_5152,N_3486,N_3683);
nor U5153 (N_5153,N_4156,N_4129);
nor U5154 (N_5154,N_3448,N_4042);
nand U5155 (N_5155,N_4494,N_4188);
nand U5156 (N_5156,N_3466,N_4092);
or U5157 (N_5157,N_4246,N_3288);
or U5158 (N_5158,N_4160,N_4272);
nand U5159 (N_5159,N_4183,N_3053);
and U5160 (N_5160,N_3208,N_3264);
and U5161 (N_5161,N_3007,N_3593);
and U5162 (N_5162,N_3081,N_3986);
nand U5163 (N_5163,N_4487,N_3156);
xnor U5164 (N_5164,N_3679,N_3098);
and U5165 (N_5165,N_4460,N_3520);
or U5166 (N_5166,N_3444,N_4125);
and U5167 (N_5167,N_3491,N_4254);
and U5168 (N_5168,N_3555,N_3524);
nand U5169 (N_5169,N_3583,N_3565);
nor U5170 (N_5170,N_3378,N_4485);
nand U5171 (N_5171,N_3618,N_3418);
nand U5172 (N_5172,N_4296,N_3529);
nor U5173 (N_5173,N_3030,N_3476);
nand U5174 (N_5174,N_3934,N_3270);
nor U5175 (N_5175,N_3338,N_3014);
nor U5176 (N_5176,N_3082,N_3015);
and U5177 (N_5177,N_4299,N_3549);
nand U5178 (N_5178,N_3462,N_3042);
and U5179 (N_5179,N_3392,N_3708);
or U5180 (N_5180,N_4483,N_3501);
nor U5181 (N_5181,N_3810,N_3060);
xnor U5182 (N_5182,N_3840,N_3890);
nor U5183 (N_5183,N_3218,N_4044);
xnor U5184 (N_5184,N_3910,N_3063);
nand U5185 (N_5185,N_3321,N_3464);
nand U5186 (N_5186,N_3149,N_4287);
and U5187 (N_5187,N_3494,N_3481);
nand U5188 (N_5188,N_4314,N_3734);
and U5189 (N_5189,N_4492,N_4331);
nand U5190 (N_5190,N_3786,N_3112);
nand U5191 (N_5191,N_3359,N_3365);
or U5192 (N_5192,N_3922,N_3245);
and U5193 (N_5193,N_3226,N_4358);
and U5194 (N_5194,N_3232,N_4111);
and U5195 (N_5195,N_4189,N_4481);
and U5196 (N_5196,N_4394,N_3093);
nor U5197 (N_5197,N_3763,N_3379);
and U5198 (N_5198,N_3423,N_4033);
nor U5199 (N_5199,N_3289,N_3836);
xor U5200 (N_5200,N_3525,N_3800);
nor U5201 (N_5201,N_3617,N_4238);
and U5202 (N_5202,N_4098,N_3296);
and U5203 (N_5203,N_4369,N_3132);
or U5204 (N_5204,N_3951,N_3965);
or U5205 (N_5205,N_3262,N_3747);
nand U5206 (N_5206,N_4105,N_4443);
xnor U5207 (N_5207,N_3518,N_4015);
and U5208 (N_5208,N_4184,N_3798);
or U5209 (N_5209,N_4151,N_3717);
nor U5210 (N_5210,N_3480,N_3212);
and U5211 (N_5211,N_3941,N_4145);
nand U5212 (N_5212,N_3202,N_3522);
nand U5213 (N_5213,N_4178,N_3441);
nor U5214 (N_5214,N_3546,N_3421);
and U5215 (N_5215,N_4114,N_3818);
and U5216 (N_5216,N_4013,N_4376);
xnor U5217 (N_5217,N_4120,N_3886);
nor U5218 (N_5218,N_3405,N_3025);
nor U5219 (N_5219,N_3089,N_3452);
xnor U5220 (N_5220,N_3608,N_3293);
nor U5221 (N_5221,N_3474,N_4134);
nand U5222 (N_5222,N_4127,N_4265);
nor U5223 (N_5223,N_3584,N_3315);
and U5224 (N_5224,N_4230,N_3537);
and U5225 (N_5225,N_4356,N_3946);
and U5226 (N_5226,N_3267,N_3855);
nor U5227 (N_5227,N_3580,N_3982);
or U5228 (N_5228,N_3545,N_3944);
nor U5229 (N_5229,N_3738,N_3766);
and U5230 (N_5230,N_3776,N_3269);
and U5231 (N_5231,N_3736,N_3762);
or U5232 (N_5232,N_3375,N_4078);
xnor U5233 (N_5233,N_4070,N_3888);
nand U5234 (N_5234,N_4076,N_3595);
and U5235 (N_5235,N_3428,N_3929);
and U5236 (N_5236,N_4201,N_3997);
and U5237 (N_5237,N_3967,N_3203);
or U5238 (N_5238,N_3241,N_3920);
and U5239 (N_5239,N_4011,N_3586);
or U5240 (N_5240,N_4303,N_4377);
and U5241 (N_5241,N_3198,N_3145);
or U5242 (N_5242,N_3272,N_4130);
nand U5243 (N_5243,N_3124,N_4244);
nand U5244 (N_5244,N_3278,N_3898);
nand U5245 (N_5245,N_4415,N_3050);
and U5246 (N_5246,N_3018,N_4239);
or U5247 (N_5247,N_3985,N_4321);
nor U5248 (N_5248,N_4095,N_3675);
nand U5249 (N_5249,N_4307,N_4478);
nand U5250 (N_5250,N_3588,N_4128);
or U5251 (N_5251,N_3343,N_4446);
and U5252 (N_5252,N_3904,N_3733);
or U5253 (N_5253,N_4002,N_3060);
nand U5254 (N_5254,N_4152,N_4302);
nor U5255 (N_5255,N_3696,N_3421);
nor U5256 (N_5256,N_4059,N_3245);
or U5257 (N_5257,N_3159,N_3285);
xnor U5258 (N_5258,N_3938,N_3163);
nor U5259 (N_5259,N_4227,N_4324);
nor U5260 (N_5260,N_3994,N_3688);
nor U5261 (N_5261,N_3689,N_3974);
and U5262 (N_5262,N_3909,N_3251);
and U5263 (N_5263,N_4263,N_3188);
and U5264 (N_5264,N_3711,N_3513);
nand U5265 (N_5265,N_3761,N_4233);
and U5266 (N_5266,N_3249,N_3845);
nor U5267 (N_5267,N_3919,N_3748);
nand U5268 (N_5268,N_3658,N_3320);
nand U5269 (N_5269,N_4354,N_4073);
xnor U5270 (N_5270,N_4233,N_3465);
or U5271 (N_5271,N_3697,N_3906);
and U5272 (N_5272,N_3366,N_3571);
or U5273 (N_5273,N_3747,N_4121);
xor U5274 (N_5274,N_4478,N_3020);
or U5275 (N_5275,N_3198,N_3690);
or U5276 (N_5276,N_3626,N_3091);
or U5277 (N_5277,N_3333,N_3448);
nand U5278 (N_5278,N_3659,N_3561);
and U5279 (N_5279,N_3780,N_4328);
and U5280 (N_5280,N_3947,N_4124);
nor U5281 (N_5281,N_3125,N_3292);
and U5282 (N_5282,N_3771,N_3429);
nand U5283 (N_5283,N_3687,N_3094);
or U5284 (N_5284,N_3728,N_3176);
and U5285 (N_5285,N_3899,N_3313);
xnor U5286 (N_5286,N_3812,N_3866);
or U5287 (N_5287,N_3912,N_3080);
nand U5288 (N_5288,N_3296,N_3258);
nor U5289 (N_5289,N_3409,N_4397);
nand U5290 (N_5290,N_3301,N_4469);
nand U5291 (N_5291,N_3007,N_3664);
nand U5292 (N_5292,N_4418,N_3215);
nand U5293 (N_5293,N_3204,N_3076);
nor U5294 (N_5294,N_3618,N_4214);
and U5295 (N_5295,N_3206,N_4212);
nor U5296 (N_5296,N_3934,N_4136);
nor U5297 (N_5297,N_3343,N_3125);
nor U5298 (N_5298,N_3473,N_3484);
or U5299 (N_5299,N_4145,N_3363);
and U5300 (N_5300,N_4076,N_3770);
and U5301 (N_5301,N_3355,N_4367);
nor U5302 (N_5302,N_3416,N_4073);
nor U5303 (N_5303,N_4269,N_4447);
nor U5304 (N_5304,N_3970,N_4026);
nand U5305 (N_5305,N_3020,N_3159);
or U5306 (N_5306,N_4023,N_3483);
and U5307 (N_5307,N_4044,N_3241);
nand U5308 (N_5308,N_3902,N_4457);
nor U5309 (N_5309,N_3437,N_3820);
nor U5310 (N_5310,N_3689,N_4155);
nand U5311 (N_5311,N_3678,N_3743);
nand U5312 (N_5312,N_3674,N_3432);
and U5313 (N_5313,N_4313,N_3763);
or U5314 (N_5314,N_4211,N_3135);
nand U5315 (N_5315,N_3294,N_3429);
and U5316 (N_5316,N_4442,N_3854);
xnor U5317 (N_5317,N_3337,N_3197);
and U5318 (N_5318,N_3490,N_3480);
xnor U5319 (N_5319,N_3258,N_4321);
xor U5320 (N_5320,N_4283,N_3605);
nor U5321 (N_5321,N_3953,N_4311);
nand U5322 (N_5322,N_4028,N_3939);
nand U5323 (N_5323,N_4456,N_3742);
or U5324 (N_5324,N_3901,N_3776);
xnor U5325 (N_5325,N_4270,N_3516);
nor U5326 (N_5326,N_3773,N_4295);
and U5327 (N_5327,N_3127,N_3546);
nor U5328 (N_5328,N_4480,N_3790);
and U5329 (N_5329,N_3616,N_3342);
or U5330 (N_5330,N_3813,N_4381);
nand U5331 (N_5331,N_3655,N_3593);
nor U5332 (N_5332,N_3725,N_4099);
or U5333 (N_5333,N_3568,N_3706);
nor U5334 (N_5334,N_3684,N_4113);
and U5335 (N_5335,N_3607,N_3116);
nor U5336 (N_5336,N_3001,N_3940);
nand U5337 (N_5337,N_3080,N_3626);
xor U5338 (N_5338,N_3575,N_3552);
nand U5339 (N_5339,N_4129,N_3176);
nor U5340 (N_5340,N_4440,N_4274);
xor U5341 (N_5341,N_4220,N_4028);
xor U5342 (N_5342,N_3272,N_3694);
nor U5343 (N_5343,N_3640,N_4256);
nand U5344 (N_5344,N_3803,N_3696);
and U5345 (N_5345,N_3488,N_4080);
nand U5346 (N_5346,N_3265,N_3370);
and U5347 (N_5347,N_3623,N_3288);
and U5348 (N_5348,N_3343,N_4473);
nand U5349 (N_5349,N_4173,N_4196);
nor U5350 (N_5350,N_3760,N_4124);
and U5351 (N_5351,N_3956,N_3339);
nor U5352 (N_5352,N_3990,N_3781);
xnor U5353 (N_5353,N_3551,N_4486);
or U5354 (N_5354,N_3734,N_4436);
or U5355 (N_5355,N_3512,N_3219);
nand U5356 (N_5356,N_4072,N_3954);
nand U5357 (N_5357,N_3010,N_3217);
and U5358 (N_5358,N_3162,N_3658);
nand U5359 (N_5359,N_3809,N_3335);
or U5360 (N_5360,N_4066,N_3314);
nor U5361 (N_5361,N_4307,N_4405);
xor U5362 (N_5362,N_3636,N_3454);
nand U5363 (N_5363,N_3241,N_3724);
xnor U5364 (N_5364,N_4220,N_4364);
or U5365 (N_5365,N_4393,N_3598);
and U5366 (N_5366,N_3524,N_3498);
or U5367 (N_5367,N_3330,N_4150);
or U5368 (N_5368,N_4288,N_3017);
or U5369 (N_5369,N_3268,N_3332);
or U5370 (N_5370,N_3793,N_4296);
and U5371 (N_5371,N_3243,N_3141);
and U5372 (N_5372,N_3854,N_3162);
nand U5373 (N_5373,N_4494,N_3419);
nand U5374 (N_5374,N_3821,N_4345);
nor U5375 (N_5375,N_3575,N_3456);
and U5376 (N_5376,N_3323,N_3100);
or U5377 (N_5377,N_3251,N_3996);
nand U5378 (N_5378,N_3435,N_4363);
or U5379 (N_5379,N_4001,N_3272);
or U5380 (N_5380,N_3963,N_3142);
nor U5381 (N_5381,N_4374,N_3225);
and U5382 (N_5382,N_4055,N_4228);
and U5383 (N_5383,N_4413,N_3192);
and U5384 (N_5384,N_3680,N_3703);
and U5385 (N_5385,N_3066,N_3301);
nor U5386 (N_5386,N_3366,N_4415);
nand U5387 (N_5387,N_3588,N_4399);
nand U5388 (N_5388,N_3807,N_3623);
and U5389 (N_5389,N_4245,N_4215);
and U5390 (N_5390,N_4039,N_3203);
xnor U5391 (N_5391,N_3465,N_3379);
nor U5392 (N_5392,N_3957,N_3136);
and U5393 (N_5393,N_3530,N_3178);
or U5394 (N_5394,N_3093,N_3201);
and U5395 (N_5395,N_3719,N_3714);
and U5396 (N_5396,N_3709,N_3501);
nand U5397 (N_5397,N_4215,N_4066);
nand U5398 (N_5398,N_3206,N_3928);
nor U5399 (N_5399,N_4465,N_3760);
nor U5400 (N_5400,N_4173,N_4495);
nor U5401 (N_5401,N_3976,N_4222);
nor U5402 (N_5402,N_4317,N_3570);
nand U5403 (N_5403,N_4059,N_4302);
nor U5404 (N_5404,N_4228,N_3384);
nor U5405 (N_5405,N_3491,N_4420);
and U5406 (N_5406,N_4083,N_4281);
nor U5407 (N_5407,N_4178,N_3356);
and U5408 (N_5408,N_3991,N_3254);
or U5409 (N_5409,N_4188,N_3365);
nand U5410 (N_5410,N_3046,N_3436);
nand U5411 (N_5411,N_3376,N_3357);
nand U5412 (N_5412,N_4237,N_4159);
and U5413 (N_5413,N_3466,N_3471);
nand U5414 (N_5414,N_3663,N_3531);
nor U5415 (N_5415,N_3489,N_4143);
or U5416 (N_5416,N_4141,N_3803);
or U5417 (N_5417,N_3709,N_3088);
and U5418 (N_5418,N_4371,N_3774);
nor U5419 (N_5419,N_4261,N_4476);
nand U5420 (N_5420,N_4205,N_3056);
or U5421 (N_5421,N_3753,N_3768);
nor U5422 (N_5422,N_4053,N_3948);
or U5423 (N_5423,N_4113,N_3493);
nand U5424 (N_5424,N_4306,N_3930);
and U5425 (N_5425,N_3257,N_3643);
nand U5426 (N_5426,N_4281,N_4372);
or U5427 (N_5427,N_3348,N_3169);
and U5428 (N_5428,N_4121,N_4010);
nand U5429 (N_5429,N_3619,N_3342);
or U5430 (N_5430,N_3178,N_3951);
and U5431 (N_5431,N_3628,N_3527);
xor U5432 (N_5432,N_4293,N_4328);
and U5433 (N_5433,N_4361,N_3985);
nand U5434 (N_5434,N_4195,N_3612);
xor U5435 (N_5435,N_3784,N_3903);
nor U5436 (N_5436,N_4254,N_3831);
xor U5437 (N_5437,N_4466,N_3259);
and U5438 (N_5438,N_4289,N_3914);
and U5439 (N_5439,N_4026,N_4269);
nand U5440 (N_5440,N_3036,N_3927);
and U5441 (N_5441,N_4102,N_3824);
nor U5442 (N_5442,N_3471,N_3839);
nor U5443 (N_5443,N_3871,N_4409);
nand U5444 (N_5444,N_3806,N_4054);
or U5445 (N_5445,N_3854,N_4472);
nor U5446 (N_5446,N_4317,N_4411);
and U5447 (N_5447,N_4461,N_3935);
xnor U5448 (N_5448,N_3776,N_3227);
nand U5449 (N_5449,N_4349,N_3757);
nor U5450 (N_5450,N_3872,N_3290);
or U5451 (N_5451,N_3659,N_4149);
xnor U5452 (N_5452,N_3011,N_4209);
or U5453 (N_5453,N_3179,N_3734);
nor U5454 (N_5454,N_4245,N_4144);
and U5455 (N_5455,N_4405,N_3968);
nor U5456 (N_5456,N_3706,N_3180);
nor U5457 (N_5457,N_4082,N_3063);
nand U5458 (N_5458,N_3147,N_4206);
nor U5459 (N_5459,N_3854,N_3458);
nor U5460 (N_5460,N_3115,N_3059);
xnor U5461 (N_5461,N_3340,N_3789);
or U5462 (N_5462,N_4287,N_3593);
nor U5463 (N_5463,N_3563,N_3343);
nand U5464 (N_5464,N_4445,N_3504);
or U5465 (N_5465,N_3337,N_4414);
nand U5466 (N_5466,N_3316,N_4327);
nand U5467 (N_5467,N_3386,N_3788);
nor U5468 (N_5468,N_3824,N_3593);
nand U5469 (N_5469,N_3942,N_3936);
or U5470 (N_5470,N_4161,N_3872);
and U5471 (N_5471,N_4069,N_3616);
nor U5472 (N_5472,N_4432,N_3519);
and U5473 (N_5473,N_4156,N_3250);
nor U5474 (N_5474,N_3945,N_3149);
xor U5475 (N_5475,N_3237,N_3863);
nand U5476 (N_5476,N_4362,N_4481);
nand U5477 (N_5477,N_3203,N_4312);
nand U5478 (N_5478,N_4134,N_3346);
or U5479 (N_5479,N_3136,N_4407);
or U5480 (N_5480,N_3830,N_3768);
and U5481 (N_5481,N_4360,N_3786);
nor U5482 (N_5482,N_3717,N_3127);
nand U5483 (N_5483,N_4366,N_3447);
nor U5484 (N_5484,N_3474,N_4304);
xnor U5485 (N_5485,N_3131,N_3597);
or U5486 (N_5486,N_4264,N_3257);
and U5487 (N_5487,N_3627,N_3294);
nor U5488 (N_5488,N_3280,N_3917);
or U5489 (N_5489,N_3477,N_3266);
or U5490 (N_5490,N_3269,N_3430);
nand U5491 (N_5491,N_3080,N_4189);
and U5492 (N_5492,N_3875,N_3761);
xor U5493 (N_5493,N_3637,N_4010);
xnor U5494 (N_5494,N_4349,N_3635);
or U5495 (N_5495,N_3569,N_3856);
nor U5496 (N_5496,N_4443,N_3413);
nand U5497 (N_5497,N_3455,N_4458);
or U5498 (N_5498,N_4483,N_4130);
nand U5499 (N_5499,N_3500,N_4262);
nand U5500 (N_5500,N_3163,N_4480);
or U5501 (N_5501,N_4444,N_4268);
and U5502 (N_5502,N_4410,N_3445);
nor U5503 (N_5503,N_3994,N_4336);
xnor U5504 (N_5504,N_4346,N_3776);
nor U5505 (N_5505,N_3222,N_3865);
and U5506 (N_5506,N_3337,N_3795);
and U5507 (N_5507,N_4047,N_4497);
or U5508 (N_5508,N_3538,N_3101);
nor U5509 (N_5509,N_4221,N_3209);
xnor U5510 (N_5510,N_4104,N_3769);
nand U5511 (N_5511,N_4203,N_4448);
and U5512 (N_5512,N_3209,N_4331);
nand U5513 (N_5513,N_3767,N_3144);
nand U5514 (N_5514,N_4415,N_3929);
and U5515 (N_5515,N_4362,N_3024);
or U5516 (N_5516,N_3701,N_3557);
and U5517 (N_5517,N_3336,N_3254);
nor U5518 (N_5518,N_3221,N_3510);
xor U5519 (N_5519,N_3731,N_4206);
nor U5520 (N_5520,N_3692,N_3196);
xnor U5521 (N_5521,N_4369,N_3821);
nand U5522 (N_5522,N_4009,N_4279);
nand U5523 (N_5523,N_3521,N_3118);
nor U5524 (N_5524,N_3614,N_3878);
and U5525 (N_5525,N_3958,N_3871);
and U5526 (N_5526,N_4402,N_4015);
or U5527 (N_5527,N_3813,N_3687);
nor U5528 (N_5528,N_4030,N_3325);
nand U5529 (N_5529,N_3181,N_4331);
and U5530 (N_5530,N_3459,N_3421);
or U5531 (N_5531,N_3520,N_4045);
nor U5532 (N_5532,N_3254,N_3782);
nand U5533 (N_5533,N_3699,N_4444);
or U5534 (N_5534,N_3594,N_3340);
or U5535 (N_5535,N_3264,N_4300);
nor U5536 (N_5536,N_3376,N_3678);
nor U5537 (N_5537,N_3536,N_3869);
nand U5538 (N_5538,N_4374,N_4412);
or U5539 (N_5539,N_3858,N_3498);
or U5540 (N_5540,N_3135,N_4194);
xor U5541 (N_5541,N_3267,N_3495);
or U5542 (N_5542,N_3067,N_4284);
and U5543 (N_5543,N_3812,N_4032);
xnor U5544 (N_5544,N_3191,N_3348);
or U5545 (N_5545,N_4113,N_4099);
nand U5546 (N_5546,N_4241,N_3434);
or U5547 (N_5547,N_3278,N_4023);
or U5548 (N_5548,N_3613,N_3601);
or U5549 (N_5549,N_3796,N_3618);
nor U5550 (N_5550,N_3107,N_3322);
or U5551 (N_5551,N_3731,N_4121);
or U5552 (N_5552,N_3607,N_3821);
or U5553 (N_5553,N_4070,N_3556);
or U5554 (N_5554,N_3816,N_4392);
nor U5555 (N_5555,N_3564,N_3839);
nand U5556 (N_5556,N_3091,N_3557);
and U5557 (N_5557,N_4248,N_4342);
and U5558 (N_5558,N_4322,N_3648);
or U5559 (N_5559,N_3327,N_3967);
and U5560 (N_5560,N_4055,N_3986);
or U5561 (N_5561,N_4197,N_3388);
nor U5562 (N_5562,N_3045,N_4335);
and U5563 (N_5563,N_3257,N_3121);
xnor U5564 (N_5564,N_4490,N_3659);
xor U5565 (N_5565,N_4104,N_4461);
nand U5566 (N_5566,N_3052,N_3973);
or U5567 (N_5567,N_3367,N_3482);
or U5568 (N_5568,N_3454,N_3031);
nor U5569 (N_5569,N_3789,N_3205);
or U5570 (N_5570,N_3272,N_3021);
nor U5571 (N_5571,N_3371,N_3001);
and U5572 (N_5572,N_3357,N_4161);
xnor U5573 (N_5573,N_4237,N_3481);
nor U5574 (N_5574,N_3379,N_3853);
xnor U5575 (N_5575,N_4137,N_4480);
or U5576 (N_5576,N_3985,N_3849);
and U5577 (N_5577,N_3222,N_3350);
or U5578 (N_5578,N_4427,N_3946);
xnor U5579 (N_5579,N_3865,N_3190);
nor U5580 (N_5580,N_3351,N_4135);
nor U5581 (N_5581,N_3305,N_4117);
and U5582 (N_5582,N_4267,N_3615);
and U5583 (N_5583,N_3383,N_3239);
or U5584 (N_5584,N_3057,N_3303);
and U5585 (N_5585,N_3469,N_3043);
nor U5586 (N_5586,N_3158,N_4339);
nor U5587 (N_5587,N_3586,N_3536);
nor U5588 (N_5588,N_4300,N_3234);
and U5589 (N_5589,N_3391,N_4161);
and U5590 (N_5590,N_4433,N_3752);
nor U5591 (N_5591,N_3646,N_3789);
and U5592 (N_5592,N_3892,N_4336);
nor U5593 (N_5593,N_3236,N_3257);
and U5594 (N_5594,N_4464,N_4160);
or U5595 (N_5595,N_3522,N_3127);
nor U5596 (N_5596,N_3208,N_4079);
nor U5597 (N_5597,N_3521,N_3280);
or U5598 (N_5598,N_3259,N_4305);
or U5599 (N_5599,N_4214,N_3786);
or U5600 (N_5600,N_4434,N_3091);
and U5601 (N_5601,N_3429,N_3589);
xor U5602 (N_5602,N_3192,N_3888);
nor U5603 (N_5603,N_4088,N_3747);
nand U5604 (N_5604,N_3225,N_4473);
nor U5605 (N_5605,N_3664,N_3720);
nand U5606 (N_5606,N_3150,N_3386);
nor U5607 (N_5607,N_3904,N_4335);
or U5608 (N_5608,N_3040,N_3760);
and U5609 (N_5609,N_3169,N_3627);
and U5610 (N_5610,N_3193,N_3715);
and U5611 (N_5611,N_4117,N_4378);
nand U5612 (N_5612,N_4315,N_3219);
or U5613 (N_5613,N_3419,N_3056);
xnor U5614 (N_5614,N_3547,N_3929);
and U5615 (N_5615,N_3639,N_3850);
and U5616 (N_5616,N_3759,N_4196);
or U5617 (N_5617,N_3248,N_4389);
nand U5618 (N_5618,N_3066,N_4254);
nand U5619 (N_5619,N_3065,N_4405);
and U5620 (N_5620,N_3016,N_3345);
and U5621 (N_5621,N_3774,N_4172);
or U5622 (N_5622,N_3502,N_4143);
or U5623 (N_5623,N_3038,N_3670);
or U5624 (N_5624,N_3139,N_3142);
nand U5625 (N_5625,N_4225,N_3825);
nor U5626 (N_5626,N_3894,N_4061);
nor U5627 (N_5627,N_3166,N_3485);
xnor U5628 (N_5628,N_3661,N_4039);
and U5629 (N_5629,N_3839,N_4293);
or U5630 (N_5630,N_4218,N_3222);
and U5631 (N_5631,N_3081,N_4379);
nor U5632 (N_5632,N_3974,N_4159);
nor U5633 (N_5633,N_4270,N_3681);
xor U5634 (N_5634,N_3016,N_3412);
xor U5635 (N_5635,N_3285,N_3027);
xor U5636 (N_5636,N_3817,N_4346);
xnor U5637 (N_5637,N_3002,N_4263);
and U5638 (N_5638,N_3125,N_3930);
nand U5639 (N_5639,N_4385,N_4365);
and U5640 (N_5640,N_3995,N_3469);
nor U5641 (N_5641,N_4213,N_4447);
nor U5642 (N_5642,N_4031,N_4186);
and U5643 (N_5643,N_4077,N_4089);
nand U5644 (N_5644,N_3465,N_4032);
xor U5645 (N_5645,N_3044,N_3870);
nand U5646 (N_5646,N_3772,N_3885);
nand U5647 (N_5647,N_4419,N_3703);
or U5648 (N_5648,N_4138,N_3358);
nand U5649 (N_5649,N_3869,N_4069);
nand U5650 (N_5650,N_4491,N_3964);
nor U5651 (N_5651,N_3816,N_3432);
and U5652 (N_5652,N_3015,N_4459);
nor U5653 (N_5653,N_3307,N_3360);
and U5654 (N_5654,N_4389,N_3257);
nor U5655 (N_5655,N_3656,N_3066);
nor U5656 (N_5656,N_4016,N_4082);
xor U5657 (N_5657,N_4086,N_3722);
nor U5658 (N_5658,N_3376,N_3285);
nor U5659 (N_5659,N_3373,N_3145);
or U5660 (N_5660,N_4007,N_4105);
or U5661 (N_5661,N_4425,N_4356);
and U5662 (N_5662,N_3510,N_3984);
nor U5663 (N_5663,N_4027,N_3855);
nor U5664 (N_5664,N_3789,N_3765);
and U5665 (N_5665,N_3219,N_3840);
nor U5666 (N_5666,N_3519,N_3606);
nor U5667 (N_5667,N_3227,N_3476);
nand U5668 (N_5668,N_3076,N_3106);
and U5669 (N_5669,N_3922,N_3605);
and U5670 (N_5670,N_3252,N_3395);
or U5671 (N_5671,N_4232,N_3223);
or U5672 (N_5672,N_4433,N_3128);
nand U5673 (N_5673,N_3922,N_4283);
and U5674 (N_5674,N_3378,N_3957);
and U5675 (N_5675,N_3633,N_3191);
or U5676 (N_5676,N_3962,N_3417);
and U5677 (N_5677,N_3554,N_3129);
or U5678 (N_5678,N_3147,N_3710);
nand U5679 (N_5679,N_3884,N_3745);
or U5680 (N_5680,N_3380,N_4076);
nor U5681 (N_5681,N_3443,N_4403);
and U5682 (N_5682,N_3453,N_4319);
and U5683 (N_5683,N_4136,N_3661);
or U5684 (N_5684,N_3479,N_3939);
nor U5685 (N_5685,N_3551,N_3093);
nor U5686 (N_5686,N_3108,N_3550);
and U5687 (N_5687,N_3602,N_3683);
or U5688 (N_5688,N_4184,N_3281);
or U5689 (N_5689,N_3390,N_3993);
or U5690 (N_5690,N_3859,N_3120);
nand U5691 (N_5691,N_3048,N_4256);
nor U5692 (N_5692,N_3091,N_3285);
and U5693 (N_5693,N_4358,N_3224);
and U5694 (N_5694,N_4427,N_3851);
nand U5695 (N_5695,N_4323,N_3611);
nand U5696 (N_5696,N_3167,N_3963);
nor U5697 (N_5697,N_3763,N_4312);
nand U5698 (N_5698,N_3770,N_3280);
nand U5699 (N_5699,N_3131,N_3009);
nand U5700 (N_5700,N_4287,N_3793);
nor U5701 (N_5701,N_4048,N_4050);
nor U5702 (N_5702,N_4134,N_4294);
and U5703 (N_5703,N_4332,N_4355);
and U5704 (N_5704,N_3037,N_4436);
and U5705 (N_5705,N_3171,N_3161);
xnor U5706 (N_5706,N_3079,N_4412);
nand U5707 (N_5707,N_3393,N_3738);
nand U5708 (N_5708,N_4446,N_3985);
or U5709 (N_5709,N_4165,N_3381);
xnor U5710 (N_5710,N_3048,N_3751);
and U5711 (N_5711,N_4385,N_3996);
and U5712 (N_5712,N_3070,N_4069);
and U5713 (N_5713,N_3833,N_4339);
and U5714 (N_5714,N_3453,N_4104);
nor U5715 (N_5715,N_3675,N_4413);
nand U5716 (N_5716,N_3502,N_4190);
or U5717 (N_5717,N_4489,N_3622);
and U5718 (N_5718,N_3094,N_3221);
nor U5719 (N_5719,N_3815,N_4287);
nand U5720 (N_5720,N_3610,N_3323);
and U5721 (N_5721,N_4151,N_4145);
nor U5722 (N_5722,N_4308,N_3707);
nand U5723 (N_5723,N_3362,N_3657);
or U5724 (N_5724,N_4114,N_3301);
or U5725 (N_5725,N_3756,N_3680);
nor U5726 (N_5726,N_3177,N_3124);
or U5727 (N_5727,N_4166,N_4052);
and U5728 (N_5728,N_3297,N_4390);
nand U5729 (N_5729,N_3765,N_3379);
xnor U5730 (N_5730,N_4143,N_4057);
or U5731 (N_5731,N_3226,N_3897);
and U5732 (N_5732,N_3047,N_4408);
or U5733 (N_5733,N_4416,N_3704);
or U5734 (N_5734,N_4406,N_3523);
or U5735 (N_5735,N_3639,N_3825);
nand U5736 (N_5736,N_3704,N_4383);
or U5737 (N_5737,N_3639,N_3671);
nor U5738 (N_5738,N_3172,N_4311);
nand U5739 (N_5739,N_3108,N_4188);
xnor U5740 (N_5740,N_4158,N_3924);
nand U5741 (N_5741,N_3190,N_4370);
nand U5742 (N_5742,N_4109,N_4006);
nor U5743 (N_5743,N_3946,N_3401);
or U5744 (N_5744,N_3453,N_3872);
and U5745 (N_5745,N_3110,N_3124);
xor U5746 (N_5746,N_3405,N_3429);
nor U5747 (N_5747,N_3172,N_4037);
or U5748 (N_5748,N_3668,N_3005);
and U5749 (N_5749,N_4054,N_3105);
and U5750 (N_5750,N_3828,N_4138);
or U5751 (N_5751,N_4219,N_3748);
nand U5752 (N_5752,N_4461,N_4429);
nand U5753 (N_5753,N_3948,N_3578);
nor U5754 (N_5754,N_4452,N_4183);
or U5755 (N_5755,N_3122,N_3602);
and U5756 (N_5756,N_3852,N_3427);
nor U5757 (N_5757,N_4206,N_4020);
and U5758 (N_5758,N_4197,N_3130);
nand U5759 (N_5759,N_3325,N_3115);
and U5760 (N_5760,N_3457,N_4222);
nand U5761 (N_5761,N_4474,N_3996);
nor U5762 (N_5762,N_3111,N_3268);
and U5763 (N_5763,N_3276,N_4050);
or U5764 (N_5764,N_3411,N_4390);
or U5765 (N_5765,N_3177,N_3495);
nor U5766 (N_5766,N_3232,N_3759);
or U5767 (N_5767,N_4311,N_4371);
or U5768 (N_5768,N_4108,N_4066);
nor U5769 (N_5769,N_3036,N_3539);
nand U5770 (N_5770,N_4265,N_3518);
or U5771 (N_5771,N_3409,N_3371);
nor U5772 (N_5772,N_3160,N_4174);
or U5773 (N_5773,N_3018,N_3100);
xor U5774 (N_5774,N_3000,N_3107);
and U5775 (N_5775,N_3307,N_3166);
or U5776 (N_5776,N_3510,N_3855);
and U5777 (N_5777,N_3123,N_3689);
and U5778 (N_5778,N_4051,N_3255);
nor U5779 (N_5779,N_4183,N_4435);
or U5780 (N_5780,N_3310,N_4460);
nand U5781 (N_5781,N_4350,N_3384);
nor U5782 (N_5782,N_3625,N_4043);
nor U5783 (N_5783,N_3417,N_3878);
nand U5784 (N_5784,N_4127,N_3343);
nand U5785 (N_5785,N_3968,N_4122);
and U5786 (N_5786,N_3010,N_3431);
and U5787 (N_5787,N_4455,N_4210);
and U5788 (N_5788,N_4265,N_3883);
nor U5789 (N_5789,N_3502,N_3894);
and U5790 (N_5790,N_4393,N_4302);
nand U5791 (N_5791,N_4439,N_4250);
nor U5792 (N_5792,N_4387,N_3568);
or U5793 (N_5793,N_3277,N_4184);
and U5794 (N_5794,N_3335,N_3448);
nand U5795 (N_5795,N_3684,N_3059);
nor U5796 (N_5796,N_3535,N_3815);
nor U5797 (N_5797,N_3147,N_3133);
nor U5798 (N_5798,N_3625,N_3530);
nor U5799 (N_5799,N_3664,N_3755);
and U5800 (N_5800,N_4048,N_4337);
or U5801 (N_5801,N_3449,N_3858);
xor U5802 (N_5802,N_3695,N_3651);
nor U5803 (N_5803,N_3890,N_3158);
or U5804 (N_5804,N_4261,N_3819);
nand U5805 (N_5805,N_3977,N_3131);
and U5806 (N_5806,N_3921,N_4385);
nand U5807 (N_5807,N_3416,N_3733);
or U5808 (N_5808,N_3686,N_4280);
or U5809 (N_5809,N_3053,N_4072);
or U5810 (N_5810,N_3334,N_4341);
or U5811 (N_5811,N_4001,N_3894);
and U5812 (N_5812,N_4452,N_3598);
nand U5813 (N_5813,N_4277,N_3930);
nor U5814 (N_5814,N_3029,N_4489);
nand U5815 (N_5815,N_4151,N_3620);
nor U5816 (N_5816,N_4228,N_3031);
or U5817 (N_5817,N_4273,N_4184);
or U5818 (N_5818,N_4084,N_3255);
nor U5819 (N_5819,N_3896,N_3448);
or U5820 (N_5820,N_3230,N_3884);
and U5821 (N_5821,N_3193,N_3743);
xnor U5822 (N_5822,N_3092,N_3700);
nor U5823 (N_5823,N_3558,N_4097);
or U5824 (N_5824,N_3422,N_3775);
and U5825 (N_5825,N_3752,N_3604);
or U5826 (N_5826,N_3130,N_4402);
or U5827 (N_5827,N_3041,N_4290);
nor U5828 (N_5828,N_3941,N_3467);
xor U5829 (N_5829,N_3561,N_3569);
or U5830 (N_5830,N_3093,N_3510);
nand U5831 (N_5831,N_3524,N_3594);
or U5832 (N_5832,N_4447,N_3377);
nor U5833 (N_5833,N_3708,N_3615);
nor U5834 (N_5834,N_3386,N_3251);
xor U5835 (N_5835,N_3339,N_4206);
and U5836 (N_5836,N_4087,N_4458);
or U5837 (N_5837,N_4174,N_3580);
nand U5838 (N_5838,N_4187,N_4124);
nor U5839 (N_5839,N_3654,N_3719);
and U5840 (N_5840,N_3474,N_3566);
nor U5841 (N_5841,N_3146,N_3427);
and U5842 (N_5842,N_3516,N_4222);
and U5843 (N_5843,N_3268,N_3005);
or U5844 (N_5844,N_3335,N_4424);
nor U5845 (N_5845,N_4393,N_3581);
xor U5846 (N_5846,N_3291,N_3140);
or U5847 (N_5847,N_3670,N_3091);
or U5848 (N_5848,N_4357,N_3896);
nor U5849 (N_5849,N_3608,N_4242);
or U5850 (N_5850,N_3969,N_3307);
and U5851 (N_5851,N_3801,N_4328);
or U5852 (N_5852,N_3364,N_3271);
and U5853 (N_5853,N_3543,N_3014);
nor U5854 (N_5854,N_3915,N_4423);
and U5855 (N_5855,N_4494,N_3304);
nand U5856 (N_5856,N_3290,N_3662);
and U5857 (N_5857,N_3083,N_3595);
nor U5858 (N_5858,N_3979,N_3632);
nor U5859 (N_5859,N_4176,N_4284);
nor U5860 (N_5860,N_3040,N_3611);
or U5861 (N_5861,N_4140,N_4111);
nor U5862 (N_5862,N_4387,N_4248);
and U5863 (N_5863,N_3249,N_3554);
xnor U5864 (N_5864,N_3763,N_3129);
nor U5865 (N_5865,N_4089,N_4174);
nand U5866 (N_5866,N_4415,N_4236);
nor U5867 (N_5867,N_4116,N_3122);
nand U5868 (N_5868,N_3785,N_3159);
and U5869 (N_5869,N_4448,N_3792);
nand U5870 (N_5870,N_3797,N_3785);
nor U5871 (N_5871,N_3212,N_3359);
and U5872 (N_5872,N_3106,N_4350);
xnor U5873 (N_5873,N_3009,N_3931);
nand U5874 (N_5874,N_3570,N_3900);
or U5875 (N_5875,N_3203,N_3608);
nand U5876 (N_5876,N_4390,N_3647);
or U5877 (N_5877,N_3700,N_4378);
xnor U5878 (N_5878,N_4438,N_3003);
nor U5879 (N_5879,N_4179,N_3174);
xnor U5880 (N_5880,N_3166,N_3359);
nor U5881 (N_5881,N_3584,N_3007);
or U5882 (N_5882,N_3526,N_4347);
nor U5883 (N_5883,N_3254,N_4317);
or U5884 (N_5884,N_3560,N_3999);
xnor U5885 (N_5885,N_3450,N_4396);
nor U5886 (N_5886,N_4371,N_3118);
or U5887 (N_5887,N_4039,N_3807);
nand U5888 (N_5888,N_3792,N_3211);
nand U5889 (N_5889,N_3780,N_4354);
xor U5890 (N_5890,N_3754,N_3558);
or U5891 (N_5891,N_3955,N_3096);
or U5892 (N_5892,N_4005,N_3554);
nor U5893 (N_5893,N_3897,N_3034);
and U5894 (N_5894,N_3421,N_3606);
xor U5895 (N_5895,N_3167,N_3289);
nand U5896 (N_5896,N_3116,N_3355);
and U5897 (N_5897,N_3239,N_3735);
nand U5898 (N_5898,N_3439,N_4452);
nor U5899 (N_5899,N_3212,N_4318);
nor U5900 (N_5900,N_3415,N_3798);
or U5901 (N_5901,N_3549,N_3913);
or U5902 (N_5902,N_4415,N_3877);
nor U5903 (N_5903,N_3749,N_3291);
nor U5904 (N_5904,N_3350,N_3294);
or U5905 (N_5905,N_4391,N_3742);
nand U5906 (N_5906,N_3622,N_3546);
nand U5907 (N_5907,N_3460,N_3528);
xor U5908 (N_5908,N_3159,N_4223);
xor U5909 (N_5909,N_3880,N_3329);
nor U5910 (N_5910,N_4152,N_4258);
nor U5911 (N_5911,N_3479,N_3232);
xor U5912 (N_5912,N_3955,N_3976);
nand U5913 (N_5913,N_3080,N_3396);
and U5914 (N_5914,N_4430,N_3818);
or U5915 (N_5915,N_3444,N_4459);
nand U5916 (N_5916,N_4232,N_4410);
nor U5917 (N_5917,N_3392,N_4220);
nor U5918 (N_5918,N_3222,N_3915);
and U5919 (N_5919,N_3052,N_3676);
and U5920 (N_5920,N_3777,N_3221);
xnor U5921 (N_5921,N_3641,N_3200);
or U5922 (N_5922,N_3104,N_4442);
or U5923 (N_5923,N_4485,N_3219);
nand U5924 (N_5924,N_4387,N_3241);
nand U5925 (N_5925,N_3092,N_3635);
or U5926 (N_5926,N_3268,N_3369);
and U5927 (N_5927,N_3729,N_3411);
or U5928 (N_5928,N_4454,N_4160);
or U5929 (N_5929,N_3772,N_4116);
xnor U5930 (N_5930,N_4336,N_3960);
or U5931 (N_5931,N_4263,N_4390);
nor U5932 (N_5932,N_3907,N_3929);
nand U5933 (N_5933,N_4163,N_4313);
and U5934 (N_5934,N_3979,N_3150);
nand U5935 (N_5935,N_3280,N_4038);
or U5936 (N_5936,N_4461,N_3052);
and U5937 (N_5937,N_3475,N_3466);
nand U5938 (N_5938,N_4013,N_3493);
xnor U5939 (N_5939,N_3150,N_3685);
nand U5940 (N_5940,N_4302,N_3975);
nor U5941 (N_5941,N_3688,N_3393);
nand U5942 (N_5942,N_4326,N_3327);
or U5943 (N_5943,N_3366,N_3625);
and U5944 (N_5944,N_3281,N_3036);
nand U5945 (N_5945,N_4301,N_4205);
nand U5946 (N_5946,N_3909,N_3895);
nor U5947 (N_5947,N_3564,N_3295);
nand U5948 (N_5948,N_3533,N_3061);
or U5949 (N_5949,N_4460,N_3358);
nand U5950 (N_5950,N_3157,N_3686);
and U5951 (N_5951,N_3190,N_3653);
or U5952 (N_5952,N_3705,N_3467);
and U5953 (N_5953,N_4101,N_3018);
or U5954 (N_5954,N_3254,N_4422);
nor U5955 (N_5955,N_3384,N_3968);
or U5956 (N_5956,N_3311,N_3328);
nor U5957 (N_5957,N_4018,N_3661);
nand U5958 (N_5958,N_3904,N_3740);
nand U5959 (N_5959,N_4261,N_3839);
or U5960 (N_5960,N_3835,N_3399);
or U5961 (N_5961,N_3704,N_3157);
and U5962 (N_5962,N_3599,N_3511);
or U5963 (N_5963,N_4373,N_3421);
nand U5964 (N_5964,N_4482,N_3706);
nand U5965 (N_5965,N_3313,N_3708);
and U5966 (N_5966,N_3487,N_3917);
nand U5967 (N_5967,N_4273,N_3380);
xor U5968 (N_5968,N_3778,N_3511);
nor U5969 (N_5969,N_4131,N_3338);
or U5970 (N_5970,N_3635,N_3965);
nand U5971 (N_5971,N_3384,N_4125);
xor U5972 (N_5972,N_3725,N_3766);
nand U5973 (N_5973,N_4194,N_3248);
and U5974 (N_5974,N_3603,N_3040);
and U5975 (N_5975,N_3711,N_3429);
or U5976 (N_5976,N_3820,N_3292);
or U5977 (N_5977,N_3841,N_3154);
nor U5978 (N_5978,N_4489,N_4268);
and U5979 (N_5979,N_3720,N_4276);
nor U5980 (N_5980,N_3085,N_3216);
nor U5981 (N_5981,N_3812,N_4472);
nor U5982 (N_5982,N_3243,N_4472);
nor U5983 (N_5983,N_4173,N_3080);
or U5984 (N_5984,N_4085,N_4488);
nor U5985 (N_5985,N_4451,N_4236);
and U5986 (N_5986,N_4334,N_3726);
or U5987 (N_5987,N_3099,N_4440);
or U5988 (N_5988,N_3325,N_3265);
xor U5989 (N_5989,N_3796,N_3518);
and U5990 (N_5990,N_4106,N_3127);
xor U5991 (N_5991,N_3487,N_4348);
or U5992 (N_5992,N_3686,N_3713);
nor U5993 (N_5993,N_4425,N_4046);
xor U5994 (N_5994,N_3057,N_4081);
nor U5995 (N_5995,N_4366,N_3994);
nand U5996 (N_5996,N_3250,N_3587);
or U5997 (N_5997,N_3661,N_3201);
nand U5998 (N_5998,N_3216,N_4478);
nand U5999 (N_5999,N_3221,N_3848);
or U6000 (N_6000,N_5125,N_5031);
nor U6001 (N_6001,N_5821,N_4723);
and U6002 (N_6002,N_4533,N_5006);
or U6003 (N_6003,N_5834,N_5176);
and U6004 (N_6004,N_5977,N_4852);
nor U6005 (N_6005,N_5955,N_5791);
and U6006 (N_6006,N_4857,N_5849);
nand U6007 (N_6007,N_5291,N_4811);
and U6008 (N_6008,N_5343,N_5133);
nor U6009 (N_6009,N_5585,N_4786);
nor U6010 (N_6010,N_4543,N_5987);
nor U6011 (N_6011,N_5757,N_5164);
or U6012 (N_6012,N_4604,N_4758);
nor U6013 (N_6013,N_5450,N_5101);
and U6014 (N_6014,N_5709,N_5926);
or U6015 (N_6015,N_5707,N_4664);
or U6016 (N_6016,N_5716,N_5517);
or U6017 (N_6017,N_5367,N_5512);
and U6018 (N_6018,N_4737,N_5676);
or U6019 (N_6019,N_5805,N_4710);
nand U6020 (N_6020,N_5300,N_5379);
nor U6021 (N_6021,N_5800,N_4762);
nor U6022 (N_6022,N_4589,N_4866);
or U6023 (N_6023,N_5168,N_5768);
and U6024 (N_6024,N_5384,N_5219);
xor U6025 (N_6025,N_4521,N_5163);
and U6026 (N_6026,N_5469,N_5761);
xor U6027 (N_6027,N_4803,N_4807);
or U6028 (N_6028,N_5232,N_5082);
nand U6029 (N_6029,N_5623,N_5932);
or U6030 (N_6030,N_4727,N_4862);
or U6031 (N_6031,N_4738,N_4554);
and U6032 (N_6032,N_5792,N_5545);
nand U6033 (N_6033,N_5643,N_5826);
or U6034 (N_6034,N_5378,N_5479);
nor U6035 (N_6035,N_4783,N_4679);
and U6036 (N_6036,N_4797,N_5533);
nand U6037 (N_6037,N_5774,N_5855);
xor U6038 (N_6038,N_5865,N_5796);
nand U6039 (N_6039,N_4986,N_4606);
nand U6040 (N_6040,N_4769,N_4962);
nand U6041 (N_6041,N_4711,N_4677);
xnor U6042 (N_6042,N_5007,N_5747);
nand U6043 (N_6043,N_4901,N_5965);
nor U6044 (N_6044,N_4657,N_5197);
or U6045 (N_6045,N_5756,N_4501);
and U6046 (N_6046,N_5595,N_5373);
xor U6047 (N_6047,N_4959,N_5655);
or U6048 (N_6048,N_5781,N_5825);
nand U6049 (N_6049,N_4970,N_4886);
nor U6050 (N_6050,N_5644,N_5346);
or U6051 (N_6051,N_4730,N_4602);
and U6052 (N_6052,N_5744,N_5257);
nand U6053 (N_6053,N_5582,N_5029);
nor U6054 (N_6054,N_4514,N_5460);
or U6055 (N_6055,N_5600,N_5397);
or U6056 (N_6056,N_5976,N_5216);
and U6057 (N_6057,N_5355,N_5348);
nor U6058 (N_6058,N_5626,N_5881);
or U6059 (N_6059,N_5454,N_5620);
xor U6060 (N_6060,N_4778,N_5952);
or U6061 (N_6061,N_5649,N_5632);
or U6062 (N_6062,N_5990,N_5698);
nand U6063 (N_6063,N_5048,N_5445);
xor U6064 (N_6064,N_4618,N_5551);
xnor U6065 (N_6065,N_4693,N_4828);
and U6066 (N_6066,N_5265,N_4814);
or U6067 (N_6067,N_5284,N_5306);
or U6068 (N_6068,N_4903,N_5844);
nor U6069 (N_6069,N_4817,N_4922);
nand U6070 (N_6070,N_5614,N_4990);
or U6071 (N_6071,N_5092,N_5763);
nand U6072 (N_6072,N_5640,N_5391);
and U6073 (N_6073,N_5058,N_5657);
nand U6074 (N_6074,N_5771,N_4920);
and U6075 (N_6075,N_4892,N_5966);
nand U6076 (N_6076,N_5960,N_5462);
and U6077 (N_6077,N_5225,N_5916);
and U6078 (N_6078,N_5631,N_4776);
nor U6079 (N_6079,N_4566,N_4721);
or U6080 (N_6080,N_4526,N_5453);
and U6081 (N_6081,N_5094,N_4592);
nor U6082 (N_6082,N_4728,N_5498);
and U6083 (N_6083,N_5458,N_5220);
or U6084 (N_6084,N_5764,N_5417);
and U6085 (N_6085,N_4957,N_5302);
nand U6086 (N_6086,N_5700,N_5557);
or U6087 (N_6087,N_5573,N_5637);
or U6088 (N_6088,N_4902,N_5576);
nand U6089 (N_6089,N_4847,N_4988);
nor U6090 (N_6090,N_5345,N_4751);
nand U6091 (N_6091,N_5194,N_5287);
or U6092 (N_6092,N_4539,N_4971);
xor U6093 (N_6093,N_5224,N_5424);
or U6094 (N_6094,N_4631,N_5119);
nand U6095 (N_6095,N_4871,N_5726);
and U6096 (N_6096,N_4932,N_5583);
and U6097 (N_6097,N_4593,N_5671);
nor U6098 (N_6098,N_5079,N_5661);
nor U6099 (N_6099,N_4582,N_4967);
and U6100 (N_6100,N_5681,N_5853);
nor U6101 (N_6101,N_5123,N_5118);
nor U6102 (N_6102,N_5374,N_4870);
nor U6103 (N_6103,N_5175,N_4872);
nand U6104 (N_6104,N_4934,N_4535);
or U6105 (N_6105,N_4795,N_4873);
nor U6106 (N_6106,N_5828,N_4598);
or U6107 (N_6107,N_5263,N_5850);
nor U6108 (N_6108,N_5239,N_5276);
nor U6109 (N_6109,N_4517,N_4599);
xnor U6110 (N_6110,N_5651,N_4757);
or U6111 (N_6111,N_4840,N_5930);
nor U6112 (N_6112,N_5913,N_4575);
nand U6113 (N_6113,N_4629,N_4729);
or U6114 (N_6114,N_4616,N_5230);
or U6115 (N_6115,N_5147,N_5096);
nor U6116 (N_6116,N_5452,N_5080);
xnor U6117 (N_6117,N_5028,N_5245);
xnor U6118 (N_6118,N_4780,N_4691);
nor U6119 (N_6119,N_4619,N_5843);
or U6120 (N_6120,N_5138,N_5605);
xor U6121 (N_6121,N_5408,N_5519);
nand U6122 (N_6122,N_5034,N_5650);
or U6123 (N_6123,N_5072,N_4890);
nor U6124 (N_6124,N_5363,N_5560);
or U6125 (N_6125,N_5003,N_4676);
nand U6126 (N_6126,N_5815,N_5196);
nor U6127 (N_6127,N_5621,N_5032);
nand U6128 (N_6128,N_5909,N_5900);
nand U6129 (N_6129,N_5552,N_5658);
or U6130 (N_6130,N_5663,N_5336);
nor U6131 (N_6131,N_5157,N_4844);
nor U6132 (N_6132,N_5019,N_5496);
or U6133 (N_6133,N_4742,N_4587);
and U6134 (N_6134,N_5038,N_4768);
nand U6135 (N_6135,N_4960,N_5301);
and U6136 (N_6136,N_5974,N_4835);
and U6137 (N_6137,N_5714,N_4996);
nor U6138 (N_6138,N_5799,N_5786);
nand U6139 (N_6139,N_5285,N_5759);
or U6140 (N_6140,N_4955,N_4538);
or U6141 (N_6141,N_5307,N_5337);
and U6142 (N_6142,N_4510,N_5782);
nand U6143 (N_6143,N_4607,N_5594);
or U6144 (N_6144,N_5622,N_4977);
and U6145 (N_6145,N_5540,N_4662);
nand U6146 (N_6146,N_5494,N_4699);
or U6147 (N_6147,N_5905,N_5213);
or U6148 (N_6148,N_5723,N_4731);
nor U6149 (N_6149,N_4788,N_5227);
nand U6150 (N_6150,N_4830,N_5735);
xnor U6151 (N_6151,N_4546,N_5470);
or U6152 (N_6152,N_5228,N_5710);
and U6153 (N_6153,N_5074,N_5968);
or U6154 (N_6154,N_5888,N_5143);
and U6155 (N_6155,N_4666,N_4658);
xor U6156 (N_6156,N_4919,N_4838);
or U6157 (N_6157,N_4573,N_5130);
nand U6158 (N_6158,N_5243,N_4725);
nor U6159 (N_6159,N_4652,N_5407);
nand U6160 (N_6160,N_5894,N_5013);
or U6161 (N_6161,N_4966,N_5639);
nand U6162 (N_6162,N_5642,N_5113);
and U6163 (N_6163,N_5515,N_5137);
or U6164 (N_6164,N_5429,N_5127);
nor U6165 (N_6165,N_5910,N_5192);
or U6166 (N_6166,N_5487,N_4692);
and U6167 (N_6167,N_4622,N_5488);
nor U6168 (N_6168,N_4669,N_4821);
xor U6169 (N_6169,N_4734,N_4802);
or U6170 (N_6170,N_5769,N_5332);
xnor U6171 (N_6171,N_4956,N_5142);
nand U6172 (N_6172,N_5288,N_5705);
xnor U6173 (N_6173,N_5702,N_4884);
nor U6174 (N_6174,N_5908,N_5914);
nand U6175 (N_6175,N_5040,N_5776);
or U6176 (N_6176,N_5953,N_4696);
and U6177 (N_6177,N_5069,N_5467);
or U6178 (N_6178,N_4686,N_5674);
xor U6179 (N_6179,N_5876,N_5489);
and U6180 (N_6180,N_5530,N_4531);
nand U6181 (N_6181,N_4946,N_4528);
nand U6182 (N_6182,N_5528,N_5158);
nor U6183 (N_6183,N_5253,N_4899);
or U6184 (N_6184,N_5720,N_5544);
nand U6185 (N_6185,N_5466,N_4644);
nor U6186 (N_6186,N_4542,N_5724);
and U6187 (N_6187,N_4614,N_5304);
xnor U6188 (N_6188,N_5693,N_5514);
nor U6189 (N_6189,N_4709,N_5588);
xor U6190 (N_6190,N_5559,N_5387);
or U6191 (N_6191,N_5793,N_4842);
nor U6192 (N_6192,N_4829,N_5247);
or U6193 (N_6193,N_5303,N_5993);
or U6194 (N_6194,N_5593,N_5633);
and U6195 (N_6195,N_5983,N_5523);
nor U6196 (N_6196,N_5235,N_5997);
nor U6197 (N_6197,N_4954,N_4815);
nand U6198 (N_6198,N_5982,N_5659);
nand U6199 (N_6199,N_5959,N_5190);
nand U6200 (N_6200,N_5110,N_4735);
nand U6201 (N_6201,N_4855,N_5410);
and U6202 (N_6202,N_5592,N_4520);
nor U6203 (N_6203,N_4944,N_5618);
or U6204 (N_6204,N_4541,N_5372);
nor U6205 (N_6205,N_5734,N_4585);
nand U6206 (N_6206,N_4524,N_4813);
and U6207 (N_6207,N_5803,N_5571);
nand U6208 (N_6208,N_5836,N_4794);
and U6209 (N_6209,N_5317,N_5087);
nor U6210 (N_6210,N_4525,N_5210);
nand U6211 (N_6211,N_4576,N_5845);
nor U6212 (N_6212,N_5956,N_5969);
nand U6213 (N_6213,N_4981,N_5824);
xor U6214 (N_6214,N_5308,N_5282);
and U6215 (N_6215,N_5043,N_5296);
nand U6216 (N_6216,N_4595,N_4621);
nand U6217 (N_6217,N_4741,N_5338);
nor U6218 (N_6218,N_5711,N_4653);
nor U6219 (N_6219,N_5677,N_5719);
and U6220 (N_6220,N_5160,N_4808);
and U6221 (N_6221,N_5508,N_4748);
nand U6222 (N_6222,N_5923,N_5963);
and U6223 (N_6223,N_4623,N_5144);
or U6224 (N_6224,N_5875,N_5922);
nor U6225 (N_6225,N_5558,N_5446);
xnor U6226 (N_6226,N_5992,N_5035);
nor U6227 (N_6227,N_5520,N_4574);
nor U6228 (N_6228,N_5026,N_5667);
nand U6229 (N_6229,N_5505,N_4639);
nand U6230 (N_6230,N_4714,N_5172);
nand U6231 (N_6231,N_5076,N_5122);
nand U6232 (N_6232,N_5510,N_4910);
nand U6233 (N_6233,N_5393,N_5773);
nor U6234 (N_6234,N_4879,N_4646);
nor U6235 (N_6235,N_5706,N_5687);
nor U6236 (N_6236,N_5527,N_5195);
nor U6237 (N_6237,N_4874,N_5179);
nand U6238 (N_6238,N_4889,N_5548);
and U6239 (N_6239,N_4854,N_5690);
nand U6240 (N_6240,N_5177,N_4583);
nor U6241 (N_6241,N_5991,N_5725);
nand U6242 (N_6242,N_4650,N_5067);
and U6243 (N_6243,N_5180,N_4605);
nor U6244 (N_6244,N_4518,N_4567);
nand U6245 (N_6245,N_4754,N_5619);
or U6246 (N_6246,N_4883,N_5145);
xnor U6247 (N_6247,N_5281,N_4880);
nand U6248 (N_6248,N_4519,N_4506);
and U6249 (N_6249,N_5750,N_4825);
nand U6250 (N_6250,N_5093,N_5349);
nand U6251 (N_6251,N_5126,N_4749);
xor U6252 (N_6252,N_5120,N_5624);
nand U6253 (N_6253,N_5617,N_5872);
and U6254 (N_6254,N_5684,N_4701);
nand U6255 (N_6255,N_4645,N_4790);
nor U6256 (N_6256,N_5537,N_5973);
and U6257 (N_6257,N_5381,N_5459);
or U6258 (N_6258,N_5717,N_5002);
or U6259 (N_6259,N_5733,N_4550);
nand U6260 (N_6260,N_4948,N_4836);
nand U6261 (N_6261,N_4881,N_4522);
and U6262 (N_6262,N_5008,N_5511);
nor U6263 (N_6263,N_5925,N_5091);
nand U6264 (N_6264,N_5327,N_5598);
nand U6265 (N_6265,N_5695,N_5423);
xnor U6266 (N_6266,N_5108,N_4824);
or U6267 (N_6267,N_5811,N_4951);
nand U6268 (N_6268,N_5440,N_5241);
and U6269 (N_6269,N_5314,N_4911);
and U6270 (N_6270,N_5935,N_4994);
and U6271 (N_6271,N_5940,N_4654);
xnor U6272 (N_6272,N_5903,N_5840);
nor U6273 (N_6273,N_5015,N_4924);
or U6274 (N_6274,N_4505,N_5516);
or U6275 (N_6275,N_5085,N_5638);
nor U6276 (N_6276,N_5679,N_5563);
nor U6277 (N_6277,N_5597,N_5708);
and U6278 (N_6278,N_5320,N_5586);
and U6279 (N_6279,N_4826,N_5689);
nor U6280 (N_6280,N_5155,N_4865);
or U6281 (N_6281,N_5541,N_5415);
nor U6282 (N_6282,N_5680,N_4635);
nand U6283 (N_6283,N_4529,N_4912);
nor U6284 (N_6284,N_4896,N_5267);
nand U6285 (N_6285,N_5493,N_5729);
and U6286 (N_6286,N_5084,N_5703);
nor U6287 (N_6287,N_4895,N_5242);
nand U6288 (N_6288,N_4800,N_5478);
nand U6289 (N_6289,N_5746,N_5859);
or U6290 (N_6290,N_4995,N_5376);
nor U6291 (N_6291,N_5670,N_5736);
nand U6292 (N_6292,N_4894,N_4552);
nor U6293 (N_6293,N_5941,N_5406);
nand U6294 (N_6294,N_5481,N_5613);
nor U6295 (N_6295,N_4939,N_5666);
nor U6296 (N_6296,N_5042,N_5686);
nor U6297 (N_6297,N_5664,N_5602);
and U6298 (N_6298,N_5864,N_4916);
xor U6299 (N_6299,N_5901,N_4570);
nand U6300 (N_6300,N_5293,N_5536);
or U6301 (N_6301,N_5139,N_5911);
and U6302 (N_6302,N_5752,N_4781);
nand U6303 (N_6303,N_5140,N_5476);
nand U6304 (N_6304,N_5004,N_5297);
nand U6305 (N_6305,N_4663,N_5753);
nor U6306 (N_6306,N_4562,N_5873);
or U6307 (N_6307,N_5463,N_5924);
nand U6308 (N_6308,N_4683,N_5731);
or U6309 (N_6309,N_4509,N_5529);
xor U6310 (N_6310,N_4885,N_5315);
nand U6311 (N_6311,N_5730,N_4551);
xnor U6312 (N_6312,N_5755,N_5813);
and U6313 (N_6313,N_4673,N_5165);
xnor U6314 (N_6314,N_5421,N_5513);
xnor U6315 (N_6315,N_4684,N_4945);
nor U6316 (N_6316,N_5857,N_5052);
or U6317 (N_6317,N_4628,N_4511);
nor U6318 (N_6318,N_5669,N_5701);
and U6319 (N_6319,N_5893,N_5036);
and U6320 (N_6320,N_5590,N_5835);
and U6321 (N_6321,N_5906,N_4841);
nor U6322 (N_6322,N_5403,N_5389);
nand U6323 (N_6323,N_4905,N_4779);
nor U6324 (N_6324,N_4561,N_5538);
nand U6325 (N_6325,N_5251,N_5057);
or U6326 (N_6326,N_4591,N_5295);
nand U6327 (N_6327,N_4702,N_5416);
nand U6328 (N_6328,N_4578,N_5570);
and U6329 (N_6329,N_5159,N_5063);
nor U6330 (N_6330,N_5823,N_5971);
or U6331 (N_6331,N_5102,N_5098);
nand U6332 (N_6332,N_4968,N_5390);
xor U6333 (N_6333,N_5205,N_5129);
and U6334 (N_6334,N_4915,N_5174);
nand U6335 (N_6335,N_4752,N_5949);
or U6336 (N_6336,N_5967,N_4633);
nand U6337 (N_6337,N_4613,N_5395);
nand U6338 (N_6338,N_5331,N_5271);
or U6339 (N_6339,N_5161,N_5854);
and U6340 (N_6340,N_4600,N_5890);
nor U6341 (N_6341,N_4888,N_5798);
nand U6342 (N_6342,N_5289,N_4914);
xnor U6343 (N_6343,N_5432,N_5556);
and U6344 (N_6344,N_5685,N_4819);
or U6345 (N_6345,N_5555,N_4827);
or U6346 (N_6346,N_5419,N_5979);
or U6347 (N_6347,N_5269,N_5049);
or U6348 (N_6348,N_4625,N_4630);
xnor U6349 (N_6349,N_4667,N_5095);
nor U6350 (N_6350,N_5173,N_5044);
nor U6351 (N_6351,N_5927,N_5249);
nand U6352 (N_6352,N_4579,N_5319);
or U6353 (N_6353,N_5068,N_4816);
nor U6354 (N_6354,N_4685,N_4512);
or U6355 (N_6355,N_5532,N_5920);
xor U6356 (N_6356,N_5964,N_5141);
or U6357 (N_6357,N_5848,N_5630);
nor U6358 (N_6358,N_5937,N_4700);
xnor U6359 (N_6359,N_4581,N_5465);
and U6360 (N_6360,N_4975,N_4926);
nor U6361 (N_6361,N_4743,N_5608);
or U6362 (N_6362,N_5616,N_5645);
nand U6363 (N_6363,N_5231,N_5311);
and U6364 (N_6364,N_5156,N_5081);
nand U6365 (N_6365,N_5264,N_4853);
and U6366 (N_6366,N_5201,N_5656);
nor U6367 (N_6367,N_5200,N_5441);
and U6368 (N_6368,N_5439,N_5229);
nand U6369 (N_6369,N_5070,N_5340);
and U6370 (N_6370,N_4627,N_5193);
or U6371 (N_6371,N_5842,N_4636);
nor U6372 (N_6372,N_5212,N_5790);
and U6373 (N_6373,N_5699,N_4864);
and U6374 (N_6374,N_5862,N_5604);
and U6375 (N_6375,N_5411,N_5103);
nor U6376 (N_6376,N_5256,N_4770);
xnor U6377 (N_6377,N_5322,N_4739);
nand U6378 (N_6378,N_5889,N_5895);
nand U6379 (N_6379,N_4672,N_5827);
nor U6380 (N_6380,N_5426,N_4637);
nor U6381 (N_6381,N_4972,N_5567);
nand U6382 (N_6382,N_5207,N_5075);
and U6383 (N_6383,N_5509,N_5341);
nor U6384 (N_6384,N_4984,N_5817);
nor U6385 (N_6385,N_5100,N_5861);
nor U6386 (N_6386,N_5178,N_5083);
nand U6387 (N_6387,N_4898,N_4882);
nand U6388 (N_6388,N_5504,N_4850);
or U6389 (N_6389,N_5783,N_4610);
nor U6390 (N_6390,N_5921,N_5754);
and U6391 (N_6391,N_4736,N_4943);
nor U6392 (N_6392,N_5045,N_5596);
nor U6393 (N_6393,N_4810,N_4564);
nand U6394 (N_6394,N_5434,N_4978);
and U6395 (N_6395,N_5182,N_5501);
xor U6396 (N_6396,N_5366,N_4942);
and U6397 (N_6397,N_5554,N_4998);
and U6398 (N_6398,N_5473,N_4860);
and U6399 (N_6399,N_5739,N_4747);
nand U6400 (N_6400,N_4722,N_5951);
or U6401 (N_6401,N_5612,N_4745);
nor U6402 (N_6402,N_5652,N_4868);
nor U6403 (N_6403,N_4964,N_4785);
nand U6404 (N_6404,N_5892,N_5778);
nand U6405 (N_6405,N_5436,N_5396);
or U6406 (N_6406,N_5060,N_5751);
and U6407 (N_6407,N_5564,N_5683);
nand U6408 (N_6408,N_5447,N_5316);
xor U6409 (N_6409,N_5443,N_5722);
and U6410 (N_6410,N_4609,N_5209);
or U6411 (N_6411,N_4818,N_4689);
nor U6412 (N_6412,N_4513,N_5115);
or U6413 (N_6413,N_5606,N_5323);
or U6414 (N_6414,N_5361,N_5246);
and U6415 (N_6415,N_5697,N_5185);
nand U6416 (N_6416,N_4806,N_5326);
or U6417 (N_6417,N_4532,N_4717);
nor U6418 (N_6418,N_4558,N_4671);
nor U6419 (N_6419,N_4965,N_5055);
xnor U6420 (N_6420,N_5627,N_4863);
and U6421 (N_6421,N_5053,N_5948);
nand U6422 (N_6422,N_5442,N_5915);
nand U6423 (N_6423,N_5342,N_4682);
and U6424 (N_6424,N_5525,N_5758);
or U6425 (N_6425,N_5305,N_5187);
nand U6426 (N_6426,N_5017,N_5678);
nor U6427 (N_6427,N_5918,N_5005);
or U6428 (N_6428,N_5898,N_4985);
nor U6429 (N_6429,N_5106,N_4974);
nand U6430 (N_6430,N_5810,N_5765);
nor U6431 (N_6431,N_5542,N_5996);
nand U6432 (N_6432,N_5694,N_4504);
nand U6433 (N_6433,N_5430,N_4507);
or U6434 (N_6434,N_5899,N_4680);
xor U6435 (N_6435,N_4715,N_4647);
nor U6436 (N_6436,N_5354,N_4839);
or U6437 (N_6437,N_5985,N_5858);
nor U6438 (N_6438,N_4831,N_5767);
and U6439 (N_6439,N_5775,N_5660);
and U6440 (N_6440,N_4568,N_5449);
and U6441 (N_6441,N_5866,N_5062);
nand U6442 (N_6442,N_5428,N_5904);
or U6443 (N_6443,N_5211,N_5673);
xor U6444 (N_6444,N_5418,N_5938);
or U6445 (N_6445,N_4856,N_5398);
and U6446 (N_6446,N_5524,N_4503);
or U6447 (N_6447,N_5981,N_4958);
and U6448 (N_6448,N_4897,N_4557);
and U6449 (N_6449,N_5989,N_4620);
and U6450 (N_6450,N_5360,N_4547);
or U6451 (N_6451,N_5388,N_5420);
nand U6452 (N_6452,N_5727,N_4668);
nor U6453 (N_6453,N_5433,N_5869);
nor U6454 (N_6454,N_5309,N_5027);
xnor U6455 (N_6455,N_4812,N_5198);
and U6456 (N_6456,N_4764,N_5492);
and U6457 (N_6457,N_5777,N_4858);
and U6458 (N_6458,N_5766,N_4549);
nand U6459 (N_6459,N_5486,N_5609);
nor U6460 (N_6460,N_5988,N_5191);
nor U6461 (N_6461,N_5237,N_4876);
nor U6462 (N_6462,N_5500,N_5785);
xnor U6463 (N_6463,N_5547,N_5012);
and U6464 (N_6464,N_5833,N_5896);
nor U6465 (N_6465,N_4718,N_5599);
nand U6466 (N_6466,N_4976,N_5648);
xor U6467 (N_6467,N_5578,N_5518);
and U6468 (N_6468,N_5064,N_5891);
and U6469 (N_6469,N_4537,N_5167);
and U6470 (N_6470,N_5290,N_5362);
nor U6471 (N_6471,N_5841,N_4921);
and U6472 (N_6472,N_5860,N_5568);
or U6473 (N_6473,N_5409,N_5377);
or U6474 (N_6474,N_5574,N_5867);
xnor U6475 (N_6475,N_5275,N_4670);
or U6476 (N_6476,N_5186,N_5359);
nor U6477 (N_6477,N_5818,N_5880);
and U6478 (N_6478,N_4792,N_5902);
nor U6479 (N_6479,N_5077,N_5279);
nor U6480 (N_6480,N_5328,N_5150);
or U6481 (N_6481,N_4724,N_5802);
xor U6482 (N_6482,N_5111,N_4641);
and U6483 (N_6483,N_5628,N_5566);
nand U6484 (N_6484,N_5882,N_4705);
nor U6485 (N_6485,N_5995,N_5692);
nand U6486 (N_6486,N_4940,N_5183);
xor U6487 (N_6487,N_5954,N_4767);
or U6488 (N_6488,N_4516,N_5772);
xnor U6489 (N_6489,N_5184,N_5413);
or U6490 (N_6490,N_5472,N_5061);
and U6491 (N_6491,N_4548,N_4963);
or U6492 (N_6492,N_4877,N_5414);
nand U6493 (N_6493,N_5665,N_5745);
nor U6494 (N_6494,N_4798,N_5051);
and U6495 (N_6495,N_5738,N_5740);
and U6496 (N_6496,N_5961,N_5485);
nor U6497 (N_6497,N_5779,N_5116);
and U6498 (N_6498,N_5254,N_4848);
nor U6499 (N_6499,N_5749,N_4867);
nand U6500 (N_6500,N_5400,N_5356);
nor U6501 (N_6501,N_5318,N_5874);
nand U6502 (N_6502,N_5589,N_5009);
and U6503 (N_6503,N_5942,N_4875);
and U6504 (N_6504,N_4572,N_4571);
nor U6505 (N_6505,N_4703,N_4713);
nor U6506 (N_6506,N_5427,N_5457);
or U6507 (N_6507,N_5696,N_4846);
and U6508 (N_6508,N_5572,N_5250);
nand U6509 (N_6509,N_4791,N_4891);
nand U6510 (N_6510,N_5046,N_5121);
and U6511 (N_6511,N_4651,N_5054);
xnor U6512 (N_6512,N_5856,N_5104);
and U6513 (N_6513,N_4675,N_5298);
xnor U6514 (N_6514,N_5422,N_5975);
nand U6515 (N_6515,N_5591,N_5401);
nor U6516 (N_6516,N_5497,N_5073);
xor U6517 (N_6517,N_5561,N_5808);
xor U6518 (N_6518,N_5531,N_4787);
or U6519 (N_6519,N_5829,N_5059);
xnor U6520 (N_6520,N_5351,N_5662);
or U6521 (N_6521,N_5831,N_4584);
nor U6522 (N_6522,N_5405,N_5713);
or U6523 (N_6523,N_4733,N_5522);
nand U6524 (N_6524,N_4923,N_4695);
and U6525 (N_6525,N_5325,N_4845);
or U6526 (N_6526,N_5748,N_5151);
or U6527 (N_6527,N_5347,N_5283);
and U6528 (N_6528,N_5939,N_5482);
nor U6529 (N_6529,N_5986,N_5128);
xor U6530 (N_6530,N_5310,N_5732);
or U6531 (N_6531,N_5721,N_5202);
and U6532 (N_6532,N_5477,N_5294);
nand U6533 (N_6533,N_4530,N_4624);
nand U6534 (N_6534,N_5030,N_5728);
nor U6535 (N_6535,N_4586,N_4805);
and U6536 (N_6536,N_5820,N_5404);
and U6537 (N_6537,N_4904,N_5350);
xor U6538 (N_6538,N_5970,N_4569);
nor U6539 (N_6539,N_5399,N_5839);
and U6540 (N_6540,N_4983,N_5236);
and U6541 (N_6541,N_5980,N_5280);
nor U6542 (N_6542,N_5371,N_4941);
or U6543 (N_6543,N_5742,N_5780);
nand U6544 (N_6544,N_5553,N_5884);
and U6545 (N_6545,N_5610,N_4809);
nor U6546 (N_6546,N_5461,N_5448);
and U6547 (N_6547,N_5575,N_4707);
and U6548 (N_6548,N_5543,N_4665);
and U6549 (N_6549,N_4590,N_4823);
nand U6550 (N_6550,N_5016,N_5838);
or U6551 (N_6551,N_4992,N_5535);
nand U6552 (N_6552,N_5611,N_4704);
or U6553 (N_6553,N_4997,N_5221);
nand U6554 (N_6554,N_4887,N_5321);
nor U6555 (N_6555,N_5770,N_5382);
nand U6556 (N_6556,N_5000,N_5490);
xor U6557 (N_6557,N_5919,N_4936);
or U6558 (N_6558,N_5392,N_4720);
and U6559 (N_6559,N_5534,N_4801);
and U6560 (N_6560,N_5025,N_4608);
and U6561 (N_6561,N_5244,N_5760);
and U6562 (N_6562,N_4750,N_5261);
nor U6563 (N_6563,N_5089,N_5584);
nor U6564 (N_6564,N_5154,N_4643);
and U6565 (N_6565,N_4740,N_5830);
or U6566 (N_6566,N_5020,N_5124);
and U6567 (N_6567,N_4931,N_5483);
or U6568 (N_6568,N_5812,N_4746);
nor U6569 (N_6569,N_5109,N_4594);
nand U6570 (N_6570,N_5999,N_5832);
xnor U6571 (N_6571,N_5870,N_4893);
and U6572 (N_6572,N_5809,N_4928);
xor U6573 (N_6573,N_4822,N_5521);
and U6574 (N_6574,N_5464,N_5741);
or U6575 (N_6575,N_5947,N_5252);
nand U6576 (N_6576,N_4648,N_5474);
nand U6577 (N_6577,N_5958,N_5217);
or U6578 (N_6578,N_5099,N_4775);
nor U6579 (N_6579,N_4612,N_5878);
xor U6580 (N_6580,N_4674,N_5743);
and U6581 (N_6581,N_5438,N_5218);
or U6582 (N_6582,N_4793,N_5936);
nor U6583 (N_6583,N_4577,N_4597);
or U6584 (N_6584,N_5712,N_4580);
or U6585 (N_6585,N_4999,N_4744);
nor U6586 (N_6586,N_5789,N_4678);
nor U6587 (N_6587,N_4982,N_5934);
nand U6588 (N_6588,N_4952,N_4989);
or U6589 (N_6589,N_4777,N_5784);
xor U6590 (N_6590,N_5672,N_4935);
nand U6591 (N_6591,N_5037,N_5189);
or U6592 (N_6592,N_5928,N_5480);
or U6593 (N_6593,N_4565,N_4706);
nor U6594 (N_6594,N_5259,N_5268);
or U6595 (N_6595,N_4927,N_4716);
or U6596 (N_6596,N_5629,N_4774);
nand U6597 (N_6597,N_5206,N_5526);
nand U6598 (N_6598,N_5364,N_4799);
nor U6599 (N_6599,N_5358,N_4961);
xnor U6600 (N_6600,N_5071,N_5386);
nand U6601 (N_6601,N_4869,N_4784);
nand U6602 (N_6602,N_5819,N_5654);
xor U6603 (N_6603,N_5682,N_4929);
or U6604 (N_6604,N_4900,N_5797);
nand U6605 (N_6605,N_5357,N_5148);
and U6606 (N_6606,N_4837,N_5056);
or U6607 (N_6607,N_5912,N_5806);
or U6608 (N_6608,N_5851,N_5199);
nor U6609 (N_6609,N_5117,N_5962);
and U6610 (N_6610,N_5370,N_5335);
nand U6611 (N_6611,N_4834,N_5233);
nor U6612 (N_6612,N_4642,N_4611);
nand U6613 (N_6613,N_4694,N_4688);
nor U6614 (N_6614,N_5383,N_5863);
or U6615 (N_6615,N_4878,N_5668);
nand U6616 (N_6616,N_4502,N_5402);
or U6617 (N_6617,N_5299,N_4656);
or U6618 (N_6618,N_5078,N_5565);
xnor U6619 (N_6619,N_4545,N_5188);
nor U6620 (N_6620,N_4536,N_5380);
nor U6621 (N_6621,N_4820,N_5066);
nor U6622 (N_6622,N_5887,N_4913);
and U6623 (N_6623,N_5871,N_4947);
nand U6624 (N_6624,N_5506,N_4804);
or U6625 (N_6625,N_5944,N_4708);
and U6626 (N_6626,N_5580,N_4756);
or U6627 (N_6627,N_5647,N_5837);
nor U6628 (N_6628,N_5041,N_5023);
or U6629 (N_6629,N_5097,N_5957);
and U6630 (N_6630,N_4937,N_5437);
or U6631 (N_6631,N_5272,N_5412);
nand U6632 (N_6632,N_4861,N_4681);
and U6633 (N_6633,N_4953,N_5984);
or U6634 (N_6634,N_5385,N_4773);
and U6635 (N_6635,N_5022,N_5877);
nor U6636 (N_6636,N_5170,N_4726);
or U6637 (N_6637,N_4993,N_5804);
or U6638 (N_6638,N_5737,N_5581);
or U6639 (N_6639,N_4979,N_5943);
or U6640 (N_6640,N_5603,N_5885);
nor U6641 (N_6641,N_5152,N_5491);
nand U6642 (N_6642,N_5762,N_5258);
nor U6643 (N_6643,N_5273,N_5577);
or U6644 (N_6644,N_4555,N_4559);
or U6645 (N_6645,N_5105,N_5248);
xnor U6646 (N_6646,N_4649,N_5607);
xor U6647 (N_6647,N_5562,N_5431);
nand U6648 (N_6648,N_5897,N_4640);
nand U6649 (N_6649,N_4789,N_5131);
xnor U6650 (N_6650,N_4907,N_5277);
or U6651 (N_6651,N_5675,N_5635);
and U6652 (N_6652,N_4534,N_4712);
or U6653 (N_6653,N_4933,N_5134);
nand U6654 (N_6654,N_5471,N_5146);
nand U6655 (N_6655,N_4849,N_5226);
and U6656 (N_6656,N_5033,N_5333);
nor U6657 (N_6657,N_5507,N_4563);
or U6658 (N_6658,N_5615,N_5208);
xnor U6659 (N_6659,N_5931,N_5569);
nand U6660 (N_6660,N_5153,N_5579);
nand U6661 (N_6661,N_4753,N_5215);
and U6662 (N_6662,N_4601,N_5181);
nand U6663 (N_6663,N_5456,N_5455);
or U6664 (N_6664,N_5330,N_5451);
xor U6665 (N_6665,N_4560,N_4527);
nor U6666 (N_6666,N_5166,N_5312);
nor U6667 (N_6667,N_5171,N_5204);
or U6668 (N_6668,N_4617,N_5203);
or U6669 (N_6669,N_4969,N_5024);
xnor U6670 (N_6670,N_4908,N_5047);
xor U6671 (N_6671,N_5634,N_5950);
nand U6672 (N_6672,N_4540,N_5353);
nor U6673 (N_6673,N_5846,N_5018);
nand U6674 (N_6674,N_4763,N_4626);
nand U6675 (N_6675,N_5468,N_5136);
nand U6676 (N_6676,N_5425,N_5050);
nand U6677 (N_6677,N_4833,N_5549);
xor U6678 (N_6678,N_4832,N_5014);
nand U6679 (N_6679,N_4515,N_4765);
and U6680 (N_6680,N_5994,N_5852);
and U6681 (N_6681,N_5369,N_4796);
and U6682 (N_6682,N_5972,N_4615);
nand U6683 (N_6683,N_5794,N_5868);
or U6684 (N_6684,N_4698,N_5503);
or U6685 (N_6685,N_4661,N_5946);
and U6686 (N_6686,N_5313,N_5907);
and U6687 (N_6687,N_5601,N_4909);
or U6688 (N_6688,N_5787,N_5814);
or U6689 (N_6689,N_5394,N_4938);
nand U6690 (N_6690,N_5169,N_5238);
and U6691 (N_6691,N_5625,N_4851);
nand U6692 (N_6692,N_4950,N_5822);
and U6693 (N_6693,N_4697,N_5886);
xor U6694 (N_6694,N_5001,N_5214);
nor U6695 (N_6695,N_4523,N_4843);
nand U6696 (N_6696,N_4782,N_4659);
or U6697 (N_6697,N_4859,N_4949);
and U6698 (N_6698,N_5266,N_4634);
or U6699 (N_6699,N_5010,N_5222);
and U6700 (N_6700,N_4553,N_5324);
nor U6701 (N_6701,N_4772,N_5255);
or U6702 (N_6702,N_5495,N_5816);
and U6703 (N_6703,N_5539,N_5039);
nor U6704 (N_6704,N_5270,N_4918);
nor U6705 (N_6705,N_5162,N_4973);
nand U6706 (N_6706,N_4755,N_5114);
or U6707 (N_6707,N_5929,N_4687);
nand U6708 (N_6708,N_5484,N_5240);
and U6709 (N_6709,N_4771,N_5883);
nor U6710 (N_6710,N_5978,N_4632);
and U6711 (N_6711,N_5274,N_4556);
nor U6712 (N_6712,N_5278,N_5223);
or U6713 (N_6713,N_5688,N_5788);
nor U6714 (N_6714,N_5262,N_5344);
or U6715 (N_6715,N_5847,N_5149);
or U6716 (N_6716,N_4761,N_4588);
or U6717 (N_6717,N_5368,N_5021);
nor U6718 (N_6718,N_5636,N_5691);
xnor U6719 (N_6719,N_5107,N_4766);
nor U6720 (N_6720,N_5945,N_5998);
nand U6721 (N_6721,N_4638,N_5365);
nor U6722 (N_6722,N_4760,N_5088);
nor U6723 (N_6723,N_5653,N_4732);
and U6724 (N_6724,N_5329,N_5011);
and U6725 (N_6725,N_5718,N_5260);
and U6726 (N_6726,N_5132,N_4660);
or U6727 (N_6727,N_5704,N_5546);
or U6728 (N_6728,N_5086,N_4603);
nand U6729 (N_6729,N_4759,N_4925);
nand U6730 (N_6730,N_4508,N_4906);
nor U6731 (N_6731,N_4980,N_5065);
nor U6732 (N_6732,N_5550,N_5917);
or U6733 (N_6733,N_5334,N_5587);
nor U6734 (N_6734,N_5646,N_4690);
or U6735 (N_6735,N_5090,N_4991);
nor U6736 (N_6736,N_4987,N_5879);
nor U6737 (N_6737,N_5112,N_5715);
xnor U6738 (N_6738,N_5502,N_4596);
nand U6739 (N_6739,N_5499,N_5135);
and U6740 (N_6740,N_5795,N_5292);
or U6741 (N_6741,N_5641,N_4544);
and U6742 (N_6742,N_5933,N_5286);
nand U6743 (N_6743,N_4930,N_5352);
and U6744 (N_6744,N_5475,N_5801);
and U6745 (N_6745,N_5339,N_5444);
or U6746 (N_6746,N_4500,N_5807);
xor U6747 (N_6747,N_4719,N_4917);
nand U6748 (N_6748,N_5234,N_5435);
and U6749 (N_6749,N_4655,N_5375);
nand U6750 (N_6750,N_5057,N_5873);
xnor U6751 (N_6751,N_5679,N_4669);
xor U6752 (N_6752,N_5406,N_5372);
nand U6753 (N_6753,N_4767,N_4615);
nand U6754 (N_6754,N_5171,N_5553);
nand U6755 (N_6755,N_4626,N_5014);
and U6756 (N_6756,N_5500,N_4625);
nor U6757 (N_6757,N_5197,N_5934);
and U6758 (N_6758,N_5914,N_5893);
nand U6759 (N_6759,N_5632,N_5491);
and U6760 (N_6760,N_5133,N_5887);
or U6761 (N_6761,N_4974,N_5977);
and U6762 (N_6762,N_5782,N_4730);
and U6763 (N_6763,N_4844,N_5346);
or U6764 (N_6764,N_4978,N_4812);
xnor U6765 (N_6765,N_5864,N_5403);
nor U6766 (N_6766,N_4776,N_4514);
nor U6767 (N_6767,N_5223,N_5192);
nand U6768 (N_6768,N_5383,N_5892);
or U6769 (N_6769,N_4853,N_5322);
and U6770 (N_6770,N_4566,N_5388);
nand U6771 (N_6771,N_5687,N_5766);
xnor U6772 (N_6772,N_5174,N_5776);
nand U6773 (N_6773,N_5962,N_5006);
nand U6774 (N_6774,N_4641,N_4542);
xnor U6775 (N_6775,N_5447,N_4801);
nor U6776 (N_6776,N_4594,N_5337);
and U6777 (N_6777,N_5102,N_5116);
nor U6778 (N_6778,N_4850,N_5106);
nor U6779 (N_6779,N_5626,N_4575);
and U6780 (N_6780,N_5259,N_5117);
and U6781 (N_6781,N_4953,N_4979);
or U6782 (N_6782,N_5572,N_5552);
and U6783 (N_6783,N_5956,N_4926);
and U6784 (N_6784,N_5191,N_5265);
nand U6785 (N_6785,N_4755,N_5418);
nor U6786 (N_6786,N_5734,N_5038);
nand U6787 (N_6787,N_5567,N_4877);
xor U6788 (N_6788,N_4637,N_5925);
nor U6789 (N_6789,N_5984,N_5729);
nand U6790 (N_6790,N_4651,N_5988);
or U6791 (N_6791,N_5394,N_5145);
and U6792 (N_6792,N_5844,N_4854);
or U6793 (N_6793,N_5346,N_4993);
and U6794 (N_6794,N_4934,N_5748);
and U6795 (N_6795,N_5270,N_5623);
nor U6796 (N_6796,N_5805,N_5011);
xor U6797 (N_6797,N_5886,N_5313);
nand U6798 (N_6798,N_5149,N_5420);
nor U6799 (N_6799,N_5382,N_4670);
nor U6800 (N_6800,N_5271,N_4681);
xnor U6801 (N_6801,N_5238,N_5870);
xnor U6802 (N_6802,N_5876,N_4664);
and U6803 (N_6803,N_5610,N_5555);
or U6804 (N_6804,N_4623,N_5207);
nand U6805 (N_6805,N_4661,N_5190);
nor U6806 (N_6806,N_4726,N_4946);
and U6807 (N_6807,N_5021,N_5475);
or U6808 (N_6808,N_5914,N_5714);
nand U6809 (N_6809,N_5252,N_5343);
and U6810 (N_6810,N_5875,N_4978);
nor U6811 (N_6811,N_4829,N_4658);
nor U6812 (N_6812,N_5916,N_5943);
and U6813 (N_6813,N_4999,N_4811);
nand U6814 (N_6814,N_4643,N_5658);
and U6815 (N_6815,N_5232,N_5884);
nor U6816 (N_6816,N_4589,N_4953);
and U6817 (N_6817,N_5865,N_5240);
and U6818 (N_6818,N_5847,N_5096);
and U6819 (N_6819,N_5376,N_5300);
nor U6820 (N_6820,N_5780,N_4951);
or U6821 (N_6821,N_5270,N_5648);
xnor U6822 (N_6822,N_5952,N_5864);
or U6823 (N_6823,N_5657,N_5277);
and U6824 (N_6824,N_4531,N_4740);
nor U6825 (N_6825,N_5183,N_5621);
nor U6826 (N_6826,N_5068,N_4856);
or U6827 (N_6827,N_5472,N_5539);
nor U6828 (N_6828,N_5833,N_4546);
and U6829 (N_6829,N_5477,N_4645);
nor U6830 (N_6830,N_5346,N_5053);
or U6831 (N_6831,N_4930,N_5703);
nor U6832 (N_6832,N_4822,N_5964);
nor U6833 (N_6833,N_4920,N_5570);
nand U6834 (N_6834,N_5742,N_5675);
nand U6835 (N_6835,N_5420,N_5937);
and U6836 (N_6836,N_4553,N_4985);
nand U6837 (N_6837,N_5121,N_5406);
and U6838 (N_6838,N_5975,N_5896);
nand U6839 (N_6839,N_5626,N_5389);
nand U6840 (N_6840,N_4529,N_5145);
or U6841 (N_6841,N_4834,N_5554);
and U6842 (N_6842,N_5834,N_4556);
or U6843 (N_6843,N_5931,N_4661);
or U6844 (N_6844,N_4902,N_4829);
and U6845 (N_6845,N_5346,N_5987);
xor U6846 (N_6846,N_4555,N_5711);
nor U6847 (N_6847,N_5529,N_5752);
nand U6848 (N_6848,N_5876,N_4944);
nor U6849 (N_6849,N_4518,N_5712);
or U6850 (N_6850,N_5133,N_4813);
xnor U6851 (N_6851,N_5866,N_5131);
nand U6852 (N_6852,N_5603,N_4637);
nor U6853 (N_6853,N_5192,N_4990);
or U6854 (N_6854,N_4718,N_4959);
xnor U6855 (N_6855,N_5234,N_5129);
xor U6856 (N_6856,N_5667,N_4655);
nand U6857 (N_6857,N_4881,N_5701);
and U6858 (N_6858,N_4985,N_5068);
or U6859 (N_6859,N_5997,N_5900);
xnor U6860 (N_6860,N_5447,N_4975);
or U6861 (N_6861,N_4650,N_5953);
nand U6862 (N_6862,N_5290,N_5861);
or U6863 (N_6863,N_5933,N_4701);
nor U6864 (N_6864,N_4829,N_5195);
nand U6865 (N_6865,N_5002,N_5608);
nand U6866 (N_6866,N_5879,N_5840);
nor U6867 (N_6867,N_4716,N_4984);
and U6868 (N_6868,N_5277,N_4841);
nand U6869 (N_6869,N_5784,N_5894);
nor U6870 (N_6870,N_4796,N_5842);
and U6871 (N_6871,N_4816,N_5884);
or U6872 (N_6872,N_4961,N_5446);
nor U6873 (N_6873,N_4955,N_5488);
or U6874 (N_6874,N_5459,N_5558);
or U6875 (N_6875,N_4916,N_4638);
and U6876 (N_6876,N_4924,N_5097);
and U6877 (N_6877,N_5635,N_5120);
xor U6878 (N_6878,N_5825,N_4749);
nor U6879 (N_6879,N_4586,N_5171);
nor U6880 (N_6880,N_5490,N_4539);
nand U6881 (N_6881,N_5799,N_4913);
and U6882 (N_6882,N_5493,N_5882);
and U6883 (N_6883,N_4908,N_5713);
or U6884 (N_6884,N_5747,N_4522);
or U6885 (N_6885,N_5945,N_4826);
and U6886 (N_6886,N_4983,N_5573);
nor U6887 (N_6887,N_5379,N_4666);
xor U6888 (N_6888,N_5621,N_4613);
nand U6889 (N_6889,N_5853,N_5302);
nand U6890 (N_6890,N_4794,N_4602);
nand U6891 (N_6891,N_4767,N_4801);
xor U6892 (N_6892,N_5549,N_5039);
nor U6893 (N_6893,N_5695,N_5819);
nand U6894 (N_6894,N_5585,N_5344);
and U6895 (N_6895,N_5578,N_4974);
nor U6896 (N_6896,N_5123,N_5689);
or U6897 (N_6897,N_5094,N_5848);
nor U6898 (N_6898,N_5692,N_4698);
nand U6899 (N_6899,N_5497,N_4643);
nand U6900 (N_6900,N_5495,N_5408);
and U6901 (N_6901,N_5536,N_5416);
and U6902 (N_6902,N_4702,N_4797);
nor U6903 (N_6903,N_5489,N_5899);
nand U6904 (N_6904,N_5953,N_4819);
and U6905 (N_6905,N_4600,N_4896);
and U6906 (N_6906,N_5960,N_5237);
and U6907 (N_6907,N_5767,N_5124);
nor U6908 (N_6908,N_5077,N_5228);
nor U6909 (N_6909,N_4512,N_4988);
and U6910 (N_6910,N_5862,N_4978);
or U6911 (N_6911,N_4877,N_4887);
nand U6912 (N_6912,N_5513,N_5961);
and U6913 (N_6913,N_5307,N_4929);
or U6914 (N_6914,N_5777,N_4676);
and U6915 (N_6915,N_5962,N_5213);
or U6916 (N_6916,N_5433,N_4974);
xnor U6917 (N_6917,N_5646,N_4962);
nor U6918 (N_6918,N_4572,N_4978);
and U6919 (N_6919,N_4594,N_4959);
xor U6920 (N_6920,N_5148,N_5311);
xor U6921 (N_6921,N_5132,N_5873);
xnor U6922 (N_6922,N_4905,N_4538);
nor U6923 (N_6923,N_5942,N_4841);
nand U6924 (N_6924,N_5225,N_4854);
nand U6925 (N_6925,N_5823,N_4871);
and U6926 (N_6926,N_5495,N_5256);
and U6927 (N_6927,N_5478,N_5983);
or U6928 (N_6928,N_4875,N_5346);
and U6929 (N_6929,N_5647,N_5870);
or U6930 (N_6930,N_5467,N_5051);
and U6931 (N_6931,N_4909,N_5471);
nand U6932 (N_6932,N_5132,N_4724);
or U6933 (N_6933,N_5075,N_4830);
nor U6934 (N_6934,N_5179,N_5676);
nor U6935 (N_6935,N_4940,N_5483);
nor U6936 (N_6936,N_4594,N_4785);
nand U6937 (N_6937,N_5278,N_4529);
nand U6938 (N_6938,N_5079,N_4691);
xor U6939 (N_6939,N_5283,N_4619);
and U6940 (N_6940,N_4688,N_5941);
or U6941 (N_6941,N_5808,N_5670);
nand U6942 (N_6942,N_5728,N_4933);
and U6943 (N_6943,N_5689,N_4750);
and U6944 (N_6944,N_4881,N_5225);
and U6945 (N_6945,N_5564,N_5181);
nand U6946 (N_6946,N_4904,N_4702);
xor U6947 (N_6947,N_5553,N_5565);
and U6948 (N_6948,N_5291,N_5104);
or U6949 (N_6949,N_5504,N_5056);
nand U6950 (N_6950,N_4784,N_4594);
and U6951 (N_6951,N_4732,N_4677);
or U6952 (N_6952,N_5085,N_5511);
and U6953 (N_6953,N_5894,N_4848);
xnor U6954 (N_6954,N_5525,N_4985);
and U6955 (N_6955,N_5342,N_5545);
nor U6956 (N_6956,N_5249,N_4720);
nor U6957 (N_6957,N_5725,N_5129);
and U6958 (N_6958,N_5902,N_5798);
nor U6959 (N_6959,N_4776,N_5805);
nand U6960 (N_6960,N_5057,N_4709);
or U6961 (N_6961,N_5188,N_4716);
nor U6962 (N_6962,N_5600,N_5929);
and U6963 (N_6963,N_5582,N_5805);
or U6964 (N_6964,N_5892,N_5372);
nand U6965 (N_6965,N_5080,N_5313);
and U6966 (N_6966,N_5669,N_4683);
and U6967 (N_6967,N_5543,N_5846);
nand U6968 (N_6968,N_5319,N_4909);
and U6969 (N_6969,N_4680,N_5519);
and U6970 (N_6970,N_4888,N_5207);
nor U6971 (N_6971,N_5581,N_5766);
nor U6972 (N_6972,N_4683,N_4688);
xor U6973 (N_6973,N_5447,N_5736);
nand U6974 (N_6974,N_5438,N_5264);
and U6975 (N_6975,N_5107,N_5757);
xnor U6976 (N_6976,N_5116,N_5250);
nand U6977 (N_6977,N_5656,N_4784);
and U6978 (N_6978,N_4845,N_4815);
and U6979 (N_6979,N_5721,N_4502);
or U6980 (N_6980,N_5997,N_5631);
nand U6981 (N_6981,N_5902,N_4542);
or U6982 (N_6982,N_4806,N_5965);
or U6983 (N_6983,N_5660,N_5678);
nor U6984 (N_6984,N_5676,N_5212);
or U6985 (N_6985,N_4601,N_4637);
nand U6986 (N_6986,N_5258,N_4507);
xnor U6987 (N_6987,N_5584,N_4504);
and U6988 (N_6988,N_4957,N_5690);
nand U6989 (N_6989,N_4921,N_5185);
nor U6990 (N_6990,N_4609,N_5018);
nor U6991 (N_6991,N_4952,N_4539);
and U6992 (N_6992,N_4684,N_4941);
and U6993 (N_6993,N_5256,N_5862);
nand U6994 (N_6994,N_5540,N_5376);
and U6995 (N_6995,N_4954,N_5528);
or U6996 (N_6996,N_4789,N_4960);
nor U6997 (N_6997,N_5457,N_5864);
or U6998 (N_6998,N_5002,N_5560);
xnor U6999 (N_6999,N_4621,N_4685);
nand U7000 (N_7000,N_5403,N_5527);
nand U7001 (N_7001,N_5257,N_4705);
nor U7002 (N_7002,N_5434,N_4829);
nand U7003 (N_7003,N_5433,N_4525);
nand U7004 (N_7004,N_5707,N_5552);
nor U7005 (N_7005,N_5740,N_4698);
and U7006 (N_7006,N_5145,N_5256);
and U7007 (N_7007,N_5506,N_5874);
or U7008 (N_7008,N_5458,N_5208);
nor U7009 (N_7009,N_5216,N_4535);
xor U7010 (N_7010,N_5624,N_5433);
or U7011 (N_7011,N_5786,N_4652);
or U7012 (N_7012,N_4914,N_5688);
and U7013 (N_7013,N_5107,N_5064);
nand U7014 (N_7014,N_4653,N_5925);
nand U7015 (N_7015,N_5012,N_4621);
nor U7016 (N_7016,N_5269,N_4862);
or U7017 (N_7017,N_5488,N_5315);
nor U7018 (N_7018,N_5889,N_4967);
and U7019 (N_7019,N_5962,N_5801);
or U7020 (N_7020,N_5492,N_5739);
or U7021 (N_7021,N_5409,N_4788);
and U7022 (N_7022,N_5483,N_4755);
nor U7023 (N_7023,N_4844,N_4792);
and U7024 (N_7024,N_4965,N_4876);
nor U7025 (N_7025,N_4702,N_5970);
nand U7026 (N_7026,N_5536,N_5128);
or U7027 (N_7027,N_5236,N_5547);
nor U7028 (N_7028,N_5359,N_4582);
nand U7029 (N_7029,N_5128,N_5908);
nand U7030 (N_7030,N_5944,N_5429);
and U7031 (N_7031,N_5156,N_5169);
or U7032 (N_7032,N_5265,N_5522);
nand U7033 (N_7033,N_5591,N_5100);
nor U7034 (N_7034,N_4971,N_5756);
nor U7035 (N_7035,N_5132,N_4733);
nand U7036 (N_7036,N_4662,N_5258);
or U7037 (N_7037,N_5426,N_5132);
nand U7038 (N_7038,N_5485,N_5381);
xnor U7039 (N_7039,N_5020,N_5234);
xor U7040 (N_7040,N_5132,N_5946);
or U7041 (N_7041,N_4802,N_4558);
or U7042 (N_7042,N_4882,N_5602);
nand U7043 (N_7043,N_5831,N_5232);
nor U7044 (N_7044,N_5992,N_4552);
or U7045 (N_7045,N_5940,N_5689);
and U7046 (N_7046,N_5517,N_4560);
or U7047 (N_7047,N_4614,N_5403);
and U7048 (N_7048,N_4842,N_4636);
nor U7049 (N_7049,N_4907,N_5774);
nor U7050 (N_7050,N_5733,N_4855);
nor U7051 (N_7051,N_4548,N_4955);
or U7052 (N_7052,N_5642,N_5035);
xnor U7053 (N_7053,N_4586,N_5983);
and U7054 (N_7054,N_5944,N_4754);
and U7055 (N_7055,N_5240,N_5802);
nand U7056 (N_7056,N_4895,N_4819);
and U7057 (N_7057,N_4716,N_5135);
xnor U7058 (N_7058,N_4978,N_5495);
xnor U7059 (N_7059,N_4743,N_5468);
and U7060 (N_7060,N_4756,N_5317);
nor U7061 (N_7061,N_5475,N_5073);
nand U7062 (N_7062,N_4836,N_5253);
nand U7063 (N_7063,N_5987,N_4848);
nor U7064 (N_7064,N_5513,N_4607);
nand U7065 (N_7065,N_4932,N_4937);
nor U7066 (N_7066,N_4919,N_5575);
nor U7067 (N_7067,N_5132,N_5752);
or U7068 (N_7068,N_4577,N_5840);
nand U7069 (N_7069,N_5462,N_4687);
or U7070 (N_7070,N_4850,N_5927);
and U7071 (N_7071,N_4658,N_5679);
or U7072 (N_7072,N_5781,N_5631);
nor U7073 (N_7073,N_5919,N_5132);
and U7074 (N_7074,N_5580,N_5478);
xnor U7075 (N_7075,N_4904,N_5525);
nand U7076 (N_7076,N_5298,N_5710);
and U7077 (N_7077,N_4722,N_5811);
nand U7078 (N_7078,N_5845,N_5403);
and U7079 (N_7079,N_5290,N_5174);
nor U7080 (N_7080,N_5049,N_5568);
or U7081 (N_7081,N_5172,N_5530);
or U7082 (N_7082,N_5594,N_5455);
nand U7083 (N_7083,N_5313,N_4556);
or U7084 (N_7084,N_5935,N_5837);
xnor U7085 (N_7085,N_4698,N_5936);
or U7086 (N_7086,N_4565,N_5192);
or U7087 (N_7087,N_5755,N_5708);
and U7088 (N_7088,N_4701,N_5802);
nor U7089 (N_7089,N_5149,N_5328);
nand U7090 (N_7090,N_5974,N_5901);
and U7091 (N_7091,N_5764,N_5691);
and U7092 (N_7092,N_4972,N_5994);
or U7093 (N_7093,N_4567,N_5347);
and U7094 (N_7094,N_5010,N_5052);
and U7095 (N_7095,N_5703,N_4737);
and U7096 (N_7096,N_5654,N_5074);
nor U7097 (N_7097,N_4700,N_5805);
nor U7098 (N_7098,N_4636,N_5924);
xor U7099 (N_7099,N_5386,N_4554);
nand U7100 (N_7100,N_4628,N_4538);
or U7101 (N_7101,N_4961,N_5315);
and U7102 (N_7102,N_4989,N_4834);
or U7103 (N_7103,N_5603,N_5053);
nor U7104 (N_7104,N_5087,N_5111);
xnor U7105 (N_7105,N_5662,N_5517);
nand U7106 (N_7106,N_5708,N_4981);
and U7107 (N_7107,N_5353,N_5456);
and U7108 (N_7108,N_5576,N_5639);
and U7109 (N_7109,N_5533,N_4839);
and U7110 (N_7110,N_5111,N_5592);
nand U7111 (N_7111,N_4905,N_4595);
and U7112 (N_7112,N_5674,N_5665);
and U7113 (N_7113,N_4914,N_4654);
nand U7114 (N_7114,N_5223,N_5127);
nor U7115 (N_7115,N_5250,N_5332);
nor U7116 (N_7116,N_5987,N_4722);
nor U7117 (N_7117,N_4884,N_5518);
or U7118 (N_7118,N_5105,N_4556);
nor U7119 (N_7119,N_5591,N_4841);
nand U7120 (N_7120,N_4916,N_4977);
nor U7121 (N_7121,N_4875,N_5010);
or U7122 (N_7122,N_5278,N_4622);
or U7123 (N_7123,N_4849,N_5955);
and U7124 (N_7124,N_5638,N_5204);
nor U7125 (N_7125,N_5173,N_4581);
xor U7126 (N_7126,N_4539,N_4739);
or U7127 (N_7127,N_4520,N_5331);
and U7128 (N_7128,N_5987,N_4546);
nor U7129 (N_7129,N_5266,N_5361);
and U7130 (N_7130,N_4817,N_5571);
nor U7131 (N_7131,N_4698,N_5577);
nand U7132 (N_7132,N_5728,N_5155);
or U7133 (N_7133,N_5147,N_5601);
and U7134 (N_7134,N_4844,N_4890);
or U7135 (N_7135,N_4571,N_5436);
xor U7136 (N_7136,N_5136,N_5648);
nand U7137 (N_7137,N_4770,N_5050);
or U7138 (N_7138,N_5077,N_4950);
xnor U7139 (N_7139,N_5349,N_4864);
and U7140 (N_7140,N_5281,N_5655);
nand U7141 (N_7141,N_5992,N_5337);
nor U7142 (N_7142,N_5775,N_5041);
nor U7143 (N_7143,N_5715,N_5119);
nor U7144 (N_7144,N_5218,N_5528);
nand U7145 (N_7145,N_5398,N_5692);
or U7146 (N_7146,N_5167,N_5492);
xor U7147 (N_7147,N_5920,N_5625);
and U7148 (N_7148,N_5418,N_4953);
nor U7149 (N_7149,N_4847,N_4813);
nor U7150 (N_7150,N_4694,N_4775);
or U7151 (N_7151,N_5365,N_4504);
nor U7152 (N_7152,N_5825,N_5712);
or U7153 (N_7153,N_4617,N_5634);
and U7154 (N_7154,N_5522,N_5944);
or U7155 (N_7155,N_4848,N_5397);
nand U7156 (N_7156,N_5350,N_4920);
nand U7157 (N_7157,N_4824,N_5716);
xnor U7158 (N_7158,N_5510,N_5963);
nor U7159 (N_7159,N_5879,N_4845);
nor U7160 (N_7160,N_5540,N_5971);
and U7161 (N_7161,N_5605,N_5820);
or U7162 (N_7162,N_5563,N_4910);
or U7163 (N_7163,N_5164,N_5707);
nand U7164 (N_7164,N_5741,N_5069);
and U7165 (N_7165,N_5907,N_4901);
or U7166 (N_7166,N_5482,N_5341);
xnor U7167 (N_7167,N_4505,N_5358);
nand U7168 (N_7168,N_5772,N_4679);
nand U7169 (N_7169,N_5525,N_4613);
and U7170 (N_7170,N_4620,N_5056);
and U7171 (N_7171,N_5558,N_5977);
nor U7172 (N_7172,N_4971,N_4957);
xnor U7173 (N_7173,N_5104,N_4736);
and U7174 (N_7174,N_5716,N_4869);
and U7175 (N_7175,N_4954,N_5102);
xor U7176 (N_7176,N_5909,N_5787);
and U7177 (N_7177,N_5111,N_5552);
or U7178 (N_7178,N_5953,N_4744);
nand U7179 (N_7179,N_5752,N_5398);
nand U7180 (N_7180,N_4951,N_4902);
and U7181 (N_7181,N_4525,N_5614);
or U7182 (N_7182,N_5085,N_4598);
and U7183 (N_7183,N_5220,N_4775);
nor U7184 (N_7184,N_4731,N_4595);
or U7185 (N_7185,N_5729,N_4554);
nor U7186 (N_7186,N_5090,N_5046);
nor U7187 (N_7187,N_5765,N_5939);
nand U7188 (N_7188,N_5232,N_5429);
nor U7189 (N_7189,N_5489,N_4858);
or U7190 (N_7190,N_4719,N_5279);
and U7191 (N_7191,N_5494,N_5917);
nand U7192 (N_7192,N_4543,N_5200);
nand U7193 (N_7193,N_4779,N_5483);
or U7194 (N_7194,N_5008,N_5376);
or U7195 (N_7195,N_5731,N_5362);
nor U7196 (N_7196,N_5204,N_5480);
nand U7197 (N_7197,N_5158,N_4822);
or U7198 (N_7198,N_5096,N_5936);
and U7199 (N_7199,N_5535,N_5328);
and U7200 (N_7200,N_5742,N_5628);
or U7201 (N_7201,N_4691,N_4703);
nand U7202 (N_7202,N_5285,N_4693);
and U7203 (N_7203,N_4704,N_4556);
nand U7204 (N_7204,N_5379,N_5839);
nand U7205 (N_7205,N_5875,N_5737);
and U7206 (N_7206,N_5820,N_5840);
nor U7207 (N_7207,N_4708,N_4798);
and U7208 (N_7208,N_5986,N_5633);
nor U7209 (N_7209,N_4796,N_5846);
nand U7210 (N_7210,N_5325,N_5597);
and U7211 (N_7211,N_5502,N_5002);
nand U7212 (N_7212,N_5170,N_4837);
nand U7213 (N_7213,N_5535,N_4844);
nor U7214 (N_7214,N_5175,N_5177);
xnor U7215 (N_7215,N_5636,N_4956);
nor U7216 (N_7216,N_5457,N_5170);
or U7217 (N_7217,N_5643,N_5769);
and U7218 (N_7218,N_5520,N_5667);
or U7219 (N_7219,N_5221,N_4521);
or U7220 (N_7220,N_5587,N_4672);
xor U7221 (N_7221,N_5407,N_5449);
and U7222 (N_7222,N_5780,N_5434);
or U7223 (N_7223,N_5022,N_5992);
nor U7224 (N_7224,N_4581,N_5178);
nor U7225 (N_7225,N_4626,N_5759);
or U7226 (N_7226,N_5003,N_4907);
nand U7227 (N_7227,N_4519,N_5684);
nor U7228 (N_7228,N_4575,N_5979);
nand U7229 (N_7229,N_5719,N_5439);
or U7230 (N_7230,N_5059,N_4836);
xor U7231 (N_7231,N_5012,N_5603);
or U7232 (N_7232,N_5126,N_4519);
or U7233 (N_7233,N_5420,N_4651);
or U7234 (N_7234,N_4844,N_4992);
and U7235 (N_7235,N_4714,N_4667);
or U7236 (N_7236,N_4875,N_5512);
and U7237 (N_7237,N_4612,N_4846);
or U7238 (N_7238,N_4951,N_5138);
xnor U7239 (N_7239,N_4873,N_5253);
nand U7240 (N_7240,N_4502,N_5477);
nand U7241 (N_7241,N_5490,N_5822);
xnor U7242 (N_7242,N_5492,N_4956);
or U7243 (N_7243,N_4801,N_4648);
or U7244 (N_7244,N_5819,N_4821);
nand U7245 (N_7245,N_5521,N_5071);
nor U7246 (N_7246,N_4725,N_5637);
nand U7247 (N_7247,N_5633,N_5060);
nor U7248 (N_7248,N_5876,N_5855);
nand U7249 (N_7249,N_5213,N_4770);
nand U7250 (N_7250,N_5523,N_4821);
and U7251 (N_7251,N_5022,N_5453);
nand U7252 (N_7252,N_5026,N_4622);
or U7253 (N_7253,N_5566,N_5328);
and U7254 (N_7254,N_5919,N_5627);
nor U7255 (N_7255,N_5433,N_5152);
and U7256 (N_7256,N_4709,N_5920);
xnor U7257 (N_7257,N_5266,N_5546);
or U7258 (N_7258,N_5840,N_4761);
xnor U7259 (N_7259,N_5345,N_5542);
xor U7260 (N_7260,N_4544,N_4968);
and U7261 (N_7261,N_5036,N_5790);
nor U7262 (N_7262,N_5731,N_5501);
and U7263 (N_7263,N_5948,N_4505);
xor U7264 (N_7264,N_5888,N_5429);
nand U7265 (N_7265,N_5828,N_5874);
and U7266 (N_7266,N_4662,N_4645);
or U7267 (N_7267,N_5322,N_5663);
or U7268 (N_7268,N_5035,N_5492);
nor U7269 (N_7269,N_5279,N_5199);
nand U7270 (N_7270,N_4987,N_5450);
nor U7271 (N_7271,N_5520,N_4552);
and U7272 (N_7272,N_4973,N_5835);
or U7273 (N_7273,N_4707,N_5305);
xor U7274 (N_7274,N_5817,N_5069);
and U7275 (N_7275,N_4732,N_5293);
nor U7276 (N_7276,N_5853,N_5996);
nor U7277 (N_7277,N_5987,N_4838);
xor U7278 (N_7278,N_5801,N_5059);
nor U7279 (N_7279,N_5997,N_5050);
nand U7280 (N_7280,N_5086,N_4854);
and U7281 (N_7281,N_4648,N_4501);
nor U7282 (N_7282,N_5612,N_5767);
and U7283 (N_7283,N_4534,N_4631);
nor U7284 (N_7284,N_5995,N_5722);
and U7285 (N_7285,N_5953,N_5569);
nor U7286 (N_7286,N_5111,N_5132);
nand U7287 (N_7287,N_5648,N_5137);
and U7288 (N_7288,N_4728,N_5985);
xor U7289 (N_7289,N_4933,N_5551);
and U7290 (N_7290,N_4765,N_5040);
or U7291 (N_7291,N_4787,N_5893);
nor U7292 (N_7292,N_5254,N_5935);
and U7293 (N_7293,N_5393,N_5273);
xnor U7294 (N_7294,N_4701,N_5408);
xnor U7295 (N_7295,N_5555,N_5604);
or U7296 (N_7296,N_5597,N_5069);
nor U7297 (N_7297,N_4778,N_4746);
nor U7298 (N_7298,N_5263,N_5256);
nand U7299 (N_7299,N_5350,N_5873);
and U7300 (N_7300,N_5056,N_5759);
nor U7301 (N_7301,N_4985,N_4737);
nor U7302 (N_7302,N_5201,N_5323);
nand U7303 (N_7303,N_5758,N_5708);
nand U7304 (N_7304,N_4859,N_4958);
or U7305 (N_7305,N_5677,N_5941);
nor U7306 (N_7306,N_4983,N_5525);
nor U7307 (N_7307,N_5350,N_5001);
nand U7308 (N_7308,N_5248,N_5604);
nor U7309 (N_7309,N_5251,N_5859);
nor U7310 (N_7310,N_4927,N_5802);
nor U7311 (N_7311,N_5758,N_5393);
or U7312 (N_7312,N_4948,N_5746);
or U7313 (N_7313,N_4813,N_5763);
nand U7314 (N_7314,N_4998,N_5275);
xnor U7315 (N_7315,N_5003,N_5007);
nand U7316 (N_7316,N_5941,N_5643);
and U7317 (N_7317,N_5600,N_4968);
nand U7318 (N_7318,N_5564,N_4717);
nor U7319 (N_7319,N_4672,N_4999);
nor U7320 (N_7320,N_4572,N_4868);
xor U7321 (N_7321,N_5039,N_5708);
nand U7322 (N_7322,N_5235,N_5899);
nand U7323 (N_7323,N_4936,N_5447);
nand U7324 (N_7324,N_4783,N_5695);
nand U7325 (N_7325,N_5673,N_5432);
and U7326 (N_7326,N_4921,N_5533);
and U7327 (N_7327,N_5388,N_5038);
nand U7328 (N_7328,N_5051,N_5351);
and U7329 (N_7329,N_5785,N_5730);
or U7330 (N_7330,N_5648,N_5042);
nor U7331 (N_7331,N_4899,N_4747);
nand U7332 (N_7332,N_5817,N_5958);
xor U7333 (N_7333,N_5865,N_5377);
xor U7334 (N_7334,N_5108,N_5325);
nand U7335 (N_7335,N_5707,N_5622);
nand U7336 (N_7336,N_5621,N_4778);
or U7337 (N_7337,N_4727,N_5696);
or U7338 (N_7338,N_5333,N_5904);
nor U7339 (N_7339,N_4872,N_5868);
nand U7340 (N_7340,N_5778,N_5708);
nand U7341 (N_7341,N_5529,N_5032);
nor U7342 (N_7342,N_5316,N_4912);
and U7343 (N_7343,N_5500,N_5374);
nor U7344 (N_7344,N_5458,N_5432);
nor U7345 (N_7345,N_5639,N_4709);
or U7346 (N_7346,N_4786,N_4923);
nor U7347 (N_7347,N_5970,N_4647);
nor U7348 (N_7348,N_4756,N_4510);
nand U7349 (N_7349,N_5096,N_4874);
or U7350 (N_7350,N_4815,N_5700);
xnor U7351 (N_7351,N_5421,N_4850);
nor U7352 (N_7352,N_5043,N_5967);
and U7353 (N_7353,N_4511,N_4570);
nor U7354 (N_7354,N_5016,N_4922);
nor U7355 (N_7355,N_5445,N_4662);
nand U7356 (N_7356,N_5900,N_5409);
nor U7357 (N_7357,N_5468,N_5741);
or U7358 (N_7358,N_5851,N_5676);
xor U7359 (N_7359,N_4692,N_4559);
nand U7360 (N_7360,N_5321,N_5585);
and U7361 (N_7361,N_4780,N_5304);
or U7362 (N_7362,N_5585,N_5937);
nor U7363 (N_7363,N_5906,N_5970);
nor U7364 (N_7364,N_5688,N_4989);
and U7365 (N_7365,N_5115,N_5076);
or U7366 (N_7366,N_4500,N_4933);
or U7367 (N_7367,N_5431,N_4919);
nand U7368 (N_7368,N_5461,N_5633);
and U7369 (N_7369,N_5311,N_5241);
or U7370 (N_7370,N_4817,N_4807);
or U7371 (N_7371,N_4799,N_4899);
nor U7372 (N_7372,N_5701,N_4964);
and U7373 (N_7373,N_4703,N_4814);
nand U7374 (N_7374,N_4820,N_4521);
nor U7375 (N_7375,N_4624,N_4927);
and U7376 (N_7376,N_4696,N_5833);
nor U7377 (N_7377,N_5060,N_5613);
and U7378 (N_7378,N_4574,N_5660);
xor U7379 (N_7379,N_5906,N_5480);
nor U7380 (N_7380,N_4928,N_4564);
xnor U7381 (N_7381,N_5910,N_5101);
and U7382 (N_7382,N_5365,N_5227);
nand U7383 (N_7383,N_5331,N_4945);
nor U7384 (N_7384,N_4909,N_4969);
nand U7385 (N_7385,N_4609,N_4962);
or U7386 (N_7386,N_4818,N_5723);
or U7387 (N_7387,N_5965,N_4755);
and U7388 (N_7388,N_4586,N_5685);
and U7389 (N_7389,N_5976,N_5816);
nand U7390 (N_7390,N_5049,N_5381);
and U7391 (N_7391,N_5420,N_4971);
or U7392 (N_7392,N_4988,N_5462);
and U7393 (N_7393,N_4657,N_5407);
nand U7394 (N_7394,N_4848,N_4952);
nor U7395 (N_7395,N_5778,N_4958);
and U7396 (N_7396,N_4838,N_5476);
nor U7397 (N_7397,N_5806,N_4688);
nand U7398 (N_7398,N_4572,N_4871);
or U7399 (N_7399,N_5960,N_5568);
and U7400 (N_7400,N_5580,N_4641);
nor U7401 (N_7401,N_4958,N_5405);
nand U7402 (N_7402,N_5280,N_5601);
and U7403 (N_7403,N_5092,N_5937);
nand U7404 (N_7404,N_5182,N_5345);
xnor U7405 (N_7405,N_5039,N_5975);
nand U7406 (N_7406,N_5597,N_5005);
and U7407 (N_7407,N_5339,N_5808);
and U7408 (N_7408,N_5149,N_5049);
nor U7409 (N_7409,N_5226,N_5292);
nand U7410 (N_7410,N_5346,N_4718);
or U7411 (N_7411,N_4807,N_5538);
xnor U7412 (N_7412,N_4698,N_5959);
xnor U7413 (N_7413,N_5883,N_5941);
and U7414 (N_7414,N_4718,N_5049);
nor U7415 (N_7415,N_5057,N_5254);
or U7416 (N_7416,N_5117,N_5113);
or U7417 (N_7417,N_4700,N_5582);
nand U7418 (N_7418,N_5023,N_5001);
nor U7419 (N_7419,N_4733,N_5006);
nor U7420 (N_7420,N_4600,N_5876);
xor U7421 (N_7421,N_5251,N_5618);
nand U7422 (N_7422,N_4892,N_4752);
or U7423 (N_7423,N_4606,N_5207);
and U7424 (N_7424,N_5156,N_5343);
nand U7425 (N_7425,N_5395,N_4734);
xnor U7426 (N_7426,N_5025,N_4744);
and U7427 (N_7427,N_5008,N_5197);
and U7428 (N_7428,N_5058,N_5460);
nand U7429 (N_7429,N_5959,N_5873);
nand U7430 (N_7430,N_5132,N_5407);
nor U7431 (N_7431,N_4759,N_5959);
nor U7432 (N_7432,N_4639,N_4715);
and U7433 (N_7433,N_5682,N_5353);
or U7434 (N_7434,N_4877,N_4829);
nand U7435 (N_7435,N_4850,N_5398);
or U7436 (N_7436,N_4724,N_5187);
xnor U7437 (N_7437,N_4764,N_5792);
nor U7438 (N_7438,N_4692,N_5804);
nor U7439 (N_7439,N_5100,N_5718);
or U7440 (N_7440,N_4531,N_4897);
nor U7441 (N_7441,N_4823,N_4630);
nand U7442 (N_7442,N_4813,N_5144);
and U7443 (N_7443,N_5973,N_4984);
or U7444 (N_7444,N_5618,N_5574);
or U7445 (N_7445,N_5123,N_4854);
and U7446 (N_7446,N_4737,N_5753);
and U7447 (N_7447,N_5480,N_5756);
xnor U7448 (N_7448,N_5367,N_4902);
nand U7449 (N_7449,N_5556,N_4917);
nor U7450 (N_7450,N_4585,N_5611);
and U7451 (N_7451,N_4943,N_5395);
and U7452 (N_7452,N_4539,N_4839);
nand U7453 (N_7453,N_4626,N_5546);
nor U7454 (N_7454,N_5438,N_4534);
nor U7455 (N_7455,N_5945,N_4866);
and U7456 (N_7456,N_5512,N_4670);
nand U7457 (N_7457,N_4610,N_5944);
or U7458 (N_7458,N_5194,N_4657);
xnor U7459 (N_7459,N_5178,N_5342);
or U7460 (N_7460,N_4719,N_5641);
nand U7461 (N_7461,N_5690,N_5639);
and U7462 (N_7462,N_5709,N_5937);
or U7463 (N_7463,N_5914,N_5100);
xor U7464 (N_7464,N_5596,N_4768);
or U7465 (N_7465,N_5550,N_5001);
and U7466 (N_7466,N_5356,N_4592);
and U7467 (N_7467,N_4935,N_5398);
nand U7468 (N_7468,N_4555,N_5286);
and U7469 (N_7469,N_5302,N_5899);
nand U7470 (N_7470,N_4907,N_4864);
or U7471 (N_7471,N_4570,N_5965);
and U7472 (N_7472,N_4822,N_5411);
nor U7473 (N_7473,N_4741,N_5946);
nor U7474 (N_7474,N_5910,N_5117);
nand U7475 (N_7475,N_5601,N_5312);
nand U7476 (N_7476,N_5778,N_5610);
nor U7477 (N_7477,N_5952,N_5137);
and U7478 (N_7478,N_5628,N_4830);
or U7479 (N_7479,N_4743,N_5289);
and U7480 (N_7480,N_5595,N_5254);
nor U7481 (N_7481,N_5393,N_5394);
xor U7482 (N_7482,N_5710,N_5568);
or U7483 (N_7483,N_5173,N_5426);
xnor U7484 (N_7484,N_5822,N_5928);
xnor U7485 (N_7485,N_4981,N_4696);
nor U7486 (N_7486,N_5705,N_5940);
nand U7487 (N_7487,N_4956,N_5330);
and U7488 (N_7488,N_5541,N_4646);
nand U7489 (N_7489,N_5446,N_5722);
xnor U7490 (N_7490,N_5963,N_5057);
nand U7491 (N_7491,N_5531,N_5754);
xnor U7492 (N_7492,N_5890,N_5560);
and U7493 (N_7493,N_5328,N_5076);
nand U7494 (N_7494,N_5878,N_4872);
nor U7495 (N_7495,N_5163,N_5305);
nand U7496 (N_7496,N_5055,N_4537);
and U7497 (N_7497,N_5766,N_5110);
nor U7498 (N_7498,N_5675,N_5187);
and U7499 (N_7499,N_5321,N_5056);
nor U7500 (N_7500,N_6285,N_6916);
nand U7501 (N_7501,N_7108,N_6010);
or U7502 (N_7502,N_6815,N_6337);
or U7503 (N_7503,N_6401,N_6839);
or U7504 (N_7504,N_6366,N_7416);
nand U7505 (N_7505,N_6968,N_6866);
or U7506 (N_7506,N_7339,N_7408);
nand U7507 (N_7507,N_6498,N_6963);
or U7508 (N_7508,N_6153,N_6579);
and U7509 (N_7509,N_6521,N_6376);
and U7510 (N_7510,N_6977,N_6900);
nor U7511 (N_7511,N_6096,N_7298);
or U7512 (N_7512,N_7326,N_7097);
or U7513 (N_7513,N_7386,N_6501);
or U7514 (N_7514,N_6591,N_6301);
or U7515 (N_7515,N_7224,N_6193);
nand U7516 (N_7516,N_6294,N_6592);
nor U7517 (N_7517,N_6621,N_6039);
xnor U7518 (N_7518,N_7016,N_6251);
nor U7519 (N_7519,N_7267,N_6713);
and U7520 (N_7520,N_7367,N_6563);
or U7521 (N_7521,N_6457,N_7289);
nor U7522 (N_7522,N_6038,N_6372);
nand U7523 (N_7523,N_6500,N_6090);
and U7524 (N_7524,N_6583,N_6092);
or U7525 (N_7525,N_6303,N_6821);
nor U7526 (N_7526,N_7182,N_6252);
nand U7527 (N_7527,N_7363,N_6857);
nor U7528 (N_7528,N_6156,N_6868);
xor U7529 (N_7529,N_6256,N_6982);
nand U7530 (N_7530,N_6031,N_6249);
xor U7531 (N_7531,N_7469,N_7472);
nand U7532 (N_7532,N_7093,N_7112);
or U7533 (N_7533,N_6912,N_6082);
nand U7534 (N_7534,N_6272,N_6177);
nor U7535 (N_7535,N_6551,N_6433);
nor U7536 (N_7536,N_7196,N_7389);
or U7537 (N_7537,N_6605,N_6195);
nand U7538 (N_7538,N_6748,N_6232);
xor U7539 (N_7539,N_6012,N_7414);
nand U7540 (N_7540,N_7448,N_6850);
xnor U7541 (N_7541,N_6679,N_6130);
or U7542 (N_7542,N_6684,N_6469);
nor U7543 (N_7543,N_7418,N_7211);
and U7544 (N_7544,N_6657,N_6577);
and U7545 (N_7545,N_7316,N_6479);
and U7546 (N_7546,N_6216,N_6336);
and U7547 (N_7547,N_7085,N_7336);
and U7548 (N_7548,N_6856,N_6844);
or U7549 (N_7549,N_6631,N_6400);
nor U7550 (N_7550,N_6833,N_6518);
nand U7551 (N_7551,N_7406,N_6851);
or U7552 (N_7552,N_6890,N_6261);
or U7553 (N_7553,N_6598,N_7475);
nor U7554 (N_7554,N_6978,N_6021);
or U7555 (N_7555,N_7137,N_6179);
nand U7556 (N_7556,N_7461,N_7338);
or U7557 (N_7557,N_7059,N_6543);
and U7558 (N_7558,N_6842,N_6753);
nand U7559 (N_7559,N_6765,N_6064);
nor U7560 (N_7560,N_7038,N_6791);
xor U7561 (N_7561,N_6192,N_7420);
and U7562 (N_7562,N_6528,N_6965);
nand U7563 (N_7563,N_7006,N_6248);
and U7564 (N_7564,N_6489,N_6594);
nor U7565 (N_7565,N_6808,N_7191);
xnor U7566 (N_7566,N_6310,N_6752);
nand U7567 (N_7567,N_6873,N_6393);
and U7568 (N_7568,N_6969,N_7307);
nand U7569 (N_7569,N_6661,N_7240);
nand U7570 (N_7570,N_6065,N_6711);
xnor U7571 (N_7571,N_6229,N_6120);
nor U7572 (N_7572,N_7319,N_6172);
or U7573 (N_7573,N_7257,N_6107);
and U7574 (N_7574,N_6874,N_6472);
or U7575 (N_7575,N_7403,N_6585);
or U7576 (N_7576,N_6214,N_6914);
nand U7577 (N_7577,N_6390,N_6576);
xnor U7578 (N_7578,N_7467,N_6690);
or U7579 (N_7579,N_6237,N_6678);
and U7580 (N_7580,N_7046,N_7165);
nor U7581 (N_7581,N_6486,N_6847);
and U7582 (N_7582,N_7050,N_6266);
or U7583 (N_7583,N_6228,N_6902);
nor U7584 (N_7584,N_7049,N_6556);
and U7585 (N_7585,N_6779,N_6204);
or U7586 (N_7586,N_7183,N_6407);
nand U7587 (N_7587,N_6328,N_6643);
and U7588 (N_7588,N_6731,N_7134);
and U7589 (N_7589,N_6616,N_6276);
and U7590 (N_7590,N_6097,N_7215);
nand U7591 (N_7591,N_6386,N_6478);
nor U7592 (N_7592,N_6801,N_6614);
xnor U7593 (N_7593,N_6320,N_7436);
or U7594 (N_7594,N_6408,N_7082);
and U7595 (N_7595,N_7306,N_6960);
nand U7596 (N_7596,N_7478,N_6812);
and U7597 (N_7597,N_6829,N_7352);
and U7598 (N_7598,N_6171,N_7263);
or U7599 (N_7599,N_6789,N_6625);
or U7600 (N_7600,N_6766,N_7299);
nor U7601 (N_7601,N_6483,N_6936);
nand U7602 (N_7602,N_6988,N_6410);
and U7603 (N_7603,N_6143,N_6298);
xnor U7604 (N_7604,N_7325,N_6203);
nand U7605 (N_7605,N_6878,N_6106);
nand U7606 (N_7606,N_6194,N_7243);
and U7607 (N_7607,N_6326,N_7491);
and U7608 (N_7608,N_7041,N_7375);
or U7609 (N_7609,N_7370,N_6609);
nand U7610 (N_7610,N_6973,N_6663);
and U7611 (N_7611,N_6206,N_6058);
xnor U7612 (N_7612,N_6072,N_7255);
nand U7613 (N_7613,N_7277,N_6324);
nor U7614 (N_7614,N_6353,N_7492);
nand U7615 (N_7615,N_6901,N_6024);
or U7616 (N_7616,N_6265,N_6370);
or U7617 (N_7617,N_7178,N_7258);
nand U7618 (N_7618,N_7139,N_6419);
and U7619 (N_7619,N_6841,N_6710);
or U7620 (N_7620,N_7479,N_6159);
nand U7621 (N_7621,N_6155,N_6702);
or U7622 (N_7622,N_6131,N_7008);
nor U7623 (N_7623,N_6539,N_6806);
and U7624 (N_7624,N_6550,N_6468);
nand U7625 (N_7625,N_7252,N_7042);
nor U7626 (N_7626,N_6638,N_6163);
and U7627 (N_7627,N_6384,N_6721);
xor U7628 (N_7628,N_7433,N_7355);
or U7629 (N_7629,N_6431,N_7162);
or U7630 (N_7630,N_6762,N_6749);
nand U7631 (N_7631,N_6552,N_7397);
nor U7632 (N_7632,N_6785,N_6420);
or U7633 (N_7633,N_6567,N_7206);
and U7634 (N_7634,N_6444,N_6746);
nand U7635 (N_7635,N_6682,N_6040);
xor U7636 (N_7636,N_6817,N_7413);
nand U7637 (N_7637,N_6819,N_7264);
and U7638 (N_7638,N_6627,N_6146);
xor U7639 (N_7639,N_7309,N_6388);
or U7640 (N_7640,N_7081,N_7466);
and U7641 (N_7641,N_7213,N_7254);
nand U7642 (N_7642,N_6102,N_6547);
nor U7643 (N_7643,N_7207,N_7174);
and U7644 (N_7644,N_6626,N_7455);
or U7645 (N_7645,N_7158,N_6707);
nand U7646 (N_7646,N_6755,N_6774);
or U7647 (N_7647,N_6473,N_6318);
and U7648 (N_7648,N_7036,N_7075);
or U7649 (N_7649,N_6076,N_7440);
and U7650 (N_7650,N_7321,N_6920);
or U7651 (N_7651,N_6818,N_7331);
and U7652 (N_7652,N_6332,N_6955);
nor U7653 (N_7653,N_6128,N_6295);
nand U7654 (N_7654,N_7171,N_7179);
or U7655 (N_7655,N_7166,N_7381);
nor U7656 (N_7656,N_6083,N_6695);
nand U7657 (N_7657,N_6828,N_6454);
nor U7658 (N_7658,N_6279,N_7320);
nand U7659 (N_7659,N_6150,N_6321);
nand U7660 (N_7660,N_6830,N_6763);
or U7661 (N_7661,N_6344,N_7281);
or U7662 (N_7662,N_6913,N_6436);
nand U7663 (N_7663,N_6079,N_6043);
nand U7664 (N_7664,N_6198,N_6964);
nand U7665 (N_7665,N_7113,N_7117);
nor U7666 (N_7666,N_6768,N_7044);
nor U7667 (N_7667,N_6549,N_6932);
xnor U7668 (N_7668,N_6933,N_6619);
nand U7669 (N_7669,N_7452,N_7067);
nand U7670 (N_7670,N_6115,N_7454);
and U7671 (N_7671,N_7032,N_6354);
and U7672 (N_7672,N_6464,N_6374);
xnor U7673 (N_7673,N_6787,N_6597);
nor U7674 (N_7674,N_6009,N_7251);
or U7675 (N_7675,N_6693,N_7157);
and U7676 (N_7676,N_7421,N_7245);
nor U7677 (N_7677,N_6554,N_6796);
nand U7678 (N_7678,N_6441,N_6425);
and U7679 (N_7679,N_6290,N_6944);
xnor U7680 (N_7680,N_7221,N_6775);
nor U7681 (N_7681,N_6646,N_7177);
nor U7682 (N_7682,N_7017,N_6906);
and U7683 (N_7683,N_6312,N_6943);
nand U7684 (N_7684,N_6300,N_7026);
nor U7685 (N_7685,N_7283,N_6673);
xnor U7686 (N_7686,N_6329,N_6217);
and U7687 (N_7687,N_6381,N_6523);
nand U7688 (N_7688,N_6529,N_7404);
nor U7689 (N_7689,N_6223,N_6896);
xor U7690 (N_7690,N_6451,N_6687);
nor U7691 (N_7691,N_7147,N_6046);
and U7692 (N_7692,N_6398,N_6101);
and U7693 (N_7693,N_6306,N_6089);
or U7694 (N_7694,N_6602,N_7099);
or U7695 (N_7695,N_6481,N_7280);
nor U7696 (N_7696,N_6289,N_7148);
nand U7697 (N_7697,N_6221,N_6729);
and U7698 (N_7698,N_6091,N_6145);
and U7699 (N_7699,N_6185,N_7344);
nor U7700 (N_7700,N_6049,N_6772);
xnor U7701 (N_7701,N_7248,N_6647);
or U7702 (N_7702,N_6377,N_6892);
or U7703 (N_7703,N_6477,N_6174);
xor U7704 (N_7704,N_7119,N_6604);
and U7705 (N_7705,N_7218,N_6509);
nor U7706 (N_7706,N_7458,N_7365);
or U7707 (N_7707,N_7069,N_6532);
and U7708 (N_7708,N_6650,N_6396);
or U7709 (N_7709,N_6971,N_6334);
or U7710 (N_7710,N_7347,N_7062);
nor U7711 (N_7711,N_7378,N_6862);
nand U7712 (N_7712,N_6720,N_6241);
or U7713 (N_7713,N_6608,N_6093);
and U7714 (N_7714,N_6582,N_6356);
or U7715 (N_7715,N_6792,N_7229);
or U7716 (N_7716,N_7031,N_6607);
nor U7717 (N_7717,N_7053,N_7285);
nor U7718 (N_7718,N_6365,N_6267);
nand U7719 (N_7719,N_6234,N_6861);
or U7720 (N_7720,N_7095,N_6846);
nor U7721 (N_7721,N_7350,N_6984);
or U7722 (N_7722,N_7393,N_6777);
nand U7723 (N_7723,N_7203,N_6181);
nand U7724 (N_7724,N_6446,N_6404);
and U7725 (N_7725,N_6149,N_6974);
or U7726 (N_7726,N_6680,N_6416);
and U7727 (N_7727,N_6235,N_6421);
or U7728 (N_7728,N_6000,N_7156);
nand U7729 (N_7729,N_7411,N_7315);
nor U7730 (N_7730,N_6210,N_7002);
nand U7731 (N_7731,N_6893,N_7223);
and U7732 (N_7732,N_6613,N_6423);
nand U7733 (N_7733,N_6593,N_7020);
xnor U7734 (N_7734,N_7018,N_6259);
xnor U7735 (N_7735,N_6013,N_6075);
or U7736 (N_7736,N_6880,N_7483);
nor U7737 (N_7737,N_7051,N_7068);
and U7738 (N_7738,N_6709,N_6599);
and U7739 (N_7739,N_6986,N_6480);
nand U7740 (N_7740,N_6200,N_6726);
nor U7741 (N_7741,N_6531,N_7482);
and U7742 (N_7742,N_7311,N_6962);
or U7743 (N_7743,N_6751,N_7402);
nor U7744 (N_7744,N_6826,N_7003);
or U7745 (N_7745,N_6907,N_6277);
or U7746 (N_7746,N_7253,N_6516);
nor U7747 (N_7747,N_6784,N_6142);
and U7748 (N_7748,N_6242,N_6471);
and U7749 (N_7749,N_6522,N_6226);
nand U7750 (N_7750,N_6827,N_6224);
and U7751 (N_7751,N_6389,N_6628);
or U7752 (N_7752,N_6568,N_6794);
nor U7753 (N_7753,N_7133,N_6692);
nand U7754 (N_7754,N_6519,N_7159);
xnor U7755 (N_7755,N_6342,N_6507);
nor U7756 (N_7756,N_6909,N_6871);
nor U7757 (N_7757,N_7300,N_6165);
nor U7758 (N_7758,N_6173,N_6849);
and U7759 (N_7759,N_7219,N_6168);
and U7760 (N_7760,N_6975,N_7040);
and U7761 (N_7761,N_6257,N_6566);
xnor U7762 (N_7762,N_6254,N_6668);
xor U7763 (N_7763,N_6526,N_6188);
or U7764 (N_7764,N_7357,N_7318);
nor U7765 (N_7765,N_7314,N_6681);
nor U7766 (N_7766,N_6315,N_6688);
nor U7767 (N_7767,N_7362,N_7324);
and U7768 (N_7768,N_6428,N_6976);
nand U7769 (N_7769,N_6855,N_6073);
or U7770 (N_7770,N_6280,N_6927);
nor U7771 (N_7771,N_7185,N_6345);
nand U7772 (N_7772,N_6028,N_7235);
or U7773 (N_7773,N_6415,N_7019);
nand U7774 (N_7774,N_7234,N_6760);
nor U7775 (N_7775,N_7197,N_6564);
and U7776 (N_7776,N_6233,N_7333);
xnor U7777 (N_7777,N_6135,N_7232);
nand U7778 (N_7778,N_7138,N_6184);
or U7779 (N_7779,N_7380,N_6080);
or U7780 (N_7780,N_6284,N_6382);
nand U7781 (N_7781,N_6026,N_6020);
and U7782 (N_7782,N_7072,N_6459);
nor U7783 (N_7783,N_7023,N_7084);
and U7784 (N_7784,N_7497,N_6050);
nand U7785 (N_7785,N_7463,N_6343);
nand U7786 (N_7786,N_6967,N_7341);
xnor U7787 (N_7787,N_6525,N_7401);
or U7788 (N_7788,N_7180,N_6595);
nor U7789 (N_7789,N_6570,N_6816);
or U7790 (N_7790,N_6439,N_6007);
nor U7791 (N_7791,N_6956,N_7163);
nand U7792 (N_7792,N_6641,N_6905);
nor U7793 (N_7793,N_6623,N_6924);
nor U7794 (N_7794,N_7494,N_6700);
and U7795 (N_7795,N_6124,N_7390);
nor U7796 (N_7796,N_6961,N_6837);
and U7797 (N_7797,N_6704,N_7190);
and U7798 (N_7798,N_6581,N_7334);
nor U7799 (N_7799,N_6744,N_6652);
or U7800 (N_7800,N_6739,N_6317);
xnor U7801 (N_7801,N_6660,N_7371);
and U7802 (N_7802,N_7110,N_7058);
and U7803 (N_7803,N_7192,N_6994);
nand U7804 (N_7804,N_6898,N_6843);
nand U7805 (N_7805,N_6771,N_6066);
xnor U7806 (N_7806,N_6085,N_6741);
nand U7807 (N_7807,N_6019,N_6948);
and U7808 (N_7808,N_7278,N_6456);
xor U7809 (N_7809,N_7122,N_6671);
nand U7810 (N_7810,N_7230,N_7426);
nor U7811 (N_7811,N_7188,N_7181);
or U7812 (N_7812,N_7290,N_6895);
nand U7813 (N_7813,N_7176,N_7091);
nand U7814 (N_7814,N_6610,N_6985);
nor U7815 (N_7815,N_6781,N_6455);
and U7816 (N_7816,N_7260,N_6848);
xnor U7817 (N_7817,N_6411,N_6716);
and U7818 (N_7818,N_6190,N_6394);
or U7819 (N_7819,N_7312,N_6574);
nor U7820 (N_7820,N_6718,N_6016);
and U7821 (N_7821,N_6998,N_7246);
nor U7822 (N_7822,N_6508,N_7425);
nor U7823 (N_7823,N_6029,N_6392);
nand U7824 (N_7824,N_6487,N_6118);
nor U7825 (N_7825,N_6001,N_6903);
nor U7826 (N_7826,N_6418,N_7202);
or U7827 (N_7827,N_7237,N_6689);
and U7828 (N_7828,N_6018,N_6653);
or U7829 (N_7829,N_7087,N_6078);
nand U7830 (N_7830,N_6575,N_6109);
and U7831 (N_7831,N_6904,N_6557);
nand U7832 (N_7832,N_6778,N_7010);
nor U7833 (N_7833,N_7037,N_6864);
or U7834 (N_7834,N_7310,N_6544);
nor U7835 (N_7835,N_6559,N_7427);
nor U7836 (N_7836,N_7111,N_6735);
or U7837 (N_7837,N_6450,N_6350);
nor U7838 (N_7838,N_6669,N_7453);
nand U7839 (N_7839,N_7399,N_6546);
nor U7840 (N_7840,N_6629,N_6644);
and U7841 (N_7841,N_6141,N_7377);
or U7842 (N_7842,N_7236,N_7129);
and U7843 (N_7843,N_6449,N_7261);
and U7844 (N_7844,N_7198,N_6447);
or U7845 (N_7845,N_7282,N_6225);
nor U7846 (N_7846,N_7445,N_6802);
and U7847 (N_7847,N_6211,N_6151);
nand U7848 (N_7848,N_6725,N_6887);
or U7849 (N_7849,N_6612,N_6513);
nand U7850 (N_7850,N_6686,N_7431);
and U7851 (N_7851,N_7275,N_7287);
nor U7852 (N_7852,N_7126,N_6283);
and U7853 (N_7853,N_6139,N_6346);
and U7854 (N_7854,N_6137,N_7106);
and U7855 (N_7855,N_7101,N_7313);
and U7856 (N_7856,N_6872,N_6160);
nor U7857 (N_7857,N_6402,N_6706);
xor U7858 (N_7858,N_6510,N_7271);
xnor U7859 (N_7859,N_6723,N_6304);
or U7860 (N_7860,N_6341,N_6852);
nand U7861 (N_7861,N_7276,N_6157);
and U7862 (N_7862,N_7410,N_7109);
and U7863 (N_7863,N_7079,N_7268);
nor U7864 (N_7864,N_6213,N_6972);
xnor U7865 (N_7865,N_6790,N_6061);
nand U7866 (N_7866,N_6877,N_7043);
nor U7867 (N_7867,N_6170,N_7142);
nand U7868 (N_7868,N_6103,N_7291);
xor U7869 (N_7869,N_7273,N_6783);
nor U7870 (N_7870,N_7173,N_7118);
xnor U7871 (N_7871,N_7439,N_6931);
nand U7872 (N_7872,N_6712,N_6536);
nor U7873 (N_7873,N_6245,N_6127);
or U7874 (N_7874,N_6732,N_6399);
nand U7875 (N_7875,N_6011,N_6297);
or U7876 (N_7876,N_6045,N_7490);
or U7877 (N_7877,N_7358,N_7394);
nand U7878 (N_7878,N_6182,N_6189);
nand U7879 (N_7879,N_6426,N_7152);
and U7880 (N_7880,N_7353,N_6558);
xnor U7881 (N_7881,N_6035,N_6077);
nand U7882 (N_7882,N_6606,N_7021);
nor U7883 (N_7883,N_6664,N_6809);
nand U7884 (N_7884,N_7373,N_6496);
xor U7885 (N_7885,N_7056,N_6520);
and U7886 (N_7886,N_6600,N_6832);
nor U7887 (N_7887,N_6201,N_6260);
nor U7888 (N_7888,N_6022,N_7356);
nor U7889 (N_7889,N_6470,N_7132);
nand U7890 (N_7890,N_6938,N_6939);
or U7891 (N_7891,N_7456,N_7214);
xnor U7892 (N_7892,N_7366,N_6957);
or U7893 (N_7893,N_6950,N_7130);
nand U7894 (N_7894,N_7167,N_6497);
or U7895 (N_7895,N_6838,N_6129);
and U7896 (N_7896,N_6351,N_6367);
or U7897 (N_7897,N_6152,N_6738);
xor U7898 (N_7898,N_6331,N_7330);
nand U7899 (N_7899,N_7028,N_6070);
and U7900 (N_7900,N_7265,N_6466);
nor U7901 (N_7901,N_6268,N_7470);
nor U7902 (N_7902,N_7337,N_6383);
or U7903 (N_7903,N_6624,N_6946);
nand U7904 (N_7904,N_6275,N_6474);
nand U7905 (N_7905,N_6349,N_6287);
nand U7906 (N_7906,N_6705,N_6067);
nand U7907 (N_7907,N_7231,N_6945);
nor U7908 (N_7908,N_6807,N_6915);
nor U7909 (N_7909,N_7462,N_7272);
and U7910 (N_7910,N_7070,N_6462);
and U7911 (N_7911,N_6959,N_7328);
or U7912 (N_7912,N_6541,N_7088);
xor U7913 (N_7913,N_6391,N_6244);
nor U7914 (N_7914,N_7136,N_7034);
xor U7915 (N_7915,N_7080,N_6074);
or U7916 (N_7916,N_6088,N_6571);
xor U7917 (N_7917,N_6236,N_6134);
nor U7918 (N_7918,N_7102,N_7493);
nand U7919 (N_7919,N_6339,N_7437);
nand U7920 (N_7920,N_7474,N_7064);
and U7921 (N_7921,N_6361,N_7189);
xnor U7922 (N_7922,N_6158,N_6288);
nand U7923 (N_7923,N_7204,N_7104);
or U7924 (N_7924,N_6656,N_6113);
nor U7925 (N_7925,N_7151,N_6999);
and U7926 (N_7926,N_6993,N_7442);
nor U7927 (N_7927,N_6348,N_6588);
nand U7928 (N_7928,N_6786,N_7061);
nor U7929 (N_7929,N_6169,N_6465);
or U7930 (N_7930,N_6798,N_6002);
nand U7931 (N_7931,N_7351,N_6799);
or U7932 (N_7932,N_6918,N_7013);
or U7933 (N_7933,N_7292,N_7077);
or U7934 (N_7934,N_6979,N_6069);
nand U7935 (N_7935,N_6413,N_7346);
xnor U7936 (N_7936,N_6769,N_7125);
nand U7937 (N_7937,N_6782,N_6869);
xor U7938 (N_7938,N_6313,N_6845);
nor U7939 (N_7939,N_7065,N_7419);
and U7940 (N_7940,N_7047,N_6330);
and U7941 (N_7941,N_6997,N_6764);
and U7942 (N_7942,N_6263,N_7488);
nor U7943 (N_7943,N_6467,N_6108);
nand U7944 (N_7944,N_6662,N_6071);
and U7945 (N_7945,N_6834,N_6730);
or U7946 (N_7946,N_6333,N_7480);
or U7947 (N_7947,N_6030,N_7301);
nor U7948 (N_7948,N_6917,N_6770);
nand U7949 (N_7949,N_6970,N_6057);
and U7950 (N_7950,N_6636,N_6590);
nand U7951 (N_7951,N_7450,N_6036);
xnor U7952 (N_7952,N_6995,N_6632);
or U7953 (N_7953,N_7195,N_6954);
or U7954 (N_7954,N_6722,N_6553);
xor U7955 (N_7955,N_6922,N_6282);
nor U7956 (N_7956,N_6814,N_6357);
nor U7957 (N_7957,N_6951,N_6630);
and U7958 (N_7958,N_7398,N_6202);
and U7959 (N_7959,N_7322,N_7295);
or U7960 (N_7960,N_6068,N_7090);
and U7961 (N_7961,N_6340,N_6911);
nand U7962 (N_7962,N_6891,N_6405);
nor U7963 (N_7963,N_7415,N_6562);
and U7964 (N_7964,N_6087,N_6055);
and U7965 (N_7965,N_6414,N_6714);
and U7966 (N_7966,N_6053,N_6187);
nand U7967 (N_7967,N_6117,N_7200);
nand U7968 (N_7968,N_6144,N_6041);
or U7969 (N_7969,N_7468,N_6443);
or U7970 (N_7970,N_6360,N_7000);
and U7971 (N_7971,N_6797,N_6452);
nand U7972 (N_7972,N_7096,N_6006);
xor U7973 (N_7973,N_7342,N_6363);
and U7974 (N_7974,N_6175,N_6534);
nor U7975 (N_7975,N_7074,N_6412);
nand U7976 (N_7976,N_7242,N_6100);
nand U7977 (N_7977,N_7015,N_6941);
and U7978 (N_7978,N_7045,N_6196);
or U7979 (N_7979,N_6757,N_6514);
xnor U7980 (N_7980,N_6996,N_6824);
nor U7981 (N_7981,N_6379,N_6347);
nand U7982 (N_7982,N_7150,N_6112);
or U7983 (N_7983,N_7270,N_6215);
or U7984 (N_7984,N_7303,N_6589);
or U7985 (N_7985,N_6453,N_6736);
and U7986 (N_7986,N_6618,N_7444);
and U7987 (N_7987,N_6654,N_7484);
or U7988 (N_7988,N_7140,N_7476);
nand U7989 (N_7989,N_6111,N_7438);
and U7990 (N_7990,N_6530,N_6086);
nand U7991 (N_7991,N_6359,N_6417);
or U7992 (N_7992,N_6060,N_6054);
and U7993 (N_7993,N_6645,N_7423);
nor U7994 (N_7994,N_6569,N_6448);
or U7995 (N_7995,N_6258,N_6742);
nand U7996 (N_7996,N_7449,N_7374);
and U7997 (N_7997,N_7385,N_6699);
nor U7998 (N_7998,N_6533,N_6293);
nor U7999 (N_7999,N_6422,N_7217);
or U8000 (N_8000,N_7107,N_6925);
nor U8001 (N_8001,N_6062,N_7441);
xnor U8002 (N_8002,N_6114,N_7220);
and U8003 (N_8003,N_7274,N_6813);
or U8004 (N_8004,N_7343,N_6987);
nor U8005 (N_8005,N_7060,N_7066);
xor U8006 (N_8006,N_6865,N_6899);
or U8007 (N_8007,N_6565,N_6637);
and U8008 (N_8008,N_6919,N_6296);
or U8009 (N_8009,N_6584,N_7128);
or U8010 (N_8010,N_7209,N_6494);
xnor U8011 (N_8011,N_6886,N_6105);
or U8012 (N_8012,N_6305,N_7446);
or U8013 (N_8013,N_7286,N_7302);
and U8014 (N_8014,N_6429,N_6804);
nand U8015 (N_8015,N_6311,N_6378);
or U8016 (N_8016,N_6499,N_7384);
and U8017 (N_8017,N_6940,N_6727);
nor U8018 (N_8018,N_6482,N_6836);
nor U8019 (N_8019,N_6008,N_7025);
or U8020 (N_8020,N_7103,N_6929);
or U8021 (N_8021,N_6140,N_6840);
and U8022 (N_8022,N_7323,N_6596);
xor U8023 (N_8023,N_7144,N_6395);
nand U8024 (N_8024,N_6364,N_6811);
xnor U8025 (N_8025,N_6894,N_6484);
nor U8026 (N_8026,N_6191,N_6147);
or U8027 (N_8027,N_6788,N_7269);
or U8028 (N_8028,N_6199,N_7073);
nor U8029 (N_8029,N_6136,N_7024);
xnor U8030 (N_8030,N_6281,N_6243);
nand U8031 (N_8031,N_6207,N_6527);
nand U8032 (N_8032,N_7039,N_6273);
and U8033 (N_8033,N_7329,N_7057);
or U8034 (N_8034,N_6325,N_6745);
nand U8035 (N_8035,N_6271,N_7011);
nand U8036 (N_8036,N_7317,N_7349);
nand U8037 (N_8037,N_6949,N_7094);
and U8038 (N_8038,N_6197,N_6368);
nor U8039 (N_8039,N_6042,N_7161);
nand U8040 (N_8040,N_6517,N_6810);
or U8041 (N_8041,N_6992,N_6250);
nand U8042 (N_8042,N_7395,N_7012);
nand U8043 (N_8043,N_7429,N_7495);
or U8044 (N_8044,N_7233,N_6611);
xnor U8045 (N_8045,N_6208,N_6867);
nand U8046 (N_8046,N_6005,N_6262);
nand U8047 (N_8047,N_6239,N_6104);
or U8048 (N_8048,N_6220,N_6362);
and U8049 (N_8049,N_6885,N_7294);
nand U8050 (N_8050,N_7443,N_7071);
xor U8051 (N_8051,N_6698,N_7143);
or U8052 (N_8052,N_7262,N_6403);
and U8053 (N_8053,N_6397,N_7496);
xnor U8054 (N_8054,N_6307,N_7086);
nand U8055 (N_8055,N_6463,N_6860);
nand U8056 (N_8056,N_6511,N_6573);
xor U8057 (N_8057,N_7305,N_6953);
nor U8058 (N_8058,N_7145,N_6222);
and U8059 (N_8059,N_6655,N_6897);
or U8060 (N_8060,N_6023,N_6437);
nand U8061 (N_8061,N_7238,N_7259);
nand U8062 (N_8062,N_7149,N_6659);
nor U8063 (N_8063,N_6492,N_7487);
nand U8064 (N_8064,N_6981,N_6502);
nand U8065 (N_8065,N_6677,N_6634);
nor U8066 (N_8066,N_6697,N_7288);
nor U8067 (N_8067,N_7141,N_6278);
or U8068 (N_8068,N_6461,N_6027);
and U8069 (N_8069,N_7199,N_7308);
xor U8070 (N_8070,N_6327,N_6375);
or U8071 (N_8071,N_7164,N_7486);
and U8072 (N_8072,N_6316,N_6675);
or U8073 (N_8073,N_6302,N_6743);
nor U8074 (N_8074,N_7186,N_6740);
or U8075 (N_8075,N_6264,N_7030);
and U8076 (N_8076,N_7369,N_7359);
nor U8077 (N_8077,N_7304,N_7114);
nand U8078 (N_8078,N_7340,N_6560);
nor U8079 (N_8079,N_6715,N_6674);
nand U8080 (N_8080,N_7428,N_7027);
nor U8081 (N_8081,N_6162,N_7222);
and U8082 (N_8082,N_6734,N_7078);
nor U8083 (N_8083,N_6047,N_6572);
or U8084 (N_8084,N_6853,N_6728);
nor U8085 (N_8085,N_6767,N_6110);
nand U8086 (N_8086,N_6227,N_6440);
or U8087 (N_8087,N_7383,N_7127);
and U8088 (N_8088,N_6133,N_6424);
or U8089 (N_8089,N_6921,N_6358);
and U8090 (N_8090,N_6319,N_7226);
or U8091 (N_8091,N_7249,N_7210);
nor U8092 (N_8092,N_6615,N_6759);
nor U8093 (N_8093,N_6323,N_6966);
and U8094 (N_8094,N_7004,N_6238);
and U8095 (N_8095,N_6186,N_6084);
or U8096 (N_8096,N_6747,N_7083);
nand U8097 (N_8097,N_6503,N_6255);
nand U8098 (N_8098,N_6037,N_6908);
or U8099 (N_8099,N_6122,N_6098);
or U8100 (N_8100,N_6991,N_6178);
nor U8101 (N_8101,N_7465,N_6314);
nand U8102 (N_8102,N_6427,N_6138);
and U8103 (N_8103,N_6776,N_6056);
nor U8104 (N_8104,N_7489,N_6942);
nor U8105 (N_8105,N_6822,N_6665);
nor U8106 (N_8106,N_6835,N_7464);
nand U8107 (N_8107,N_7135,N_7434);
nand U8108 (N_8108,N_6989,N_6475);
or U8109 (N_8109,N_6717,N_6888);
nor U8110 (N_8110,N_7052,N_6432);
nor U8111 (N_8111,N_6274,N_7412);
or U8112 (N_8112,N_6033,N_6603);
xnor U8113 (N_8113,N_6635,N_6338);
or U8114 (N_8114,N_7089,N_7477);
or U8115 (N_8115,N_6052,N_6642);
nor U8116 (N_8116,N_6148,N_6773);
nand U8117 (N_8117,N_6123,N_7187);
nand U8118 (N_8118,N_7424,N_6524);
and U8119 (N_8119,N_6126,N_6212);
nor U8120 (N_8120,N_7360,N_6676);
nand U8121 (N_8121,N_6803,N_7354);
and U8122 (N_8122,N_6032,N_6164);
nor U8123 (N_8123,N_6651,N_6445);
or U8124 (N_8124,N_7368,N_7239);
nand U8125 (N_8125,N_6870,N_7048);
or U8126 (N_8126,N_6733,N_6044);
and U8127 (N_8127,N_6270,N_7332);
nand U8128 (N_8128,N_7212,N_7400);
and U8129 (N_8129,N_6240,N_6132);
xor U8130 (N_8130,N_6504,N_6758);
nor U8131 (N_8131,N_7055,N_7457);
nand U8132 (N_8132,N_7435,N_6291);
and U8133 (N_8133,N_7471,N_6561);
xnor U8134 (N_8134,N_7228,N_7033);
nand U8135 (N_8135,N_7422,N_6491);
and U8136 (N_8136,N_6121,N_6535);
nor U8137 (N_8137,N_7432,N_7014);
or U8138 (N_8138,N_6537,N_7120);
nand U8139 (N_8139,N_6719,N_6934);
and U8140 (N_8140,N_6003,N_7154);
and U8141 (N_8141,N_6831,N_7451);
nor U8142 (N_8142,N_7131,N_6490);
nor U8143 (N_8143,N_6176,N_6116);
or U8144 (N_8144,N_6696,N_6691);
nor U8145 (N_8145,N_7392,N_7123);
and U8146 (N_8146,N_6875,N_7293);
nor U8147 (N_8147,N_6658,N_7327);
or U8148 (N_8148,N_7116,N_6081);
or U8149 (N_8149,N_7409,N_6183);
and U8150 (N_8150,N_6004,N_7029);
nand U8151 (N_8151,N_7153,N_7396);
nand U8152 (N_8152,N_6269,N_7430);
and U8153 (N_8153,N_6434,N_6694);
xor U8154 (N_8154,N_7175,N_6476);
and U8155 (N_8155,N_6048,N_6883);
or U8156 (N_8156,N_7348,N_7225);
nand U8157 (N_8157,N_6930,N_7247);
or U8158 (N_8158,N_6219,N_7100);
or U8159 (N_8159,N_6034,N_6854);
and U8160 (N_8160,N_6352,N_6672);
nor U8161 (N_8161,N_7009,N_6292);
nand U8162 (N_8162,N_7205,N_7241);
or U8163 (N_8163,N_6859,N_6876);
or U8164 (N_8164,N_6015,N_7297);
or U8165 (N_8165,N_6369,N_6309);
and U8166 (N_8166,N_7256,N_7447);
and U8167 (N_8167,N_6371,N_6406);
nand U8168 (N_8168,N_7168,N_6863);
nand U8169 (N_8169,N_7485,N_6701);
or U8170 (N_8170,N_7098,N_6685);
and U8171 (N_8171,N_7092,N_6409);
or U8172 (N_8172,N_7184,N_6063);
xor U8173 (N_8173,N_6884,N_6545);
nand U8174 (N_8174,N_7335,N_6493);
xnor U8175 (N_8175,N_7146,N_6820);
nand U8176 (N_8176,N_6180,N_6387);
or U8177 (N_8177,N_6059,N_7216);
or U8178 (N_8178,N_7387,N_7405);
nor U8179 (N_8179,N_6708,N_6230);
or U8180 (N_8180,N_6485,N_6014);
nor U8181 (N_8181,N_6666,N_7201);
nor U8182 (N_8182,N_7379,N_6980);
nor U8183 (N_8183,N_6308,N_7063);
or U8184 (N_8184,N_7266,N_6025);
or U8185 (N_8185,N_6505,N_7382);
or U8186 (N_8186,N_7244,N_7499);
nand U8187 (N_8187,N_6793,N_6800);
or U8188 (N_8188,N_6442,N_7296);
and U8189 (N_8189,N_6952,N_6780);
nor U8190 (N_8190,N_6587,N_7155);
nor U8191 (N_8191,N_6724,N_6094);
nand U8192 (N_8192,N_6099,N_6683);
and U8193 (N_8193,N_6542,N_7007);
or U8194 (N_8194,N_6335,N_6246);
nand U8195 (N_8195,N_7481,N_6299);
xor U8196 (N_8196,N_7105,N_6737);
and U8197 (N_8197,N_7372,N_6512);
xnor U8198 (N_8198,N_6435,N_6231);
and U8199 (N_8199,N_6640,N_7193);
nand U8200 (N_8200,N_6154,N_6380);
xor U8201 (N_8201,N_7160,N_6253);
nand U8202 (N_8202,N_6617,N_6538);
nand U8203 (N_8203,N_6548,N_6889);
xnor U8204 (N_8204,N_7172,N_6506);
or U8205 (N_8205,N_7170,N_6754);
and U8206 (N_8206,N_6355,N_7005);
and U8207 (N_8207,N_6430,N_7169);
or U8208 (N_8208,N_6286,N_6515);
and U8209 (N_8209,N_6580,N_6923);
nand U8210 (N_8210,N_6205,N_6935);
and U8211 (N_8211,N_7459,N_6385);
xnor U8212 (N_8212,N_6947,N_6540);
nor U8213 (N_8213,N_6879,N_6622);
or U8214 (N_8214,N_7473,N_6247);
nor U8215 (N_8215,N_6639,N_7460);
or U8216 (N_8216,N_6095,N_6881);
nor U8217 (N_8217,N_7364,N_6438);
or U8218 (N_8218,N_6761,N_6858);
and U8219 (N_8219,N_6017,N_6983);
nor U8220 (N_8220,N_6218,N_7124);
nand U8221 (N_8221,N_7194,N_6458);
or U8222 (N_8222,N_6649,N_7121);
or U8223 (N_8223,N_6125,N_7250);
nor U8224 (N_8224,N_6209,N_7498);
and U8225 (N_8225,N_6488,N_7279);
or U8226 (N_8226,N_6926,N_6825);
or U8227 (N_8227,N_6495,N_6670);
xnor U8228 (N_8228,N_6460,N_6166);
and U8229 (N_8229,N_6578,N_6928);
nor U8230 (N_8230,N_6750,N_6620);
or U8231 (N_8231,N_6667,N_7407);
nand U8232 (N_8232,N_6910,N_6633);
xnor U8233 (N_8233,N_7054,N_6119);
or U8234 (N_8234,N_7035,N_6882);
nand U8235 (N_8235,N_6958,N_7001);
nor U8236 (N_8236,N_6161,N_6322);
nor U8237 (N_8237,N_7391,N_7417);
and U8238 (N_8238,N_7388,N_6795);
and U8239 (N_8239,N_6373,N_6586);
nor U8240 (N_8240,N_7115,N_7227);
or U8241 (N_8241,N_6805,N_7376);
nor U8242 (N_8242,N_6051,N_6937);
and U8243 (N_8243,N_6555,N_6823);
and U8244 (N_8244,N_7022,N_7208);
nand U8245 (N_8245,N_6990,N_7284);
or U8246 (N_8246,N_7361,N_6601);
or U8247 (N_8247,N_7345,N_6756);
or U8248 (N_8248,N_7076,N_6648);
or U8249 (N_8249,N_6167,N_6703);
and U8250 (N_8250,N_7480,N_6000);
nand U8251 (N_8251,N_6752,N_6838);
nor U8252 (N_8252,N_6451,N_7187);
or U8253 (N_8253,N_6733,N_7072);
and U8254 (N_8254,N_6732,N_7480);
and U8255 (N_8255,N_6305,N_6293);
nor U8256 (N_8256,N_6718,N_6810);
nor U8257 (N_8257,N_6510,N_6715);
xnor U8258 (N_8258,N_6139,N_6355);
and U8259 (N_8259,N_6787,N_6884);
and U8260 (N_8260,N_7451,N_7322);
nand U8261 (N_8261,N_7442,N_7461);
xor U8262 (N_8262,N_7138,N_7375);
nor U8263 (N_8263,N_7203,N_7351);
xor U8264 (N_8264,N_7296,N_6762);
and U8265 (N_8265,N_6080,N_7014);
nor U8266 (N_8266,N_6225,N_6143);
or U8267 (N_8267,N_6303,N_7093);
or U8268 (N_8268,N_6970,N_6459);
nand U8269 (N_8269,N_7290,N_7335);
xnor U8270 (N_8270,N_6057,N_7173);
xor U8271 (N_8271,N_6293,N_6188);
or U8272 (N_8272,N_6858,N_7299);
nand U8273 (N_8273,N_7299,N_7318);
xor U8274 (N_8274,N_6008,N_7432);
or U8275 (N_8275,N_7171,N_6365);
nor U8276 (N_8276,N_7473,N_6193);
nand U8277 (N_8277,N_6876,N_6896);
nor U8278 (N_8278,N_7207,N_6548);
and U8279 (N_8279,N_6503,N_6565);
nor U8280 (N_8280,N_6841,N_6658);
and U8281 (N_8281,N_7190,N_7498);
or U8282 (N_8282,N_7201,N_6095);
or U8283 (N_8283,N_6053,N_6548);
nor U8284 (N_8284,N_7357,N_6767);
nor U8285 (N_8285,N_6884,N_7080);
nor U8286 (N_8286,N_6690,N_7389);
nand U8287 (N_8287,N_6884,N_6494);
nor U8288 (N_8288,N_6037,N_6008);
and U8289 (N_8289,N_6948,N_6090);
nand U8290 (N_8290,N_7249,N_6151);
nor U8291 (N_8291,N_7281,N_6126);
or U8292 (N_8292,N_6412,N_6881);
or U8293 (N_8293,N_6765,N_6758);
and U8294 (N_8294,N_6690,N_6533);
nand U8295 (N_8295,N_6081,N_7053);
or U8296 (N_8296,N_6721,N_6022);
nand U8297 (N_8297,N_6544,N_7376);
and U8298 (N_8298,N_6260,N_6437);
or U8299 (N_8299,N_6724,N_7481);
nor U8300 (N_8300,N_6611,N_6037);
or U8301 (N_8301,N_7099,N_6284);
or U8302 (N_8302,N_7115,N_6333);
nor U8303 (N_8303,N_7231,N_7164);
nand U8304 (N_8304,N_6675,N_7142);
nand U8305 (N_8305,N_6091,N_7209);
and U8306 (N_8306,N_6336,N_6107);
and U8307 (N_8307,N_6920,N_6720);
and U8308 (N_8308,N_7165,N_6801);
nand U8309 (N_8309,N_7390,N_6125);
nand U8310 (N_8310,N_6849,N_6893);
xnor U8311 (N_8311,N_6091,N_6208);
xnor U8312 (N_8312,N_7279,N_7028);
nor U8313 (N_8313,N_7033,N_6615);
and U8314 (N_8314,N_6913,N_6270);
nor U8315 (N_8315,N_6333,N_7444);
and U8316 (N_8316,N_6751,N_6145);
nor U8317 (N_8317,N_6464,N_6072);
nand U8318 (N_8318,N_6754,N_6181);
and U8319 (N_8319,N_6014,N_6200);
nor U8320 (N_8320,N_6163,N_7346);
nor U8321 (N_8321,N_6545,N_6327);
or U8322 (N_8322,N_6245,N_6209);
nor U8323 (N_8323,N_6206,N_7321);
nand U8324 (N_8324,N_6449,N_7286);
and U8325 (N_8325,N_6835,N_7006);
nor U8326 (N_8326,N_6011,N_6635);
nand U8327 (N_8327,N_6767,N_6237);
and U8328 (N_8328,N_6543,N_7431);
nand U8329 (N_8329,N_7169,N_6284);
and U8330 (N_8330,N_6078,N_6367);
nand U8331 (N_8331,N_6073,N_6225);
and U8332 (N_8332,N_7330,N_7384);
nor U8333 (N_8333,N_6746,N_6344);
and U8334 (N_8334,N_7157,N_6192);
xor U8335 (N_8335,N_6813,N_6519);
nor U8336 (N_8336,N_6087,N_6168);
nor U8337 (N_8337,N_6799,N_6267);
nor U8338 (N_8338,N_7001,N_7105);
nand U8339 (N_8339,N_6021,N_7408);
and U8340 (N_8340,N_6086,N_7223);
nand U8341 (N_8341,N_6864,N_6519);
nand U8342 (N_8342,N_7474,N_6030);
nand U8343 (N_8343,N_6935,N_6101);
or U8344 (N_8344,N_6969,N_6106);
nor U8345 (N_8345,N_6184,N_7184);
nor U8346 (N_8346,N_6695,N_6068);
nor U8347 (N_8347,N_6121,N_7122);
or U8348 (N_8348,N_6555,N_6170);
and U8349 (N_8349,N_6380,N_7012);
nor U8350 (N_8350,N_7029,N_6624);
and U8351 (N_8351,N_7415,N_6969);
nor U8352 (N_8352,N_6086,N_6123);
and U8353 (N_8353,N_7214,N_6022);
nand U8354 (N_8354,N_6835,N_6713);
and U8355 (N_8355,N_6175,N_6174);
and U8356 (N_8356,N_7074,N_6886);
xor U8357 (N_8357,N_6029,N_6976);
or U8358 (N_8358,N_7188,N_6317);
nor U8359 (N_8359,N_6564,N_7313);
nand U8360 (N_8360,N_6576,N_6463);
nor U8361 (N_8361,N_6314,N_6810);
or U8362 (N_8362,N_6835,N_7115);
or U8363 (N_8363,N_6421,N_6660);
xnor U8364 (N_8364,N_6426,N_7166);
nor U8365 (N_8365,N_7240,N_6464);
or U8366 (N_8366,N_7208,N_6050);
nor U8367 (N_8367,N_7100,N_7470);
nand U8368 (N_8368,N_7384,N_6792);
nor U8369 (N_8369,N_7495,N_7236);
nand U8370 (N_8370,N_6657,N_7460);
or U8371 (N_8371,N_6177,N_6672);
or U8372 (N_8372,N_7171,N_6657);
nor U8373 (N_8373,N_7076,N_6735);
nand U8374 (N_8374,N_6580,N_7493);
nor U8375 (N_8375,N_6764,N_6039);
and U8376 (N_8376,N_7206,N_7471);
or U8377 (N_8377,N_7249,N_6687);
or U8378 (N_8378,N_6876,N_6922);
nand U8379 (N_8379,N_7483,N_7331);
and U8380 (N_8380,N_6760,N_6498);
and U8381 (N_8381,N_6992,N_6773);
or U8382 (N_8382,N_7469,N_7150);
nor U8383 (N_8383,N_7165,N_6156);
and U8384 (N_8384,N_6595,N_7378);
or U8385 (N_8385,N_6046,N_6401);
and U8386 (N_8386,N_6937,N_6049);
or U8387 (N_8387,N_7218,N_6251);
nor U8388 (N_8388,N_6984,N_7263);
nand U8389 (N_8389,N_7365,N_6885);
xor U8390 (N_8390,N_6314,N_6367);
nor U8391 (N_8391,N_7135,N_6856);
and U8392 (N_8392,N_6956,N_7191);
xor U8393 (N_8393,N_6905,N_6703);
or U8394 (N_8394,N_6023,N_7158);
nand U8395 (N_8395,N_6244,N_7150);
nor U8396 (N_8396,N_7483,N_6054);
xor U8397 (N_8397,N_6891,N_6314);
nand U8398 (N_8398,N_6492,N_6254);
nor U8399 (N_8399,N_6448,N_6492);
nand U8400 (N_8400,N_6326,N_6751);
nand U8401 (N_8401,N_6856,N_6056);
or U8402 (N_8402,N_6928,N_7016);
and U8403 (N_8403,N_7263,N_7256);
nor U8404 (N_8404,N_6380,N_6086);
or U8405 (N_8405,N_6382,N_7398);
xor U8406 (N_8406,N_7023,N_6329);
and U8407 (N_8407,N_7375,N_6037);
or U8408 (N_8408,N_6361,N_6126);
xnor U8409 (N_8409,N_7183,N_7184);
nand U8410 (N_8410,N_6694,N_6714);
and U8411 (N_8411,N_6760,N_6686);
or U8412 (N_8412,N_6737,N_7013);
nand U8413 (N_8413,N_6290,N_7249);
xor U8414 (N_8414,N_6193,N_7357);
xor U8415 (N_8415,N_6903,N_6804);
nand U8416 (N_8416,N_6916,N_6888);
nor U8417 (N_8417,N_6604,N_7216);
nor U8418 (N_8418,N_7377,N_6012);
nand U8419 (N_8419,N_6528,N_6306);
nand U8420 (N_8420,N_6250,N_7486);
xor U8421 (N_8421,N_6349,N_6940);
and U8422 (N_8422,N_6990,N_6736);
or U8423 (N_8423,N_6699,N_6129);
nand U8424 (N_8424,N_6040,N_6769);
and U8425 (N_8425,N_7178,N_6877);
and U8426 (N_8426,N_6576,N_6612);
nor U8427 (N_8427,N_7050,N_6322);
and U8428 (N_8428,N_6965,N_6369);
nor U8429 (N_8429,N_6267,N_7309);
or U8430 (N_8430,N_6270,N_6279);
nor U8431 (N_8431,N_6078,N_7072);
or U8432 (N_8432,N_6929,N_7334);
nor U8433 (N_8433,N_7122,N_7431);
nor U8434 (N_8434,N_6817,N_6268);
nor U8435 (N_8435,N_6140,N_6058);
or U8436 (N_8436,N_6031,N_6033);
nand U8437 (N_8437,N_6396,N_6086);
and U8438 (N_8438,N_6068,N_7277);
nor U8439 (N_8439,N_6362,N_6056);
xor U8440 (N_8440,N_6027,N_6031);
xnor U8441 (N_8441,N_6778,N_6004);
and U8442 (N_8442,N_7141,N_7076);
or U8443 (N_8443,N_7239,N_6420);
or U8444 (N_8444,N_6766,N_7388);
or U8445 (N_8445,N_7148,N_6788);
and U8446 (N_8446,N_6489,N_7222);
and U8447 (N_8447,N_7436,N_6464);
nor U8448 (N_8448,N_6719,N_6174);
xor U8449 (N_8449,N_6634,N_6254);
nor U8450 (N_8450,N_6590,N_6348);
and U8451 (N_8451,N_6222,N_7340);
or U8452 (N_8452,N_6506,N_6815);
nand U8453 (N_8453,N_7111,N_6131);
xnor U8454 (N_8454,N_7274,N_7435);
nor U8455 (N_8455,N_6590,N_7495);
or U8456 (N_8456,N_6367,N_7008);
nand U8457 (N_8457,N_6263,N_7083);
nor U8458 (N_8458,N_6782,N_7359);
nor U8459 (N_8459,N_6605,N_6653);
xor U8460 (N_8460,N_6068,N_6998);
nand U8461 (N_8461,N_6948,N_7338);
nand U8462 (N_8462,N_6789,N_7457);
nor U8463 (N_8463,N_6404,N_7184);
and U8464 (N_8464,N_6387,N_7330);
nor U8465 (N_8465,N_7397,N_6384);
and U8466 (N_8466,N_6483,N_7446);
nand U8467 (N_8467,N_6549,N_7276);
and U8468 (N_8468,N_6990,N_6391);
and U8469 (N_8469,N_6990,N_7236);
nand U8470 (N_8470,N_6066,N_6318);
or U8471 (N_8471,N_6250,N_6891);
or U8472 (N_8472,N_6258,N_7239);
and U8473 (N_8473,N_6642,N_6558);
nand U8474 (N_8474,N_6538,N_6674);
nor U8475 (N_8475,N_6368,N_6741);
or U8476 (N_8476,N_6280,N_6285);
or U8477 (N_8477,N_7124,N_6824);
nor U8478 (N_8478,N_6710,N_6919);
nand U8479 (N_8479,N_7279,N_6228);
nor U8480 (N_8480,N_6041,N_7422);
and U8481 (N_8481,N_6760,N_6428);
nor U8482 (N_8482,N_6825,N_6387);
and U8483 (N_8483,N_6608,N_6193);
or U8484 (N_8484,N_7430,N_7492);
nand U8485 (N_8485,N_6306,N_6868);
and U8486 (N_8486,N_7111,N_7048);
and U8487 (N_8487,N_7311,N_6161);
nor U8488 (N_8488,N_6601,N_6752);
nor U8489 (N_8489,N_6295,N_6571);
nand U8490 (N_8490,N_6626,N_7444);
nor U8491 (N_8491,N_6625,N_6904);
nand U8492 (N_8492,N_6540,N_7474);
nand U8493 (N_8493,N_6739,N_7415);
nand U8494 (N_8494,N_6702,N_7218);
and U8495 (N_8495,N_7444,N_6531);
nand U8496 (N_8496,N_6219,N_7129);
nor U8497 (N_8497,N_6085,N_7031);
nand U8498 (N_8498,N_6968,N_7376);
or U8499 (N_8499,N_6479,N_6087);
and U8500 (N_8500,N_6607,N_7067);
nand U8501 (N_8501,N_6387,N_7334);
and U8502 (N_8502,N_6087,N_7201);
or U8503 (N_8503,N_6343,N_7025);
or U8504 (N_8504,N_7129,N_7227);
or U8505 (N_8505,N_6580,N_6654);
or U8506 (N_8506,N_6549,N_7164);
and U8507 (N_8507,N_6339,N_7225);
or U8508 (N_8508,N_7266,N_6316);
nand U8509 (N_8509,N_7372,N_6876);
nand U8510 (N_8510,N_7241,N_6079);
and U8511 (N_8511,N_7120,N_6273);
nand U8512 (N_8512,N_6058,N_6763);
nor U8513 (N_8513,N_6736,N_7479);
nand U8514 (N_8514,N_6325,N_6758);
nor U8515 (N_8515,N_7437,N_7001);
or U8516 (N_8516,N_6693,N_6030);
or U8517 (N_8517,N_6630,N_6483);
xor U8518 (N_8518,N_7002,N_6943);
xnor U8519 (N_8519,N_6614,N_7482);
xnor U8520 (N_8520,N_7266,N_6291);
and U8521 (N_8521,N_7129,N_7115);
or U8522 (N_8522,N_6960,N_7291);
and U8523 (N_8523,N_6846,N_6138);
or U8524 (N_8524,N_7254,N_6498);
nand U8525 (N_8525,N_6694,N_7092);
xnor U8526 (N_8526,N_6133,N_6091);
xor U8527 (N_8527,N_6551,N_7306);
nand U8528 (N_8528,N_6306,N_6927);
xnor U8529 (N_8529,N_6679,N_7313);
nand U8530 (N_8530,N_7075,N_6321);
nor U8531 (N_8531,N_6312,N_7375);
xor U8532 (N_8532,N_6598,N_6241);
and U8533 (N_8533,N_6636,N_6492);
or U8534 (N_8534,N_6114,N_6292);
nand U8535 (N_8535,N_7018,N_6265);
and U8536 (N_8536,N_6407,N_7390);
nand U8537 (N_8537,N_7148,N_6189);
nand U8538 (N_8538,N_7313,N_6411);
or U8539 (N_8539,N_7200,N_6613);
xor U8540 (N_8540,N_6775,N_7020);
nand U8541 (N_8541,N_6979,N_7388);
and U8542 (N_8542,N_6980,N_6415);
and U8543 (N_8543,N_6034,N_7389);
and U8544 (N_8544,N_6439,N_7346);
or U8545 (N_8545,N_6967,N_6788);
and U8546 (N_8546,N_6486,N_7005);
xnor U8547 (N_8547,N_6044,N_6474);
or U8548 (N_8548,N_6685,N_6670);
or U8549 (N_8549,N_7417,N_6914);
and U8550 (N_8550,N_7305,N_6724);
xnor U8551 (N_8551,N_6573,N_6766);
nor U8552 (N_8552,N_6065,N_7035);
nand U8553 (N_8553,N_6696,N_7314);
nor U8554 (N_8554,N_7154,N_6367);
nor U8555 (N_8555,N_6654,N_7317);
nand U8556 (N_8556,N_6694,N_7412);
nor U8557 (N_8557,N_7033,N_7252);
nor U8558 (N_8558,N_6018,N_6117);
nor U8559 (N_8559,N_7342,N_6743);
and U8560 (N_8560,N_6067,N_6772);
and U8561 (N_8561,N_6094,N_7120);
nor U8562 (N_8562,N_6796,N_6806);
nor U8563 (N_8563,N_6262,N_7009);
nor U8564 (N_8564,N_6259,N_7378);
or U8565 (N_8565,N_7078,N_6749);
and U8566 (N_8566,N_6260,N_6269);
nand U8567 (N_8567,N_7055,N_7095);
or U8568 (N_8568,N_6281,N_7334);
or U8569 (N_8569,N_7116,N_6740);
nand U8570 (N_8570,N_7136,N_6731);
or U8571 (N_8571,N_6572,N_6917);
xor U8572 (N_8572,N_7476,N_6139);
nor U8573 (N_8573,N_6027,N_7279);
and U8574 (N_8574,N_7053,N_7246);
nand U8575 (N_8575,N_7228,N_6315);
or U8576 (N_8576,N_7001,N_6046);
or U8577 (N_8577,N_6566,N_6351);
xor U8578 (N_8578,N_7040,N_7107);
nor U8579 (N_8579,N_6736,N_6745);
nor U8580 (N_8580,N_6382,N_7256);
nand U8581 (N_8581,N_7025,N_7499);
or U8582 (N_8582,N_7027,N_6419);
xnor U8583 (N_8583,N_6079,N_7107);
and U8584 (N_8584,N_6480,N_7290);
xor U8585 (N_8585,N_6119,N_6683);
nand U8586 (N_8586,N_6309,N_6431);
nand U8587 (N_8587,N_6980,N_7094);
nor U8588 (N_8588,N_6149,N_6226);
nor U8589 (N_8589,N_7168,N_6492);
nor U8590 (N_8590,N_7127,N_6382);
nand U8591 (N_8591,N_6086,N_6217);
xnor U8592 (N_8592,N_6069,N_6304);
and U8593 (N_8593,N_6965,N_7173);
nand U8594 (N_8594,N_7106,N_7095);
nor U8595 (N_8595,N_6915,N_6189);
nand U8596 (N_8596,N_6952,N_6339);
or U8597 (N_8597,N_6116,N_6909);
nor U8598 (N_8598,N_6038,N_6026);
or U8599 (N_8599,N_7119,N_6532);
xor U8600 (N_8600,N_7148,N_7127);
and U8601 (N_8601,N_6465,N_7163);
nand U8602 (N_8602,N_7137,N_6281);
or U8603 (N_8603,N_6859,N_6806);
and U8604 (N_8604,N_6888,N_6541);
or U8605 (N_8605,N_7398,N_6043);
or U8606 (N_8606,N_6245,N_6923);
xor U8607 (N_8607,N_6233,N_6164);
xnor U8608 (N_8608,N_6913,N_7257);
nor U8609 (N_8609,N_7141,N_6396);
or U8610 (N_8610,N_6841,N_7472);
or U8611 (N_8611,N_6128,N_6943);
or U8612 (N_8612,N_6531,N_6897);
or U8613 (N_8613,N_6236,N_6373);
or U8614 (N_8614,N_6418,N_7207);
and U8615 (N_8615,N_6021,N_6689);
or U8616 (N_8616,N_7130,N_6955);
nand U8617 (N_8617,N_6101,N_7441);
xnor U8618 (N_8618,N_6978,N_6880);
or U8619 (N_8619,N_6076,N_7152);
nand U8620 (N_8620,N_6902,N_6813);
and U8621 (N_8621,N_7175,N_6253);
nor U8622 (N_8622,N_6366,N_7061);
nand U8623 (N_8623,N_6846,N_6069);
nor U8624 (N_8624,N_7348,N_6405);
and U8625 (N_8625,N_6036,N_6066);
nand U8626 (N_8626,N_6815,N_7283);
xor U8627 (N_8627,N_6083,N_6030);
nand U8628 (N_8628,N_7082,N_7450);
and U8629 (N_8629,N_6339,N_6302);
and U8630 (N_8630,N_6138,N_6710);
and U8631 (N_8631,N_6378,N_6886);
or U8632 (N_8632,N_7454,N_6444);
nand U8633 (N_8633,N_6663,N_6606);
nor U8634 (N_8634,N_7312,N_7130);
xnor U8635 (N_8635,N_6229,N_7283);
and U8636 (N_8636,N_6250,N_6833);
nor U8637 (N_8637,N_6192,N_6684);
nor U8638 (N_8638,N_7330,N_6848);
or U8639 (N_8639,N_7413,N_7280);
xnor U8640 (N_8640,N_6740,N_6713);
and U8641 (N_8641,N_6593,N_6425);
nand U8642 (N_8642,N_6554,N_6631);
and U8643 (N_8643,N_6491,N_7431);
nor U8644 (N_8644,N_7355,N_6906);
or U8645 (N_8645,N_6663,N_6653);
and U8646 (N_8646,N_7343,N_7388);
or U8647 (N_8647,N_7150,N_6559);
or U8648 (N_8648,N_6680,N_7106);
or U8649 (N_8649,N_7038,N_6824);
nor U8650 (N_8650,N_6434,N_6460);
nor U8651 (N_8651,N_6297,N_6783);
nor U8652 (N_8652,N_6411,N_6428);
nor U8653 (N_8653,N_6453,N_6086);
or U8654 (N_8654,N_6201,N_6239);
and U8655 (N_8655,N_6100,N_6894);
and U8656 (N_8656,N_7145,N_6762);
or U8657 (N_8657,N_6136,N_7042);
or U8658 (N_8658,N_7287,N_6890);
nand U8659 (N_8659,N_6188,N_6753);
nand U8660 (N_8660,N_7127,N_6496);
and U8661 (N_8661,N_6742,N_7237);
nor U8662 (N_8662,N_7139,N_7180);
or U8663 (N_8663,N_6072,N_6441);
or U8664 (N_8664,N_7020,N_7135);
or U8665 (N_8665,N_6211,N_6718);
and U8666 (N_8666,N_6725,N_6716);
nand U8667 (N_8667,N_7410,N_6506);
xnor U8668 (N_8668,N_6130,N_6906);
and U8669 (N_8669,N_6450,N_6107);
and U8670 (N_8670,N_6822,N_6132);
or U8671 (N_8671,N_6169,N_6003);
or U8672 (N_8672,N_6064,N_7310);
or U8673 (N_8673,N_7223,N_6281);
nor U8674 (N_8674,N_6325,N_7241);
and U8675 (N_8675,N_7410,N_7105);
nor U8676 (N_8676,N_6903,N_6516);
or U8677 (N_8677,N_6847,N_6204);
and U8678 (N_8678,N_6595,N_6369);
xor U8679 (N_8679,N_6516,N_6229);
xor U8680 (N_8680,N_7063,N_7157);
nor U8681 (N_8681,N_7422,N_6187);
nand U8682 (N_8682,N_6587,N_7030);
and U8683 (N_8683,N_6424,N_6529);
xnor U8684 (N_8684,N_6566,N_7420);
nor U8685 (N_8685,N_7310,N_6542);
and U8686 (N_8686,N_6976,N_6618);
xor U8687 (N_8687,N_6462,N_6322);
xnor U8688 (N_8688,N_7129,N_6702);
nand U8689 (N_8689,N_7231,N_6338);
nor U8690 (N_8690,N_6034,N_7406);
or U8691 (N_8691,N_6661,N_7371);
xor U8692 (N_8692,N_6167,N_7269);
or U8693 (N_8693,N_6960,N_6431);
xnor U8694 (N_8694,N_6895,N_6805);
nor U8695 (N_8695,N_6853,N_7214);
or U8696 (N_8696,N_7064,N_7250);
nor U8697 (N_8697,N_6060,N_6151);
xnor U8698 (N_8698,N_7384,N_7302);
nor U8699 (N_8699,N_7137,N_6241);
and U8700 (N_8700,N_6247,N_6864);
xor U8701 (N_8701,N_6034,N_6448);
nand U8702 (N_8702,N_6023,N_6529);
or U8703 (N_8703,N_7406,N_6138);
and U8704 (N_8704,N_6782,N_6245);
nor U8705 (N_8705,N_6120,N_6100);
nor U8706 (N_8706,N_6794,N_7491);
nand U8707 (N_8707,N_6108,N_6854);
nor U8708 (N_8708,N_7357,N_6396);
nor U8709 (N_8709,N_6813,N_6498);
and U8710 (N_8710,N_6568,N_6134);
nor U8711 (N_8711,N_6101,N_6933);
nor U8712 (N_8712,N_6303,N_7126);
or U8713 (N_8713,N_7184,N_7050);
or U8714 (N_8714,N_6630,N_6017);
nor U8715 (N_8715,N_7146,N_6761);
and U8716 (N_8716,N_6937,N_6838);
and U8717 (N_8717,N_6244,N_6701);
or U8718 (N_8718,N_6613,N_6580);
nor U8719 (N_8719,N_7013,N_6864);
nand U8720 (N_8720,N_6293,N_7473);
or U8721 (N_8721,N_7330,N_6940);
or U8722 (N_8722,N_6769,N_7123);
and U8723 (N_8723,N_6649,N_6774);
nand U8724 (N_8724,N_7103,N_6759);
nor U8725 (N_8725,N_6484,N_7360);
nor U8726 (N_8726,N_7109,N_6435);
xnor U8727 (N_8727,N_6583,N_6199);
and U8728 (N_8728,N_6243,N_6446);
or U8729 (N_8729,N_6533,N_7266);
nand U8730 (N_8730,N_6498,N_6764);
and U8731 (N_8731,N_6792,N_6804);
and U8732 (N_8732,N_6381,N_7170);
nor U8733 (N_8733,N_6552,N_7143);
or U8734 (N_8734,N_6725,N_6398);
xnor U8735 (N_8735,N_7199,N_6810);
and U8736 (N_8736,N_6300,N_6090);
and U8737 (N_8737,N_6984,N_6367);
nor U8738 (N_8738,N_6915,N_7048);
and U8739 (N_8739,N_6261,N_6341);
nor U8740 (N_8740,N_6839,N_6020);
nand U8741 (N_8741,N_6190,N_6999);
or U8742 (N_8742,N_6499,N_6766);
nand U8743 (N_8743,N_6811,N_6444);
nor U8744 (N_8744,N_6766,N_7072);
nor U8745 (N_8745,N_7142,N_6534);
and U8746 (N_8746,N_6610,N_7367);
nand U8747 (N_8747,N_7337,N_6600);
nand U8748 (N_8748,N_7369,N_7394);
nand U8749 (N_8749,N_7483,N_7137);
xnor U8750 (N_8750,N_7254,N_7454);
nand U8751 (N_8751,N_6375,N_6908);
nor U8752 (N_8752,N_7231,N_6470);
and U8753 (N_8753,N_6375,N_6459);
xnor U8754 (N_8754,N_6370,N_6081);
nand U8755 (N_8755,N_6133,N_6079);
or U8756 (N_8756,N_6424,N_6361);
and U8757 (N_8757,N_6576,N_6467);
nand U8758 (N_8758,N_7019,N_6428);
nor U8759 (N_8759,N_6346,N_6250);
nand U8760 (N_8760,N_6327,N_6337);
and U8761 (N_8761,N_6571,N_6981);
nand U8762 (N_8762,N_7121,N_7283);
and U8763 (N_8763,N_6877,N_6954);
nand U8764 (N_8764,N_6899,N_6188);
nor U8765 (N_8765,N_6346,N_7008);
nand U8766 (N_8766,N_7070,N_7011);
nand U8767 (N_8767,N_7194,N_6220);
nor U8768 (N_8768,N_7175,N_6931);
nand U8769 (N_8769,N_6146,N_6061);
or U8770 (N_8770,N_6984,N_7348);
nor U8771 (N_8771,N_7083,N_7333);
nand U8772 (N_8772,N_7102,N_6792);
or U8773 (N_8773,N_6679,N_6299);
nand U8774 (N_8774,N_6366,N_6796);
nand U8775 (N_8775,N_7342,N_6560);
nand U8776 (N_8776,N_7439,N_6484);
xnor U8777 (N_8777,N_6179,N_6398);
and U8778 (N_8778,N_6842,N_7255);
nand U8779 (N_8779,N_6390,N_6101);
nor U8780 (N_8780,N_6213,N_6473);
and U8781 (N_8781,N_7039,N_6342);
nor U8782 (N_8782,N_6350,N_7383);
nand U8783 (N_8783,N_6240,N_7193);
or U8784 (N_8784,N_6764,N_7046);
or U8785 (N_8785,N_6387,N_7025);
or U8786 (N_8786,N_7460,N_6327);
nand U8787 (N_8787,N_6578,N_7024);
nand U8788 (N_8788,N_6198,N_6352);
nor U8789 (N_8789,N_6426,N_6154);
and U8790 (N_8790,N_7056,N_7284);
and U8791 (N_8791,N_6796,N_6099);
nand U8792 (N_8792,N_6084,N_7347);
nand U8793 (N_8793,N_6261,N_6724);
nor U8794 (N_8794,N_6205,N_7420);
and U8795 (N_8795,N_6488,N_7338);
nand U8796 (N_8796,N_6076,N_6620);
or U8797 (N_8797,N_7338,N_6394);
nand U8798 (N_8798,N_6133,N_6924);
nor U8799 (N_8799,N_7043,N_7258);
nand U8800 (N_8800,N_6359,N_6480);
nand U8801 (N_8801,N_6641,N_7262);
or U8802 (N_8802,N_6260,N_6598);
nor U8803 (N_8803,N_6194,N_7180);
and U8804 (N_8804,N_6965,N_6753);
and U8805 (N_8805,N_6127,N_7255);
nor U8806 (N_8806,N_6031,N_7316);
nand U8807 (N_8807,N_7477,N_6689);
or U8808 (N_8808,N_6559,N_7168);
nand U8809 (N_8809,N_7089,N_6264);
and U8810 (N_8810,N_6206,N_6828);
nor U8811 (N_8811,N_6351,N_6895);
nor U8812 (N_8812,N_7057,N_6509);
nand U8813 (N_8813,N_6147,N_7389);
nand U8814 (N_8814,N_6717,N_6654);
or U8815 (N_8815,N_6109,N_6623);
nor U8816 (N_8816,N_6482,N_6813);
or U8817 (N_8817,N_7260,N_7012);
nand U8818 (N_8818,N_6174,N_6721);
nor U8819 (N_8819,N_6119,N_6502);
or U8820 (N_8820,N_6449,N_7193);
or U8821 (N_8821,N_6553,N_6497);
nand U8822 (N_8822,N_7402,N_6277);
nand U8823 (N_8823,N_6214,N_6386);
nor U8824 (N_8824,N_7286,N_7096);
and U8825 (N_8825,N_6110,N_6634);
and U8826 (N_8826,N_7454,N_6999);
and U8827 (N_8827,N_7443,N_7425);
xnor U8828 (N_8828,N_6453,N_7325);
nand U8829 (N_8829,N_6882,N_7180);
nand U8830 (N_8830,N_6827,N_7238);
nor U8831 (N_8831,N_6130,N_6564);
or U8832 (N_8832,N_7087,N_6134);
or U8833 (N_8833,N_7257,N_6501);
or U8834 (N_8834,N_6727,N_6501);
and U8835 (N_8835,N_6469,N_6115);
or U8836 (N_8836,N_6758,N_6211);
or U8837 (N_8837,N_7319,N_6666);
or U8838 (N_8838,N_6338,N_7237);
or U8839 (N_8839,N_6213,N_7006);
and U8840 (N_8840,N_7093,N_7314);
or U8841 (N_8841,N_6177,N_6879);
xor U8842 (N_8842,N_6549,N_6747);
and U8843 (N_8843,N_6968,N_6036);
nand U8844 (N_8844,N_6117,N_6751);
nand U8845 (N_8845,N_6649,N_6040);
and U8846 (N_8846,N_7010,N_7005);
and U8847 (N_8847,N_6619,N_6439);
nand U8848 (N_8848,N_6534,N_6676);
or U8849 (N_8849,N_6597,N_6486);
and U8850 (N_8850,N_7157,N_7094);
and U8851 (N_8851,N_6795,N_7055);
nand U8852 (N_8852,N_6278,N_6174);
nand U8853 (N_8853,N_6293,N_6676);
and U8854 (N_8854,N_6432,N_6766);
and U8855 (N_8855,N_7488,N_7083);
and U8856 (N_8856,N_6193,N_7409);
nor U8857 (N_8857,N_6992,N_7333);
nand U8858 (N_8858,N_7388,N_6364);
or U8859 (N_8859,N_6623,N_6710);
or U8860 (N_8860,N_6227,N_6535);
or U8861 (N_8861,N_7307,N_6049);
xnor U8862 (N_8862,N_7339,N_6190);
xor U8863 (N_8863,N_6491,N_6383);
or U8864 (N_8864,N_7441,N_6721);
nor U8865 (N_8865,N_6301,N_6238);
and U8866 (N_8866,N_7425,N_6784);
nand U8867 (N_8867,N_6449,N_6841);
or U8868 (N_8868,N_6272,N_7391);
or U8869 (N_8869,N_6895,N_6336);
nor U8870 (N_8870,N_6986,N_6517);
nand U8871 (N_8871,N_6820,N_6758);
or U8872 (N_8872,N_7460,N_6008);
nand U8873 (N_8873,N_7313,N_7350);
nand U8874 (N_8874,N_6196,N_7042);
nor U8875 (N_8875,N_7341,N_7351);
or U8876 (N_8876,N_6445,N_6846);
and U8877 (N_8877,N_6354,N_7117);
xnor U8878 (N_8878,N_6933,N_7159);
nor U8879 (N_8879,N_6663,N_6731);
or U8880 (N_8880,N_7104,N_6441);
nor U8881 (N_8881,N_6597,N_7174);
and U8882 (N_8882,N_6224,N_7137);
xnor U8883 (N_8883,N_7223,N_7322);
nand U8884 (N_8884,N_6774,N_6191);
nand U8885 (N_8885,N_6023,N_7175);
nand U8886 (N_8886,N_6923,N_7463);
and U8887 (N_8887,N_6880,N_6533);
and U8888 (N_8888,N_7066,N_7008);
nor U8889 (N_8889,N_6117,N_7064);
nor U8890 (N_8890,N_6463,N_7016);
or U8891 (N_8891,N_7450,N_6324);
nand U8892 (N_8892,N_6079,N_6551);
or U8893 (N_8893,N_6506,N_7214);
or U8894 (N_8894,N_6376,N_7145);
nor U8895 (N_8895,N_7256,N_6134);
xor U8896 (N_8896,N_6278,N_7459);
and U8897 (N_8897,N_6534,N_6828);
nand U8898 (N_8898,N_6979,N_6297);
nand U8899 (N_8899,N_6847,N_6604);
and U8900 (N_8900,N_7206,N_6514);
or U8901 (N_8901,N_7218,N_6340);
nand U8902 (N_8902,N_6196,N_6423);
and U8903 (N_8903,N_6567,N_6264);
nor U8904 (N_8904,N_7353,N_6677);
nor U8905 (N_8905,N_7207,N_6049);
and U8906 (N_8906,N_7353,N_7293);
nor U8907 (N_8907,N_7254,N_6915);
nand U8908 (N_8908,N_7005,N_6969);
nor U8909 (N_8909,N_7409,N_6360);
nand U8910 (N_8910,N_6441,N_6168);
xnor U8911 (N_8911,N_6906,N_7136);
nor U8912 (N_8912,N_7414,N_7292);
nor U8913 (N_8913,N_6424,N_6431);
nand U8914 (N_8914,N_7472,N_6431);
and U8915 (N_8915,N_6163,N_6639);
nand U8916 (N_8916,N_6989,N_6090);
or U8917 (N_8917,N_6301,N_7376);
nand U8918 (N_8918,N_7033,N_7498);
nor U8919 (N_8919,N_7234,N_7455);
nor U8920 (N_8920,N_6799,N_6180);
xnor U8921 (N_8921,N_6686,N_7147);
and U8922 (N_8922,N_6665,N_7276);
nor U8923 (N_8923,N_6205,N_6556);
nor U8924 (N_8924,N_7424,N_6689);
nor U8925 (N_8925,N_7003,N_6724);
xor U8926 (N_8926,N_7175,N_6519);
nor U8927 (N_8927,N_6191,N_6979);
nand U8928 (N_8928,N_6882,N_6365);
nand U8929 (N_8929,N_7363,N_6348);
and U8930 (N_8930,N_6059,N_6488);
nand U8931 (N_8931,N_7300,N_6033);
nand U8932 (N_8932,N_6792,N_7213);
or U8933 (N_8933,N_6705,N_7355);
nand U8934 (N_8934,N_7022,N_7178);
nand U8935 (N_8935,N_7276,N_6591);
or U8936 (N_8936,N_6329,N_7110);
nand U8937 (N_8937,N_7391,N_6787);
and U8938 (N_8938,N_6958,N_6937);
nand U8939 (N_8939,N_6826,N_6616);
nand U8940 (N_8940,N_6021,N_7336);
or U8941 (N_8941,N_6199,N_6492);
and U8942 (N_8942,N_7086,N_6562);
nor U8943 (N_8943,N_6832,N_7275);
nor U8944 (N_8944,N_6510,N_6333);
or U8945 (N_8945,N_6522,N_6811);
nor U8946 (N_8946,N_6219,N_7219);
and U8947 (N_8947,N_7134,N_7257);
nand U8948 (N_8948,N_7078,N_6086);
and U8949 (N_8949,N_6674,N_6503);
and U8950 (N_8950,N_7434,N_6798);
and U8951 (N_8951,N_6114,N_6712);
nand U8952 (N_8952,N_6393,N_6512);
and U8953 (N_8953,N_7348,N_6378);
or U8954 (N_8954,N_6102,N_7437);
or U8955 (N_8955,N_6411,N_7195);
and U8956 (N_8956,N_6024,N_6277);
or U8957 (N_8957,N_6172,N_6448);
nor U8958 (N_8958,N_6966,N_6217);
nand U8959 (N_8959,N_7439,N_6158);
nor U8960 (N_8960,N_6666,N_6670);
nand U8961 (N_8961,N_6311,N_6747);
or U8962 (N_8962,N_6238,N_6395);
or U8963 (N_8963,N_6602,N_6465);
or U8964 (N_8964,N_6206,N_7261);
nor U8965 (N_8965,N_7085,N_6951);
nor U8966 (N_8966,N_6188,N_6652);
or U8967 (N_8967,N_7104,N_6808);
nand U8968 (N_8968,N_7159,N_7094);
or U8969 (N_8969,N_7375,N_6627);
nand U8970 (N_8970,N_6630,N_6992);
or U8971 (N_8971,N_7228,N_7176);
nor U8972 (N_8972,N_6556,N_7429);
and U8973 (N_8973,N_6570,N_6974);
xor U8974 (N_8974,N_6145,N_7142);
nor U8975 (N_8975,N_6798,N_6440);
and U8976 (N_8976,N_6764,N_7345);
and U8977 (N_8977,N_6942,N_7135);
xor U8978 (N_8978,N_7258,N_7435);
nand U8979 (N_8979,N_6371,N_7027);
nand U8980 (N_8980,N_7349,N_6977);
nand U8981 (N_8981,N_6584,N_6268);
or U8982 (N_8982,N_7028,N_6406);
or U8983 (N_8983,N_6692,N_6834);
nand U8984 (N_8984,N_7267,N_7341);
or U8985 (N_8985,N_6251,N_6930);
nand U8986 (N_8986,N_6368,N_6291);
nand U8987 (N_8987,N_6242,N_7477);
nand U8988 (N_8988,N_7128,N_6129);
xor U8989 (N_8989,N_6307,N_6987);
nor U8990 (N_8990,N_6502,N_6674);
and U8991 (N_8991,N_6553,N_6672);
nor U8992 (N_8992,N_7111,N_7195);
and U8993 (N_8993,N_6728,N_6334);
nor U8994 (N_8994,N_7236,N_6195);
or U8995 (N_8995,N_6459,N_6622);
xor U8996 (N_8996,N_7075,N_7473);
and U8997 (N_8997,N_6553,N_6733);
and U8998 (N_8998,N_6354,N_6650);
nand U8999 (N_8999,N_7193,N_6946);
xor U9000 (N_9000,N_8420,N_8833);
nand U9001 (N_9001,N_7907,N_8057);
and U9002 (N_9002,N_7980,N_8434);
nor U9003 (N_9003,N_8291,N_7555);
xnor U9004 (N_9004,N_8148,N_8152);
nand U9005 (N_9005,N_8363,N_8820);
and U9006 (N_9006,N_7977,N_7634);
and U9007 (N_9007,N_8428,N_8711);
nor U9008 (N_9008,N_7516,N_7870);
nand U9009 (N_9009,N_8108,N_7881);
or U9010 (N_9010,N_8872,N_8464);
nand U9011 (N_9011,N_8981,N_7524);
or U9012 (N_9012,N_8260,N_8520);
nor U9013 (N_9013,N_7591,N_7791);
nand U9014 (N_9014,N_8048,N_8914);
and U9015 (N_9015,N_8760,N_8731);
nor U9016 (N_9016,N_8145,N_7878);
or U9017 (N_9017,N_8812,N_8065);
nand U9018 (N_9018,N_8450,N_8063);
or U9019 (N_9019,N_8021,N_7617);
and U9020 (N_9020,N_8446,N_8839);
or U9021 (N_9021,N_8422,N_8730);
nand U9022 (N_9022,N_8800,N_8697);
nand U9023 (N_9023,N_7646,N_7859);
or U9024 (N_9024,N_7974,N_8873);
nor U9025 (N_9025,N_8763,N_8512);
nor U9026 (N_9026,N_8311,N_8451);
nand U9027 (N_9027,N_8320,N_8902);
or U9028 (N_9028,N_7582,N_7904);
nor U9029 (N_9029,N_8782,N_7540);
nor U9030 (N_9030,N_8991,N_8777);
and U9031 (N_9031,N_8824,N_8398);
or U9032 (N_9032,N_7528,N_8035);
nand U9033 (N_9033,N_7626,N_7560);
nand U9034 (N_9034,N_8047,N_8941);
nor U9035 (N_9035,N_8208,N_8727);
and U9036 (N_9036,N_7811,N_8085);
or U9037 (N_9037,N_8556,N_7542);
xnor U9038 (N_9038,N_8948,N_8427);
or U9039 (N_9039,N_8429,N_8765);
nand U9040 (N_9040,N_8792,N_7586);
nand U9041 (N_9041,N_8261,N_7619);
nor U9042 (N_9042,N_7906,N_7843);
and U9043 (N_9043,N_7603,N_8983);
nand U9044 (N_9044,N_8814,N_8678);
and U9045 (N_9045,N_7761,N_8789);
nor U9046 (N_9046,N_8665,N_7537);
nand U9047 (N_9047,N_8139,N_8971);
nor U9048 (N_9048,N_8210,N_8615);
and U9049 (N_9049,N_8005,N_8608);
or U9050 (N_9050,N_8436,N_8146);
xor U9051 (N_9051,N_8797,N_7664);
nand U9052 (N_9052,N_8595,N_8612);
nand U9053 (N_9053,N_8070,N_8942);
nor U9054 (N_9054,N_8135,N_8857);
nor U9055 (N_9055,N_8172,N_8356);
nand U9056 (N_9056,N_8091,N_7650);
nand U9057 (N_9057,N_8387,N_8099);
nor U9058 (N_9058,N_8424,N_8967);
nand U9059 (N_9059,N_8488,N_8321);
and U9060 (N_9060,N_8028,N_8610);
nand U9061 (N_9061,N_7958,N_8822);
nand U9062 (N_9062,N_8324,N_8004);
nor U9063 (N_9063,N_8658,N_8372);
or U9064 (N_9064,N_8755,N_7564);
nor U9065 (N_9065,N_8354,N_7680);
nand U9066 (N_9066,N_8875,N_8032);
nand U9067 (N_9067,N_8623,N_7598);
or U9068 (N_9068,N_8346,N_8771);
nand U9069 (N_9069,N_8200,N_8044);
or U9070 (N_9070,N_7658,N_8323);
and U9071 (N_9071,N_7822,N_8911);
nand U9072 (N_9072,N_7709,N_8160);
nor U9073 (N_9073,N_7877,N_7563);
nor U9074 (N_9074,N_7995,N_8523);
and U9075 (N_9075,N_7826,N_8856);
or U9076 (N_9076,N_8564,N_8717);
or U9077 (N_9077,N_7857,N_7799);
xor U9078 (N_9078,N_8607,N_8114);
nand U9079 (N_9079,N_8205,N_8423);
xor U9080 (N_9080,N_8897,N_8600);
xor U9081 (N_9081,N_8851,N_7611);
xor U9082 (N_9082,N_7728,N_8507);
and U9083 (N_9083,N_7814,N_8453);
nand U9084 (N_9084,N_8509,N_8670);
nand U9085 (N_9085,N_7831,N_7796);
or U9086 (N_9086,N_7817,N_7840);
or U9087 (N_9087,N_8554,N_8953);
xor U9088 (N_9088,N_8435,N_8278);
xnor U9089 (N_9089,N_8449,N_7994);
and U9090 (N_9090,N_8233,N_8051);
nor U9091 (N_9091,N_8790,N_7723);
nand U9092 (N_9092,N_7970,N_8891);
nand U9093 (N_9093,N_8050,N_7635);
nand U9094 (N_9094,N_8632,N_8505);
nand U9095 (N_9095,N_7729,N_8781);
nor U9096 (N_9096,N_8475,N_8006);
or U9097 (N_9097,N_8325,N_8076);
xnor U9098 (N_9098,N_8293,N_8042);
nor U9099 (N_9099,N_8965,N_8784);
or U9100 (N_9100,N_8893,N_8534);
xnor U9101 (N_9101,N_7957,N_8726);
or U9102 (N_9102,N_8132,N_8212);
nand U9103 (N_9103,N_8750,N_8438);
nand U9104 (N_9104,N_8932,N_8654);
nor U9105 (N_9105,N_7866,N_8191);
nand U9106 (N_9106,N_8111,N_7942);
nand U9107 (N_9107,N_8740,N_8134);
xor U9108 (N_9108,N_8280,N_8604);
xor U9109 (N_9109,N_8588,N_8136);
and U9110 (N_9110,N_8131,N_7876);
nor U9111 (N_9111,N_8769,N_8343);
and U9112 (N_9112,N_8606,N_7851);
nor U9113 (N_9113,N_7987,N_7771);
nor U9114 (N_9114,N_7543,N_7825);
and U9115 (N_9115,N_8133,N_8796);
xnor U9116 (N_9116,N_8980,N_7684);
nand U9117 (N_9117,N_8213,N_7532);
and U9118 (N_9118,N_8360,N_7522);
or U9119 (N_9119,N_8494,N_7726);
or U9120 (N_9120,N_8227,N_8883);
nor U9121 (N_9121,N_7504,N_8926);
or U9122 (N_9122,N_8657,N_8586);
and U9123 (N_9123,N_7687,N_8409);
or U9124 (N_9124,N_7845,N_8445);
nor U9125 (N_9125,N_8403,N_8575);
or U9126 (N_9126,N_8371,N_7701);
and U9127 (N_9127,N_7861,N_7629);
nand U9128 (N_9128,N_8544,N_7609);
or U9129 (N_9129,N_8170,N_7679);
nor U9130 (N_9130,N_8164,N_8561);
and U9131 (N_9131,N_8693,N_7828);
nand U9132 (N_9132,N_8310,N_7571);
nor U9133 (N_9133,N_8976,N_8517);
nand U9134 (N_9134,N_8754,N_7640);
xnor U9135 (N_9135,N_8823,N_8269);
nor U9136 (N_9136,N_7940,N_8306);
nor U9137 (N_9137,N_7961,N_8444);
nand U9138 (N_9138,N_8794,N_8752);
and U9139 (N_9139,N_7715,N_8467);
or U9140 (N_9140,N_7765,N_7694);
and U9141 (N_9141,N_8033,N_8748);
and U9142 (N_9142,N_8110,N_8876);
and U9143 (N_9143,N_8843,N_8813);
nand U9144 (N_9144,N_7926,N_8944);
and U9145 (N_9145,N_7979,N_8892);
nand U9146 (N_9146,N_7931,N_7722);
nand U9147 (N_9147,N_8228,N_8602);
and U9148 (N_9148,N_8811,N_7772);
or U9149 (N_9149,N_8109,N_8737);
and U9150 (N_9150,N_7959,N_8799);
nand U9151 (N_9151,N_8120,N_8447);
and U9152 (N_9152,N_8836,N_7557);
or U9153 (N_9153,N_8027,N_8954);
xnor U9154 (N_9154,N_7782,N_8698);
and U9155 (N_9155,N_7523,N_8550);
nand U9156 (N_9156,N_8835,N_8441);
nor U9157 (N_9157,N_8772,N_8783);
and U9158 (N_9158,N_8008,N_8204);
and U9159 (N_9159,N_7850,N_8312);
and U9160 (N_9160,N_8171,N_7963);
and U9161 (N_9161,N_8583,N_7601);
or U9162 (N_9162,N_8142,N_8990);
and U9163 (N_9163,N_8405,N_8266);
and U9164 (N_9164,N_8530,N_7784);
nor U9165 (N_9165,N_7686,N_8045);
nor U9166 (N_9166,N_8055,N_7879);
and U9167 (N_9167,N_8504,N_7508);
and U9168 (N_9168,N_7746,N_8985);
nand U9169 (N_9169,N_8557,N_8679);
nor U9170 (N_9170,N_7880,N_8117);
or U9171 (N_9171,N_8770,N_7946);
and U9172 (N_9172,N_8921,N_8952);
xor U9173 (N_9173,N_8459,N_7518);
nand U9174 (N_9174,N_7808,N_8605);
xnor U9175 (N_9175,N_7804,N_8758);
xor U9176 (N_9176,N_8974,N_7887);
or U9177 (N_9177,N_7649,N_8179);
nand U9178 (N_9178,N_7741,N_8161);
nand U9179 (N_9179,N_8849,N_8756);
xnor U9180 (N_9180,N_7743,N_8244);
nand U9181 (N_9181,N_8531,N_7633);
nor U9182 (N_9182,N_7570,N_7777);
xnor U9183 (N_9183,N_8068,N_8469);
nand U9184 (N_9184,N_8270,N_8125);
or U9185 (N_9185,N_8041,N_8949);
or U9186 (N_9186,N_8098,N_8889);
and U9187 (N_9187,N_8964,N_8181);
or U9188 (N_9188,N_7872,N_8997);
nor U9189 (N_9189,N_8359,N_8620);
nand U9190 (N_9190,N_8089,N_7645);
or U9191 (N_9191,N_8102,N_8318);
nor U9192 (N_9192,N_7832,N_8513);
xor U9193 (N_9193,N_7602,N_8924);
and U9194 (N_9194,N_8274,N_8355);
or U9195 (N_9195,N_7975,N_7699);
and U9196 (N_9196,N_8712,N_8439);
nor U9197 (N_9197,N_8425,N_7769);
or U9198 (N_9198,N_8598,N_7574);
nor U9199 (N_9199,N_8353,N_7618);
nor U9200 (N_9200,N_7875,N_8844);
nor U9201 (N_9201,N_8576,N_7747);
nor U9202 (N_9202,N_7507,N_8681);
and U9203 (N_9203,N_8452,N_8518);
and U9204 (N_9204,N_8118,N_7717);
nand U9205 (N_9205,N_7930,N_7721);
and U9206 (N_9206,N_7889,N_7731);
nand U9207 (N_9207,N_7853,N_7565);
or U9208 (N_9208,N_8945,N_8675);
and U9209 (N_9209,N_7550,N_7541);
nor U9210 (N_9210,N_7984,N_7689);
nor U9211 (N_9211,N_8202,N_8484);
nor U9212 (N_9212,N_8336,N_7501);
nand U9213 (N_9213,N_7954,N_7763);
or U9214 (N_9214,N_8417,N_7939);
or U9215 (N_9215,N_8018,N_7670);
nand U9216 (N_9216,N_7801,N_8918);
or U9217 (N_9217,N_8448,N_7526);
nor U9218 (N_9218,N_8762,N_7732);
and U9219 (N_9219,N_8219,N_7667);
nand U9220 (N_9220,N_8377,N_8947);
or U9221 (N_9221,N_8471,N_7923);
nor U9222 (N_9222,N_8487,N_8618);
or U9223 (N_9223,N_8502,N_7632);
nor U9224 (N_9224,N_7669,N_8548);
xnor U9225 (N_9225,N_8049,N_7727);
nor U9226 (N_9226,N_8500,N_8128);
and U9227 (N_9227,N_8516,N_7512);
nor U9228 (N_9228,N_8072,N_8616);
or U9229 (N_9229,N_8286,N_7638);
or U9230 (N_9230,N_8011,N_7647);
nor U9231 (N_9231,N_7599,N_7860);
and U9232 (N_9232,N_8305,N_7554);
nand U9233 (N_9233,N_8759,N_7585);
and U9234 (N_9234,N_7841,N_8587);
nor U9235 (N_9235,N_8097,N_8087);
and U9236 (N_9236,N_8268,N_7606);
xor U9237 (N_9237,N_7558,N_8749);
or U9238 (N_9238,N_8719,N_7553);
nand U9239 (N_9239,N_7533,N_7909);
nor U9240 (N_9240,N_8014,N_8903);
or U9241 (N_9241,N_8309,N_7833);
and U9242 (N_9242,N_8388,N_8455);
or U9243 (N_9243,N_8662,N_8023);
xor U9244 (N_9244,N_8669,N_8722);
or U9245 (N_9245,N_7815,N_7973);
or U9246 (N_9246,N_8369,N_7648);
or U9247 (N_9247,N_8300,N_8601);
or U9248 (N_9248,N_8061,N_8144);
nand U9249 (N_9249,N_8106,N_7756);
nand U9250 (N_9250,N_8351,N_8887);
nand U9251 (N_9251,N_8637,N_7932);
and U9252 (N_9252,N_7884,N_7983);
nor U9253 (N_9253,N_8768,N_8565);
and U9254 (N_9254,N_7624,N_7823);
and U9255 (N_9255,N_8870,N_8721);
nand U9256 (N_9256,N_7581,N_8514);
or U9257 (N_9257,N_8700,N_7636);
nand U9258 (N_9258,N_8495,N_8246);
nor U9259 (N_9259,N_8252,N_7759);
xnor U9260 (N_9260,N_8592,N_8303);
nand U9261 (N_9261,N_8767,N_7625);
or U9262 (N_9262,N_7608,N_8243);
or U9263 (N_9263,N_7678,N_7613);
or U9264 (N_9264,N_7621,N_7999);
and U9265 (N_9265,N_8705,N_8378);
and U9266 (N_9266,N_7894,N_7842);
nor U9267 (N_9267,N_8928,N_7754);
and U9268 (N_9268,N_8101,N_8478);
or U9269 (N_9269,N_7534,N_8793);
xor U9270 (N_9270,N_7682,N_7527);
nand U9271 (N_9271,N_7837,N_7775);
and U9272 (N_9272,N_8828,N_8643);
nand U9273 (N_9273,N_8521,N_8651);
and U9274 (N_9274,N_8473,N_8358);
nand U9275 (N_9275,N_7673,N_8593);
nand U9276 (N_9276,N_8543,N_8066);
nand U9277 (N_9277,N_8294,N_7762);
nand U9278 (N_9278,N_8809,N_8374);
or U9279 (N_9279,N_8326,N_8810);
nor U9280 (N_9280,N_8163,N_8655);
or U9281 (N_9281,N_8166,N_8482);
nand U9282 (N_9282,N_8264,N_8284);
nand U9283 (N_9283,N_7949,N_7951);
nand U9284 (N_9284,N_8255,N_8638);
nand U9285 (N_9285,N_7720,N_7869);
nand U9286 (N_9286,N_8344,N_8054);
and U9287 (N_9287,N_7675,N_8385);
nor U9288 (N_9288,N_8720,N_8614);
or U9289 (N_9289,N_8939,N_7651);
nand U9290 (N_9290,N_7929,N_7862);
and U9291 (N_9291,N_7978,N_8716);
nor U9292 (N_9292,N_7655,N_8533);
and U9293 (N_9293,N_8150,N_7768);
nor U9294 (N_9294,N_8331,N_8126);
nand U9295 (N_9295,N_7604,N_7748);
xor U9296 (N_9296,N_7665,N_8515);
nand U9297 (N_9297,N_7852,N_7992);
nand U9298 (N_9298,N_7776,N_7578);
or U9299 (N_9299,N_7674,N_7924);
and U9300 (N_9300,N_8585,N_8297);
and U9301 (N_9301,N_7685,N_8682);
and U9302 (N_9302,N_7816,N_8639);
and U9303 (N_9303,N_8250,N_8563);
and U9304 (N_9304,N_7637,N_7809);
nand U9305 (N_9305,N_8242,N_8538);
nor U9306 (N_9306,N_8915,N_7751);
and U9307 (N_9307,N_8400,N_8677);
nor U9308 (N_9308,N_8917,N_7916);
or U9309 (N_9309,N_8113,N_7736);
nor U9310 (N_9310,N_8989,N_8203);
nand U9311 (N_9311,N_7967,N_8966);
and U9312 (N_9312,N_7780,N_8370);
or U9313 (N_9313,N_8725,N_8577);
xor U9314 (N_9314,N_8282,N_7838);
nand U9315 (N_9315,N_8062,N_8871);
nand U9316 (N_9316,N_8979,N_8619);
or U9317 (N_9317,N_7821,N_8993);
xnor U9318 (N_9318,N_8649,N_8265);
and U9319 (N_9319,N_8015,N_8982);
nand U9320 (N_9320,N_8798,N_8874);
or U9321 (N_9321,N_7500,N_8570);
and U9322 (N_9322,N_8086,N_7506);
and U9323 (N_9323,N_8396,N_8978);
nand U9324 (N_9324,N_8194,N_8723);
nor U9325 (N_9325,N_8256,N_7883);
nand U9326 (N_9326,N_8753,N_8036);
and U9327 (N_9327,N_7901,N_8234);
xnor U9328 (N_9328,N_8078,N_8847);
or U9329 (N_9329,N_8248,N_8263);
or U9330 (N_9330,N_8931,N_8082);
xor U9331 (N_9331,N_7536,N_7971);
and U9332 (N_9332,N_8165,N_7614);
and U9333 (N_9333,N_8462,N_7918);
or U9334 (N_9334,N_8906,N_7935);
or U9335 (N_9335,N_8640,N_8861);
nor U9336 (N_9336,N_8850,N_8551);
or U9337 (N_9337,N_8216,N_7538);
or U9338 (N_9338,N_8186,N_8776);
xnor U9339 (N_9339,N_8338,N_8877);
and U9340 (N_9340,N_8271,N_7797);
and U9341 (N_9341,N_8671,N_7903);
or U9342 (N_9342,N_7594,N_8384);
xor U9343 (N_9343,N_7631,N_7738);
nor U9344 (N_9344,N_7740,N_7810);
nand U9345 (N_9345,N_7713,N_8345);
nand U9346 (N_9346,N_8333,N_7703);
nand U9347 (N_9347,N_8829,N_8339);
and U9348 (N_9348,N_7937,N_8830);
and U9349 (N_9349,N_7596,N_8925);
nand U9350 (N_9350,N_8560,N_7610);
and U9351 (N_9351,N_8819,N_7583);
and U9352 (N_9352,N_8667,N_8237);
and U9353 (N_9353,N_8687,N_7864);
or U9354 (N_9354,N_7690,N_7734);
nand U9355 (N_9355,N_8340,N_8408);
and U9356 (N_9356,N_7915,N_8691);
or U9357 (N_9357,N_8149,N_7829);
nand U9358 (N_9358,N_7868,N_7724);
or U9359 (N_9359,N_7927,N_8259);
nor U9360 (N_9360,N_8209,N_8886);
nand U9361 (N_9361,N_8898,N_7998);
or U9362 (N_9362,N_8996,N_7652);
and U9363 (N_9363,N_8977,N_8157);
nor U9364 (N_9364,N_8295,N_7639);
or U9365 (N_9365,N_8332,N_7745);
or U9366 (N_9366,N_8580,N_8366);
or U9367 (N_9367,N_8104,N_7630);
nor U9368 (N_9368,N_7752,N_8442);
nand U9369 (N_9369,N_7529,N_8189);
nor U9370 (N_9370,N_8553,N_8454);
nand U9371 (N_9371,N_8650,N_8696);
and U9372 (N_9372,N_7579,N_8831);
nand U9373 (N_9373,N_8416,N_7891);
or U9374 (N_9374,N_8973,N_7712);
nand U9375 (N_9375,N_8406,N_7794);
xor U9376 (N_9376,N_8328,N_8468);
nand U9377 (N_9377,N_8426,N_7849);
or U9378 (N_9378,N_8421,N_7573);
or U9379 (N_9379,N_7600,N_7535);
nor U9380 (N_9380,N_8483,N_8497);
nand U9381 (N_9381,N_7502,N_8415);
or U9382 (N_9382,N_7695,N_8373);
nand U9383 (N_9383,N_8221,N_7917);
nor U9384 (N_9384,N_8704,N_8573);
xor U9385 (N_9385,N_8927,N_8167);
and U9386 (N_9386,N_8742,N_7662);
or U9387 (N_9387,N_8815,N_8433);
nand U9388 (N_9388,N_7642,N_7750);
nand U9389 (N_9389,N_8555,N_7530);
or U9390 (N_9390,N_7716,N_8791);
nand U9391 (N_9391,N_8357,N_8007);
or U9392 (N_9392,N_8672,N_7774);
and U9393 (N_9393,N_7925,N_8838);
xor U9394 (N_9394,N_7806,N_7749);
nand U9395 (N_9395,N_8214,N_8020);
nand U9396 (N_9396,N_7654,N_8489);
nand U9397 (N_9397,N_8506,N_8786);
nor U9398 (N_9398,N_7575,N_7990);
nor U9399 (N_9399,N_7911,N_7943);
nor U9400 (N_9400,N_8536,N_8192);
nand U9401 (N_9401,N_8361,N_8196);
nand U9402 (N_9402,N_7584,N_8147);
nand U9403 (N_9403,N_8298,N_7789);
nor U9404 (N_9404,N_7962,N_7834);
and U9405 (N_9405,N_8472,N_7547);
and U9406 (N_9406,N_8071,N_8702);
nor U9407 (N_9407,N_8825,N_8081);
and U9408 (N_9408,N_8582,N_8735);
and U9409 (N_9409,N_8100,N_8391);
nor U9410 (N_9410,N_8183,N_8714);
nand U9411 (N_9411,N_7525,N_8253);
nor U9412 (N_9412,N_8951,N_8092);
nand U9413 (N_9413,N_7548,N_7913);
nand U9414 (N_9414,N_7562,N_8404);
or U9415 (N_9415,N_8524,N_7733);
nor U9416 (N_9416,N_8056,N_7739);
nor U9417 (N_9417,N_7770,N_8955);
nor U9418 (N_9418,N_8162,N_7813);
or U9419 (N_9419,N_7890,N_8012);
nand U9420 (N_9420,N_7661,N_8962);
xnor U9421 (N_9421,N_8626,N_7793);
nor U9422 (N_9422,N_8067,N_8666);
or U9423 (N_9423,N_7790,N_8302);
or U9424 (N_9424,N_8413,N_7902);
nor U9425 (N_9425,N_8112,N_8090);
nand U9426 (N_9426,N_7580,N_7539);
nor U9427 (N_9427,N_8477,N_7844);
or U9428 (N_9428,N_8019,N_8412);
nor U9429 (N_9429,N_8910,N_8362);
nor U9430 (N_9430,N_8633,N_8493);
and U9431 (N_9431,N_8460,N_7965);
and U9432 (N_9432,N_8597,N_8900);
and U9433 (N_9433,N_8862,N_7892);
and U9434 (N_9434,N_8868,N_8349);
or U9435 (N_9435,N_8584,N_8299);
nor U9436 (N_9436,N_8708,N_8093);
nor U9437 (N_9437,N_7641,N_7921);
or U9438 (N_9438,N_7628,N_7515);
or U9439 (N_9439,N_8817,N_7824);
xnor U9440 (N_9440,N_7802,N_8046);
xnor U9441 (N_9441,N_7855,N_8074);
nand U9442 (N_9442,N_8549,N_8865);
and U9443 (N_9443,N_8491,N_7786);
and U9444 (N_9444,N_7783,N_7693);
or U9445 (N_9445,N_8138,N_8217);
nor U9446 (N_9446,N_8443,N_8578);
or U9447 (N_9447,N_8929,N_7947);
nor U9448 (N_9448,N_7672,N_8909);
and U9449 (N_9449,N_7663,N_8364);
or U9450 (N_9450,N_8958,N_8970);
and U9451 (N_9451,N_8972,N_8571);
or U9452 (N_9452,N_8375,N_8218);
nor U9453 (N_9453,N_7505,N_8201);
nand U9454 (N_9454,N_8207,N_8899);
or U9455 (N_9455,N_8279,N_8552);
nor U9456 (N_9456,N_8342,N_8567);
nor U9457 (N_9457,N_7950,N_7589);
and U9458 (N_9458,N_7847,N_8137);
and U9459 (N_9459,N_7800,N_8936);
nand U9460 (N_9460,N_8775,N_7960);
or U9461 (N_9461,N_7520,N_7659);
or U9462 (N_9462,N_7968,N_8431);
and U9463 (N_9463,N_8198,N_7854);
or U9464 (N_9464,N_8635,N_7807);
nor U9465 (N_9465,N_8852,N_8854);
and U9466 (N_9466,N_8394,N_8251);
or U9467 (N_9467,N_7873,N_8129);
and U9468 (N_9468,N_8465,N_8395);
nor U9469 (N_9469,N_8528,N_8627);
nand U9470 (N_9470,N_8766,N_8778);
nor U9471 (N_9471,N_7615,N_8846);
xor U9472 (N_9472,N_8069,N_8804);
and U9473 (N_9473,N_8743,N_8151);
nand U9474 (N_9474,N_8629,N_8540);
and U9475 (N_9475,N_8119,N_8330);
nand U9476 (N_9476,N_8457,N_8880);
nor U9477 (N_9477,N_7511,N_8154);
nor U9478 (N_9478,N_8501,N_8946);
nor U9479 (N_9479,N_8631,N_8624);
nor U9480 (N_9480,N_8296,N_8511);
nor U9481 (N_9481,N_7757,N_7556);
nand U9482 (N_9482,N_8231,N_8277);
or U9483 (N_9483,N_8289,N_7737);
nand U9484 (N_9484,N_8187,N_7900);
nor U9485 (N_9485,N_8940,N_7908);
or U9486 (N_9486,N_7773,N_8001);
nor U9487 (N_9487,N_7976,N_7711);
nand U9488 (N_9488,N_7944,N_8695);
nand U9489 (N_9489,N_8199,N_8002);
nand U9490 (N_9490,N_8881,N_7592);
nand U9491 (N_9491,N_7934,N_8747);
and U9492 (N_9492,N_8116,N_8184);
nor U9493 (N_9493,N_7702,N_7576);
and U9494 (N_9494,N_8519,N_7744);
nand U9495 (N_9495,N_8079,N_7595);
nand U9496 (N_9496,N_8175,N_8896);
or U9497 (N_9497,N_8827,N_7788);
or U9498 (N_9498,N_7572,N_8692);
and U9499 (N_9499,N_8807,N_8922);
nor U9500 (N_9500,N_8636,N_7865);
nand U9501 (N_9501,N_7830,N_8984);
nand U9502 (N_9502,N_8058,N_8392);
nor U9503 (N_9503,N_8879,N_8840);
nor U9504 (N_9504,N_8821,N_8016);
or U9505 (N_9505,N_7544,N_8314);
and U9506 (N_9506,N_8864,N_8647);
nor U9507 (N_9507,N_8476,N_7919);
nand U9508 (N_9508,N_8741,N_8975);
or U9509 (N_9509,N_8037,N_8327);
nor U9510 (N_9510,N_8569,N_8913);
nor U9511 (N_9511,N_8481,N_7820);
nor U9512 (N_9512,N_7714,N_8890);
xor U9513 (N_9513,N_8525,N_7707);
nand U9514 (N_9514,N_8030,N_8337);
xor U9515 (N_9515,N_7710,N_8188);
xnor U9516 (N_9516,N_8499,N_8155);
and U9517 (N_9517,N_8998,N_7945);
nor U9518 (N_9518,N_7899,N_7938);
or U9519 (N_9519,N_8867,N_7514);
nand U9520 (N_9520,N_8628,N_8229);
nand U9521 (N_9521,N_8130,N_8287);
or U9522 (N_9522,N_7566,N_8590);
or U9523 (N_9523,N_8646,N_8664);
and U9524 (N_9524,N_7835,N_7991);
or U9525 (N_9525,N_8316,N_8699);
nor U9526 (N_9526,N_8223,N_8096);
and U9527 (N_9527,N_8458,N_8961);
nor U9528 (N_9528,N_8818,N_8034);
nor U9529 (N_9529,N_8053,N_8674);
nor U9530 (N_9530,N_8845,N_7779);
nand U9531 (N_9531,N_8994,N_8774);
nor U9532 (N_9532,N_7567,N_8283);
nand U9533 (N_9533,N_7510,N_8292);
or U9534 (N_9534,N_7753,N_8411);
nor U9535 (N_9535,N_8919,N_8498);
and U9536 (N_9536,N_8103,N_7792);
and U9537 (N_9537,N_8661,N_8226);
nor U9538 (N_9538,N_8381,N_8878);
nor U9539 (N_9539,N_8934,N_8432);
nand U9540 (N_9540,N_8235,N_7607);
nand U9541 (N_9541,N_8841,N_8176);
nor U9542 (N_9542,N_7988,N_8043);
xnor U9543 (N_9543,N_8414,N_7982);
nor U9544 (N_9544,N_8609,N_8779);
or U9545 (N_9545,N_8140,N_7597);
nand U9546 (N_9546,N_8480,N_8938);
or U9547 (N_9547,N_7692,N_8652);
and U9548 (N_9548,N_7910,N_8684);
and U9549 (N_9549,N_8059,N_8676);
nand U9550 (N_9550,N_8322,N_7513);
xor U9551 (N_9551,N_7708,N_8738);
or U9552 (N_9552,N_8668,N_8795);
and U9553 (N_9553,N_7969,N_8347);
nor U9554 (N_9554,N_8220,N_8245);
nor U9555 (N_9555,N_7781,N_8503);
nor U9556 (N_9556,N_8622,N_8115);
nor U9557 (N_9557,N_7819,N_8240);
xnor U9558 (N_9558,N_7922,N_8574);
nor U9559 (N_9559,N_8143,N_8905);
and U9560 (N_9560,N_8174,N_8785);
and U9561 (N_9561,N_8642,N_8159);
and U9562 (N_9562,N_8156,N_8437);
nor U9563 (N_9563,N_8808,N_8526);
or U9564 (N_9564,N_8273,N_7798);
or U9565 (N_9565,N_7920,N_8386);
nor U9566 (N_9566,N_8496,N_8379);
or U9567 (N_9567,N_8764,N_7551);
xor U9568 (N_9568,N_7778,N_8732);
nand U9569 (N_9569,N_8486,N_8987);
or U9570 (N_9570,N_8780,N_8935);
xor U9571 (N_9571,N_7644,N_8197);
nor U9572 (N_9572,N_7668,N_7552);
and U9573 (N_9573,N_7964,N_8084);
or U9574 (N_9574,N_8690,N_8859);
or U9575 (N_9575,N_7897,N_8319);
or U9576 (N_9576,N_7795,N_8853);
or U9577 (N_9577,N_8566,N_7719);
nand U9578 (N_9578,N_8211,N_8461);
and U9579 (N_9579,N_8095,N_8430);
nand U9580 (N_9580,N_7966,N_8393);
or U9581 (N_9581,N_8224,N_8930);
nor U9582 (N_9582,N_7989,N_7593);
nand U9583 (N_9583,N_8383,N_7677);
and U9584 (N_9584,N_8083,N_7590);
nand U9585 (N_9585,N_8884,N_7888);
xor U9586 (N_9586,N_8680,N_8052);
nand U9587 (N_9587,N_8222,N_8158);
nand U9588 (N_9588,N_8744,N_8508);
nor U9589 (N_9589,N_8547,N_8895);
and U9590 (N_9590,N_7803,N_7764);
and U9591 (N_9591,N_8599,N_7561);
nand U9592 (N_9592,N_8645,N_8591);
and U9593 (N_9593,N_8539,N_7616);
or U9594 (N_9594,N_8805,N_7981);
nand U9595 (N_9595,N_8660,N_8689);
or U9596 (N_9596,N_7871,N_8912);
nand U9597 (N_9597,N_7858,N_8064);
and U9598 (N_9598,N_8399,N_8401);
nand U9599 (N_9599,N_8713,N_8995);
nor U9600 (N_9600,N_7742,N_7827);
nor U9601 (N_9601,N_8285,N_7905);
nand U9602 (N_9602,N_8621,N_8535);
and U9603 (N_9603,N_8267,N_7941);
nor U9604 (N_9604,N_8236,N_8329);
and U9605 (N_9605,N_8788,N_8040);
nor U9606 (N_9606,N_7812,N_7568);
and U9607 (N_9607,N_7569,N_7886);
or U9608 (N_9608,N_7688,N_8290);
nor U9609 (N_9609,N_8073,N_7766);
nand U9610 (N_9610,N_8916,N_7706);
nand U9611 (N_9611,N_8773,N_8123);
nor U9612 (N_9612,N_8734,N_8562);
nor U9613 (N_9613,N_8933,N_8532);
xnor U9614 (N_9614,N_8736,N_7993);
nor U9615 (N_9615,N_8348,N_7986);
and U9616 (N_9616,N_8380,N_8334);
and U9617 (N_9617,N_7683,N_7698);
nand U9618 (N_9618,N_7517,N_7867);
nand U9619 (N_9619,N_8960,N_7705);
and U9620 (N_9620,N_8656,N_8307);
and U9621 (N_9621,N_8950,N_8746);
and U9622 (N_9622,N_8963,N_8456);
or U9623 (N_9623,N_8683,N_7519);
and U9624 (N_9624,N_8195,N_8968);
and U9625 (N_9625,N_8182,N_8673);
nor U9626 (N_9626,N_7885,N_8241);
nand U9627 (N_9627,N_7933,N_8703);
nor U9628 (N_9628,N_7953,N_8545);
or U9629 (N_9629,N_8335,N_8659);
nor U9630 (N_9630,N_8959,N_8888);
nor U9631 (N_9631,N_8022,N_8479);
nor U9632 (N_9632,N_8988,N_8710);
and U9633 (N_9633,N_8024,N_8986);
and U9634 (N_9634,N_7839,N_7697);
nor U9635 (N_9635,N_8603,N_8634);
or U9636 (N_9636,N_8173,N_8003);
nand U9637 (N_9637,N_8648,N_8863);
or U9638 (N_9638,N_8522,N_8376);
xor U9639 (N_9639,N_8301,N_7559);
nand U9640 (N_9640,N_7848,N_7696);
nor U9641 (N_9641,N_8923,N_8304);
and U9642 (N_9642,N_8247,N_8510);
nor U9643 (N_9643,N_8031,N_8193);
and U9644 (N_9644,N_8122,N_8943);
nand U9645 (N_9645,N_7588,N_7996);
or U9646 (N_9646,N_8238,N_8542);
and U9647 (N_9647,N_7767,N_8739);
and U9648 (N_9648,N_7836,N_8826);
and U9649 (N_9649,N_8907,N_8801);
nor U9650 (N_9650,N_8956,N_8694);
nand U9651 (N_9651,N_8190,N_7657);
nor U9652 (N_9652,N_8490,N_8937);
or U9653 (N_9653,N_8026,N_8168);
and U9654 (N_9654,N_7653,N_8397);
xor U9655 (N_9655,N_7928,N_8281);
nor U9656 (N_9656,N_8546,N_8206);
or U9657 (N_9657,N_8470,N_7681);
nor U9658 (N_9658,N_8802,N_8860);
and U9659 (N_9659,N_8230,N_7735);
and U9660 (N_9660,N_7643,N_8834);
nand U9661 (N_9661,N_7718,N_8806);
xor U9662 (N_9662,N_8761,N_8707);
nor U9663 (N_9663,N_7656,N_7805);
or U9664 (N_9664,N_8706,N_8920);
xnor U9665 (N_9665,N_8402,N_8169);
and U9666 (N_9666,N_7895,N_8013);
and U9667 (N_9667,N_7620,N_8869);
nand U9668 (N_9668,N_8185,N_8418);
or U9669 (N_9669,N_8733,N_7948);
nand U9670 (N_9670,N_8060,N_8177);
nor U9671 (N_9671,N_7577,N_7912);
nor U9672 (N_9672,N_8258,N_8816);
nor U9673 (N_9673,N_8848,N_8029);
and U9674 (N_9674,N_8088,N_7623);
nand U9675 (N_9675,N_8249,N_8389);
nor U9676 (N_9676,N_8686,N_8077);
nand U9677 (N_9677,N_8701,N_8075);
and U9678 (N_9678,N_7896,N_8308);
and U9679 (N_9679,N_7622,N_8885);
or U9680 (N_9680,N_8625,N_7545);
nor U9681 (N_9681,N_7893,N_8832);
nor U9682 (N_9682,N_7605,N_8541);
nor U9683 (N_9683,N_8572,N_8581);
or U9684 (N_9684,N_8558,N_7863);
or U9685 (N_9685,N_8232,N_8239);
and U9686 (N_9686,N_7882,N_7846);
nor U9687 (N_9687,N_8407,N_8718);
and U9688 (N_9688,N_7787,N_8663);
nor U9689 (N_9689,N_8474,N_8644);
nor U9690 (N_9690,N_8904,N_8009);
nor U9691 (N_9691,N_7952,N_7956);
and U9692 (N_9692,N_7730,N_8025);
nor U9693 (N_9693,N_8215,N_8039);
or U9694 (N_9694,N_8365,N_8094);
nor U9695 (N_9695,N_7985,N_7671);
or U9696 (N_9696,N_8262,N_8751);
and U9697 (N_9697,N_8757,N_8288);
or U9698 (N_9698,N_7856,N_7955);
or U9699 (N_9699,N_8803,N_8596);
nor U9700 (N_9700,N_8419,N_8124);
nor U9701 (N_9701,N_7760,N_8272);
or U9702 (N_9702,N_8908,N_8653);
and U9703 (N_9703,N_8017,N_7587);
nand U9704 (N_9704,N_8313,N_7612);
or U9705 (N_9705,N_8894,N_8315);
nor U9706 (N_9706,N_8254,N_8529);
nand U9707 (N_9707,N_8685,N_8180);
xnor U9708 (N_9708,N_7725,N_8178);
nor U9709 (N_9709,N_7531,N_8969);
and U9710 (N_9710,N_8368,N_8350);
or U9711 (N_9711,N_8745,N_8466);
nand U9712 (N_9712,N_7549,N_8688);
nor U9713 (N_9713,N_8341,N_8080);
nand U9714 (N_9714,N_8038,N_8275);
nor U9715 (N_9715,N_8641,N_8257);
nand U9716 (N_9716,N_7936,N_8709);
and U9717 (N_9717,N_7704,N_7758);
and U9718 (N_9718,N_8527,N_8589);
and U9719 (N_9719,N_7874,N_8317);
xor U9720 (N_9720,N_8382,N_8276);
nand U9721 (N_9721,N_7521,N_8127);
nand U9722 (N_9722,N_8866,N_8617);
nor U9723 (N_9723,N_8440,N_7785);
nor U9724 (N_9724,N_7676,N_8837);
xor U9725 (N_9725,N_7546,N_8352);
nor U9726 (N_9726,N_8000,N_8787);
and U9727 (N_9727,N_8594,N_8715);
nor U9728 (N_9728,N_7898,N_8882);
or U9729 (N_9729,N_7627,N_8724);
nand U9730 (N_9730,N_8842,N_8367);
nor U9731 (N_9731,N_7818,N_8107);
nor U9732 (N_9732,N_8463,N_8121);
nand U9733 (N_9733,N_7914,N_8579);
or U9734 (N_9734,N_8153,N_7666);
or U9735 (N_9735,N_7509,N_7691);
nand U9736 (N_9736,N_7997,N_8855);
nor U9737 (N_9737,N_8613,N_8559);
nor U9738 (N_9738,N_8105,N_8999);
or U9739 (N_9739,N_8537,N_8492);
or U9740 (N_9740,N_8729,N_8611);
nor U9741 (N_9741,N_8630,N_8957);
or U9742 (N_9742,N_8901,N_8728);
and U9743 (N_9743,N_8225,N_8485);
nand U9744 (N_9744,N_8010,N_7660);
nand U9745 (N_9745,N_8410,N_7700);
or U9746 (N_9746,N_7755,N_8141);
and U9747 (N_9747,N_8568,N_7503);
or U9748 (N_9748,N_8390,N_8858);
or U9749 (N_9749,N_8992,N_7972);
nor U9750 (N_9750,N_8223,N_8641);
nor U9751 (N_9751,N_7974,N_7866);
nor U9752 (N_9752,N_7580,N_7617);
and U9753 (N_9753,N_8393,N_8271);
nor U9754 (N_9754,N_8294,N_7561);
nor U9755 (N_9755,N_8168,N_8619);
and U9756 (N_9756,N_8440,N_8266);
and U9757 (N_9757,N_8680,N_8820);
nor U9758 (N_9758,N_8746,N_8328);
and U9759 (N_9759,N_7650,N_8043);
nor U9760 (N_9760,N_8371,N_7692);
nand U9761 (N_9761,N_8834,N_7596);
nor U9762 (N_9762,N_7666,N_8862);
nor U9763 (N_9763,N_7958,N_8316);
and U9764 (N_9764,N_7987,N_8889);
and U9765 (N_9765,N_8056,N_8014);
or U9766 (N_9766,N_7843,N_8129);
nand U9767 (N_9767,N_8980,N_8250);
nor U9768 (N_9768,N_8888,N_8126);
nand U9769 (N_9769,N_8868,N_8452);
and U9770 (N_9770,N_7906,N_7801);
xnor U9771 (N_9771,N_7539,N_8909);
and U9772 (N_9772,N_7781,N_7757);
or U9773 (N_9773,N_7670,N_7528);
or U9774 (N_9774,N_8032,N_8915);
or U9775 (N_9775,N_8606,N_8316);
nor U9776 (N_9776,N_7777,N_7970);
and U9777 (N_9777,N_8061,N_8027);
nor U9778 (N_9778,N_8220,N_7918);
or U9779 (N_9779,N_8980,N_8349);
and U9780 (N_9780,N_8202,N_8151);
or U9781 (N_9781,N_7794,N_8302);
or U9782 (N_9782,N_8212,N_8840);
and U9783 (N_9783,N_8018,N_7775);
nor U9784 (N_9784,N_8582,N_7686);
xnor U9785 (N_9785,N_8227,N_8347);
nor U9786 (N_9786,N_8220,N_8587);
and U9787 (N_9787,N_7608,N_7741);
nand U9788 (N_9788,N_8660,N_8659);
nand U9789 (N_9789,N_8726,N_7719);
and U9790 (N_9790,N_7986,N_7937);
or U9791 (N_9791,N_8756,N_8793);
nor U9792 (N_9792,N_8553,N_7634);
nand U9793 (N_9793,N_8001,N_8763);
or U9794 (N_9794,N_8821,N_7715);
and U9795 (N_9795,N_8395,N_8310);
and U9796 (N_9796,N_8907,N_8002);
nand U9797 (N_9797,N_7888,N_7636);
and U9798 (N_9798,N_8889,N_8045);
xnor U9799 (N_9799,N_7723,N_8891);
and U9800 (N_9800,N_8858,N_8138);
nand U9801 (N_9801,N_8149,N_7630);
and U9802 (N_9802,N_8284,N_8674);
or U9803 (N_9803,N_8233,N_8806);
nand U9804 (N_9804,N_8073,N_7948);
nand U9805 (N_9805,N_8116,N_8095);
or U9806 (N_9806,N_7582,N_8129);
nor U9807 (N_9807,N_8790,N_8044);
or U9808 (N_9808,N_8932,N_8164);
or U9809 (N_9809,N_8918,N_8211);
xnor U9810 (N_9810,N_8220,N_8939);
nand U9811 (N_9811,N_7923,N_7648);
or U9812 (N_9812,N_8296,N_8493);
and U9813 (N_9813,N_7916,N_7621);
and U9814 (N_9814,N_7831,N_7503);
and U9815 (N_9815,N_8284,N_8214);
nor U9816 (N_9816,N_7614,N_8543);
xnor U9817 (N_9817,N_7665,N_7895);
and U9818 (N_9818,N_8264,N_8841);
nor U9819 (N_9819,N_8549,N_7795);
or U9820 (N_9820,N_8710,N_8496);
or U9821 (N_9821,N_8749,N_7685);
and U9822 (N_9822,N_8471,N_8054);
nand U9823 (N_9823,N_7970,N_8576);
nor U9824 (N_9824,N_8543,N_7647);
or U9825 (N_9825,N_7618,N_7583);
or U9826 (N_9826,N_8676,N_8954);
nor U9827 (N_9827,N_8523,N_7965);
and U9828 (N_9828,N_8135,N_8302);
nor U9829 (N_9829,N_7740,N_7871);
nand U9830 (N_9830,N_7955,N_8302);
nor U9831 (N_9831,N_8409,N_8679);
and U9832 (N_9832,N_7944,N_8684);
nor U9833 (N_9833,N_8957,N_7712);
and U9834 (N_9834,N_8287,N_8783);
and U9835 (N_9835,N_8848,N_8067);
and U9836 (N_9836,N_8098,N_8600);
nand U9837 (N_9837,N_8999,N_7955);
or U9838 (N_9838,N_8816,N_8287);
and U9839 (N_9839,N_7995,N_7927);
and U9840 (N_9840,N_8010,N_7757);
nor U9841 (N_9841,N_7571,N_7634);
nor U9842 (N_9842,N_8993,N_7801);
and U9843 (N_9843,N_7623,N_8468);
nand U9844 (N_9844,N_7672,N_8073);
nor U9845 (N_9845,N_8326,N_8119);
nor U9846 (N_9846,N_7858,N_8853);
and U9847 (N_9847,N_8094,N_8977);
nand U9848 (N_9848,N_8789,N_7916);
or U9849 (N_9849,N_8640,N_8707);
nand U9850 (N_9850,N_8875,N_8505);
and U9851 (N_9851,N_7999,N_8734);
nor U9852 (N_9852,N_8393,N_7909);
or U9853 (N_9853,N_8223,N_8194);
and U9854 (N_9854,N_8561,N_8180);
or U9855 (N_9855,N_8878,N_8073);
nor U9856 (N_9856,N_7653,N_8358);
or U9857 (N_9857,N_8644,N_8280);
nor U9858 (N_9858,N_7809,N_7978);
and U9859 (N_9859,N_7883,N_7688);
xor U9860 (N_9860,N_7971,N_8870);
or U9861 (N_9861,N_8110,N_8099);
and U9862 (N_9862,N_8280,N_7810);
nand U9863 (N_9863,N_7525,N_7656);
nand U9864 (N_9864,N_8042,N_8705);
and U9865 (N_9865,N_8616,N_8330);
or U9866 (N_9866,N_8021,N_8784);
xor U9867 (N_9867,N_8865,N_7975);
and U9868 (N_9868,N_8855,N_8875);
nand U9869 (N_9869,N_7726,N_8862);
nor U9870 (N_9870,N_7935,N_8659);
nand U9871 (N_9871,N_8802,N_8943);
or U9872 (N_9872,N_8095,N_8021);
and U9873 (N_9873,N_7592,N_8794);
nand U9874 (N_9874,N_7891,N_8892);
or U9875 (N_9875,N_7931,N_8335);
or U9876 (N_9876,N_8905,N_8371);
or U9877 (N_9877,N_8082,N_8587);
and U9878 (N_9878,N_7888,N_7949);
nor U9879 (N_9879,N_8198,N_7892);
or U9880 (N_9880,N_7824,N_8507);
nor U9881 (N_9881,N_8290,N_8841);
and U9882 (N_9882,N_8997,N_8145);
nor U9883 (N_9883,N_8423,N_8095);
nand U9884 (N_9884,N_8785,N_8776);
nand U9885 (N_9885,N_8096,N_8273);
or U9886 (N_9886,N_8579,N_8874);
nand U9887 (N_9887,N_8311,N_8212);
nor U9888 (N_9888,N_8208,N_8189);
or U9889 (N_9889,N_7752,N_8883);
nor U9890 (N_9890,N_8165,N_7784);
nor U9891 (N_9891,N_8459,N_7782);
or U9892 (N_9892,N_8323,N_8661);
or U9893 (N_9893,N_8500,N_7797);
and U9894 (N_9894,N_7789,N_7686);
xor U9895 (N_9895,N_8080,N_7603);
or U9896 (N_9896,N_8292,N_7820);
or U9897 (N_9897,N_8703,N_8460);
and U9898 (N_9898,N_8185,N_7525);
and U9899 (N_9899,N_7559,N_8595);
and U9900 (N_9900,N_7908,N_7572);
nor U9901 (N_9901,N_7562,N_8724);
and U9902 (N_9902,N_8362,N_8737);
and U9903 (N_9903,N_7848,N_7527);
xnor U9904 (N_9904,N_8580,N_7809);
nand U9905 (N_9905,N_7758,N_8242);
nor U9906 (N_9906,N_7917,N_8703);
nor U9907 (N_9907,N_7879,N_7546);
nand U9908 (N_9908,N_7833,N_8063);
and U9909 (N_9909,N_8898,N_8631);
and U9910 (N_9910,N_7952,N_8122);
nand U9911 (N_9911,N_8572,N_8461);
xor U9912 (N_9912,N_8301,N_8175);
and U9913 (N_9913,N_8183,N_8343);
nor U9914 (N_9914,N_8350,N_8789);
and U9915 (N_9915,N_8352,N_7588);
nand U9916 (N_9916,N_8039,N_7937);
and U9917 (N_9917,N_7763,N_8684);
and U9918 (N_9918,N_7903,N_7743);
and U9919 (N_9919,N_8902,N_8258);
nand U9920 (N_9920,N_7891,N_8082);
and U9921 (N_9921,N_7884,N_7616);
and U9922 (N_9922,N_8761,N_7976);
and U9923 (N_9923,N_8503,N_8160);
or U9924 (N_9924,N_8000,N_8094);
nor U9925 (N_9925,N_8649,N_8851);
nor U9926 (N_9926,N_8614,N_8964);
or U9927 (N_9927,N_8328,N_7502);
nand U9928 (N_9928,N_8516,N_7636);
and U9929 (N_9929,N_8609,N_8204);
nor U9930 (N_9930,N_8043,N_8897);
nor U9931 (N_9931,N_8674,N_8693);
and U9932 (N_9932,N_8324,N_8112);
and U9933 (N_9933,N_8415,N_8972);
nand U9934 (N_9934,N_8814,N_7552);
nor U9935 (N_9935,N_8004,N_7902);
xor U9936 (N_9936,N_8015,N_8429);
xnor U9937 (N_9937,N_8793,N_7670);
nor U9938 (N_9938,N_8037,N_8656);
nand U9939 (N_9939,N_8233,N_7684);
xor U9940 (N_9940,N_8010,N_7769);
nand U9941 (N_9941,N_7738,N_8310);
or U9942 (N_9942,N_7952,N_8693);
nand U9943 (N_9943,N_8497,N_7907);
or U9944 (N_9944,N_8667,N_7758);
and U9945 (N_9945,N_8413,N_8006);
nand U9946 (N_9946,N_8685,N_8426);
nand U9947 (N_9947,N_8680,N_8678);
and U9948 (N_9948,N_7918,N_8651);
nor U9949 (N_9949,N_8274,N_8042);
or U9950 (N_9950,N_8982,N_8442);
nand U9951 (N_9951,N_8403,N_8941);
nand U9952 (N_9952,N_7550,N_8282);
and U9953 (N_9953,N_8838,N_8670);
nand U9954 (N_9954,N_7617,N_8241);
and U9955 (N_9955,N_8897,N_8653);
nand U9956 (N_9956,N_8950,N_8159);
nor U9957 (N_9957,N_8408,N_8637);
nor U9958 (N_9958,N_8240,N_8882);
and U9959 (N_9959,N_8042,N_7728);
xnor U9960 (N_9960,N_7758,N_7626);
nand U9961 (N_9961,N_7968,N_8194);
nor U9962 (N_9962,N_8611,N_8107);
nor U9963 (N_9963,N_8586,N_8503);
and U9964 (N_9964,N_8169,N_8794);
or U9965 (N_9965,N_7632,N_7739);
or U9966 (N_9966,N_7699,N_8371);
xor U9967 (N_9967,N_8427,N_7517);
nand U9968 (N_9968,N_8863,N_7596);
or U9969 (N_9969,N_8408,N_7572);
or U9970 (N_9970,N_8937,N_8505);
or U9971 (N_9971,N_8457,N_8209);
or U9972 (N_9972,N_8017,N_8522);
or U9973 (N_9973,N_8763,N_8648);
or U9974 (N_9974,N_8947,N_8430);
nand U9975 (N_9975,N_7972,N_7668);
or U9976 (N_9976,N_7942,N_7665);
or U9977 (N_9977,N_7965,N_8632);
nand U9978 (N_9978,N_8102,N_7505);
nand U9979 (N_9979,N_8309,N_7934);
nor U9980 (N_9980,N_8810,N_8490);
nor U9981 (N_9981,N_8329,N_8155);
nand U9982 (N_9982,N_8995,N_8802);
nor U9983 (N_9983,N_8756,N_8214);
or U9984 (N_9984,N_7504,N_8985);
or U9985 (N_9985,N_8200,N_8598);
and U9986 (N_9986,N_7840,N_8951);
nand U9987 (N_9987,N_8505,N_8408);
nand U9988 (N_9988,N_8192,N_7653);
or U9989 (N_9989,N_7988,N_8678);
or U9990 (N_9990,N_8251,N_7877);
nor U9991 (N_9991,N_8609,N_8848);
and U9992 (N_9992,N_7752,N_7672);
or U9993 (N_9993,N_7790,N_7791);
nor U9994 (N_9994,N_8060,N_7816);
or U9995 (N_9995,N_7968,N_7958);
and U9996 (N_9996,N_7553,N_8884);
or U9997 (N_9997,N_8104,N_8903);
or U9998 (N_9998,N_8227,N_8890);
nand U9999 (N_9999,N_8461,N_7783);
xnor U10000 (N_10000,N_7886,N_8378);
xnor U10001 (N_10001,N_8653,N_7738);
xnor U10002 (N_10002,N_7630,N_8913);
or U10003 (N_10003,N_8498,N_8367);
or U10004 (N_10004,N_7674,N_8081);
xor U10005 (N_10005,N_8406,N_8027);
xor U10006 (N_10006,N_8711,N_8802);
and U10007 (N_10007,N_8469,N_8709);
nand U10008 (N_10008,N_8839,N_8583);
or U10009 (N_10009,N_7621,N_8838);
or U10010 (N_10010,N_8375,N_7726);
nand U10011 (N_10011,N_7766,N_8010);
nor U10012 (N_10012,N_7975,N_8272);
nand U10013 (N_10013,N_7557,N_7706);
and U10014 (N_10014,N_7507,N_8863);
nor U10015 (N_10015,N_7820,N_7501);
xnor U10016 (N_10016,N_8723,N_8346);
nand U10017 (N_10017,N_8491,N_8426);
xor U10018 (N_10018,N_8102,N_8228);
or U10019 (N_10019,N_7549,N_8058);
and U10020 (N_10020,N_8971,N_8625);
nand U10021 (N_10021,N_8199,N_8874);
and U10022 (N_10022,N_8699,N_8938);
nand U10023 (N_10023,N_7836,N_8321);
or U10024 (N_10024,N_7893,N_8390);
nand U10025 (N_10025,N_8114,N_8146);
nor U10026 (N_10026,N_7812,N_8935);
nand U10027 (N_10027,N_8238,N_8516);
or U10028 (N_10028,N_8971,N_8263);
nand U10029 (N_10029,N_8506,N_8953);
and U10030 (N_10030,N_7548,N_8148);
and U10031 (N_10031,N_8969,N_8761);
and U10032 (N_10032,N_7780,N_7979);
xor U10033 (N_10033,N_7658,N_8685);
or U10034 (N_10034,N_8115,N_8422);
xor U10035 (N_10035,N_8058,N_8840);
nand U10036 (N_10036,N_8016,N_8167);
nand U10037 (N_10037,N_8473,N_8228);
or U10038 (N_10038,N_8190,N_8408);
and U10039 (N_10039,N_8315,N_8743);
or U10040 (N_10040,N_8063,N_8963);
or U10041 (N_10041,N_8625,N_8105);
nor U10042 (N_10042,N_8540,N_7763);
or U10043 (N_10043,N_8445,N_7956);
or U10044 (N_10044,N_8104,N_7768);
and U10045 (N_10045,N_8594,N_8986);
xnor U10046 (N_10046,N_7692,N_7542);
and U10047 (N_10047,N_8355,N_7982);
nand U10048 (N_10048,N_8153,N_8885);
nor U10049 (N_10049,N_8863,N_8668);
nor U10050 (N_10050,N_7849,N_8910);
nor U10051 (N_10051,N_7718,N_7814);
and U10052 (N_10052,N_7978,N_7800);
and U10053 (N_10053,N_7621,N_8382);
and U10054 (N_10054,N_8179,N_7576);
xnor U10055 (N_10055,N_8485,N_8758);
or U10056 (N_10056,N_7581,N_8720);
and U10057 (N_10057,N_8050,N_8131);
or U10058 (N_10058,N_7516,N_8849);
xor U10059 (N_10059,N_8851,N_8803);
or U10060 (N_10060,N_8697,N_8396);
nor U10061 (N_10061,N_8254,N_7570);
or U10062 (N_10062,N_7529,N_7837);
nand U10063 (N_10063,N_7718,N_7692);
and U10064 (N_10064,N_8581,N_8627);
xnor U10065 (N_10065,N_8980,N_8233);
or U10066 (N_10066,N_8143,N_8718);
or U10067 (N_10067,N_8077,N_7817);
and U10068 (N_10068,N_7575,N_8856);
nand U10069 (N_10069,N_8353,N_7902);
nand U10070 (N_10070,N_7565,N_8188);
xnor U10071 (N_10071,N_7690,N_8994);
and U10072 (N_10072,N_8040,N_8047);
nand U10073 (N_10073,N_8325,N_8158);
nor U10074 (N_10074,N_8407,N_7986);
or U10075 (N_10075,N_7840,N_7845);
or U10076 (N_10076,N_8909,N_8492);
or U10077 (N_10077,N_7530,N_8401);
nand U10078 (N_10078,N_8178,N_8511);
and U10079 (N_10079,N_8323,N_8351);
nand U10080 (N_10080,N_7906,N_7758);
nand U10081 (N_10081,N_8200,N_8538);
or U10082 (N_10082,N_8447,N_7747);
or U10083 (N_10083,N_8450,N_8322);
xor U10084 (N_10084,N_8036,N_7514);
and U10085 (N_10085,N_8549,N_7637);
nand U10086 (N_10086,N_8465,N_7885);
nand U10087 (N_10087,N_8582,N_8476);
xor U10088 (N_10088,N_8230,N_7833);
nor U10089 (N_10089,N_7891,N_8708);
nor U10090 (N_10090,N_7619,N_7658);
or U10091 (N_10091,N_7756,N_7849);
nand U10092 (N_10092,N_8344,N_8601);
and U10093 (N_10093,N_8382,N_8595);
xnor U10094 (N_10094,N_7598,N_8022);
nor U10095 (N_10095,N_8721,N_8402);
and U10096 (N_10096,N_8518,N_8110);
nor U10097 (N_10097,N_8516,N_8275);
and U10098 (N_10098,N_8914,N_8074);
or U10099 (N_10099,N_7598,N_8142);
nor U10100 (N_10100,N_7872,N_8080);
nor U10101 (N_10101,N_8249,N_8180);
nor U10102 (N_10102,N_8108,N_8596);
nand U10103 (N_10103,N_8110,N_8806);
and U10104 (N_10104,N_8570,N_7981);
nand U10105 (N_10105,N_8891,N_7899);
and U10106 (N_10106,N_8196,N_7843);
and U10107 (N_10107,N_8953,N_7575);
nor U10108 (N_10108,N_8149,N_8361);
and U10109 (N_10109,N_8666,N_8537);
nor U10110 (N_10110,N_7857,N_8806);
nor U10111 (N_10111,N_8711,N_8900);
and U10112 (N_10112,N_8378,N_8367);
and U10113 (N_10113,N_7646,N_8778);
or U10114 (N_10114,N_8161,N_8267);
nor U10115 (N_10115,N_8086,N_8528);
or U10116 (N_10116,N_7573,N_8523);
nor U10117 (N_10117,N_7824,N_8282);
nand U10118 (N_10118,N_8059,N_8468);
or U10119 (N_10119,N_7944,N_8501);
nor U10120 (N_10120,N_8798,N_8132);
nand U10121 (N_10121,N_7537,N_8504);
or U10122 (N_10122,N_7653,N_7955);
nor U10123 (N_10123,N_8080,N_8822);
xnor U10124 (N_10124,N_8614,N_8001);
nand U10125 (N_10125,N_8192,N_8927);
and U10126 (N_10126,N_8864,N_8429);
and U10127 (N_10127,N_8161,N_7606);
nand U10128 (N_10128,N_8193,N_7627);
xor U10129 (N_10129,N_8057,N_8532);
nand U10130 (N_10130,N_7960,N_7598);
and U10131 (N_10131,N_8130,N_7915);
or U10132 (N_10132,N_8271,N_8103);
and U10133 (N_10133,N_8169,N_8685);
nor U10134 (N_10134,N_8193,N_8686);
or U10135 (N_10135,N_8652,N_8663);
or U10136 (N_10136,N_7661,N_8345);
and U10137 (N_10137,N_8560,N_8985);
nor U10138 (N_10138,N_8793,N_8308);
nor U10139 (N_10139,N_8417,N_8788);
and U10140 (N_10140,N_8820,N_7930);
nand U10141 (N_10141,N_8004,N_7617);
nor U10142 (N_10142,N_8060,N_8668);
and U10143 (N_10143,N_7837,N_8225);
or U10144 (N_10144,N_8530,N_8177);
nand U10145 (N_10145,N_7817,N_8041);
nand U10146 (N_10146,N_8723,N_8832);
nor U10147 (N_10147,N_8503,N_8793);
nand U10148 (N_10148,N_7764,N_7965);
nor U10149 (N_10149,N_7806,N_8741);
nor U10150 (N_10150,N_7890,N_8030);
and U10151 (N_10151,N_8403,N_8003);
and U10152 (N_10152,N_7540,N_8260);
xnor U10153 (N_10153,N_7833,N_8755);
nand U10154 (N_10154,N_7862,N_7584);
nor U10155 (N_10155,N_7532,N_7836);
nand U10156 (N_10156,N_8055,N_7875);
xor U10157 (N_10157,N_8073,N_7523);
or U10158 (N_10158,N_8159,N_8794);
or U10159 (N_10159,N_7993,N_8373);
xnor U10160 (N_10160,N_8899,N_7743);
nor U10161 (N_10161,N_8149,N_8718);
or U10162 (N_10162,N_8927,N_7819);
xnor U10163 (N_10163,N_7580,N_7839);
xor U10164 (N_10164,N_8127,N_8079);
and U10165 (N_10165,N_8263,N_8199);
nor U10166 (N_10166,N_8004,N_8274);
xor U10167 (N_10167,N_8332,N_8337);
and U10168 (N_10168,N_8996,N_7513);
and U10169 (N_10169,N_8802,N_8849);
and U10170 (N_10170,N_8428,N_7756);
or U10171 (N_10171,N_8707,N_8019);
and U10172 (N_10172,N_8364,N_8402);
and U10173 (N_10173,N_8784,N_8227);
xnor U10174 (N_10174,N_8112,N_8214);
and U10175 (N_10175,N_7847,N_8448);
nor U10176 (N_10176,N_8365,N_7598);
or U10177 (N_10177,N_7853,N_8637);
nand U10178 (N_10178,N_7560,N_8723);
or U10179 (N_10179,N_8895,N_7680);
nor U10180 (N_10180,N_8501,N_7987);
or U10181 (N_10181,N_8241,N_7921);
and U10182 (N_10182,N_8699,N_7750);
or U10183 (N_10183,N_7731,N_7946);
or U10184 (N_10184,N_8514,N_8423);
xnor U10185 (N_10185,N_7505,N_8006);
nand U10186 (N_10186,N_7600,N_7959);
or U10187 (N_10187,N_7612,N_7990);
xor U10188 (N_10188,N_8677,N_8112);
nand U10189 (N_10189,N_8898,N_8135);
or U10190 (N_10190,N_7931,N_7600);
or U10191 (N_10191,N_8676,N_8142);
or U10192 (N_10192,N_8696,N_7821);
and U10193 (N_10193,N_8891,N_8404);
nor U10194 (N_10194,N_8755,N_8801);
nor U10195 (N_10195,N_8627,N_7630);
nand U10196 (N_10196,N_8063,N_7988);
nand U10197 (N_10197,N_8464,N_8721);
or U10198 (N_10198,N_7548,N_7776);
nand U10199 (N_10199,N_8892,N_7598);
or U10200 (N_10200,N_8852,N_8931);
or U10201 (N_10201,N_8993,N_7664);
and U10202 (N_10202,N_8601,N_7787);
nor U10203 (N_10203,N_8021,N_8137);
or U10204 (N_10204,N_7678,N_8006);
xnor U10205 (N_10205,N_8994,N_7692);
or U10206 (N_10206,N_8230,N_8996);
nand U10207 (N_10207,N_8497,N_7848);
nand U10208 (N_10208,N_7526,N_7577);
nor U10209 (N_10209,N_8338,N_8644);
or U10210 (N_10210,N_8089,N_8535);
nand U10211 (N_10211,N_7954,N_8977);
nand U10212 (N_10212,N_8554,N_7796);
and U10213 (N_10213,N_8107,N_8232);
or U10214 (N_10214,N_8636,N_7678);
nor U10215 (N_10215,N_8371,N_8016);
or U10216 (N_10216,N_7892,N_8976);
xor U10217 (N_10217,N_8381,N_7515);
and U10218 (N_10218,N_8904,N_7903);
xor U10219 (N_10219,N_8968,N_7839);
nand U10220 (N_10220,N_8707,N_7922);
and U10221 (N_10221,N_8039,N_8613);
and U10222 (N_10222,N_8925,N_8022);
and U10223 (N_10223,N_7895,N_8391);
and U10224 (N_10224,N_8916,N_8099);
nor U10225 (N_10225,N_7766,N_8472);
nand U10226 (N_10226,N_8095,N_7528);
and U10227 (N_10227,N_8223,N_8354);
and U10228 (N_10228,N_8781,N_7979);
nand U10229 (N_10229,N_8498,N_7522);
or U10230 (N_10230,N_8954,N_7900);
nor U10231 (N_10231,N_7696,N_8240);
and U10232 (N_10232,N_8096,N_8191);
nor U10233 (N_10233,N_8835,N_8150);
or U10234 (N_10234,N_8507,N_8266);
or U10235 (N_10235,N_7899,N_8412);
nand U10236 (N_10236,N_8251,N_8897);
and U10237 (N_10237,N_8993,N_8561);
and U10238 (N_10238,N_8291,N_8709);
nand U10239 (N_10239,N_7769,N_7833);
and U10240 (N_10240,N_7886,N_8636);
or U10241 (N_10241,N_7603,N_8402);
or U10242 (N_10242,N_8470,N_8104);
xor U10243 (N_10243,N_8292,N_8160);
nor U10244 (N_10244,N_8228,N_7970);
and U10245 (N_10245,N_7891,N_8936);
and U10246 (N_10246,N_8688,N_8578);
nand U10247 (N_10247,N_8396,N_8519);
and U10248 (N_10248,N_8858,N_8416);
and U10249 (N_10249,N_8196,N_8429);
nor U10250 (N_10250,N_8878,N_7517);
or U10251 (N_10251,N_8848,N_8224);
or U10252 (N_10252,N_8270,N_8812);
and U10253 (N_10253,N_8195,N_7529);
or U10254 (N_10254,N_7988,N_8971);
and U10255 (N_10255,N_8421,N_8592);
nor U10256 (N_10256,N_7531,N_7633);
nor U10257 (N_10257,N_8772,N_8094);
or U10258 (N_10258,N_8970,N_8161);
or U10259 (N_10259,N_8990,N_7889);
or U10260 (N_10260,N_7597,N_7999);
and U10261 (N_10261,N_7507,N_8394);
and U10262 (N_10262,N_8626,N_7770);
and U10263 (N_10263,N_7662,N_7501);
nor U10264 (N_10264,N_8580,N_8756);
nor U10265 (N_10265,N_8833,N_8953);
xnor U10266 (N_10266,N_7899,N_7729);
or U10267 (N_10267,N_8705,N_8186);
xnor U10268 (N_10268,N_8244,N_8333);
and U10269 (N_10269,N_8479,N_7783);
and U10270 (N_10270,N_7761,N_8054);
or U10271 (N_10271,N_8029,N_8597);
nor U10272 (N_10272,N_8838,N_8321);
nor U10273 (N_10273,N_7868,N_8113);
or U10274 (N_10274,N_8314,N_8128);
or U10275 (N_10275,N_7814,N_8668);
and U10276 (N_10276,N_8194,N_7675);
and U10277 (N_10277,N_8122,N_8408);
nand U10278 (N_10278,N_7678,N_8576);
and U10279 (N_10279,N_8767,N_8232);
and U10280 (N_10280,N_8013,N_8361);
nand U10281 (N_10281,N_8172,N_8765);
nor U10282 (N_10282,N_8360,N_8645);
or U10283 (N_10283,N_8157,N_8651);
nand U10284 (N_10284,N_8669,N_8261);
nor U10285 (N_10285,N_7647,N_8494);
and U10286 (N_10286,N_8740,N_8876);
nand U10287 (N_10287,N_8789,N_8006);
nand U10288 (N_10288,N_7698,N_8850);
nor U10289 (N_10289,N_8613,N_8679);
or U10290 (N_10290,N_8791,N_8496);
or U10291 (N_10291,N_7856,N_8535);
xor U10292 (N_10292,N_7742,N_8483);
or U10293 (N_10293,N_8449,N_8791);
and U10294 (N_10294,N_7713,N_8589);
nand U10295 (N_10295,N_7672,N_8191);
or U10296 (N_10296,N_8972,N_7869);
nor U10297 (N_10297,N_7914,N_7658);
and U10298 (N_10298,N_7818,N_8949);
xnor U10299 (N_10299,N_8388,N_8124);
and U10300 (N_10300,N_7605,N_8257);
or U10301 (N_10301,N_8022,N_7635);
and U10302 (N_10302,N_7860,N_8392);
nor U10303 (N_10303,N_8798,N_8106);
or U10304 (N_10304,N_7986,N_8117);
and U10305 (N_10305,N_8771,N_8384);
or U10306 (N_10306,N_8770,N_8852);
or U10307 (N_10307,N_8025,N_7783);
and U10308 (N_10308,N_8637,N_7611);
nor U10309 (N_10309,N_7826,N_7625);
xor U10310 (N_10310,N_8384,N_8742);
xnor U10311 (N_10311,N_7780,N_8506);
nand U10312 (N_10312,N_8168,N_8938);
or U10313 (N_10313,N_8488,N_7506);
nor U10314 (N_10314,N_8939,N_7509);
nand U10315 (N_10315,N_8181,N_8464);
and U10316 (N_10316,N_7616,N_7585);
or U10317 (N_10317,N_8793,N_8770);
nand U10318 (N_10318,N_8470,N_7539);
xnor U10319 (N_10319,N_8259,N_7544);
or U10320 (N_10320,N_8786,N_8327);
nand U10321 (N_10321,N_8542,N_8905);
or U10322 (N_10322,N_8065,N_8091);
or U10323 (N_10323,N_8603,N_8654);
nand U10324 (N_10324,N_8749,N_8634);
and U10325 (N_10325,N_8477,N_8157);
nand U10326 (N_10326,N_8136,N_8188);
or U10327 (N_10327,N_8714,N_8048);
nor U10328 (N_10328,N_8391,N_8007);
xnor U10329 (N_10329,N_7552,N_8968);
or U10330 (N_10330,N_7510,N_8011);
nand U10331 (N_10331,N_8669,N_8839);
xor U10332 (N_10332,N_7709,N_8933);
nor U10333 (N_10333,N_7723,N_8948);
or U10334 (N_10334,N_7827,N_8059);
or U10335 (N_10335,N_8320,N_8693);
nand U10336 (N_10336,N_8912,N_7934);
nor U10337 (N_10337,N_7526,N_8794);
nor U10338 (N_10338,N_8671,N_8189);
or U10339 (N_10339,N_8902,N_8704);
nor U10340 (N_10340,N_7717,N_7782);
or U10341 (N_10341,N_8643,N_8117);
or U10342 (N_10342,N_8351,N_8484);
nor U10343 (N_10343,N_8876,N_8430);
or U10344 (N_10344,N_7713,N_8066);
nor U10345 (N_10345,N_7644,N_8746);
xnor U10346 (N_10346,N_8489,N_7857);
or U10347 (N_10347,N_8565,N_8560);
or U10348 (N_10348,N_7622,N_7508);
or U10349 (N_10349,N_8817,N_8066);
or U10350 (N_10350,N_7845,N_7764);
or U10351 (N_10351,N_8268,N_7697);
or U10352 (N_10352,N_7740,N_7845);
nand U10353 (N_10353,N_8604,N_8047);
nor U10354 (N_10354,N_8723,N_8657);
and U10355 (N_10355,N_7752,N_7665);
and U10356 (N_10356,N_7696,N_8646);
nand U10357 (N_10357,N_7972,N_7968);
nand U10358 (N_10358,N_7684,N_8214);
or U10359 (N_10359,N_8448,N_8951);
and U10360 (N_10360,N_8052,N_8368);
nand U10361 (N_10361,N_7826,N_8835);
and U10362 (N_10362,N_8876,N_7775);
and U10363 (N_10363,N_7612,N_7953);
xnor U10364 (N_10364,N_8050,N_8883);
nor U10365 (N_10365,N_8648,N_8116);
nand U10366 (N_10366,N_7877,N_8132);
and U10367 (N_10367,N_8945,N_8030);
or U10368 (N_10368,N_8555,N_8172);
nor U10369 (N_10369,N_8451,N_8541);
or U10370 (N_10370,N_8277,N_8528);
or U10371 (N_10371,N_8135,N_8936);
and U10372 (N_10372,N_8731,N_7569);
and U10373 (N_10373,N_8495,N_7900);
xnor U10374 (N_10374,N_7660,N_7581);
nand U10375 (N_10375,N_7802,N_7748);
and U10376 (N_10376,N_7631,N_8887);
and U10377 (N_10377,N_7742,N_8182);
or U10378 (N_10378,N_8615,N_7540);
or U10379 (N_10379,N_8667,N_8087);
or U10380 (N_10380,N_8651,N_7962);
and U10381 (N_10381,N_8357,N_7685);
and U10382 (N_10382,N_8381,N_8882);
nand U10383 (N_10383,N_7886,N_8735);
and U10384 (N_10384,N_7663,N_7856);
nand U10385 (N_10385,N_7896,N_8370);
and U10386 (N_10386,N_8039,N_7983);
and U10387 (N_10387,N_7524,N_8796);
nand U10388 (N_10388,N_8528,N_8106);
xnor U10389 (N_10389,N_8919,N_8864);
and U10390 (N_10390,N_8792,N_7887);
nor U10391 (N_10391,N_8172,N_8844);
or U10392 (N_10392,N_7865,N_8993);
and U10393 (N_10393,N_7985,N_7504);
and U10394 (N_10394,N_8621,N_8515);
and U10395 (N_10395,N_8177,N_7620);
nand U10396 (N_10396,N_8455,N_7711);
nor U10397 (N_10397,N_8261,N_8868);
nand U10398 (N_10398,N_8817,N_8295);
xor U10399 (N_10399,N_8697,N_7522);
nand U10400 (N_10400,N_8682,N_8561);
and U10401 (N_10401,N_8775,N_8905);
or U10402 (N_10402,N_8348,N_8383);
and U10403 (N_10403,N_8114,N_7745);
nor U10404 (N_10404,N_8843,N_8223);
nor U10405 (N_10405,N_8675,N_7911);
or U10406 (N_10406,N_7997,N_8911);
or U10407 (N_10407,N_8084,N_7512);
or U10408 (N_10408,N_8191,N_8677);
and U10409 (N_10409,N_7888,N_8262);
nand U10410 (N_10410,N_8934,N_8846);
and U10411 (N_10411,N_8936,N_8251);
nor U10412 (N_10412,N_8293,N_8562);
nand U10413 (N_10413,N_7847,N_8639);
nand U10414 (N_10414,N_8114,N_8667);
nand U10415 (N_10415,N_8019,N_7628);
xor U10416 (N_10416,N_8197,N_8426);
or U10417 (N_10417,N_7614,N_7861);
and U10418 (N_10418,N_8564,N_7938);
nor U10419 (N_10419,N_8711,N_8834);
nand U10420 (N_10420,N_8714,N_8842);
or U10421 (N_10421,N_8147,N_8600);
and U10422 (N_10422,N_8003,N_8259);
or U10423 (N_10423,N_8854,N_7596);
and U10424 (N_10424,N_7937,N_8527);
and U10425 (N_10425,N_8721,N_8319);
nand U10426 (N_10426,N_7819,N_7533);
or U10427 (N_10427,N_8069,N_8739);
and U10428 (N_10428,N_7969,N_7958);
nor U10429 (N_10429,N_8893,N_8905);
or U10430 (N_10430,N_8723,N_7926);
nor U10431 (N_10431,N_8146,N_8565);
and U10432 (N_10432,N_8386,N_7710);
nor U10433 (N_10433,N_8978,N_8726);
or U10434 (N_10434,N_8558,N_7684);
and U10435 (N_10435,N_8649,N_7882);
nand U10436 (N_10436,N_8144,N_8803);
nand U10437 (N_10437,N_8878,N_8431);
nor U10438 (N_10438,N_8456,N_7793);
nor U10439 (N_10439,N_8475,N_8986);
nor U10440 (N_10440,N_8012,N_8614);
or U10441 (N_10441,N_7964,N_8270);
nand U10442 (N_10442,N_8678,N_8496);
and U10443 (N_10443,N_7531,N_7855);
nor U10444 (N_10444,N_7515,N_7928);
and U10445 (N_10445,N_8345,N_8476);
and U10446 (N_10446,N_8531,N_8688);
nor U10447 (N_10447,N_8055,N_8490);
nand U10448 (N_10448,N_8727,N_8037);
nand U10449 (N_10449,N_7724,N_8661);
or U10450 (N_10450,N_7514,N_8696);
nand U10451 (N_10451,N_7570,N_8960);
xor U10452 (N_10452,N_8244,N_7713);
or U10453 (N_10453,N_7554,N_8055);
nand U10454 (N_10454,N_8091,N_8926);
and U10455 (N_10455,N_8483,N_7830);
nor U10456 (N_10456,N_8317,N_8323);
nand U10457 (N_10457,N_8391,N_8562);
xor U10458 (N_10458,N_8367,N_8986);
nand U10459 (N_10459,N_8544,N_8343);
and U10460 (N_10460,N_8882,N_7789);
xnor U10461 (N_10461,N_8800,N_8163);
nor U10462 (N_10462,N_8189,N_8306);
nor U10463 (N_10463,N_8527,N_8425);
nand U10464 (N_10464,N_7968,N_7918);
and U10465 (N_10465,N_8382,N_8579);
nor U10466 (N_10466,N_8099,N_8985);
nand U10467 (N_10467,N_7952,N_8338);
or U10468 (N_10468,N_8915,N_8085);
nor U10469 (N_10469,N_8582,N_8330);
and U10470 (N_10470,N_8558,N_8269);
nand U10471 (N_10471,N_8284,N_8986);
and U10472 (N_10472,N_8702,N_8107);
or U10473 (N_10473,N_8585,N_7933);
and U10474 (N_10474,N_8342,N_8194);
and U10475 (N_10475,N_7811,N_8486);
xnor U10476 (N_10476,N_8183,N_8279);
and U10477 (N_10477,N_7662,N_8218);
nand U10478 (N_10478,N_8151,N_7621);
and U10479 (N_10479,N_7543,N_8016);
nand U10480 (N_10480,N_8995,N_7521);
xnor U10481 (N_10481,N_8098,N_8367);
and U10482 (N_10482,N_8360,N_7915);
nor U10483 (N_10483,N_8243,N_7690);
nor U10484 (N_10484,N_8560,N_8334);
nand U10485 (N_10485,N_8332,N_8778);
or U10486 (N_10486,N_8991,N_8694);
or U10487 (N_10487,N_7532,N_7725);
nand U10488 (N_10488,N_7564,N_8645);
and U10489 (N_10489,N_7951,N_8561);
nor U10490 (N_10490,N_8246,N_8462);
or U10491 (N_10491,N_7527,N_8115);
or U10492 (N_10492,N_8265,N_8311);
or U10493 (N_10493,N_8535,N_7635);
nor U10494 (N_10494,N_8679,N_8968);
or U10495 (N_10495,N_8521,N_8067);
nand U10496 (N_10496,N_8230,N_7789);
nand U10497 (N_10497,N_8958,N_8013);
nor U10498 (N_10498,N_8459,N_8536);
nand U10499 (N_10499,N_7920,N_7713);
and U10500 (N_10500,N_9011,N_10217);
or U10501 (N_10501,N_9534,N_10036);
or U10502 (N_10502,N_9943,N_10301);
nor U10503 (N_10503,N_9009,N_9296);
or U10504 (N_10504,N_9406,N_9300);
nor U10505 (N_10505,N_10427,N_9561);
nor U10506 (N_10506,N_9007,N_10133);
xor U10507 (N_10507,N_9759,N_10314);
or U10508 (N_10508,N_10222,N_10086);
nand U10509 (N_10509,N_9301,N_10077);
or U10510 (N_10510,N_9717,N_10138);
and U10511 (N_10511,N_9680,N_10363);
and U10512 (N_10512,N_9601,N_9085);
nor U10513 (N_10513,N_9062,N_10078);
nor U10514 (N_10514,N_10203,N_10058);
nand U10515 (N_10515,N_9971,N_9151);
nor U10516 (N_10516,N_9161,N_9502);
or U10517 (N_10517,N_9849,N_10475);
and U10518 (N_10518,N_9469,N_9321);
nor U10519 (N_10519,N_9729,N_10052);
nor U10520 (N_10520,N_10282,N_9076);
nor U10521 (N_10521,N_10247,N_9059);
nand U10522 (N_10522,N_9380,N_9565);
nand U10523 (N_10523,N_9265,N_9612);
nand U10524 (N_10524,N_10229,N_10408);
and U10525 (N_10525,N_9579,N_9042);
or U10526 (N_10526,N_10180,N_9397);
nand U10527 (N_10527,N_9533,N_9434);
nand U10528 (N_10528,N_10249,N_9274);
or U10529 (N_10529,N_9547,N_9412);
or U10530 (N_10530,N_10371,N_10354);
and U10531 (N_10531,N_10070,N_9213);
nor U10532 (N_10532,N_9550,N_9889);
or U10533 (N_10533,N_9431,N_9463);
or U10534 (N_10534,N_9825,N_9629);
nor U10535 (N_10535,N_9168,N_10144);
nor U10536 (N_10536,N_9900,N_9086);
nand U10537 (N_10537,N_9493,N_10392);
and U10538 (N_10538,N_9836,N_9455);
and U10539 (N_10539,N_10029,N_9883);
xor U10540 (N_10540,N_9590,N_9003);
and U10541 (N_10541,N_10009,N_9818);
nand U10542 (N_10542,N_10318,N_9134);
nor U10543 (N_10543,N_10104,N_10380);
or U10544 (N_10544,N_9553,N_9722);
and U10545 (N_10545,N_9893,N_10485);
and U10546 (N_10546,N_10178,N_10147);
nor U10547 (N_10547,N_10093,N_10400);
nor U10548 (N_10548,N_10121,N_10342);
nand U10549 (N_10549,N_9145,N_9864);
nand U10550 (N_10550,N_9284,N_9154);
and U10551 (N_10551,N_10436,N_10228);
nor U10552 (N_10552,N_10462,N_9377);
and U10553 (N_10553,N_10418,N_10351);
nand U10554 (N_10554,N_10328,N_10098);
xor U10555 (N_10555,N_9555,N_9255);
and U10556 (N_10556,N_9277,N_9209);
and U10557 (N_10557,N_9813,N_9230);
nand U10558 (N_10558,N_10488,N_9593);
nand U10559 (N_10559,N_9211,N_10304);
nand U10560 (N_10560,N_9551,N_9904);
nor U10561 (N_10561,N_9030,N_10306);
or U10562 (N_10562,N_9917,N_9994);
and U10563 (N_10563,N_9395,N_9914);
nor U10564 (N_10564,N_9632,N_9851);
or U10565 (N_10565,N_10442,N_9583);
nand U10566 (N_10566,N_10346,N_9846);
xor U10567 (N_10567,N_10125,N_9665);
and U10568 (N_10568,N_10022,N_9790);
xor U10569 (N_10569,N_10456,N_10375);
xnor U10570 (N_10570,N_9381,N_9794);
nand U10571 (N_10571,N_10031,N_10466);
xor U10572 (N_10572,N_9111,N_9570);
nand U10573 (N_10573,N_9985,N_10013);
nand U10574 (N_10574,N_9270,N_9298);
and U10575 (N_10575,N_9787,N_10006);
and U10576 (N_10576,N_10263,N_10429);
nor U10577 (N_10577,N_9107,N_9389);
or U10578 (N_10578,N_9051,N_10194);
xor U10579 (N_10579,N_10177,N_9054);
and U10580 (N_10580,N_9542,N_9529);
nor U10581 (N_10581,N_9282,N_9528);
or U10582 (N_10582,N_9567,N_9564);
nor U10583 (N_10583,N_9407,N_9267);
nand U10584 (N_10584,N_10057,N_9067);
nor U10585 (N_10585,N_10124,N_10295);
nand U10586 (N_10586,N_9188,N_9289);
nor U10587 (N_10587,N_10421,N_9718);
or U10588 (N_10588,N_9682,N_9637);
xnor U10589 (N_10589,N_9667,N_9388);
or U10590 (N_10590,N_9242,N_9205);
nand U10591 (N_10591,N_9201,N_9870);
nand U10592 (N_10592,N_9236,N_9024);
nor U10593 (N_10593,N_9322,N_9472);
or U10594 (N_10594,N_10407,N_10333);
and U10595 (N_10595,N_9952,N_9753);
and U10596 (N_10596,N_9854,N_9105);
nand U10597 (N_10597,N_10051,N_10437);
nand U10598 (N_10598,N_9095,N_10327);
or U10599 (N_10599,N_9987,N_9878);
nand U10600 (N_10600,N_10186,N_10184);
and U10601 (N_10601,N_9113,N_9064);
nand U10602 (N_10602,N_10017,N_9304);
nor U10603 (N_10603,N_9786,N_10498);
or U10604 (N_10604,N_9853,N_9083);
and U10605 (N_10605,N_10298,N_10444);
nor U10606 (N_10606,N_9766,N_9191);
nor U10607 (N_10607,N_9998,N_9369);
nor U10608 (N_10608,N_9137,N_9231);
and U10609 (N_10609,N_9924,N_9166);
or U10610 (N_10610,N_10120,N_10198);
nor U10611 (N_10611,N_10291,N_9452);
nor U10612 (N_10612,N_10486,N_9225);
xnor U10613 (N_10613,N_9148,N_10463);
nand U10614 (N_10614,N_9713,N_10310);
or U10615 (N_10615,N_9285,N_9396);
nor U10616 (N_10616,N_9109,N_10092);
or U10617 (N_10617,N_9752,N_9873);
nand U10618 (N_10618,N_9700,N_9275);
nor U10619 (N_10619,N_9807,N_10182);
and U10620 (N_10620,N_10353,N_9781);
or U10621 (N_10621,N_10479,N_9822);
and U10622 (N_10622,N_9088,N_10069);
xnor U10623 (N_10623,N_10361,N_9358);
nand U10624 (N_10624,N_9709,N_10060);
nand U10625 (N_10625,N_9457,N_10382);
and U10626 (N_10626,N_9147,N_9892);
and U10627 (N_10627,N_9200,N_10303);
nor U10628 (N_10628,N_9416,N_9081);
nor U10629 (N_10629,N_10299,N_9256);
xnor U10630 (N_10630,N_9509,N_9538);
nor U10631 (N_10631,N_9848,N_10487);
xor U10632 (N_10632,N_9750,N_10240);
nand U10633 (N_10633,N_9645,N_9664);
nor U10634 (N_10634,N_10330,N_9756);
nand U10635 (N_10635,N_9910,N_9863);
xnor U10636 (N_10636,N_10202,N_9726);
nand U10637 (N_10637,N_9847,N_9784);
nand U10638 (N_10638,N_10205,N_10096);
or U10639 (N_10639,N_9075,N_9581);
nor U10640 (N_10640,N_9675,N_9830);
or U10641 (N_10641,N_10085,N_9424);
nor U10642 (N_10642,N_10484,N_9536);
or U10643 (N_10643,N_10336,N_10317);
or U10644 (N_10644,N_9293,N_10350);
nand U10645 (N_10645,N_9999,N_9535);
xor U10646 (N_10646,N_9356,N_9053);
and U10647 (N_10647,N_10434,N_9643);
nor U10648 (N_10648,N_9876,N_10416);
xor U10649 (N_10649,N_9678,N_9335);
or U10650 (N_10650,N_9996,N_9268);
or U10651 (N_10651,N_9571,N_9340);
nor U10652 (N_10652,N_9809,N_9410);
and U10653 (N_10653,N_10037,N_9520);
or U10654 (N_10654,N_10467,N_9526);
or U10655 (N_10655,N_9888,N_9391);
or U10656 (N_10656,N_9033,N_9648);
and U10657 (N_10657,N_9869,N_9762);
or U10658 (N_10658,N_9865,N_9370);
xor U10659 (N_10659,N_9744,N_9855);
or U10660 (N_10660,N_9441,N_9026);
nand U10661 (N_10661,N_9221,N_9760);
nor U10662 (N_10662,N_9641,N_9723);
and U10663 (N_10663,N_9939,N_9186);
xor U10664 (N_10664,N_9886,N_9361);
nor U10665 (N_10665,N_10253,N_9898);
and U10666 (N_10666,N_9945,N_10329);
nor U10667 (N_10667,N_9946,N_10403);
or U10668 (N_10668,N_10493,N_9650);
nand U10669 (N_10669,N_9208,N_9458);
nand U10670 (N_10670,N_9110,N_9922);
nor U10671 (N_10671,N_9012,N_9896);
or U10672 (N_10672,N_10196,N_9165);
nor U10673 (N_10673,N_9069,N_10173);
nor U10674 (N_10674,N_10084,N_9367);
and U10675 (N_10675,N_10206,N_9004);
nor U10676 (N_10676,N_10204,N_9913);
nor U10677 (N_10677,N_9811,N_9785);
nand U10678 (N_10678,N_9384,N_9019);
nand U10679 (N_10679,N_9280,N_10045);
or U10680 (N_10680,N_9585,N_10388);
nor U10681 (N_10681,N_9131,N_9038);
xor U10682 (N_10682,N_9184,N_9710);
nand U10683 (N_10683,N_10459,N_10034);
and U10684 (N_10684,N_10016,N_9278);
or U10685 (N_10685,N_10080,N_10075);
nor U10686 (N_10686,N_10137,N_9919);
nor U10687 (N_10687,N_9291,N_10344);
nand U10688 (N_10688,N_10119,N_9348);
xor U10689 (N_10689,N_9039,N_9491);
and U10690 (N_10690,N_9938,N_10162);
nand U10691 (N_10691,N_10073,N_10453);
nor U10692 (N_10692,N_9378,N_9239);
and U10693 (N_10693,N_9828,N_9118);
nor U10694 (N_10694,N_10471,N_9479);
nor U10695 (N_10695,N_9730,N_10103);
or U10696 (N_10696,N_10142,N_9731);
nor U10697 (N_10697,N_9951,N_9511);
nor U10698 (N_10698,N_9959,N_9228);
and U10699 (N_10699,N_9102,N_10116);
nor U10700 (N_10700,N_10130,N_10218);
or U10701 (N_10701,N_10391,N_9568);
and U10702 (N_10702,N_9516,N_10366);
nor U10703 (N_10703,N_9634,N_10386);
or U10704 (N_10704,N_9016,N_10050);
nor U10705 (N_10705,N_10258,N_9115);
nor U10706 (N_10706,N_9963,N_9329);
nand U10707 (N_10707,N_10132,N_9185);
xnor U10708 (N_10708,N_9449,N_9606);
nand U10709 (N_10709,N_9383,N_10422);
and U10710 (N_10710,N_9195,N_9465);
nor U10711 (N_10711,N_10113,N_9198);
xnor U10712 (N_10712,N_9988,N_10071);
nand U10713 (N_10713,N_10101,N_9841);
nand U10714 (N_10714,N_9136,N_10308);
nand U10715 (N_10715,N_9591,N_10131);
and U10716 (N_10716,N_10215,N_9049);
or U10717 (N_10717,N_9474,N_9143);
or U10718 (N_10718,N_9513,N_9313);
or U10719 (N_10719,N_9418,N_10449);
nor U10720 (N_10720,N_9360,N_9798);
nor U10721 (N_10721,N_9975,N_9927);
nand U10722 (N_10722,N_9600,N_9577);
nand U10723 (N_10723,N_9464,N_9912);
and U10724 (N_10724,N_9487,N_9852);
nand U10725 (N_10725,N_9932,N_9087);
nor U10726 (N_10726,N_10220,N_9099);
and U10727 (N_10727,N_10067,N_10090);
nand U10728 (N_10728,N_9349,N_10250);
nand U10729 (N_10729,N_9057,N_10123);
nor U10730 (N_10730,N_9034,N_9953);
nand U10731 (N_10731,N_9721,N_10043);
nor U10732 (N_10732,N_9557,N_10094);
xnor U10733 (N_10733,N_10149,N_9793);
and U10734 (N_10734,N_10476,N_9832);
or U10735 (N_10735,N_9379,N_9877);
nor U10736 (N_10736,N_9023,N_10244);
nand U10737 (N_10737,N_9725,N_10225);
nor U10738 (N_10738,N_9192,N_9860);
nand U10739 (N_10739,N_10039,N_9252);
and U10740 (N_10740,N_9341,N_10213);
or U10741 (N_10741,N_9937,N_10193);
nand U10742 (N_10742,N_9394,N_9310);
nor U10743 (N_10743,N_9925,N_9029);
and U10744 (N_10744,N_9202,N_10266);
and U10745 (N_10745,N_9408,N_9651);
nand U10746 (N_10746,N_10431,N_10231);
or U10747 (N_10747,N_9940,N_10134);
or U10748 (N_10748,N_10181,N_9470);
nor U10749 (N_10749,N_9690,N_9505);
nor U10750 (N_10750,N_9164,N_9751);
and U10751 (N_10751,N_10200,N_9554);
nor U10752 (N_10752,N_10325,N_9114);
and U10753 (N_10753,N_10270,N_10259);
nand U10754 (N_10754,N_10188,N_9531);
nand U10755 (N_10755,N_9598,N_9498);
nand U10756 (N_10756,N_9631,N_9778);
or U10757 (N_10757,N_9626,N_9646);
nor U10758 (N_10758,N_9618,N_9838);
and U10759 (N_10759,N_9749,N_10042);
nor U10760 (N_10760,N_9354,N_9001);
or U10761 (N_10761,N_10242,N_10345);
nor U10762 (N_10762,N_9219,N_9303);
or U10763 (N_10763,N_10316,N_9628);
and U10764 (N_10764,N_9810,N_9544);
nand U10765 (N_10765,N_9915,N_9158);
or U10766 (N_10766,N_9814,N_9290);
and U10767 (N_10767,N_10292,N_9180);
and U10768 (N_10768,N_10324,N_9442);
or U10769 (N_10769,N_9005,N_9989);
nor U10770 (N_10770,N_9764,N_9500);
and U10771 (N_10771,N_9868,N_9679);
nor U10772 (N_10772,N_10197,N_9797);
or U10773 (N_10773,N_9783,N_10003);
nand U10774 (N_10774,N_10183,N_9592);
and U10775 (N_10775,N_10271,N_9548);
xor U10776 (N_10776,N_9492,N_9918);
nor U10777 (N_10777,N_10404,N_9302);
or U10778 (N_10778,N_10338,N_9041);
nand U10779 (N_10779,N_9903,N_10396);
and U10780 (N_10780,N_9362,N_9139);
or U10781 (N_10781,N_9171,N_9234);
or U10782 (N_10782,N_9385,N_9639);
or U10783 (N_10783,N_9803,N_10102);
nand U10784 (N_10784,N_10157,N_9417);
nor U10785 (N_10785,N_9050,N_9132);
nor U10786 (N_10786,N_9485,N_10390);
xor U10787 (N_10787,N_9991,N_9776);
nor U10788 (N_10788,N_10251,N_9124);
or U10789 (N_10789,N_9446,N_9572);
and U10790 (N_10790,N_9672,N_9357);
or U10791 (N_10791,N_9043,N_9758);
or U10792 (N_10792,N_9642,N_9140);
nor U10793 (N_10793,N_10163,N_9328);
and U10794 (N_10794,N_10011,N_9539);
nand U10795 (N_10795,N_9711,N_10237);
nor U10796 (N_10796,N_9748,N_9459);
and U10797 (N_10797,N_9061,N_10236);
or U10798 (N_10798,N_10428,N_9902);
or U10799 (N_10799,N_9871,N_9414);
xor U10800 (N_10800,N_9401,N_9415);
nor U10801 (N_10801,N_9587,N_9507);
nor U10802 (N_10802,N_10339,N_10072);
or U10803 (N_10803,N_9443,N_9524);
and U10804 (N_10804,N_9821,N_9177);
and U10805 (N_10805,N_10461,N_10021);
nor U10806 (N_10806,N_10277,N_9036);
nor U10807 (N_10807,N_9541,N_9018);
nor U10808 (N_10808,N_9220,N_9856);
nor U10809 (N_10809,N_10469,N_9684);
or U10810 (N_10810,N_9022,N_9887);
and U10811 (N_10811,N_10141,N_9556);
or U10812 (N_10812,N_9248,N_9325);
or U10813 (N_10813,N_9494,N_9506);
nand U10814 (N_10814,N_9695,N_9704);
and U10815 (N_10815,N_10383,N_10246);
nor U10816 (N_10816,N_10414,N_9673);
nand U10817 (N_10817,N_10384,N_9866);
and U10818 (N_10818,N_9279,N_9233);
or U10819 (N_10819,N_10447,N_9060);
nand U10820 (N_10820,N_9392,N_9295);
nand U10821 (N_10821,N_9677,N_9272);
or U10822 (N_10822,N_10076,N_9190);
nand U10823 (N_10823,N_10309,N_10285);
and U10824 (N_10824,N_9331,N_9499);
and U10825 (N_10825,N_10114,N_9826);
nor U10826 (N_10826,N_10281,N_9966);
xnor U10827 (N_10827,N_9405,N_9747);
nand U10828 (N_10828,N_10401,N_9112);
nand U10829 (N_10829,N_9961,N_10235);
or U10830 (N_10830,N_9983,N_9259);
nand U10831 (N_10831,N_9210,N_10473);
or U10832 (N_10832,N_9142,N_9837);
xor U10833 (N_10833,N_10038,N_9537);
or U10834 (N_10834,N_9696,N_9635);
nor U10835 (N_10835,N_9624,N_9194);
nand U10836 (N_10836,N_9092,N_9817);
nor U10837 (N_10837,N_10274,N_9880);
and U10838 (N_10838,N_10106,N_9400);
or U10839 (N_10839,N_10441,N_9454);
and U10840 (N_10840,N_9128,N_9373);
nand U10841 (N_10841,N_9578,N_9438);
or U10842 (N_10842,N_9834,N_9074);
nand U10843 (N_10843,N_9347,N_10364);
or U10844 (N_10844,N_10458,N_9674);
or U10845 (N_10845,N_9420,N_9573);
nor U10846 (N_10846,N_10059,N_9742);
or U10847 (N_10847,N_9497,N_10257);
or U10848 (N_10848,N_9920,N_10323);
and U10849 (N_10849,N_10100,N_10082);
or U10850 (N_10850,N_9032,N_9174);
or U10851 (N_10851,N_10430,N_10413);
or U10852 (N_10852,N_9286,N_10152);
and U10853 (N_10853,N_9653,N_10439);
nand U10854 (N_10854,N_10097,N_9839);
and U10855 (N_10855,N_10288,N_9345);
nor U10856 (N_10856,N_10111,N_10239);
nor U10857 (N_10857,N_9517,N_10049);
nor U10858 (N_10858,N_9859,N_9525);
xnor U10859 (N_10859,N_9596,N_9398);
or U10860 (N_10860,N_9720,N_9167);
nor U10861 (N_10861,N_9668,N_9897);
and U10862 (N_10862,N_9563,N_10191);
nand U10863 (N_10863,N_9163,N_10047);
xnor U10864 (N_10864,N_9144,N_9566);
nand U10865 (N_10865,N_9580,N_9299);
xnor U10866 (N_10866,N_10481,N_10169);
nand U10867 (N_10867,N_10424,N_9037);
nor U10868 (N_10868,N_10008,N_9843);
nor U10869 (N_10869,N_9546,N_9217);
and U10870 (N_10870,N_9477,N_9436);
and U10871 (N_10871,N_10372,N_9906);
or U10872 (N_10872,N_10450,N_10457);
or U10873 (N_10873,N_9768,N_9805);
nand U10874 (N_10874,N_9676,N_9736);
nor U10875 (N_10875,N_9402,N_9215);
and U10876 (N_10876,N_10061,N_10305);
nand U10877 (N_10877,N_10275,N_9595);
nand U10878 (N_10878,N_9224,N_10472);
and U10879 (N_10879,N_9104,N_9488);
and U10880 (N_10880,N_10255,N_10495);
nor U10881 (N_10881,N_9972,N_9404);
or U10882 (N_10882,N_9948,N_10219);
and U10883 (N_10883,N_9035,N_9343);
nor U10884 (N_10884,N_9599,N_9250);
and U10885 (N_10885,N_10440,N_9895);
or U10886 (N_10886,N_10393,N_9597);
nand U10887 (N_10887,N_9882,N_9617);
nand U10888 (N_10888,N_9956,N_10454);
or U10889 (N_10889,N_9376,N_9657);
and U10890 (N_10890,N_9604,N_10083);
and U10891 (N_10891,N_9135,N_9375);
or U10892 (N_10892,N_9371,N_9514);
or U10893 (N_10893,N_9350,N_9992);
nand U10894 (N_10894,N_9117,N_10341);
or U10895 (N_10895,N_9152,N_10112);
nand U10896 (N_10896,N_9519,N_9281);
nand U10897 (N_10897,N_10286,N_9779);
and U10898 (N_10898,N_10252,N_9691);
nor U10899 (N_10899,N_9656,N_10207);
or U10900 (N_10900,N_10452,N_10234);
nand U10901 (N_10901,N_9755,N_9745);
and U10902 (N_10902,N_10348,N_9079);
or U10903 (N_10903,N_9782,N_10358);
nand U10904 (N_10904,N_10041,N_9072);
nor U10905 (N_10905,N_10280,N_10066);
or U10906 (N_10906,N_9253,N_9045);
nor U10907 (N_10907,N_10175,N_9739);
nand U10908 (N_10908,N_9048,N_9501);
and U10909 (N_10909,N_9346,N_9512);
and U10910 (N_10910,N_9411,N_10283);
xnor U10911 (N_10911,N_9271,N_9263);
nor U10912 (N_10912,N_10232,N_9719);
or U10913 (N_10913,N_9521,N_9489);
and U10914 (N_10914,N_9767,N_9387);
nand U10915 (N_10915,N_9965,N_9448);
and U10916 (N_10916,N_10012,N_9316);
nor U10917 (N_10917,N_9247,N_9052);
nand U10918 (N_10918,N_10296,N_10068);
nor U10919 (N_10919,N_9780,N_9771);
and U10920 (N_10920,N_9978,N_9495);
and U10921 (N_10921,N_9101,N_9671);
or U10922 (N_10922,N_10004,N_10368);
nand U10923 (N_10923,N_10294,N_9881);
and U10924 (N_10924,N_9160,N_10322);
nor U10925 (N_10925,N_9941,N_10489);
nor U10926 (N_10926,N_10208,N_9942);
and U10927 (N_10927,N_9342,N_10492);
or U10928 (N_10928,N_9911,N_9307);
and U10929 (N_10929,N_10312,N_9614);
nand U10930 (N_10930,N_9947,N_10381);
nor U10931 (N_10931,N_9984,N_9108);
xnor U10932 (N_10932,N_10035,N_9040);
and U10933 (N_10933,N_9423,N_10397);
nor U10934 (N_10934,N_9842,N_9586);
nand U10935 (N_10935,N_9703,N_9334);
and U10936 (N_10936,N_9769,N_10435);
and U10937 (N_10937,N_10482,N_9475);
nand U10938 (N_10938,N_9850,N_9046);
and U10939 (N_10939,N_9337,N_9801);
nand U10940 (N_10940,N_9312,N_10126);
nor U10941 (N_10941,N_10265,N_10010);
and U10942 (N_10942,N_10150,N_9025);
nand U10943 (N_10943,N_10478,N_9120);
and U10944 (N_10944,N_9603,N_10377);
xnor U10945 (N_10945,N_9727,N_9435);
nor U10946 (N_10946,N_9245,N_9047);
or U10947 (N_10947,N_9808,N_10201);
nor U10948 (N_10948,N_10032,N_9508);
and U10949 (N_10949,N_9788,N_9123);
and U10950 (N_10950,N_9044,N_9738);
and U10951 (N_10951,N_9235,N_10107);
nand U10952 (N_10952,N_9958,N_10272);
nand U10953 (N_10953,N_9610,N_9181);
nor U10954 (N_10954,N_9071,N_9461);
nor U10955 (N_10955,N_10446,N_10089);
or U10956 (N_10956,N_9804,N_9241);
and U10957 (N_10957,N_10018,N_9000);
nor U10958 (N_10958,N_9861,N_9659);
nand U10959 (N_10959,N_10356,N_10343);
or U10960 (N_10960,N_9020,N_9698);
xnor U10961 (N_10961,N_9240,N_9169);
nand U10962 (N_10962,N_10445,N_9269);
xnor U10963 (N_10963,N_10129,N_10211);
and U10964 (N_10964,N_9106,N_9266);
nor U10965 (N_10965,N_9309,N_9662);
and U10966 (N_10966,N_10154,N_10405);
nand U10967 (N_10967,N_10331,N_10189);
or U10968 (N_10968,N_9757,N_9504);
nand U10969 (N_10969,N_9827,N_9276);
nor U10970 (N_10970,N_9066,N_10040);
or U10971 (N_10971,N_9562,N_10195);
or U10972 (N_10972,N_10477,N_10118);
or U10973 (N_10973,N_9243,N_9615);
and U10974 (N_10974,N_9390,N_9616);
nand U10975 (N_10975,N_9789,N_10238);
or U10976 (N_10976,N_9715,N_9928);
and U10977 (N_10977,N_10158,N_9950);
xnor U10978 (N_10978,N_10374,N_9440);
nand U10979 (N_10979,N_10389,N_9365);
or U10980 (N_10980,N_9260,N_10245);
nand U10981 (N_10981,N_10001,N_10307);
nand U10982 (N_10982,N_10199,N_10367);
or U10983 (N_10983,N_9478,N_9182);
nor U10984 (N_10984,N_10053,N_9254);
nand U10985 (N_10985,N_10095,N_9437);
nand U10986 (N_10986,N_9737,N_10321);
and U10987 (N_10987,N_10046,N_9944);
xor U10988 (N_10988,N_9353,N_9559);
nor U10989 (N_10989,N_9481,N_9823);
nand U10990 (N_10990,N_9264,N_9661);
xnor U10991 (N_10991,N_9249,N_9393);
nor U10992 (N_10992,N_9339,N_9352);
xor U10993 (N_10993,N_9323,N_9908);
and U10994 (N_10994,N_9133,N_10369);
or U10995 (N_10995,N_9921,N_10319);
xor U10996 (N_10996,N_9486,N_9824);
or U10997 (N_10997,N_10464,N_10499);
nor U10998 (N_10998,N_9970,N_10256);
nor U10999 (N_10999,N_10474,N_9179);
xnor U11000 (N_11000,N_9319,N_9763);
and U11001 (N_11001,N_9430,N_9874);
nor U11002 (N_11002,N_9355,N_9403);
and U11003 (N_11003,N_9885,N_10027);
nor U11004 (N_11004,N_10115,N_10128);
or U11005 (N_11005,N_9777,N_9063);
and U11006 (N_11006,N_9916,N_9466);
or U11007 (N_11007,N_10349,N_9973);
nor U11008 (N_11008,N_9607,N_9216);
nor U11009 (N_11009,N_9125,N_9294);
nand U11010 (N_11010,N_9223,N_10494);
nor U11011 (N_11011,N_9122,N_9031);
or U11012 (N_11012,N_9157,N_9451);
and U11013 (N_11013,N_9705,N_9483);
nand U11014 (N_11014,N_10337,N_9608);
nor U11015 (N_11015,N_10233,N_9336);
and U11016 (N_11016,N_9476,N_9138);
nand U11017 (N_11017,N_10451,N_10326);
nor U11018 (N_11018,N_10024,N_9620);
xnor U11019 (N_11019,N_10332,N_9735);
and U11020 (N_11020,N_9532,N_9251);
nand U11021 (N_11021,N_9933,N_10026);
nor U11022 (N_11022,N_9706,N_9625);
and U11023 (N_11023,N_9707,N_10171);
nor U11024 (N_11024,N_9708,N_9288);
xor U11025 (N_11025,N_9318,N_9320);
xor U11026 (N_11026,N_9936,N_9426);
nand U11027 (N_11027,N_10168,N_9317);
or U11028 (N_11028,N_10497,N_10365);
nor U11029 (N_11029,N_10230,N_10300);
nand U11030 (N_11030,N_10273,N_10302);
and U11031 (N_11031,N_9652,N_9287);
or U11032 (N_11032,N_9589,N_9929);
nor U11033 (N_11033,N_9518,N_9008);
nor U11034 (N_11034,N_10143,N_9444);
or U11035 (N_11035,N_9746,N_10438);
and U11036 (N_11036,N_9611,N_9197);
and U11037 (N_11037,N_9582,N_10019);
nand U11038 (N_11038,N_10320,N_9701);
nor U11039 (N_11039,N_10216,N_9619);
and U11040 (N_11040,N_10293,N_9829);
nand U11041 (N_11041,N_9986,N_9522);
xnor U11042 (N_11042,N_9068,N_9630);
nor U11043 (N_11043,N_9670,N_9574);
nor U11044 (N_11044,N_9199,N_10108);
or U11045 (N_11045,N_9351,N_9292);
xnor U11046 (N_11046,N_10468,N_9773);
xor U11047 (N_11047,N_9327,N_9774);
and U11048 (N_11048,N_10023,N_10385);
and U11049 (N_11049,N_10015,N_10264);
nor U11050 (N_11050,N_10410,N_9419);
nand U11051 (N_11051,N_9433,N_9058);
nand U11052 (N_11052,N_9070,N_10311);
or U11053 (N_11053,N_9995,N_9890);
and U11054 (N_11054,N_10284,N_9980);
nand U11055 (N_11055,N_10491,N_10415);
nor U11056 (N_11056,N_10432,N_10185);
and U11057 (N_11057,N_9716,N_10412);
or U11058 (N_11058,N_9368,N_9196);
or U11059 (N_11059,N_10161,N_9229);
and U11060 (N_11060,N_9979,N_9802);
nor U11061 (N_11061,N_9982,N_9344);
nor U11062 (N_11062,N_9366,N_9078);
xor U11063 (N_11063,N_9427,N_10399);
xor U11064 (N_11064,N_9153,N_10223);
or U11065 (N_11065,N_9332,N_9761);
xor U11066 (N_11066,N_9155,N_9314);
xor U11067 (N_11067,N_9728,N_9644);
nand U11068 (N_11068,N_9840,N_9116);
nor U11069 (N_11069,N_9934,N_9692);
and U11070 (N_11070,N_9480,N_9697);
nor U11071 (N_11071,N_9311,N_9627);
or U11072 (N_11072,N_10261,N_10087);
xor U11073 (N_11073,N_10151,N_9689);
nand U11074 (N_11074,N_9096,N_10370);
nand U11075 (N_11075,N_10334,N_9014);
or U11076 (N_11076,N_10267,N_10423);
or U11077 (N_11077,N_9413,N_9660);
and U11078 (N_11078,N_9330,N_9178);
and U11079 (N_11079,N_10387,N_9257);
nor U11080 (N_11080,N_9421,N_9694);
and U11081 (N_11081,N_9867,N_9121);
nor U11082 (N_11082,N_9258,N_9006);
nand U11083 (N_11083,N_9002,N_9584);
xor U11084 (N_11084,N_9862,N_9923);
nand U11085 (N_11085,N_9954,N_9090);
xnor U11086 (N_11086,N_9712,N_9382);
nand U11087 (N_11087,N_9796,N_9207);
and U11088 (N_11088,N_9364,N_10062);
or U11089 (N_11089,N_10470,N_9232);
or U11090 (N_11090,N_10340,N_9569);
nor U11091 (N_11091,N_9702,N_9326);
or U11092 (N_11092,N_9594,N_9432);
nand U11093 (N_11093,N_9262,N_10088);
or U11094 (N_11094,N_9858,N_9891);
xnor U11095 (N_11095,N_9655,N_9100);
nand U11096 (N_11096,N_9576,N_9409);
or U11097 (N_11097,N_9149,N_9453);
nor U11098 (N_11098,N_9901,N_9636);
nand U11099 (N_11099,N_9605,N_9183);
or U11100 (N_11100,N_9905,N_9089);
nand U11101 (N_11101,N_9097,N_10105);
nand U11102 (N_11102,N_9386,N_9170);
or U11103 (N_11103,N_10170,N_9175);
nand U11104 (N_11104,N_9543,N_9549);
or U11105 (N_11105,N_9926,N_10362);
and U11106 (N_11106,N_9206,N_9669);
nor U11107 (N_11107,N_10419,N_10483);
or U11108 (N_11108,N_9428,N_9103);
or U11109 (N_11109,N_10433,N_10167);
nor U11110 (N_11110,N_9819,N_9990);
xnor U11111 (N_11111,N_9324,N_9315);
nor U11112 (N_11112,N_10443,N_10214);
and U11113 (N_11113,N_9425,N_9150);
or U11114 (N_11114,N_9816,N_9082);
and U11115 (N_11115,N_10287,N_10379);
or U11116 (N_11116,N_9844,N_10166);
and U11117 (N_11117,N_10176,N_9468);
and U11118 (N_11118,N_10425,N_9203);
xnor U11119 (N_11119,N_9094,N_9176);
or U11120 (N_11120,N_10360,N_10465);
and U11121 (N_11121,N_10402,N_10347);
nor U11122 (N_11122,N_10406,N_10044);
nand U11123 (N_11123,N_10276,N_9754);
nand U11124 (N_11124,N_9772,N_10063);
and U11125 (N_11125,N_10376,N_9214);
nor U11126 (N_11126,N_9056,N_9935);
or U11127 (N_11127,N_10192,N_10033);
nand U11128 (N_11128,N_9482,N_9510);
nor U11129 (N_11129,N_9146,N_10426);
nand U11130 (N_11130,N_10164,N_10005);
nor U11131 (N_11131,N_9724,N_9931);
and U11132 (N_11132,N_9338,N_10146);
and U11133 (N_11133,N_9484,N_9957);
or U11134 (N_11134,N_9899,N_9222);
and U11135 (N_11135,N_9812,N_9015);
nand U11136 (N_11136,N_9993,N_10160);
or U11137 (N_11137,N_9741,N_10064);
nand U11138 (N_11138,N_9770,N_10352);
xnor U11139 (N_11139,N_10395,N_10480);
nor U11140 (N_11140,N_10122,N_9306);
nor U11141 (N_11141,N_10297,N_9173);
or U11142 (N_11142,N_10000,N_9977);
and U11143 (N_11143,N_9884,N_9997);
or U11144 (N_11144,N_9080,N_9490);
xor U11145 (N_11145,N_9685,N_10190);
nand U11146 (N_11146,N_9799,N_10359);
nor U11147 (N_11147,N_10490,N_9967);
nor U11148 (N_11148,N_9212,N_9460);
or U11149 (N_11149,N_9552,N_9833);
nand U11150 (N_11150,N_9084,N_9226);
and U11151 (N_11151,N_10156,N_10136);
nand U11152 (N_11152,N_9845,N_9238);
nor U11153 (N_11153,N_9447,N_9613);
nand U11154 (N_11154,N_9471,N_9647);
nand U11155 (N_11155,N_9162,N_10174);
and U11156 (N_11156,N_9129,N_10002);
and U11157 (N_11157,N_9077,N_9649);
nor U11158 (N_11158,N_10140,N_9227);
nor U11159 (N_11159,N_10153,N_9714);
or U11160 (N_11160,N_9623,N_9065);
nor U11161 (N_11161,N_9021,N_9969);
or U11162 (N_11162,N_9273,N_10241);
nor U11163 (N_11163,N_10248,N_9732);
nand U11164 (N_11164,N_9686,N_10278);
or U11165 (N_11165,N_9831,N_9976);
nand U11166 (N_11166,N_9093,N_10209);
and U11167 (N_11167,N_10411,N_10099);
or U11168 (N_11168,N_9261,N_9633);
nor U11169 (N_11169,N_10055,N_9028);
nor U11170 (N_11170,N_10187,N_9968);
or U11171 (N_11171,N_9359,N_9496);
nor U11172 (N_11172,N_10355,N_9964);
nor U11173 (N_11173,N_9333,N_9640);
or U11174 (N_11174,N_10335,N_9462);
nor U11175 (N_11175,N_10081,N_9681);
nand U11176 (N_11176,N_10117,N_10165);
xor U11177 (N_11177,N_10148,N_9374);
and U11178 (N_11178,N_10020,N_9073);
or U11179 (N_11179,N_9560,N_9815);
xor U11180 (N_11180,N_10315,N_10074);
nor U11181 (N_11181,N_10290,N_10109);
or U11182 (N_11182,N_10417,N_9399);
or U11183 (N_11183,N_10079,N_9189);
and U11184 (N_11184,N_10054,N_10155);
nor U11185 (N_11185,N_10221,N_10226);
or U11186 (N_11186,N_10048,N_9791);
or U11187 (N_11187,N_10398,N_9467);
nand U11188 (N_11188,N_9835,N_9027);
xor U11189 (N_11189,N_9237,N_9693);
xnor U11190 (N_11190,N_10269,N_9218);
xor U11191 (N_11191,N_10135,N_9806);
xnor U11192 (N_11192,N_9445,N_9456);
nand U11193 (N_11193,N_9013,N_9654);
and U11194 (N_11194,N_10357,N_9244);
nor U11195 (N_11195,N_9055,N_10210);
nor U11196 (N_11196,N_10409,N_10212);
nand U11197 (N_11197,N_9503,N_9666);
nor U11198 (N_11198,N_9422,N_10028);
nand U11199 (N_11199,N_10014,N_10159);
nor U11200 (N_11200,N_10056,N_10139);
nand U11201 (N_11201,N_9515,N_9960);
nand U11202 (N_11202,N_9575,N_9974);
nand U11203 (N_11203,N_9429,N_9743);
nor U11204 (N_11204,N_9875,N_9699);
nor U11205 (N_11205,N_9687,N_9187);
and U11206 (N_11206,N_10224,N_9820);
and U11207 (N_11207,N_9558,N_10394);
and U11208 (N_11208,N_9879,N_9372);
nor U11209 (N_11209,N_10378,N_10110);
nand U11210 (N_11210,N_10448,N_10007);
nor U11211 (N_11211,N_9930,N_10145);
or U11212 (N_11212,N_9872,N_10127);
nor U11213 (N_11213,N_9545,N_9740);
and U11214 (N_11214,N_10373,N_9119);
xnor U11215 (N_11215,N_9792,N_9949);
nand U11216 (N_11216,N_9523,N_9857);
and U11217 (N_11217,N_9204,N_10172);
and U11218 (N_11218,N_10455,N_9800);
nand U11219 (N_11219,N_9733,N_9909);
nor U11220 (N_11220,N_9775,N_9010);
and U11221 (N_11221,N_9688,N_10254);
xor U11222 (N_11222,N_9091,N_10260);
or U11223 (N_11223,N_9683,N_9981);
nand U11224 (N_11224,N_10262,N_9193);
nand U11225 (N_11225,N_9159,N_9962);
and U11226 (N_11226,N_9439,N_10091);
or U11227 (N_11227,N_10268,N_9894);
nor U11228 (N_11228,N_9609,N_9473);
nor U11229 (N_11229,N_9098,N_10030);
xor U11230 (N_11230,N_9602,N_9283);
nand U11231 (N_11231,N_9527,N_9363);
nand U11232 (N_11232,N_9126,N_10313);
nor U11233 (N_11233,N_10289,N_10179);
and U11234 (N_11234,N_9305,N_9308);
or U11235 (N_11235,N_10279,N_9795);
or U11236 (N_11236,N_9638,N_9172);
xor U11237 (N_11237,N_10025,N_9907);
nand U11238 (N_11238,N_9622,N_9530);
nor U11239 (N_11239,N_9156,N_9658);
nor U11240 (N_11240,N_9734,N_9130);
and U11241 (N_11241,N_9663,N_10420);
nor U11242 (N_11242,N_9127,N_9621);
and U11243 (N_11243,N_9297,N_10243);
nand U11244 (N_11244,N_10496,N_9246);
nand U11245 (N_11245,N_9765,N_9588);
nor U11246 (N_11246,N_10065,N_9017);
nor U11247 (N_11247,N_9540,N_9955);
nor U11248 (N_11248,N_10227,N_10460);
nor U11249 (N_11249,N_9141,N_9450);
nand U11250 (N_11250,N_10288,N_10206);
xnor U11251 (N_11251,N_10321,N_9067);
and U11252 (N_11252,N_9343,N_10287);
and U11253 (N_11253,N_10443,N_9300);
or U11254 (N_11254,N_9508,N_9312);
or U11255 (N_11255,N_10397,N_9662);
nand U11256 (N_11256,N_9302,N_9590);
nor U11257 (N_11257,N_9870,N_9719);
nor U11258 (N_11258,N_9163,N_10433);
nor U11259 (N_11259,N_10391,N_9607);
nor U11260 (N_11260,N_9339,N_10231);
or U11261 (N_11261,N_9965,N_9128);
and U11262 (N_11262,N_10156,N_9770);
and U11263 (N_11263,N_9562,N_9872);
nand U11264 (N_11264,N_9350,N_10219);
or U11265 (N_11265,N_9646,N_9890);
nor U11266 (N_11266,N_9360,N_9217);
xor U11267 (N_11267,N_9653,N_9915);
nand U11268 (N_11268,N_10020,N_10093);
nor U11269 (N_11269,N_9047,N_9169);
or U11270 (N_11270,N_9997,N_10270);
xnor U11271 (N_11271,N_9149,N_9189);
xor U11272 (N_11272,N_10332,N_10401);
or U11273 (N_11273,N_10181,N_9215);
or U11274 (N_11274,N_9033,N_10346);
and U11275 (N_11275,N_10348,N_9868);
or U11276 (N_11276,N_9228,N_9847);
and U11277 (N_11277,N_9461,N_9206);
xor U11278 (N_11278,N_10360,N_9684);
nand U11279 (N_11279,N_10037,N_9257);
or U11280 (N_11280,N_9826,N_10293);
nand U11281 (N_11281,N_10372,N_9696);
nor U11282 (N_11282,N_9797,N_9463);
and U11283 (N_11283,N_9610,N_10368);
and U11284 (N_11284,N_9500,N_10242);
nor U11285 (N_11285,N_9486,N_9519);
and U11286 (N_11286,N_9501,N_10281);
nand U11287 (N_11287,N_10053,N_10121);
or U11288 (N_11288,N_10184,N_9458);
nand U11289 (N_11289,N_9316,N_10040);
and U11290 (N_11290,N_9343,N_10110);
and U11291 (N_11291,N_10344,N_10482);
or U11292 (N_11292,N_9322,N_10086);
or U11293 (N_11293,N_9185,N_9572);
nand U11294 (N_11294,N_9427,N_9824);
or U11295 (N_11295,N_9887,N_9720);
nand U11296 (N_11296,N_9883,N_10056);
nand U11297 (N_11297,N_9845,N_9789);
xnor U11298 (N_11298,N_9745,N_9065);
nand U11299 (N_11299,N_9813,N_9884);
and U11300 (N_11300,N_9613,N_9820);
xor U11301 (N_11301,N_10124,N_9811);
and U11302 (N_11302,N_9085,N_10117);
nand U11303 (N_11303,N_9395,N_9611);
and U11304 (N_11304,N_9081,N_9359);
nor U11305 (N_11305,N_9330,N_9593);
xor U11306 (N_11306,N_9069,N_9366);
or U11307 (N_11307,N_9990,N_9165);
and U11308 (N_11308,N_9461,N_9396);
and U11309 (N_11309,N_9053,N_9823);
nand U11310 (N_11310,N_9346,N_9836);
or U11311 (N_11311,N_9780,N_9532);
and U11312 (N_11312,N_9012,N_10075);
xnor U11313 (N_11313,N_10081,N_10373);
nor U11314 (N_11314,N_10059,N_9335);
xnor U11315 (N_11315,N_9896,N_10192);
nor U11316 (N_11316,N_10496,N_9688);
nor U11317 (N_11317,N_9869,N_10215);
nand U11318 (N_11318,N_9577,N_9199);
nor U11319 (N_11319,N_9149,N_9839);
nand U11320 (N_11320,N_10069,N_10080);
xor U11321 (N_11321,N_9493,N_9265);
or U11322 (N_11322,N_10181,N_9171);
xor U11323 (N_11323,N_9395,N_9092);
nand U11324 (N_11324,N_9367,N_9057);
nand U11325 (N_11325,N_10075,N_9376);
or U11326 (N_11326,N_10495,N_9056);
nor U11327 (N_11327,N_9791,N_10071);
and U11328 (N_11328,N_10071,N_9565);
nand U11329 (N_11329,N_10401,N_9949);
nand U11330 (N_11330,N_9813,N_10268);
xor U11331 (N_11331,N_9763,N_9728);
nand U11332 (N_11332,N_10179,N_9916);
nand U11333 (N_11333,N_9422,N_10094);
nor U11334 (N_11334,N_10184,N_10132);
or U11335 (N_11335,N_9581,N_9182);
xnor U11336 (N_11336,N_9326,N_9900);
or U11337 (N_11337,N_9332,N_9082);
xor U11338 (N_11338,N_9799,N_9751);
nand U11339 (N_11339,N_9451,N_9717);
nand U11340 (N_11340,N_9181,N_10011);
nor U11341 (N_11341,N_9499,N_9786);
or U11342 (N_11342,N_9286,N_9342);
xor U11343 (N_11343,N_9467,N_10060);
nor U11344 (N_11344,N_9727,N_9805);
nand U11345 (N_11345,N_10069,N_9866);
and U11346 (N_11346,N_9719,N_9161);
and U11347 (N_11347,N_10294,N_10242);
or U11348 (N_11348,N_9637,N_9500);
nand U11349 (N_11349,N_9724,N_9677);
xor U11350 (N_11350,N_10018,N_9813);
or U11351 (N_11351,N_9328,N_9394);
and U11352 (N_11352,N_9376,N_9024);
and U11353 (N_11353,N_9852,N_10271);
or U11354 (N_11354,N_9671,N_9798);
nor U11355 (N_11355,N_9243,N_9658);
nand U11356 (N_11356,N_9546,N_9361);
nor U11357 (N_11357,N_10201,N_9110);
nor U11358 (N_11358,N_10223,N_9943);
nor U11359 (N_11359,N_10332,N_9821);
and U11360 (N_11360,N_9555,N_9955);
nor U11361 (N_11361,N_10271,N_9344);
nor U11362 (N_11362,N_10038,N_10115);
nor U11363 (N_11363,N_9601,N_10433);
nor U11364 (N_11364,N_10414,N_9406);
nor U11365 (N_11365,N_10079,N_9959);
and U11366 (N_11366,N_9486,N_10003);
and U11367 (N_11367,N_9029,N_9601);
nand U11368 (N_11368,N_9212,N_9832);
and U11369 (N_11369,N_10285,N_10459);
xnor U11370 (N_11370,N_9422,N_9828);
nor U11371 (N_11371,N_9466,N_9392);
xnor U11372 (N_11372,N_10322,N_10429);
and U11373 (N_11373,N_10089,N_9898);
and U11374 (N_11374,N_9797,N_9047);
nand U11375 (N_11375,N_9873,N_9739);
nand U11376 (N_11376,N_10361,N_10200);
or U11377 (N_11377,N_10378,N_9980);
nor U11378 (N_11378,N_9287,N_9550);
nor U11379 (N_11379,N_9345,N_9915);
nand U11380 (N_11380,N_9944,N_10325);
and U11381 (N_11381,N_9488,N_10241);
xnor U11382 (N_11382,N_9905,N_9186);
or U11383 (N_11383,N_10223,N_9783);
nand U11384 (N_11384,N_9214,N_9361);
xnor U11385 (N_11385,N_10382,N_10478);
nor U11386 (N_11386,N_9363,N_9161);
nor U11387 (N_11387,N_9680,N_9473);
nand U11388 (N_11388,N_10202,N_10249);
nor U11389 (N_11389,N_9820,N_10403);
nor U11390 (N_11390,N_9010,N_9318);
nand U11391 (N_11391,N_9930,N_10154);
xnor U11392 (N_11392,N_9454,N_9647);
and U11393 (N_11393,N_10217,N_10079);
xnor U11394 (N_11394,N_9107,N_9559);
and U11395 (N_11395,N_10101,N_9505);
nand U11396 (N_11396,N_9471,N_9482);
nand U11397 (N_11397,N_10058,N_9972);
nand U11398 (N_11398,N_10013,N_10006);
nor U11399 (N_11399,N_9286,N_9326);
nand U11400 (N_11400,N_9526,N_9850);
or U11401 (N_11401,N_9112,N_9470);
nor U11402 (N_11402,N_9778,N_9395);
nor U11403 (N_11403,N_10008,N_9694);
nor U11404 (N_11404,N_9448,N_10231);
nand U11405 (N_11405,N_9105,N_9448);
nor U11406 (N_11406,N_10170,N_9988);
nand U11407 (N_11407,N_10164,N_9807);
and U11408 (N_11408,N_10118,N_9038);
xor U11409 (N_11409,N_10460,N_10297);
and U11410 (N_11410,N_10418,N_10363);
nand U11411 (N_11411,N_9883,N_9986);
or U11412 (N_11412,N_10352,N_9902);
or U11413 (N_11413,N_9775,N_9294);
nand U11414 (N_11414,N_10168,N_10204);
nor U11415 (N_11415,N_9979,N_9599);
or U11416 (N_11416,N_10239,N_10194);
nor U11417 (N_11417,N_9397,N_10229);
nor U11418 (N_11418,N_10461,N_9412);
and U11419 (N_11419,N_10198,N_9661);
nor U11420 (N_11420,N_9676,N_10382);
xnor U11421 (N_11421,N_9939,N_9259);
nor U11422 (N_11422,N_10126,N_9447);
and U11423 (N_11423,N_9688,N_10361);
or U11424 (N_11424,N_10448,N_9215);
nand U11425 (N_11425,N_9532,N_9596);
and U11426 (N_11426,N_9804,N_9696);
or U11427 (N_11427,N_9448,N_9250);
and U11428 (N_11428,N_9758,N_9807);
or U11429 (N_11429,N_9995,N_9882);
xor U11430 (N_11430,N_9297,N_9248);
or U11431 (N_11431,N_9206,N_9955);
or U11432 (N_11432,N_9322,N_9143);
or U11433 (N_11433,N_9605,N_9994);
and U11434 (N_11434,N_9989,N_9035);
and U11435 (N_11435,N_9482,N_9460);
and U11436 (N_11436,N_10144,N_9607);
nand U11437 (N_11437,N_9822,N_10088);
nand U11438 (N_11438,N_9906,N_9362);
nand U11439 (N_11439,N_9509,N_9475);
and U11440 (N_11440,N_9488,N_9050);
and U11441 (N_11441,N_10325,N_10319);
and U11442 (N_11442,N_9847,N_9017);
or U11443 (N_11443,N_9131,N_10002);
nand U11444 (N_11444,N_9253,N_9939);
nand U11445 (N_11445,N_9654,N_9336);
xnor U11446 (N_11446,N_10172,N_10215);
or U11447 (N_11447,N_9126,N_10103);
nor U11448 (N_11448,N_10216,N_10076);
xnor U11449 (N_11449,N_9293,N_9135);
or U11450 (N_11450,N_9349,N_9361);
xnor U11451 (N_11451,N_9386,N_10373);
nand U11452 (N_11452,N_10067,N_10295);
or U11453 (N_11453,N_9056,N_9075);
nand U11454 (N_11454,N_9540,N_9811);
nor U11455 (N_11455,N_10370,N_9841);
or U11456 (N_11456,N_9031,N_10335);
nor U11457 (N_11457,N_9086,N_9831);
or U11458 (N_11458,N_9643,N_9468);
or U11459 (N_11459,N_9840,N_10327);
and U11460 (N_11460,N_9106,N_10001);
nor U11461 (N_11461,N_9552,N_9619);
or U11462 (N_11462,N_9457,N_9618);
or U11463 (N_11463,N_9637,N_9703);
nor U11464 (N_11464,N_9433,N_9679);
nand U11465 (N_11465,N_9455,N_9185);
nand U11466 (N_11466,N_9383,N_9187);
nor U11467 (N_11467,N_10439,N_10435);
and U11468 (N_11468,N_10330,N_9802);
and U11469 (N_11469,N_10141,N_10002);
nor U11470 (N_11470,N_9693,N_10168);
nand U11471 (N_11471,N_9478,N_9265);
nand U11472 (N_11472,N_9222,N_9178);
or U11473 (N_11473,N_9443,N_10448);
nor U11474 (N_11474,N_9237,N_9560);
or U11475 (N_11475,N_10160,N_10267);
or U11476 (N_11476,N_10053,N_9515);
nand U11477 (N_11477,N_9740,N_9769);
nand U11478 (N_11478,N_9495,N_10211);
or U11479 (N_11479,N_9242,N_9050);
nor U11480 (N_11480,N_9896,N_9387);
and U11481 (N_11481,N_9374,N_9553);
nand U11482 (N_11482,N_9417,N_9894);
and U11483 (N_11483,N_10279,N_10438);
nor U11484 (N_11484,N_9783,N_9007);
and U11485 (N_11485,N_9066,N_9217);
nand U11486 (N_11486,N_10100,N_9564);
xor U11487 (N_11487,N_10100,N_9555);
and U11488 (N_11488,N_9392,N_9551);
xor U11489 (N_11489,N_9543,N_10151);
and U11490 (N_11490,N_9914,N_10462);
or U11491 (N_11491,N_10312,N_10310);
nor U11492 (N_11492,N_9747,N_10268);
nand U11493 (N_11493,N_10353,N_10488);
nand U11494 (N_11494,N_9183,N_9358);
or U11495 (N_11495,N_9789,N_9126);
nand U11496 (N_11496,N_10444,N_9309);
or U11497 (N_11497,N_9530,N_9647);
or U11498 (N_11498,N_9074,N_9785);
nand U11499 (N_11499,N_10117,N_9914);
nand U11500 (N_11500,N_9363,N_10235);
nor U11501 (N_11501,N_9141,N_10135);
or U11502 (N_11502,N_10058,N_9450);
nor U11503 (N_11503,N_9273,N_10356);
nand U11504 (N_11504,N_10102,N_9751);
nor U11505 (N_11505,N_9483,N_9060);
or U11506 (N_11506,N_10178,N_9911);
or U11507 (N_11507,N_9199,N_9693);
or U11508 (N_11508,N_9833,N_10346);
and U11509 (N_11509,N_9050,N_10049);
nor U11510 (N_11510,N_10196,N_9962);
and U11511 (N_11511,N_9631,N_10255);
and U11512 (N_11512,N_9797,N_9720);
nand U11513 (N_11513,N_9052,N_9689);
and U11514 (N_11514,N_9834,N_9208);
and U11515 (N_11515,N_10270,N_9485);
nand U11516 (N_11516,N_9579,N_10095);
nand U11517 (N_11517,N_10267,N_9073);
nand U11518 (N_11518,N_9867,N_10245);
or U11519 (N_11519,N_10186,N_9621);
nor U11520 (N_11520,N_9824,N_10361);
nor U11521 (N_11521,N_10481,N_9640);
nand U11522 (N_11522,N_10336,N_9255);
nor U11523 (N_11523,N_9501,N_10221);
or U11524 (N_11524,N_9183,N_10343);
or U11525 (N_11525,N_9514,N_10157);
nand U11526 (N_11526,N_9193,N_10329);
nor U11527 (N_11527,N_9757,N_10242);
nand U11528 (N_11528,N_9571,N_10454);
and U11529 (N_11529,N_9342,N_9199);
and U11530 (N_11530,N_9063,N_10266);
xor U11531 (N_11531,N_10178,N_9724);
nor U11532 (N_11532,N_9861,N_9451);
and U11533 (N_11533,N_9729,N_10490);
or U11534 (N_11534,N_10102,N_9499);
nand U11535 (N_11535,N_9395,N_9219);
xnor U11536 (N_11536,N_9055,N_10278);
nand U11537 (N_11537,N_9073,N_10088);
or U11538 (N_11538,N_9385,N_9490);
nand U11539 (N_11539,N_9636,N_10247);
or U11540 (N_11540,N_10425,N_9228);
nand U11541 (N_11541,N_9149,N_10498);
or U11542 (N_11542,N_9322,N_10433);
nor U11543 (N_11543,N_9434,N_10370);
or U11544 (N_11544,N_10126,N_9719);
or U11545 (N_11545,N_9581,N_9307);
and U11546 (N_11546,N_10132,N_9463);
nor U11547 (N_11547,N_10485,N_9618);
or U11548 (N_11548,N_10391,N_10093);
and U11549 (N_11549,N_9960,N_9069);
or U11550 (N_11550,N_9704,N_9055);
nand U11551 (N_11551,N_10030,N_10139);
nand U11552 (N_11552,N_10321,N_9291);
nand U11553 (N_11553,N_9365,N_9910);
and U11554 (N_11554,N_10348,N_10279);
and U11555 (N_11555,N_9472,N_9105);
or U11556 (N_11556,N_9003,N_9459);
nor U11557 (N_11557,N_10260,N_10499);
or U11558 (N_11558,N_10413,N_9075);
and U11559 (N_11559,N_9399,N_9584);
or U11560 (N_11560,N_10230,N_9078);
or U11561 (N_11561,N_10161,N_9786);
or U11562 (N_11562,N_9788,N_10400);
nor U11563 (N_11563,N_10023,N_10269);
or U11564 (N_11564,N_9729,N_9416);
or U11565 (N_11565,N_9837,N_10379);
or U11566 (N_11566,N_9849,N_9416);
and U11567 (N_11567,N_9533,N_10462);
or U11568 (N_11568,N_9458,N_9327);
and U11569 (N_11569,N_9457,N_10496);
xnor U11570 (N_11570,N_9325,N_10429);
nor U11571 (N_11571,N_9411,N_9690);
or U11572 (N_11572,N_10180,N_9995);
and U11573 (N_11573,N_9735,N_9065);
xor U11574 (N_11574,N_9552,N_9667);
and U11575 (N_11575,N_9157,N_9853);
nand U11576 (N_11576,N_9036,N_10194);
nor U11577 (N_11577,N_9673,N_10215);
xnor U11578 (N_11578,N_10113,N_9963);
nand U11579 (N_11579,N_10015,N_10341);
and U11580 (N_11580,N_9046,N_10182);
nor U11581 (N_11581,N_9128,N_10366);
nor U11582 (N_11582,N_9620,N_10289);
nand U11583 (N_11583,N_10147,N_9199);
nor U11584 (N_11584,N_9646,N_9405);
nor U11585 (N_11585,N_10358,N_10442);
nor U11586 (N_11586,N_9450,N_9241);
xnor U11587 (N_11587,N_9806,N_10178);
nand U11588 (N_11588,N_9241,N_9487);
or U11589 (N_11589,N_9224,N_10447);
xnor U11590 (N_11590,N_10335,N_9701);
xnor U11591 (N_11591,N_9657,N_9828);
nand U11592 (N_11592,N_9157,N_10094);
nand U11593 (N_11593,N_10189,N_9463);
nor U11594 (N_11594,N_10474,N_9739);
and U11595 (N_11595,N_10043,N_9693);
nand U11596 (N_11596,N_10225,N_9254);
and U11597 (N_11597,N_9685,N_9973);
or U11598 (N_11598,N_10356,N_9445);
nor U11599 (N_11599,N_10388,N_10274);
or U11600 (N_11600,N_9811,N_9416);
xor U11601 (N_11601,N_9306,N_10420);
xor U11602 (N_11602,N_9699,N_9562);
nor U11603 (N_11603,N_10300,N_10021);
nand U11604 (N_11604,N_9083,N_9541);
nor U11605 (N_11605,N_9348,N_10116);
nor U11606 (N_11606,N_10401,N_10126);
nor U11607 (N_11607,N_10369,N_9000);
nand U11608 (N_11608,N_9864,N_9514);
or U11609 (N_11609,N_9949,N_10410);
xor U11610 (N_11610,N_9484,N_10277);
nor U11611 (N_11611,N_9365,N_10080);
nor U11612 (N_11612,N_10007,N_10010);
and U11613 (N_11613,N_10363,N_10459);
or U11614 (N_11614,N_10392,N_9714);
and U11615 (N_11615,N_9048,N_10126);
or U11616 (N_11616,N_9072,N_9333);
nand U11617 (N_11617,N_9042,N_10251);
and U11618 (N_11618,N_9006,N_9104);
nor U11619 (N_11619,N_10138,N_9886);
or U11620 (N_11620,N_9885,N_9139);
or U11621 (N_11621,N_10470,N_9329);
nand U11622 (N_11622,N_10172,N_9654);
or U11623 (N_11623,N_10176,N_9141);
xor U11624 (N_11624,N_9494,N_9232);
nor U11625 (N_11625,N_9218,N_9645);
nand U11626 (N_11626,N_9639,N_10441);
or U11627 (N_11627,N_9155,N_9241);
or U11628 (N_11628,N_9013,N_10246);
nor U11629 (N_11629,N_10063,N_9901);
xor U11630 (N_11630,N_10222,N_10337);
nor U11631 (N_11631,N_10034,N_9753);
or U11632 (N_11632,N_10241,N_9800);
or U11633 (N_11633,N_9787,N_9382);
and U11634 (N_11634,N_10100,N_10208);
nor U11635 (N_11635,N_9321,N_9374);
nor U11636 (N_11636,N_9745,N_10076);
nand U11637 (N_11637,N_10406,N_9394);
xnor U11638 (N_11638,N_9132,N_10031);
xor U11639 (N_11639,N_9045,N_9905);
nand U11640 (N_11640,N_9225,N_9575);
nand U11641 (N_11641,N_9609,N_9289);
nor U11642 (N_11642,N_10483,N_9394);
nor U11643 (N_11643,N_9899,N_9154);
or U11644 (N_11644,N_9906,N_9300);
xor U11645 (N_11645,N_9873,N_10181);
and U11646 (N_11646,N_10064,N_9706);
and U11647 (N_11647,N_9551,N_9403);
or U11648 (N_11648,N_9114,N_9002);
and U11649 (N_11649,N_9823,N_9340);
xor U11650 (N_11650,N_10424,N_9524);
xnor U11651 (N_11651,N_10228,N_9515);
and U11652 (N_11652,N_10256,N_9732);
and U11653 (N_11653,N_9797,N_9172);
nand U11654 (N_11654,N_10247,N_10453);
xnor U11655 (N_11655,N_10251,N_9556);
and U11656 (N_11656,N_10349,N_10341);
nor U11657 (N_11657,N_9656,N_10260);
and U11658 (N_11658,N_9431,N_10241);
nand U11659 (N_11659,N_9974,N_9339);
nor U11660 (N_11660,N_10446,N_9121);
nor U11661 (N_11661,N_9399,N_10086);
nor U11662 (N_11662,N_9938,N_10329);
nand U11663 (N_11663,N_10246,N_9450);
or U11664 (N_11664,N_10392,N_9172);
or U11665 (N_11665,N_10434,N_10109);
xnor U11666 (N_11666,N_10475,N_10493);
nor U11667 (N_11667,N_9316,N_10471);
and U11668 (N_11668,N_9139,N_10123);
and U11669 (N_11669,N_9299,N_9865);
nand U11670 (N_11670,N_10374,N_10253);
nand U11671 (N_11671,N_9861,N_9554);
xnor U11672 (N_11672,N_9577,N_9422);
nor U11673 (N_11673,N_9291,N_9913);
or U11674 (N_11674,N_9054,N_9616);
xnor U11675 (N_11675,N_9494,N_9411);
xnor U11676 (N_11676,N_9002,N_9903);
nor U11677 (N_11677,N_9679,N_10232);
and U11678 (N_11678,N_10000,N_10263);
and U11679 (N_11679,N_10122,N_9874);
or U11680 (N_11680,N_9335,N_9177);
or U11681 (N_11681,N_9103,N_10152);
nor U11682 (N_11682,N_9920,N_10230);
xnor U11683 (N_11683,N_9896,N_9769);
and U11684 (N_11684,N_9882,N_9368);
or U11685 (N_11685,N_9615,N_9011);
and U11686 (N_11686,N_9172,N_9194);
nand U11687 (N_11687,N_9743,N_9737);
nand U11688 (N_11688,N_9530,N_9625);
nand U11689 (N_11689,N_9868,N_9236);
and U11690 (N_11690,N_9430,N_9206);
nand U11691 (N_11691,N_9547,N_10314);
or U11692 (N_11692,N_10265,N_10409);
nand U11693 (N_11693,N_10198,N_9769);
and U11694 (N_11694,N_9554,N_9725);
nand U11695 (N_11695,N_10116,N_10012);
nand U11696 (N_11696,N_10455,N_9805);
and U11697 (N_11697,N_9002,N_10170);
nor U11698 (N_11698,N_9129,N_10104);
nor U11699 (N_11699,N_9734,N_10032);
and U11700 (N_11700,N_9993,N_9987);
nor U11701 (N_11701,N_9260,N_10016);
or U11702 (N_11702,N_10010,N_10055);
nor U11703 (N_11703,N_10110,N_9417);
and U11704 (N_11704,N_9903,N_9639);
nor U11705 (N_11705,N_9376,N_9142);
nand U11706 (N_11706,N_9223,N_9231);
and U11707 (N_11707,N_9463,N_10427);
nand U11708 (N_11708,N_10035,N_9867);
or U11709 (N_11709,N_10429,N_9271);
nor U11710 (N_11710,N_9355,N_9024);
xnor U11711 (N_11711,N_9973,N_9720);
or U11712 (N_11712,N_9701,N_9417);
xnor U11713 (N_11713,N_10098,N_9125);
and U11714 (N_11714,N_9744,N_9421);
nand U11715 (N_11715,N_10034,N_9675);
or U11716 (N_11716,N_10485,N_10472);
and U11717 (N_11717,N_9084,N_9055);
nand U11718 (N_11718,N_9993,N_9523);
nand U11719 (N_11719,N_10447,N_9852);
nor U11720 (N_11720,N_9985,N_10372);
nor U11721 (N_11721,N_9597,N_10104);
and U11722 (N_11722,N_9518,N_9344);
nand U11723 (N_11723,N_10150,N_9625);
nor U11724 (N_11724,N_9297,N_10489);
and U11725 (N_11725,N_10149,N_10354);
or U11726 (N_11726,N_9721,N_10361);
or U11727 (N_11727,N_9309,N_10275);
nor U11728 (N_11728,N_9605,N_9667);
or U11729 (N_11729,N_9032,N_9894);
and U11730 (N_11730,N_9774,N_9577);
nand U11731 (N_11731,N_9100,N_10013);
nor U11732 (N_11732,N_10440,N_10384);
nand U11733 (N_11733,N_9871,N_10381);
or U11734 (N_11734,N_9314,N_9351);
nand U11735 (N_11735,N_10004,N_9502);
nor U11736 (N_11736,N_10420,N_10389);
nand U11737 (N_11737,N_9194,N_10228);
nor U11738 (N_11738,N_9312,N_9042);
nor U11739 (N_11739,N_10461,N_9474);
nand U11740 (N_11740,N_10278,N_10044);
and U11741 (N_11741,N_10458,N_9341);
or U11742 (N_11742,N_9946,N_9844);
nand U11743 (N_11743,N_10038,N_9372);
nand U11744 (N_11744,N_9979,N_9469);
xor U11745 (N_11745,N_10167,N_10233);
nand U11746 (N_11746,N_9527,N_9388);
or U11747 (N_11747,N_10062,N_9981);
and U11748 (N_11748,N_9225,N_10222);
xnor U11749 (N_11749,N_9855,N_9214);
nor U11750 (N_11750,N_9120,N_10383);
nor U11751 (N_11751,N_10196,N_10412);
or U11752 (N_11752,N_9140,N_9325);
or U11753 (N_11753,N_9021,N_9376);
nor U11754 (N_11754,N_10281,N_10039);
nor U11755 (N_11755,N_10124,N_9466);
nor U11756 (N_11756,N_10364,N_9204);
and U11757 (N_11757,N_10490,N_9035);
or U11758 (N_11758,N_9576,N_9152);
or U11759 (N_11759,N_10452,N_10307);
nor U11760 (N_11760,N_10383,N_9081);
nand U11761 (N_11761,N_10117,N_10330);
xnor U11762 (N_11762,N_10216,N_9783);
or U11763 (N_11763,N_9921,N_9711);
nor U11764 (N_11764,N_9429,N_9537);
nor U11765 (N_11765,N_9597,N_10017);
nor U11766 (N_11766,N_9592,N_10282);
or U11767 (N_11767,N_9322,N_9030);
or U11768 (N_11768,N_10412,N_10335);
and U11769 (N_11769,N_9679,N_10060);
nor U11770 (N_11770,N_9261,N_10285);
nor U11771 (N_11771,N_9565,N_10138);
nand U11772 (N_11772,N_10295,N_10261);
nor U11773 (N_11773,N_9119,N_9384);
nor U11774 (N_11774,N_9636,N_9669);
nand U11775 (N_11775,N_10323,N_10137);
and U11776 (N_11776,N_9363,N_10069);
xor U11777 (N_11777,N_10309,N_9778);
and U11778 (N_11778,N_9933,N_9273);
and U11779 (N_11779,N_9880,N_9561);
nand U11780 (N_11780,N_9759,N_9815);
and U11781 (N_11781,N_9473,N_9318);
nand U11782 (N_11782,N_9462,N_10470);
and U11783 (N_11783,N_9555,N_9398);
and U11784 (N_11784,N_10197,N_9949);
nand U11785 (N_11785,N_9968,N_9627);
or U11786 (N_11786,N_9083,N_9993);
nor U11787 (N_11787,N_10371,N_9260);
and U11788 (N_11788,N_9417,N_9468);
nor U11789 (N_11789,N_9440,N_9553);
and U11790 (N_11790,N_9932,N_10071);
nor U11791 (N_11791,N_9804,N_10290);
and U11792 (N_11792,N_10091,N_10022);
nor U11793 (N_11793,N_10096,N_9597);
or U11794 (N_11794,N_10127,N_10356);
and U11795 (N_11795,N_9430,N_9375);
nor U11796 (N_11796,N_10005,N_9904);
nand U11797 (N_11797,N_9527,N_9309);
or U11798 (N_11798,N_10155,N_9111);
nor U11799 (N_11799,N_9153,N_9768);
nor U11800 (N_11800,N_10422,N_10485);
nor U11801 (N_11801,N_9444,N_9631);
nor U11802 (N_11802,N_10323,N_9604);
nand U11803 (N_11803,N_9457,N_10384);
nand U11804 (N_11804,N_9106,N_9633);
and U11805 (N_11805,N_9251,N_10372);
or U11806 (N_11806,N_9436,N_9209);
nor U11807 (N_11807,N_10139,N_9146);
and U11808 (N_11808,N_10395,N_10266);
nor U11809 (N_11809,N_9478,N_10412);
nand U11810 (N_11810,N_9658,N_9530);
and U11811 (N_11811,N_9059,N_9108);
nand U11812 (N_11812,N_10079,N_10496);
xor U11813 (N_11813,N_10057,N_9230);
or U11814 (N_11814,N_10100,N_9738);
and U11815 (N_11815,N_9331,N_9734);
and U11816 (N_11816,N_9234,N_9551);
or U11817 (N_11817,N_9524,N_9395);
nand U11818 (N_11818,N_10213,N_9059);
or U11819 (N_11819,N_9276,N_9715);
and U11820 (N_11820,N_9440,N_10483);
or U11821 (N_11821,N_9355,N_9116);
xor U11822 (N_11822,N_9458,N_9318);
nor U11823 (N_11823,N_9247,N_9453);
nor U11824 (N_11824,N_10428,N_10013);
and U11825 (N_11825,N_9508,N_9385);
nor U11826 (N_11826,N_9893,N_9495);
nand U11827 (N_11827,N_9817,N_10299);
nor U11828 (N_11828,N_9231,N_9382);
and U11829 (N_11829,N_9751,N_9995);
and U11830 (N_11830,N_9341,N_9432);
or U11831 (N_11831,N_9191,N_10475);
nand U11832 (N_11832,N_10413,N_9319);
and U11833 (N_11833,N_9368,N_9565);
nand U11834 (N_11834,N_10218,N_9923);
nor U11835 (N_11835,N_9579,N_9945);
and U11836 (N_11836,N_10447,N_9586);
xnor U11837 (N_11837,N_9525,N_9189);
or U11838 (N_11838,N_9888,N_9050);
xnor U11839 (N_11839,N_9266,N_10224);
nand U11840 (N_11840,N_9316,N_10484);
and U11841 (N_11841,N_9836,N_10162);
xor U11842 (N_11842,N_10349,N_9064);
or U11843 (N_11843,N_9251,N_9014);
nand U11844 (N_11844,N_9714,N_10439);
and U11845 (N_11845,N_10237,N_10016);
nor U11846 (N_11846,N_9303,N_9355);
nand U11847 (N_11847,N_10140,N_9765);
nand U11848 (N_11848,N_9091,N_9631);
nand U11849 (N_11849,N_9674,N_9993);
and U11850 (N_11850,N_9708,N_10238);
nand U11851 (N_11851,N_9732,N_9316);
and U11852 (N_11852,N_10344,N_9491);
or U11853 (N_11853,N_9074,N_10335);
and U11854 (N_11854,N_10498,N_9485);
nor U11855 (N_11855,N_9309,N_10096);
xor U11856 (N_11856,N_10391,N_10057);
and U11857 (N_11857,N_10192,N_9361);
and U11858 (N_11858,N_9966,N_9770);
or U11859 (N_11859,N_9771,N_9709);
or U11860 (N_11860,N_9641,N_10096);
and U11861 (N_11861,N_9199,N_9096);
or U11862 (N_11862,N_10074,N_10289);
nor U11863 (N_11863,N_9816,N_9346);
and U11864 (N_11864,N_9046,N_10481);
nand U11865 (N_11865,N_10167,N_10469);
nor U11866 (N_11866,N_10116,N_9493);
nor U11867 (N_11867,N_9386,N_9879);
nor U11868 (N_11868,N_9988,N_10140);
nand U11869 (N_11869,N_10463,N_9221);
nor U11870 (N_11870,N_9087,N_9900);
nand U11871 (N_11871,N_10496,N_9238);
nand U11872 (N_11872,N_9244,N_9267);
and U11873 (N_11873,N_9664,N_9393);
nand U11874 (N_11874,N_9255,N_9217);
and U11875 (N_11875,N_9592,N_9777);
or U11876 (N_11876,N_10161,N_9524);
nor U11877 (N_11877,N_9816,N_9736);
nor U11878 (N_11878,N_9525,N_9826);
xnor U11879 (N_11879,N_9403,N_9953);
and U11880 (N_11880,N_9317,N_9838);
nand U11881 (N_11881,N_10071,N_10115);
nor U11882 (N_11882,N_9886,N_9740);
nor U11883 (N_11883,N_9591,N_10036);
or U11884 (N_11884,N_9229,N_10375);
or U11885 (N_11885,N_10052,N_10224);
or U11886 (N_11886,N_9317,N_10272);
nand U11887 (N_11887,N_10328,N_9385);
nand U11888 (N_11888,N_9558,N_9778);
or U11889 (N_11889,N_9517,N_10197);
nor U11890 (N_11890,N_9848,N_9443);
nand U11891 (N_11891,N_9575,N_9788);
or U11892 (N_11892,N_10247,N_10386);
or U11893 (N_11893,N_9741,N_9597);
nand U11894 (N_11894,N_9017,N_9708);
nand U11895 (N_11895,N_9480,N_10490);
nand U11896 (N_11896,N_9802,N_9635);
or U11897 (N_11897,N_9560,N_9214);
and U11898 (N_11898,N_9387,N_9305);
nor U11899 (N_11899,N_10367,N_10391);
nand U11900 (N_11900,N_9838,N_9339);
and U11901 (N_11901,N_10132,N_9566);
and U11902 (N_11902,N_9597,N_9785);
xor U11903 (N_11903,N_9704,N_10208);
or U11904 (N_11904,N_9469,N_10375);
or U11905 (N_11905,N_10283,N_9500);
or U11906 (N_11906,N_10493,N_9010);
or U11907 (N_11907,N_9790,N_9727);
or U11908 (N_11908,N_10494,N_9143);
nand U11909 (N_11909,N_9546,N_10292);
nand U11910 (N_11910,N_10187,N_9669);
and U11911 (N_11911,N_10390,N_10443);
and U11912 (N_11912,N_10365,N_10263);
nand U11913 (N_11913,N_9782,N_9793);
nand U11914 (N_11914,N_9027,N_9271);
or U11915 (N_11915,N_10059,N_10305);
nor U11916 (N_11916,N_9177,N_10112);
nand U11917 (N_11917,N_9829,N_10042);
and U11918 (N_11918,N_9496,N_10151);
and U11919 (N_11919,N_9816,N_9269);
nor U11920 (N_11920,N_10307,N_9294);
nor U11921 (N_11921,N_9049,N_9755);
or U11922 (N_11922,N_9869,N_9903);
and U11923 (N_11923,N_10053,N_9163);
nor U11924 (N_11924,N_9187,N_10160);
nor U11925 (N_11925,N_9733,N_9616);
xnor U11926 (N_11926,N_10366,N_9063);
nand U11927 (N_11927,N_9764,N_9373);
and U11928 (N_11928,N_9306,N_9089);
nand U11929 (N_11929,N_9027,N_9390);
and U11930 (N_11930,N_9642,N_10214);
nor U11931 (N_11931,N_9575,N_9530);
and U11932 (N_11932,N_9392,N_9624);
nor U11933 (N_11933,N_10385,N_10492);
and U11934 (N_11934,N_10379,N_9787);
nor U11935 (N_11935,N_10341,N_9968);
and U11936 (N_11936,N_9683,N_10244);
nor U11937 (N_11937,N_9046,N_10149);
nand U11938 (N_11938,N_9830,N_9946);
nand U11939 (N_11939,N_9584,N_10337);
and U11940 (N_11940,N_10400,N_9481);
or U11941 (N_11941,N_9632,N_9982);
and U11942 (N_11942,N_9615,N_9878);
and U11943 (N_11943,N_10476,N_9216);
nor U11944 (N_11944,N_10277,N_9002);
nand U11945 (N_11945,N_9118,N_9789);
and U11946 (N_11946,N_9212,N_10089);
nor U11947 (N_11947,N_10123,N_9887);
and U11948 (N_11948,N_9210,N_10203);
or U11949 (N_11949,N_10479,N_9178);
nand U11950 (N_11950,N_9156,N_9129);
xor U11951 (N_11951,N_10078,N_9315);
nand U11952 (N_11952,N_9467,N_9055);
nor U11953 (N_11953,N_9091,N_10374);
nand U11954 (N_11954,N_9682,N_9846);
and U11955 (N_11955,N_9839,N_10226);
nor U11956 (N_11956,N_9163,N_9613);
and U11957 (N_11957,N_9076,N_10006);
nand U11958 (N_11958,N_10253,N_10000);
or U11959 (N_11959,N_9141,N_9075);
nor U11960 (N_11960,N_10458,N_10392);
nor U11961 (N_11961,N_9735,N_9778);
xnor U11962 (N_11962,N_9099,N_9218);
nand U11963 (N_11963,N_10106,N_9792);
or U11964 (N_11964,N_10371,N_9113);
nor U11965 (N_11965,N_9685,N_9105);
or U11966 (N_11966,N_10483,N_9511);
or U11967 (N_11967,N_9224,N_9128);
or U11968 (N_11968,N_9960,N_9874);
or U11969 (N_11969,N_10456,N_9492);
or U11970 (N_11970,N_9813,N_9097);
nor U11971 (N_11971,N_10082,N_10483);
and U11972 (N_11972,N_10143,N_10452);
and U11973 (N_11973,N_9884,N_9213);
xor U11974 (N_11974,N_9088,N_9827);
nand U11975 (N_11975,N_9337,N_9736);
or U11976 (N_11976,N_9921,N_10013);
nand U11977 (N_11977,N_9515,N_9972);
and U11978 (N_11978,N_9360,N_9470);
nand U11979 (N_11979,N_9531,N_9207);
and U11980 (N_11980,N_10246,N_9481);
nand U11981 (N_11981,N_9514,N_10184);
nor U11982 (N_11982,N_9075,N_9199);
or U11983 (N_11983,N_9625,N_9614);
nor U11984 (N_11984,N_9416,N_9199);
or U11985 (N_11985,N_9842,N_9668);
or U11986 (N_11986,N_9751,N_9320);
or U11987 (N_11987,N_9463,N_9874);
nor U11988 (N_11988,N_10207,N_9299);
nand U11989 (N_11989,N_9663,N_9784);
or U11990 (N_11990,N_10475,N_10346);
or U11991 (N_11991,N_10106,N_10115);
nor U11992 (N_11992,N_10331,N_9951);
and U11993 (N_11993,N_10194,N_9438);
nor U11994 (N_11994,N_9345,N_9756);
nor U11995 (N_11995,N_10474,N_9164);
or U11996 (N_11996,N_9667,N_10349);
nor U11997 (N_11997,N_10351,N_10264);
and U11998 (N_11998,N_9634,N_10297);
nand U11999 (N_11999,N_9942,N_9615);
nor U12000 (N_12000,N_11501,N_11460);
or U12001 (N_12001,N_11352,N_11058);
or U12002 (N_12002,N_11739,N_10994);
and U12003 (N_12003,N_10590,N_10610);
nor U12004 (N_12004,N_11286,N_11988);
and U12005 (N_12005,N_11504,N_10622);
nor U12006 (N_12006,N_11257,N_11600);
nor U12007 (N_12007,N_11836,N_11455);
nor U12008 (N_12008,N_11278,N_11081);
and U12009 (N_12009,N_10624,N_10714);
nor U12010 (N_12010,N_11473,N_11125);
or U12011 (N_12011,N_10914,N_11420);
or U12012 (N_12012,N_11881,N_11467);
nand U12013 (N_12013,N_11395,N_11032);
and U12014 (N_12014,N_10794,N_11475);
nor U12015 (N_12015,N_10619,N_11775);
and U12016 (N_12016,N_10996,N_11583);
and U12017 (N_12017,N_11917,N_11176);
or U12018 (N_12018,N_10621,N_11969);
nand U12019 (N_12019,N_10685,N_11985);
xor U12020 (N_12020,N_11172,N_10552);
and U12021 (N_12021,N_10861,N_11790);
or U12022 (N_12022,N_10859,N_11797);
xor U12023 (N_12023,N_10691,N_11750);
or U12024 (N_12024,N_11579,N_11535);
xor U12025 (N_12025,N_11412,N_11464);
xor U12026 (N_12026,N_11159,N_11134);
and U12027 (N_12027,N_11981,N_11347);
and U12028 (N_12028,N_11670,N_11288);
and U12029 (N_12029,N_11823,N_11009);
and U12030 (N_12030,N_10952,N_11121);
or U12031 (N_12031,N_10586,N_10733);
xor U12032 (N_12032,N_10991,N_11962);
or U12033 (N_12033,N_11503,N_11841);
nand U12034 (N_12034,N_10767,N_10814);
nor U12035 (N_12035,N_11915,N_11530);
or U12036 (N_12036,N_11242,N_11760);
nand U12037 (N_12037,N_10611,N_10900);
nor U12038 (N_12038,N_10742,N_11961);
nor U12039 (N_12039,N_11371,N_10908);
or U12040 (N_12040,N_11366,N_11311);
nand U12041 (N_12041,N_11472,N_11163);
nand U12042 (N_12042,N_11238,N_11339);
or U12043 (N_12043,N_10819,N_11997);
and U12044 (N_12044,N_10762,N_10632);
nand U12045 (N_12045,N_11629,N_11118);
nor U12046 (N_12046,N_10508,N_11213);
or U12047 (N_12047,N_10707,N_11633);
and U12048 (N_12048,N_11882,N_11338);
nor U12049 (N_12049,N_11859,N_11798);
and U12050 (N_12050,N_11306,N_11016);
xnor U12051 (N_12051,N_10573,N_10647);
xor U12052 (N_12052,N_11335,N_11830);
nor U12053 (N_12053,N_11914,N_11133);
nand U12054 (N_12054,N_11035,N_11452);
and U12055 (N_12055,N_11280,N_10515);
nand U12056 (N_12056,N_10858,N_10982);
or U12057 (N_12057,N_10744,N_10846);
xnor U12058 (N_12058,N_10974,N_10957);
and U12059 (N_12059,N_11062,N_11314);
or U12060 (N_12060,N_10516,N_11324);
or U12061 (N_12061,N_10678,N_11142);
nand U12062 (N_12062,N_11768,N_11619);
nand U12063 (N_12063,N_10787,N_11900);
nand U12064 (N_12064,N_10877,N_11196);
nand U12065 (N_12065,N_11792,N_11965);
nor U12066 (N_12066,N_11038,N_11814);
or U12067 (N_12067,N_11104,N_11466);
or U12068 (N_12068,N_11683,N_10972);
or U12069 (N_12069,N_11788,N_10514);
nor U12070 (N_12070,N_10860,N_11899);
nor U12071 (N_12071,N_10944,N_11313);
or U12072 (N_12072,N_11514,N_10580);
nand U12073 (N_12073,N_11766,N_11291);
or U12074 (N_12074,N_11774,N_10776);
and U12075 (N_12075,N_10725,N_10689);
or U12076 (N_12076,N_11640,N_10649);
nor U12077 (N_12077,N_11363,N_11487);
and U12078 (N_12078,N_10571,N_10987);
nand U12079 (N_12079,N_11853,N_11974);
xnor U12080 (N_12080,N_10539,N_10953);
nor U12081 (N_12081,N_10576,N_11925);
and U12082 (N_12082,N_11883,N_11236);
nor U12083 (N_12083,N_11270,N_11254);
nand U12084 (N_12084,N_10839,N_11046);
nor U12085 (N_12085,N_10793,N_11920);
nor U12086 (N_12086,N_10640,N_11543);
nor U12087 (N_12087,N_11717,N_11239);
and U12088 (N_12088,N_11012,N_11279);
and U12089 (N_12089,N_10663,N_11197);
xnor U12090 (N_12090,N_10880,N_11927);
nor U12091 (N_12091,N_11327,N_10889);
nand U12092 (N_12092,N_10977,N_11827);
xnor U12093 (N_12093,N_11409,N_10894);
or U12094 (N_12094,N_11036,N_11672);
nor U12095 (N_12095,N_10631,N_11716);
nand U12096 (N_12096,N_10822,N_10706);
or U12097 (N_12097,N_11800,N_11701);
nand U12098 (N_12098,N_11442,N_11843);
or U12099 (N_12099,N_11525,N_11993);
nor U12100 (N_12100,N_11382,N_11357);
nand U12101 (N_12101,N_11975,N_10556);
nand U12102 (N_12102,N_11676,N_11149);
or U12103 (N_12103,N_11088,N_11305);
and U12104 (N_12104,N_11607,N_11057);
and U12105 (N_12105,N_11041,N_10739);
xnor U12106 (N_12106,N_10560,N_10921);
and U12107 (N_12107,N_11761,N_10710);
and U12108 (N_12108,N_11734,N_10965);
or U12109 (N_12109,N_10716,N_11650);
and U12110 (N_12110,N_10599,N_11942);
or U12111 (N_12111,N_11065,N_11707);
nor U12112 (N_12112,N_10978,N_11093);
xor U12113 (N_12113,N_10916,N_11937);
or U12114 (N_12114,N_11740,N_10713);
and U12115 (N_12115,N_11317,N_11253);
nor U12116 (N_12116,N_11381,N_11918);
xnor U12117 (N_12117,N_11434,N_10764);
nand U12118 (N_12118,N_10973,N_10771);
nor U12119 (N_12119,N_11380,N_10786);
or U12120 (N_12120,N_10595,N_11591);
or U12121 (N_12121,N_11580,N_11101);
or U12122 (N_12122,N_10934,N_11665);
or U12123 (N_12123,N_11470,N_11561);
nor U12124 (N_12124,N_10785,N_11850);
xnor U12125 (N_12125,N_11052,N_10761);
nand U12126 (N_12126,N_11906,N_11803);
nor U12127 (N_12127,N_11166,N_11778);
nor U12128 (N_12128,N_11938,N_10538);
and U12129 (N_12129,N_11231,N_11515);
nor U12130 (N_12130,N_10630,N_10734);
and U12131 (N_12131,N_10643,N_11560);
and U12132 (N_12132,N_11916,N_11256);
nand U12133 (N_12133,N_10768,N_11073);
nor U12134 (N_12134,N_11621,N_11978);
xor U12135 (N_12135,N_11705,N_11789);
nor U12136 (N_12136,N_11287,N_11384);
and U12137 (N_12137,N_11154,N_11893);
or U12138 (N_12138,N_11471,N_11011);
nor U12139 (N_12139,N_11932,N_11128);
or U12140 (N_12140,N_11982,N_11903);
nor U12141 (N_12141,N_10812,N_10728);
or U12142 (N_12142,N_11980,N_11266);
nand U12143 (N_12143,N_11043,N_11725);
or U12144 (N_12144,N_11263,N_11599);
nor U12145 (N_12145,N_11265,N_10535);
nand U12146 (N_12146,N_11753,N_11871);
and U12147 (N_12147,N_10789,N_11585);
and U12148 (N_12148,N_11763,N_10993);
xnor U12149 (N_12149,N_11811,N_11341);
nor U12150 (N_12150,N_11603,N_10703);
or U12151 (N_12151,N_11427,N_11576);
and U12152 (N_12152,N_11838,N_11158);
or U12153 (N_12153,N_11553,N_11877);
nor U12154 (N_12154,N_10844,N_11330);
or U12155 (N_12155,N_11542,N_11520);
or U12156 (N_12156,N_11641,N_11414);
nand U12157 (N_12157,N_11546,N_10718);
nand U12158 (N_12158,N_10740,N_11379);
nor U12159 (N_12159,N_10567,N_11747);
nand U12160 (N_12160,N_11564,N_10989);
nor U12161 (N_12161,N_11069,N_11879);
and U12162 (N_12162,N_10808,N_10667);
nor U12163 (N_12163,N_10682,N_10796);
and U12164 (N_12164,N_10609,N_11976);
and U12165 (N_12165,N_10801,N_10605);
xnor U12166 (N_12166,N_11157,N_10745);
and U12167 (N_12167,N_10532,N_11923);
or U12168 (N_12168,N_10960,N_11067);
nand U12169 (N_12169,N_11512,N_10543);
or U12170 (N_12170,N_10887,N_11730);
nor U12171 (N_12171,N_10730,N_11781);
or U12172 (N_12172,N_11084,N_10520);
or U12173 (N_12173,N_11362,N_11572);
and U12174 (N_12174,N_11365,N_11096);
or U12175 (N_12175,N_11094,N_11147);
or U12176 (N_12176,N_11887,N_11557);
nand U12177 (N_12177,N_11675,N_10709);
or U12178 (N_12178,N_11541,N_11044);
nor U12179 (N_12179,N_10705,N_10855);
nor U12180 (N_12180,N_10522,N_11198);
xnor U12181 (N_12181,N_11489,N_10815);
nand U12182 (N_12182,N_10980,N_10551);
and U12183 (N_12183,N_11200,N_11548);
nor U12184 (N_12184,N_10866,N_11045);
or U12185 (N_12185,N_11889,N_11934);
nand U12186 (N_12186,N_10760,N_10988);
and U12187 (N_12187,N_11419,N_11521);
nand U12188 (N_12188,N_10669,N_11224);
nor U12189 (N_12189,N_10747,N_10902);
and U12190 (N_12190,N_10909,N_10884);
xnor U12191 (N_12191,N_11397,N_11894);
xnor U12192 (N_12192,N_11896,N_10969);
nand U12193 (N_12193,N_11491,N_11060);
xor U12194 (N_12194,N_10506,N_11223);
and U12195 (N_12195,N_11483,N_11657);
nand U12196 (N_12196,N_11168,N_10911);
nor U12197 (N_12197,N_10658,N_11804);
nor U12198 (N_12198,N_11193,N_11951);
and U12199 (N_12199,N_11430,N_11644);
and U12200 (N_12200,N_10806,N_11960);
or U12201 (N_12201,N_11114,N_11596);
and U12202 (N_12202,N_11465,N_11661);
and U12203 (N_12203,N_10672,N_11127);
nor U12204 (N_12204,N_11486,N_10869);
nand U12205 (N_12205,N_11769,N_11735);
and U12206 (N_12206,N_11589,N_11669);
nor U12207 (N_12207,N_11729,N_11570);
nand U12208 (N_12208,N_11010,N_10687);
and U12209 (N_12209,N_11275,N_11972);
nand U12210 (N_12210,N_10698,N_11271);
or U12211 (N_12211,N_11303,N_11639);
nor U12212 (N_12212,N_11642,N_10601);
and U12213 (N_12213,N_11048,N_11684);
or U12214 (N_12214,N_11428,N_10804);
nor U12215 (N_12215,N_10995,N_11711);
nand U12216 (N_12216,N_10545,N_10606);
and U12217 (N_12217,N_10939,N_11499);
xnor U12218 (N_12218,N_11526,N_11777);
or U12219 (N_12219,N_11137,N_11849);
nand U12220 (N_12220,N_11040,N_11416);
nor U12221 (N_12221,N_11097,N_11724);
and U12222 (N_12222,N_11261,N_11034);
nand U12223 (N_12223,N_11214,N_11531);
nor U12224 (N_12224,N_11723,N_11813);
nand U12225 (N_12225,N_11353,N_10961);
or U12226 (N_12226,N_11374,N_11631);
and U12227 (N_12227,N_11174,N_11481);
nor U12228 (N_12228,N_11952,N_10942);
nand U12229 (N_12229,N_11156,N_11431);
nor U12230 (N_12230,N_10779,N_11108);
and U12231 (N_12231,N_11630,N_10549);
and U12232 (N_12232,N_11605,N_10526);
nor U12233 (N_12233,N_11354,N_11226);
nor U12234 (N_12234,N_11516,N_11581);
and U12235 (N_12235,N_11806,N_10655);
and U12236 (N_12236,N_11979,N_11232);
and U12237 (N_12237,N_11150,N_11139);
nand U12238 (N_12238,N_11839,N_11245);
or U12239 (N_12239,N_11574,N_11819);
nor U12240 (N_12240,N_11569,N_11398);
or U12241 (N_12241,N_11540,N_10583);
and U12242 (N_12242,N_11905,N_11064);
or U12243 (N_12243,N_11228,N_11234);
nand U12244 (N_12244,N_11578,N_10507);
nor U12245 (N_12245,N_11875,N_11722);
nor U12246 (N_12246,N_11418,N_11926);
xor U12247 (N_12247,N_10818,N_11904);
and U12248 (N_12248,N_11396,N_10845);
xor U12249 (N_12249,N_11169,N_11831);
nand U12250 (N_12250,N_11528,N_11872);
and U12251 (N_12251,N_11008,N_11003);
nor U12252 (N_12252,N_11854,N_10770);
xor U12253 (N_12253,N_10907,N_11162);
xor U12254 (N_12254,N_10755,N_11509);
and U12255 (N_12255,N_10616,N_11647);
nand U12256 (N_12256,N_11216,N_11756);
or U12257 (N_12257,N_10736,N_11664);
or U12258 (N_12258,N_10662,N_11293);
nand U12259 (N_12259,N_11924,N_11217);
and U12260 (N_12260,N_10751,N_10603);
nand U12261 (N_12261,N_10842,N_10854);
or U12262 (N_12262,N_10863,N_11229);
or U12263 (N_12263,N_11241,N_11493);
and U12264 (N_12264,N_11623,N_10851);
nor U12265 (N_12265,N_11613,N_11911);
and U12266 (N_12266,N_11129,N_11828);
or U12267 (N_12267,N_10829,N_11113);
or U12268 (N_12268,N_11793,N_10912);
nand U12269 (N_12269,N_11026,N_11055);
and U12270 (N_12270,N_11674,N_11340);
or U12271 (N_12271,N_11592,N_11334);
nor U12272 (N_12272,N_11205,N_11891);
nor U12273 (N_12273,N_11696,N_11289);
or U12274 (N_12274,N_11145,N_11654);
and U12275 (N_12275,N_11506,N_10864);
or U12276 (N_12276,N_10541,N_11086);
and U12277 (N_12277,N_10935,N_10857);
xor U12278 (N_12278,N_11435,N_11143);
and U12279 (N_12279,N_10901,N_11402);
nor U12280 (N_12280,N_11627,N_11267);
xnor U12281 (N_12281,N_10671,N_11651);
nor U12282 (N_12282,N_11290,N_11689);
nand U12283 (N_12283,N_11207,N_11533);
nand U12284 (N_12284,N_10597,N_10686);
nand U12285 (N_12285,N_11555,N_11700);
nand U12286 (N_12286,N_11594,N_11027);
and U12287 (N_12287,N_11868,N_11710);
nor U12288 (N_12288,N_10849,N_10546);
nor U12289 (N_12289,N_10651,N_11861);
and U12290 (N_12290,N_11478,N_11999);
and U12291 (N_12291,N_10588,N_11480);
or U12292 (N_12292,N_10654,N_11105);
and U12293 (N_12293,N_11954,N_10653);
and U12294 (N_12294,N_11047,N_11461);
nand U12295 (N_12295,N_10749,N_11928);
nor U12296 (N_12296,N_10743,N_11636);
nor U12297 (N_12297,N_11070,N_11780);
and U12298 (N_12298,N_11549,N_11856);
nand U12299 (N_12299,N_11686,N_11488);
nor U12300 (N_12300,N_11391,N_10676);
or U12301 (N_12301,N_11946,N_11712);
nand U12302 (N_12302,N_11869,N_10578);
nand U12303 (N_12303,N_11325,N_10906);
or U12304 (N_12304,N_11106,N_11862);
nor U12305 (N_12305,N_10668,N_11744);
or U12306 (N_12306,N_11100,N_10792);
and U12307 (N_12307,N_10592,N_10711);
and U12308 (N_12308,N_11930,N_10915);
nand U12309 (N_12309,N_11706,N_10614);
and U12310 (N_12310,N_11272,N_10838);
xnor U12311 (N_12311,N_10598,N_11816);
and U12312 (N_12312,N_11837,N_11643);
nor U12313 (N_12313,N_11237,N_11323);
nor U12314 (N_12314,N_10579,N_10505);
nand U12315 (N_12315,N_10874,N_11588);
xor U12316 (N_12316,N_10945,N_11179);
nor U12317 (N_12317,N_11028,N_11273);
or U12318 (N_12318,N_11929,N_11551);
nor U12319 (N_12319,N_11662,N_10847);
or U12320 (N_12320,N_10832,N_11160);
or U12321 (N_12321,N_11678,N_11109);
nor U12322 (N_12322,N_11984,N_10738);
nand U12323 (N_12323,N_11146,N_10811);
nor U12324 (N_12324,N_11948,N_11746);
and U12325 (N_12325,N_11848,N_10600);
nor U12326 (N_12326,N_11191,N_11264);
xnor U12327 (N_12327,N_11945,N_11284);
nor U12328 (N_12328,N_10502,N_10523);
nor U12329 (N_12329,N_11072,N_11112);
and U12330 (N_12330,N_11593,N_10753);
and U12331 (N_12331,N_10897,N_11310);
or U12332 (N_12332,N_10544,N_10783);
and U12333 (N_12333,N_11815,N_10591);
nor U12334 (N_12334,N_11298,N_11632);
nor U12335 (N_12335,N_11614,N_10958);
nor U12336 (N_12336,N_10639,N_11233);
and U12337 (N_12337,N_11152,N_11616);
and U12338 (N_12338,N_10809,N_11500);
or U12339 (N_12339,N_10841,N_11649);
nand U12340 (N_12340,N_10999,N_10719);
nand U12341 (N_12341,N_11567,N_11620);
or U12342 (N_12342,N_11292,N_11646);
nand U12343 (N_12343,N_11453,N_10636);
nand U12344 (N_12344,N_10959,N_11971);
and U12345 (N_12345,N_11846,N_11751);
xnor U12346 (N_12346,N_11755,N_10984);
and U12347 (N_12347,N_11405,N_10879);
and U12348 (N_12348,N_11731,N_10933);
xor U12349 (N_12349,N_11030,N_11432);
nor U12350 (N_12350,N_10823,N_11385);
and U12351 (N_12351,N_10848,N_11022);
and U12352 (N_12352,N_11359,N_11429);
nor U12353 (N_12353,N_10593,N_11004);
or U12354 (N_12354,N_11252,N_10670);
nand U12355 (N_12355,N_11776,N_11206);
or U12356 (N_12356,N_11155,N_11822);
nor U12357 (N_12357,N_11842,N_11824);
xnor U12358 (N_12358,N_11496,N_10941);
nor U12359 (N_12359,N_10684,N_11860);
nand U12360 (N_12360,N_10701,N_11728);
nand U12361 (N_12361,N_10585,N_10873);
nor U12362 (N_12362,N_11652,N_10582);
and U12363 (N_12363,N_10641,N_11437);
nand U12364 (N_12364,N_11110,N_11350);
nor U12365 (N_12365,N_10704,N_11433);
nor U12366 (N_12366,N_10550,N_10837);
nor U12367 (N_12367,N_10681,N_10910);
and U12368 (N_12368,N_10850,N_11508);
nor U12369 (N_12369,N_10964,N_11536);
nand U12370 (N_12370,N_11818,N_10553);
xor U12371 (N_12371,N_11054,N_11699);
or U12372 (N_12372,N_11994,N_11167);
or U12373 (N_12373,N_10778,N_11328);
or U12374 (N_12374,N_11469,N_10635);
or U12375 (N_12375,N_11864,N_11099);
or U12376 (N_12376,N_11941,N_10803);
and U12377 (N_12377,N_11645,N_11527);
and U12378 (N_12378,N_10975,N_11741);
nor U12379 (N_12379,N_11377,N_11477);
nand U12380 (N_12380,N_11181,N_11595);
nand U12381 (N_12381,N_11857,N_11079);
and U12382 (N_12382,N_10628,N_11785);
and U12383 (N_12383,N_11243,N_11635);
nand U12384 (N_12384,N_11656,N_11117);
nand U12385 (N_12385,N_11681,N_11691);
or U12386 (N_12386,N_11378,N_11655);
or U12387 (N_12387,N_11376,N_11436);
and U12388 (N_12388,N_10540,N_11690);
xnor U12389 (N_12389,N_10834,N_11014);
nand U12390 (N_12390,N_11111,N_10634);
or U12391 (N_12391,N_11413,N_11522);
nor U12392 (N_12392,N_11212,N_11727);
nor U12393 (N_12393,N_11092,N_11608);
nand U12394 (N_12394,N_11025,N_11817);
nand U12395 (N_12395,N_11479,N_11051);
nand U12396 (N_12396,N_10518,N_10642);
or U12397 (N_12397,N_10559,N_11124);
and U12398 (N_12398,N_11130,N_11020);
and U12399 (N_12399,N_10615,N_10816);
xnor U12400 (N_12400,N_11996,N_10830);
nor U12401 (N_12401,N_11666,N_11448);
nand U12402 (N_12402,N_11713,N_11299);
nor U12403 (N_12403,N_10620,N_11821);
or U12404 (N_12404,N_11301,N_11534);
or U12405 (N_12405,N_11936,N_10917);
or U12406 (N_12406,N_10920,N_11421);
or U12407 (N_12407,N_11227,N_10990);
nor U12408 (N_12408,N_11852,N_11178);
nor U12409 (N_12409,N_10766,N_10922);
and U12410 (N_12410,N_11919,N_11966);
nand U12411 (N_12411,N_10528,N_11957);
or U12412 (N_12412,N_11922,N_11805);
or U12413 (N_12413,N_11175,N_11463);
and U12414 (N_12414,N_10602,N_10765);
and U12415 (N_12415,N_10569,N_11468);
and U12416 (N_12416,N_11582,N_11424);
nor U12417 (N_12417,N_10512,N_11141);
nand U12418 (N_12418,N_10565,N_11029);
nand U12419 (N_12419,N_10510,N_10644);
nand U12420 (N_12420,N_11485,N_10756);
or U12421 (N_12421,N_10898,N_10937);
nor U12422 (N_12422,N_11454,N_10693);
or U12423 (N_12423,N_10835,N_11844);
and U12424 (N_12424,N_11387,N_11745);
and U12425 (N_12425,N_11302,N_11947);
xnor U12426 (N_12426,N_10913,N_11680);
nor U12427 (N_12427,N_11577,N_10677);
and U12428 (N_12428,N_10949,N_11210);
nand U12429 (N_12429,N_11276,N_11845);
or U12430 (N_12430,N_11329,N_11692);
and U12431 (N_12431,N_11532,N_11991);
nand U12432 (N_12432,N_11119,N_11006);
nand U12433 (N_12433,N_11794,N_11829);
and U12434 (N_12434,N_11474,N_11886);
nor U12435 (N_12435,N_10613,N_11476);
or U12436 (N_12436,N_10825,N_11001);
xnor U12437 (N_12437,N_11399,N_11095);
nor U12438 (N_12438,N_11415,N_11726);
or U12439 (N_12439,N_10876,N_11322);
nand U12440 (N_12440,N_11230,N_10797);
or U12441 (N_12441,N_10905,N_11736);
and U12442 (N_12442,N_11895,N_11565);
and U12443 (N_12443,N_11987,N_11523);
xnor U12444 (N_12444,N_11407,N_11078);
or U12445 (N_12445,N_10554,N_11539);
and U12446 (N_12446,N_10536,N_10903);
and U12447 (N_12447,N_11990,N_10971);
xor U12448 (N_12448,N_11890,N_11074);
nand U12449 (N_12449,N_10629,N_11495);
nand U12450 (N_12450,N_11795,N_10795);
nor U12451 (N_12451,N_11878,N_11375);
and U12452 (N_12452,N_10732,N_11738);
or U12453 (N_12453,N_11122,N_11708);
nor U12454 (N_12454,N_10712,N_11312);
and U12455 (N_12455,N_10694,N_11601);
or U12456 (N_12456,N_10517,N_11083);
or U12457 (N_12457,N_11714,N_11719);
or U12458 (N_12458,N_10775,N_10503);
xor U12459 (N_12459,N_10542,N_11018);
nand U12460 (N_12460,N_11066,N_10650);
xor U12461 (N_12461,N_10577,N_10773);
nand U12462 (N_12462,N_10826,N_10895);
nor U12463 (N_12463,N_10843,N_11931);
or U12464 (N_12464,N_11590,N_11132);
nand U12465 (N_12465,N_11693,N_11183);
and U12466 (N_12466,N_10781,N_11344);
nor U12467 (N_12467,N_11316,N_11449);
or U12468 (N_12468,N_11185,N_10986);
and U12469 (N_12469,N_10925,N_11809);
nor U12470 (N_12470,N_11423,N_10918);
and U12471 (N_12471,N_10752,N_10660);
xor U12472 (N_12472,N_10790,N_11211);
nor U12473 (N_12473,N_11524,N_10926);
nand U12474 (N_12474,N_11337,N_11007);
nand U12475 (N_12475,N_10534,N_11484);
or U12476 (N_12476,N_10992,N_11203);
nand U12477 (N_12477,N_11444,N_11388);
nor U12478 (N_12478,N_11274,N_11367);
xnor U12479 (N_12479,N_10527,N_10853);
and U12480 (N_12480,N_11884,N_10533);
and U12481 (N_12481,N_10904,N_11743);
and U12482 (N_12482,N_10805,N_11372);
nand U12483 (N_12483,N_11184,N_10574);
xor U12484 (N_12484,N_10575,N_10501);
or U12485 (N_12485,N_11782,N_10967);
nand U12486 (N_12486,N_10633,N_11400);
and U12487 (N_12487,N_11342,N_11562);
nand U12488 (N_12488,N_11510,N_11135);
xnor U12489 (N_12489,N_10791,N_11968);
nand U12490 (N_12490,N_11138,N_10930);
nand U12491 (N_12491,N_11783,N_11459);
and U12492 (N_12492,N_10625,N_10637);
nor U12493 (N_12493,N_11695,N_11558);
nand U12494 (N_12494,N_11194,N_11089);
xor U12495 (N_12495,N_11116,N_10923);
and U12496 (N_12496,N_11956,N_11959);
or U12497 (N_12497,N_11867,N_11682);
nand U12498 (N_12498,N_10998,N_10699);
xnor U12499 (N_12499,N_11115,N_11492);
xor U12500 (N_12500,N_11702,N_11024);
nand U12501 (N_12501,N_10570,N_11170);
and U12502 (N_12502,N_11277,N_10870);
nor U12503 (N_12503,N_11336,N_10511);
or U12504 (N_12504,N_11218,N_11733);
or U12505 (N_12505,N_11720,N_11346);
and U12506 (N_12506,N_10883,N_11573);
nand U12507 (N_12507,N_10813,N_11787);
and U12508 (N_12508,N_11408,N_11939);
or U12509 (N_12509,N_10557,N_11295);
or U12510 (N_12510,N_11189,N_11718);
nor U12511 (N_12511,N_10664,N_10700);
or U12512 (N_12512,N_11358,N_11494);
nand U12513 (N_12513,N_10932,N_10924);
or U12514 (N_12514,N_10782,N_11225);
xnor U12515 (N_12515,N_11575,N_10954);
nor U12516 (N_12516,N_10548,N_11360);
and U12517 (N_12517,N_11820,N_11807);
and U12518 (N_12518,N_10638,N_10652);
xor U12519 (N_12519,N_11995,N_11186);
nor U12520 (N_12520,N_11742,N_11754);
and U12521 (N_12521,N_11219,N_10584);
or U12522 (N_12522,N_11977,N_10680);
or U12523 (N_12523,N_10673,N_11606);
nand U12524 (N_12524,N_11611,N_10697);
nor U12525 (N_12525,N_11511,N_11015);
nor U12526 (N_12526,N_10872,N_11552);
nand U12527 (N_12527,N_11772,N_11441);
and U12528 (N_12528,N_10737,N_11897);
and U12529 (N_12529,N_10840,N_10899);
and U12530 (N_12530,N_11973,N_10513);
nand U12531 (N_12531,N_10715,N_10951);
and U12532 (N_12532,N_10763,N_10589);
and U12533 (N_12533,N_11440,N_11858);
nand U12534 (N_12534,N_11544,N_11876);
xor U12535 (N_12535,N_11865,N_11023);
and U12536 (N_12536,N_11282,N_11671);
xnor U12537 (N_12537,N_10757,N_11244);
and U12538 (N_12538,N_10524,N_11296);
nand U12539 (N_12539,N_11457,N_11571);
or U12540 (N_12540,N_11173,N_11091);
and U12541 (N_12541,N_10799,N_10608);
xnor U12542 (N_12542,N_11497,N_11808);
nand U12543 (N_12543,N_10679,N_11615);
or U12544 (N_12544,N_11773,N_11355);
or U12545 (N_12545,N_11556,N_11153);
nor U12546 (N_12546,N_11568,N_11071);
nor U12547 (N_12547,N_10675,N_10833);
nand U12548 (N_12548,N_11053,N_11732);
or U12549 (N_12549,N_11131,N_11762);
or U12550 (N_12550,N_11637,N_10623);
nor U12551 (N_12551,N_10798,N_10836);
nand U12552 (N_12552,N_11039,N_11679);
nand U12553 (N_12553,N_11618,N_10893);
or U12554 (N_12554,N_11584,N_10862);
and U12555 (N_12555,N_11625,N_11538);
or U12556 (N_12556,N_10831,N_11786);
nand U12557 (N_12557,N_10885,N_11285);
nor U12558 (N_12558,N_11709,N_11202);
xnor U12559 (N_12559,N_11518,N_11126);
nor U12560 (N_12560,N_11326,N_11076);
and U12561 (N_12561,N_11902,N_11759);
nand U12562 (N_12562,N_11749,N_10731);
xor U12563 (N_12563,N_11545,N_11660);
nand U12564 (N_12564,N_11704,N_11438);
nand U12565 (N_12565,N_10891,N_10529);
nor U12566 (N_12566,N_11368,N_10943);
or U12567 (N_12567,N_10722,N_10878);
nor U12568 (N_12568,N_11502,N_11404);
and U12569 (N_12569,N_11222,N_11812);
nand U12570 (N_12570,N_11983,N_10547);
or U12571 (N_12571,N_11369,N_10802);
xnor U12572 (N_12572,N_11042,N_11258);
and U12573 (N_12573,N_11304,N_11410);
and U12574 (N_12574,N_11624,N_10758);
and U12575 (N_12575,N_10674,N_11240);
and U12576 (N_12576,N_11507,N_10871);
or U12577 (N_12577,N_10821,N_11259);
nand U12578 (N_12578,N_10950,N_10856);
nor U12579 (N_12579,N_11598,N_11446);
or U12580 (N_12580,N_11386,N_10566);
nand U12581 (N_12581,N_11810,N_10690);
or U12582 (N_12582,N_10723,N_11554);
nor U12583 (N_12583,N_11950,N_10892);
xnor U12584 (N_12584,N_10692,N_11949);
and U12585 (N_12585,N_11913,N_10788);
nand U12586 (N_12586,N_11294,N_11752);
and U12587 (N_12587,N_10500,N_10696);
and U12588 (N_12588,N_11874,N_10645);
or U12589 (N_12589,N_10970,N_11251);
nor U12590 (N_12590,N_11333,N_10618);
nand U12591 (N_12591,N_10810,N_11080);
and U12592 (N_12592,N_11005,N_10890);
or U12593 (N_12593,N_11953,N_11703);
and U12594 (N_12594,N_10563,N_11249);
and U12595 (N_12595,N_11663,N_10868);
nand U12596 (N_12596,N_11425,N_10587);
nand U12597 (N_12597,N_10735,N_10772);
and U12598 (N_12598,N_11685,N_11017);
xnor U12599 (N_12599,N_10882,N_11220);
or U12600 (N_12600,N_11833,N_10509);
nand U12601 (N_12601,N_10648,N_11443);
and U12602 (N_12602,N_11059,N_11361);
nor U12603 (N_12603,N_11199,N_11393);
and U12604 (N_12604,N_10596,N_11935);
and U12605 (N_12605,N_11049,N_10946);
or U12606 (N_12606,N_11796,N_11873);
and U12607 (N_12607,N_10983,N_10695);
nor U12608 (N_12608,N_10750,N_10561);
nand U12609 (N_12609,N_10865,N_11190);
nand U12610 (N_12610,N_10968,N_11221);
nand U12611 (N_12611,N_11204,N_10800);
and U12612 (N_12612,N_11748,N_11826);
or U12613 (N_12613,N_10963,N_11075);
nor U12614 (N_12614,N_10572,N_11033);
or U12615 (N_12615,N_11364,N_11389);
nand U12616 (N_12616,N_10657,N_11866);
nand U12617 (N_12617,N_11451,N_11513);
nor U12618 (N_12618,N_11610,N_10780);
or U12619 (N_12619,N_11458,N_11622);
and U12620 (N_12620,N_10666,N_11320);
and U12621 (N_12621,N_11770,N_10754);
and U12622 (N_12622,N_10947,N_10827);
nor U12623 (N_12623,N_11697,N_11002);
and U12624 (N_12624,N_11319,N_11192);
nand U12625 (N_12625,N_10936,N_11944);
and U12626 (N_12626,N_11602,N_11801);
nand U12627 (N_12627,N_10659,N_11687);
or U12628 (N_12628,N_10828,N_10525);
or U12629 (N_12629,N_10746,N_11077);
nand U12630 (N_12630,N_11090,N_11107);
nand U12631 (N_12631,N_11880,N_11825);
nor U12632 (N_12632,N_11550,N_10769);
nand U12633 (N_12633,N_11767,N_11586);
nand U12634 (N_12634,N_11309,N_10721);
xnor U12635 (N_12635,N_11832,N_11648);
or U12636 (N_12636,N_10555,N_11587);
or U12637 (N_12637,N_11955,N_10537);
xor U12638 (N_12638,N_11182,N_10948);
and U12639 (N_12639,N_11161,N_11658);
or U12640 (N_12640,N_10519,N_11771);
nand U12641 (N_12641,N_11673,N_11390);
and U12642 (N_12642,N_11255,N_11281);
nand U12643 (N_12643,N_10955,N_11964);
nor U12644 (N_12644,N_10928,N_11123);
and U12645 (N_12645,N_10564,N_11268);
nor U12646 (N_12646,N_11863,N_11349);
and U12647 (N_12647,N_11417,N_11758);
nor U12648 (N_12648,N_10824,N_11208);
and U12649 (N_12649,N_11910,N_11260);
and U12650 (N_12650,N_11356,N_10940);
and U12651 (N_12651,N_11667,N_11348);
and U12652 (N_12652,N_10748,N_11855);
nand U12653 (N_12653,N_10617,N_10962);
xnor U12654 (N_12654,N_11909,N_10807);
nor U12655 (N_12655,N_11970,N_10708);
nand U12656 (N_12656,N_11986,N_11098);
or U12657 (N_12657,N_11698,N_11343);
nand U12658 (N_12658,N_11547,N_11307);
and U12659 (N_12659,N_11351,N_11021);
xnor U12660 (N_12660,N_10774,N_10604);
nand U12661 (N_12661,N_11688,N_10919);
nor U12662 (N_12662,N_10607,N_11517);
or U12663 (N_12663,N_11300,N_10724);
or U12664 (N_12664,N_11426,N_11694);
or U12665 (N_12665,N_10741,N_10966);
nand U12666 (N_12666,N_11401,N_10646);
nand U12667 (N_12667,N_11345,N_11912);
and U12668 (N_12668,N_11085,N_11537);
and U12669 (N_12669,N_11332,N_10820);
or U12670 (N_12670,N_11559,N_11000);
or U12671 (N_12671,N_10612,N_11031);
and U12672 (N_12672,N_11201,N_10688);
nor U12673 (N_12673,N_11315,N_11851);
nor U12674 (N_12674,N_11715,N_11784);
and U12675 (N_12675,N_11737,N_11250);
or U12676 (N_12676,N_11597,N_11612);
or U12677 (N_12677,N_11888,N_10981);
nand U12678 (N_12678,N_10881,N_11462);
and U12679 (N_12679,N_11370,N_11563);
or U12680 (N_12680,N_10504,N_10530);
or U12681 (N_12681,N_11490,N_11120);
nor U12682 (N_12682,N_10927,N_11779);
or U12683 (N_12683,N_11297,N_11422);
and U12684 (N_12684,N_10626,N_10727);
and U12685 (N_12685,N_11609,N_11171);
nand U12686 (N_12686,N_11802,N_11403);
nand U12687 (N_12687,N_11102,N_11215);
and U12688 (N_12688,N_10997,N_11406);
or U12689 (N_12689,N_11963,N_11321);
nor U12690 (N_12690,N_11757,N_10956);
or U12691 (N_12691,N_11617,N_11764);
xnor U12692 (N_12692,N_10665,N_10979);
or U12693 (N_12693,N_11653,N_11799);
and U12694 (N_12694,N_11892,N_11056);
nand U12695 (N_12695,N_11765,N_11187);
nor U12696 (N_12696,N_10817,N_11151);
or U12697 (N_12697,N_11050,N_10720);
nand U12698 (N_12698,N_11721,N_11604);
nand U12699 (N_12699,N_10888,N_11103);
or U12700 (N_12700,N_11634,N_11235);
nor U12701 (N_12701,N_10581,N_11037);
or U12702 (N_12702,N_11262,N_11450);
and U12703 (N_12703,N_11373,N_11659);
nor U12704 (N_12704,N_11677,N_11835);
nor U12705 (N_12705,N_11165,N_10929);
nor U12706 (N_12706,N_11907,N_11638);
nand U12707 (N_12707,N_11908,N_11248);
or U12708 (N_12708,N_11068,N_11061);
xor U12709 (N_12709,N_11087,N_10717);
or U12710 (N_12710,N_11082,N_11394);
nor U12711 (N_12711,N_10702,N_11013);
or U12712 (N_12712,N_11628,N_11505);
nand U12713 (N_12713,N_11967,N_11989);
and U12714 (N_12714,N_11456,N_10521);
nor U12715 (N_12715,N_10938,N_11180);
and U12716 (N_12716,N_11885,N_11177);
or U12717 (N_12717,N_10784,N_11943);
nor U12718 (N_12718,N_11445,N_11519);
and U12719 (N_12719,N_11283,N_11921);
nand U12720 (N_12720,N_10726,N_11668);
nand U12721 (N_12721,N_11791,N_10886);
and U12722 (N_12722,N_11331,N_11308);
nor U12723 (N_12723,N_10852,N_11940);
or U12724 (N_12724,N_11447,N_11318);
nor U12725 (N_12725,N_10627,N_11992);
xor U12726 (N_12726,N_11958,N_11144);
nor U12727 (N_12727,N_11269,N_11136);
nand U12728 (N_12728,N_11140,N_11383);
nand U12729 (N_12729,N_11834,N_10985);
xnor U12730 (N_12730,N_11566,N_10896);
nand U12731 (N_12731,N_10931,N_10759);
nor U12732 (N_12732,N_10683,N_11209);
nand U12733 (N_12733,N_11847,N_11998);
xnor U12734 (N_12734,N_10558,N_11482);
or U12735 (N_12735,N_11529,N_10656);
nand U12736 (N_12736,N_10777,N_11246);
or U12737 (N_12737,N_11188,N_11498);
or U12738 (N_12738,N_11063,N_11898);
nor U12739 (N_12739,N_10976,N_10568);
and U12740 (N_12740,N_11870,N_11164);
or U12741 (N_12741,N_11626,N_11019);
and U12742 (N_12742,N_11901,N_11933);
or U12743 (N_12743,N_10729,N_10867);
nor U12744 (N_12744,N_10562,N_11392);
xnor U12745 (N_12745,N_11840,N_11195);
and U12746 (N_12746,N_10661,N_11247);
and U12747 (N_12747,N_10594,N_11411);
nand U12748 (N_12748,N_10875,N_10531);
nor U12749 (N_12749,N_11439,N_11148);
nor U12750 (N_12750,N_11907,N_10699);
nand U12751 (N_12751,N_11031,N_11064);
nand U12752 (N_12752,N_10971,N_11126);
or U12753 (N_12753,N_11012,N_11639);
or U12754 (N_12754,N_11663,N_10855);
xnor U12755 (N_12755,N_11656,N_11399);
xnor U12756 (N_12756,N_11056,N_11682);
nor U12757 (N_12757,N_11614,N_10896);
and U12758 (N_12758,N_11235,N_11827);
or U12759 (N_12759,N_10572,N_11387);
or U12760 (N_12760,N_11154,N_10586);
nor U12761 (N_12761,N_11317,N_11408);
nand U12762 (N_12762,N_11071,N_11016);
xor U12763 (N_12763,N_11951,N_10537);
nand U12764 (N_12764,N_11606,N_10866);
and U12765 (N_12765,N_11182,N_10601);
and U12766 (N_12766,N_11654,N_11740);
xnor U12767 (N_12767,N_11528,N_11986);
nor U12768 (N_12768,N_10541,N_11800);
nor U12769 (N_12769,N_10730,N_10736);
nor U12770 (N_12770,N_11928,N_10846);
and U12771 (N_12771,N_11634,N_11932);
or U12772 (N_12772,N_10979,N_11369);
or U12773 (N_12773,N_11139,N_11886);
nor U12774 (N_12774,N_10691,N_11985);
or U12775 (N_12775,N_11888,N_11216);
and U12776 (N_12776,N_11601,N_11667);
nand U12777 (N_12777,N_11873,N_10666);
nor U12778 (N_12778,N_11970,N_11155);
nand U12779 (N_12779,N_10824,N_11087);
and U12780 (N_12780,N_11305,N_11174);
nor U12781 (N_12781,N_10554,N_11845);
and U12782 (N_12782,N_10639,N_11937);
nand U12783 (N_12783,N_10708,N_10687);
or U12784 (N_12784,N_11381,N_10653);
nor U12785 (N_12785,N_11819,N_11380);
and U12786 (N_12786,N_11089,N_11877);
nand U12787 (N_12787,N_10635,N_11719);
xnor U12788 (N_12788,N_11136,N_11344);
nor U12789 (N_12789,N_11879,N_11340);
nor U12790 (N_12790,N_11603,N_11574);
nand U12791 (N_12791,N_11454,N_10873);
xor U12792 (N_12792,N_10630,N_11455);
and U12793 (N_12793,N_11989,N_11699);
nor U12794 (N_12794,N_11023,N_10845);
nand U12795 (N_12795,N_11667,N_10631);
xnor U12796 (N_12796,N_10670,N_11783);
and U12797 (N_12797,N_10990,N_11949);
and U12798 (N_12798,N_11991,N_10747);
nand U12799 (N_12799,N_10645,N_11116);
or U12800 (N_12800,N_11564,N_11505);
and U12801 (N_12801,N_10964,N_11465);
and U12802 (N_12802,N_11028,N_10877);
or U12803 (N_12803,N_10758,N_10825);
nand U12804 (N_12804,N_10789,N_10719);
nor U12805 (N_12805,N_11021,N_10627);
or U12806 (N_12806,N_10640,N_11951);
and U12807 (N_12807,N_11582,N_11741);
or U12808 (N_12808,N_10755,N_11004);
nor U12809 (N_12809,N_11828,N_10560);
and U12810 (N_12810,N_10688,N_11954);
or U12811 (N_12811,N_11335,N_11317);
or U12812 (N_12812,N_11763,N_10646);
and U12813 (N_12813,N_10900,N_10591);
or U12814 (N_12814,N_11075,N_11647);
and U12815 (N_12815,N_10951,N_11233);
nand U12816 (N_12816,N_10620,N_11074);
and U12817 (N_12817,N_11252,N_11631);
or U12818 (N_12818,N_11273,N_10890);
nor U12819 (N_12819,N_10972,N_11128);
nor U12820 (N_12820,N_11071,N_10586);
xnor U12821 (N_12821,N_10566,N_11606);
or U12822 (N_12822,N_11458,N_11875);
and U12823 (N_12823,N_11391,N_11764);
and U12824 (N_12824,N_11733,N_11193);
or U12825 (N_12825,N_10801,N_11362);
or U12826 (N_12826,N_11764,N_11707);
nand U12827 (N_12827,N_10829,N_11130);
nand U12828 (N_12828,N_11587,N_10855);
nand U12829 (N_12829,N_11540,N_11088);
or U12830 (N_12830,N_11424,N_11893);
or U12831 (N_12831,N_11775,N_11086);
xnor U12832 (N_12832,N_11606,N_10572);
nand U12833 (N_12833,N_11956,N_10929);
nand U12834 (N_12834,N_11779,N_10632);
nand U12835 (N_12835,N_11214,N_11387);
nand U12836 (N_12836,N_11024,N_10561);
or U12837 (N_12837,N_11505,N_11898);
and U12838 (N_12838,N_11326,N_10931);
or U12839 (N_12839,N_10807,N_11817);
or U12840 (N_12840,N_11510,N_11294);
or U12841 (N_12841,N_11811,N_11434);
nand U12842 (N_12842,N_11666,N_10604);
nor U12843 (N_12843,N_11983,N_10866);
or U12844 (N_12844,N_11505,N_10953);
or U12845 (N_12845,N_11973,N_10794);
and U12846 (N_12846,N_11489,N_11351);
and U12847 (N_12847,N_11713,N_10769);
xor U12848 (N_12848,N_10868,N_11950);
xnor U12849 (N_12849,N_11960,N_11237);
or U12850 (N_12850,N_10893,N_11449);
xor U12851 (N_12851,N_11013,N_11879);
nor U12852 (N_12852,N_11456,N_11554);
or U12853 (N_12853,N_11719,N_10700);
or U12854 (N_12854,N_10575,N_10918);
nand U12855 (N_12855,N_10761,N_10949);
xnor U12856 (N_12856,N_11014,N_11803);
nand U12857 (N_12857,N_11493,N_11204);
or U12858 (N_12858,N_10721,N_10612);
or U12859 (N_12859,N_10661,N_10729);
or U12860 (N_12860,N_11489,N_10863);
or U12861 (N_12861,N_11502,N_10862);
nor U12862 (N_12862,N_11026,N_10674);
nor U12863 (N_12863,N_10534,N_11531);
and U12864 (N_12864,N_11142,N_11982);
nand U12865 (N_12865,N_11734,N_11338);
nand U12866 (N_12866,N_11769,N_11976);
xnor U12867 (N_12867,N_11815,N_10759);
xor U12868 (N_12868,N_11851,N_11618);
and U12869 (N_12869,N_11036,N_11157);
and U12870 (N_12870,N_11845,N_11510);
nand U12871 (N_12871,N_10619,N_11856);
nand U12872 (N_12872,N_10782,N_11884);
nand U12873 (N_12873,N_11206,N_10606);
nand U12874 (N_12874,N_10544,N_11371);
nor U12875 (N_12875,N_11211,N_11412);
xor U12876 (N_12876,N_10529,N_11741);
nand U12877 (N_12877,N_10956,N_11449);
nor U12878 (N_12878,N_10927,N_11595);
and U12879 (N_12879,N_11799,N_11154);
and U12880 (N_12880,N_10991,N_11242);
nand U12881 (N_12881,N_11253,N_11512);
nand U12882 (N_12882,N_10921,N_10657);
and U12883 (N_12883,N_11538,N_10669);
nand U12884 (N_12884,N_11944,N_11070);
nand U12885 (N_12885,N_11482,N_11972);
or U12886 (N_12886,N_10622,N_11031);
and U12887 (N_12887,N_10929,N_10799);
nor U12888 (N_12888,N_10665,N_11356);
and U12889 (N_12889,N_10903,N_10893);
and U12890 (N_12890,N_10629,N_11505);
nand U12891 (N_12891,N_11719,N_11145);
nand U12892 (N_12892,N_11338,N_10508);
nand U12893 (N_12893,N_11325,N_11735);
nor U12894 (N_12894,N_11401,N_11353);
or U12895 (N_12895,N_11551,N_11357);
nor U12896 (N_12896,N_11823,N_11974);
and U12897 (N_12897,N_11455,N_11391);
nor U12898 (N_12898,N_10655,N_10537);
or U12899 (N_12899,N_11239,N_10876);
nand U12900 (N_12900,N_10917,N_10507);
xor U12901 (N_12901,N_10736,N_11862);
nor U12902 (N_12902,N_11151,N_10680);
or U12903 (N_12903,N_11714,N_11005);
nand U12904 (N_12904,N_11866,N_11070);
nor U12905 (N_12905,N_11268,N_11899);
nor U12906 (N_12906,N_11221,N_11767);
nand U12907 (N_12907,N_11038,N_11079);
and U12908 (N_12908,N_10735,N_10675);
nand U12909 (N_12909,N_11161,N_11522);
xnor U12910 (N_12910,N_11190,N_10568);
nor U12911 (N_12911,N_10895,N_10897);
and U12912 (N_12912,N_11000,N_11370);
xnor U12913 (N_12913,N_11963,N_11611);
or U12914 (N_12914,N_11976,N_11921);
and U12915 (N_12915,N_11228,N_10851);
or U12916 (N_12916,N_11099,N_10669);
and U12917 (N_12917,N_11423,N_10694);
xor U12918 (N_12918,N_10760,N_11303);
nand U12919 (N_12919,N_11065,N_10658);
or U12920 (N_12920,N_11893,N_11938);
nor U12921 (N_12921,N_10955,N_10872);
or U12922 (N_12922,N_11866,N_10589);
and U12923 (N_12923,N_11023,N_10647);
nor U12924 (N_12924,N_11603,N_11646);
nor U12925 (N_12925,N_10849,N_10694);
or U12926 (N_12926,N_11238,N_10629);
nand U12927 (N_12927,N_11719,N_11903);
and U12928 (N_12928,N_10792,N_11659);
nand U12929 (N_12929,N_11298,N_11938);
and U12930 (N_12930,N_11380,N_10797);
nor U12931 (N_12931,N_11194,N_11440);
or U12932 (N_12932,N_11969,N_10729);
and U12933 (N_12933,N_10581,N_10526);
nand U12934 (N_12934,N_11622,N_10695);
xor U12935 (N_12935,N_11132,N_11121);
or U12936 (N_12936,N_11123,N_10593);
or U12937 (N_12937,N_11614,N_10972);
or U12938 (N_12938,N_10614,N_10519);
or U12939 (N_12939,N_10867,N_11705);
nand U12940 (N_12940,N_11368,N_11750);
nor U12941 (N_12941,N_10972,N_11315);
and U12942 (N_12942,N_11087,N_11940);
or U12943 (N_12943,N_11356,N_11146);
nand U12944 (N_12944,N_11604,N_11314);
or U12945 (N_12945,N_11582,N_11413);
and U12946 (N_12946,N_11710,N_11469);
and U12947 (N_12947,N_11981,N_11026);
and U12948 (N_12948,N_11430,N_11746);
xnor U12949 (N_12949,N_10838,N_11258);
nor U12950 (N_12950,N_11154,N_11943);
xor U12951 (N_12951,N_10997,N_11699);
and U12952 (N_12952,N_11904,N_11240);
nand U12953 (N_12953,N_11598,N_10705);
or U12954 (N_12954,N_10638,N_11874);
nand U12955 (N_12955,N_11224,N_11814);
nor U12956 (N_12956,N_10789,N_11289);
nand U12957 (N_12957,N_10617,N_10804);
or U12958 (N_12958,N_11903,N_11217);
and U12959 (N_12959,N_11724,N_11885);
nand U12960 (N_12960,N_11100,N_11214);
xor U12961 (N_12961,N_11591,N_11360);
or U12962 (N_12962,N_11496,N_10556);
or U12963 (N_12963,N_11207,N_11911);
or U12964 (N_12964,N_10816,N_10811);
or U12965 (N_12965,N_11075,N_11233);
nand U12966 (N_12966,N_11147,N_11315);
nand U12967 (N_12967,N_11621,N_10900);
xor U12968 (N_12968,N_11411,N_11763);
nor U12969 (N_12969,N_11842,N_11402);
nor U12970 (N_12970,N_11556,N_11193);
nor U12971 (N_12971,N_10715,N_11037);
nand U12972 (N_12972,N_10794,N_10512);
or U12973 (N_12973,N_11055,N_10889);
or U12974 (N_12974,N_11110,N_11323);
xor U12975 (N_12975,N_11884,N_10646);
xnor U12976 (N_12976,N_11004,N_11347);
nand U12977 (N_12977,N_11820,N_11016);
xnor U12978 (N_12978,N_10592,N_11243);
xnor U12979 (N_12979,N_10705,N_11851);
or U12980 (N_12980,N_10946,N_11913);
nand U12981 (N_12981,N_11331,N_10734);
nand U12982 (N_12982,N_11925,N_10596);
nand U12983 (N_12983,N_11413,N_11950);
or U12984 (N_12984,N_11140,N_10733);
or U12985 (N_12985,N_11869,N_11598);
nand U12986 (N_12986,N_11479,N_11031);
and U12987 (N_12987,N_10738,N_10923);
or U12988 (N_12988,N_10562,N_10956);
xnor U12989 (N_12989,N_11769,N_10690);
or U12990 (N_12990,N_10624,N_11187);
and U12991 (N_12991,N_11293,N_11666);
nor U12992 (N_12992,N_10554,N_10805);
and U12993 (N_12993,N_11681,N_11526);
nor U12994 (N_12994,N_10727,N_10604);
nand U12995 (N_12995,N_10734,N_11379);
or U12996 (N_12996,N_10590,N_11740);
or U12997 (N_12997,N_11455,N_10742);
nand U12998 (N_12998,N_10927,N_11671);
nor U12999 (N_12999,N_11631,N_10631);
nand U13000 (N_13000,N_10612,N_11903);
nand U13001 (N_13001,N_11786,N_10776);
nor U13002 (N_13002,N_11910,N_11078);
nand U13003 (N_13003,N_11531,N_11244);
nor U13004 (N_13004,N_11279,N_11813);
nor U13005 (N_13005,N_10746,N_10560);
nor U13006 (N_13006,N_11101,N_11924);
nor U13007 (N_13007,N_10871,N_11140);
or U13008 (N_13008,N_11743,N_11447);
nand U13009 (N_13009,N_11161,N_11324);
xor U13010 (N_13010,N_11737,N_11491);
and U13011 (N_13011,N_11396,N_10694);
nand U13012 (N_13012,N_11296,N_10515);
or U13013 (N_13013,N_11073,N_10750);
nor U13014 (N_13014,N_11509,N_11485);
xnor U13015 (N_13015,N_11261,N_11015);
or U13016 (N_13016,N_11518,N_11940);
nor U13017 (N_13017,N_10819,N_11402);
or U13018 (N_13018,N_11012,N_10981);
and U13019 (N_13019,N_10918,N_11120);
and U13020 (N_13020,N_11936,N_11358);
nor U13021 (N_13021,N_10664,N_10774);
and U13022 (N_13022,N_11026,N_11268);
nand U13023 (N_13023,N_10740,N_11981);
nand U13024 (N_13024,N_11316,N_11532);
and U13025 (N_13025,N_11176,N_11107);
and U13026 (N_13026,N_11205,N_11310);
or U13027 (N_13027,N_11421,N_11582);
nand U13028 (N_13028,N_11564,N_10717);
or U13029 (N_13029,N_11433,N_11298);
nand U13030 (N_13030,N_10580,N_11290);
and U13031 (N_13031,N_11816,N_10995);
xor U13032 (N_13032,N_11124,N_11997);
and U13033 (N_13033,N_10560,N_11203);
xnor U13034 (N_13034,N_11260,N_11639);
nor U13035 (N_13035,N_10842,N_11450);
nand U13036 (N_13036,N_10666,N_11799);
nand U13037 (N_13037,N_10701,N_11276);
nand U13038 (N_13038,N_11039,N_10596);
and U13039 (N_13039,N_11851,N_10964);
or U13040 (N_13040,N_11847,N_11646);
nand U13041 (N_13041,N_10600,N_11965);
or U13042 (N_13042,N_11075,N_11320);
or U13043 (N_13043,N_11583,N_11935);
and U13044 (N_13044,N_11044,N_11494);
or U13045 (N_13045,N_11587,N_11930);
nand U13046 (N_13046,N_11976,N_11937);
nand U13047 (N_13047,N_10789,N_11291);
and U13048 (N_13048,N_10727,N_11652);
nor U13049 (N_13049,N_11445,N_11651);
nor U13050 (N_13050,N_11770,N_11234);
nor U13051 (N_13051,N_11394,N_10745);
nor U13052 (N_13052,N_10583,N_11714);
nand U13053 (N_13053,N_10508,N_10962);
or U13054 (N_13054,N_11797,N_10623);
and U13055 (N_13055,N_10892,N_10511);
xnor U13056 (N_13056,N_11241,N_11429);
nand U13057 (N_13057,N_10870,N_11244);
nor U13058 (N_13058,N_11009,N_11691);
nor U13059 (N_13059,N_11524,N_10790);
nand U13060 (N_13060,N_10601,N_10761);
or U13061 (N_13061,N_11906,N_11395);
xor U13062 (N_13062,N_10994,N_11130);
nand U13063 (N_13063,N_11559,N_11638);
and U13064 (N_13064,N_11459,N_10987);
and U13065 (N_13065,N_10902,N_11303);
or U13066 (N_13066,N_11358,N_10585);
nand U13067 (N_13067,N_11584,N_11737);
nor U13068 (N_13068,N_11066,N_10533);
or U13069 (N_13069,N_11201,N_11007);
xnor U13070 (N_13070,N_11040,N_11623);
xnor U13071 (N_13071,N_11552,N_11769);
nor U13072 (N_13072,N_11305,N_11594);
and U13073 (N_13073,N_11579,N_11583);
nand U13074 (N_13074,N_11843,N_10803);
and U13075 (N_13075,N_11312,N_11905);
and U13076 (N_13076,N_11761,N_10548);
nand U13077 (N_13077,N_11588,N_11624);
nand U13078 (N_13078,N_11064,N_10679);
or U13079 (N_13079,N_11466,N_11162);
or U13080 (N_13080,N_10687,N_10593);
and U13081 (N_13081,N_11217,N_10897);
nor U13082 (N_13082,N_11158,N_10543);
and U13083 (N_13083,N_11539,N_11754);
nand U13084 (N_13084,N_10803,N_11755);
or U13085 (N_13085,N_10840,N_11133);
nand U13086 (N_13086,N_10704,N_11666);
or U13087 (N_13087,N_10662,N_11668);
xor U13088 (N_13088,N_11673,N_11383);
or U13089 (N_13089,N_11406,N_11438);
or U13090 (N_13090,N_11644,N_10944);
and U13091 (N_13091,N_10862,N_10550);
nor U13092 (N_13092,N_10768,N_11594);
nand U13093 (N_13093,N_11514,N_11065);
nor U13094 (N_13094,N_11016,N_11611);
or U13095 (N_13095,N_11842,N_11041);
nor U13096 (N_13096,N_10920,N_11625);
and U13097 (N_13097,N_11276,N_11984);
or U13098 (N_13098,N_10567,N_10509);
nor U13099 (N_13099,N_11144,N_10907);
nand U13100 (N_13100,N_11011,N_10548);
xnor U13101 (N_13101,N_10986,N_11276);
and U13102 (N_13102,N_11667,N_11999);
nand U13103 (N_13103,N_11087,N_10535);
nor U13104 (N_13104,N_11773,N_11302);
nand U13105 (N_13105,N_11015,N_11218);
xor U13106 (N_13106,N_11531,N_11550);
or U13107 (N_13107,N_11595,N_11169);
nor U13108 (N_13108,N_10543,N_11685);
and U13109 (N_13109,N_10998,N_11677);
and U13110 (N_13110,N_11305,N_10555);
and U13111 (N_13111,N_10765,N_11543);
nor U13112 (N_13112,N_11167,N_10981);
or U13113 (N_13113,N_10872,N_11378);
and U13114 (N_13114,N_10953,N_10724);
nand U13115 (N_13115,N_11888,N_11767);
nand U13116 (N_13116,N_11522,N_11875);
nor U13117 (N_13117,N_10936,N_11494);
nand U13118 (N_13118,N_11711,N_11927);
nor U13119 (N_13119,N_11253,N_11333);
nand U13120 (N_13120,N_11014,N_10926);
and U13121 (N_13121,N_10765,N_10638);
or U13122 (N_13122,N_10755,N_11378);
nand U13123 (N_13123,N_10754,N_11983);
xor U13124 (N_13124,N_10612,N_11106);
xnor U13125 (N_13125,N_10862,N_10974);
nor U13126 (N_13126,N_11621,N_10881);
or U13127 (N_13127,N_11320,N_11603);
and U13128 (N_13128,N_11143,N_11569);
or U13129 (N_13129,N_10574,N_11237);
nand U13130 (N_13130,N_11146,N_11168);
or U13131 (N_13131,N_11480,N_10982);
and U13132 (N_13132,N_11356,N_10786);
nor U13133 (N_13133,N_10948,N_11066);
nand U13134 (N_13134,N_10513,N_10705);
nor U13135 (N_13135,N_11286,N_11828);
or U13136 (N_13136,N_11226,N_11432);
nor U13137 (N_13137,N_10981,N_11638);
xor U13138 (N_13138,N_11735,N_10813);
nand U13139 (N_13139,N_10509,N_11495);
nand U13140 (N_13140,N_11285,N_11123);
or U13141 (N_13141,N_10542,N_10690);
nand U13142 (N_13142,N_10597,N_10803);
or U13143 (N_13143,N_11009,N_11556);
nand U13144 (N_13144,N_11851,N_11756);
xnor U13145 (N_13145,N_11405,N_10619);
or U13146 (N_13146,N_11908,N_11975);
nor U13147 (N_13147,N_10768,N_11666);
xor U13148 (N_13148,N_11038,N_10565);
nand U13149 (N_13149,N_11252,N_11651);
nand U13150 (N_13150,N_11892,N_11274);
xor U13151 (N_13151,N_11607,N_11817);
nand U13152 (N_13152,N_11969,N_10706);
and U13153 (N_13153,N_11466,N_11308);
or U13154 (N_13154,N_11152,N_10649);
nand U13155 (N_13155,N_10929,N_11844);
and U13156 (N_13156,N_11717,N_11547);
or U13157 (N_13157,N_11769,N_11229);
or U13158 (N_13158,N_10582,N_11357);
nor U13159 (N_13159,N_10552,N_11023);
or U13160 (N_13160,N_10662,N_10770);
nand U13161 (N_13161,N_11239,N_10631);
xnor U13162 (N_13162,N_11533,N_11441);
or U13163 (N_13163,N_10644,N_11430);
and U13164 (N_13164,N_10824,N_10756);
xnor U13165 (N_13165,N_11514,N_11679);
and U13166 (N_13166,N_10910,N_11656);
and U13167 (N_13167,N_11401,N_10776);
or U13168 (N_13168,N_11245,N_10504);
nor U13169 (N_13169,N_11236,N_11900);
nor U13170 (N_13170,N_10978,N_11400);
nand U13171 (N_13171,N_10730,N_11445);
and U13172 (N_13172,N_11960,N_11950);
nor U13173 (N_13173,N_11646,N_11936);
and U13174 (N_13174,N_10652,N_11273);
or U13175 (N_13175,N_11014,N_10558);
or U13176 (N_13176,N_10577,N_11455);
nand U13177 (N_13177,N_11488,N_11704);
and U13178 (N_13178,N_11370,N_11233);
or U13179 (N_13179,N_11281,N_11925);
and U13180 (N_13180,N_10921,N_11294);
or U13181 (N_13181,N_10619,N_10797);
and U13182 (N_13182,N_11921,N_11263);
nand U13183 (N_13183,N_11277,N_10834);
or U13184 (N_13184,N_10938,N_11191);
and U13185 (N_13185,N_11771,N_11378);
nor U13186 (N_13186,N_10602,N_11447);
and U13187 (N_13187,N_10915,N_11655);
nor U13188 (N_13188,N_11161,N_10635);
or U13189 (N_13189,N_10770,N_10843);
nor U13190 (N_13190,N_11759,N_10557);
nand U13191 (N_13191,N_11141,N_10694);
nand U13192 (N_13192,N_11946,N_11883);
and U13193 (N_13193,N_11918,N_10615);
nand U13194 (N_13194,N_10685,N_11388);
nand U13195 (N_13195,N_11460,N_11533);
or U13196 (N_13196,N_11944,N_10993);
nor U13197 (N_13197,N_10544,N_11378);
or U13198 (N_13198,N_10617,N_10774);
xor U13199 (N_13199,N_10634,N_11943);
nand U13200 (N_13200,N_11907,N_11343);
and U13201 (N_13201,N_11443,N_11744);
nand U13202 (N_13202,N_11775,N_10707);
nand U13203 (N_13203,N_10745,N_11817);
nor U13204 (N_13204,N_11178,N_10758);
and U13205 (N_13205,N_11987,N_11058);
nor U13206 (N_13206,N_10821,N_11945);
and U13207 (N_13207,N_11684,N_11353);
nand U13208 (N_13208,N_11832,N_10753);
and U13209 (N_13209,N_11769,N_11322);
and U13210 (N_13210,N_11569,N_11220);
or U13211 (N_13211,N_10759,N_11489);
or U13212 (N_13212,N_10963,N_10970);
nand U13213 (N_13213,N_11836,N_10501);
nand U13214 (N_13214,N_10813,N_10767);
and U13215 (N_13215,N_10510,N_11027);
and U13216 (N_13216,N_10948,N_11134);
or U13217 (N_13217,N_11495,N_11878);
nand U13218 (N_13218,N_10956,N_11289);
or U13219 (N_13219,N_10718,N_11409);
or U13220 (N_13220,N_10677,N_11781);
nand U13221 (N_13221,N_10632,N_10752);
or U13222 (N_13222,N_10872,N_11809);
xnor U13223 (N_13223,N_11139,N_11792);
and U13224 (N_13224,N_10695,N_10616);
xnor U13225 (N_13225,N_11828,N_11086);
nor U13226 (N_13226,N_11058,N_11264);
or U13227 (N_13227,N_11923,N_11633);
and U13228 (N_13228,N_11230,N_11922);
xor U13229 (N_13229,N_11544,N_11805);
and U13230 (N_13230,N_11060,N_11801);
and U13231 (N_13231,N_10852,N_11403);
nand U13232 (N_13232,N_11754,N_11018);
nor U13233 (N_13233,N_11503,N_11174);
nor U13234 (N_13234,N_11065,N_11942);
nand U13235 (N_13235,N_11623,N_11586);
and U13236 (N_13236,N_11330,N_10645);
xnor U13237 (N_13237,N_11304,N_10556);
nor U13238 (N_13238,N_10758,N_10540);
or U13239 (N_13239,N_11332,N_11499);
xor U13240 (N_13240,N_11013,N_10510);
and U13241 (N_13241,N_11849,N_11101);
nand U13242 (N_13242,N_11709,N_11936);
xor U13243 (N_13243,N_11131,N_10807);
nand U13244 (N_13244,N_10739,N_11029);
nand U13245 (N_13245,N_11132,N_10988);
nand U13246 (N_13246,N_10538,N_10602);
or U13247 (N_13247,N_10890,N_11198);
and U13248 (N_13248,N_11039,N_10942);
or U13249 (N_13249,N_10812,N_11811);
and U13250 (N_13250,N_11614,N_11405);
and U13251 (N_13251,N_11564,N_11529);
and U13252 (N_13252,N_11281,N_10827);
and U13253 (N_13253,N_11402,N_11580);
and U13254 (N_13254,N_10888,N_11466);
or U13255 (N_13255,N_11317,N_11176);
nor U13256 (N_13256,N_11249,N_10636);
nor U13257 (N_13257,N_10508,N_11628);
or U13258 (N_13258,N_10672,N_10983);
and U13259 (N_13259,N_11566,N_11224);
nand U13260 (N_13260,N_11053,N_11275);
nor U13261 (N_13261,N_11123,N_11716);
nand U13262 (N_13262,N_11163,N_11194);
nor U13263 (N_13263,N_11752,N_10506);
nor U13264 (N_13264,N_11752,N_10897);
nor U13265 (N_13265,N_11595,N_11380);
nand U13266 (N_13266,N_11566,N_10521);
nor U13267 (N_13267,N_10751,N_11398);
nand U13268 (N_13268,N_11096,N_11323);
xnor U13269 (N_13269,N_11071,N_10836);
and U13270 (N_13270,N_10835,N_10792);
and U13271 (N_13271,N_11191,N_10511);
or U13272 (N_13272,N_11068,N_11414);
and U13273 (N_13273,N_11550,N_10974);
nand U13274 (N_13274,N_10515,N_11675);
nor U13275 (N_13275,N_11388,N_11849);
xor U13276 (N_13276,N_11751,N_10860);
or U13277 (N_13277,N_11262,N_11785);
xnor U13278 (N_13278,N_11653,N_11245);
or U13279 (N_13279,N_11805,N_10534);
nor U13280 (N_13280,N_10980,N_11751);
or U13281 (N_13281,N_10776,N_11356);
xnor U13282 (N_13282,N_11550,N_11949);
nor U13283 (N_13283,N_11752,N_11087);
nor U13284 (N_13284,N_11567,N_11702);
and U13285 (N_13285,N_11094,N_10621);
and U13286 (N_13286,N_10756,N_11153);
or U13287 (N_13287,N_11947,N_11156);
nor U13288 (N_13288,N_11028,N_11292);
or U13289 (N_13289,N_10851,N_11251);
and U13290 (N_13290,N_10699,N_10562);
and U13291 (N_13291,N_11382,N_10870);
nor U13292 (N_13292,N_10857,N_11593);
nor U13293 (N_13293,N_11693,N_11050);
nor U13294 (N_13294,N_11098,N_10760);
nor U13295 (N_13295,N_11462,N_11623);
and U13296 (N_13296,N_11456,N_11103);
nor U13297 (N_13297,N_11274,N_11500);
or U13298 (N_13298,N_10813,N_11218);
and U13299 (N_13299,N_11937,N_11115);
nor U13300 (N_13300,N_11334,N_10825);
nand U13301 (N_13301,N_10890,N_11913);
xnor U13302 (N_13302,N_10616,N_11602);
nor U13303 (N_13303,N_10944,N_10876);
or U13304 (N_13304,N_11340,N_11031);
nand U13305 (N_13305,N_10957,N_11949);
or U13306 (N_13306,N_10800,N_10830);
nand U13307 (N_13307,N_11809,N_11105);
or U13308 (N_13308,N_11950,N_10649);
and U13309 (N_13309,N_11274,N_11543);
nor U13310 (N_13310,N_11368,N_10710);
nand U13311 (N_13311,N_10946,N_11763);
nor U13312 (N_13312,N_10866,N_11964);
and U13313 (N_13313,N_11447,N_11109);
nor U13314 (N_13314,N_11291,N_10581);
nand U13315 (N_13315,N_10612,N_11659);
nor U13316 (N_13316,N_11353,N_10734);
and U13317 (N_13317,N_11328,N_11274);
nand U13318 (N_13318,N_11004,N_10762);
nand U13319 (N_13319,N_11790,N_11793);
xor U13320 (N_13320,N_11474,N_11601);
or U13321 (N_13321,N_11348,N_10562);
nand U13322 (N_13322,N_11932,N_10866);
nand U13323 (N_13323,N_10840,N_11509);
or U13324 (N_13324,N_11183,N_11050);
or U13325 (N_13325,N_10906,N_11566);
xnor U13326 (N_13326,N_11327,N_11655);
or U13327 (N_13327,N_11329,N_11942);
or U13328 (N_13328,N_11494,N_11768);
or U13329 (N_13329,N_11381,N_11175);
and U13330 (N_13330,N_10645,N_11653);
nor U13331 (N_13331,N_10925,N_10706);
nor U13332 (N_13332,N_11642,N_11504);
nor U13333 (N_13333,N_11821,N_11839);
or U13334 (N_13334,N_11856,N_10866);
and U13335 (N_13335,N_11132,N_10570);
xor U13336 (N_13336,N_10992,N_10790);
and U13337 (N_13337,N_11990,N_11248);
xnor U13338 (N_13338,N_10586,N_10821);
nor U13339 (N_13339,N_11793,N_11616);
or U13340 (N_13340,N_11929,N_10590);
nor U13341 (N_13341,N_11749,N_10976);
and U13342 (N_13342,N_11657,N_10807);
and U13343 (N_13343,N_10541,N_11718);
and U13344 (N_13344,N_11279,N_10966);
nand U13345 (N_13345,N_10595,N_11666);
and U13346 (N_13346,N_11804,N_10874);
nand U13347 (N_13347,N_11694,N_11696);
and U13348 (N_13348,N_11554,N_11058);
nand U13349 (N_13349,N_10715,N_11589);
and U13350 (N_13350,N_11136,N_11664);
or U13351 (N_13351,N_11280,N_11825);
or U13352 (N_13352,N_11917,N_11667);
or U13353 (N_13353,N_11027,N_11126);
and U13354 (N_13354,N_10836,N_11910);
nand U13355 (N_13355,N_11605,N_11735);
or U13356 (N_13356,N_11552,N_10994);
nor U13357 (N_13357,N_11087,N_11208);
nor U13358 (N_13358,N_11850,N_10878);
or U13359 (N_13359,N_10881,N_10756);
or U13360 (N_13360,N_10560,N_11604);
and U13361 (N_13361,N_11722,N_11274);
nand U13362 (N_13362,N_10772,N_11422);
and U13363 (N_13363,N_11778,N_10658);
and U13364 (N_13364,N_11543,N_11813);
or U13365 (N_13365,N_11885,N_11261);
nand U13366 (N_13366,N_11662,N_11305);
nand U13367 (N_13367,N_11790,N_10937);
nor U13368 (N_13368,N_11735,N_11079);
xnor U13369 (N_13369,N_10731,N_10803);
and U13370 (N_13370,N_11660,N_11059);
nand U13371 (N_13371,N_11494,N_11662);
and U13372 (N_13372,N_11647,N_11491);
xnor U13373 (N_13373,N_11287,N_10998);
and U13374 (N_13374,N_11118,N_11772);
nand U13375 (N_13375,N_11478,N_10728);
and U13376 (N_13376,N_10523,N_11082);
and U13377 (N_13377,N_10828,N_10648);
nor U13378 (N_13378,N_11125,N_11592);
or U13379 (N_13379,N_11516,N_11153);
or U13380 (N_13380,N_11832,N_11424);
and U13381 (N_13381,N_11364,N_10618);
nor U13382 (N_13382,N_10685,N_11943);
nor U13383 (N_13383,N_11861,N_11663);
nand U13384 (N_13384,N_11781,N_11025);
nor U13385 (N_13385,N_10564,N_10928);
nand U13386 (N_13386,N_10957,N_11428);
nand U13387 (N_13387,N_11938,N_11800);
and U13388 (N_13388,N_11021,N_11763);
nor U13389 (N_13389,N_11372,N_11187);
nor U13390 (N_13390,N_11732,N_11280);
nand U13391 (N_13391,N_11420,N_11429);
xor U13392 (N_13392,N_10950,N_11500);
and U13393 (N_13393,N_11833,N_11366);
and U13394 (N_13394,N_11520,N_11600);
nand U13395 (N_13395,N_11006,N_11830);
and U13396 (N_13396,N_11324,N_11497);
nor U13397 (N_13397,N_11308,N_10740);
and U13398 (N_13398,N_11832,N_10977);
nand U13399 (N_13399,N_10581,N_10788);
or U13400 (N_13400,N_10730,N_11664);
nand U13401 (N_13401,N_10514,N_11022);
nor U13402 (N_13402,N_11668,N_10572);
nor U13403 (N_13403,N_11348,N_11468);
and U13404 (N_13404,N_11025,N_11733);
or U13405 (N_13405,N_11405,N_11211);
nor U13406 (N_13406,N_10759,N_10986);
nor U13407 (N_13407,N_10728,N_11095);
nor U13408 (N_13408,N_10826,N_11284);
or U13409 (N_13409,N_11695,N_10712);
and U13410 (N_13410,N_11268,N_10608);
or U13411 (N_13411,N_10982,N_11064);
nor U13412 (N_13412,N_10538,N_11463);
nand U13413 (N_13413,N_11145,N_11186);
nor U13414 (N_13414,N_11728,N_11878);
nand U13415 (N_13415,N_11825,N_10900);
nand U13416 (N_13416,N_11199,N_11645);
nand U13417 (N_13417,N_11970,N_11370);
or U13418 (N_13418,N_10633,N_11886);
nand U13419 (N_13419,N_11228,N_11370);
xnor U13420 (N_13420,N_11538,N_10564);
nor U13421 (N_13421,N_10951,N_11325);
nor U13422 (N_13422,N_11448,N_11333);
nor U13423 (N_13423,N_11497,N_11639);
xnor U13424 (N_13424,N_11014,N_10588);
or U13425 (N_13425,N_11443,N_11073);
nand U13426 (N_13426,N_10895,N_10511);
and U13427 (N_13427,N_11025,N_11408);
or U13428 (N_13428,N_11768,N_11742);
and U13429 (N_13429,N_10643,N_10811);
nor U13430 (N_13430,N_11384,N_10686);
and U13431 (N_13431,N_11388,N_10828);
or U13432 (N_13432,N_10661,N_10951);
and U13433 (N_13433,N_11438,N_11140);
and U13434 (N_13434,N_11974,N_11452);
or U13435 (N_13435,N_11211,N_11521);
nand U13436 (N_13436,N_11041,N_11402);
nor U13437 (N_13437,N_11105,N_11034);
and U13438 (N_13438,N_11210,N_11273);
nand U13439 (N_13439,N_11651,N_10691);
nor U13440 (N_13440,N_11286,N_10500);
nand U13441 (N_13441,N_10536,N_11907);
and U13442 (N_13442,N_11509,N_11490);
nor U13443 (N_13443,N_10683,N_10812);
nand U13444 (N_13444,N_11075,N_10714);
and U13445 (N_13445,N_11332,N_11666);
nand U13446 (N_13446,N_11882,N_11564);
and U13447 (N_13447,N_11006,N_10632);
and U13448 (N_13448,N_11694,N_10976);
or U13449 (N_13449,N_11417,N_11826);
nor U13450 (N_13450,N_11576,N_11738);
and U13451 (N_13451,N_11614,N_11775);
nand U13452 (N_13452,N_11667,N_11332);
xnor U13453 (N_13453,N_10879,N_11643);
and U13454 (N_13454,N_11505,N_10676);
and U13455 (N_13455,N_11325,N_11036);
nand U13456 (N_13456,N_11022,N_11934);
nand U13457 (N_13457,N_10813,N_11388);
nand U13458 (N_13458,N_10598,N_11167);
nand U13459 (N_13459,N_11584,N_11211);
nand U13460 (N_13460,N_11791,N_11164);
nor U13461 (N_13461,N_11683,N_11059);
xnor U13462 (N_13462,N_10700,N_11579);
nor U13463 (N_13463,N_11441,N_11828);
or U13464 (N_13464,N_10628,N_11034);
nand U13465 (N_13465,N_10904,N_10645);
and U13466 (N_13466,N_11610,N_11103);
and U13467 (N_13467,N_11947,N_10703);
nand U13468 (N_13468,N_11553,N_10613);
or U13469 (N_13469,N_10776,N_11832);
and U13470 (N_13470,N_11075,N_11821);
and U13471 (N_13471,N_11436,N_10505);
nor U13472 (N_13472,N_10987,N_11023);
nor U13473 (N_13473,N_10805,N_11678);
nand U13474 (N_13474,N_11723,N_11013);
and U13475 (N_13475,N_11533,N_11149);
nand U13476 (N_13476,N_10553,N_10784);
and U13477 (N_13477,N_11895,N_11634);
and U13478 (N_13478,N_11253,N_11833);
and U13479 (N_13479,N_11732,N_11198);
nand U13480 (N_13480,N_11710,N_10571);
and U13481 (N_13481,N_11328,N_11723);
nor U13482 (N_13482,N_11539,N_10538);
nand U13483 (N_13483,N_11018,N_10882);
or U13484 (N_13484,N_11711,N_11024);
nand U13485 (N_13485,N_11635,N_11424);
or U13486 (N_13486,N_11965,N_11404);
xnor U13487 (N_13487,N_10966,N_10583);
and U13488 (N_13488,N_10876,N_11251);
nand U13489 (N_13489,N_11990,N_11679);
nand U13490 (N_13490,N_11302,N_10812);
nor U13491 (N_13491,N_11158,N_11690);
nand U13492 (N_13492,N_11897,N_11736);
nand U13493 (N_13493,N_11529,N_11283);
and U13494 (N_13494,N_10735,N_10511);
nand U13495 (N_13495,N_10799,N_10951);
and U13496 (N_13496,N_11694,N_10739);
and U13497 (N_13497,N_11181,N_10542);
nand U13498 (N_13498,N_11601,N_11308);
nor U13499 (N_13499,N_11632,N_10600);
xnor U13500 (N_13500,N_13398,N_12396);
nor U13501 (N_13501,N_13091,N_12285);
xor U13502 (N_13502,N_12872,N_12564);
or U13503 (N_13503,N_13057,N_12777);
or U13504 (N_13504,N_12211,N_12014);
nand U13505 (N_13505,N_12834,N_13331);
nand U13506 (N_13506,N_12560,N_13148);
or U13507 (N_13507,N_12798,N_12429);
or U13508 (N_13508,N_12679,N_13442);
nor U13509 (N_13509,N_13154,N_12613);
and U13510 (N_13510,N_13487,N_12929);
and U13511 (N_13511,N_12862,N_12704);
nand U13512 (N_13512,N_12382,N_12258);
nand U13513 (N_13513,N_12216,N_12267);
xor U13514 (N_13514,N_12774,N_13160);
nand U13515 (N_13515,N_12203,N_12128);
nand U13516 (N_13516,N_13413,N_12562);
nand U13517 (N_13517,N_12176,N_12260);
or U13518 (N_13518,N_12551,N_13299);
or U13519 (N_13519,N_12197,N_13462);
and U13520 (N_13520,N_12545,N_12845);
and U13521 (N_13521,N_12257,N_12603);
xor U13522 (N_13522,N_13086,N_13395);
nor U13523 (N_13523,N_12893,N_12379);
and U13524 (N_13524,N_12409,N_12702);
and U13525 (N_13525,N_12940,N_13447);
nand U13526 (N_13526,N_12754,N_12312);
nand U13527 (N_13527,N_12087,N_12620);
and U13528 (N_13528,N_13129,N_12601);
and U13529 (N_13529,N_13417,N_12424);
and U13530 (N_13530,N_12393,N_12277);
and U13531 (N_13531,N_13052,N_12824);
or U13532 (N_13532,N_12935,N_12838);
or U13533 (N_13533,N_13096,N_12237);
or U13534 (N_13534,N_12671,N_12638);
nand U13535 (N_13535,N_13290,N_12650);
nand U13536 (N_13536,N_12062,N_13268);
or U13537 (N_13537,N_12363,N_12591);
nand U13538 (N_13538,N_12991,N_13240);
xnor U13539 (N_13539,N_13062,N_12817);
nand U13540 (N_13540,N_13326,N_12522);
or U13541 (N_13541,N_13341,N_12222);
nand U13542 (N_13542,N_12959,N_12595);
nand U13543 (N_13543,N_13283,N_12544);
and U13544 (N_13544,N_12651,N_12200);
and U13545 (N_13545,N_13370,N_13421);
nand U13546 (N_13546,N_13213,N_12346);
xnor U13547 (N_13547,N_12910,N_12172);
nand U13548 (N_13548,N_12981,N_12292);
and U13549 (N_13549,N_12626,N_12144);
or U13550 (N_13550,N_12367,N_12863);
and U13551 (N_13551,N_12828,N_12303);
and U13552 (N_13552,N_13015,N_13353);
or U13553 (N_13553,N_12673,N_13409);
nand U13554 (N_13554,N_12475,N_12201);
or U13555 (N_13555,N_12892,N_12808);
xor U13556 (N_13556,N_13220,N_13403);
nor U13557 (N_13557,N_13125,N_12787);
nor U13558 (N_13558,N_13031,N_12415);
nand U13559 (N_13559,N_12231,N_12460);
or U13560 (N_13560,N_12670,N_12607);
or U13561 (N_13561,N_12107,N_13435);
and U13562 (N_13562,N_12625,N_13378);
xnor U13563 (N_13563,N_12871,N_13272);
and U13564 (N_13564,N_12778,N_12189);
xnor U13565 (N_13565,N_12581,N_13262);
or U13566 (N_13566,N_12122,N_12851);
or U13567 (N_13567,N_13004,N_13387);
nand U13568 (N_13568,N_13209,N_12814);
and U13569 (N_13569,N_13484,N_12282);
nor U13570 (N_13570,N_12448,N_12063);
nor U13571 (N_13571,N_12680,N_12842);
nor U13572 (N_13572,N_12686,N_13222);
and U13573 (N_13573,N_13118,N_12476);
nand U13574 (N_13574,N_12232,N_12726);
or U13575 (N_13575,N_12706,N_12012);
or U13576 (N_13576,N_12614,N_12406);
or U13577 (N_13577,N_12470,N_12677);
and U13578 (N_13578,N_12191,N_12418);
nand U13579 (N_13579,N_12199,N_12349);
and U13580 (N_13580,N_12903,N_12352);
nor U13581 (N_13581,N_13126,N_12002);
or U13582 (N_13582,N_12813,N_12752);
nor U13583 (N_13583,N_13279,N_12473);
nor U13584 (N_13584,N_13274,N_13266);
xor U13585 (N_13585,N_12345,N_13494);
xnor U13586 (N_13586,N_12032,N_12779);
nor U13587 (N_13587,N_13269,N_12598);
nor U13588 (N_13588,N_12036,N_13214);
and U13589 (N_13589,N_12207,N_12129);
nand U13590 (N_13590,N_12244,N_12105);
and U13591 (N_13591,N_12648,N_13249);
xnor U13592 (N_13592,N_13495,N_12286);
or U13593 (N_13593,N_12064,N_12442);
nor U13594 (N_13594,N_13349,N_12426);
or U13595 (N_13595,N_12117,N_12042);
or U13596 (N_13596,N_13168,N_12605);
nand U13597 (N_13597,N_12279,N_12511);
nor U13598 (N_13598,N_12536,N_13040);
and U13599 (N_13599,N_12717,N_13253);
or U13600 (N_13600,N_12274,N_12362);
nand U13601 (N_13601,N_12873,N_12775);
and U13602 (N_13602,N_12925,N_12293);
xor U13603 (N_13603,N_13431,N_12986);
nand U13604 (N_13604,N_13360,N_12301);
xor U13605 (N_13605,N_12911,N_13210);
xnor U13606 (N_13606,N_13449,N_13248);
nand U13607 (N_13607,N_12147,N_12302);
nand U13608 (N_13608,N_12633,N_13100);
and U13609 (N_13609,N_12608,N_12789);
or U13610 (N_13610,N_13282,N_12384);
or U13611 (N_13611,N_13109,N_13061);
xnor U13612 (N_13612,N_13416,N_12526);
nor U13613 (N_13613,N_12112,N_12322);
and U13614 (N_13614,N_12377,N_12185);
and U13615 (N_13615,N_12462,N_12395);
and U13616 (N_13616,N_12157,N_12832);
nor U13617 (N_13617,N_13055,N_13013);
or U13618 (N_13618,N_12988,N_12996);
nand U13619 (N_13619,N_12785,N_13362);
nand U13620 (N_13620,N_12289,N_12836);
xor U13621 (N_13621,N_12075,N_12241);
or U13622 (N_13622,N_12948,N_12950);
and U13623 (N_13623,N_13205,N_12657);
nor U13624 (N_13624,N_12103,N_12043);
or U13625 (N_13625,N_12655,N_12969);
or U13626 (N_13626,N_12849,N_12080);
and U13627 (N_13627,N_13485,N_12400);
and U13628 (N_13628,N_13489,N_12439);
nand U13629 (N_13629,N_13028,N_13263);
or U13630 (N_13630,N_12329,N_12891);
nand U13631 (N_13631,N_12599,N_13309);
or U13632 (N_13632,N_13173,N_13196);
or U13633 (N_13633,N_13251,N_12085);
or U13634 (N_13634,N_13415,N_12416);
or U13635 (N_13635,N_13161,N_12943);
and U13636 (N_13636,N_13250,N_13458);
and U13637 (N_13637,N_12719,N_12255);
nand U13638 (N_13638,N_13023,N_12627);
or U13639 (N_13639,N_13321,N_12003);
nor U13640 (N_13640,N_12713,N_12835);
nand U13641 (N_13641,N_12243,N_12529);
and U13642 (N_13642,N_13386,N_12983);
and U13643 (N_13643,N_12389,N_13008);
xnor U13644 (N_13644,N_12049,N_12746);
and U13645 (N_13645,N_12877,N_12446);
nor U13646 (N_13646,N_13034,N_12576);
and U13647 (N_13647,N_12639,N_12226);
or U13648 (N_13648,N_13163,N_12310);
xnor U13649 (N_13649,N_12502,N_12965);
xor U13650 (N_13650,N_12116,N_13418);
or U13651 (N_13651,N_13318,N_13158);
nor U13652 (N_13652,N_12963,N_12498);
nor U13653 (N_13653,N_13069,N_12005);
or U13654 (N_13654,N_12435,N_12334);
nand U13655 (N_13655,N_12166,N_13334);
nand U13656 (N_13656,N_12693,N_13448);
nor U13657 (N_13657,N_12033,N_12763);
nand U13658 (N_13658,N_12577,N_13133);
or U13659 (N_13659,N_12223,N_13373);
or U13660 (N_13660,N_12934,N_12356);
nor U13661 (N_13661,N_12177,N_12833);
nor U13662 (N_13662,N_12127,N_12390);
nand U13663 (N_13663,N_13192,N_12931);
and U13664 (N_13664,N_13037,N_13184);
nor U13665 (N_13665,N_13369,N_12812);
nand U13666 (N_13666,N_13146,N_12995);
and U13667 (N_13667,N_12060,N_13312);
xnor U13668 (N_13668,N_13194,N_13423);
nor U13669 (N_13669,N_12450,N_12245);
nor U13670 (N_13670,N_12654,N_12734);
or U13671 (N_13671,N_12913,N_12811);
and U13672 (N_13672,N_12205,N_13389);
or U13673 (N_13673,N_12699,N_13490);
and U13674 (N_13674,N_13344,N_12090);
nor U13675 (N_13675,N_13419,N_12731);
or U13676 (N_13676,N_12264,N_12610);
xor U13677 (N_13677,N_12490,N_12477);
nor U13678 (N_13678,N_12850,N_12521);
or U13679 (N_13679,N_12807,N_12797);
nand U13680 (N_13680,N_13257,N_12268);
nand U13681 (N_13681,N_12816,N_12664);
nor U13682 (N_13682,N_13228,N_13032);
nor U13683 (N_13683,N_13271,N_12479);
xor U13684 (N_13684,N_12410,N_12124);
nand U13685 (N_13685,N_13256,N_12436);
nand U13686 (N_13686,N_12408,N_12271);
nand U13687 (N_13687,N_13195,N_12380);
and U13688 (N_13688,N_12535,N_13367);
and U13689 (N_13689,N_12474,N_12993);
and U13690 (N_13690,N_12632,N_13302);
or U13691 (N_13691,N_13343,N_12839);
nor U13692 (N_13692,N_13451,N_12987);
or U13693 (N_13693,N_12137,N_12372);
and U13694 (N_13694,N_13217,N_12841);
nor U13695 (N_13695,N_12252,N_12451);
nand U13696 (N_13696,N_12433,N_12361);
and U13697 (N_13697,N_12924,N_12636);
xor U13698 (N_13698,N_12947,N_13258);
or U13699 (N_13699,N_12070,N_12484);
nand U13700 (N_13700,N_12558,N_13342);
and U13701 (N_13701,N_12360,N_12034);
nor U13702 (N_13702,N_12898,N_13443);
nor U13703 (N_13703,N_12242,N_12698);
and U13704 (N_13704,N_12944,N_13330);
nand U13705 (N_13705,N_12167,N_13246);
nor U13706 (N_13706,N_12159,N_12419);
or U13707 (N_13707,N_12154,N_13460);
nand U13708 (N_13708,N_12720,N_12325);
and U13709 (N_13709,N_13374,N_13012);
nand U13710 (N_13710,N_12238,N_13167);
and U13711 (N_13711,N_12121,N_13208);
nor U13712 (N_13712,N_13394,N_13223);
or U13713 (N_13713,N_12729,N_13313);
nor U13714 (N_13714,N_13426,N_13070);
nor U13715 (N_13715,N_12765,N_13292);
nor U13716 (N_13716,N_12273,N_12283);
nor U13717 (N_13717,N_13151,N_13306);
nand U13718 (N_13718,N_13245,N_12645);
or U13719 (N_13719,N_12974,N_12852);
or U13720 (N_13720,N_12151,N_12694);
xnor U13721 (N_13721,N_13232,N_12915);
and U13722 (N_13722,N_13317,N_13106);
nand U13723 (N_13723,N_12123,N_12051);
nor U13724 (N_13724,N_12964,N_12229);
nand U13725 (N_13725,N_12989,N_12617);
nor U13726 (N_13726,N_12888,N_13043);
and U13727 (N_13727,N_13089,N_13479);
nand U13728 (N_13728,N_13492,N_12225);
nand U13729 (N_13729,N_13138,N_12885);
nor U13730 (N_13730,N_12432,N_12027);
nand U13731 (N_13731,N_13017,N_13041);
or U13732 (N_13732,N_13322,N_13346);
nor U13733 (N_13733,N_13436,N_12712);
nand U13734 (N_13734,N_13095,N_13270);
nor U13735 (N_13735,N_12642,N_12593);
nor U13736 (N_13736,N_12708,N_12161);
and U13737 (N_13737,N_12879,N_12262);
xnor U13738 (N_13738,N_13388,N_13325);
or U13739 (N_13739,N_12725,N_12695);
nand U13740 (N_13740,N_12459,N_13345);
or U13741 (N_13741,N_12132,N_13265);
xor U13742 (N_13742,N_13324,N_12021);
or U13743 (N_13743,N_12554,N_12188);
nor U13744 (N_13744,N_13035,N_13390);
and U13745 (N_13745,N_13113,N_12641);
and U13746 (N_13746,N_12570,N_12826);
and U13747 (N_13747,N_13193,N_12737);
nand U13748 (N_13748,N_12643,N_12468);
nor U13749 (N_13749,N_12582,N_12357);
nand U13750 (N_13750,N_12198,N_13088);
nand U13751 (N_13751,N_12278,N_12170);
and U13752 (N_13752,N_12023,N_12004);
and U13753 (N_13753,N_12383,N_13082);
or U13754 (N_13754,N_13047,N_13131);
or U13755 (N_13755,N_13338,N_12156);
or U13756 (N_13756,N_12139,N_12256);
nand U13757 (N_13757,N_12882,N_13468);
and U13758 (N_13758,N_12365,N_12342);
or U13759 (N_13759,N_12876,N_12853);
xor U13760 (N_13760,N_13304,N_12316);
and U13761 (N_13761,N_12532,N_12456);
and U13762 (N_13762,N_12227,N_12573);
xor U13763 (N_13763,N_12392,N_12973);
and U13764 (N_13764,N_12295,N_12196);
xor U13765 (N_13765,N_13073,N_13289);
nor U13766 (N_13766,N_12982,N_12423);
or U13767 (N_13767,N_13284,N_13219);
nor U13768 (N_13768,N_12210,N_13459);
or U13769 (N_13769,N_13122,N_12584);
xnor U13770 (N_13770,N_12829,N_12482);
and U13771 (N_13771,N_12495,N_12319);
or U13772 (N_13772,N_12250,N_12594);
nor U13773 (N_13773,N_12178,N_13347);
nand U13774 (N_13774,N_12815,N_12097);
nor U13775 (N_13775,N_12369,N_12119);
or U13776 (N_13776,N_12135,N_12743);
and U13777 (N_13777,N_12452,N_12331);
and U13778 (N_13778,N_12492,N_12848);
nor U13779 (N_13779,N_12855,N_13049);
or U13780 (N_13780,N_12733,N_12703);
nand U13781 (N_13781,N_12265,N_12588);
nor U13782 (N_13782,N_13293,N_13036);
and U13783 (N_13783,N_12984,N_13110);
or U13784 (N_13784,N_13066,N_12761);
nand U13785 (N_13785,N_12762,N_13018);
nor U13786 (N_13786,N_12045,N_13156);
nand U13787 (N_13787,N_13359,N_12985);
or U13788 (N_13788,N_12275,N_12722);
nor U13789 (N_13789,N_13024,N_12221);
and U13790 (N_13790,N_12514,N_12634);
nand U13791 (N_13791,N_12220,N_12094);
nor U13792 (N_13792,N_12168,N_13111);
nor U13793 (N_13793,N_12736,N_13166);
xnor U13794 (N_13794,N_12402,N_13428);
nand U13795 (N_13795,N_12281,N_13425);
xor U13796 (N_13796,N_12270,N_13124);
nor U13797 (N_13797,N_12247,N_12209);
and U13798 (N_13798,N_12953,N_12854);
and U13799 (N_13799,N_12592,N_12269);
and U13800 (N_13800,N_12760,N_13296);
nor U13801 (N_13801,N_13307,N_12263);
or U13802 (N_13802,N_13169,N_12276);
or U13803 (N_13803,N_13164,N_12101);
or U13804 (N_13804,N_12037,N_12202);
and U13805 (N_13805,N_12580,N_13261);
and U13806 (N_13806,N_13295,N_12516);
and U13807 (N_13807,N_13237,N_12010);
and U13808 (N_13808,N_12745,N_12715);
nand U13809 (N_13809,N_12518,N_12542);
nand U13810 (N_13810,N_13420,N_12024);
xor U13811 (N_13811,N_13243,N_12099);
nor U13812 (N_13812,N_12174,N_12933);
and U13813 (N_13813,N_12669,N_13379);
or U13814 (N_13814,N_12134,N_12388);
or U13815 (N_13815,N_12351,N_13084);
and U13816 (N_13816,N_12895,N_12149);
and U13817 (N_13817,N_12297,N_13352);
nand U13818 (N_13818,N_13456,N_12425);
and U13819 (N_13819,N_12148,N_13044);
nand U13820 (N_13820,N_12249,N_13215);
nor U13821 (N_13821,N_12773,N_12102);
xnor U13822 (N_13822,N_12011,N_12016);
nor U13823 (N_13823,N_13063,N_12224);
or U13824 (N_13824,N_13189,N_13328);
or U13825 (N_13825,N_13337,N_12818);
xor U13826 (N_13826,N_13132,N_12524);
or U13827 (N_13827,N_12215,N_12530);
nor U13828 (N_13828,N_13402,N_13333);
and U13829 (N_13829,N_12788,N_12441);
nor U13830 (N_13830,N_12054,N_12674);
xnor U13831 (N_13831,N_12411,N_13311);
and U13832 (N_13832,N_12029,N_12538);
or U13833 (N_13833,N_13238,N_13368);
nand U13834 (N_13834,N_12055,N_12866);
nand U13835 (N_13835,N_13392,N_12730);
or U13836 (N_13836,N_12481,N_12748);
and U13837 (N_13837,N_12039,N_12398);
or U13838 (N_13838,N_12234,N_13310);
nand U13839 (N_13839,N_12096,N_13039);
nand U13840 (N_13840,N_12688,N_12098);
xnor U13841 (N_13841,N_12251,N_13178);
nor U13842 (N_13842,N_12772,N_12946);
or U13843 (N_13843,N_12799,N_13074);
nor U13844 (N_13844,N_12875,N_12653);
nand U13845 (N_13845,N_12485,N_12407);
nand U13846 (N_13846,N_12540,N_12480);
nor U13847 (N_13847,N_12978,N_12757);
xor U13848 (N_13848,N_12074,N_12696);
nor U13849 (N_13849,N_12022,N_13080);
or U13850 (N_13850,N_12507,N_12975);
and U13851 (N_13851,N_12195,N_12926);
or U13852 (N_13852,N_12528,N_12368);
xnor U13853 (N_13853,N_13050,N_12971);
and U13854 (N_13854,N_12496,N_13117);
and U13855 (N_13855,N_13134,N_12806);
or U13856 (N_13856,N_12072,N_13336);
and U13857 (N_13857,N_13446,N_13139);
nand U13858 (N_13858,N_13236,N_12077);
or U13859 (N_13859,N_12404,N_12317);
or U13860 (N_13860,N_12307,N_12999);
nor U13861 (N_13861,N_12864,N_12923);
nor U13862 (N_13862,N_12635,N_12510);
nor U13863 (N_13863,N_12488,N_13021);
nand U13864 (N_13864,N_13026,N_12458);
or U13865 (N_13865,N_12019,N_12445);
xor U13866 (N_13866,N_13294,N_12727);
and U13867 (N_13867,N_12505,N_12897);
and U13868 (N_13868,N_12192,N_13308);
and U13869 (N_13869,N_12878,N_12449);
or U13870 (N_13870,N_13059,N_12909);
nand U13871 (N_13871,N_12533,N_12417);
and U13872 (N_13872,N_12537,N_13065);
nand U13873 (N_13873,N_12881,N_13281);
xor U13874 (N_13874,N_12930,N_12823);
nand U13875 (N_13875,N_12942,N_13339);
or U13876 (N_13876,N_13083,N_12683);
xnor U13877 (N_13877,N_12115,N_13048);
xnor U13878 (N_13878,N_13497,N_13499);
or U13879 (N_13879,N_12682,N_13252);
nor U13880 (N_13880,N_12304,N_12714);
nor U13881 (N_13881,N_12574,N_12187);
nand U13882 (N_13882,N_12637,N_13198);
nor U13883 (N_13883,N_12499,N_13174);
nor U13884 (N_13884,N_12792,N_12171);
and U13885 (N_13885,N_12313,N_12628);
and U13886 (N_13886,N_12314,N_12622);
and U13887 (N_13887,N_12338,N_12755);
or U13888 (N_13888,N_13385,N_12579);
nor U13889 (N_13889,N_12454,N_13006);
or U13890 (N_13890,N_13212,N_12291);
nor U13891 (N_13891,N_12158,N_12596);
nor U13892 (N_13892,N_12018,N_13076);
nand U13893 (N_13893,N_12966,N_12932);
nand U13894 (N_13894,N_12515,N_12837);
nand U13895 (N_13895,N_13099,N_13022);
nand U13896 (N_13896,N_12890,N_12219);
and U13897 (N_13897,N_12728,N_13000);
or U13898 (N_13898,N_12284,N_12486);
and U13899 (N_13899,N_12880,N_12697);
nor U13900 (N_13900,N_13211,N_12658);
or U13901 (N_13901,N_13206,N_12769);
nor U13902 (N_13902,N_12443,N_13121);
nor U13903 (N_13903,N_13165,N_12753);
or U13904 (N_13904,N_13465,N_12901);
nor U13905 (N_13905,N_13014,N_12155);
xnor U13906 (N_13906,N_12527,N_12374);
and U13907 (N_13907,N_12391,N_12309);
and U13908 (N_13908,N_13473,N_12353);
nor U13909 (N_13909,N_13203,N_12186);
or U13910 (N_13910,N_13463,N_12548);
nand U13911 (N_13911,N_13051,N_12358);
and U13912 (N_13912,N_12457,N_12348);
and U13913 (N_13913,N_12615,N_12491);
nand U13914 (N_13914,N_13453,N_12142);
or U13915 (N_13915,N_12744,N_12444);
and U13916 (N_13916,N_13199,N_12681);
and U13917 (N_13917,N_13277,N_12434);
or U13918 (N_13918,N_13010,N_12689);
nor U13919 (N_13919,N_13285,N_12938);
nor U13920 (N_13920,N_13445,N_13332);
nor U13921 (N_13921,N_12290,N_13297);
xor U13922 (N_13922,N_12738,N_12870);
nor U13923 (N_13923,N_13365,N_12604);
nand U13924 (N_13924,N_12179,N_12071);
nand U13925 (N_13925,N_13414,N_13135);
or U13926 (N_13926,N_13241,N_12519);
and U13927 (N_13927,N_13225,N_13185);
nor U13928 (N_13928,N_12413,N_12906);
nor U13929 (N_13929,N_13244,N_12246);
or U13930 (N_13930,N_13016,N_13187);
nor U13931 (N_13931,N_12233,N_13234);
xor U13932 (N_13932,N_13033,N_12990);
and U13933 (N_13933,N_13108,N_12500);
nor U13934 (N_13934,N_13483,N_12568);
nand U13935 (N_13935,N_13119,N_12563);
and U13936 (N_13936,N_12919,N_12578);
nor U13937 (N_13937,N_12623,N_12387);
nand U13938 (N_13938,N_12958,N_13137);
nor U13939 (N_13939,N_12130,N_13183);
or U13940 (N_13940,N_12028,N_12184);
nand U13941 (N_13941,N_13221,N_13377);
and U13942 (N_13942,N_12937,N_12865);
nand U13943 (N_13943,N_12764,N_13072);
nor U13944 (N_13944,N_12489,N_12253);
nand U13945 (N_13945,N_12711,N_12742);
nand U13946 (N_13946,N_12861,N_12684);
nand U13947 (N_13947,N_12050,N_12204);
or U13948 (N_13948,N_13384,N_12165);
or U13949 (N_13949,N_12649,N_13375);
nor U13950 (N_13950,N_13071,N_13315);
and U13951 (N_13951,N_12206,N_12503);
xor U13952 (N_13952,N_12026,N_13439);
and U13953 (N_13953,N_12145,N_12666);
or U13954 (N_13954,N_12464,N_13218);
nand U13955 (N_13955,N_12756,N_12376);
or U13956 (N_13956,N_12618,N_12180);
and U13957 (N_13957,N_13280,N_12668);
nor U13958 (N_13958,N_12954,N_13247);
or U13959 (N_13959,N_13466,N_12455);
nand U13960 (N_13960,N_12830,N_12979);
nor U13961 (N_13961,N_12401,N_12998);
and U13962 (N_13962,N_12970,N_12336);
nand U13963 (N_13963,N_12905,N_13438);
and U13964 (N_13964,N_13475,N_13180);
nand U13965 (N_13965,N_13363,N_13254);
and U13966 (N_13966,N_13481,N_13090);
and U13967 (N_13967,N_12952,N_12869);
and U13968 (N_13968,N_12556,N_13042);
or U13969 (N_13969,N_12859,N_12751);
nand U13970 (N_13970,N_12371,N_12254);
and U13971 (N_13971,N_13396,N_12108);
or U13972 (N_13972,N_12431,N_12732);
and U13973 (N_13973,N_13058,N_13201);
or U13974 (N_13974,N_12506,N_12333);
nor U13975 (N_13975,N_12800,N_12553);
and U13976 (N_13976,N_13441,N_12136);
or U13977 (N_13977,N_12784,N_13354);
xnor U13978 (N_13978,N_12525,N_12575);
and U13979 (N_13979,N_13153,N_12889);
nand U13980 (N_13980,N_12083,N_12945);
and U13981 (N_13981,N_12093,N_12821);
and U13982 (N_13982,N_12927,N_12914);
and U13983 (N_13983,N_12046,N_13364);
nor U13984 (N_13984,N_12860,N_12631);
nand U13985 (N_13985,N_12710,N_12447);
nor U13986 (N_13986,N_13276,N_13207);
or U13987 (N_13987,N_12587,N_12550);
nor U13988 (N_13988,N_13202,N_12339);
or U13989 (N_13989,N_12126,N_12110);
or U13990 (N_13990,N_12118,N_13170);
nor U13991 (N_13991,N_12796,N_12053);
and U13992 (N_13992,N_13319,N_12175);
xnor U13993 (N_13993,N_12790,N_12543);
or U13994 (N_13994,N_13476,N_12163);
nor U13995 (N_13995,N_13176,N_13029);
and U13996 (N_13996,N_12463,N_13371);
xor U13997 (N_13997,N_12955,N_13382);
or U13998 (N_13998,N_12076,N_13397);
or U13999 (N_13999,N_12678,N_12230);
xor U14000 (N_14000,N_13162,N_13393);
or U14001 (N_14001,N_12164,N_12483);
nor U14002 (N_14002,N_12287,N_13060);
nand U14003 (N_14003,N_12771,N_12768);
or U14004 (N_14004,N_12918,N_12822);
nand U14005 (N_14005,N_12138,N_12058);
nand U14006 (N_14006,N_13019,N_13340);
and U14007 (N_14007,N_13452,N_12106);
nand U14008 (N_14008,N_13025,N_12335);
and U14009 (N_14009,N_12846,N_12068);
nand U14010 (N_14010,N_12009,N_13054);
and U14011 (N_14011,N_12856,N_12359);
nor U14012 (N_14012,N_12646,N_12700);
and U14013 (N_14013,N_13102,N_12364);
nor U14014 (N_14014,N_12373,N_12957);
or U14015 (N_14015,N_12612,N_12193);
nor U14016 (N_14016,N_12378,N_13300);
nand U14017 (N_14017,N_13114,N_12044);
nor U14018 (N_14018,N_12960,N_13235);
and U14019 (N_14019,N_13401,N_12968);
nor U14020 (N_14020,N_13191,N_13348);
and U14021 (N_14021,N_12504,N_13150);
nor U14022 (N_14022,N_12904,N_12723);
or U14023 (N_14023,N_12802,N_12173);
nor U14024 (N_14024,N_13155,N_13491);
and U14025 (N_14025,N_13188,N_13406);
nand U14026 (N_14026,N_13464,N_13087);
and U14027 (N_14027,N_12992,N_13093);
nor U14028 (N_14028,N_13200,N_12735);
nand U14029 (N_14029,N_12555,N_12624);
and U14030 (N_14030,N_12217,N_12041);
or U14031 (N_14031,N_12261,N_12513);
nand U14032 (N_14032,N_12111,N_12386);
and U14033 (N_14033,N_12782,N_13305);
and U14034 (N_14034,N_12472,N_12017);
or U14035 (N_14035,N_12056,N_12493);
or U14036 (N_14036,N_12619,N_12665);
nor U14037 (N_14037,N_13467,N_12541);
xnor U14038 (N_14038,N_12928,N_12977);
nand U14039 (N_14039,N_12299,N_12208);
nor U14040 (N_14040,N_12059,N_12810);
and U14041 (N_14041,N_13381,N_13242);
or U14042 (N_14042,N_12825,N_12994);
nand U14043 (N_14043,N_13190,N_13461);
nor U14044 (N_14044,N_13267,N_12652);
nand U14045 (N_14045,N_12921,N_13264);
nand U14046 (N_14046,N_13112,N_12323);
nor U14047 (N_14047,N_12586,N_12381);
or U14048 (N_14048,N_12660,N_12520);
xnor U14049 (N_14049,N_12494,N_13077);
nand U14050 (N_14050,N_12428,N_13030);
nand U14051 (N_14051,N_12770,N_12330);
and U14052 (N_14052,N_13329,N_12793);
nand U14053 (N_14053,N_13301,N_13287);
xnor U14054 (N_14054,N_12015,N_12061);
and U14055 (N_14055,N_12235,N_13278);
or U14056 (N_14056,N_12565,N_13255);
nand U14057 (N_14057,N_13434,N_12427);
or U14058 (N_14058,N_13260,N_13229);
nor U14059 (N_14059,N_12962,N_13437);
and U14060 (N_14060,N_12306,N_13009);
or U14061 (N_14061,N_13496,N_12236);
nor U14062 (N_14062,N_13275,N_12557);
and U14063 (N_14063,N_12886,N_13227);
nand U14064 (N_14064,N_12583,N_12585);
xor U14065 (N_14065,N_12355,N_13147);
xnor U14066 (N_14066,N_12162,N_12440);
nor U14067 (N_14067,N_12160,N_12766);
or U14068 (N_14068,N_12844,N_12939);
xnor U14069 (N_14069,N_13303,N_12294);
nor U14070 (N_14070,N_12095,N_13433);
nor U14071 (N_14071,N_13358,N_13157);
nor U14072 (N_14072,N_13107,N_12767);
xnor U14073 (N_14073,N_13273,N_12883);
and U14074 (N_14074,N_13186,N_12340);
and U14075 (N_14075,N_12212,N_12786);
and U14076 (N_14076,N_12916,N_12405);
xor U14077 (N_14077,N_13092,N_13141);
or U14078 (N_14078,N_12783,N_13046);
and U14079 (N_14079,N_12438,N_12153);
nor U14080 (N_14080,N_12676,N_12917);
nand U14081 (N_14081,N_12847,N_12397);
or U14082 (N_14082,N_13179,N_13079);
nor U14083 (N_14083,N_12315,N_12795);
nand U14084 (N_14084,N_12794,N_13335);
and U14085 (N_14085,N_13357,N_13470);
nor U14086 (N_14086,N_13471,N_13440);
nand U14087 (N_14087,N_12190,N_12350);
nor U14088 (N_14088,N_12858,N_12240);
nand U14089 (N_14089,N_12741,N_12600);
and U14090 (N_14090,N_12920,N_13411);
nor U14091 (N_14091,N_13410,N_13064);
nand U14092 (N_14092,N_12001,N_12549);
and U14093 (N_14093,N_13038,N_13078);
or U14094 (N_14094,N_13020,N_12394);
xnor U14095 (N_14095,N_13053,N_12716);
nor U14096 (N_14096,N_13430,N_13323);
nand U14097 (N_14097,N_12567,N_13314);
or U14098 (N_14098,N_12508,N_12182);
nor U14099 (N_14099,N_12248,N_12311);
nand U14100 (N_14100,N_12038,N_12308);
xor U14101 (N_14101,N_13444,N_13288);
or U14102 (N_14102,N_13298,N_12332);
nand U14103 (N_14103,N_12709,N_12531);
xor U14104 (N_14104,N_12228,N_13075);
or U14105 (N_14105,N_12092,N_12214);
and U14106 (N_14106,N_12354,N_12692);
nand U14107 (N_14107,N_12467,N_12820);
nand U14108 (N_14108,N_12907,N_12104);
and U14109 (N_14109,N_12894,N_12073);
or U14110 (N_14110,N_13120,N_12663);
xnor U14111 (N_14111,N_12366,N_12296);
nand U14112 (N_14112,N_12320,N_13136);
and U14113 (N_14113,N_12086,N_13005);
nor U14114 (N_14114,N_12422,N_12078);
and U14115 (N_14115,N_12280,N_12412);
or U14116 (N_14116,N_12512,N_12884);
xnor U14117 (N_14117,N_13472,N_13366);
nand U14118 (N_14118,N_12239,N_13376);
and U14119 (N_14119,N_12747,N_12066);
nand U14120 (N_14120,N_13159,N_13493);
and U14121 (N_14121,N_12375,N_12120);
nand U14122 (N_14122,N_13488,N_13182);
nand U14123 (N_14123,N_13400,N_12899);
and U14124 (N_14124,N_13454,N_13391);
and U14125 (N_14125,N_12081,N_12724);
or U14126 (N_14126,N_12659,N_12052);
nor U14127 (N_14127,N_12082,N_13380);
xnor U14128 (N_14128,N_12672,N_12749);
and U14129 (N_14129,N_12067,N_13101);
nor U14130 (N_14130,N_13144,N_12469);
and U14131 (N_14131,N_12125,N_12150);
and U14132 (N_14132,N_12133,N_12152);
nand U14133 (N_14133,N_12656,N_13327);
nand U14134 (N_14134,N_12566,N_12007);
xnor U14135 (N_14135,N_13003,N_12000);
and U14136 (N_14136,N_13177,N_13412);
nand U14137 (N_14137,N_13351,N_12571);
xnor U14138 (N_14138,N_13097,N_12194);
and U14139 (N_14139,N_12759,N_12647);
nor U14140 (N_14140,N_13286,N_13478);
or U14141 (N_14141,N_12896,N_13098);
or U14142 (N_14142,N_13143,N_12569);
and U14143 (N_14143,N_12874,N_13007);
or U14144 (N_14144,N_12084,N_12547);
nand U14145 (N_14145,N_12661,N_12140);
xnor U14146 (N_14146,N_12501,N_12047);
nand U14147 (N_14147,N_12146,N_12035);
and U14148 (N_14148,N_13056,N_12539);
and U14149 (N_14149,N_12403,N_12385);
and U14150 (N_14150,N_12561,N_13011);
nor U14151 (N_14151,N_13045,N_12809);
and U14152 (N_14152,N_12590,N_12272);
nand U14153 (N_14153,N_13424,N_13068);
and U14154 (N_14154,N_13152,N_13239);
nand U14155 (N_14155,N_12523,N_12288);
and U14156 (N_14156,N_12305,N_12065);
and U14157 (N_14157,N_13422,N_12008);
or U14158 (N_14158,N_12318,N_13067);
nand U14159 (N_14159,N_12675,N_12300);
nand U14160 (N_14160,N_12347,N_12776);
nand U14161 (N_14161,N_13356,N_12109);
or U14162 (N_14162,N_12509,N_12621);
nor U14163 (N_14163,N_12956,N_12819);
or U14164 (N_14164,N_12025,N_12804);
xnor U14165 (N_14165,N_12517,N_12143);
nand U14166 (N_14166,N_13480,N_13127);
nor U14167 (N_14167,N_12606,N_13320);
and U14168 (N_14168,N_13316,N_13130);
xor U14169 (N_14169,N_12478,N_13145);
nand U14170 (N_14170,N_12707,N_13427);
nand U14171 (N_14171,N_13094,N_12031);
nor U14172 (N_14172,N_12687,N_12420);
or U14173 (N_14173,N_12370,N_13457);
nand U14174 (N_14174,N_12629,N_12739);
and U14175 (N_14175,N_12900,N_12857);
or U14176 (N_14176,N_12465,N_13105);
nand U14177 (N_14177,N_13085,N_12972);
nor U14178 (N_14178,N_12980,N_12867);
xor U14179 (N_14179,N_12298,N_12213);
or U14180 (N_14180,N_12069,N_12902);
and U14181 (N_14181,N_13123,N_13405);
or U14182 (N_14182,N_12967,N_12337);
nor U14183 (N_14183,N_13350,N_12718);
xnor U14184 (N_14184,N_12266,N_12006);
nor U14185 (N_14185,N_12597,N_12430);
and U14186 (N_14186,N_12805,N_12951);
xor U14187 (N_14187,N_12326,N_13455);
or U14188 (N_14188,N_12327,N_12572);
or U14189 (N_14189,N_13172,N_12114);
nor U14190 (N_14190,N_12602,N_12644);
xor U14191 (N_14191,N_13128,N_12831);
nand U14192 (N_14192,N_13482,N_12487);
and U14193 (N_14193,N_12721,N_12559);
nor U14194 (N_14194,N_12113,N_12801);
nand U14195 (N_14195,N_12780,N_12259);
or U14196 (N_14196,N_12183,N_12091);
or U14197 (N_14197,N_13197,N_12497);
and U14198 (N_14198,N_13486,N_12534);
and U14199 (N_14199,N_13103,N_13259);
and U14200 (N_14200,N_12936,N_13477);
or U14201 (N_14201,N_12912,N_13116);
and U14202 (N_14202,N_13230,N_12827);
and U14203 (N_14203,N_12040,N_12908);
and U14204 (N_14204,N_12758,N_12701);
or U14205 (N_14205,N_12868,N_12088);
and U14206 (N_14206,N_12079,N_13226);
nand U14207 (N_14207,N_13027,N_13142);
and U14208 (N_14208,N_13429,N_13171);
nand U14209 (N_14209,N_13216,N_13474);
xnor U14210 (N_14210,N_13399,N_12690);
nor U14211 (N_14211,N_13498,N_12750);
xor U14212 (N_14212,N_12616,N_13372);
or U14213 (N_14213,N_12181,N_12781);
or U14214 (N_14214,N_12328,N_12843);
nand U14215 (N_14215,N_13001,N_12840);
and U14216 (N_14216,N_12630,N_12611);
nand U14217 (N_14217,N_12321,N_13081);
and U14218 (N_14218,N_13149,N_12399);
or U14219 (N_14219,N_13002,N_13291);
nor U14220 (N_14220,N_12100,N_12941);
nand U14221 (N_14221,N_13383,N_12013);
nor U14222 (N_14222,N_12437,N_12048);
nand U14223 (N_14223,N_13175,N_13355);
nand U14224 (N_14224,N_12453,N_13469);
nand U14225 (N_14225,N_12922,N_12997);
and U14226 (N_14226,N_12141,N_12705);
and U14227 (N_14227,N_13404,N_13204);
or U14228 (N_14228,N_12640,N_13115);
and U14229 (N_14229,N_12791,N_13450);
nand U14230 (N_14230,N_12218,N_12344);
and U14231 (N_14231,N_13407,N_12740);
nor U14232 (N_14232,N_12471,N_12961);
or U14233 (N_14233,N_12461,N_13140);
nor U14234 (N_14234,N_12466,N_12169);
nor U14235 (N_14235,N_12949,N_13432);
and U14236 (N_14236,N_12803,N_12020);
and U14237 (N_14237,N_12414,N_13231);
nor U14238 (N_14238,N_13233,N_13224);
or U14239 (N_14239,N_12089,N_12691);
nor U14240 (N_14240,N_12667,N_12030);
and U14241 (N_14241,N_13361,N_12131);
and U14242 (N_14242,N_13408,N_12976);
nor U14243 (N_14243,N_12685,N_12887);
nor U14244 (N_14244,N_13104,N_12609);
nor U14245 (N_14245,N_12057,N_12546);
and U14246 (N_14246,N_12343,N_12341);
nand U14247 (N_14247,N_12662,N_13181);
nor U14248 (N_14248,N_12589,N_12324);
and U14249 (N_14249,N_12421,N_12552);
nor U14250 (N_14250,N_12963,N_12177);
nand U14251 (N_14251,N_12957,N_12432);
nand U14252 (N_14252,N_12231,N_13065);
nor U14253 (N_14253,N_13150,N_12004);
and U14254 (N_14254,N_12332,N_13212);
and U14255 (N_14255,N_12574,N_12529);
nor U14256 (N_14256,N_12537,N_13241);
and U14257 (N_14257,N_12423,N_13255);
xor U14258 (N_14258,N_12433,N_12717);
or U14259 (N_14259,N_13093,N_12491);
xnor U14260 (N_14260,N_13081,N_12822);
and U14261 (N_14261,N_12294,N_12125);
nor U14262 (N_14262,N_12056,N_12776);
or U14263 (N_14263,N_12744,N_12510);
nand U14264 (N_14264,N_13411,N_13484);
nand U14265 (N_14265,N_12328,N_13325);
nor U14266 (N_14266,N_12552,N_12634);
and U14267 (N_14267,N_12529,N_13197);
or U14268 (N_14268,N_12451,N_12522);
and U14269 (N_14269,N_13499,N_12583);
or U14270 (N_14270,N_13483,N_12029);
nand U14271 (N_14271,N_12900,N_12311);
nor U14272 (N_14272,N_13045,N_12390);
or U14273 (N_14273,N_12940,N_13105);
xnor U14274 (N_14274,N_13420,N_12017);
or U14275 (N_14275,N_12024,N_12744);
nand U14276 (N_14276,N_13274,N_12247);
and U14277 (N_14277,N_12619,N_12653);
or U14278 (N_14278,N_12649,N_12069);
and U14279 (N_14279,N_12894,N_12456);
xor U14280 (N_14280,N_12551,N_12783);
or U14281 (N_14281,N_13257,N_12861);
nor U14282 (N_14282,N_12628,N_12508);
and U14283 (N_14283,N_12088,N_13128);
or U14284 (N_14284,N_12231,N_13353);
nor U14285 (N_14285,N_12890,N_12861);
nor U14286 (N_14286,N_12463,N_12619);
nor U14287 (N_14287,N_12947,N_13494);
or U14288 (N_14288,N_13101,N_12103);
nor U14289 (N_14289,N_12796,N_12428);
xor U14290 (N_14290,N_12966,N_12857);
nor U14291 (N_14291,N_13238,N_12718);
nand U14292 (N_14292,N_12134,N_12898);
nor U14293 (N_14293,N_12326,N_13305);
or U14294 (N_14294,N_12696,N_12911);
nor U14295 (N_14295,N_12300,N_12933);
or U14296 (N_14296,N_12321,N_13219);
and U14297 (N_14297,N_13351,N_12826);
nor U14298 (N_14298,N_12746,N_12441);
nand U14299 (N_14299,N_12552,N_12555);
and U14300 (N_14300,N_12496,N_12281);
nor U14301 (N_14301,N_12740,N_12382);
nand U14302 (N_14302,N_12414,N_13006);
xnor U14303 (N_14303,N_13180,N_12028);
nor U14304 (N_14304,N_12911,N_12791);
nor U14305 (N_14305,N_12710,N_12765);
xnor U14306 (N_14306,N_12100,N_12136);
xnor U14307 (N_14307,N_12645,N_12656);
nor U14308 (N_14308,N_13040,N_12738);
and U14309 (N_14309,N_13157,N_13349);
or U14310 (N_14310,N_12649,N_12080);
xor U14311 (N_14311,N_13325,N_13265);
and U14312 (N_14312,N_12182,N_12377);
xor U14313 (N_14313,N_12643,N_13489);
xnor U14314 (N_14314,N_13264,N_12449);
nor U14315 (N_14315,N_12185,N_13076);
xnor U14316 (N_14316,N_12164,N_12153);
and U14317 (N_14317,N_12653,N_12308);
nand U14318 (N_14318,N_13151,N_12342);
nand U14319 (N_14319,N_12697,N_12337);
nand U14320 (N_14320,N_12959,N_12539);
and U14321 (N_14321,N_12925,N_13466);
xnor U14322 (N_14322,N_13409,N_12100);
and U14323 (N_14323,N_12109,N_12105);
and U14324 (N_14324,N_12155,N_12780);
nor U14325 (N_14325,N_12739,N_12483);
xor U14326 (N_14326,N_13415,N_12467);
nand U14327 (N_14327,N_12251,N_12180);
nor U14328 (N_14328,N_13332,N_13002);
xor U14329 (N_14329,N_12698,N_13443);
or U14330 (N_14330,N_12727,N_12495);
nand U14331 (N_14331,N_13051,N_12463);
xnor U14332 (N_14332,N_12872,N_13472);
or U14333 (N_14333,N_12180,N_12093);
nor U14334 (N_14334,N_12441,N_12311);
nor U14335 (N_14335,N_12848,N_12927);
nand U14336 (N_14336,N_13040,N_13316);
nand U14337 (N_14337,N_12436,N_13037);
and U14338 (N_14338,N_12101,N_12785);
and U14339 (N_14339,N_12515,N_13310);
nand U14340 (N_14340,N_13049,N_12473);
nand U14341 (N_14341,N_12937,N_12267);
nand U14342 (N_14342,N_12396,N_12080);
nor U14343 (N_14343,N_13006,N_13041);
nor U14344 (N_14344,N_12923,N_12057);
and U14345 (N_14345,N_13049,N_12535);
and U14346 (N_14346,N_12261,N_12220);
nor U14347 (N_14347,N_12788,N_12320);
or U14348 (N_14348,N_12045,N_12950);
and U14349 (N_14349,N_12565,N_12136);
nand U14350 (N_14350,N_12767,N_13239);
and U14351 (N_14351,N_13384,N_13019);
or U14352 (N_14352,N_13497,N_12530);
and U14353 (N_14353,N_12174,N_12882);
xnor U14354 (N_14354,N_12153,N_12440);
nand U14355 (N_14355,N_12118,N_13460);
nand U14356 (N_14356,N_12567,N_13384);
nand U14357 (N_14357,N_12059,N_13294);
nand U14358 (N_14358,N_12766,N_12880);
or U14359 (N_14359,N_12106,N_12157);
nand U14360 (N_14360,N_13121,N_12387);
and U14361 (N_14361,N_13324,N_12301);
xnor U14362 (N_14362,N_12759,N_12567);
nand U14363 (N_14363,N_12192,N_12073);
nor U14364 (N_14364,N_12753,N_13285);
xnor U14365 (N_14365,N_12076,N_13041);
xor U14366 (N_14366,N_12132,N_12152);
xor U14367 (N_14367,N_12988,N_13075);
nand U14368 (N_14368,N_12547,N_13150);
or U14369 (N_14369,N_12913,N_12556);
nor U14370 (N_14370,N_12661,N_12301);
nand U14371 (N_14371,N_12402,N_12834);
or U14372 (N_14372,N_13248,N_13486);
and U14373 (N_14373,N_12763,N_12431);
or U14374 (N_14374,N_13287,N_12932);
or U14375 (N_14375,N_12154,N_13149);
and U14376 (N_14376,N_12559,N_12877);
or U14377 (N_14377,N_12231,N_12197);
or U14378 (N_14378,N_12651,N_12289);
or U14379 (N_14379,N_12168,N_13047);
or U14380 (N_14380,N_12525,N_12288);
nor U14381 (N_14381,N_13348,N_12088);
xnor U14382 (N_14382,N_13026,N_13233);
or U14383 (N_14383,N_12685,N_12436);
and U14384 (N_14384,N_12119,N_12648);
or U14385 (N_14385,N_12000,N_12077);
nor U14386 (N_14386,N_13065,N_12306);
nand U14387 (N_14387,N_12941,N_12691);
nor U14388 (N_14388,N_13226,N_12614);
nor U14389 (N_14389,N_12999,N_12130);
or U14390 (N_14390,N_13357,N_12722);
nand U14391 (N_14391,N_12378,N_13390);
nor U14392 (N_14392,N_12492,N_12300);
and U14393 (N_14393,N_12366,N_13223);
nand U14394 (N_14394,N_12320,N_13064);
nor U14395 (N_14395,N_12749,N_12170);
or U14396 (N_14396,N_13020,N_12913);
nor U14397 (N_14397,N_13246,N_13082);
nand U14398 (N_14398,N_12506,N_12223);
nand U14399 (N_14399,N_13412,N_12864);
nand U14400 (N_14400,N_13025,N_13217);
xor U14401 (N_14401,N_12492,N_12811);
and U14402 (N_14402,N_12973,N_12399);
or U14403 (N_14403,N_12252,N_12535);
or U14404 (N_14404,N_12043,N_12973);
nand U14405 (N_14405,N_12785,N_12018);
xor U14406 (N_14406,N_12993,N_13056);
and U14407 (N_14407,N_12378,N_13364);
or U14408 (N_14408,N_12496,N_12594);
or U14409 (N_14409,N_12646,N_13088);
and U14410 (N_14410,N_12077,N_13005);
nand U14411 (N_14411,N_13411,N_12217);
nand U14412 (N_14412,N_12673,N_12046);
xor U14413 (N_14413,N_13485,N_12992);
or U14414 (N_14414,N_12905,N_13240);
or U14415 (N_14415,N_12212,N_13371);
and U14416 (N_14416,N_12551,N_13362);
and U14417 (N_14417,N_12040,N_13134);
and U14418 (N_14418,N_12315,N_12834);
nor U14419 (N_14419,N_12015,N_12395);
nand U14420 (N_14420,N_13287,N_12260);
nor U14421 (N_14421,N_12398,N_12104);
or U14422 (N_14422,N_13237,N_12989);
and U14423 (N_14423,N_12618,N_12113);
or U14424 (N_14424,N_12460,N_12899);
xnor U14425 (N_14425,N_12750,N_12587);
or U14426 (N_14426,N_12027,N_12401);
and U14427 (N_14427,N_12979,N_12726);
nand U14428 (N_14428,N_12866,N_13376);
nor U14429 (N_14429,N_12768,N_13189);
nor U14430 (N_14430,N_12104,N_13119);
nand U14431 (N_14431,N_13212,N_12962);
and U14432 (N_14432,N_12267,N_12977);
or U14433 (N_14433,N_12011,N_13224);
nor U14434 (N_14434,N_13443,N_13390);
and U14435 (N_14435,N_12219,N_12453);
xnor U14436 (N_14436,N_12887,N_12241);
and U14437 (N_14437,N_12174,N_12098);
or U14438 (N_14438,N_12082,N_13340);
and U14439 (N_14439,N_13253,N_13371);
and U14440 (N_14440,N_12002,N_12956);
or U14441 (N_14441,N_12231,N_13104);
and U14442 (N_14442,N_12755,N_12402);
or U14443 (N_14443,N_12194,N_12190);
nor U14444 (N_14444,N_12125,N_12888);
nor U14445 (N_14445,N_12601,N_13031);
and U14446 (N_14446,N_13033,N_12367);
and U14447 (N_14447,N_12245,N_13190);
or U14448 (N_14448,N_12597,N_12839);
and U14449 (N_14449,N_12768,N_13143);
nand U14450 (N_14450,N_12210,N_12618);
xnor U14451 (N_14451,N_12467,N_12773);
or U14452 (N_14452,N_12452,N_13359);
nor U14453 (N_14453,N_12321,N_13042);
xor U14454 (N_14454,N_12711,N_13130);
xor U14455 (N_14455,N_13009,N_13137);
or U14456 (N_14456,N_12589,N_12035);
and U14457 (N_14457,N_13394,N_12650);
nor U14458 (N_14458,N_13237,N_12634);
or U14459 (N_14459,N_12268,N_12103);
and U14460 (N_14460,N_12649,N_13330);
xor U14461 (N_14461,N_13333,N_12552);
and U14462 (N_14462,N_13178,N_12897);
nand U14463 (N_14463,N_12212,N_12481);
or U14464 (N_14464,N_12411,N_12363);
or U14465 (N_14465,N_12875,N_12407);
or U14466 (N_14466,N_12487,N_12094);
nand U14467 (N_14467,N_12648,N_12376);
xor U14468 (N_14468,N_13048,N_12666);
and U14469 (N_14469,N_13469,N_12058);
xnor U14470 (N_14470,N_12056,N_13486);
or U14471 (N_14471,N_13169,N_12637);
and U14472 (N_14472,N_13405,N_12178);
and U14473 (N_14473,N_12563,N_12792);
xor U14474 (N_14474,N_13095,N_13253);
and U14475 (N_14475,N_12293,N_13400);
and U14476 (N_14476,N_12476,N_13087);
xnor U14477 (N_14477,N_13069,N_12878);
nor U14478 (N_14478,N_13459,N_12166);
nor U14479 (N_14479,N_13073,N_13176);
or U14480 (N_14480,N_12997,N_12142);
or U14481 (N_14481,N_12169,N_13043);
and U14482 (N_14482,N_13000,N_12178);
and U14483 (N_14483,N_13157,N_12526);
and U14484 (N_14484,N_12191,N_12030);
nand U14485 (N_14485,N_13074,N_12385);
nand U14486 (N_14486,N_12805,N_13269);
nand U14487 (N_14487,N_12416,N_12442);
nor U14488 (N_14488,N_12776,N_12414);
nand U14489 (N_14489,N_13368,N_12459);
or U14490 (N_14490,N_12540,N_12341);
xnor U14491 (N_14491,N_13319,N_12114);
or U14492 (N_14492,N_13459,N_12724);
nor U14493 (N_14493,N_13020,N_12340);
nand U14494 (N_14494,N_13249,N_13077);
nand U14495 (N_14495,N_12018,N_12062);
and U14496 (N_14496,N_13417,N_12502);
nor U14497 (N_14497,N_13129,N_13230);
or U14498 (N_14498,N_13027,N_13320);
nor U14499 (N_14499,N_12570,N_12002);
or U14500 (N_14500,N_12346,N_13496);
xor U14501 (N_14501,N_12420,N_12077);
nand U14502 (N_14502,N_13256,N_12839);
or U14503 (N_14503,N_12802,N_12667);
or U14504 (N_14504,N_12741,N_12008);
or U14505 (N_14505,N_13360,N_12428);
nand U14506 (N_14506,N_12513,N_12508);
nor U14507 (N_14507,N_12312,N_13295);
nor U14508 (N_14508,N_12462,N_12808);
nand U14509 (N_14509,N_12396,N_12984);
nor U14510 (N_14510,N_12705,N_12769);
nand U14511 (N_14511,N_13477,N_13356);
nor U14512 (N_14512,N_12931,N_12401);
nor U14513 (N_14513,N_13224,N_13029);
and U14514 (N_14514,N_12830,N_12045);
nand U14515 (N_14515,N_13278,N_13004);
nor U14516 (N_14516,N_13079,N_12644);
and U14517 (N_14517,N_12668,N_12527);
xnor U14518 (N_14518,N_12951,N_13303);
and U14519 (N_14519,N_13077,N_12173);
nand U14520 (N_14520,N_12466,N_13169);
xor U14521 (N_14521,N_12634,N_12257);
nand U14522 (N_14522,N_13075,N_13392);
or U14523 (N_14523,N_12347,N_13313);
nand U14524 (N_14524,N_13036,N_12764);
or U14525 (N_14525,N_12319,N_13200);
and U14526 (N_14526,N_12660,N_12307);
and U14527 (N_14527,N_13140,N_12811);
and U14528 (N_14528,N_13035,N_12223);
nor U14529 (N_14529,N_12472,N_12572);
or U14530 (N_14530,N_12529,N_12655);
or U14531 (N_14531,N_12667,N_12411);
and U14532 (N_14532,N_13479,N_13395);
or U14533 (N_14533,N_12273,N_13336);
nor U14534 (N_14534,N_12402,N_12520);
nand U14535 (N_14535,N_12857,N_13009);
or U14536 (N_14536,N_13256,N_12432);
and U14537 (N_14537,N_12083,N_13182);
nor U14538 (N_14538,N_12223,N_12335);
nor U14539 (N_14539,N_13255,N_13089);
nor U14540 (N_14540,N_12051,N_12101);
nor U14541 (N_14541,N_13290,N_12130);
or U14542 (N_14542,N_12245,N_13311);
nor U14543 (N_14543,N_13448,N_12636);
nand U14544 (N_14544,N_12004,N_12742);
nand U14545 (N_14545,N_12378,N_12487);
or U14546 (N_14546,N_13436,N_12604);
nor U14547 (N_14547,N_12367,N_12021);
or U14548 (N_14548,N_12524,N_13214);
and U14549 (N_14549,N_12646,N_13039);
or U14550 (N_14550,N_12196,N_12548);
nor U14551 (N_14551,N_12004,N_12739);
nor U14552 (N_14552,N_13346,N_12153);
xor U14553 (N_14553,N_13117,N_13294);
and U14554 (N_14554,N_12108,N_12775);
and U14555 (N_14555,N_13227,N_12404);
nor U14556 (N_14556,N_12075,N_12914);
xor U14557 (N_14557,N_13443,N_12122);
or U14558 (N_14558,N_13238,N_13130);
nand U14559 (N_14559,N_13004,N_12498);
or U14560 (N_14560,N_12136,N_12187);
nand U14561 (N_14561,N_12690,N_12758);
or U14562 (N_14562,N_12051,N_12751);
and U14563 (N_14563,N_13148,N_13073);
or U14564 (N_14564,N_12982,N_12531);
or U14565 (N_14565,N_12906,N_12321);
nand U14566 (N_14566,N_12833,N_13489);
nor U14567 (N_14567,N_13068,N_12608);
nand U14568 (N_14568,N_12156,N_12448);
and U14569 (N_14569,N_12309,N_13310);
nand U14570 (N_14570,N_12394,N_12756);
nor U14571 (N_14571,N_12683,N_12506);
and U14572 (N_14572,N_13323,N_12470);
or U14573 (N_14573,N_12845,N_13149);
and U14574 (N_14574,N_13145,N_12308);
xnor U14575 (N_14575,N_12306,N_13410);
and U14576 (N_14576,N_12208,N_12430);
or U14577 (N_14577,N_12555,N_13284);
xor U14578 (N_14578,N_12753,N_13388);
and U14579 (N_14579,N_12168,N_13112);
nor U14580 (N_14580,N_12569,N_12109);
or U14581 (N_14581,N_13109,N_13457);
or U14582 (N_14582,N_12661,N_12205);
and U14583 (N_14583,N_12610,N_13486);
nor U14584 (N_14584,N_13235,N_12045);
nand U14585 (N_14585,N_12976,N_12235);
xor U14586 (N_14586,N_12297,N_12273);
xnor U14587 (N_14587,N_12771,N_12493);
xnor U14588 (N_14588,N_13332,N_12210);
nand U14589 (N_14589,N_12866,N_13149);
nand U14590 (N_14590,N_12360,N_12747);
nand U14591 (N_14591,N_13134,N_12864);
nor U14592 (N_14592,N_12779,N_13257);
xor U14593 (N_14593,N_13108,N_13158);
nor U14594 (N_14594,N_12345,N_12149);
or U14595 (N_14595,N_13007,N_12158);
and U14596 (N_14596,N_12454,N_13151);
nor U14597 (N_14597,N_12379,N_12955);
nor U14598 (N_14598,N_13388,N_12539);
nand U14599 (N_14599,N_13086,N_13130);
and U14600 (N_14600,N_13374,N_13045);
or U14601 (N_14601,N_12304,N_12046);
nor U14602 (N_14602,N_12072,N_12252);
or U14603 (N_14603,N_12509,N_12951);
xnor U14604 (N_14604,N_12174,N_12924);
nor U14605 (N_14605,N_12137,N_12242);
nand U14606 (N_14606,N_13085,N_12108);
nand U14607 (N_14607,N_13230,N_12308);
or U14608 (N_14608,N_12847,N_12785);
nor U14609 (N_14609,N_12643,N_12896);
xnor U14610 (N_14610,N_12435,N_12510);
and U14611 (N_14611,N_12305,N_13340);
or U14612 (N_14612,N_12656,N_12621);
or U14613 (N_14613,N_13175,N_12609);
and U14614 (N_14614,N_13426,N_12215);
and U14615 (N_14615,N_12321,N_13083);
and U14616 (N_14616,N_12795,N_12835);
nor U14617 (N_14617,N_12598,N_12995);
and U14618 (N_14618,N_13250,N_13290);
nor U14619 (N_14619,N_13409,N_12384);
nand U14620 (N_14620,N_12579,N_12992);
nand U14621 (N_14621,N_12262,N_12805);
nor U14622 (N_14622,N_12855,N_12109);
nand U14623 (N_14623,N_12876,N_12679);
nand U14624 (N_14624,N_12137,N_12850);
or U14625 (N_14625,N_12131,N_12646);
nand U14626 (N_14626,N_12163,N_12645);
nand U14627 (N_14627,N_12628,N_12084);
nand U14628 (N_14628,N_13263,N_12918);
or U14629 (N_14629,N_12201,N_13306);
and U14630 (N_14630,N_12447,N_12090);
nor U14631 (N_14631,N_12239,N_12771);
nand U14632 (N_14632,N_12401,N_12776);
or U14633 (N_14633,N_13161,N_12444);
xnor U14634 (N_14634,N_12525,N_13053);
xor U14635 (N_14635,N_12819,N_12087);
or U14636 (N_14636,N_13158,N_12605);
or U14637 (N_14637,N_13126,N_13041);
and U14638 (N_14638,N_13376,N_13091);
xnor U14639 (N_14639,N_12344,N_12419);
and U14640 (N_14640,N_13217,N_13304);
or U14641 (N_14641,N_12554,N_13034);
and U14642 (N_14642,N_12212,N_12593);
nor U14643 (N_14643,N_12267,N_12849);
xor U14644 (N_14644,N_13251,N_12350);
and U14645 (N_14645,N_13400,N_13467);
nor U14646 (N_14646,N_13149,N_12087);
and U14647 (N_14647,N_12299,N_12852);
and U14648 (N_14648,N_12948,N_13381);
nand U14649 (N_14649,N_12907,N_12295);
nand U14650 (N_14650,N_13015,N_12776);
and U14651 (N_14651,N_12853,N_13008);
and U14652 (N_14652,N_13044,N_12207);
and U14653 (N_14653,N_12497,N_12879);
and U14654 (N_14654,N_12916,N_12601);
or U14655 (N_14655,N_12629,N_12638);
nand U14656 (N_14656,N_12617,N_12838);
and U14657 (N_14657,N_12934,N_12760);
and U14658 (N_14658,N_13026,N_12864);
xnor U14659 (N_14659,N_12035,N_12522);
and U14660 (N_14660,N_13458,N_12712);
or U14661 (N_14661,N_12879,N_13238);
nand U14662 (N_14662,N_12127,N_13468);
xnor U14663 (N_14663,N_12006,N_13182);
nand U14664 (N_14664,N_12012,N_12919);
nor U14665 (N_14665,N_12232,N_12171);
nor U14666 (N_14666,N_12683,N_12292);
or U14667 (N_14667,N_12362,N_12773);
nor U14668 (N_14668,N_13373,N_13431);
and U14669 (N_14669,N_12603,N_13001);
nand U14670 (N_14670,N_12091,N_13096);
xor U14671 (N_14671,N_12312,N_13442);
nor U14672 (N_14672,N_12147,N_13455);
or U14673 (N_14673,N_12337,N_12331);
nor U14674 (N_14674,N_12179,N_12415);
or U14675 (N_14675,N_12840,N_12959);
and U14676 (N_14676,N_12740,N_13240);
and U14677 (N_14677,N_12910,N_12998);
xor U14678 (N_14678,N_12097,N_12005);
xnor U14679 (N_14679,N_13445,N_12077);
and U14680 (N_14680,N_12848,N_12282);
xnor U14681 (N_14681,N_12954,N_13349);
nor U14682 (N_14682,N_13104,N_12125);
nand U14683 (N_14683,N_12588,N_12524);
nand U14684 (N_14684,N_13189,N_12854);
nor U14685 (N_14685,N_12381,N_12951);
nand U14686 (N_14686,N_13438,N_13453);
or U14687 (N_14687,N_12913,N_13345);
nor U14688 (N_14688,N_12942,N_12090);
nand U14689 (N_14689,N_12518,N_13164);
or U14690 (N_14690,N_12392,N_12137);
nand U14691 (N_14691,N_12828,N_12504);
nor U14692 (N_14692,N_12969,N_12187);
xnor U14693 (N_14693,N_12290,N_12408);
nand U14694 (N_14694,N_12816,N_13419);
nor U14695 (N_14695,N_12625,N_12773);
nand U14696 (N_14696,N_13105,N_13399);
xor U14697 (N_14697,N_13290,N_12556);
and U14698 (N_14698,N_12489,N_12764);
nand U14699 (N_14699,N_13023,N_13279);
and U14700 (N_14700,N_13155,N_12976);
nand U14701 (N_14701,N_13236,N_12621);
nor U14702 (N_14702,N_12393,N_12843);
and U14703 (N_14703,N_12162,N_12716);
nor U14704 (N_14704,N_12140,N_12173);
xnor U14705 (N_14705,N_12868,N_13352);
nand U14706 (N_14706,N_13246,N_12649);
xor U14707 (N_14707,N_12945,N_12017);
and U14708 (N_14708,N_12142,N_12394);
nor U14709 (N_14709,N_13022,N_12534);
and U14710 (N_14710,N_12412,N_13096);
nor U14711 (N_14711,N_12064,N_12471);
or U14712 (N_14712,N_12177,N_12729);
or U14713 (N_14713,N_12086,N_12139);
nor U14714 (N_14714,N_13077,N_12676);
and U14715 (N_14715,N_12211,N_13462);
or U14716 (N_14716,N_12631,N_12278);
and U14717 (N_14717,N_13285,N_12117);
nand U14718 (N_14718,N_13452,N_13463);
nor U14719 (N_14719,N_12050,N_12834);
nor U14720 (N_14720,N_12650,N_13094);
and U14721 (N_14721,N_13055,N_12078);
nand U14722 (N_14722,N_12206,N_12337);
nor U14723 (N_14723,N_13180,N_12478);
and U14724 (N_14724,N_12220,N_12167);
nand U14725 (N_14725,N_12088,N_12282);
xor U14726 (N_14726,N_12697,N_13251);
xor U14727 (N_14727,N_12474,N_13397);
or U14728 (N_14728,N_12472,N_12257);
nor U14729 (N_14729,N_12861,N_12934);
nor U14730 (N_14730,N_12558,N_13395);
nor U14731 (N_14731,N_12977,N_12672);
and U14732 (N_14732,N_12090,N_12988);
and U14733 (N_14733,N_13497,N_12628);
and U14734 (N_14734,N_12883,N_12544);
nor U14735 (N_14735,N_13134,N_13301);
nand U14736 (N_14736,N_13119,N_12508);
or U14737 (N_14737,N_13435,N_12768);
nor U14738 (N_14738,N_13481,N_13453);
or U14739 (N_14739,N_12279,N_13013);
nand U14740 (N_14740,N_13208,N_12812);
and U14741 (N_14741,N_13127,N_13103);
and U14742 (N_14742,N_12339,N_13362);
nor U14743 (N_14743,N_12356,N_12293);
or U14744 (N_14744,N_12786,N_13209);
and U14745 (N_14745,N_12321,N_12934);
and U14746 (N_14746,N_12626,N_12402);
nand U14747 (N_14747,N_12098,N_13446);
nor U14748 (N_14748,N_12062,N_13269);
xor U14749 (N_14749,N_12334,N_12306);
nor U14750 (N_14750,N_12869,N_12332);
nor U14751 (N_14751,N_12435,N_13251);
and U14752 (N_14752,N_12792,N_12689);
nor U14753 (N_14753,N_12135,N_13060);
xnor U14754 (N_14754,N_12496,N_12981);
nand U14755 (N_14755,N_13398,N_12466);
and U14756 (N_14756,N_12641,N_12452);
or U14757 (N_14757,N_12326,N_12744);
nand U14758 (N_14758,N_12729,N_13488);
xnor U14759 (N_14759,N_12093,N_12417);
and U14760 (N_14760,N_13076,N_12168);
or U14761 (N_14761,N_12218,N_12641);
and U14762 (N_14762,N_12903,N_13213);
and U14763 (N_14763,N_12170,N_12998);
and U14764 (N_14764,N_12273,N_12928);
nor U14765 (N_14765,N_12437,N_12764);
and U14766 (N_14766,N_13037,N_12475);
and U14767 (N_14767,N_12566,N_12132);
nor U14768 (N_14768,N_13262,N_12775);
nor U14769 (N_14769,N_13042,N_12716);
nor U14770 (N_14770,N_13348,N_12948);
or U14771 (N_14771,N_12830,N_12929);
and U14772 (N_14772,N_12945,N_12818);
or U14773 (N_14773,N_13366,N_12696);
and U14774 (N_14774,N_12084,N_12658);
nand U14775 (N_14775,N_13034,N_12820);
xnor U14776 (N_14776,N_12845,N_13297);
or U14777 (N_14777,N_12138,N_12413);
or U14778 (N_14778,N_13251,N_13400);
nor U14779 (N_14779,N_13211,N_13247);
or U14780 (N_14780,N_12892,N_13277);
nor U14781 (N_14781,N_13348,N_13286);
and U14782 (N_14782,N_12824,N_12711);
or U14783 (N_14783,N_13296,N_13274);
and U14784 (N_14784,N_12572,N_13336);
xnor U14785 (N_14785,N_12655,N_12683);
nor U14786 (N_14786,N_12150,N_12079);
nand U14787 (N_14787,N_12966,N_12812);
xnor U14788 (N_14788,N_12994,N_12284);
and U14789 (N_14789,N_13381,N_13447);
nor U14790 (N_14790,N_13206,N_12087);
xnor U14791 (N_14791,N_13365,N_12854);
or U14792 (N_14792,N_12343,N_13107);
nand U14793 (N_14793,N_13296,N_12254);
nand U14794 (N_14794,N_12748,N_12853);
or U14795 (N_14795,N_13037,N_13073);
nand U14796 (N_14796,N_12067,N_12418);
or U14797 (N_14797,N_13423,N_12508);
nor U14798 (N_14798,N_12432,N_12915);
xnor U14799 (N_14799,N_12815,N_12847);
and U14800 (N_14800,N_12917,N_12653);
or U14801 (N_14801,N_12102,N_13178);
or U14802 (N_14802,N_13401,N_12643);
nor U14803 (N_14803,N_12197,N_13261);
nand U14804 (N_14804,N_13429,N_13132);
and U14805 (N_14805,N_12231,N_12654);
nand U14806 (N_14806,N_12836,N_12527);
nand U14807 (N_14807,N_12479,N_12611);
and U14808 (N_14808,N_12589,N_12988);
or U14809 (N_14809,N_12267,N_12818);
xor U14810 (N_14810,N_12500,N_12213);
xnor U14811 (N_14811,N_12400,N_12805);
xnor U14812 (N_14812,N_12233,N_13479);
or U14813 (N_14813,N_12049,N_13248);
xor U14814 (N_14814,N_13152,N_12526);
and U14815 (N_14815,N_13316,N_13198);
or U14816 (N_14816,N_12707,N_13293);
nand U14817 (N_14817,N_12952,N_12349);
and U14818 (N_14818,N_12192,N_12137);
and U14819 (N_14819,N_12255,N_13191);
nand U14820 (N_14820,N_13497,N_12936);
nand U14821 (N_14821,N_12261,N_12452);
nand U14822 (N_14822,N_13087,N_12439);
nor U14823 (N_14823,N_12539,N_13436);
and U14824 (N_14824,N_12579,N_13186);
or U14825 (N_14825,N_12567,N_12273);
xor U14826 (N_14826,N_12179,N_13266);
or U14827 (N_14827,N_12228,N_12869);
nor U14828 (N_14828,N_12249,N_12985);
or U14829 (N_14829,N_12490,N_12440);
nand U14830 (N_14830,N_12361,N_12984);
and U14831 (N_14831,N_12129,N_12218);
nor U14832 (N_14832,N_13366,N_12181);
nand U14833 (N_14833,N_12896,N_12816);
nor U14834 (N_14834,N_12709,N_12926);
nand U14835 (N_14835,N_12369,N_12344);
nor U14836 (N_14836,N_12982,N_12250);
or U14837 (N_14837,N_12486,N_13272);
or U14838 (N_14838,N_12433,N_13080);
nand U14839 (N_14839,N_13429,N_12989);
and U14840 (N_14840,N_12373,N_13370);
or U14841 (N_14841,N_13027,N_12133);
nand U14842 (N_14842,N_12413,N_12204);
nand U14843 (N_14843,N_13427,N_13217);
nand U14844 (N_14844,N_13466,N_12904);
nor U14845 (N_14845,N_12936,N_12424);
and U14846 (N_14846,N_12217,N_12362);
nand U14847 (N_14847,N_13179,N_12690);
or U14848 (N_14848,N_12203,N_13468);
and U14849 (N_14849,N_13110,N_12151);
or U14850 (N_14850,N_12578,N_12191);
and U14851 (N_14851,N_12921,N_13340);
or U14852 (N_14852,N_12048,N_13471);
or U14853 (N_14853,N_12650,N_12624);
xnor U14854 (N_14854,N_13352,N_12019);
nand U14855 (N_14855,N_12737,N_12652);
nand U14856 (N_14856,N_12183,N_12835);
nand U14857 (N_14857,N_12032,N_13017);
and U14858 (N_14858,N_12381,N_13298);
or U14859 (N_14859,N_13271,N_12546);
and U14860 (N_14860,N_12289,N_13138);
and U14861 (N_14861,N_12672,N_12995);
nor U14862 (N_14862,N_13080,N_12589);
and U14863 (N_14863,N_12608,N_12240);
nand U14864 (N_14864,N_12934,N_12700);
and U14865 (N_14865,N_12757,N_12622);
nor U14866 (N_14866,N_12584,N_13088);
or U14867 (N_14867,N_13021,N_12244);
nand U14868 (N_14868,N_13087,N_13473);
nand U14869 (N_14869,N_13275,N_12171);
or U14870 (N_14870,N_12817,N_13233);
xnor U14871 (N_14871,N_13000,N_12480);
nand U14872 (N_14872,N_13480,N_12612);
and U14873 (N_14873,N_13234,N_13010);
nor U14874 (N_14874,N_12147,N_13236);
and U14875 (N_14875,N_13220,N_12572);
and U14876 (N_14876,N_13460,N_12909);
and U14877 (N_14877,N_12784,N_12876);
xor U14878 (N_14878,N_12862,N_13201);
or U14879 (N_14879,N_12142,N_12786);
or U14880 (N_14880,N_12755,N_13465);
and U14881 (N_14881,N_13076,N_13187);
nand U14882 (N_14882,N_13085,N_12660);
nor U14883 (N_14883,N_13105,N_12001);
nand U14884 (N_14884,N_12262,N_13419);
or U14885 (N_14885,N_12816,N_12284);
or U14886 (N_14886,N_13267,N_12272);
nand U14887 (N_14887,N_13293,N_12356);
and U14888 (N_14888,N_13470,N_13273);
and U14889 (N_14889,N_12111,N_12453);
nand U14890 (N_14890,N_12831,N_12327);
and U14891 (N_14891,N_12939,N_13351);
xnor U14892 (N_14892,N_13293,N_12980);
xnor U14893 (N_14893,N_12604,N_12982);
xnor U14894 (N_14894,N_12974,N_12687);
or U14895 (N_14895,N_13217,N_12811);
or U14896 (N_14896,N_12710,N_12850);
nand U14897 (N_14897,N_12852,N_12881);
or U14898 (N_14898,N_12406,N_12220);
and U14899 (N_14899,N_12043,N_12132);
xnor U14900 (N_14900,N_12334,N_13309);
xnor U14901 (N_14901,N_12836,N_13055);
or U14902 (N_14902,N_13444,N_12327);
nand U14903 (N_14903,N_12636,N_12199);
xor U14904 (N_14904,N_13210,N_13256);
nor U14905 (N_14905,N_13100,N_13296);
nand U14906 (N_14906,N_12734,N_12249);
or U14907 (N_14907,N_12872,N_13190);
xor U14908 (N_14908,N_12724,N_12493);
or U14909 (N_14909,N_12874,N_12932);
and U14910 (N_14910,N_12304,N_12264);
nor U14911 (N_14911,N_12808,N_12703);
nand U14912 (N_14912,N_13436,N_12511);
and U14913 (N_14913,N_12451,N_13353);
or U14914 (N_14914,N_13074,N_13462);
nand U14915 (N_14915,N_12669,N_12649);
and U14916 (N_14916,N_13257,N_13220);
nand U14917 (N_14917,N_13095,N_12873);
nor U14918 (N_14918,N_12091,N_12239);
nand U14919 (N_14919,N_12781,N_12497);
or U14920 (N_14920,N_13259,N_12795);
and U14921 (N_14921,N_13238,N_12340);
nand U14922 (N_14922,N_12290,N_12634);
and U14923 (N_14923,N_12054,N_12004);
or U14924 (N_14924,N_12288,N_12356);
or U14925 (N_14925,N_12271,N_12470);
or U14926 (N_14926,N_12197,N_12409);
or U14927 (N_14927,N_12160,N_12833);
xnor U14928 (N_14928,N_12893,N_13405);
xor U14929 (N_14929,N_12059,N_12243);
and U14930 (N_14930,N_12741,N_12238);
nor U14931 (N_14931,N_12108,N_12919);
nand U14932 (N_14932,N_13320,N_13360);
or U14933 (N_14933,N_12151,N_12531);
or U14934 (N_14934,N_13012,N_13046);
and U14935 (N_14935,N_12865,N_12834);
and U14936 (N_14936,N_12279,N_12792);
and U14937 (N_14937,N_12429,N_12011);
and U14938 (N_14938,N_12219,N_12646);
or U14939 (N_14939,N_12836,N_12815);
xor U14940 (N_14940,N_12244,N_12973);
and U14941 (N_14941,N_12794,N_12128);
nor U14942 (N_14942,N_12673,N_12304);
nand U14943 (N_14943,N_12815,N_13466);
or U14944 (N_14944,N_12901,N_13189);
nand U14945 (N_14945,N_13054,N_12671);
and U14946 (N_14946,N_13100,N_12973);
and U14947 (N_14947,N_12657,N_12009);
nor U14948 (N_14948,N_12348,N_12951);
or U14949 (N_14949,N_12149,N_13345);
xnor U14950 (N_14950,N_12902,N_12782);
nand U14951 (N_14951,N_13486,N_13479);
and U14952 (N_14952,N_12728,N_12202);
or U14953 (N_14953,N_12432,N_12515);
nand U14954 (N_14954,N_12930,N_13076);
nor U14955 (N_14955,N_13228,N_12602);
nor U14956 (N_14956,N_12378,N_13252);
nor U14957 (N_14957,N_13083,N_13219);
nor U14958 (N_14958,N_13245,N_12024);
xnor U14959 (N_14959,N_12009,N_13041);
nor U14960 (N_14960,N_13498,N_12398);
nor U14961 (N_14961,N_13323,N_12785);
and U14962 (N_14962,N_12245,N_12795);
nor U14963 (N_14963,N_12525,N_12811);
xor U14964 (N_14964,N_12369,N_12304);
nor U14965 (N_14965,N_12527,N_13206);
nand U14966 (N_14966,N_13270,N_13317);
nand U14967 (N_14967,N_12742,N_13348);
nand U14968 (N_14968,N_13244,N_12148);
nand U14969 (N_14969,N_12038,N_12805);
nor U14970 (N_14970,N_12763,N_12160);
and U14971 (N_14971,N_12184,N_12788);
xor U14972 (N_14972,N_13289,N_13030);
nand U14973 (N_14973,N_13156,N_13224);
and U14974 (N_14974,N_12073,N_12869);
and U14975 (N_14975,N_12638,N_12341);
nand U14976 (N_14976,N_13054,N_12135);
or U14977 (N_14977,N_12385,N_12414);
and U14978 (N_14978,N_13414,N_12280);
nor U14979 (N_14979,N_12769,N_12067);
nand U14980 (N_14980,N_12870,N_12944);
nand U14981 (N_14981,N_12659,N_12036);
xnor U14982 (N_14982,N_13165,N_12364);
nor U14983 (N_14983,N_13037,N_12591);
xnor U14984 (N_14984,N_12813,N_13139);
or U14985 (N_14985,N_13453,N_12272);
nand U14986 (N_14986,N_12861,N_12879);
nand U14987 (N_14987,N_13265,N_12171);
or U14988 (N_14988,N_12677,N_12745);
or U14989 (N_14989,N_12323,N_13065);
nand U14990 (N_14990,N_13104,N_13432);
nor U14991 (N_14991,N_12130,N_12241);
xnor U14992 (N_14992,N_12188,N_12366);
xnor U14993 (N_14993,N_12188,N_12836);
xor U14994 (N_14994,N_12891,N_12739);
and U14995 (N_14995,N_13109,N_13434);
nor U14996 (N_14996,N_12855,N_13208);
nor U14997 (N_14997,N_12623,N_12978);
nor U14998 (N_14998,N_13044,N_12758);
nor U14999 (N_14999,N_12566,N_12110);
and UO_0 (O_0,N_14867,N_13621);
or UO_1 (O_1,N_14876,N_14277);
nand UO_2 (O_2,N_14213,N_13963);
and UO_3 (O_3,N_14336,N_14424);
nand UO_4 (O_4,N_14159,N_13526);
nand UO_5 (O_5,N_14802,N_14353);
nor UO_6 (O_6,N_14979,N_13893);
nand UO_7 (O_7,N_13620,N_14015);
nor UO_8 (O_8,N_14448,N_13966);
or UO_9 (O_9,N_14124,N_14634);
xnor UO_10 (O_10,N_13528,N_14436);
nand UO_11 (O_11,N_13656,N_13684);
nand UO_12 (O_12,N_14117,N_14589);
and UO_13 (O_13,N_14997,N_13922);
xnor UO_14 (O_14,N_14434,N_13662);
nand UO_15 (O_15,N_13578,N_13548);
or UO_16 (O_16,N_14536,N_14706);
or UO_17 (O_17,N_14507,N_13653);
or UO_18 (O_18,N_13686,N_14269);
and UO_19 (O_19,N_14119,N_13892);
xnor UO_20 (O_20,N_14000,N_13984);
and UO_21 (O_21,N_14279,N_14477);
or UO_22 (O_22,N_13557,N_14446);
nor UO_23 (O_23,N_14447,N_14560);
nor UO_24 (O_24,N_13552,N_13756);
xor UO_25 (O_25,N_14440,N_13775);
nor UO_26 (O_26,N_14325,N_13981);
nor UO_27 (O_27,N_13946,N_14268);
nand UO_28 (O_28,N_14397,N_14454);
or UO_29 (O_29,N_14254,N_13827);
xor UO_30 (O_30,N_13865,N_13742);
xor UO_31 (O_31,N_14501,N_14090);
or UO_32 (O_32,N_14415,N_14452);
or UO_33 (O_33,N_14994,N_14737);
and UO_34 (O_34,N_14999,N_14239);
or UO_35 (O_35,N_13983,N_13729);
and UO_36 (O_36,N_14741,N_14635);
and UO_37 (O_37,N_14420,N_13625);
or UO_38 (O_38,N_14684,N_13670);
nand UO_39 (O_39,N_14464,N_14272);
xor UO_40 (O_40,N_14458,N_13875);
nor UO_41 (O_41,N_14054,N_14895);
nor UO_42 (O_42,N_13673,N_14941);
xnor UO_43 (O_43,N_14045,N_14130);
nand UO_44 (O_44,N_14386,N_14855);
nand UO_45 (O_45,N_14658,N_13795);
and UO_46 (O_46,N_14717,N_14813);
and UO_47 (O_47,N_14746,N_13530);
and UO_48 (O_48,N_13926,N_14870);
and UO_49 (O_49,N_14363,N_14579);
nand UO_50 (O_50,N_13560,N_14647);
nor UO_51 (O_51,N_13772,N_14531);
nor UO_52 (O_52,N_14361,N_13900);
xnor UO_53 (O_53,N_13968,N_14487);
and UO_54 (O_54,N_13898,N_13868);
and UO_55 (O_55,N_13715,N_14222);
xor UO_56 (O_56,N_14591,N_14413);
and UO_57 (O_57,N_14567,N_14396);
xor UO_58 (O_58,N_14598,N_13937);
nand UO_59 (O_59,N_14334,N_14187);
or UO_60 (O_60,N_14766,N_14935);
nor UO_61 (O_61,N_14486,N_13839);
or UO_62 (O_62,N_13899,N_13733);
or UO_63 (O_63,N_13743,N_13592);
and UO_64 (O_64,N_14996,N_13699);
or UO_65 (O_65,N_14449,N_13864);
or UO_66 (O_66,N_13609,N_13734);
nand UO_67 (O_67,N_14557,N_14688);
nand UO_68 (O_68,N_14644,N_14760);
and UO_69 (O_69,N_13681,N_14077);
or UO_70 (O_70,N_14733,N_14586);
and UO_71 (O_71,N_13757,N_13543);
and UO_72 (O_72,N_14341,N_14535);
or UO_73 (O_73,N_13830,N_13654);
nor UO_74 (O_74,N_13655,N_13822);
nand UO_75 (O_75,N_13542,N_13998);
xor UO_76 (O_76,N_14603,N_14835);
or UO_77 (O_77,N_14580,N_14221);
and UO_78 (O_78,N_14463,N_14340);
and UO_79 (O_79,N_13546,N_14692);
or UO_80 (O_80,N_14437,N_14066);
nand UO_81 (O_81,N_14089,N_14711);
nand UO_82 (O_82,N_13515,N_14196);
nor UO_83 (O_83,N_13750,N_13845);
xnor UO_84 (O_84,N_14236,N_14652);
nor UO_85 (O_85,N_13726,N_13944);
nor UO_86 (O_86,N_14701,N_14956);
xnor UO_87 (O_87,N_14663,N_13836);
xnor UO_88 (O_88,N_14190,N_14484);
nand UO_89 (O_89,N_14837,N_14590);
nor UO_90 (O_90,N_14393,N_14808);
nand UO_91 (O_91,N_13501,N_13918);
nor UO_92 (O_92,N_13793,N_14178);
nand UO_93 (O_93,N_14520,N_14332);
xor UO_94 (O_94,N_14314,N_14248);
nand UO_95 (O_95,N_13708,N_14443);
nand UO_96 (O_96,N_14964,N_14351);
nand UO_97 (O_97,N_14127,N_13763);
nor UO_98 (O_98,N_14683,N_13611);
and UO_99 (O_99,N_14005,N_13996);
or UO_100 (O_100,N_14925,N_14331);
nand UO_101 (O_101,N_14110,N_14249);
or UO_102 (O_102,N_14722,N_13646);
or UO_103 (O_103,N_14508,N_13940);
nor UO_104 (O_104,N_13506,N_14076);
or UO_105 (O_105,N_14920,N_13901);
and UO_106 (O_106,N_14262,N_14576);
nand UO_107 (O_107,N_13829,N_14553);
nor UO_108 (O_108,N_13718,N_14461);
or UO_109 (O_109,N_13985,N_14223);
nor UO_110 (O_110,N_14990,N_14662);
nand UO_111 (O_111,N_13999,N_14244);
or UO_112 (O_112,N_14201,N_14329);
xor UO_113 (O_113,N_14150,N_14655);
or UO_114 (O_114,N_14946,N_13623);
and UO_115 (O_115,N_14969,N_13687);
and UO_116 (O_116,N_14164,N_14742);
nand UO_117 (O_117,N_14624,N_14073);
nand UO_118 (O_118,N_14237,N_14842);
nand UO_119 (O_119,N_14206,N_14227);
nor UO_120 (O_120,N_13789,N_14521);
and UO_121 (O_121,N_14273,N_13848);
nor UO_122 (O_122,N_14034,N_14756);
nand UO_123 (O_123,N_14856,N_14305);
nor UO_124 (O_124,N_13693,N_14451);
and UO_125 (O_125,N_14229,N_13907);
or UO_126 (O_126,N_14356,N_14412);
and UO_127 (O_127,N_14904,N_13645);
and UO_128 (O_128,N_13852,N_14417);
or UO_129 (O_129,N_13919,N_14632);
nand UO_130 (O_130,N_14983,N_14065);
and UO_131 (O_131,N_14499,N_14071);
nand UO_132 (O_132,N_14271,N_14901);
nor UO_133 (O_133,N_13558,N_14093);
nand UO_134 (O_134,N_13914,N_13751);
or UO_135 (O_135,N_14184,N_13967);
or UO_136 (O_136,N_13897,N_14167);
or UO_137 (O_137,N_14707,N_14646);
or UO_138 (O_138,N_14369,N_14405);
or UO_139 (O_139,N_13923,N_13711);
or UO_140 (O_140,N_14062,N_14795);
nand UO_141 (O_141,N_14787,N_14051);
xor UO_142 (O_142,N_13881,N_14800);
nor UO_143 (O_143,N_14027,N_13694);
nor UO_144 (O_144,N_14324,N_13814);
and UO_145 (O_145,N_14354,N_13870);
nand UO_146 (O_146,N_14350,N_14182);
nand UO_147 (O_147,N_14654,N_14028);
and UO_148 (O_148,N_14615,N_14659);
nand UO_149 (O_149,N_14980,N_13579);
and UO_150 (O_150,N_14299,N_14940);
nand UO_151 (O_151,N_14714,N_14147);
nand UO_152 (O_152,N_14612,N_14530);
nor UO_153 (O_153,N_14761,N_13706);
and UO_154 (O_154,N_14322,N_14828);
or UO_155 (O_155,N_14165,N_14181);
or UO_156 (O_156,N_13713,N_14109);
and UO_157 (O_157,N_14952,N_13976);
nand UO_158 (O_158,N_13509,N_13631);
or UO_159 (O_159,N_14786,N_14004);
nand UO_160 (O_160,N_14561,N_14665);
and UO_161 (O_161,N_14383,N_14522);
nand UO_162 (O_162,N_14562,N_14200);
nand UO_163 (O_163,N_14376,N_13634);
nor UO_164 (O_164,N_14719,N_14754);
nand UO_165 (O_165,N_13666,N_14650);
or UO_166 (O_166,N_13585,N_14991);
nor UO_167 (O_167,N_13682,N_14774);
nor UO_168 (O_168,N_14911,N_13748);
or UO_169 (O_169,N_14623,N_14748);
or UO_170 (O_170,N_13633,N_13951);
or UO_171 (O_171,N_13770,N_14421);
nand UO_172 (O_172,N_13785,N_13819);
xnor UO_173 (O_173,N_13692,N_13811);
and UO_174 (O_174,N_14040,N_14265);
or UO_175 (O_175,N_13929,N_13920);
and UO_176 (O_176,N_14661,N_13502);
and UO_177 (O_177,N_13791,N_14745);
and UO_178 (O_178,N_13947,N_14868);
or UO_179 (O_179,N_14620,N_14466);
nor UO_180 (O_180,N_14723,N_13735);
nor UO_181 (O_181,N_14605,N_14317);
nand UO_182 (O_182,N_14394,N_14948);
nor UO_183 (O_183,N_14003,N_14203);
and UO_184 (O_184,N_14315,N_14366);
and UO_185 (O_185,N_14116,N_14335);
nand UO_186 (O_186,N_14432,N_13618);
or UO_187 (O_187,N_14479,N_13934);
or UO_188 (O_188,N_14263,N_14713);
nand UO_189 (O_189,N_14462,N_14427);
xnor UO_190 (O_190,N_13752,N_13594);
or UO_191 (O_191,N_14850,N_14505);
nand UO_192 (O_192,N_14129,N_14571);
nor UO_193 (O_193,N_14836,N_14481);
or UO_194 (O_194,N_14512,N_13950);
nand UO_195 (O_195,N_14798,N_13603);
nand UO_196 (O_196,N_14138,N_13941);
and UO_197 (O_197,N_14140,N_13874);
nand UO_198 (O_198,N_13863,N_14465);
or UO_199 (O_199,N_14389,N_13938);
nand UO_200 (O_200,N_14379,N_13608);
and UO_201 (O_201,N_13825,N_14801);
nor UO_202 (O_202,N_14538,N_14725);
or UO_203 (O_203,N_13606,N_14112);
and UO_204 (O_204,N_14215,N_14715);
nand UO_205 (O_205,N_13849,N_14957);
nor UO_206 (O_206,N_13927,N_14482);
nor UO_207 (O_207,N_13664,N_13851);
and UO_208 (O_208,N_14891,N_14298);
nand UO_209 (O_209,N_13943,N_14762);
nor UO_210 (O_210,N_14695,N_14170);
nor UO_211 (O_211,N_14549,N_13590);
and UO_212 (O_212,N_13601,N_14136);
or UO_213 (O_213,N_14998,N_14735);
nor UO_214 (O_214,N_14976,N_13816);
xnor UO_215 (O_215,N_14936,N_14156);
nand UO_216 (O_216,N_14144,N_13761);
or UO_217 (O_217,N_14617,N_13888);
xnor UO_218 (O_218,N_14008,N_13806);
nand UO_219 (O_219,N_14846,N_14653);
or UO_220 (O_220,N_14310,N_14916);
nand UO_221 (O_221,N_14931,N_14540);
xnor UO_222 (O_222,N_14230,N_14260);
nand UO_223 (O_223,N_14671,N_13524);
and UO_224 (O_224,N_14491,N_14799);
nor UO_225 (O_225,N_13774,N_14664);
and UO_226 (O_226,N_14243,N_13913);
nor UO_227 (O_227,N_14960,N_14036);
or UO_228 (O_228,N_14026,N_13615);
and UO_229 (O_229,N_13568,N_13958);
nand UO_230 (O_230,N_14772,N_14416);
nand UO_231 (O_231,N_13828,N_14987);
and UO_232 (O_232,N_14975,N_13826);
nand UO_233 (O_233,N_13702,N_13564);
and UO_234 (O_234,N_13639,N_13841);
xnor UO_235 (O_235,N_14057,N_13513);
nand UO_236 (O_236,N_14785,N_14172);
nor UO_237 (O_237,N_13768,N_14300);
nand UO_238 (O_238,N_14488,N_14552);
nand UO_239 (O_239,N_14729,N_14543);
nand UO_240 (O_240,N_13518,N_14968);
or UO_241 (O_241,N_13628,N_14824);
and UO_242 (O_242,N_14668,N_13799);
nor UO_243 (O_243,N_14608,N_14438);
and UO_244 (O_244,N_14545,N_14890);
nand UO_245 (O_245,N_14199,N_13755);
nand UO_246 (O_246,N_13689,N_13691);
or UO_247 (O_247,N_14294,N_14018);
nor UO_248 (O_248,N_14306,N_14595);
and UO_249 (O_249,N_14510,N_14506);
nor UO_250 (O_250,N_13837,N_14985);
and UO_251 (O_251,N_14803,N_14764);
nor UO_252 (O_252,N_14086,N_14217);
nor UO_253 (O_253,N_13962,N_13847);
or UO_254 (O_254,N_14592,N_14922);
xor UO_255 (O_255,N_14915,N_14607);
nand UO_256 (O_256,N_14233,N_14207);
and UO_257 (O_257,N_14084,N_14641);
nor UO_258 (O_258,N_14905,N_14459);
or UO_259 (O_259,N_14826,N_14024);
nand UO_260 (O_260,N_14881,N_14739);
or UO_261 (O_261,N_13665,N_14872);
xor UO_262 (O_262,N_14435,N_13741);
nand UO_263 (O_263,N_13866,N_14834);
or UO_264 (O_264,N_13760,N_13771);
nand UO_265 (O_265,N_14873,N_13571);
and UO_266 (O_266,N_14053,N_14319);
or UO_267 (O_267,N_13720,N_14814);
nor UO_268 (O_268,N_14455,N_13957);
nor UO_269 (O_269,N_14118,N_14154);
or UO_270 (O_270,N_13555,N_14788);
or UO_271 (O_271,N_14953,N_13857);
and UO_272 (O_272,N_13942,N_14963);
and UO_273 (O_273,N_14977,N_14853);
and UO_274 (O_274,N_13613,N_13889);
and UO_275 (O_275,N_14778,N_13904);
and UO_276 (O_276,N_14686,N_14894);
nand UO_277 (O_277,N_14472,N_14407);
or UO_278 (O_278,N_14295,N_13707);
and UO_279 (O_279,N_13973,N_14770);
and UO_280 (O_280,N_14281,N_14049);
xor UO_281 (O_281,N_14480,N_14186);
nor UO_282 (O_282,N_14564,N_13820);
nand UO_283 (O_283,N_14578,N_14747);
nand UO_284 (O_284,N_14691,N_13562);
nand UO_285 (O_285,N_14330,N_14555);
nand UO_286 (O_286,N_14255,N_14145);
or UO_287 (O_287,N_14710,N_14757);
nand UO_288 (O_288,N_13635,N_14947);
nor UO_289 (O_289,N_14070,N_13593);
or UO_290 (O_290,N_14986,N_14175);
nor UO_291 (O_291,N_13636,N_13978);
nand UO_292 (O_292,N_14485,N_14681);
nand UO_293 (O_293,N_14068,N_13717);
or UO_294 (O_294,N_13710,N_14515);
nand UO_295 (O_295,N_14886,N_14284);
xnor UO_296 (O_296,N_13658,N_13876);
or UO_297 (O_297,N_14541,N_14544);
nor UO_298 (O_298,N_14738,N_14556);
or UO_299 (O_299,N_13727,N_14431);
and UO_300 (O_300,N_14879,N_14301);
nand UO_301 (O_301,N_14374,N_14048);
xnor UO_302 (O_302,N_13887,N_14352);
nor UO_303 (O_303,N_13778,N_14694);
xor UO_304 (O_304,N_13604,N_14736);
or UO_305 (O_305,N_14425,N_13732);
and UO_306 (O_306,N_13986,N_13896);
and UO_307 (O_307,N_13910,N_13780);
and UO_308 (O_308,N_13832,N_14716);
nor UO_309 (O_309,N_14958,N_13796);
nor UO_310 (O_310,N_13858,N_13672);
or UO_311 (O_311,N_14767,N_14102);
nand UO_312 (O_312,N_14075,N_14489);
or UO_313 (O_313,N_13818,N_14318);
xnor UO_314 (O_314,N_14157,N_14442);
or UO_315 (O_315,N_13627,N_14470);
or UO_316 (O_316,N_14573,N_14875);
nand UO_317 (O_317,N_13522,N_13790);
nor UO_318 (O_318,N_13583,N_14583);
nand UO_319 (O_319,N_14385,N_14108);
or UO_320 (O_320,N_14587,N_14669);
xor UO_321 (O_321,N_14871,N_13731);
nand UO_322 (O_322,N_14765,N_14582);
nand UO_323 (O_323,N_13959,N_14860);
nand UO_324 (O_324,N_14844,N_14107);
xor UO_325 (O_325,N_14061,N_14493);
or UO_326 (O_326,N_14794,N_14337);
or UO_327 (O_327,N_13992,N_14132);
or UO_328 (O_328,N_14078,N_14651);
and UO_329 (O_329,N_14818,N_14547);
or UO_330 (O_330,N_14640,N_14899);
xor UO_331 (O_331,N_14577,N_13925);
and UO_332 (O_332,N_14313,N_13703);
or UO_333 (O_333,N_13669,N_13648);
nor UO_334 (O_334,N_13994,N_13644);
or UO_335 (O_335,N_14815,N_14095);
and UO_336 (O_336,N_13667,N_13801);
or UO_337 (O_337,N_14569,N_14457);
nand UO_338 (O_338,N_14893,N_14115);
or UO_339 (O_339,N_14469,N_13700);
nor UO_340 (O_340,N_13948,N_14032);
nor UO_341 (O_341,N_14282,N_14029);
or UO_342 (O_342,N_14606,N_13749);
nand UO_343 (O_343,N_14546,N_13572);
or UO_344 (O_344,N_13800,N_14791);
or UO_345 (O_345,N_13917,N_13643);
and UO_346 (O_346,N_13574,N_14198);
and UO_347 (O_347,N_14627,N_14398);
nand UO_348 (O_348,N_13647,N_14283);
nand UO_349 (O_349,N_14373,N_14810);
and UO_350 (O_350,N_14670,N_14174);
and UO_351 (O_351,N_13619,N_13612);
and UO_352 (O_352,N_14498,N_14266);
xor UO_353 (O_353,N_13758,N_14563);
nor UO_354 (O_354,N_13663,N_13598);
and UO_355 (O_355,N_13817,N_14967);
and UO_356 (O_356,N_14993,N_13565);
and UO_357 (O_357,N_14906,N_14529);
nor UO_358 (O_358,N_13738,N_13709);
and UO_359 (O_359,N_14072,N_14995);
nand UO_360 (O_360,N_14224,N_14637);
nor UO_361 (O_361,N_13529,N_14046);
nor UO_362 (O_362,N_13840,N_14193);
nand UO_363 (O_363,N_14192,N_13792);
and UO_364 (O_364,N_13834,N_14020);
nor UO_365 (O_365,N_14897,N_13971);
nor UO_366 (O_366,N_14047,N_14568);
or UO_367 (O_367,N_14082,N_14289);
nor UO_368 (O_368,N_14690,N_13997);
nor UO_369 (O_369,N_13885,N_14471);
nand UO_370 (O_370,N_13508,N_13591);
nand UO_371 (O_371,N_14101,N_13674);
nand UO_372 (O_372,N_13690,N_14588);
and UO_373 (O_373,N_13545,N_14751);
nand UO_374 (O_374,N_14702,N_14126);
nor UO_375 (O_375,N_13906,N_13519);
xor UO_376 (O_376,N_13764,N_13617);
and UO_377 (O_377,N_14323,N_13652);
nor UO_378 (O_378,N_14418,N_14320);
nand UO_379 (O_379,N_13566,N_14749);
nand UO_380 (O_380,N_14938,N_13746);
or UO_381 (O_381,N_14682,N_14149);
nor UO_382 (O_382,N_14402,N_14992);
nand UO_383 (O_383,N_14974,N_13535);
and UO_384 (O_384,N_14220,N_14400);
and UO_385 (O_385,N_14019,N_14316);
nand UO_386 (O_386,N_13895,N_14513);
and UO_387 (O_387,N_14504,N_14278);
nor UO_388 (O_388,N_13504,N_14423);
nor UO_389 (O_389,N_13928,N_14308);
and UO_390 (O_390,N_14050,N_13668);
nor UO_391 (O_391,N_13714,N_14378);
or UO_392 (O_392,N_13517,N_14291);
nand UO_393 (O_393,N_14104,N_13979);
and UO_394 (O_394,N_14247,N_13831);
or UO_395 (O_395,N_14514,N_14534);
nand UO_396 (O_396,N_14173,N_13777);
and UO_397 (O_397,N_13879,N_13532);
and UO_398 (O_398,N_14518,N_13964);
or UO_399 (O_399,N_14759,N_14209);
and UO_400 (O_400,N_14918,N_14779);
nand UO_401 (O_401,N_13776,N_14091);
nand UO_402 (O_402,N_14044,N_14861);
or UO_403 (O_403,N_13784,N_14932);
nand UO_404 (O_404,N_14011,N_14264);
or UO_405 (O_405,N_14368,N_14554);
and UO_406 (O_406,N_14642,N_13730);
and UO_407 (O_407,N_13544,N_14025);
nand UO_408 (O_408,N_14055,N_14473);
xnor UO_409 (O_409,N_14296,N_14395);
nor UO_410 (O_410,N_14763,N_14384);
nor UO_411 (O_411,N_13838,N_14648);
or UO_412 (O_412,N_14253,N_13823);
or UO_413 (O_413,N_14945,N_14769);
and UO_414 (O_414,N_14923,N_14618);
or UO_415 (O_415,N_14348,N_13728);
xor UO_416 (O_416,N_13576,N_14111);
and UO_417 (O_417,N_13523,N_13626);
xnor UO_418 (O_418,N_14414,N_14478);
or UO_419 (O_419,N_14185,N_14825);
nor UO_420 (O_420,N_14083,N_14371);
or UO_421 (O_421,N_14143,N_14445);
nor UO_422 (O_422,N_13802,N_13953);
nor UO_423 (O_423,N_14246,N_14252);
and UO_424 (O_424,N_14558,N_14240);
and UO_425 (O_425,N_14001,N_14581);
nor UO_426 (O_426,N_13605,N_14476);
or UO_427 (O_427,N_14806,N_14430);
or UO_428 (O_428,N_14060,N_13556);
and UO_429 (O_429,N_14849,N_14900);
nor UO_430 (O_430,N_14841,N_14516);
xnor UO_431 (O_431,N_13807,N_13722);
nand UO_432 (O_432,N_13853,N_14625);
or UO_433 (O_433,N_13961,N_14913);
nand UO_434 (O_434,N_14596,N_14724);
and UO_435 (O_435,N_14845,N_13980);
nand UO_436 (O_436,N_14851,N_14017);
nor UO_437 (O_437,N_14527,N_14257);
nor UO_438 (O_438,N_14226,N_14344);
or UO_439 (O_439,N_14358,N_14619);
nor UO_440 (O_440,N_14775,N_14929);
or UO_441 (O_441,N_14796,N_14892);
nor UO_442 (O_442,N_14467,N_13846);
nor UO_443 (O_443,N_14188,N_14205);
or UO_444 (O_444,N_14888,N_13859);
xnor UO_445 (O_445,N_14303,N_13933);
nor UO_446 (O_446,N_13769,N_14212);
nand UO_447 (O_447,N_14933,N_14832);
nand UO_448 (O_448,N_13582,N_14021);
nand UO_449 (O_449,N_14730,N_14858);
or UO_450 (O_450,N_14633,N_14864);
and UO_451 (O_451,N_14857,N_13642);
nand UO_452 (O_452,N_13527,N_13507);
nor UO_453 (O_453,N_14755,N_14565);
or UO_454 (O_454,N_13581,N_14302);
and UO_455 (O_455,N_14194,N_14866);
or UO_456 (O_456,N_14602,N_14098);
and UO_457 (O_457,N_13854,N_14792);
and UO_458 (O_458,N_14509,N_14307);
or UO_459 (O_459,N_14645,N_13577);
nand UO_460 (O_460,N_14258,N_14820);
nand UO_461 (O_461,N_14539,N_14597);
or UO_462 (O_462,N_14410,N_14697);
and UO_463 (O_463,N_14622,N_14033);
nor UO_464 (O_464,N_14345,N_13659);
or UO_465 (O_465,N_14570,N_13787);
and UO_466 (O_466,N_14016,N_14880);
or UO_467 (O_467,N_13597,N_13931);
nand UO_468 (O_468,N_14636,N_13872);
nor UO_469 (O_469,N_13739,N_13765);
or UO_470 (O_470,N_14146,N_14189);
or UO_471 (O_471,N_14752,N_14649);
nand UO_472 (O_472,N_14208,N_14256);
nor UO_473 (O_473,N_14609,N_13873);
nor UO_474 (O_474,N_13525,N_14532);
and UO_475 (O_475,N_13632,N_13982);
xor UO_476 (O_476,N_14720,N_14013);
nand UO_477 (O_477,N_13930,N_14377);
xnor UO_478 (O_478,N_14962,N_13797);
xnor UO_479 (O_479,N_14698,N_13640);
or UO_480 (O_480,N_14370,N_14153);
nand UO_481 (O_481,N_13835,N_14270);
nand UO_482 (O_482,N_14503,N_14610);
or UO_483 (O_483,N_14492,N_14286);
nor UO_484 (O_484,N_13563,N_14169);
or UO_485 (O_485,N_14882,N_13783);
and UO_486 (O_486,N_14038,N_13924);
and UO_487 (O_487,N_13815,N_14903);
nand UO_488 (O_488,N_14103,N_13745);
nor UO_489 (O_489,N_14495,N_14574);
nand UO_490 (O_490,N_14689,N_13553);
nor UO_491 (O_491,N_13638,N_14099);
nand UO_492 (O_492,N_14460,N_14228);
xnor UO_493 (O_493,N_13610,N_13512);
or UO_494 (O_494,N_13740,N_13891);
nand UO_495 (O_495,N_13736,N_14784);
xor UO_496 (O_496,N_14907,N_14926);
xnor UO_497 (O_497,N_14180,N_14023);
and UO_498 (O_498,N_14183,N_14950);
and UO_499 (O_499,N_14274,N_13683);
or UO_500 (O_500,N_14548,N_14629);
xor UO_501 (O_501,N_14639,N_14843);
xnor UO_502 (O_502,N_14100,N_14972);
nor UO_503 (O_503,N_14081,N_13894);
or UO_504 (O_504,N_13622,N_14357);
nor UO_505 (O_505,N_14128,N_14981);
or UO_506 (O_506,N_14197,N_13676);
nor UO_507 (O_507,N_14304,N_14261);
and UO_508 (O_508,N_14411,N_13936);
nand UO_509 (O_509,N_14638,N_14984);
or UO_510 (O_510,N_13550,N_14456);
nor UO_511 (O_511,N_14359,N_14910);
and UO_512 (O_512,N_14744,N_14106);
nor UO_513 (O_513,N_14327,N_13956);
xor UO_514 (O_514,N_13505,N_13514);
xnor UO_515 (O_515,N_14951,N_14312);
nor UO_516 (O_516,N_14542,N_14789);
or UO_517 (O_517,N_14056,N_14982);
nor UO_518 (O_518,N_14293,N_14811);
nor UO_519 (O_519,N_13878,N_14195);
or UO_520 (O_520,N_14245,N_14219);
xor UO_521 (O_521,N_13599,N_13580);
and UO_522 (O_522,N_14693,N_13698);
nor UO_523 (O_523,N_13551,N_14919);
or UO_524 (O_524,N_14973,N_13890);
xor UO_525 (O_525,N_14666,N_14680);
nor UO_526 (O_526,N_14776,N_14218);
nor UO_527 (O_527,N_13723,N_13861);
xnor UO_528 (O_528,N_13510,N_13701);
or UO_529 (O_529,N_14584,N_14242);
nor UO_530 (O_530,N_13905,N_14444);
nor UO_531 (O_531,N_13909,N_13805);
nor UO_532 (O_532,N_14063,N_14601);
xnor UO_533 (O_533,N_14924,N_14041);
nor UO_534 (O_534,N_14753,N_14902);
nand UO_535 (O_535,N_13503,N_14677);
and UO_536 (O_536,N_14092,N_14380);
and UO_537 (O_537,N_14403,N_13716);
and UO_538 (O_538,N_14210,N_13935);
nand UO_539 (O_539,N_14216,N_13766);
or UO_540 (O_540,N_13880,N_13641);
nor UO_541 (O_541,N_14202,N_14781);
or UO_542 (O_542,N_14777,N_13867);
or UO_543 (O_543,N_13536,N_14022);
and UO_544 (O_544,N_14537,N_13970);
xnor UO_545 (O_545,N_13883,N_14678);
nand UO_546 (O_546,N_13630,N_13675);
and UO_547 (O_547,N_13719,N_14134);
nand UO_548 (O_548,N_13657,N_13697);
nand UO_549 (O_549,N_13549,N_14064);
nor UO_550 (O_550,N_14819,N_13779);
nor UO_551 (O_551,N_14575,N_13902);
or UO_552 (O_552,N_14812,N_14250);
nand UO_553 (O_553,N_14852,N_13573);
nand UO_554 (O_554,N_13680,N_14817);
nand UO_555 (O_555,N_13809,N_13781);
xor UO_556 (O_556,N_13804,N_13843);
and UO_557 (O_557,N_13965,N_14037);
and UO_558 (O_558,N_13559,N_14885);
and UO_559 (O_559,N_14928,N_13725);
or UO_560 (O_560,N_14333,N_14927);
nor UO_561 (O_561,N_14614,N_13767);
and UO_562 (O_562,N_14657,N_14559);
nor UO_563 (O_563,N_14288,N_14042);
xor UO_564 (O_564,N_13788,N_13531);
nor UO_565 (O_565,N_13747,N_13824);
or UO_566 (O_566,N_13537,N_13540);
nand UO_567 (O_567,N_14500,N_14673);
or UO_568 (O_568,N_14404,N_14367);
xnor UO_569 (O_569,N_13637,N_14524);
and UO_570 (O_570,N_14978,N_14816);
nand UO_571 (O_571,N_14321,N_13808);
xnor UO_572 (O_572,N_14593,N_14821);
or UO_573 (O_573,N_14088,N_13915);
nand UO_574 (O_574,N_14162,N_14838);
nand UO_575 (O_575,N_14840,N_13975);
nand UO_576 (O_576,N_13539,N_14827);
and UO_577 (O_577,N_14863,N_13685);
xor UO_578 (O_578,N_14889,N_14631);
nand UO_579 (O_579,N_14703,N_14238);
or UO_580 (O_580,N_14232,N_14059);
or UO_581 (O_581,N_14039,N_13886);
or UO_582 (O_582,N_14912,N_13649);
nand UO_583 (O_583,N_13569,N_13803);
or UO_584 (O_584,N_14704,N_14388);
nand UO_585 (O_585,N_13561,N_14676);
nor UO_586 (O_586,N_14921,N_14783);
xor UO_587 (O_587,N_13547,N_14643);
nor UO_588 (O_588,N_13602,N_14551);
or UO_589 (O_589,N_14087,N_14526);
nand UO_590 (O_590,N_14151,N_14939);
xor UO_591 (O_591,N_13678,N_13520);
or UO_592 (O_592,N_14010,N_14275);
or UO_593 (O_593,N_14667,N_13762);
and UO_594 (O_594,N_14793,N_13952);
nor UO_595 (O_595,N_14177,N_13810);
nor UO_596 (O_596,N_13990,N_14519);
and UO_597 (O_597,N_13833,N_14365);
nand UO_598 (O_598,N_14497,N_13567);
nand UO_599 (O_599,N_14372,N_13737);
nor UO_600 (O_600,N_14490,N_14214);
and UO_601 (O_601,N_14672,N_13993);
or UO_602 (O_602,N_14731,N_14930);
and UO_603 (O_603,N_14166,N_14342);
xnor UO_604 (O_604,N_14347,N_14155);
and UO_605 (O_605,N_14085,N_14750);
or UO_606 (O_606,N_14831,N_13903);
or UO_607 (O_607,N_14626,N_14483);
nand UO_608 (O_608,N_14988,N_14297);
and UO_609 (O_609,N_14934,N_14708);
nor UO_610 (O_610,N_14161,N_14406);
xor UO_611 (O_611,N_14475,N_14758);
or UO_612 (O_612,N_13844,N_13554);
nand UO_613 (O_613,N_13588,N_13908);
nand UO_614 (O_614,N_14728,N_13995);
and UO_615 (O_615,N_13705,N_13589);
and UO_616 (O_616,N_14511,N_14621);
or UO_617 (O_617,N_13533,N_14280);
or UO_618 (O_618,N_14865,N_14171);
and UO_619 (O_619,N_14517,N_14251);
and UO_620 (O_620,N_14080,N_13534);
nor UO_621 (O_621,N_14862,N_14426);
or UO_622 (O_622,N_14734,N_14399);
xor UO_623 (O_623,N_13586,N_14152);
and UO_624 (O_624,N_14031,N_13912);
nor UO_625 (O_625,N_14139,N_13511);
nand UO_626 (O_626,N_13587,N_13538);
or UO_627 (O_627,N_13798,N_14848);
or UO_628 (O_628,N_14113,N_14494);
and UO_629 (O_629,N_14343,N_13989);
or UO_630 (O_630,N_13974,N_14674);
or UO_631 (O_631,N_14869,N_14326);
or UO_632 (O_632,N_13786,N_13945);
xnor UO_633 (O_633,N_14877,N_14768);
nor UO_634 (O_634,N_14699,N_14097);
or UO_635 (O_635,N_14675,N_14830);
nand UO_636 (O_636,N_14392,N_14599);
xor UO_637 (O_637,N_13712,N_13972);
nand UO_638 (O_638,N_14292,N_13860);
nor UO_639 (O_639,N_14959,N_13570);
and UO_640 (O_640,N_14628,N_13724);
nor UO_641 (O_641,N_13575,N_14401);
and UO_642 (O_642,N_13629,N_14285);
and UO_643 (O_643,N_13882,N_14349);
nor UO_644 (O_644,N_14163,N_14450);
and UO_645 (O_645,N_14550,N_14012);
nor UO_646 (O_646,N_14809,N_14566);
and UO_647 (O_647,N_14006,N_14375);
xnor UO_648 (O_648,N_14961,N_13782);
or UO_649 (O_649,N_14009,N_14600);
nor UO_650 (O_650,N_14211,N_14381);
nor UO_651 (O_651,N_14943,N_14179);
xnor UO_652 (O_652,N_14105,N_13856);
and UO_653 (O_653,N_13794,N_14854);
or UO_654 (O_654,N_14259,N_13921);
and UO_655 (O_655,N_14726,N_14533);
or UO_656 (O_656,N_13721,N_14721);
nand UO_657 (O_657,N_13862,N_13869);
and UO_658 (O_658,N_13677,N_14133);
or UO_659 (O_659,N_14884,N_13773);
nor UO_660 (O_660,N_14030,N_14122);
or UO_661 (O_661,N_14771,N_13651);
nand UO_662 (O_662,N_13500,N_14074);
nor UO_663 (O_663,N_14896,N_14656);
nand UO_664 (O_664,N_14409,N_13884);
and UO_665 (O_665,N_14131,N_14362);
or UO_666 (O_666,N_14328,N_13516);
nor UO_667 (O_667,N_13877,N_14712);
xor UO_668 (O_668,N_14727,N_14035);
nor UO_669 (O_669,N_14058,N_14276);
nor UO_670 (O_670,N_14502,N_14887);
or UO_671 (O_671,N_14160,N_14859);
or UO_672 (O_672,N_14267,N_14433);
nor UO_673 (O_673,N_14822,N_13813);
and UO_674 (O_674,N_13704,N_14528);
and UO_675 (O_675,N_13688,N_14740);
nand UO_676 (O_676,N_14382,N_14231);
and UO_677 (O_677,N_14441,N_14338);
nand UO_678 (O_678,N_14829,N_14660);
nand UO_679 (O_679,N_14954,N_13596);
nand UO_680 (O_680,N_13855,N_14613);
and UO_681 (O_681,N_14067,N_14955);
or UO_682 (O_682,N_14096,N_14874);
nor UO_683 (O_683,N_14878,N_14121);
and UO_684 (O_684,N_13595,N_14311);
or UO_685 (O_685,N_14525,N_14287);
and UO_686 (O_686,N_13916,N_14007);
nand UO_687 (O_687,N_14705,N_13696);
nor UO_688 (O_688,N_14696,N_13660);
nand UO_689 (O_689,N_14225,N_14002);
nand UO_690 (O_690,N_14234,N_14782);
or UO_691 (O_691,N_14585,N_13624);
and UO_692 (O_692,N_13614,N_14804);
and UO_693 (O_693,N_14176,N_13871);
and UO_694 (O_694,N_13949,N_14718);
nand UO_695 (O_695,N_14807,N_14474);
nor UO_696 (O_696,N_14141,N_14709);
nor UO_697 (O_697,N_13754,N_14797);
or UO_698 (O_698,N_14355,N_13661);
nor UO_699 (O_699,N_14422,N_14937);
and UO_700 (O_700,N_14429,N_14339);
or UO_701 (O_701,N_13600,N_14158);
nand UO_702 (O_702,N_13679,N_13671);
xor UO_703 (O_703,N_14428,N_13812);
nand UO_704 (O_704,N_14616,N_14914);
nor UO_705 (O_705,N_14790,N_14391);
and UO_706 (O_706,N_14685,N_14043);
xor UO_707 (O_707,N_13759,N_14966);
and UO_708 (O_708,N_14135,N_14079);
nand UO_709 (O_709,N_13988,N_14125);
nor UO_710 (O_710,N_14123,N_14970);
nor UO_711 (O_711,N_14419,N_14360);
nor UO_712 (O_712,N_13987,N_14290);
nand UO_713 (O_713,N_14780,N_14743);
or UO_714 (O_714,N_14908,N_14687);
nand UO_715 (O_715,N_14611,N_14944);
nor UO_716 (O_716,N_13821,N_13695);
or UO_717 (O_717,N_14971,N_14949);
and UO_718 (O_718,N_14094,N_14052);
nor UO_719 (O_719,N_13977,N_14523);
or UO_720 (O_720,N_14839,N_14364);
nor UO_721 (O_721,N_14847,N_14732);
xor UO_722 (O_722,N_13932,N_14439);
nand UO_723 (O_723,N_14468,N_14965);
xor UO_724 (O_724,N_14142,N_13521);
nor UO_725 (O_725,N_14594,N_14917);
or UO_726 (O_726,N_13850,N_13969);
and UO_727 (O_727,N_14309,N_13939);
nand UO_728 (O_728,N_13753,N_13650);
nand UO_729 (O_729,N_14390,N_13842);
nor UO_730 (O_730,N_14604,N_13607);
nand UO_731 (O_731,N_14120,N_14700);
xor UO_732 (O_732,N_14014,N_14241);
nand UO_733 (O_733,N_14630,N_14235);
and UO_734 (O_734,N_14453,N_13954);
nor UO_735 (O_735,N_14805,N_14069);
nand UO_736 (O_736,N_13991,N_14679);
nand UO_737 (O_737,N_14114,N_14496);
and UO_738 (O_738,N_13616,N_14833);
xnor UO_739 (O_739,N_14823,N_14773);
xor UO_740 (O_740,N_14168,N_13960);
and UO_741 (O_741,N_13541,N_13911);
and UO_742 (O_742,N_14898,N_13584);
and UO_743 (O_743,N_14387,N_14883);
and UO_744 (O_744,N_13744,N_14572);
and UO_745 (O_745,N_14191,N_14148);
nor UO_746 (O_746,N_14346,N_14989);
xnor UO_747 (O_747,N_14909,N_14408);
and UO_748 (O_748,N_14942,N_14137);
or UO_749 (O_749,N_13955,N_14204);
nand UO_750 (O_750,N_13517,N_14938);
and UO_751 (O_751,N_14558,N_14641);
nand UO_752 (O_752,N_14013,N_14204);
nor UO_753 (O_753,N_14723,N_14563);
and UO_754 (O_754,N_14841,N_13610);
and UO_755 (O_755,N_14591,N_14374);
and UO_756 (O_756,N_14595,N_13754);
nand UO_757 (O_757,N_14828,N_13847);
nor UO_758 (O_758,N_14122,N_14038);
nor UO_759 (O_759,N_13819,N_13581);
nand UO_760 (O_760,N_13746,N_14475);
or UO_761 (O_761,N_13783,N_14571);
nor UO_762 (O_762,N_13670,N_14836);
nand UO_763 (O_763,N_14399,N_14611);
nand UO_764 (O_764,N_14284,N_14911);
nor UO_765 (O_765,N_14069,N_14515);
nor UO_766 (O_766,N_14782,N_14650);
or UO_767 (O_767,N_14396,N_14268);
nor UO_768 (O_768,N_14215,N_13544);
or UO_769 (O_769,N_14583,N_13726);
xnor UO_770 (O_770,N_14344,N_14933);
nand UO_771 (O_771,N_14454,N_13509);
nor UO_772 (O_772,N_13689,N_14112);
and UO_773 (O_773,N_13767,N_14771);
nand UO_774 (O_774,N_14891,N_14875);
and UO_775 (O_775,N_13725,N_14718);
or UO_776 (O_776,N_14855,N_13511);
or UO_777 (O_777,N_14982,N_14894);
nor UO_778 (O_778,N_14971,N_14403);
nand UO_779 (O_779,N_14255,N_14124);
or UO_780 (O_780,N_14192,N_14110);
and UO_781 (O_781,N_14121,N_13614);
and UO_782 (O_782,N_14242,N_14459);
or UO_783 (O_783,N_14957,N_14377);
nand UO_784 (O_784,N_13503,N_13842);
and UO_785 (O_785,N_13917,N_14791);
nor UO_786 (O_786,N_14156,N_14851);
or UO_787 (O_787,N_14906,N_14153);
nor UO_788 (O_788,N_14438,N_14995);
or UO_789 (O_789,N_14475,N_14295);
xor UO_790 (O_790,N_14689,N_14237);
xnor UO_791 (O_791,N_14774,N_14631);
nand UO_792 (O_792,N_14492,N_14463);
or UO_793 (O_793,N_13989,N_13854);
and UO_794 (O_794,N_13814,N_13955);
nor UO_795 (O_795,N_14666,N_14669);
nor UO_796 (O_796,N_13854,N_14998);
xnor UO_797 (O_797,N_14655,N_14783);
or UO_798 (O_798,N_14477,N_14467);
nand UO_799 (O_799,N_14501,N_13868);
or UO_800 (O_800,N_14958,N_13801);
nor UO_801 (O_801,N_14304,N_13689);
xnor UO_802 (O_802,N_14170,N_14450);
nor UO_803 (O_803,N_14639,N_14201);
and UO_804 (O_804,N_14633,N_14025);
and UO_805 (O_805,N_14796,N_14853);
and UO_806 (O_806,N_14966,N_14397);
nor UO_807 (O_807,N_13826,N_13513);
or UO_808 (O_808,N_14637,N_14307);
and UO_809 (O_809,N_14415,N_13561);
nor UO_810 (O_810,N_14529,N_14966);
nor UO_811 (O_811,N_14460,N_14151);
and UO_812 (O_812,N_13836,N_13526);
or UO_813 (O_813,N_14765,N_14456);
and UO_814 (O_814,N_13740,N_13712);
nor UO_815 (O_815,N_14163,N_13835);
nor UO_816 (O_816,N_14660,N_13871);
and UO_817 (O_817,N_13755,N_13840);
nor UO_818 (O_818,N_14306,N_13665);
and UO_819 (O_819,N_14195,N_14853);
or UO_820 (O_820,N_13668,N_14931);
or UO_821 (O_821,N_14806,N_13554);
nand UO_822 (O_822,N_14738,N_14223);
nand UO_823 (O_823,N_14710,N_14711);
and UO_824 (O_824,N_14958,N_14589);
nand UO_825 (O_825,N_13785,N_13853);
nand UO_826 (O_826,N_14569,N_14761);
nor UO_827 (O_827,N_14127,N_13933);
nor UO_828 (O_828,N_14919,N_14518);
nor UO_829 (O_829,N_14626,N_14450);
xnor UO_830 (O_830,N_14996,N_14444);
and UO_831 (O_831,N_14806,N_14901);
or UO_832 (O_832,N_14648,N_13526);
nand UO_833 (O_833,N_13561,N_14679);
or UO_834 (O_834,N_14666,N_14864);
nand UO_835 (O_835,N_14976,N_13613);
or UO_836 (O_836,N_14572,N_14764);
nor UO_837 (O_837,N_14480,N_13910);
nor UO_838 (O_838,N_13605,N_14553);
nand UO_839 (O_839,N_13611,N_14276);
and UO_840 (O_840,N_13726,N_14423);
or UO_841 (O_841,N_13861,N_13714);
xor UO_842 (O_842,N_13594,N_13505);
and UO_843 (O_843,N_13931,N_13967);
or UO_844 (O_844,N_13848,N_14959);
and UO_845 (O_845,N_13658,N_14029);
and UO_846 (O_846,N_14523,N_14293);
nand UO_847 (O_847,N_13904,N_14394);
or UO_848 (O_848,N_14530,N_14448);
nor UO_849 (O_849,N_14125,N_13560);
or UO_850 (O_850,N_14351,N_14321);
nand UO_851 (O_851,N_13970,N_14108);
or UO_852 (O_852,N_13875,N_14484);
or UO_853 (O_853,N_14449,N_14725);
nor UO_854 (O_854,N_13826,N_14470);
nor UO_855 (O_855,N_14178,N_14536);
nor UO_856 (O_856,N_13629,N_14502);
or UO_857 (O_857,N_14448,N_14381);
and UO_858 (O_858,N_14525,N_14405);
or UO_859 (O_859,N_14430,N_14877);
or UO_860 (O_860,N_14184,N_14763);
nand UO_861 (O_861,N_13903,N_14244);
nand UO_862 (O_862,N_14401,N_14173);
nand UO_863 (O_863,N_13688,N_14881);
nand UO_864 (O_864,N_14264,N_13570);
nand UO_865 (O_865,N_14245,N_14173);
or UO_866 (O_866,N_13526,N_14755);
nor UO_867 (O_867,N_14914,N_13842);
nor UO_868 (O_868,N_14720,N_14180);
and UO_869 (O_869,N_13930,N_14166);
nor UO_870 (O_870,N_14770,N_13786);
or UO_871 (O_871,N_13888,N_14610);
nand UO_872 (O_872,N_14590,N_14353);
nand UO_873 (O_873,N_14905,N_13945);
nor UO_874 (O_874,N_13852,N_13998);
nor UO_875 (O_875,N_14770,N_13916);
or UO_876 (O_876,N_14191,N_14760);
nand UO_877 (O_877,N_14539,N_14236);
and UO_878 (O_878,N_14349,N_14931);
xnor UO_879 (O_879,N_14873,N_13874);
and UO_880 (O_880,N_14753,N_13994);
nand UO_881 (O_881,N_14804,N_14215);
nor UO_882 (O_882,N_13762,N_14696);
and UO_883 (O_883,N_14626,N_13843);
and UO_884 (O_884,N_14341,N_14440);
and UO_885 (O_885,N_14613,N_14299);
nand UO_886 (O_886,N_14283,N_13998);
xnor UO_887 (O_887,N_13992,N_13636);
and UO_888 (O_888,N_14831,N_14280);
xor UO_889 (O_889,N_14799,N_13766);
or UO_890 (O_890,N_13580,N_14427);
or UO_891 (O_891,N_13747,N_14501);
nor UO_892 (O_892,N_14674,N_14966);
or UO_893 (O_893,N_14275,N_13929);
xor UO_894 (O_894,N_14103,N_13596);
nor UO_895 (O_895,N_13535,N_14705);
or UO_896 (O_896,N_14588,N_14093);
and UO_897 (O_897,N_14570,N_14403);
or UO_898 (O_898,N_14438,N_14893);
and UO_899 (O_899,N_13931,N_13875);
nand UO_900 (O_900,N_13681,N_14525);
nand UO_901 (O_901,N_13549,N_13819);
xor UO_902 (O_902,N_13731,N_13935);
or UO_903 (O_903,N_14390,N_14640);
nand UO_904 (O_904,N_14266,N_14742);
xnor UO_905 (O_905,N_13588,N_14441);
or UO_906 (O_906,N_14682,N_14417);
nand UO_907 (O_907,N_14589,N_14606);
nand UO_908 (O_908,N_14062,N_14088);
and UO_909 (O_909,N_13702,N_14658);
or UO_910 (O_910,N_14496,N_13675);
and UO_911 (O_911,N_14773,N_14830);
nor UO_912 (O_912,N_13769,N_13841);
nand UO_913 (O_913,N_14378,N_14805);
and UO_914 (O_914,N_14085,N_14712);
and UO_915 (O_915,N_14027,N_14161);
nand UO_916 (O_916,N_13759,N_14430);
nor UO_917 (O_917,N_14147,N_13570);
nor UO_918 (O_918,N_13521,N_14899);
nor UO_919 (O_919,N_14630,N_14397);
nand UO_920 (O_920,N_13667,N_14756);
nand UO_921 (O_921,N_13809,N_14877);
nor UO_922 (O_922,N_14493,N_14283);
or UO_923 (O_923,N_13598,N_13696);
xor UO_924 (O_924,N_14353,N_14693);
nand UO_925 (O_925,N_13642,N_14095);
and UO_926 (O_926,N_14200,N_14640);
and UO_927 (O_927,N_14711,N_13706);
or UO_928 (O_928,N_13760,N_14274);
and UO_929 (O_929,N_13649,N_14793);
nand UO_930 (O_930,N_14940,N_14221);
nand UO_931 (O_931,N_14098,N_14286);
or UO_932 (O_932,N_14025,N_14671);
nand UO_933 (O_933,N_14032,N_14589);
nand UO_934 (O_934,N_13921,N_14521);
or UO_935 (O_935,N_14947,N_14843);
nand UO_936 (O_936,N_14904,N_14045);
nor UO_937 (O_937,N_14251,N_13867);
nand UO_938 (O_938,N_13602,N_13873);
nor UO_939 (O_939,N_13790,N_14926);
nand UO_940 (O_940,N_13921,N_14287);
or UO_941 (O_941,N_14237,N_13852);
or UO_942 (O_942,N_13869,N_13659);
or UO_943 (O_943,N_14839,N_14687);
or UO_944 (O_944,N_14532,N_14930);
nand UO_945 (O_945,N_14704,N_14916);
and UO_946 (O_946,N_14271,N_14203);
and UO_947 (O_947,N_13686,N_13694);
nor UO_948 (O_948,N_13595,N_13518);
nand UO_949 (O_949,N_14221,N_13601);
and UO_950 (O_950,N_14738,N_14434);
nor UO_951 (O_951,N_14273,N_14782);
or UO_952 (O_952,N_13847,N_14577);
xor UO_953 (O_953,N_13816,N_14914);
or UO_954 (O_954,N_14681,N_14357);
and UO_955 (O_955,N_14881,N_14564);
nand UO_956 (O_956,N_13767,N_14565);
nor UO_957 (O_957,N_14406,N_14019);
xnor UO_958 (O_958,N_14972,N_14440);
and UO_959 (O_959,N_13733,N_14956);
or UO_960 (O_960,N_13847,N_14981);
xor UO_961 (O_961,N_13530,N_14220);
nor UO_962 (O_962,N_13814,N_14110);
nand UO_963 (O_963,N_13500,N_14659);
nand UO_964 (O_964,N_14864,N_14211);
or UO_965 (O_965,N_14848,N_14838);
nand UO_966 (O_966,N_14595,N_13615);
nand UO_967 (O_967,N_14540,N_14587);
xor UO_968 (O_968,N_13656,N_13526);
nand UO_969 (O_969,N_14586,N_14179);
nand UO_970 (O_970,N_13703,N_14117);
and UO_971 (O_971,N_14384,N_13532);
and UO_972 (O_972,N_13766,N_13796);
nand UO_973 (O_973,N_14070,N_14216);
nor UO_974 (O_974,N_14747,N_13949);
and UO_975 (O_975,N_14706,N_13679);
nor UO_976 (O_976,N_14156,N_13683);
nand UO_977 (O_977,N_13662,N_14627);
and UO_978 (O_978,N_14934,N_13935);
nor UO_979 (O_979,N_14574,N_14608);
or UO_980 (O_980,N_14905,N_13722);
nor UO_981 (O_981,N_13930,N_13624);
or UO_982 (O_982,N_14037,N_13709);
nor UO_983 (O_983,N_14000,N_14206);
and UO_984 (O_984,N_14299,N_14044);
and UO_985 (O_985,N_14661,N_14225);
nand UO_986 (O_986,N_14202,N_14708);
nor UO_987 (O_987,N_13755,N_14249);
nor UO_988 (O_988,N_13985,N_14461);
xor UO_989 (O_989,N_13699,N_14665);
nand UO_990 (O_990,N_14329,N_14139);
nor UO_991 (O_991,N_14735,N_13979);
and UO_992 (O_992,N_14408,N_14749);
nand UO_993 (O_993,N_13843,N_14844);
xnor UO_994 (O_994,N_14875,N_13646);
or UO_995 (O_995,N_14518,N_14830);
and UO_996 (O_996,N_13995,N_13713);
and UO_997 (O_997,N_14708,N_14684);
nand UO_998 (O_998,N_14625,N_14028);
and UO_999 (O_999,N_14305,N_14649);
or UO_1000 (O_1000,N_14420,N_13720);
and UO_1001 (O_1001,N_13997,N_14536);
and UO_1002 (O_1002,N_14174,N_13615);
and UO_1003 (O_1003,N_13921,N_13504);
and UO_1004 (O_1004,N_14635,N_13901);
nand UO_1005 (O_1005,N_13719,N_14921);
and UO_1006 (O_1006,N_14074,N_14574);
nand UO_1007 (O_1007,N_14994,N_14705);
and UO_1008 (O_1008,N_14713,N_14832);
xor UO_1009 (O_1009,N_14238,N_14959);
and UO_1010 (O_1010,N_14141,N_14910);
xnor UO_1011 (O_1011,N_14343,N_13919);
nor UO_1012 (O_1012,N_13533,N_13965);
nand UO_1013 (O_1013,N_13506,N_14516);
nor UO_1014 (O_1014,N_14389,N_14196);
nor UO_1015 (O_1015,N_14235,N_13720);
or UO_1016 (O_1016,N_13796,N_14013);
and UO_1017 (O_1017,N_14021,N_14297);
or UO_1018 (O_1018,N_13780,N_14048);
nand UO_1019 (O_1019,N_13794,N_14017);
and UO_1020 (O_1020,N_14021,N_13750);
and UO_1021 (O_1021,N_13894,N_13962);
xnor UO_1022 (O_1022,N_13590,N_13884);
or UO_1023 (O_1023,N_14280,N_14332);
nor UO_1024 (O_1024,N_13746,N_14355);
and UO_1025 (O_1025,N_14631,N_14376);
nand UO_1026 (O_1026,N_14655,N_13988);
or UO_1027 (O_1027,N_14853,N_14443);
nand UO_1028 (O_1028,N_14395,N_14284);
and UO_1029 (O_1029,N_13566,N_13923);
nand UO_1030 (O_1030,N_14814,N_14321);
or UO_1031 (O_1031,N_13809,N_13817);
or UO_1032 (O_1032,N_13877,N_14412);
nand UO_1033 (O_1033,N_14211,N_14618);
nor UO_1034 (O_1034,N_14775,N_13913);
and UO_1035 (O_1035,N_14223,N_14144);
nor UO_1036 (O_1036,N_14730,N_14443);
nand UO_1037 (O_1037,N_14030,N_14256);
and UO_1038 (O_1038,N_13907,N_13745);
nand UO_1039 (O_1039,N_14290,N_14379);
or UO_1040 (O_1040,N_14476,N_14805);
xnor UO_1041 (O_1041,N_14574,N_14768);
or UO_1042 (O_1042,N_14177,N_14028);
or UO_1043 (O_1043,N_13822,N_14521);
or UO_1044 (O_1044,N_14778,N_13771);
nor UO_1045 (O_1045,N_14695,N_13951);
nor UO_1046 (O_1046,N_13776,N_14856);
and UO_1047 (O_1047,N_14901,N_13607);
nor UO_1048 (O_1048,N_14950,N_13534);
or UO_1049 (O_1049,N_14622,N_14062);
xnor UO_1050 (O_1050,N_14689,N_13725);
or UO_1051 (O_1051,N_13697,N_13512);
nor UO_1052 (O_1052,N_14405,N_14392);
nand UO_1053 (O_1053,N_13593,N_13581);
nand UO_1054 (O_1054,N_14154,N_14780);
nor UO_1055 (O_1055,N_14570,N_14178);
or UO_1056 (O_1056,N_14302,N_14621);
and UO_1057 (O_1057,N_14844,N_14700);
xor UO_1058 (O_1058,N_14816,N_13707);
or UO_1059 (O_1059,N_14086,N_14665);
nand UO_1060 (O_1060,N_13660,N_13800);
xor UO_1061 (O_1061,N_14219,N_14354);
and UO_1062 (O_1062,N_14246,N_13886);
nor UO_1063 (O_1063,N_13805,N_14573);
xnor UO_1064 (O_1064,N_13587,N_14779);
xor UO_1065 (O_1065,N_14282,N_14858);
nor UO_1066 (O_1066,N_13639,N_14798);
and UO_1067 (O_1067,N_13930,N_13829);
nor UO_1068 (O_1068,N_14844,N_14522);
and UO_1069 (O_1069,N_14487,N_14249);
nand UO_1070 (O_1070,N_14597,N_14426);
nand UO_1071 (O_1071,N_13943,N_13957);
xnor UO_1072 (O_1072,N_13520,N_14228);
and UO_1073 (O_1073,N_14310,N_14285);
and UO_1074 (O_1074,N_14920,N_13552);
nand UO_1075 (O_1075,N_13868,N_13766);
nand UO_1076 (O_1076,N_14961,N_14670);
or UO_1077 (O_1077,N_14951,N_14266);
nor UO_1078 (O_1078,N_14584,N_14113);
nor UO_1079 (O_1079,N_13936,N_14670);
or UO_1080 (O_1080,N_14694,N_14698);
and UO_1081 (O_1081,N_13953,N_14568);
and UO_1082 (O_1082,N_13567,N_14301);
or UO_1083 (O_1083,N_14120,N_13597);
and UO_1084 (O_1084,N_14342,N_13508);
or UO_1085 (O_1085,N_14001,N_14087);
nor UO_1086 (O_1086,N_14634,N_14089);
or UO_1087 (O_1087,N_13966,N_13587);
and UO_1088 (O_1088,N_14391,N_14981);
nand UO_1089 (O_1089,N_14484,N_13863);
and UO_1090 (O_1090,N_14906,N_14201);
xor UO_1091 (O_1091,N_14047,N_14736);
nand UO_1092 (O_1092,N_13554,N_13907);
and UO_1093 (O_1093,N_13548,N_13519);
nor UO_1094 (O_1094,N_13747,N_13553);
nand UO_1095 (O_1095,N_13756,N_13551);
xnor UO_1096 (O_1096,N_14848,N_14941);
or UO_1097 (O_1097,N_14840,N_14000);
or UO_1098 (O_1098,N_13506,N_14084);
nand UO_1099 (O_1099,N_14940,N_13940);
nor UO_1100 (O_1100,N_13873,N_13516);
or UO_1101 (O_1101,N_14771,N_14629);
xnor UO_1102 (O_1102,N_13911,N_14000);
nand UO_1103 (O_1103,N_14160,N_13630);
nor UO_1104 (O_1104,N_14491,N_13678);
nor UO_1105 (O_1105,N_13616,N_14163);
and UO_1106 (O_1106,N_14726,N_13693);
nor UO_1107 (O_1107,N_13835,N_14870);
xor UO_1108 (O_1108,N_14685,N_14240);
or UO_1109 (O_1109,N_14384,N_14657);
or UO_1110 (O_1110,N_14291,N_13685);
xor UO_1111 (O_1111,N_14729,N_14822);
xnor UO_1112 (O_1112,N_13672,N_14723);
and UO_1113 (O_1113,N_14360,N_14774);
or UO_1114 (O_1114,N_14238,N_14289);
nor UO_1115 (O_1115,N_14333,N_14412);
and UO_1116 (O_1116,N_14803,N_14428);
nand UO_1117 (O_1117,N_14689,N_14597);
xnor UO_1118 (O_1118,N_13831,N_13671);
nand UO_1119 (O_1119,N_14735,N_14425);
nand UO_1120 (O_1120,N_13994,N_13731);
nor UO_1121 (O_1121,N_14023,N_13846);
and UO_1122 (O_1122,N_14800,N_14685);
and UO_1123 (O_1123,N_13934,N_14114);
or UO_1124 (O_1124,N_13923,N_13958);
or UO_1125 (O_1125,N_13881,N_13940);
nor UO_1126 (O_1126,N_13611,N_13553);
xor UO_1127 (O_1127,N_14474,N_14205);
and UO_1128 (O_1128,N_14976,N_14684);
nand UO_1129 (O_1129,N_14310,N_14020);
nor UO_1130 (O_1130,N_14864,N_13967);
nor UO_1131 (O_1131,N_13865,N_13706);
and UO_1132 (O_1132,N_14878,N_13618);
or UO_1133 (O_1133,N_14243,N_13807);
or UO_1134 (O_1134,N_13699,N_14985);
nor UO_1135 (O_1135,N_14558,N_14769);
and UO_1136 (O_1136,N_14096,N_13742);
nor UO_1137 (O_1137,N_13750,N_14658);
and UO_1138 (O_1138,N_14219,N_14429);
nor UO_1139 (O_1139,N_14428,N_13970);
nor UO_1140 (O_1140,N_14103,N_14964);
nor UO_1141 (O_1141,N_14634,N_14408);
nand UO_1142 (O_1142,N_13849,N_14282);
nand UO_1143 (O_1143,N_13653,N_14687);
nand UO_1144 (O_1144,N_14860,N_13991);
and UO_1145 (O_1145,N_14139,N_13677);
nand UO_1146 (O_1146,N_13556,N_14624);
or UO_1147 (O_1147,N_13557,N_13821);
nor UO_1148 (O_1148,N_14638,N_14471);
or UO_1149 (O_1149,N_14648,N_14024);
or UO_1150 (O_1150,N_13955,N_13610);
nand UO_1151 (O_1151,N_14854,N_14138);
nor UO_1152 (O_1152,N_14382,N_13807);
or UO_1153 (O_1153,N_14144,N_14491);
or UO_1154 (O_1154,N_14286,N_13954);
nand UO_1155 (O_1155,N_13612,N_13988);
nor UO_1156 (O_1156,N_14201,N_13754);
nor UO_1157 (O_1157,N_13794,N_14307);
nand UO_1158 (O_1158,N_14592,N_13998);
or UO_1159 (O_1159,N_13837,N_14376);
nor UO_1160 (O_1160,N_14902,N_13966);
and UO_1161 (O_1161,N_14592,N_14128);
nor UO_1162 (O_1162,N_13548,N_14485);
and UO_1163 (O_1163,N_13697,N_14038);
nand UO_1164 (O_1164,N_14614,N_14138);
and UO_1165 (O_1165,N_13583,N_14679);
and UO_1166 (O_1166,N_13984,N_14081);
and UO_1167 (O_1167,N_14257,N_14626);
nand UO_1168 (O_1168,N_14713,N_14022);
and UO_1169 (O_1169,N_13811,N_13780);
xnor UO_1170 (O_1170,N_14951,N_13992);
nor UO_1171 (O_1171,N_13847,N_13824);
or UO_1172 (O_1172,N_14993,N_14614);
nand UO_1173 (O_1173,N_14216,N_14553);
nand UO_1174 (O_1174,N_13796,N_14468);
and UO_1175 (O_1175,N_13750,N_14180);
or UO_1176 (O_1176,N_14543,N_14125);
and UO_1177 (O_1177,N_14754,N_14749);
nand UO_1178 (O_1178,N_14913,N_14587);
nor UO_1179 (O_1179,N_13866,N_14995);
nand UO_1180 (O_1180,N_13974,N_14583);
or UO_1181 (O_1181,N_14187,N_13687);
and UO_1182 (O_1182,N_13972,N_14464);
nand UO_1183 (O_1183,N_13847,N_14952);
nand UO_1184 (O_1184,N_14546,N_13767);
nand UO_1185 (O_1185,N_14949,N_13650);
or UO_1186 (O_1186,N_14129,N_13575);
xnor UO_1187 (O_1187,N_14107,N_13825);
nand UO_1188 (O_1188,N_14109,N_14856);
or UO_1189 (O_1189,N_14655,N_13631);
and UO_1190 (O_1190,N_14398,N_13823);
or UO_1191 (O_1191,N_14819,N_13671);
nor UO_1192 (O_1192,N_13860,N_14972);
and UO_1193 (O_1193,N_13547,N_14064);
and UO_1194 (O_1194,N_13811,N_14191);
nand UO_1195 (O_1195,N_14510,N_14800);
nor UO_1196 (O_1196,N_14842,N_13751);
xor UO_1197 (O_1197,N_14969,N_14106);
and UO_1198 (O_1198,N_14472,N_13650);
nand UO_1199 (O_1199,N_14468,N_14129);
nor UO_1200 (O_1200,N_14825,N_14767);
xor UO_1201 (O_1201,N_14745,N_13614);
and UO_1202 (O_1202,N_13630,N_14007);
or UO_1203 (O_1203,N_14358,N_13559);
nand UO_1204 (O_1204,N_14674,N_13649);
xor UO_1205 (O_1205,N_13947,N_14558);
and UO_1206 (O_1206,N_14347,N_13608);
or UO_1207 (O_1207,N_13598,N_14418);
nor UO_1208 (O_1208,N_14825,N_14053);
nor UO_1209 (O_1209,N_13806,N_14821);
and UO_1210 (O_1210,N_14841,N_13669);
and UO_1211 (O_1211,N_14418,N_14481);
nand UO_1212 (O_1212,N_14302,N_14171);
or UO_1213 (O_1213,N_14264,N_14677);
or UO_1214 (O_1214,N_13943,N_14903);
and UO_1215 (O_1215,N_13633,N_13701);
and UO_1216 (O_1216,N_14395,N_13913);
nand UO_1217 (O_1217,N_14621,N_14822);
nor UO_1218 (O_1218,N_14772,N_14129);
nand UO_1219 (O_1219,N_13994,N_14422);
and UO_1220 (O_1220,N_13665,N_14128);
nand UO_1221 (O_1221,N_13966,N_13683);
nor UO_1222 (O_1222,N_14662,N_13662);
nor UO_1223 (O_1223,N_13516,N_14465);
nand UO_1224 (O_1224,N_13664,N_14859);
or UO_1225 (O_1225,N_13544,N_14730);
nand UO_1226 (O_1226,N_14277,N_14306);
nor UO_1227 (O_1227,N_14704,N_14926);
nor UO_1228 (O_1228,N_13573,N_13922);
nor UO_1229 (O_1229,N_14826,N_14609);
and UO_1230 (O_1230,N_13976,N_14921);
nor UO_1231 (O_1231,N_14332,N_14943);
nand UO_1232 (O_1232,N_14709,N_14580);
nor UO_1233 (O_1233,N_13502,N_13641);
and UO_1234 (O_1234,N_14112,N_14956);
and UO_1235 (O_1235,N_13802,N_13814);
nand UO_1236 (O_1236,N_13535,N_14384);
and UO_1237 (O_1237,N_14006,N_14607);
and UO_1238 (O_1238,N_14474,N_14156);
nand UO_1239 (O_1239,N_14026,N_14205);
nor UO_1240 (O_1240,N_14610,N_13980);
or UO_1241 (O_1241,N_13612,N_14319);
nand UO_1242 (O_1242,N_14676,N_13815);
xnor UO_1243 (O_1243,N_14578,N_14494);
nor UO_1244 (O_1244,N_14673,N_13708);
and UO_1245 (O_1245,N_14845,N_13768);
and UO_1246 (O_1246,N_13880,N_14893);
nand UO_1247 (O_1247,N_13704,N_14331);
or UO_1248 (O_1248,N_13587,N_14685);
or UO_1249 (O_1249,N_14886,N_14343);
xor UO_1250 (O_1250,N_14715,N_14678);
xnor UO_1251 (O_1251,N_14072,N_13768);
or UO_1252 (O_1252,N_14638,N_14160);
nand UO_1253 (O_1253,N_14990,N_14327);
or UO_1254 (O_1254,N_14340,N_14203);
or UO_1255 (O_1255,N_14621,N_14594);
nor UO_1256 (O_1256,N_14802,N_13547);
nor UO_1257 (O_1257,N_13555,N_14998);
nand UO_1258 (O_1258,N_13862,N_14213);
nor UO_1259 (O_1259,N_14634,N_14663);
or UO_1260 (O_1260,N_14711,N_14863);
or UO_1261 (O_1261,N_13656,N_14334);
nand UO_1262 (O_1262,N_14316,N_14783);
nand UO_1263 (O_1263,N_14895,N_13885);
nor UO_1264 (O_1264,N_13517,N_13853);
nor UO_1265 (O_1265,N_14227,N_13981);
nor UO_1266 (O_1266,N_14634,N_13701);
or UO_1267 (O_1267,N_14874,N_14905);
and UO_1268 (O_1268,N_14149,N_14800);
nor UO_1269 (O_1269,N_14569,N_13833);
nand UO_1270 (O_1270,N_14462,N_14160);
and UO_1271 (O_1271,N_13889,N_14773);
nor UO_1272 (O_1272,N_14414,N_14325);
nand UO_1273 (O_1273,N_13999,N_13891);
nor UO_1274 (O_1274,N_14635,N_14336);
nor UO_1275 (O_1275,N_14673,N_14368);
or UO_1276 (O_1276,N_14478,N_13717);
or UO_1277 (O_1277,N_13673,N_14751);
and UO_1278 (O_1278,N_13882,N_14167);
nor UO_1279 (O_1279,N_14516,N_14548);
nand UO_1280 (O_1280,N_13567,N_13980);
or UO_1281 (O_1281,N_14887,N_14769);
xor UO_1282 (O_1282,N_14668,N_14200);
nor UO_1283 (O_1283,N_13990,N_13751);
or UO_1284 (O_1284,N_13930,N_13857);
nand UO_1285 (O_1285,N_13729,N_14086);
nor UO_1286 (O_1286,N_13545,N_14383);
nor UO_1287 (O_1287,N_14423,N_13685);
and UO_1288 (O_1288,N_13790,N_14688);
or UO_1289 (O_1289,N_14620,N_14923);
and UO_1290 (O_1290,N_14544,N_14585);
nor UO_1291 (O_1291,N_14426,N_14666);
nor UO_1292 (O_1292,N_14334,N_14589);
and UO_1293 (O_1293,N_13645,N_14704);
xnor UO_1294 (O_1294,N_14997,N_13871);
and UO_1295 (O_1295,N_14682,N_14619);
or UO_1296 (O_1296,N_14557,N_13813);
xor UO_1297 (O_1297,N_13738,N_13784);
nor UO_1298 (O_1298,N_13820,N_13806);
nor UO_1299 (O_1299,N_14905,N_14675);
nor UO_1300 (O_1300,N_14632,N_14400);
or UO_1301 (O_1301,N_14213,N_14168);
or UO_1302 (O_1302,N_14397,N_14814);
xor UO_1303 (O_1303,N_14786,N_14310);
or UO_1304 (O_1304,N_14106,N_14817);
xnor UO_1305 (O_1305,N_13546,N_13858);
and UO_1306 (O_1306,N_13786,N_14489);
and UO_1307 (O_1307,N_14030,N_13723);
nand UO_1308 (O_1308,N_13907,N_14588);
xor UO_1309 (O_1309,N_14314,N_14006);
xor UO_1310 (O_1310,N_14841,N_14281);
and UO_1311 (O_1311,N_14527,N_14378);
and UO_1312 (O_1312,N_14835,N_13664);
nand UO_1313 (O_1313,N_14750,N_14600);
nor UO_1314 (O_1314,N_13588,N_13975);
and UO_1315 (O_1315,N_14577,N_13598);
nor UO_1316 (O_1316,N_13690,N_13595);
and UO_1317 (O_1317,N_14656,N_14527);
nor UO_1318 (O_1318,N_14299,N_13658);
or UO_1319 (O_1319,N_14166,N_14970);
or UO_1320 (O_1320,N_13777,N_13920);
or UO_1321 (O_1321,N_13657,N_14883);
and UO_1322 (O_1322,N_14647,N_14407);
xnor UO_1323 (O_1323,N_14369,N_14732);
nand UO_1324 (O_1324,N_13702,N_13756);
and UO_1325 (O_1325,N_13508,N_14165);
and UO_1326 (O_1326,N_14650,N_14771);
nand UO_1327 (O_1327,N_13528,N_14164);
and UO_1328 (O_1328,N_14595,N_13785);
nand UO_1329 (O_1329,N_14100,N_14652);
nor UO_1330 (O_1330,N_13974,N_13945);
nor UO_1331 (O_1331,N_14573,N_14374);
xor UO_1332 (O_1332,N_14818,N_14308);
nand UO_1333 (O_1333,N_14285,N_14014);
and UO_1334 (O_1334,N_14735,N_14559);
xor UO_1335 (O_1335,N_14018,N_13675);
nor UO_1336 (O_1336,N_14388,N_14479);
and UO_1337 (O_1337,N_14364,N_13539);
nor UO_1338 (O_1338,N_13936,N_14892);
nand UO_1339 (O_1339,N_14140,N_14149);
nand UO_1340 (O_1340,N_14767,N_14382);
nand UO_1341 (O_1341,N_14064,N_14995);
nand UO_1342 (O_1342,N_14638,N_14559);
nand UO_1343 (O_1343,N_13984,N_13860);
and UO_1344 (O_1344,N_14376,N_14065);
nor UO_1345 (O_1345,N_14902,N_14935);
nor UO_1346 (O_1346,N_14318,N_13912);
nand UO_1347 (O_1347,N_14527,N_14118);
xor UO_1348 (O_1348,N_14623,N_14240);
and UO_1349 (O_1349,N_14679,N_14057);
or UO_1350 (O_1350,N_14932,N_14102);
or UO_1351 (O_1351,N_14181,N_14922);
nor UO_1352 (O_1352,N_14625,N_14744);
nand UO_1353 (O_1353,N_14919,N_14327);
nor UO_1354 (O_1354,N_14753,N_13678);
nand UO_1355 (O_1355,N_14902,N_13578);
or UO_1356 (O_1356,N_14852,N_13621);
nand UO_1357 (O_1357,N_13775,N_14301);
nor UO_1358 (O_1358,N_13843,N_14678);
nand UO_1359 (O_1359,N_14286,N_14320);
and UO_1360 (O_1360,N_14578,N_14988);
or UO_1361 (O_1361,N_14943,N_13966);
nand UO_1362 (O_1362,N_13648,N_13982);
nand UO_1363 (O_1363,N_14353,N_14869);
or UO_1364 (O_1364,N_14441,N_14201);
nand UO_1365 (O_1365,N_14117,N_14878);
nor UO_1366 (O_1366,N_14209,N_13996);
nor UO_1367 (O_1367,N_14418,N_14373);
or UO_1368 (O_1368,N_13778,N_14243);
nand UO_1369 (O_1369,N_14387,N_14203);
nor UO_1370 (O_1370,N_14033,N_14951);
nor UO_1371 (O_1371,N_14528,N_14891);
and UO_1372 (O_1372,N_13631,N_14861);
xor UO_1373 (O_1373,N_14368,N_14214);
nand UO_1374 (O_1374,N_14779,N_13545);
nor UO_1375 (O_1375,N_14618,N_14032);
and UO_1376 (O_1376,N_14534,N_14490);
nor UO_1377 (O_1377,N_14205,N_14371);
or UO_1378 (O_1378,N_13942,N_14341);
nor UO_1379 (O_1379,N_13986,N_14724);
nand UO_1380 (O_1380,N_14423,N_14547);
nand UO_1381 (O_1381,N_14038,N_13945);
nor UO_1382 (O_1382,N_14483,N_14047);
and UO_1383 (O_1383,N_14423,N_13713);
and UO_1384 (O_1384,N_14953,N_14553);
or UO_1385 (O_1385,N_14779,N_13818);
and UO_1386 (O_1386,N_13807,N_14548);
nand UO_1387 (O_1387,N_13522,N_13971);
nand UO_1388 (O_1388,N_14917,N_14023);
nor UO_1389 (O_1389,N_14561,N_14441);
nand UO_1390 (O_1390,N_13901,N_13774);
or UO_1391 (O_1391,N_14127,N_13502);
xnor UO_1392 (O_1392,N_14196,N_14899);
and UO_1393 (O_1393,N_14540,N_14854);
nor UO_1394 (O_1394,N_13666,N_13820);
nor UO_1395 (O_1395,N_14899,N_14110);
or UO_1396 (O_1396,N_13703,N_14475);
nand UO_1397 (O_1397,N_14998,N_14425);
nand UO_1398 (O_1398,N_14501,N_14458);
xor UO_1399 (O_1399,N_13652,N_14278);
nand UO_1400 (O_1400,N_13620,N_14694);
xor UO_1401 (O_1401,N_14486,N_13973);
nand UO_1402 (O_1402,N_14713,N_14141);
nand UO_1403 (O_1403,N_14195,N_14917);
nand UO_1404 (O_1404,N_13542,N_14735);
nor UO_1405 (O_1405,N_14687,N_13963);
xor UO_1406 (O_1406,N_14650,N_14681);
or UO_1407 (O_1407,N_14389,N_14624);
and UO_1408 (O_1408,N_14940,N_14836);
and UO_1409 (O_1409,N_14318,N_14033);
nor UO_1410 (O_1410,N_13830,N_14150);
and UO_1411 (O_1411,N_13631,N_13554);
nand UO_1412 (O_1412,N_14967,N_14558);
or UO_1413 (O_1413,N_14855,N_13527);
nand UO_1414 (O_1414,N_14080,N_14717);
or UO_1415 (O_1415,N_14715,N_14400);
and UO_1416 (O_1416,N_13708,N_14391);
xnor UO_1417 (O_1417,N_14418,N_14704);
nand UO_1418 (O_1418,N_14783,N_14923);
nand UO_1419 (O_1419,N_14321,N_14979);
or UO_1420 (O_1420,N_13735,N_14899);
or UO_1421 (O_1421,N_14422,N_14221);
or UO_1422 (O_1422,N_14465,N_14033);
xor UO_1423 (O_1423,N_13870,N_14339);
and UO_1424 (O_1424,N_14722,N_14783);
or UO_1425 (O_1425,N_13993,N_14438);
and UO_1426 (O_1426,N_14461,N_14131);
or UO_1427 (O_1427,N_14178,N_13841);
or UO_1428 (O_1428,N_14125,N_14371);
nand UO_1429 (O_1429,N_13807,N_14929);
nand UO_1430 (O_1430,N_14321,N_14005);
and UO_1431 (O_1431,N_14648,N_14653);
and UO_1432 (O_1432,N_14450,N_13957);
nand UO_1433 (O_1433,N_13549,N_14327);
nand UO_1434 (O_1434,N_13572,N_14300);
nand UO_1435 (O_1435,N_13721,N_14187);
xnor UO_1436 (O_1436,N_14949,N_13546);
nand UO_1437 (O_1437,N_13946,N_13698);
and UO_1438 (O_1438,N_14819,N_13815);
and UO_1439 (O_1439,N_14567,N_13828);
xor UO_1440 (O_1440,N_14167,N_13852);
nand UO_1441 (O_1441,N_14267,N_13967);
nor UO_1442 (O_1442,N_14701,N_14006);
xor UO_1443 (O_1443,N_14244,N_13507);
nor UO_1444 (O_1444,N_13948,N_14253);
or UO_1445 (O_1445,N_13562,N_14046);
or UO_1446 (O_1446,N_14999,N_13657);
nand UO_1447 (O_1447,N_13710,N_13857);
nor UO_1448 (O_1448,N_14071,N_14730);
nor UO_1449 (O_1449,N_14876,N_14929);
nand UO_1450 (O_1450,N_14346,N_13604);
or UO_1451 (O_1451,N_14893,N_14859);
nand UO_1452 (O_1452,N_13643,N_13563);
xnor UO_1453 (O_1453,N_14063,N_14246);
and UO_1454 (O_1454,N_14230,N_13648);
nand UO_1455 (O_1455,N_14787,N_13580);
nor UO_1456 (O_1456,N_14676,N_14495);
nor UO_1457 (O_1457,N_14939,N_13571);
nand UO_1458 (O_1458,N_14119,N_13722);
nor UO_1459 (O_1459,N_13532,N_13764);
or UO_1460 (O_1460,N_14277,N_13930);
and UO_1461 (O_1461,N_13890,N_14330);
nand UO_1462 (O_1462,N_14728,N_13975);
and UO_1463 (O_1463,N_14144,N_14509);
nor UO_1464 (O_1464,N_14639,N_14313);
and UO_1465 (O_1465,N_14297,N_14504);
nor UO_1466 (O_1466,N_14303,N_13942);
nand UO_1467 (O_1467,N_14079,N_14214);
and UO_1468 (O_1468,N_13860,N_13781);
and UO_1469 (O_1469,N_14695,N_14530);
nand UO_1470 (O_1470,N_14088,N_13681);
nor UO_1471 (O_1471,N_14689,N_14562);
nand UO_1472 (O_1472,N_14325,N_14629);
nor UO_1473 (O_1473,N_13847,N_14701);
nor UO_1474 (O_1474,N_13647,N_14781);
and UO_1475 (O_1475,N_13877,N_13580);
and UO_1476 (O_1476,N_14290,N_13528);
nand UO_1477 (O_1477,N_14955,N_14273);
or UO_1478 (O_1478,N_13969,N_14689);
nand UO_1479 (O_1479,N_13803,N_13712);
and UO_1480 (O_1480,N_14560,N_13830);
or UO_1481 (O_1481,N_14801,N_13999);
nor UO_1482 (O_1482,N_14893,N_13606);
and UO_1483 (O_1483,N_13780,N_14640);
and UO_1484 (O_1484,N_14879,N_14390);
or UO_1485 (O_1485,N_14458,N_14013);
xnor UO_1486 (O_1486,N_14884,N_14313);
nand UO_1487 (O_1487,N_14298,N_14429);
or UO_1488 (O_1488,N_13562,N_14669);
nor UO_1489 (O_1489,N_13558,N_13820);
and UO_1490 (O_1490,N_14517,N_14122);
or UO_1491 (O_1491,N_14543,N_14144);
nor UO_1492 (O_1492,N_14105,N_14168);
nand UO_1493 (O_1493,N_13679,N_13961);
and UO_1494 (O_1494,N_13628,N_14929);
nor UO_1495 (O_1495,N_14213,N_13906);
nor UO_1496 (O_1496,N_14660,N_13730);
nor UO_1497 (O_1497,N_13759,N_13508);
or UO_1498 (O_1498,N_14192,N_14799);
nor UO_1499 (O_1499,N_14713,N_14821);
and UO_1500 (O_1500,N_14733,N_14125);
or UO_1501 (O_1501,N_14630,N_14456);
nand UO_1502 (O_1502,N_14840,N_14451);
nor UO_1503 (O_1503,N_14166,N_13546);
nand UO_1504 (O_1504,N_14517,N_13600);
nor UO_1505 (O_1505,N_14806,N_14407);
or UO_1506 (O_1506,N_13564,N_14660);
nand UO_1507 (O_1507,N_13802,N_13806);
or UO_1508 (O_1508,N_14507,N_13806);
or UO_1509 (O_1509,N_13683,N_14464);
and UO_1510 (O_1510,N_13932,N_14808);
nor UO_1511 (O_1511,N_14697,N_14216);
or UO_1512 (O_1512,N_13544,N_13976);
nor UO_1513 (O_1513,N_14220,N_14227);
nand UO_1514 (O_1514,N_14992,N_14944);
and UO_1515 (O_1515,N_14231,N_13877);
nand UO_1516 (O_1516,N_14013,N_13859);
or UO_1517 (O_1517,N_14641,N_14923);
nor UO_1518 (O_1518,N_14689,N_13985);
xnor UO_1519 (O_1519,N_14516,N_14899);
nand UO_1520 (O_1520,N_14630,N_14035);
or UO_1521 (O_1521,N_14858,N_14447);
nand UO_1522 (O_1522,N_14282,N_13751);
and UO_1523 (O_1523,N_14551,N_14287);
or UO_1524 (O_1524,N_13672,N_14007);
nor UO_1525 (O_1525,N_13542,N_14081);
and UO_1526 (O_1526,N_13835,N_14067);
and UO_1527 (O_1527,N_13610,N_14864);
nor UO_1528 (O_1528,N_14047,N_14805);
nand UO_1529 (O_1529,N_13729,N_13675);
nor UO_1530 (O_1530,N_14743,N_13562);
and UO_1531 (O_1531,N_14259,N_14945);
or UO_1532 (O_1532,N_14839,N_13873);
nor UO_1533 (O_1533,N_14575,N_14363);
and UO_1534 (O_1534,N_14509,N_14985);
nor UO_1535 (O_1535,N_13599,N_14273);
or UO_1536 (O_1536,N_14992,N_14631);
xnor UO_1537 (O_1537,N_14230,N_14277);
nand UO_1538 (O_1538,N_14138,N_14545);
nand UO_1539 (O_1539,N_14009,N_14181);
or UO_1540 (O_1540,N_14575,N_13586);
and UO_1541 (O_1541,N_14483,N_14388);
or UO_1542 (O_1542,N_13817,N_13740);
nand UO_1543 (O_1543,N_13522,N_14608);
and UO_1544 (O_1544,N_14877,N_14594);
nand UO_1545 (O_1545,N_14668,N_14263);
or UO_1546 (O_1546,N_13602,N_14779);
xor UO_1547 (O_1547,N_14290,N_14436);
and UO_1548 (O_1548,N_13512,N_14916);
nand UO_1549 (O_1549,N_14183,N_14317);
nor UO_1550 (O_1550,N_13516,N_13872);
nand UO_1551 (O_1551,N_13717,N_13897);
nand UO_1552 (O_1552,N_13926,N_13802);
and UO_1553 (O_1553,N_14263,N_13957);
nand UO_1554 (O_1554,N_14112,N_14551);
xor UO_1555 (O_1555,N_13642,N_14784);
nand UO_1556 (O_1556,N_14899,N_13691);
or UO_1557 (O_1557,N_14889,N_14651);
nand UO_1558 (O_1558,N_14044,N_13782);
and UO_1559 (O_1559,N_14378,N_14516);
or UO_1560 (O_1560,N_14571,N_14657);
or UO_1561 (O_1561,N_14602,N_14524);
or UO_1562 (O_1562,N_13818,N_14054);
and UO_1563 (O_1563,N_14848,N_14645);
nand UO_1564 (O_1564,N_14996,N_14024);
nand UO_1565 (O_1565,N_13869,N_14189);
and UO_1566 (O_1566,N_14664,N_14430);
nor UO_1567 (O_1567,N_14826,N_14545);
nor UO_1568 (O_1568,N_13650,N_14358);
nor UO_1569 (O_1569,N_13646,N_14281);
nand UO_1570 (O_1570,N_14949,N_14387);
nand UO_1571 (O_1571,N_14837,N_14966);
nor UO_1572 (O_1572,N_13754,N_14587);
xnor UO_1573 (O_1573,N_14678,N_14063);
nand UO_1574 (O_1574,N_14627,N_14182);
nand UO_1575 (O_1575,N_14253,N_14135);
nor UO_1576 (O_1576,N_14310,N_14021);
nand UO_1577 (O_1577,N_14074,N_13944);
nand UO_1578 (O_1578,N_14372,N_14602);
and UO_1579 (O_1579,N_13791,N_14285);
or UO_1580 (O_1580,N_13965,N_13562);
and UO_1581 (O_1581,N_14512,N_14837);
and UO_1582 (O_1582,N_14564,N_14610);
xnor UO_1583 (O_1583,N_14825,N_14923);
or UO_1584 (O_1584,N_13550,N_13786);
and UO_1585 (O_1585,N_14932,N_14402);
or UO_1586 (O_1586,N_13512,N_14283);
nand UO_1587 (O_1587,N_14187,N_14546);
nand UO_1588 (O_1588,N_14251,N_13894);
nand UO_1589 (O_1589,N_14326,N_14430);
and UO_1590 (O_1590,N_14012,N_14353);
or UO_1591 (O_1591,N_13781,N_14694);
nor UO_1592 (O_1592,N_14849,N_13502);
and UO_1593 (O_1593,N_14635,N_14499);
and UO_1594 (O_1594,N_14883,N_13858);
and UO_1595 (O_1595,N_14227,N_13901);
and UO_1596 (O_1596,N_13822,N_13684);
xor UO_1597 (O_1597,N_14075,N_13741);
nor UO_1598 (O_1598,N_14683,N_14907);
and UO_1599 (O_1599,N_14137,N_13548);
nand UO_1600 (O_1600,N_14118,N_14585);
nor UO_1601 (O_1601,N_14218,N_13584);
nand UO_1602 (O_1602,N_14570,N_13756);
xor UO_1603 (O_1603,N_14099,N_14146);
nor UO_1604 (O_1604,N_14885,N_14188);
or UO_1605 (O_1605,N_14288,N_14405);
nand UO_1606 (O_1606,N_14020,N_13624);
and UO_1607 (O_1607,N_14402,N_13631);
nor UO_1608 (O_1608,N_14478,N_13692);
and UO_1609 (O_1609,N_14267,N_14657);
nand UO_1610 (O_1610,N_14029,N_13605);
or UO_1611 (O_1611,N_14505,N_14052);
xnor UO_1612 (O_1612,N_13546,N_14684);
nand UO_1613 (O_1613,N_14675,N_14737);
nand UO_1614 (O_1614,N_14084,N_13835);
nor UO_1615 (O_1615,N_13537,N_14775);
xor UO_1616 (O_1616,N_14830,N_13875);
or UO_1617 (O_1617,N_13984,N_13935);
nand UO_1618 (O_1618,N_13963,N_13804);
nor UO_1619 (O_1619,N_14007,N_13886);
or UO_1620 (O_1620,N_13511,N_14134);
xnor UO_1621 (O_1621,N_14704,N_14858);
and UO_1622 (O_1622,N_14319,N_14264);
nand UO_1623 (O_1623,N_13632,N_13778);
nand UO_1624 (O_1624,N_14998,N_14665);
nor UO_1625 (O_1625,N_14880,N_14733);
and UO_1626 (O_1626,N_14814,N_13568);
nor UO_1627 (O_1627,N_14669,N_14651);
nor UO_1628 (O_1628,N_14428,N_14745);
or UO_1629 (O_1629,N_14108,N_14155);
nor UO_1630 (O_1630,N_14487,N_14296);
or UO_1631 (O_1631,N_13843,N_14672);
nor UO_1632 (O_1632,N_14894,N_13608);
xnor UO_1633 (O_1633,N_14982,N_13992);
nand UO_1634 (O_1634,N_13840,N_14923);
nor UO_1635 (O_1635,N_14067,N_14204);
nand UO_1636 (O_1636,N_14487,N_13573);
or UO_1637 (O_1637,N_14094,N_13954);
nand UO_1638 (O_1638,N_14447,N_14717);
nor UO_1639 (O_1639,N_14981,N_14404);
or UO_1640 (O_1640,N_14586,N_13974);
and UO_1641 (O_1641,N_14885,N_14529);
nand UO_1642 (O_1642,N_14327,N_14545);
nand UO_1643 (O_1643,N_14407,N_13588);
nand UO_1644 (O_1644,N_13740,N_14446);
or UO_1645 (O_1645,N_14389,N_14157);
nor UO_1646 (O_1646,N_13892,N_14120);
xnor UO_1647 (O_1647,N_13861,N_13502);
xor UO_1648 (O_1648,N_14564,N_13790);
or UO_1649 (O_1649,N_14616,N_13801);
xnor UO_1650 (O_1650,N_14502,N_13677);
nand UO_1651 (O_1651,N_14844,N_14225);
xnor UO_1652 (O_1652,N_14192,N_14945);
and UO_1653 (O_1653,N_14887,N_14977);
nand UO_1654 (O_1654,N_14478,N_14127);
xor UO_1655 (O_1655,N_14113,N_13656);
nand UO_1656 (O_1656,N_14560,N_14934);
nor UO_1657 (O_1657,N_14840,N_14787);
or UO_1658 (O_1658,N_13527,N_14309);
or UO_1659 (O_1659,N_14110,N_14146);
and UO_1660 (O_1660,N_14026,N_14624);
nand UO_1661 (O_1661,N_13928,N_14116);
or UO_1662 (O_1662,N_14307,N_14991);
nand UO_1663 (O_1663,N_13962,N_14045);
or UO_1664 (O_1664,N_13970,N_14339);
or UO_1665 (O_1665,N_14094,N_14616);
or UO_1666 (O_1666,N_14370,N_13843);
nor UO_1667 (O_1667,N_14774,N_14814);
or UO_1668 (O_1668,N_13851,N_13918);
or UO_1669 (O_1669,N_13799,N_13614);
or UO_1670 (O_1670,N_13593,N_14354);
xnor UO_1671 (O_1671,N_14935,N_14457);
and UO_1672 (O_1672,N_14190,N_13575);
nand UO_1673 (O_1673,N_14808,N_14507);
and UO_1674 (O_1674,N_14767,N_13818);
or UO_1675 (O_1675,N_14254,N_13994);
or UO_1676 (O_1676,N_13835,N_14374);
or UO_1677 (O_1677,N_14378,N_14293);
and UO_1678 (O_1678,N_14766,N_14608);
nor UO_1679 (O_1679,N_13577,N_13536);
nor UO_1680 (O_1680,N_14469,N_14650);
nor UO_1681 (O_1681,N_14423,N_13834);
nor UO_1682 (O_1682,N_14608,N_14580);
or UO_1683 (O_1683,N_13943,N_14738);
or UO_1684 (O_1684,N_14884,N_14398);
nor UO_1685 (O_1685,N_14154,N_14226);
nand UO_1686 (O_1686,N_14457,N_14602);
or UO_1687 (O_1687,N_13604,N_14686);
or UO_1688 (O_1688,N_14877,N_14040);
nor UO_1689 (O_1689,N_13820,N_13925);
or UO_1690 (O_1690,N_13579,N_13963);
nor UO_1691 (O_1691,N_14206,N_13777);
and UO_1692 (O_1692,N_13781,N_13975);
nand UO_1693 (O_1693,N_14500,N_14815);
or UO_1694 (O_1694,N_14673,N_14185);
xnor UO_1695 (O_1695,N_14858,N_14996);
or UO_1696 (O_1696,N_14442,N_13651);
nand UO_1697 (O_1697,N_13710,N_14707);
or UO_1698 (O_1698,N_13549,N_13930);
nand UO_1699 (O_1699,N_13967,N_14833);
or UO_1700 (O_1700,N_14310,N_14859);
nand UO_1701 (O_1701,N_13729,N_14308);
nand UO_1702 (O_1702,N_14209,N_14520);
xor UO_1703 (O_1703,N_13712,N_14000);
or UO_1704 (O_1704,N_14930,N_13951);
or UO_1705 (O_1705,N_14225,N_14613);
nor UO_1706 (O_1706,N_14756,N_14827);
or UO_1707 (O_1707,N_14486,N_14749);
nand UO_1708 (O_1708,N_13852,N_13615);
nand UO_1709 (O_1709,N_14811,N_13658);
and UO_1710 (O_1710,N_14222,N_14384);
nor UO_1711 (O_1711,N_13771,N_13882);
or UO_1712 (O_1712,N_14694,N_13688);
or UO_1713 (O_1713,N_14782,N_14047);
nand UO_1714 (O_1714,N_13659,N_14413);
and UO_1715 (O_1715,N_14280,N_14972);
nand UO_1716 (O_1716,N_14723,N_14323);
xnor UO_1717 (O_1717,N_13572,N_14842);
nor UO_1718 (O_1718,N_13553,N_14706);
or UO_1719 (O_1719,N_13833,N_14327);
xor UO_1720 (O_1720,N_14376,N_13692);
nand UO_1721 (O_1721,N_14740,N_13521);
and UO_1722 (O_1722,N_14230,N_14215);
or UO_1723 (O_1723,N_14087,N_13558);
or UO_1724 (O_1724,N_13798,N_14953);
or UO_1725 (O_1725,N_13881,N_14016);
nand UO_1726 (O_1726,N_14118,N_13550);
nor UO_1727 (O_1727,N_14919,N_14775);
nand UO_1728 (O_1728,N_14034,N_14349);
nor UO_1729 (O_1729,N_14477,N_13994);
nand UO_1730 (O_1730,N_13897,N_14089);
nor UO_1731 (O_1731,N_14053,N_14709);
and UO_1732 (O_1732,N_13693,N_14835);
and UO_1733 (O_1733,N_14068,N_13670);
nand UO_1734 (O_1734,N_14250,N_13503);
or UO_1735 (O_1735,N_14000,N_14548);
and UO_1736 (O_1736,N_14879,N_13669);
or UO_1737 (O_1737,N_13830,N_13653);
nor UO_1738 (O_1738,N_13603,N_13680);
nand UO_1739 (O_1739,N_13981,N_14342);
nand UO_1740 (O_1740,N_13680,N_14386);
nor UO_1741 (O_1741,N_14424,N_14370);
or UO_1742 (O_1742,N_14370,N_14226);
or UO_1743 (O_1743,N_14687,N_14346);
or UO_1744 (O_1744,N_14780,N_14923);
nor UO_1745 (O_1745,N_13629,N_14554);
or UO_1746 (O_1746,N_14495,N_14587);
and UO_1747 (O_1747,N_14155,N_14121);
nand UO_1748 (O_1748,N_14292,N_14917);
and UO_1749 (O_1749,N_14003,N_14122);
nor UO_1750 (O_1750,N_13547,N_14461);
and UO_1751 (O_1751,N_14880,N_14505);
and UO_1752 (O_1752,N_13500,N_14763);
nor UO_1753 (O_1753,N_13773,N_14583);
nor UO_1754 (O_1754,N_14122,N_13810);
nor UO_1755 (O_1755,N_14366,N_13531);
and UO_1756 (O_1756,N_13604,N_14289);
xor UO_1757 (O_1757,N_14598,N_14001);
or UO_1758 (O_1758,N_14390,N_14125);
nand UO_1759 (O_1759,N_13898,N_14499);
nor UO_1760 (O_1760,N_14580,N_14692);
xor UO_1761 (O_1761,N_14743,N_13793);
xnor UO_1762 (O_1762,N_14919,N_14152);
xnor UO_1763 (O_1763,N_14265,N_13738);
or UO_1764 (O_1764,N_14319,N_14590);
and UO_1765 (O_1765,N_14969,N_13577);
nand UO_1766 (O_1766,N_14222,N_14940);
or UO_1767 (O_1767,N_14833,N_14449);
nand UO_1768 (O_1768,N_14811,N_14006);
nor UO_1769 (O_1769,N_14123,N_14232);
nand UO_1770 (O_1770,N_14248,N_14913);
nor UO_1771 (O_1771,N_14186,N_14960);
nand UO_1772 (O_1772,N_14599,N_14904);
xor UO_1773 (O_1773,N_14993,N_14438);
or UO_1774 (O_1774,N_14020,N_14559);
nor UO_1775 (O_1775,N_14386,N_14999);
nor UO_1776 (O_1776,N_13782,N_14080);
nor UO_1777 (O_1777,N_14353,N_14189);
nor UO_1778 (O_1778,N_14073,N_13607);
nand UO_1779 (O_1779,N_14148,N_13501);
and UO_1780 (O_1780,N_14896,N_13501);
nand UO_1781 (O_1781,N_14242,N_13756);
and UO_1782 (O_1782,N_14276,N_13891);
and UO_1783 (O_1783,N_14569,N_14444);
or UO_1784 (O_1784,N_14283,N_14314);
nor UO_1785 (O_1785,N_14903,N_13756);
nand UO_1786 (O_1786,N_14621,N_13593);
and UO_1787 (O_1787,N_14117,N_14676);
and UO_1788 (O_1788,N_13885,N_14785);
or UO_1789 (O_1789,N_14109,N_14435);
or UO_1790 (O_1790,N_14985,N_14979);
and UO_1791 (O_1791,N_13635,N_14434);
nor UO_1792 (O_1792,N_14204,N_14300);
xor UO_1793 (O_1793,N_13943,N_13586);
xnor UO_1794 (O_1794,N_14535,N_14349);
and UO_1795 (O_1795,N_13576,N_14808);
nand UO_1796 (O_1796,N_14190,N_14373);
nor UO_1797 (O_1797,N_14100,N_14400);
nand UO_1798 (O_1798,N_14273,N_14836);
nor UO_1799 (O_1799,N_13700,N_13831);
nand UO_1800 (O_1800,N_14922,N_14881);
nor UO_1801 (O_1801,N_14713,N_14413);
nor UO_1802 (O_1802,N_13604,N_14409);
nand UO_1803 (O_1803,N_14063,N_14126);
and UO_1804 (O_1804,N_13775,N_14420);
nor UO_1805 (O_1805,N_13968,N_14979);
nor UO_1806 (O_1806,N_14571,N_14636);
and UO_1807 (O_1807,N_14653,N_13606);
and UO_1808 (O_1808,N_14649,N_14646);
nor UO_1809 (O_1809,N_14096,N_14157);
nor UO_1810 (O_1810,N_14484,N_14242);
nor UO_1811 (O_1811,N_13951,N_14666);
nand UO_1812 (O_1812,N_13745,N_14708);
or UO_1813 (O_1813,N_14792,N_14633);
xor UO_1814 (O_1814,N_13772,N_14362);
or UO_1815 (O_1815,N_14413,N_14447);
xor UO_1816 (O_1816,N_13784,N_13624);
nand UO_1817 (O_1817,N_14394,N_14142);
and UO_1818 (O_1818,N_14406,N_13519);
nand UO_1819 (O_1819,N_13900,N_14335);
nand UO_1820 (O_1820,N_14485,N_13629);
or UO_1821 (O_1821,N_13552,N_14938);
nand UO_1822 (O_1822,N_14435,N_14701);
or UO_1823 (O_1823,N_13647,N_14862);
nor UO_1824 (O_1824,N_14007,N_13901);
xnor UO_1825 (O_1825,N_13995,N_13572);
and UO_1826 (O_1826,N_14105,N_14471);
xor UO_1827 (O_1827,N_13545,N_14491);
nor UO_1828 (O_1828,N_14712,N_13887);
nor UO_1829 (O_1829,N_14468,N_14470);
nor UO_1830 (O_1830,N_14994,N_13531);
and UO_1831 (O_1831,N_14848,N_13941);
xor UO_1832 (O_1832,N_14286,N_14161);
or UO_1833 (O_1833,N_14137,N_14916);
nor UO_1834 (O_1834,N_14811,N_13979);
and UO_1835 (O_1835,N_14773,N_14046);
and UO_1836 (O_1836,N_13531,N_14764);
nor UO_1837 (O_1837,N_14366,N_14451);
or UO_1838 (O_1838,N_13949,N_14782);
nand UO_1839 (O_1839,N_14113,N_13704);
or UO_1840 (O_1840,N_13788,N_13703);
and UO_1841 (O_1841,N_14443,N_13772);
nand UO_1842 (O_1842,N_14565,N_14303);
or UO_1843 (O_1843,N_13705,N_13867);
nor UO_1844 (O_1844,N_14129,N_14536);
and UO_1845 (O_1845,N_14985,N_13888);
xor UO_1846 (O_1846,N_13513,N_14092);
nor UO_1847 (O_1847,N_13984,N_14800);
or UO_1848 (O_1848,N_14099,N_14609);
and UO_1849 (O_1849,N_14075,N_14795);
nand UO_1850 (O_1850,N_14443,N_14739);
and UO_1851 (O_1851,N_14734,N_14284);
nand UO_1852 (O_1852,N_14310,N_13848);
nor UO_1853 (O_1853,N_14255,N_14575);
nor UO_1854 (O_1854,N_14485,N_14180);
xor UO_1855 (O_1855,N_14382,N_14698);
nand UO_1856 (O_1856,N_14830,N_14892);
nand UO_1857 (O_1857,N_13813,N_14027);
nand UO_1858 (O_1858,N_13899,N_13848);
and UO_1859 (O_1859,N_13568,N_13803);
and UO_1860 (O_1860,N_14916,N_14566);
nand UO_1861 (O_1861,N_13736,N_14498);
and UO_1862 (O_1862,N_14933,N_14450);
and UO_1863 (O_1863,N_14877,N_13617);
nor UO_1864 (O_1864,N_13967,N_13773);
and UO_1865 (O_1865,N_13824,N_14905);
or UO_1866 (O_1866,N_14406,N_14621);
and UO_1867 (O_1867,N_14271,N_14925);
or UO_1868 (O_1868,N_13823,N_13966);
and UO_1869 (O_1869,N_13779,N_14513);
or UO_1870 (O_1870,N_14691,N_13667);
xnor UO_1871 (O_1871,N_13950,N_13765);
nand UO_1872 (O_1872,N_13774,N_13990);
nor UO_1873 (O_1873,N_14003,N_14991);
nor UO_1874 (O_1874,N_14790,N_14648);
or UO_1875 (O_1875,N_14362,N_13524);
nand UO_1876 (O_1876,N_14103,N_13529);
nand UO_1877 (O_1877,N_14808,N_14420);
or UO_1878 (O_1878,N_14589,N_14053);
nand UO_1879 (O_1879,N_14067,N_14713);
and UO_1880 (O_1880,N_13653,N_13577);
xor UO_1881 (O_1881,N_14001,N_13891);
and UO_1882 (O_1882,N_14268,N_14413);
nand UO_1883 (O_1883,N_14919,N_14143);
xnor UO_1884 (O_1884,N_14044,N_14835);
xor UO_1885 (O_1885,N_14662,N_14015);
xor UO_1886 (O_1886,N_14335,N_13863);
nand UO_1887 (O_1887,N_14646,N_13659);
and UO_1888 (O_1888,N_14738,N_14905);
nor UO_1889 (O_1889,N_14754,N_13987);
and UO_1890 (O_1890,N_13857,N_13703);
and UO_1891 (O_1891,N_13530,N_14502);
or UO_1892 (O_1892,N_14346,N_14216);
xnor UO_1893 (O_1893,N_14803,N_14747);
nand UO_1894 (O_1894,N_14194,N_14030);
xor UO_1895 (O_1895,N_14343,N_13792);
nor UO_1896 (O_1896,N_14996,N_13570);
or UO_1897 (O_1897,N_14770,N_14145);
or UO_1898 (O_1898,N_14752,N_14135);
nor UO_1899 (O_1899,N_14248,N_14627);
or UO_1900 (O_1900,N_13701,N_14571);
nand UO_1901 (O_1901,N_13698,N_13548);
nor UO_1902 (O_1902,N_14679,N_14489);
nand UO_1903 (O_1903,N_13887,N_14983);
nand UO_1904 (O_1904,N_14278,N_14799);
and UO_1905 (O_1905,N_14144,N_14356);
nor UO_1906 (O_1906,N_13594,N_13650);
and UO_1907 (O_1907,N_13697,N_14503);
nand UO_1908 (O_1908,N_13565,N_13714);
and UO_1909 (O_1909,N_13761,N_14211);
nand UO_1910 (O_1910,N_14342,N_13826);
nand UO_1911 (O_1911,N_14963,N_14269);
xor UO_1912 (O_1912,N_14094,N_14231);
and UO_1913 (O_1913,N_14723,N_13865);
or UO_1914 (O_1914,N_13870,N_14483);
or UO_1915 (O_1915,N_14845,N_14085);
or UO_1916 (O_1916,N_13609,N_14079);
or UO_1917 (O_1917,N_13935,N_13605);
or UO_1918 (O_1918,N_14105,N_13903);
or UO_1919 (O_1919,N_13719,N_14663);
nand UO_1920 (O_1920,N_14263,N_14380);
or UO_1921 (O_1921,N_14146,N_13906);
or UO_1922 (O_1922,N_14863,N_14305);
xnor UO_1923 (O_1923,N_14268,N_14968);
or UO_1924 (O_1924,N_14606,N_14658);
nor UO_1925 (O_1925,N_14847,N_14088);
nor UO_1926 (O_1926,N_13978,N_14172);
nor UO_1927 (O_1927,N_14858,N_14272);
nand UO_1928 (O_1928,N_13607,N_14790);
nor UO_1929 (O_1929,N_14869,N_13694);
nand UO_1930 (O_1930,N_14525,N_14008);
nand UO_1931 (O_1931,N_14143,N_14766);
nor UO_1932 (O_1932,N_13617,N_13709);
and UO_1933 (O_1933,N_14998,N_13859);
and UO_1934 (O_1934,N_13543,N_14651);
xor UO_1935 (O_1935,N_13583,N_13544);
nand UO_1936 (O_1936,N_14453,N_13786);
nor UO_1937 (O_1937,N_14998,N_14914);
and UO_1938 (O_1938,N_14258,N_13612);
nor UO_1939 (O_1939,N_14083,N_14568);
and UO_1940 (O_1940,N_14401,N_13692);
xnor UO_1941 (O_1941,N_13958,N_14446);
or UO_1942 (O_1942,N_13649,N_14738);
nand UO_1943 (O_1943,N_14324,N_14874);
nor UO_1944 (O_1944,N_14331,N_14599);
or UO_1945 (O_1945,N_14223,N_14965);
or UO_1946 (O_1946,N_14622,N_13533);
or UO_1947 (O_1947,N_13626,N_14070);
and UO_1948 (O_1948,N_14530,N_14678);
xnor UO_1949 (O_1949,N_14478,N_14081);
nor UO_1950 (O_1950,N_13790,N_13717);
or UO_1951 (O_1951,N_14563,N_14739);
and UO_1952 (O_1952,N_13810,N_14441);
xor UO_1953 (O_1953,N_13512,N_14102);
or UO_1954 (O_1954,N_14981,N_14832);
or UO_1955 (O_1955,N_14620,N_14603);
or UO_1956 (O_1956,N_14743,N_14155);
and UO_1957 (O_1957,N_14529,N_14071);
nor UO_1958 (O_1958,N_14666,N_14479);
and UO_1959 (O_1959,N_13527,N_14919);
and UO_1960 (O_1960,N_13572,N_13725);
nor UO_1961 (O_1961,N_14286,N_13944);
or UO_1962 (O_1962,N_14280,N_13670);
and UO_1963 (O_1963,N_13788,N_14864);
nand UO_1964 (O_1964,N_14295,N_14243);
nand UO_1965 (O_1965,N_14716,N_14310);
or UO_1966 (O_1966,N_13790,N_14712);
nor UO_1967 (O_1967,N_14520,N_13792);
xor UO_1968 (O_1968,N_14289,N_14008);
nand UO_1969 (O_1969,N_14592,N_14790);
nand UO_1970 (O_1970,N_14662,N_13704);
nand UO_1971 (O_1971,N_14890,N_14513);
or UO_1972 (O_1972,N_14517,N_14847);
nor UO_1973 (O_1973,N_14243,N_14450);
nand UO_1974 (O_1974,N_14160,N_14893);
and UO_1975 (O_1975,N_14500,N_13806);
or UO_1976 (O_1976,N_13924,N_13616);
nor UO_1977 (O_1977,N_13730,N_13718);
nand UO_1978 (O_1978,N_13890,N_13673);
nor UO_1979 (O_1979,N_14768,N_13756);
and UO_1980 (O_1980,N_13767,N_13985);
nor UO_1981 (O_1981,N_14726,N_13894);
nor UO_1982 (O_1982,N_14284,N_13660);
nor UO_1983 (O_1983,N_14637,N_14379);
and UO_1984 (O_1984,N_13752,N_14527);
xor UO_1985 (O_1985,N_14162,N_13555);
and UO_1986 (O_1986,N_14837,N_13731);
nor UO_1987 (O_1987,N_14043,N_13728);
and UO_1988 (O_1988,N_13930,N_14243);
or UO_1989 (O_1989,N_13797,N_14922);
or UO_1990 (O_1990,N_13631,N_14210);
nor UO_1991 (O_1991,N_14606,N_14272);
or UO_1992 (O_1992,N_14198,N_14945);
nor UO_1993 (O_1993,N_13984,N_14586);
nor UO_1994 (O_1994,N_14144,N_14324);
nand UO_1995 (O_1995,N_14158,N_13687);
or UO_1996 (O_1996,N_13694,N_13778);
nor UO_1997 (O_1997,N_13719,N_13502);
nor UO_1998 (O_1998,N_14980,N_13648);
and UO_1999 (O_1999,N_14989,N_14356);
endmodule